module VLMultiplier ();

endmodule
