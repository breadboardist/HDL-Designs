
module g16Arbitrator ( \clock.sysClk , \clock.rst , \m00.need , \m00.YouGotIt , 
        \m00.addrM , \m00.DoutM , \m00.DinMast , \m00.Clast_mstr , \s00.Adr , 
        \s00.dbus_in , \s00.dataOut , \s00.tarActive , \s00.Clast , \m01.need , 
        \m01.YouGotIt , \m01.addrM , \m01.DoutM , \m01.DinMast , 
        \m01.Clast_mstr , \s01.Adr , \s01.dbus_in , \s01.dataOut , 
        \s01.tarActive , \s01.Clast , \m02.need , \m02.YouGotIt , \m02.addrM , 
        \m02.DoutM , \m02.DinMast , \m02.Clast_mstr , \s02.Adr , \s02.dbus_in , 
        \s02.dataOut , \s02.tarActive , \s02.Clast , \m03.need , 
        \m03.YouGotIt , \m03.addrM , \m03.DoutM , \m03.DinMast , 
        \m03.Clast_mstr , \s03.Adr , \s03.dbus_in , \s03.dataOut , 
        \s03.tarActive , \s03.Clast , \m04.need , \m04.YouGotIt , \m04.addrM , 
        \m04.DoutM , \m04.DinMast , \m04.Clast_mstr , \s04.Adr , \s04.dbus_in , 
        \s04.dataOut , \s04.tarActive , \s04.Clast , \m05.need , 
        \m05.YouGotIt , \m05.addrM , \m05.DoutM , \m05.DinMast , 
        \m05.Clast_mstr , \s05.Adr , \s05.dbus_in , \s05.dataOut , 
        \s05.tarActive , \s05.Clast , \m06.need , \m06.YouGotIt , \m06.addrM , 
        \m06.DoutM , \m06.DinMast , \m06.Clast_mstr , \s06.Adr , \s06.dbus_in , 
        \s06.dataOut , \s06.tarActive , \s06.Clast , \s07.Adr , \s07.dbus_in , 
        \s07.dataOut , \s07.tarActive , \s07.Clast , \s08.Adr , \s08.dbus_in , 
        \s08.dataOut , \s08.tarActive , \s08.Clast , \s09.Adr , \s09.dbus_in , 
        \s09.dataOut , \s09.tarActive , \s09.Clast , \s10.Adr , \s10.dbus_in , 
        \s10.dataOut , \s10.tarActive , \s10.Clast , \s11.Adr , \s11.dbus_in , 
        \s11.dataOut , \s11.tarActive , \s11.Clast , \s12.Adr , \s12.dbus_in , 
        \s12.dataOut , \s12.tarActive , \s12.Clast , \s13.Adr , \s13.dbus_in , 
        \s13.dataOut , \s13.tarActive , \s13.Clast  );
  input [47:0] \m00.addrM ;
  input [15:0] \m00.DoutM ;
  output [15:0] \m00.DinMast ;
  output [47:0] \s00.Adr ;
  output [15:0] \s00.dbus_in ;
  input [15:0] \s00.dataOut ;
  input [47:0] \m01.addrM ;
  input [15:0] \m01.DoutM ;
  output [15:0] \m01.DinMast ;
  output [47:0] \s01.Adr ;
  output [15:0] \s01.dbus_in ;
  input [15:0] \s01.dataOut ;
  input [47:0] \m02.addrM ;
  input [15:0] \m02.DoutM ;
  output [15:0] \m02.DinMast ;
  output [47:0] \s02.Adr ;
  output [15:0] \s02.dbus_in ;
  input [15:0] \s02.dataOut ;
  input [47:0] \m03.addrM ;
  input [15:0] \m03.DoutM ;
  output [15:0] \m03.DinMast ;
  output [47:0] \s03.Adr ;
  output [15:0] \s03.dbus_in ;
  input [15:0] \s03.dataOut ;
  input [47:0] \m04.addrM ;
  input [15:0] \m04.DoutM ;
  output [15:0] \m04.DinMast ;
  output [47:0] \s04.Adr ;
  output [15:0] \s04.dbus_in ;
  input [15:0] \s04.dataOut ;
  input [47:0] \m05.addrM ;
  input [15:0] \m05.DoutM ;
  output [15:0] \m05.DinMast ;
  output [47:0] \s05.Adr ;
  output [15:0] \s05.dbus_in ;
  input [15:0] \s05.dataOut ;
  input [47:0] \m06.addrM ;
  input [15:0] \m06.DoutM ;
  output [15:0] \m06.DinMast ;
  output [47:0] \s06.Adr ;
  output [15:0] \s06.dbus_in ;
  input [15:0] \s06.dataOut ;
  output [47:0] \s07.Adr ;
  output [15:0] \s07.dbus_in ;
  input [15:0] \s07.dataOut ;
  output [47:0] \s08.Adr ;
  output [15:0] \s08.dbus_in ;
  input [15:0] \s08.dataOut ;
  output [47:0] \s09.Adr ;
  output [15:0] \s09.dbus_in ;
  input [15:0] \s09.dataOut ;
  output [47:0] \s10.Adr ;
  output [15:0] \s10.dbus_in ;
  input [15:0] \s10.dataOut ;
  output [47:0] \s11.Adr ;
  output [15:0] \s11.dbus_in ;
  input [15:0] \s11.dataOut ;
  output [47:0] \s12.Adr ;
  output [15:0] \s12.dbus_in ;
  input [15:0] \s12.dataOut ;
  output [47:0] \s13.Adr ;
  output [15:0] \s13.dbus_in ;
  input [15:0] \s13.dataOut ;
  input \clock.sysClk , \clock.rst , \m00.need , \m01.need , \m02.need ,
         \m03.need , \m04.need , \m05.need , \m06.need ;
  output \m00.YouGotIt , \m00.Clast_mstr , \s00.tarActive , \s00.Clast ,
         \m01.YouGotIt , \m01.Clast_mstr , \s01.tarActive , \s01.Clast ,
         \m02.YouGotIt , \m02.Clast_mstr , \s02.tarActive , \s02.Clast ,
         \m03.YouGotIt , \m03.Clast_mstr , \s03.tarActive , \s03.Clast ,
         \m04.YouGotIt , \m04.Clast_mstr , \s04.tarActive , \s04.Clast ,
         \m05.YouGotIt , \m05.Clast_mstr , \s05.tarActive , \s05.Clast ,
         \m06.YouGotIt , \m06.Clast_mstr , \s06.tarActive , \s06.Clast ,
         \s07.tarActive , \s07.Clast , \s08.tarActive , \s08.Clast ,
         \s09.tarActive , \s09.Clast , \s10.tarActive , \s10.Clast ,
         \s11.tarActive , \s11.Clast , \s12.tarActive , \s12.Clast ,
         \s13.tarActive , \s13.Clast ;
  wire   n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5224,
         n5225, n5235, n5245, n5255, n5265, n5275, n5285, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746;
  assign \s00.Adr  [47] = 1'b0;
  assign \s00.Adr  [46] = 1'b0;
  assign \s00.Adr  [45] = 1'b0;
  assign \s00.Adr  [44] = 1'b0;
  assign \s00.Adr  [43] = 1'b0;
  assign \s00.Adr  [42] = 1'b0;
  assign \s00.Adr  [41] = 1'b0;
  assign \s00.Adr  [40] = 1'b0;
  assign \s00.Adr  [39] = 1'b0;
  assign \s00.Adr  [38] = 1'b0;
  assign \s00.Adr  [37] = 1'b0;
  assign \s00.Adr  [36] = 1'b0;
  assign \s00.Adr  [35] = 1'b0;
  assign \s00.Adr  [34] = 1'b0;
  assign \s00.Adr  [33] = 1'b0;
  assign \s00.Adr  [32] = 1'b0;
  assign \s00.Adr  [31] = 1'b0;
  assign \s00.Adr  [30] = 1'b0;
  assign \s00.Adr  [29] = 1'b0;
  assign \s00.Adr  [28] = 1'b0;
  assign \s00.Adr  [27] = 1'b0;
  assign \s00.Adr  [26] = 1'b0;
  assign \s00.Adr  [25] = 1'b0;
  assign \s00.Adr  [24] = 1'b0;
  assign \s00.Adr  [23] = 1'b1;
  assign \s00.Adr  [22] = 1'b1;
  assign \s00.Adr  [21] = 1'b1;
  assign \s00.Adr  [20] = 1'b1;
  assign \s00.Adr  [19] = 1'b1;
  assign \s00.Adr  [18] = 1'b1;
  assign \s00.Adr  [17] = 1'b1;
  assign \s00.Adr  [16] = 1'b1;
  assign \s00.Adr  [15] = 1'b1;
  assign \s00.Adr  [14] = 1'b0;
  assign \s00.Adr  [13] = 1'b0;
  assign \s00.Adr  [12] = 1'b0;
  assign \s00.Adr  [11] = 1'b1;
  assign \s00.Adr  [10] = 1'b1;
  assign \s01.Adr  [47] = 1'b0;
  assign \s01.Adr  [46] = 1'b0;
  assign \s01.Adr  [45] = 1'b0;
  assign \s01.Adr  [44] = 1'b0;
  assign \s01.Adr  [43] = 1'b0;
  assign \s01.Adr  [42] = 1'b0;
  assign \s01.Adr  [41] = 1'b0;
  assign \s01.Adr  [40] = 1'b0;
  assign \s01.Adr  [39] = 1'b0;
  assign \s01.Adr  [38] = 1'b0;
  assign \s01.Adr  [37] = 1'b0;
  assign \s01.Adr  [36] = 1'b0;
  assign \s01.Adr  [35] = 1'b0;
  assign \s01.Adr  [34] = 1'b0;
  assign \s01.Adr  [33] = 1'b0;
  assign \s01.Adr  [32] = 1'b0;
  assign \s01.Adr  [31] = 1'b0;
  assign \s01.Adr  [30] = 1'b0;
  assign \s01.Adr  [29] = 1'b0;
  assign \s01.Adr  [28] = 1'b0;
  assign \s01.Adr  [27] = 1'b0;
  assign \s01.Adr  [26] = 1'b0;
  assign \s01.Adr  [25] = 1'b0;
  assign \s01.Adr  [24] = 1'b0;
  assign \s01.Adr  [23] = 1'b1;
  assign \s01.Adr  [22] = 1'b1;
  assign \s01.Adr  [21] = 1'b1;
  assign \s01.Adr  [20] = 1'b1;
  assign \s01.Adr  [19] = 1'b1;
  assign \s01.Adr  [18] = 1'b1;
  assign \s01.Adr  [17] = 1'b1;
  assign \s01.Adr  [16] = 1'b1;
  assign \s01.Adr  [15] = 1'b0;
  assign \s01.Adr  [14] = 1'b1;
  assign \s01.Adr  [13] = 1'b1;
  assign \s01.Adr  [12] = 1'b1;
  assign \s01.Adr  [11] = 1'b0;
  assign \s01.Adr  [10] = 1'b0;
  assign \s01.Adr  [9] = 1'b0;
  assign \s01.Adr  [8] = 1'b0;
  assign \s02.Adr  [47] = 1'b0;
  assign \s02.Adr  [46] = 1'b0;
  assign \s02.Adr  [45] = 1'b0;
  assign \s02.Adr  [44] = 1'b0;
  assign \s02.Adr  [43] = 1'b0;
  assign \s02.Adr  [42] = 1'b0;
  assign \s02.Adr  [41] = 1'b0;
  assign \s02.Adr  [40] = 1'b0;
  assign \s02.Adr  [39] = 1'b0;
  assign \s02.Adr  [38] = 1'b0;
  assign \s02.Adr  [37] = 1'b0;
  assign \s02.Adr  [36] = 1'b0;
  assign \s02.Adr  [35] = 1'b0;
  assign \s02.Adr  [34] = 1'b0;
  assign \s02.Adr  [33] = 1'b0;
  assign \s02.Adr  [32] = 1'b0;
  assign \s02.Adr  [31] = 1'b0;
  assign \s02.Adr  [30] = 1'b0;
  assign \s02.Adr  [29] = 1'b0;
  assign \s02.Adr  [28] = 1'b0;
  assign \s02.Adr  [27] = 1'b0;
  assign \s02.Adr  [26] = 1'b0;
  assign \s02.Adr  [25] = 1'b0;
  assign \s02.Adr  [24] = 1'b0;
  assign \s02.Adr  [23] = 1'b1;
  assign \s02.Adr  [22] = 1'b1;
  assign \s02.Adr  [21] = 1'b1;
  assign \s02.Adr  [20] = 1'b1;
  assign \s02.Adr  [19] = 1'b1;
  assign \s02.Adr  [18] = 1'b1;
  assign \s02.Adr  [17] = 1'b1;
  assign \s02.Adr  [16] = 1'b1;
  assign \s02.Adr  [15] = 1'b0;
  assign \s02.Adr  [14] = 1'b1;
  assign \s02.Adr  [13] = 1'b0;
  assign \s02.Adr  [12] = 1'b1;
  assign \s02.Adr  [11] = 1'b1;
  assign \s02.Adr  [10] = 1'b0;
  assign \s02.Adr  [9] = 1'b0;
  assign \s02.Adr  [8] = 1'b0;
  assign \s02.Adr  [7] = 1'b1;
  assign \s02.Adr  [6] = 1'b1;
  assign \s02.Adr  [5] = 1'b0;
  assign \s03.Adr  [47] = 1'b0;
  assign \s03.Adr  [46] = 1'b0;
  assign \s03.Adr  [45] = 1'b0;
  assign \s03.Adr  [44] = 1'b0;
  assign \s03.Adr  [43] = 1'b0;
  assign \s03.Adr  [42] = 1'b0;
  assign \s03.Adr  [41] = 1'b0;
  assign \s03.Adr  [40] = 1'b0;
  assign \s03.Adr  [39] = 1'b0;
  assign \s03.Adr  [38] = 1'b0;
  assign \s03.Adr  [37] = 1'b0;
  assign \s03.Adr  [36] = 1'b0;
  assign \s03.Adr  [35] = 1'b0;
  assign \s03.Adr  [34] = 1'b0;
  assign \s03.Adr  [33] = 1'b0;
  assign \s03.Adr  [32] = 1'b0;
  assign \s03.Adr  [31] = 1'b0;
  assign \s03.Adr  [30] = 1'b0;
  assign \s03.Adr  [29] = 1'b0;
  assign \s03.Adr  [28] = 1'b0;
  assign \s03.Adr  [27] = 1'b0;
  assign \s03.Adr  [26] = 1'b0;
  assign \s03.Adr  [25] = 1'b0;
  assign \s03.Adr  [24] = 1'b0;
  assign \s03.Adr  [23] = 1'b1;
  assign \s03.Adr  [22] = 1'b1;
  assign \s03.Adr  [21] = 1'b1;
  assign \s03.Adr  [20] = 1'b1;
  assign \s03.Adr  [19] = 1'b1;
  assign \s03.Adr  [18] = 1'b1;
  assign \s03.Adr  [17] = 1'b1;
  assign \s03.Adr  [16] = 1'b1;
  assign \s03.Adr  [15] = 1'b0;
  assign \s03.Adr  [14] = 1'b0;
  assign \s03.Adr  [13] = 1'b1;
  assign \s03.Adr  [12] = 1'b1;
  assign \s03.Adr  [11] = 1'b1;
  assign \s03.Adr  [10] = 1'b1;
  assign \s03.Adr  [9] = 1'b0;
  assign \s04.Adr  [47] = 1'b0;
  assign \s04.Adr  [46] = 1'b0;
  assign \s04.Adr  [45] = 1'b0;
  assign \s04.Adr  [44] = 1'b0;
  assign \s04.Adr  [43] = 1'b0;
  assign \s04.Adr  [42] = 1'b0;
  assign \s04.Adr  [41] = 1'b0;
  assign \s04.Adr  [40] = 1'b0;
  assign \s04.Adr  [39] = 1'b0;
  assign \s04.Adr  [38] = 1'b0;
  assign \s04.Adr  [37] = 1'b0;
  assign \s04.Adr  [36] = 1'b0;
  assign \s04.Adr  [35] = 1'b0;
  assign \s04.Adr  [34] = 1'b0;
  assign \s04.Adr  [33] = 1'b0;
  assign \s04.Adr  [32] = 1'b0;
  assign \s04.Adr  [31] = 1'b0;
  assign \s04.Adr  [30] = 1'b0;
  assign \s04.Adr  [29] = 1'b0;
  assign \s04.Adr  [28] = 1'b0;
  assign \s04.Adr  [27] = 1'b0;
  assign \s04.Adr  [26] = 1'b0;
  assign \s04.Adr  [25] = 1'b0;
  assign \s04.Adr  [24] = 1'b0;
  assign \s04.Adr  [23] = 1'b1;
  assign \s04.Adr  [22] = 1'b1;
  assign \s04.Adr  [21] = 1'b1;
  assign \s04.Adr  [20] = 1'b1;
  assign \s04.Adr  [19] = 1'b1;
  assign \s04.Adr  [18] = 1'b1;
  assign \s04.Adr  [17] = 1'b1;
  assign \s04.Adr  [16] = 1'b0;
  assign \s04.Adr  [15] = 1'b1;
  assign \s04.Adr  [14] = 1'b0;
  assign \s04.Adr  [13] = 1'b0;
  assign \s04.Adr  [12] = 1'b1;
  assign \s04.Adr  [11] = 1'b0;
  assign \s04.Adr  [10] = 1'b1;
  assign \s04.Adr  [9] = 1'b0;
  assign \s04.Adr  [8] = 1'b1;
  assign \s04.Adr  [7] = 1'b0;
  assign \s05.Adr  [47] = 1'b0;
  assign \s05.Adr  [46] = 1'b0;
  assign \s05.Adr  [45] = 1'b0;
  assign \s05.Adr  [44] = 1'b0;
  assign \s05.Adr  [43] = 1'b0;
  assign \s05.Adr  [42] = 1'b0;
  assign \s05.Adr  [41] = 1'b0;
  assign \s05.Adr  [40] = 1'b0;
  assign \s05.Adr  [39] = 1'b0;
  assign \s05.Adr  [38] = 1'b0;
  assign \s05.Adr  [37] = 1'b0;
  assign \s05.Adr  [36] = 1'b0;
  assign \s05.Adr  [35] = 1'b0;
  assign \s05.Adr  [34] = 1'b0;
  assign \s05.Adr  [33] = 1'b0;
  assign \s05.Adr  [32] = 1'b0;
  assign \s05.Adr  [31] = 1'b0;
  assign \s05.Adr  [30] = 1'b0;
  assign \s05.Adr  [29] = 1'b0;
  assign \s05.Adr  [28] = 1'b0;
  assign \s05.Adr  [27] = 1'b0;
  assign \s05.Adr  [26] = 1'b0;
  assign \s05.Adr  [25] = 1'b0;
  assign \s05.Adr  [24] = 1'b0;
  assign \s05.Adr  [23] = 1'b1;
  assign \s05.Adr  [22] = 1'b1;
  assign \s05.Adr  [21] = 1'b1;
  assign \s05.Adr  [20] = 1'b1;
  assign \s05.Adr  [19] = 1'b1;
  assign \s05.Adr  [18] = 1'b1;
  assign \s05.Adr  [17] = 1'b1;
  assign \s05.Adr  [16] = 1'b0;
  assign \s05.Adr  [15] = 1'b1;
  assign \s05.Adr  [14] = 1'b0;
  assign \s05.Adr  [13] = 1'b0;
  assign \s05.Adr  [12] = 1'b1;
  assign \s05.Adr  [11] = 1'b0;
  assign \s05.Adr  [10] = 1'b0;
  assign \s05.Adr  [9] = 1'b1;
  assign \s05.Adr  [8] = 1'b1;
  assign \s05.Adr  [7] = 1'b1;
  assign \s05.Adr  [6] = 1'b1;
  assign \s05.Adr  [5] = 1'b1;
  assign \s06.Adr  [47] = 1'b0;
  assign \s06.Adr  [46] = 1'b0;
  assign \s06.Adr  [45] = 1'b0;
  assign \s06.Adr  [44] = 1'b0;
  assign \s06.Adr  [43] = 1'b0;
  assign \s06.Adr  [42] = 1'b0;
  assign \s06.Adr  [41] = 1'b0;
  assign \s06.Adr  [40] = 1'b0;
  assign \s06.Adr  [39] = 1'b0;
  assign \s06.Adr  [38] = 1'b0;
  assign \s06.Adr  [37] = 1'b0;
  assign \s06.Adr  [36] = 1'b0;
  assign \s06.Adr  [35] = 1'b0;
  assign \s06.Adr  [34] = 1'b0;
  assign \s06.Adr  [33] = 1'b0;
  assign \s06.Adr  [32] = 1'b0;
  assign \s06.Adr  [31] = 1'b0;
  assign \s06.Adr  [30] = 1'b0;
  assign \s06.Adr  [29] = 1'b0;
  assign \s06.Adr  [28] = 1'b0;
  assign \s06.Adr  [27] = 1'b0;
  assign \s06.Adr  [26] = 1'b0;
  assign \s06.Adr  [25] = 1'b0;
  assign \s06.Adr  [24] = 1'b0;
  assign \s06.Adr  [23] = 1'b1;
  assign \s06.Adr  [22] = 1'b1;
  assign \s06.Adr  [21] = 1'b1;
  assign \s06.Adr  [20] = 1'b1;
  assign \s06.Adr  [19] = 1'b1;
  assign \s06.Adr  [18] = 1'b1;
  assign \s06.Adr  [17] = 1'b1;
  assign \s06.Adr  [16] = 1'b1;
  assign \s06.Adr  [15] = 1'b0;
  assign \s06.Adr  [14] = 1'b1;
  assign \s06.Adr  [13] = 1'b0;
  assign \s06.Adr  [12] = 1'b1;
  assign \s06.Adr  [11] = 1'b0;
  assign \s06.Adr  [10] = 1'b0;
  assign \s06.Adr  [9] = 1'b1;
  assign \s06.Adr  [8] = 1'b1;
  assign \s06.Adr  [7] = 1'b0;
  assign \s06.Adr  [6] = 1'b1;
  assign \s07.Adr  [47] = 1'b0;
  assign \s07.Adr  [46] = 1'b0;
  assign \s07.Adr  [45] = 1'b0;
  assign \s07.Adr  [44] = 1'b0;
  assign \s07.Adr  [43] = 1'b0;
  assign \s07.Adr  [42] = 1'b0;
  assign \s07.Adr  [41] = 1'b0;
  assign \s07.Adr  [40] = 1'b0;
  assign \s07.Adr  [39] = 1'b0;
  assign \s07.Adr  [38] = 1'b0;
  assign \s07.Adr  [37] = 1'b0;
  assign \s07.Adr  [36] = 1'b0;
  assign \s07.Adr  [35] = 1'b0;
  assign \s07.Adr  [34] = 1'b0;
  assign \s07.Adr  [33] = 1'b0;
  assign \s07.Adr  [32] = 1'b0;
  assign \s07.Adr  [31] = 1'b0;
  assign \s07.Adr  [30] = 1'b0;
  assign \s07.Adr  [29] = 1'b0;
  assign \s07.Adr  [28] = 1'b0;
  assign \s07.Adr  [27] = 1'b0;
  assign \s07.Adr  [26] = 1'b0;
  assign \s07.Adr  [25] = 1'b0;
  assign \s07.Adr  [24] = 1'b0;
  assign \s07.Adr  [23] = 1'b1;
  assign \s07.Adr  [22] = 1'b1;
  assign \s07.Adr  [21] = 1'b1;
  assign \s07.Adr  [20] = 1'b1;
  assign \s07.Adr  [19] = 1'b1;
  assign \s07.Adr  [18] = 1'b1;
  assign \s07.Adr  [17] = 1'b1;
  assign \s07.Adr  [16] = 1'b1;
  assign \s07.Adr  [15] = 1'b1;
  assign \s07.Adr  [14] = 1'b1;
  assign \s07.Adr  [13] = 1'b1;
  assign \s07.Adr  [12] = 1'b1;
  assign \s07.Adr  [11] = 1'b1;
  assign \s07.Adr  [10] = 1'b1;
  assign \s07.Adr  [9] = 1'b0;
  assign \s08.Adr  [47] = 1'b0;
  assign \s08.Adr  [46] = 1'b0;
  assign \s08.Adr  [45] = 1'b0;
  assign \s08.Adr  [44] = 1'b0;
  assign \s08.Adr  [43] = 1'b0;
  assign \s08.Adr  [42] = 1'b0;
  assign \s08.Adr  [41] = 1'b0;
  assign \s08.Adr  [40] = 1'b0;
  assign \s08.Adr  [39] = 1'b0;
  assign \s08.Adr  [38] = 1'b0;
  assign \s08.Adr  [37] = 1'b0;
  assign \s08.Adr  [36] = 1'b0;
  assign \s08.Adr  [35] = 1'b0;
  assign \s08.Adr  [34] = 1'b0;
  assign \s08.Adr  [33] = 1'b0;
  assign \s08.Adr  [32] = 1'b0;
  assign \s08.Adr  [31] = 1'b0;
  assign \s08.Adr  [30] = 1'b0;
  assign \s08.Adr  [29] = 1'b0;
  assign \s08.Adr  [28] = 1'b0;
  assign \s08.Adr  [27] = 1'b0;
  assign \s08.Adr  [26] = 1'b0;
  assign \s08.Adr  [25] = 1'b0;
  assign \s08.Adr  [24] = 1'b0;
  assign \s08.Adr  [23] = 1'b1;
  assign \s08.Adr  [22] = 1'b1;
  assign \s08.Adr  [21] = 1'b1;
  assign \s08.Adr  [20] = 1'b1;
  assign \s08.Adr  [19] = 1'b1;
  assign \s08.Adr  [18] = 1'b1;
  assign \s08.Adr  [17] = 1'b1;
  assign \s08.Adr  [16] = 1'b1;
  assign \s08.Adr  [15] = 1'b0;
  assign \s08.Adr  [14] = 1'b0;
  assign \s08.Adr  [13] = 1'b1;
  assign \s08.Adr  [12] = 1'b1;
  assign \s08.Adr  [11] = 1'b0;
  assign \s08.Adr  [10] = 1'b0;
  assign \s08.Adr  [9] = 1'b0;
  assign \s09.Adr  [47] = 1'b0;
  assign \s09.Adr  [46] = 1'b0;
  assign \s09.Adr  [45] = 1'b0;
  assign \s09.Adr  [44] = 1'b0;
  assign \s09.Adr  [43] = 1'b0;
  assign \s09.Adr  [42] = 1'b0;
  assign \s09.Adr  [41] = 1'b0;
  assign \s09.Adr  [40] = 1'b0;
  assign \s09.Adr  [39] = 1'b0;
  assign \s09.Adr  [38] = 1'b0;
  assign \s09.Adr  [37] = 1'b0;
  assign \s09.Adr  [36] = 1'b0;
  assign \s09.Adr  [35] = 1'b0;
  assign \s09.Adr  [34] = 1'b0;
  assign \s09.Adr  [33] = 1'b0;
  assign \s09.Adr  [32] = 1'b0;
  assign \s09.Adr  [31] = 1'b0;
  assign \s09.Adr  [30] = 1'b0;
  assign \s09.Adr  [29] = 1'b0;
  assign \s09.Adr  [28] = 1'b0;
  assign \s09.Adr  [27] = 1'b0;
  assign \s09.Adr  [26] = 1'b0;
  assign \s09.Adr  [25] = 1'b0;
  assign \s09.Adr  [24] = 1'b0;
  assign \s09.Adr  [23] = 1'b1;
  assign \s09.Adr  [22] = 1'b1;
  assign \s09.Adr  [21] = 1'b1;
  assign \s09.Adr  [20] = 1'b1;
  assign \s09.Adr  [19] = 1'b1;
  assign \s09.Adr  [18] = 1'b1;
  assign \s09.Adr  [17] = 1'b1;
  assign \s09.Adr  [16] = 1'b1;
  assign \s09.Adr  [15] = 1'b0;
  assign \s09.Adr  [14] = 1'b1;
  assign \s09.Adr  [13] = 1'b1;
  assign \s09.Adr  [12] = 1'b1;
  assign \s09.Adr  [11] = 1'b1;
  assign \s09.Adr  [10] = 1'b1;
  assign \s09.Adr  [9] = 1'b0;
  assign \s09.Adr  [8] = 1'b1;
  assign \s10.Adr  [47] = 1'b0;
  assign \s10.Adr  [46] = 1'b0;
  assign \s10.Adr  [45] = 1'b0;
  assign \s10.Adr  [44] = 1'b0;
  assign \s10.Adr  [43] = 1'b0;
  assign \s10.Adr  [42] = 1'b0;
  assign \s10.Adr  [41] = 1'b0;
  assign \s10.Adr  [40] = 1'b0;
  assign \s10.Adr  [39] = 1'b0;
  assign \s10.Adr  [38] = 1'b0;
  assign \s10.Adr  [37] = 1'b0;
  assign \s10.Adr  [36] = 1'b0;
  assign \s10.Adr  [35] = 1'b0;
  assign \s10.Adr  [34] = 1'b0;
  assign \s10.Adr  [33] = 1'b0;
  assign \s10.Adr  [32] = 1'b0;
  assign \s10.Adr  [31] = 1'b0;
  assign \s10.Adr  [30] = 1'b0;
  assign \s10.Adr  [29] = 1'b0;
  assign \s10.Adr  [28] = 1'b0;
  assign \s10.Adr  [27] = 1'b0;
  assign \s10.Adr  [26] = 1'b0;
  assign \s10.Adr  [25] = 1'b0;
  assign \s10.Adr  [24] = 1'b0;
  assign \s10.Adr  [23] = 1'b1;
  assign \s10.Adr  [22] = 1'b1;
  assign \s10.Adr  [21] = 1'b1;
  assign \s10.Adr  [20] = 1'b1;
  assign \s10.Adr  [19] = 1'b1;
  assign \s10.Adr  [18] = 1'b1;
  assign \s10.Adr  [17] = 1'b1;
  assign \s10.Adr  [16] = 1'b1;
  assign \s10.Adr  [15] = 1'b0;
  assign \s10.Adr  [14] = 1'b1;
  assign \s10.Adr  [13] = 1'b1;
  assign \s10.Adr  [12] = 1'b0;
  assign \s10.Adr  [11] = 1'b0;
  assign \s10.Adr  [10] = 1'b1;
  assign \s10.Adr  [9] = 1'b0;
  assign \s10.Adr  [8] = 1'b1;
  assign \s10.Adr  [7] = 1'b0;
  assign \s11.Adr  [47] = 1'b0;
  assign \s11.Adr  [46] = 1'b0;
  assign \s11.Adr  [45] = 1'b0;
  assign \s11.Adr  [44] = 1'b0;
  assign \s11.Adr  [43] = 1'b0;
  assign \s11.Adr  [42] = 1'b0;
  assign \s11.Adr  [41] = 1'b0;
  assign \s11.Adr  [40] = 1'b0;
  assign \s11.Adr  [39] = 1'b0;
  assign \s11.Adr  [38] = 1'b0;
  assign \s11.Adr  [37] = 1'b0;
  assign \s11.Adr  [36] = 1'b0;
  assign \s11.Adr  [35] = 1'b0;
  assign \s11.Adr  [34] = 1'b0;
  assign \s11.Adr  [33] = 1'b0;
  assign \s11.Adr  [32] = 1'b0;
  assign \s11.Adr  [31] = 1'b0;
  assign \s11.Adr  [30] = 1'b0;
  assign \s11.Adr  [29] = 1'b0;
  assign \s11.Adr  [28] = 1'b0;
  assign \s11.Adr  [27] = 1'b0;
  assign \s11.Adr  [26] = 1'b0;
  assign \s11.Adr  [25] = 1'b0;
  assign \s11.Adr  [24] = 1'b0;
  assign \s11.Adr  [23] = 1'b1;
  assign \s11.Adr  [22] = 1'b1;
  assign \s11.Adr  [21] = 1'b1;
  assign \s11.Adr  [20] = 1'b1;
  assign \s11.Adr  [19] = 1'b1;
  assign \s11.Adr  [18] = 1'b1;
  assign \s11.Adr  [17] = 1'b1;
  assign \s11.Adr  [16] = 1'b1;
  assign \s11.Adr  [15] = 1'b0;
  assign \s11.Adr  [14] = 1'b1;
  assign \s11.Adr  [13] = 1'b0;
  assign \s11.Adr  [12] = 1'b0;
  assign \s11.Adr  [11] = 1'b0;
  assign \s11.Adr  [10] = 1'b0;
  assign \s11.Adr  [9] = 1'b0;
  assign \s12.Adr  [47] = 1'b0;
  assign \s12.Adr  [46] = 1'b0;
  assign \s12.Adr  [45] = 1'b0;
  assign \s12.Adr  [44] = 1'b0;
  assign \s12.Adr  [43] = 1'b0;
  assign \s12.Adr  [42] = 1'b0;
  assign \s12.Adr  [41] = 1'b0;
  assign \s12.Adr  [40] = 1'b0;
  assign \s12.Adr  [39] = 1'b0;
  assign \s12.Adr  [38] = 1'b0;
  assign \s12.Adr  [37] = 1'b0;
  assign \s12.Adr  [36] = 1'b0;
  assign \s12.Adr  [35] = 1'b0;
  assign \s12.Adr  [34] = 1'b0;
  assign \s12.Adr  [33] = 1'b0;
  assign \s12.Adr  [32] = 1'b0;
  assign \s12.Adr  [31] = 1'b0;
  assign \s12.Adr  [30] = 1'b0;
  assign \s12.Adr  [29] = 1'b0;
  assign \s12.Adr  [28] = 1'b0;
  assign \s12.Adr  [27] = 1'b0;
  assign \s12.Adr  [26] = 1'b0;
  assign \s12.Adr  [25] = 1'b0;
  assign \s12.Adr  [24] = 1'b0;
  assign \s12.Adr  [23] = 1'b1;
  assign \s12.Adr  [22] = 1'b1;
  assign \s12.Adr  [21] = 1'b1;
  assign \s12.Adr  [20] = 1'b1;
  assign \s12.Adr  [19] = 1'b1;
  assign \s12.Adr  [18] = 1'b1;
  assign \s12.Adr  [17] = 1'b1;
  assign \s12.Adr  [16] = 1'b1;
  assign \s12.Adr  [15] = 1'b1;
  assign \s12.Adr  [14] = 1'b0;
  assign \s12.Adr  [13] = 1'b1;
  assign \s12.Adr  [12] = 1'b0;
  assign \s12.Adr  [11] = 1'b1;
  assign \s12.Adr  [10] = 1'b0;
  assign \s12.Adr  [9] = 1'b1;
  assign \s13.Adr  [47] = 1'b0;
  assign \s13.Adr  [46] = 1'b0;
  assign \s13.Adr  [45] = 1'b0;
  assign \s13.Adr  [44] = 1'b0;
  assign \s13.Adr  [43] = 1'b0;
  assign \s13.Adr  [42] = 1'b0;
  assign \s13.Adr  [41] = 1'b0;
  assign \s13.Adr  [40] = 1'b0;
  assign \s13.Adr  [39] = 1'b0;
  assign \s13.Adr  [38] = 1'b0;
  assign \s13.Adr  [37] = 1'b0;
  assign \s13.Adr  [36] = 1'b0;
  assign \s13.Adr  [35] = 1'b0;
  assign \s13.Adr  [34] = 1'b0;
  assign \s13.Adr  [33] = 1'b0;
  assign \s13.Adr  [32] = 1'b0;
  assign \s13.Adr  [31] = 1'b0;
  assign \s13.Adr  [30] = 1'b0;
  assign \s13.Adr  [29] = 1'b0;
  assign \s13.Adr  [28] = 1'b0;
  assign \s13.Adr  [27] = 1'b0;
  assign \s13.Adr  [26] = 1'b0;
  assign \s13.Adr  [25] = 1'b0;
  assign \s13.Adr  [24] = 1'b0;
  assign \s13.Adr  [23] = 1'b1;
  assign \s13.Adr  [22] = 1'b1;
  assign \s13.Adr  [21] = 1'b1;
  assign \s13.Adr  [20] = 1'b1;
  assign \s13.Adr  [19] = 1'b1;
  assign \s13.Adr  [18] = 1'b1;
  assign \s13.Adr  [17] = 1'b1;
  assign \s13.Adr  [16] = 1'b1;
  assign \s13.Adr  [15] = 1'b0;
  assign \s13.Adr  [14] = 1'b1;
  assign \s13.Adr  [13] = 1'b1;
  assign \s13.Adr  [12] = 1'b0;
  assign \s13.Adr  [11] = 1'b0;
  assign \s13.Adr  [10] = 1'b0;
  assign \s13.Adr  [9] = 1'b0;

  CFD1QXL \s12.dbus_in_reg[15]  ( .D(n5185), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [15]) );
  CFD1QXL \s12.dbus_in_reg[14]  ( .D(n5184), .CP(n7740), .Q(\s12.dbus_in [14])
         );
  CFD1QXL \s12.dbus_in_reg[13]  ( .D(n5183), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [13]) );
  CFD1QXL \s12.dbus_in_reg[12]  ( .D(n5182), .CP(n7740), .Q(\s12.dbus_in [12])
         );
  CFD1QXL \s12.dbus_in_reg[11]  ( .D(n5181), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [11]) );
  CFD1QXL \s12.dbus_in_reg[10]  ( .D(n5180), .CP(n7740), .Q(\s12.dbus_in [10])
         );
  CFD1QXL \s12.dbus_in_reg[9]  ( .D(n5179), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [9]) );
  CFD1QXL \s12.dbus_in_reg[8]  ( .D(n5178), .CP(n7740), .Q(\s12.dbus_in [8])
         );
  CFD1QXL \s12.dbus_in_reg[7]  ( .D(n5177), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [7]) );
  CFD1QXL \s12.dbus_in_reg[6]  ( .D(n5176), .CP(n7740), .Q(\s12.dbus_in [6])
         );
  CFD1QXL \s12.dbus_in_reg[5]  ( .D(n5175), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [5]) );
  CFD1QXL \s12.dbus_in_reg[4]  ( .D(n5174), .CP(n7740), .Q(\s12.dbus_in [4])
         );
  CFD1QXL \s12.dbus_in_reg[3]  ( .D(n5173), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [3]) );
  CFD1QXL \s12.dbus_in_reg[2]  ( .D(n5172), .CP(n7740), .Q(\s12.dbus_in [2])
         );
  CFD1QXL \s12.dbus_in_reg[1]  ( .D(n5171), .CP(\clock.sysClk ), .Q(
        \s12.dbus_in [1]) );
  CFD1QXL \s12.dbus_in_reg[0]  ( .D(n5170), .CP(n7740), .Q(\s12.dbus_in [0])
         );
  CFD1QXL \s13.Adr_reg[8]  ( .D(n5130), .CP(\clock.sysClk ), .Q(\s13.Adr [8])
         );
  CFD1QXL \s13.Adr_reg[7]  ( .D(n5129), .CP(\clock.sysClk ), .Q(\s13.Adr [7])
         );
  CFD1QXL \s13.Adr_reg[6]  ( .D(n5128), .CP(n7739), .Q(\s13.Adr [6]) );
  CFD1QXL \s13.Adr_reg[5]  ( .D(n5127), .CP(\clock.sysClk ), .Q(\s13.Adr [5])
         );
  CFD1QXL \s13.Adr_reg[4]  ( .D(n5126), .CP(n7739), .Q(\s13.Adr [4]) );
  CFD1QXL \s13.Adr_reg[3]  ( .D(n5125), .CP(n7739), .Q(\s13.Adr [3]) );
  CFD1QXL \s13.Adr_reg[2]  ( .D(n5124), .CP(\clock.sysClk ), .Q(\s13.Adr [2])
         );
  CFD1QXL \s13.Adr_reg[1]  ( .D(n5123), .CP(n7739), .Q(\s13.Adr [1]) );
  CFD1QXL \s13.Adr_reg[0]  ( .D(n5122), .CP(n7739), .Q(\s13.Adr [0]) );
  CFD1QXL \s13.dbus_in_reg[15]  ( .D(n5121), .CP(\clock.sysClk ), .Q(
        \s13.dbus_in [15]) );
  CFD1QXL \s13.dbus_in_reg[14]  ( .D(n5120), .CP(n7739), .Q(\s13.dbus_in [14])
         );
  CFD1QXL \s13.dbus_in_reg[13]  ( .D(n5119), .CP(n7739), .Q(\s13.dbus_in [13])
         );
  CFD1QXL \s13.dbus_in_reg[12]  ( .D(n5118), .CP(\clock.sysClk ), .Q(
        \s13.dbus_in [12]) );
  CFD1QXL \s13.dbus_in_reg[11]  ( .D(n5117), .CP(n7738), .Q(\s13.dbus_in [11])
         );
  CFD1QXL \s13.dbus_in_reg[10]  ( .D(n5116), .CP(n7738), .Q(\s13.dbus_in [10])
         );
  CFD1QXL \s13.dbus_in_reg[9]  ( .D(n5115), .CP(n7738), .Q(\s13.dbus_in [9])
         );
  CFD1QXL \s13.dbus_in_reg[8]  ( .D(n5114), .CP(n7738), .Q(\s13.dbus_in [8])
         );
  CFD1QXL \s13.dbus_in_reg[7]  ( .D(n5113), .CP(n7738), .Q(\s13.dbus_in [7])
         );
  CFD1QXL \s13.dbus_in_reg[6]  ( .D(n5112), .CP(n7738), .Q(\s13.dbus_in [6])
         );
  CFD1QXL \s13.dbus_in_reg[5]  ( .D(n5111), .CP(n7738), .Q(\s13.dbus_in [5])
         );
  CFD1QXL \s13.dbus_in_reg[4]  ( .D(n5110), .CP(n7738), .Q(\s13.dbus_in [4])
         );
  CFD1QXL \s13.dbus_in_reg[3]  ( .D(n5109), .CP(n7738), .Q(\s13.dbus_in [3])
         );
  CFD1QXL \s13.dbus_in_reg[2]  ( .D(n5108), .CP(n7738), .Q(\s13.dbus_in [2])
         );
  CFD1QXL \s13.dbus_in_reg[1]  ( .D(n5107), .CP(n7738), .Q(\s13.dbus_in [1])
         );
  CFD1QXL \s13.dbus_in_reg[0]  ( .D(n5106), .CP(n7738), .Q(\s13.dbus_in [0])
         );
  CFD1QXL \s00.Adr_reg[8]  ( .D(n5066), .CP(n7746), .Q(\s00.Adr [8]) );
  CFD1QXL \s00.Adr_reg[7]  ( .D(n5065), .CP(n7746), .Q(\s00.Adr [7]) );
  CFD1QXL \s00.Adr_reg[6]  ( .D(n5064), .CP(n7746), .Q(\s00.Adr [6]) );
  CFD1QXL \s00.Adr_reg[5]  ( .D(n5063), .CP(n7744), .Q(\s00.Adr [5]) );
  CFD1QXL \s00.Adr_reg[4]  ( .D(n5062), .CP(n7745), .Q(\s00.Adr [4]) );
  CFD1QXL \s00.Adr_reg[3]  ( .D(n5061), .CP(n7739), .Q(\s00.Adr [3]) );
  CFD1QXL \s00.Adr_reg[2]  ( .D(n5060), .CP(n7746), .Q(\s00.Adr [2]) );
  CFD1QXL \s00.Adr_reg[1]  ( .D(n5059), .CP(n7741), .Q(\s00.Adr [1]) );
  CFD1QXL \s00.Adr_reg[0]  ( .D(n5058), .CP(n7742), .Q(\s00.Adr [0]) );
  CFD1QXL \s00.dbus_in_reg[15]  ( .D(n5057), .CP(n7737), .Q(\s00.dbus_in [15])
         );
  CFD1QXL \s00.dbus_in_reg[14]  ( .D(n5056), .CP(n7737), .Q(\s00.dbus_in [14])
         );
  CFD1QXL \s00.dbus_in_reg[13]  ( .D(n5055), .CP(n7737), .Q(\s00.dbus_in [13])
         );
  CFD1QXL \s00.dbus_in_reg[12]  ( .D(n5054), .CP(n7737), .Q(\s00.dbus_in [12])
         );
  CFD1QXL \s00.dbus_in_reg[11]  ( .D(n5053), .CP(n7737), .Q(\s00.dbus_in [11])
         );
  CFD1QXL \s00.dbus_in_reg[10]  ( .D(n5052), .CP(n7743), .Q(\s00.dbus_in [10])
         );
  CFD1QXL \s00.dbus_in_reg[9]  ( .D(n5051), .CP(n7737), .Q(\s00.dbus_in [9])
         );
  CFD1QXL \s00.dbus_in_reg[8]  ( .D(n5050), .CP(n7737), .Q(\s00.dbus_in [8])
         );
  CFD1QXL \s00.dbus_in_reg[7]  ( .D(n5049), .CP(n7744), .Q(\s00.dbus_in [7])
         );
  CFD1QXL \s00.dbus_in_reg[6]  ( .D(n5048), .CP(n7737), .Q(\s00.dbus_in [6])
         );
  CFD1QXL \s00.dbus_in_reg[5]  ( .D(n5047), .CP(n7745), .Q(\s00.dbus_in [5])
         );
  CFD1QXL \s00.dbus_in_reg[4]  ( .D(n5046), .CP(n7737), .Q(\s00.dbus_in [4])
         );
  CFD1QXL \s00.dbus_in_reg[3]  ( .D(n5045), .CP(n7745), .Q(\s00.dbus_in [3])
         );
  CFD1QXL \s00.dbus_in_reg[2]  ( .D(n5044), .CP(n7737), .Q(\s00.dbus_in [2])
         );
  CFD1QXL \s00.dbus_in_reg[1]  ( .D(n5043), .CP(n7736), .Q(\s00.dbus_in [1])
         );
  CFD1QXL \s00.dbus_in_reg[0]  ( .D(n5042), .CP(n7739), .Q(\s00.dbus_in [0])
         );
  CFD1QXL \s01.Adr_reg[7]  ( .D(n4985), .CP(n7745), .Q(\s01.Adr [7]) );
  CFD1QXL \s01.Adr_reg[6]  ( .D(n4984), .CP(n7745), .Q(\s01.Adr [6]) );
  CFD1QXL \s01.Adr_reg[5]  ( .D(n4983), .CP(n7745), .Q(\s01.Adr [5]) );
  CFD1QXL \s01.Adr_reg[4]  ( .D(n4982), .CP(n7745), .Q(\s01.Adr [4]) );
  CFD1QXL \s01.Adr_reg[3]  ( .D(n4981), .CP(n7745), .Q(\s01.Adr [3]) );
  CFD1QXL \s01.Adr_reg[2]  ( .D(n4980), .CP(n7745), .Q(\s01.Adr [2]) );
  CFD1QXL \s01.Adr_reg[1]  ( .D(n4979), .CP(n7744), .Q(\s01.Adr [1]) );
  CFD1QXL \s01.Adr_reg[0]  ( .D(n4978), .CP(n7744), .Q(\s01.Adr [0]) );
  CFD1QXL \s01.dbus_in_reg[15]  ( .D(n4977), .CP(n7744), .Q(\s01.dbus_in [15])
         );
  CFD1QXL \s01.dbus_in_reg[14]  ( .D(n4976), .CP(n7744), .Q(\s01.dbus_in [14])
         );
  CFD1QXL \s01.dbus_in_reg[13]  ( .D(n4975), .CP(n7744), .Q(\s01.dbus_in [13])
         );
  CFD1QXL \s01.dbus_in_reg[12]  ( .D(n4974), .CP(n7744), .Q(\s01.dbus_in [12])
         );
  CFD1QXL \s01.dbus_in_reg[11]  ( .D(n4973), .CP(n7743), .Q(\s01.dbus_in [11])
         );
  CFD1QXL \s01.dbus_in_reg[10]  ( .D(n4972), .CP(n7743), .Q(\s01.dbus_in [10])
         );
  CFD1QXL \s01.dbus_in_reg[9]  ( .D(n4971), .CP(n7743), .Q(\s01.dbus_in [9])
         );
  CFD1QXL \s01.dbus_in_reg[8]  ( .D(n4970), .CP(n7743), .Q(\s01.dbus_in [8])
         );
  CFD1QXL \s01.dbus_in_reg[7]  ( .D(n4969), .CP(n7743), .Q(\s01.dbus_in [7])
         );
  CFD1QXL \s01.dbus_in_reg[6]  ( .D(n4968), .CP(n7743), .Q(\s01.dbus_in [6])
         );
  CFD1QXL \s01.dbus_in_reg[5]  ( .D(n4967), .CP(n7742), .Q(\s01.dbus_in [5])
         );
  CFD1QXL \s01.dbus_in_reg[4]  ( .D(n4966), .CP(n7742), .Q(\s01.dbus_in [4])
         );
  CFD1QXL \s01.dbus_in_reg[3]  ( .D(n4965), .CP(n7742), .Q(\s01.dbus_in [3])
         );
  CFD1QXL \s01.dbus_in_reg[2]  ( .D(n4964), .CP(n7742), .Q(\s01.dbus_in [2])
         );
  CFD1QXL \s01.dbus_in_reg[1]  ( .D(n4963), .CP(n7742), .Q(\s01.dbus_in [1])
         );
  CFD1QXL \s01.dbus_in_reg[0]  ( .D(n4962), .CP(n7742), .Q(\s01.dbus_in [0])
         );
  CFD1QXL \s02.Adr_reg[4]  ( .D(n4918), .CP(n7746), .Q(\s02.Adr [4]) );
  CFD1QXL \s02.Adr_reg[3]  ( .D(n4917), .CP(n7741), .Q(\s02.Adr [3]) );
  CFD1QXL \s02.Adr_reg[2]  ( .D(n4916), .CP(n7732), .Q(\s02.Adr [2]) );
  CFD1QXL \s02.Adr_reg[1]  ( .D(n4915), .CP(n7740), .Q(\s02.Adr [1]) );
  CFD1QXL \s02.Adr_reg[0]  ( .D(n4914), .CP(n7742), .Q(\s02.Adr [0]) );
  CFD1QXL \s02.dbus_in_reg[15]  ( .D(n4913), .CP(n7735), .Q(\s02.dbus_in [15])
         );
  CFD1QXL \s02.dbus_in_reg[14]  ( .D(n4912), .CP(n7735), .Q(\s02.dbus_in [14])
         );
  CFD1QXL \s02.dbus_in_reg[13]  ( .D(n4911), .CP(n7735), .Q(\s02.dbus_in [13])
         );
  CFD1QXL \s02.dbus_in_reg[12]  ( .D(n4910), .CP(n7735), .Q(\s02.dbus_in [12])
         );
  CFD1QXL \s02.dbus_in_reg[11]  ( .D(n4909), .CP(n7743), .Q(\s02.dbus_in [11])
         );
  CFD1QXL \s02.dbus_in_reg[10]  ( .D(n4908), .CP(n7735), .Q(\s02.dbus_in [10])
         );
  CFD1QXL \s02.dbus_in_reg[9]  ( .D(n4907), .CP(n7735), .Q(\s02.dbus_in [9])
         );
  CFD1QXL \s02.dbus_in_reg[8]  ( .D(n4906), .CP(n7744), .Q(\s02.dbus_in [8])
         );
  CFD1QXL \s02.dbus_in_reg[7]  ( .D(n4905), .CP(n7735), .Q(\s02.dbus_in [7])
         );
  CFD1QXL \s02.dbus_in_reg[6]  ( .D(n4904), .CP(n7735), .Q(\s02.dbus_in [6])
         );
  CFD1QXL \s02.dbus_in_reg[5]  ( .D(n4903), .CP(n7735), .Q(\s02.dbus_in [5])
         );
  CFD1QXL \s02.dbus_in_reg[4]  ( .D(n4902), .CP(n7735), .Q(\s02.dbus_in [4])
         );
  CFD1QXL \s02.dbus_in_reg[3]  ( .D(n4901), .CP(n7741), .Q(\s02.dbus_in [3])
         );
  CFD1QXL \s02.dbus_in_reg[2]  ( .D(n4900), .CP(n7741), .Q(\s02.dbus_in [2])
         );
  CFD1QXL \s02.dbus_in_reg[1]  ( .D(n4899), .CP(n7741), .Q(\s02.dbus_in [1])
         );
  CFD1QXL \s02.dbus_in_reg[0]  ( .D(n4898), .CP(n7741), .Q(\s02.dbus_in [0])
         );
  CFD1QXL \s03.Adr_reg[8]  ( .D(n4858), .CP(n7726), .Q(\s03.Adr [8]) );
  CFD1QXL \s03.Adr_reg[7]  ( .D(n4857), .CP(n7733), .Q(\s03.Adr [7]) );
  CFD1QXL \s03.Adr_reg[6]  ( .D(n4856), .CP(n7738), .Q(\s03.Adr [6]) );
  CFD1QXL \s03.Adr_reg[5]  ( .D(n4855), .CP(n7739), .Q(\s03.Adr [5]) );
  CFD1QXL \s03.Adr_reg[4]  ( .D(n4854), .CP(n7746), .Q(\s03.Adr [4]) );
  CFD1QXL \s03.Adr_reg[3]  ( .D(n4853), .CP(n7741), .Q(\s03.Adr [3]) );
  CFD1QXL \s03.Adr_reg[2]  ( .D(n4852), .CP(n7736), .Q(\s03.Adr [2]) );
  CFD1QXL \s03.Adr_reg[1]  ( .D(n4851), .CP(n7731), .Q(\s03.Adr [1]) );
  CFD1QXL \s03.Adr_reg[0]  ( .D(n4850), .CP(n7732), .Q(\s03.Adr [0]) );
  CFD1QXL \s03.dbus_in_reg[15]  ( .D(n4849), .CP(n7740), .Q(\s03.dbus_in [15])
         );
  CFD1QXL \s03.dbus_in_reg[14]  ( .D(n4848), .CP(n7727), .Q(\s03.dbus_in [14])
         );
  CFD1QXL \s03.dbus_in_reg[13]  ( .D(n4847), .CP(n7728), .Q(\s03.dbus_in [13])
         );
  CFD1QXL \s03.dbus_in_reg[12]  ( .D(n4846), .CP(n7729), .Q(\s03.dbus_in [12])
         );
  CFD1QXL \s03.dbus_in_reg[11]  ( .D(n4845), .CP(n7730), .Q(\s03.dbus_in [11])
         );
  CFD1QXL \s03.dbus_in_reg[10]  ( .D(n4844), .CP(n7735), .Q(\s03.dbus_in [10])
         );
  CFD1QXL \s03.dbus_in_reg[9]  ( .D(n4843), .CP(n7742), .Q(\s03.dbus_in [9])
         );
  CFD1QXL \s03.dbus_in_reg[8]  ( .D(n4842), .CP(n7743), .Q(\s03.dbus_in [8])
         );
  CFD1QXL \s03.dbus_in_reg[7]  ( .D(n4841), .CP(n7744), .Q(\s03.dbus_in [7])
         );
  CFD1QXL \s03.dbus_in_reg[6]  ( .D(n4840), .CP(n7745), .Q(\s03.dbus_in [6])
         );
  CFD1QXL \s03.dbus_in_reg[5]  ( .D(n4839), .CP(n7737), .Q(\s03.dbus_in [5])
         );
  CFD1QXL \s03.dbus_in_reg[4]  ( .D(n4838), .CP(n7740), .Q(\s03.dbus_in [4])
         );
  CFD1QXL \s03.dbus_in_reg[3]  ( .D(n4837), .CP(n7734), .Q(\s03.dbus_in [3])
         );
  CFD1QXL \s03.dbus_in_reg[2]  ( .D(n4836), .CP(n7726), .Q(\s03.dbus_in [2])
         );
  CFD1QXL \s03.dbus_in_reg[1]  ( .D(n4835), .CP(n7733), .Q(\s03.dbus_in [1])
         );
  CFD1QXL \s03.dbus_in_reg[0]  ( .D(n4834), .CP(n7738), .Q(\s03.dbus_in [0])
         );
  CFD1QXL \s04.Adr_reg[6]  ( .D(n4792), .CP(n7740), .Q(\s04.Adr [6]) );
  CFD1QXL \s04.Adr_reg[5]  ( .D(n4791), .CP(n7740), .Q(\s04.Adr [5]) );
  CFD1QXL \s04.Adr_reg[4]  ( .D(n4790), .CP(n7740), .Q(\s04.Adr [4]) );
  CFD1QXL \s04.Adr_reg[3]  ( .D(n4789), .CP(n7740), .Q(\s04.Adr [3]) );
  CFD1QXL \s04.Adr_reg[2]  ( .D(n4788), .CP(n7740), .Q(\s04.Adr [2]) );
  CFD1QXL \s04.Adr_reg[1]  ( .D(n4787), .CP(n7734), .Q(\s04.Adr [1]) );
  CFD1QXL \s04.Adr_reg[0]  ( .D(n4786), .CP(n7734), .Q(\s04.Adr [0]) );
  CFD1QXL \s04.dbus_in_reg[15]  ( .D(n4785), .CP(n7734), .Q(\s04.dbus_in [15])
         );
  CFD1QXL \s04.dbus_in_reg[14]  ( .D(n4784), .CP(n7734), .Q(\s04.dbus_in [14])
         );
  CFD1QXL \s04.dbus_in_reg[13]  ( .D(n4783), .CP(n7740), .Q(\s04.dbus_in [13])
         );
  CFD1QXL \s04.dbus_in_reg[12]  ( .D(n4782), .CP(n7734), .Q(\s04.dbus_in [12])
         );
  CFD1QXL \s04.dbus_in_reg[11]  ( .D(n4781), .CP(n7734), .Q(\s04.dbus_in [11])
         );
  CFD1QXL \s04.dbus_in_reg[10]  ( .D(n4780), .CP(n7740), .Q(\s04.dbus_in [10])
         );
  CFD1QXL \s04.dbus_in_reg[9]  ( .D(n4779), .CP(n7734), .Q(\s04.dbus_in [9])
         );
  CFD1QXL \s04.dbus_in_reg[8]  ( .D(n4778), .CP(n7740), .Q(\s04.dbus_in [8])
         );
  CFD1QXL \s04.dbus_in_reg[7]  ( .D(n4777), .CP(n7734), .Q(\s04.dbus_in [7])
         );
  CFD1QXL \s04.dbus_in_reg[6]  ( .D(n4776), .CP(n7740), .Q(\s04.dbus_in [6])
         );
  CFD1QXL \s04.dbus_in_reg[5]  ( .D(n4775), .CP(n7733), .Q(\s04.dbus_in [5])
         );
  CFD1QXL \s04.dbus_in_reg[4]  ( .D(n4774), .CP(n7733), .Q(\s04.dbus_in [4])
         );
  CFD1QXL \s04.dbus_in_reg[3]  ( .D(n4773), .CP(n7733), .Q(\s04.dbus_in [3])
         );
  CFD1QXL \s04.dbus_in_reg[2]  ( .D(n4772), .CP(n7733), .Q(\s04.dbus_in [2])
         );
  CFD1QXL \s04.dbus_in_reg[1]  ( .D(n4771), .CP(n7733), .Q(\s04.dbus_in [1])
         );
  CFD1QXL \s04.dbus_in_reg[0]  ( .D(n4770), .CP(n7733), .Q(\s04.dbus_in [0])
         );
  CFD1QXL \s05.Adr_reg[4]  ( .D(n4726), .CP(n7733), .Q(\s05.Adr [4]) );
  CFD1QXL \s05.Adr_reg[3]  ( .D(n4725), .CP(n7733), .Q(\s05.Adr [3]) );
  CFD1QXL \s05.Adr_reg[2]  ( .D(n4724), .CP(n7733), .Q(\s05.Adr [2]) );
  CFD1QXL \s05.Adr_reg[1]  ( .D(n4723), .CP(n7733), .Q(\s05.Adr [1]) );
  CFD1QXL \s05.Adr_reg[0]  ( .D(n4722), .CP(n7733), .Q(\s05.Adr [0]) );
  CFD1QXL \s05.dbus_in_reg[15]  ( .D(n4721), .CP(n7732), .Q(\s05.dbus_in [15])
         );
  CFD1QXL \s05.dbus_in_reg[14]  ( .D(n4720), .CP(n7732), .Q(\s05.dbus_in [14])
         );
  CFD1QXL \s05.dbus_in_reg[13]  ( .D(n4719), .CP(n7732), .Q(\s05.dbus_in [13])
         );
  CFD1QXL \s05.dbus_in_reg[12]  ( .D(n4718), .CP(n7746), .Q(\s05.dbus_in [12])
         );
  CFD1QXL \s05.dbus_in_reg[11]  ( .D(n4717), .CP(n7732), .Q(\s05.dbus_in [11])
         );
  CFD1QXL \s05.dbus_in_reg[10]  ( .D(n4716), .CP(n7741), .Q(\s05.dbus_in [10])
         );
  CFD1QXL \s05.dbus_in_reg[9]  ( .D(n4715), .CP(n7732), .Q(\s05.dbus_in [9])
         );
  CFD1QXL \s05.dbus_in_reg[8]  ( .D(n4714), .CP(n7732), .Q(\s05.dbus_in [8])
         );
  CFD1QXL \s05.dbus_in_reg[7]  ( .D(n4713), .CP(n7742), .Q(\s05.dbus_in [7])
         );
  CFD1QXL \s05.dbus_in_reg[6]  ( .D(n4712), .CP(n7732), .Q(\s05.dbus_in [6])
         );
  CFD1QXL \s05.dbus_in_reg[5]  ( .D(n4711), .CP(n7743), .Q(\s05.dbus_in [5])
         );
  CFD1QXL \s05.dbus_in_reg[4]  ( .D(n4710), .CP(n7732), .Q(\s05.dbus_in [4])
         );
  CFD1QXL \s05.dbus_in_reg[3]  ( .D(n4709), .CP(n7744), .Q(\s05.dbus_in [3])
         );
  CFD1QXL \s05.dbus_in_reg[2]  ( .D(n4708), .CP(n7745), .Q(\s05.dbus_in [2])
         );
  CFD1QXL \s05.dbus_in_reg[1]  ( .D(n4707), .CP(n7746), .Q(\s05.dbus_in [1])
         );
  CFD1QXL \s05.dbus_in_reg[0]  ( .D(n4706), .CP(n7741), .Q(\s05.dbus_in [0])
         );
  CFD1QXL \s06.Adr_reg[5]  ( .D(n4663), .CP(n7729), .Q(\s06.Adr [5]) );
  CFD1QXL \s06.Adr_reg[4]  ( .D(n4662), .CP(n7730), .Q(\s06.Adr [4]) );
  CFD1QXL \s06.Adr_reg[3]  ( .D(n4661), .CP(n7735), .Q(\s06.Adr [3]) );
  CFD1QXL \s06.Adr_reg[2]  ( .D(n4660), .CP(n7742), .Q(\s06.Adr [2]) );
  CFD1QXL \s06.Adr_reg[1]  ( .D(n4659), .CP(n7743), .Q(\s06.Adr [1]) );
  CFD1QXL \s06.Adr_reg[0]  ( .D(n4658), .CP(n7744), .Q(\s06.Adr [0]) );
  CFD1QXL \s06.dbus_in_reg[15]  ( .D(n4657), .CP(n7745), .Q(\s06.dbus_in [15])
         );
  CFD1QXL \s06.dbus_in_reg[14]  ( .D(n4656), .CP(n7737), .Q(\s06.dbus_in [14])
         );
  CFD1QXL \s06.dbus_in_reg[13]  ( .D(n4655), .CP(n7734), .Q(\s06.dbus_in [13])
         );
  CFD1QXL \s06.dbus_in_reg[12]  ( .D(n4654), .CP(n7733), .Q(\s06.dbus_in [12])
         );
  CFD1QXL \s06.dbus_in_reg[11]  ( .D(n4653), .CP(n7738), .Q(\s06.dbus_in [11])
         );
  CFD1QXL \s06.dbus_in_reg[10]  ( .D(n4652), .CP(n7739), .Q(\s06.dbus_in [10])
         );
  CFD1QXL \s06.dbus_in_reg[9]  ( .D(n4651), .CP(n7746), .Q(\s06.dbus_in [9])
         );
  CFD1QXL \s06.dbus_in_reg[8]  ( .D(n4650), .CP(n7741), .Q(\s06.dbus_in [8])
         );
  CFD1QXL \s06.dbus_in_reg[7]  ( .D(n4649), .CP(n7736), .Q(\s06.dbus_in [7])
         );
  CFD1QXL \s06.dbus_in_reg[6]  ( .D(n4648), .CP(n7732), .Q(\s06.dbus_in [6])
         );
  CFD1QXL \s06.dbus_in_reg[5]  ( .D(n4647), .CP(n7740), .Q(\s06.dbus_in [5])
         );
  CFD1QXL \s06.dbus_in_reg[4]  ( .D(n4646), .CP(n7727), .Q(\s06.dbus_in [4])
         );
  CFD1QXL \s06.dbus_in_reg[3]  ( .D(n4645), .CP(n7730), .Q(\s06.dbus_in [3])
         );
  CFD1QXL \s06.dbus_in_reg[2]  ( .D(n4644), .CP(n7735), .Q(\s06.dbus_in [2])
         );
  CFD1QXL \s06.dbus_in_reg[1]  ( .D(n4643), .CP(n7742), .Q(\s06.dbus_in [1])
         );
  CFD1QXL \s06.dbus_in_reg[0]  ( .D(n4642), .CP(n7743), .Q(\s06.dbus_in [0])
         );
  CFD1QXL \s07.Adr_reg[8]  ( .D(n4602), .CP(n7731), .Q(\s07.Adr [8]) );
  CFD1QXL \s07.Adr_reg[7]  ( .D(n4601), .CP(n7744), .Q(\s07.Adr [7]) );
  CFD1QXL \s07.Adr_reg[6]  ( .D(n4600), .CP(n7745), .Q(\s07.Adr [6]) );
  CFD1QXL \s07.Adr_reg[5]  ( .D(n4599), .CP(n7731), .Q(\s07.Adr [5]) );
  CFD1QXL \s07.Adr_reg[4]  ( .D(n4598), .CP(n7737), .Q(\s07.Adr [4]) );
  CFD1QXL \s07.Adr_reg[3]  ( .D(n4597), .CP(n7731), .Q(\s07.Adr [3]) );
  CFD1QXL \s07.Adr_reg[2]  ( .D(n4596), .CP(n7731), .Q(\s07.Adr [2]) );
  CFD1QXL \s07.Adr_reg[1]  ( .D(n4595), .CP(n7734), .Q(\s07.Adr [1]) );
  CFD1QXL \s07.Adr_reg[0]  ( .D(n4594), .CP(n7731), .Q(\s07.Adr [0]) );
  CFD1QXL \s07.dbus_in_reg[15]  ( .D(n4593), .CP(n7733), .Q(\s07.dbus_in [15])
         );
  CFD1QXL \s07.dbus_in_reg[14]  ( .D(n4592), .CP(n7731), .Q(\s07.dbus_in [14])
         );
  CFD1QXL \s07.dbus_in_reg[13]  ( .D(n4591), .CP(n7739), .Q(\s07.dbus_in [13])
         );
  CFD1QXL \s07.dbus_in_reg[12]  ( .D(n4590), .CP(n7731), .Q(\s07.dbus_in [12])
         );
  CFD1QXL \s07.dbus_in_reg[11]  ( .D(n4589), .CP(n7746), .Q(\s07.dbus_in [11])
         );
  CFD1QXL \s07.dbus_in_reg[10]  ( .D(n4588), .CP(n7731), .Q(\s07.dbus_in [10])
         );
  CFD1QXL \s07.dbus_in_reg[9]  ( .D(n4587), .CP(n7741), .Q(\s07.dbus_in [9])
         );
  CFD1QXL \s07.dbus_in_reg[8]  ( .D(n4586), .CP(n7731), .Q(\s07.dbus_in [8])
         );
  CFD1QXL \s07.dbus_in_reg[7]  ( .D(n4585), .CP(n7731), .Q(\s07.dbus_in [7])
         );
  CFD1QXL \s07.dbus_in_reg[6]  ( .D(n4584), .CP(n7736), .Q(\s07.dbus_in [6])
         );
  CFD1QXL \s07.dbus_in_reg[5]  ( .D(n4583), .CP(n7732), .Q(\s07.dbus_in [5])
         );
  CFD1QXL \s07.dbus_in_reg[4]  ( .D(n4582), .CP(n7731), .Q(\s07.dbus_in [4])
         );
  CFD1QXL \s07.dbus_in_reg[3]  ( .D(n4581), .CP(n7740), .Q(\s07.dbus_in [3])
         );
  CFD1QXL \s07.dbus_in_reg[2]  ( .D(n4580), .CP(n7730), .Q(\s07.dbus_in [2])
         );
  CFD1QXL \s07.dbus_in_reg[1]  ( .D(n4579), .CP(n7731), .Q(\s07.dbus_in [1])
         );
  CFD1QXL \s07.dbus_in_reg[0]  ( .D(n4578), .CP(n7731), .Q(\s07.dbus_in [0])
         );
  CFD1QXL \s08.Adr_reg[8]  ( .D(n4538), .CP(n7737), .Q(\s08.Adr [8]) );
  CFD1QXL \s08.Adr_reg[7]  ( .D(n4537), .CP(\clock.sysClk ), .Q(\s08.Adr [7])
         );
  CFD1QXL \s08.Adr_reg[6]  ( .D(n4536), .CP(n7734), .Q(\s08.Adr [6]) );
  CFD1QXL \s08.Adr_reg[5]  ( .D(n4535), .CP(n7726), .Q(\s08.Adr [5]) );
  CFD1QXL \s08.Adr_reg[4]  ( .D(n4534), .CP(n7733), .Q(\s08.Adr [4]) );
  CFD1QXL \s08.Adr_reg[3]  ( .D(n4533), .CP(n7738), .Q(\s08.Adr [3]) );
  CFD1QXL \s08.Adr_reg[2]  ( .D(n4532), .CP(n7739), .Q(\s08.Adr [2]) );
  CFD1QXL \s08.Adr_reg[1]  ( .D(n4531), .CP(n7746), .Q(\s08.Adr [1]) );
  CFD1QXL \s08.Adr_reg[0]  ( .D(n4530), .CP(n7741), .Q(\s08.Adr [0]) );
  CFD1QXL \s08.dbus_in_reg[15]  ( .D(n4529), .CP(n7736), .Q(\s08.dbus_in [15])
         );
  CFD1QXL \s08.dbus_in_reg[14]  ( .D(n4528), .CP(n7731), .Q(\s08.dbus_in [14])
         );
  CFD1QXL \s08.dbus_in_reg[13]  ( .D(n4527), .CP(n7732), .Q(\s08.dbus_in [13])
         );
  CFD1QXL \s08.dbus_in_reg[12]  ( .D(n4526), .CP(n7740), .Q(\s08.dbus_in [12])
         );
  CFD1QXL \s08.dbus_in_reg[11]  ( .D(n4525), .CP(n7727), .Q(\s08.dbus_in [11])
         );
  CFD1QXL \s08.dbus_in_reg[10]  ( .D(n4524), .CP(n7728), .Q(\s08.dbus_in [10])
         );
  CFD1QXL \s08.dbus_in_reg[9]  ( .D(n4523), .CP(n7729), .Q(\s08.dbus_in [9])
         );
  CFD1QXL \s08.dbus_in_reg[8]  ( .D(n4522), .CP(n7730), .Q(\s08.dbus_in [8])
         );
  CFD1QXL \s08.dbus_in_reg[7]  ( .D(n4521), .CP(n7735), .Q(\s08.dbus_in [7])
         );
  CFD1QXL \s08.dbus_in_reg[6]  ( .D(n4520), .CP(n7742), .Q(\s08.dbus_in [6])
         );
  CFD1QXL \s08.dbus_in_reg[5]  ( .D(n4519), .CP(n7743), .Q(\s08.dbus_in [5])
         );
  CFD1QXL \s08.dbus_in_reg[4]  ( .D(n4518), .CP(n7744), .Q(\s08.dbus_in [4])
         );
  CFD1QXL \s08.dbus_in_reg[3]  ( .D(n4517), .CP(n7745), .Q(\s08.dbus_in [3])
         );
  CFD1QXL \s08.dbus_in_reg[2]  ( .D(n4516), .CP(n7737), .Q(\s08.dbus_in [2])
         );
  CFD1QXL \s08.dbus_in_reg[1]  ( .D(n4515), .CP(n7740), .Q(\s08.dbus_in [1])
         );
  CFD1QXL \s08.dbus_in_reg[0]  ( .D(n4514), .CP(n7734), .Q(\s08.dbus_in [0])
         );
  CFD1QXL \s09.Adr_reg[7]  ( .D(n4473), .CP(n7736), .Q(\s09.Adr [7]) );
  CFD1QXL \s09.Adr_reg[6]  ( .D(n4472), .CP(n7732), .Q(\s09.Adr [6]) );
  CFD1QXL \s09.Adr_reg[5]  ( .D(n4471), .CP(n7740), .Q(\s09.Adr [5]) );
  CFD1QXL \s09.Adr_reg[4]  ( .D(n4470), .CP(n7735), .Q(\s09.Adr [4]) );
  CFD1QXL \s09.Adr_reg[3]  ( .D(n4469), .CP(n7730), .Q(\s09.Adr [3]) );
  CFD1QXL \s09.Adr_reg[2]  ( .D(n4468), .CP(n7730), .Q(\s09.Adr [2]) );
  CFD1QXL \s09.Adr_reg[1]  ( .D(n4467), .CP(n7742), .Q(\s09.Adr [1]) );
  CFD1QXL \s09.Adr_reg[0]  ( .D(n4466), .CP(n7730), .Q(\s09.Adr [0]) );
  CFD1QXL \s09.dbus_in_reg[15]  ( .D(n4465), .CP(n7743), .Q(\s09.dbus_in [15])
         );
  CFD1QXL \s09.dbus_in_reg[14]  ( .D(n4464), .CP(n7730), .Q(\s09.dbus_in [14])
         );
  CFD1QXL \s09.dbus_in_reg[13]  ( .D(n4463), .CP(n7730), .Q(\s09.dbus_in [13])
         );
  CFD1QXL \s09.dbus_in_reg[12]  ( .D(n4462), .CP(n7744), .Q(\s09.dbus_in [12])
         );
  CFD1QXL \s09.dbus_in_reg[11]  ( .D(n4461), .CP(n7745), .Q(\s09.dbus_in [11])
         );
  CFD1QXL \s09.dbus_in_reg[10]  ( .D(n4460), .CP(n7730), .Q(\s09.dbus_in [10])
         );
  CFD1QXL \s09.dbus_in_reg[9]  ( .D(n4459), .CP(n7737), .Q(\s09.dbus_in [9])
         );
  CFD1QXL \s09.dbus_in_reg[8]  ( .D(n4458), .CP(n7730), .Q(\s09.dbus_in [8])
         );
  CFD1QXL \s09.dbus_in_reg[7]  ( .D(n4457), .CP(n7730), .Q(\s09.dbus_in [7])
         );
  CFD1QXL \s09.dbus_in_reg[6]  ( .D(n4456), .CP(n7730), .Q(\s09.dbus_in [6])
         );
  CFD1QXL \s09.dbus_in_reg[5]  ( .D(n4455), .CP(n7734), .Q(\s09.dbus_in [5])
         );
  CFD1QXL \s09.dbus_in_reg[4]  ( .D(n4454), .CP(n7730), .Q(\s09.dbus_in [4])
         );
  CFD1QXL \s09.dbus_in_reg[3]  ( .D(n4453), .CP(n7739), .Q(\s09.dbus_in [3])
         );
  CFD1QXL \s09.dbus_in_reg[2]  ( .D(n4452), .CP(n7730), .Q(\s09.dbus_in [2])
         );
  CFD1QXL \s09.dbus_in_reg[1]  ( .D(n4451), .CP(n7729), .Q(\s09.dbus_in [1])
         );
  CFD1QXL \s09.dbus_in_reg[0]  ( .D(n4450), .CP(n7729), .Q(\s09.dbus_in [0])
         );
  CFD1QXL \s10.Adr_reg[6]  ( .D(n4408), .CP(n7729), .Q(\s10.Adr [6]) );
  CFD1QXL \s10.Adr_reg[5]  ( .D(n4407), .CP(n7729), .Q(\s10.Adr [5]) );
  CFD1QXL \s10.Adr_reg[4]  ( .D(n4406), .CP(n7729), .Q(\s10.Adr [4]) );
  CFD1QXL \s10.Adr_reg[3]  ( .D(n4405), .CP(n7729), .Q(\s10.Adr [3]) );
  CFD1QXL \s10.Adr_reg[2]  ( .D(n4404), .CP(n7729), .Q(\s10.Adr [2]) );
  CFD1QXL \s10.Adr_reg[1]  ( .D(n4403), .CP(n7729), .Q(\s10.Adr [1]) );
  CFD1QXL \s10.Adr_reg[0]  ( .D(n4402), .CP(n7729), .Q(\s10.Adr [0]) );
  CFD1QXL \s10.dbus_in_reg[15]  ( .D(n4401), .CP(n7729), .Q(\s10.dbus_in [15])
         );
  CFD1QXL \s10.dbus_in_reg[14]  ( .D(n4400), .CP(n7729), .Q(\s10.dbus_in [14])
         );
  CFD1QXL \s10.dbus_in_reg[13]  ( .D(n4399), .CP(n7729), .Q(\s10.dbus_in [13])
         );
  CFD1QXL \s10.dbus_in_reg[12]  ( .D(n4398), .CP(n7729), .Q(\s10.dbus_in [12])
         );
  CFD1QXL \s10.dbus_in_reg[11]  ( .D(n4397), .CP(n7728), .Q(\s10.dbus_in [11])
         );
  CFD1QXL \s10.dbus_in_reg[10]  ( .D(n4396), .CP(n7728), .Q(\s10.dbus_in [10])
         );
  CFD1QXL \s10.dbus_in_reg[9]  ( .D(n4395), .CP(n7728), .Q(\s10.dbus_in [9])
         );
  CFD1QXL \s10.dbus_in_reg[8]  ( .D(n4394), .CP(n7728), .Q(\s10.dbus_in [8])
         );
  CFD1QXL \s10.dbus_in_reg[7]  ( .D(n4393), .CP(n7728), .Q(\s10.dbus_in [7])
         );
  CFD1QXL \s10.dbus_in_reg[6]  ( .D(n4392), .CP(n7728), .Q(\s10.dbus_in [6])
         );
  CFD1QXL \s10.dbus_in_reg[5]  ( .D(n4391), .CP(n7728), .Q(\s10.dbus_in [5])
         );
  CFD1QXL \s10.dbus_in_reg[4]  ( .D(n4390), .CP(n7728), .Q(\s10.dbus_in [4])
         );
  CFD1QXL \s10.dbus_in_reg[3]  ( .D(n4389), .CP(n7728), .Q(\s10.dbus_in [3])
         );
  CFD1QXL \s10.dbus_in_reg[2]  ( .D(n4388), .CP(n7728), .Q(\s10.dbus_in [2])
         );
  CFD1QXL \s10.dbus_in_reg[1]  ( .D(n4387), .CP(n7728), .Q(\s10.dbus_in [1])
         );
  CFD1QXL \s10.dbus_in_reg[0]  ( .D(n4386), .CP(n7728), .Q(\s10.dbus_in [0])
         );
  CFD1QXL \s11.Adr_reg[8]  ( .D(n4346), .CP(n7728), .Q(\s11.Adr [8]) );
  CFD1QXL \s11.Adr_reg[7]  ( .D(n4345), .CP(n7728), .Q(\s11.Adr [7]) );
  CFD1QXL \s11.Adr_reg[6]  ( .D(n4344), .CP(n7728), .Q(\s11.Adr [6]) );
  CFD1QXL \s11.Adr_reg[5]  ( .D(n4343), .CP(n7727), .Q(\s11.Adr [5]) );
  CFD1QXL \s11.Adr_reg[4]  ( .D(n4342), .CP(n7727), .Q(\s11.Adr [4]) );
  CFD1QXL \s11.Adr_reg[3]  ( .D(n4341), .CP(n7735), .Q(\s11.Adr [3]) );
  CFD1QXL \s11.Adr_reg[2]  ( .D(n4340), .CP(n7727), .Q(\s11.Adr [2]) );
  CFD1QXL \s11.Adr_reg[1]  ( .D(n4339), .CP(n7742), .Q(\s11.Adr [1]) );
  CFD1QXL \s11.Adr_reg[0]  ( .D(n4338), .CP(n7727), .Q(\s11.Adr [0]) );
  CFD1QXL \s11.dbus_in_reg[15]  ( .D(n4337), .CP(n7727), .Q(\s11.dbus_in [15])
         );
  CFD1QXL \s11.dbus_in_reg[14]  ( .D(n4336), .CP(n7743), .Q(\s11.dbus_in [14])
         );
  CFD1QXL \s11.dbus_in_reg[13]  ( .D(n4335), .CP(n7744), .Q(\s11.dbus_in [13])
         );
  CFD1QXL \s11.dbus_in_reg[12]  ( .D(n4334), .CP(n7727), .Q(\s11.dbus_in [12])
         );
  CFD1QXL \s11.dbus_in_reg[11]  ( .D(n4333), .CP(n7745), .Q(\s11.dbus_in [11])
         );
  CFD1QXL \s11.dbus_in_reg[10]  ( .D(n4332), .CP(n7727), .Q(\s11.dbus_in [10])
         );
  CFD1QXL \s11.dbus_in_reg[9]  ( .D(n4331), .CP(n7727), .Q(\s11.dbus_in [9])
         );
  CFD1QXL \s11.dbus_in_reg[8]  ( .D(n4330), .CP(n7727), .Q(\s11.dbus_in [8])
         );
  CFD1QXL \s11.dbus_in_reg[7]  ( .D(n4329), .CP(n7737), .Q(\s11.dbus_in [7])
         );
  CFD1QXL \s11.dbus_in_reg[6]  ( .D(n4328), .CP(n7727), .Q(\s11.dbus_in [6])
         );
  CFD1QXL \s11.dbus_in_reg[5]  ( .D(n4327), .CP(n7727), .Q(\s11.dbus_in [5])
         );
  CFD1QXL \s11.dbus_in_reg[4]  ( .D(n4326), .CP(n7727), .Q(\s11.dbus_in [4])
         );
  CFD1QXL \s11.dbus_in_reg[3]  ( .D(n4325), .CP(n7734), .Q(\s11.dbus_in [3])
         );
  CFD1QXL \s11.dbus_in_reg[2]  ( .D(n4324), .CP(n7739), .Q(\s11.dbus_in [2])
         );
  CFD1QXL \s11.dbus_in_reg[1]  ( .D(n4323), .CP(n7746), .Q(\s11.dbus_in [1])
         );
  CFD1QXL \s11.dbus_in_reg[0]  ( .D(n4322), .CP(n7741), .Q(\s11.dbus_in [0])
         );
  CFD1QXL \s12.Adr_reg[8]  ( .D(n4282), .CP(n7736), .Q(\s12.Adr [8]) );
  CFD1QXL \s12.Adr_reg[7]  ( .D(n4281), .CP(n7731), .Q(\s12.Adr [7]) );
  CFD1QXL \s12.Adr_reg[6]  ( .D(n4280), .CP(n7732), .Q(\s12.Adr [6]) );
  CFD1QXL \s12.Adr_reg[5]  ( .D(n4279), .CP(n7740), .Q(\s12.Adr [5]) );
  CFD1QXL \s12.Adr_reg[4]  ( .D(n4278), .CP(n7727), .Q(\s12.Adr [4]) );
  CFD1QXL \s12.Adr_reg[3]  ( .D(n4277), .CP(n7739), .Q(\s12.Adr [3]) );
  CFD1QXL \s12.Adr_reg[2]  ( .D(n4276), .CP(n7729), .Q(\s12.Adr [2]) );
  CFD1QXL \s12.Adr_reg[1]  ( .D(n4275), .CP(n7746), .Q(\s12.Adr [1]) );
  CFD1QXL \s12.Adr_reg[0]  ( .D(n4274), .CP(n7730), .Q(\s12.Adr [0]) );
  CFD1QXL \m06.DinMast_reg[15]  ( .D(n5201), .CP(n7740), .Q(\m06.DinMast [15])
         );
  CFD1QXL \m06.DinMast_reg[14]  ( .D(n5200), .CP(n7740), .Q(\m06.DinMast [14])
         );
  CFD1QXL \m06.DinMast_reg[13]  ( .D(n5199), .CP(n7740), .Q(\m06.DinMast [13])
         );
  CFD1QXL \m06.DinMast_reg[12]  ( .D(n5198), .CP(n7740), .Q(\m06.DinMast [12])
         );
  CFD1QXL \m06.DinMast_reg[11]  ( .D(n5197), .CP(n7740), .Q(\m06.DinMast [11])
         );
  CFD1QXL \m06.DinMast_reg[10]  ( .D(n5196), .CP(n7740), .Q(\m06.DinMast [10])
         );
  CFD1QXL \m06.DinMast_reg[9]  ( .D(n5195), .CP(n7740), .Q(\m06.DinMast [9])
         );
  CFD1QXL \m06.DinMast_reg[7]  ( .D(n5193), .CP(n7740), .Q(\m06.DinMast [7])
         );
  CFD1QXL \m06.DinMast_reg[6]  ( .D(n5192), .CP(n7733), .Q(\m06.DinMast [6])
         );
  CFD1QXL \m06.DinMast_reg[5]  ( .D(n5191), .CP(n7738), .Q(\m06.DinMast [5])
         );
  CFD1QXL \m06.DinMast_reg[4]  ( .D(n5190), .CP(n7739), .Q(\m06.DinMast [4])
         );
  CFD1QXL \m06.DinMast_reg[3]  ( .D(n5189), .CP(n7746), .Q(\m06.DinMast [3])
         );
  CFD1QXL \m06.DinMast_reg[2]  ( .D(n5188), .CP(n7741), .Q(\m06.DinMast [2])
         );
  CFD1QXL \m06.DinMast_reg[1]  ( .D(n5187), .CP(n7736), .Q(\m06.DinMast [1])
         );
  CFD1QXL \m06.DinMast_reg[0]  ( .D(n5186), .CP(n7731), .Q(\m06.DinMast [0])
         );
  CFD1QXL \m00.DinMast_reg[15]  ( .D(n5041), .CP(n7746), .Q(\m00.DinMast [15])
         );
  CFD1QXL \m00.DinMast_reg[14]  ( .D(n5040), .CP(n7741), .Q(\m00.DinMast [14])
         );
  CFD1QXL \m00.DinMast_reg[13]  ( .D(n5039), .CP(n7736), .Q(\m00.DinMast [13])
         );
  CFD1QXL \m00.DinMast_reg[12]  ( .D(n5038), .CP(n7736), .Q(\m00.DinMast [12])
         );
  CFD1QXL \m00.DinMast_reg[11]  ( .D(n5037), .CP(n7736), .Q(\m00.DinMast [11])
         );
  CFD1QXL \m00.DinMast_reg[10]  ( .D(n5036), .CP(n7736), .Q(\m00.DinMast [10])
         );
  CFD1QXL \m00.DinMast_reg[9]  ( .D(n5035), .CP(n7736), .Q(\m00.DinMast [9])
         );
  CFD1QXL \m00.DinMast_reg[8]  ( .D(n5034), .CP(n7732), .Q(\m00.DinMast [8])
         );
  CFD1QXL \m00.DinMast_reg[7]  ( .D(n5033), .CP(n7736), .Q(\m00.DinMast [7])
         );
  CFD1QXL \m00.DinMast_reg[6]  ( .D(n5032), .CP(n7736), .Q(\m00.DinMast [6])
         );
  CFD1QXL \m00.DinMast_reg[5]  ( .D(n5031), .CP(n7742), .Q(\m00.DinMast [5])
         );
  CFD1QXL \m00.DinMast_reg[4]  ( .D(n5030), .CP(n7736), .Q(\m00.DinMast [4])
         );
  CFD1QXL \m00.DinMast_reg[3]  ( .D(n5029), .CP(n7743), .Q(\m00.DinMast [3])
         );
  CFD1QXL \m00.DinMast_reg[2]  ( .D(n5028), .CP(n7736), .Q(\m00.DinMast [2])
         );
  CFD1QXL \m00.DinMast_reg[1]  ( .D(n5027), .CP(n7746), .Q(\m00.DinMast [1])
         );
  CFD1QXL \m00.DinMast_reg[0]  ( .D(n5026), .CP(n7741), .Q(\m00.DinMast [0])
         );
  CFD1QXL \m01.DinMast_reg[15]  ( .D(n4273), .CP(n7741), .Q(\m01.DinMast [15])
         );
  CFD1QXL \m01.DinMast_reg[14]  ( .D(n4272), .CP(n7735), .Q(\m01.DinMast [14])
         );
  CFD1QXL \m01.DinMast_reg[13]  ( .D(n4271), .CP(n7742), .Q(\m01.DinMast [13])
         );
  CFD1QXL \m01.DinMast_reg[12]  ( .D(n4270), .CP(n7736), .Q(\m01.DinMast [12])
         );
  CFD1QXL \m01.DinMast_reg[11]  ( .D(n4269), .CP(n7743), .Q(\m01.DinMast [11])
         );
  CFD1QXL \m01.DinMast_reg[10]  ( .D(n4268), .CP(n7731), .Q(\m01.DinMast [10])
         );
  CFD1QXL \m01.DinMast_reg[9]  ( .D(n4267), .CP(n7732), .Q(\m01.DinMast [9])
         );
  CFD1QXL \m01.DinMast_reg[8]  ( .D(n4266), .CP(n7740), .Q(\m01.DinMast [8])
         );
  CFD1QXL \m01.DinMast_reg[7]  ( .D(n4265), .CP(n7727), .Q(\m01.DinMast [7])
         );
  CFD1QXL \m01.DinMast_reg[6]  ( .D(n4264), .CP(n7728), .Q(\m01.DinMast [6])
         );
  CFD1QXL \m01.DinMast_reg[5]  ( .D(n4263), .CP(n7729), .Q(\m01.DinMast [5])
         );
  CFD1QXL \m01.DinMast_reg[4]  ( .D(n4262), .CP(n7744), .Q(\m01.DinMast [4])
         );
  CFD1QXL \m01.DinMast_reg[3]  ( .D(n4261), .CP(n7745), .Q(\m01.DinMast [3])
         );
  CFD1QXL \m01.DinMast_reg[2]  ( .D(n4260), .CP(n7730), .Q(\m01.DinMast [2])
         );
  CFD1QXL \m01.DinMast_reg[1]  ( .D(n4259), .CP(n7737), .Q(\m01.DinMast [1])
         );
  CFD1QXL \m01.DinMast_reg[0]  ( .D(n4258), .CP(n7734), .Q(\m01.DinMast [0])
         );
  CFD1QXL \m02.DinMast_reg[15]  ( .D(n4257), .CP(n7735), .Q(\m02.DinMast [15])
         );
  CFD1QXL \m02.DinMast_reg[14]  ( .D(n4256), .CP(n7733), .Q(\m02.DinMast [14])
         );
  CFD1QXL \m02.DinMast_reg[13]  ( .D(n4255), .CP(n7742), .Q(\m02.DinMast [13])
         );
  CFD1QXL \m02.DinMast_reg[12]  ( .D(n4254), .CP(n7743), .Q(\m02.DinMast [12])
         );
  CFD1QXL \m02.DinMast_reg[11]  ( .D(n4253), .CP(n7744), .Q(\m02.DinMast [11])
         );
  CFD1QXL \m02.DinMast_reg[10]  ( .D(n4252), .CP(n7738), .Q(\m02.DinMast [10])
         );
  CFD1QXL \m02.DinMast_reg[9]  ( .D(n4251), .CP(n7739), .Q(\m02.DinMast [9])
         );
  CFD1QXL \m02.DinMast_reg[8]  ( .D(n4250), .CP(n7746), .Q(\m02.DinMast [8])
         );
  CFD1QXL \m02.DinMast_reg[7]  ( .D(n4249), .CP(n7745), .Q(\m02.DinMast [7])
         );
  CFD1QXL \m02.DinMast_reg[6]  ( .D(n4248), .CP(n7737), .Q(\m02.DinMast [6])
         );
  CFD1QXL \m02.DinMast_reg[5]  ( .D(n4247), .CP(n7734), .Q(\m02.DinMast [5])
         );
  CFD1QXL \m02.DinMast_reg[4]  ( .D(n4246), .CP(n7741), .Q(\m02.DinMast [4])
         );
  CFD1QXL \m02.DinMast_reg[3]  ( .D(n4245), .CP(n7736), .Q(\m02.DinMast [3])
         );
  CFD1QXL \m02.DinMast_reg[2]  ( .D(n4244), .CP(n7733), .Q(\m02.DinMast [2])
         );
  CFD1QXL \m02.DinMast_reg[1]  ( .D(n4243), .CP(n7738), .Q(\m02.DinMast [1])
         );
  CFD1QXL \m02.DinMast_reg[0]  ( .D(n4242), .CP(n7731), .Q(\m02.DinMast [0])
         );
  CFD1QXL \m03.DinMast_reg[15]  ( .D(n4241), .CP(n7732), .Q(\m03.DinMast [15])
         );
  CFD1QXL \m03.DinMast_reg[14]  ( .D(n4240), .CP(n7739), .Q(\m03.DinMast [14])
         );
  CFD1QXL \m03.DinMast_reg[13]  ( .D(n4239), .CP(n7746), .Q(\m03.DinMast [13])
         );
  CFD1QXL \m03.DinMast_reg[12]  ( .D(n4238), .CP(n7740), .Q(\m03.DinMast [12])
         );
  CFD1QXL \m03.DinMast_reg[11]  ( .D(n4237), .CP(n7727), .Q(\m03.DinMast [11])
         );
  CFD1QXL \m03.DinMast_reg[10]  ( .D(n4236), .CP(n7741), .Q(\m03.DinMast [10])
         );
  CFD1QXL \m03.DinMast_reg[9]  ( .D(n4235), .CP(n7742), .Q(\m03.DinMast [9])
         );
  CFD1QXL \m03.DinMast_reg[8]  ( .D(n4234), .CP(n7743), .Q(\m03.DinMast [8])
         );
  CFD1QXL \m03.DinMast_reg[7]  ( .D(n4233), .CP(n7744), .Q(\m03.DinMast [7])
         );
  CFD1QXL \m03.DinMast_reg[6]  ( .D(n4232), .CP(n7745), .Q(\m03.DinMast [6])
         );
  CFD1QXL \m03.DinMast_reg[5]  ( .D(n4231), .CP(n7737), .Q(\m03.DinMast [5])
         );
  CFD1QXL \m03.DinMast_reg[4]  ( .D(n4230), .CP(n7726), .Q(\m03.DinMast [4])
         );
  CFD1QXL \m03.DinMast_reg[3]  ( .D(n4229), .CP(n7740), .Q(\m03.DinMast [3])
         );
  CFD1QXL \m03.DinMast_reg[2]  ( .D(n4228), .CP(n7734), .Q(\m03.DinMast [2])
         );
  CFD1QXL \m03.DinMast_reg[1]  ( .D(n4227), .CP(n7733), .Q(\m03.DinMast [1])
         );
  CFD1QXL \m03.DinMast_reg[0]  ( .D(n4226), .CP(n7738), .Q(\m03.DinMast [0])
         );
  CFD1QXL \m04.DinMast_reg[15]  ( .D(n4225), .CP(n7739), .Q(\m04.DinMast [15])
         );
  CFD1QXL \m04.DinMast_reg[14]  ( .D(n4224), .CP(n7746), .Q(\m04.DinMast [14])
         );
  CFD1QXL \m04.DinMast_reg[13]  ( .D(n4223), .CP(n7741), .Q(\m04.DinMast [13])
         );
  CFD1QXL \m04.DinMast_reg[12]  ( .D(n4222), .CP(n7726), .Q(\m04.DinMast [12])
         );
  CFD1QXL \m04.DinMast_reg[11]  ( .D(n4221), .CP(n7736), .Q(\m04.DinMast [11])
         );
  CFD1QXL \m04.DinMast_reg[10]  ( .D(n4220), .CP(n7731), .Q(\m04.DinMast [10])
         );
  CFD1QXL \m04.DinMast_reg[9]  ( .D(n4219), .CP(n7726), .Q(\m04.DinMast [9])
         );
  CFD1QXL \m04.DinMast_reg[8]  ( .D(n4218), .CP(n7732), .Q(\m04.DinMast [8])
         );
  CFD1QXL \m04.DinMast_reg[7]  ( .D(n4217), .CP(n7726), .Q(\m04.DinMast [7])
         );
  CFD1QXL \m04.DinMast_reg[6]  ( .D(n4216), .CP(n7726), .Q(\m04.DinMast [6])
         );
  CFD1QXL \m04.DinMast_reg[5]  ( .D(n4215), .CP(n7740), .Q(\m04.DinMast [5])
         );
  CFD1QXL \m04.DinMast_reg[4]  ( .D(n4214), .CP(n7726), .Q(\m04.DinMast [4])
         );
  CFD1QXL \m04.DinMast_reg[3]  ( .D(n4213), .CP(n7726), .Q(\m04.DinMast [3])
         );
  CFD1QXL \m04.DinMast_reg[2]  ( .D(n4212), .CP(n7726), .Q(\m04.DinMast [2])
         );
  CFD1QXL \m04.DinMast_reg[1]  ( .D(n4211), .CP(n7726), .Q(\m04.DinMast [1])
         );
  CFD1QXL \m04.DinMast_reg[0]  ( .D(n4210), .CP(n7726), .Q(\m04.DinMast [0])
         );
  CFD1QXL \m05.DinMast_reg[15]  ( .D(n4209), .CP(n7727), .Q(\m05.DinMast [15])
         );
  CFD1QXL \m05.DinMast_reg[14]  ( .D(n4208), .CP(n7728), .Q(\m05.DinMast [14])
         );
  CFD1QXL \m05.DinMast_reg[13]  ( .D(n4207), .CP(n7729), .Q(\m05.DinMast [13])
         );
  CFD1QXL \m05.DinMast_reg[12]  ( .D(n4206), .CP(n7730), .Q(\m05.DinMast [12])
         );
  CFD1QXL \m05.DinMast_reg[11]  ( .D(n4205), .CP(n7726), .Q(\m05.DinMast [11])
         );
  CFD1QXL \m05.DinMast_reg[10]  ( .D(n4204), .CP(n7735), .Q(\m05.DinMast [10])
         );
  CFD1QXL \m05.DinMast_reg[9]  ( .D(n4203), .CP(n7742), .Q(\m05.DinMast [9])
         );
  CFD1QXL \m05.DinMast_reg[8]  ( .D(n4202), .CP(n7743), .Q(\m05.DinMast [8])
         );
  CFD1QXL \m05.DinMast_reg[7]  ( .D(n4201), .CP(n7744), .Q(\m05.DinMast [7])
         );
  CFD1QXL \m05.DinMast_reg[6]  ( .D(n4200), .CP(n7726), .Q(\m05.DinMast [6])
         );
  CFD1QXL \m05.DinMast_reg[5]  ( .D(n4199), .CP(n7726), .Q(\m05.DinMast [5])
         );
  CFD1QXL \m05.DinMast_reg[4]  ( .D(n4198), .CP(n7726), .Q(\m05.DinMast [4])
         );
  CFD1QXL \m05.DinMast_reg[3]  ( .D(n4197), .CP(n7745), .Q(\m05.DinMast [3])
         );
  CFD1QXL \m05.DinMast_reg[2]  ( .D(n4196), .CP(n7726), .Q(\m05.DinMast [2])
         );
  CFD1QXL \m05.DinMast_reg[1]  ( .D(n4195), .CP(n7726), .Q(\m05.DinMast [1])
         );
  CFD1QXL \m05.DinMast_reg[0]  ( .D(n4194), .CP(n7726), .Q(\m05.DinMast [0])
         );
  CFD1QXL \s02.tarActive_reg  ( .D(n5212), .CP(n7740), .Q(\s02.tarActive ) );
  CFD1QXL \s00.Adr_reg[9]  ( .D(n5067), .CP(n7746), .Q(\s00.Adr [9]) );
  CFD1QXL \s13.tarActive_reg  ( .D(n5224), .CP(n7740), .Q(\s13.tarActive ) );
  CFD1QXL \s00.tarActive_reg  ( .D(n5214), .CP(n7740), .Q(\s00.tarActive ) );
  CFD1QXL \s01.tarActive_reg  ( .D(n5213), .CP(n7740), .Q(\s01.tarActive ) );
  CFD1QXL \s03.tarActive_reg  ( .D(n5211), .CP(n7740), .Q(\s03.tarActive ) );
  CFD1QXL \s04.tarActive_reg  ( .D(n5210), .CP(n7740), .Q(\s04.tarActive ) );
  CFD1QXL \s05.tarActive_reg  ( .D(n5209), .CP(n7740), .Q(\s05.tarActive ) );
  CFD1QXL \s06.tarActive_reg  ( .D(n5208), .CP(n7740), .Q(\s06.tarActive ) );
  CFD1QXL \s07.tarActive_reg  ( .D(n5207), .CP(n7732), .Q(\s07.tarActive ) );
  CFD1QXL \s08.tarActive_reg  ( .D(n5206), .CP(n7740), .Q(\s08.tarActive ) );
  CFD1QXL \s09.tarActive_reg  ( .D(n5205), .CP(n7727), .Q(\s09.tarActive ) );
  CFD1QXL \s10.tarActive_reg  ( .D(n5204), .CP(n7728), .Q(\s10.tarActive ) );
  CFD1QXL \s11.tarActive_reg  ( .D(n5203), .CP(n7729), .Q(\s11.tarActive ) );
  CFD1QXL \s12.tarActive_reg  ( .D(n5202), .CP(n7730), .Q(\s12.tarActive ) );
  CFD1QXL \m06.DinMast_reg[8]  ( .D(n5194), .CP(n7735), .Q(\m06.DinMast [8])
         );
  CFD1QXL \m02.YouGotIt_reg  ( .D(n5275), .CP(\clock.sysClk ), .Q(
        \m02.YouGotIt ) );
  CFD1QXL \m05.YouGotIt_reg  ( .D(n5245), .CP(n7740), .Q(\m05.YouGotIt ) );
  CFD1QXL \m06.YouGotIt_reg  ( .D(n5285), .CP(n7740), .Q(\m06.YouGotIt ) );
  CFD1QXL \m04.YouGotIt_reg  ( .D(n5235), .CP(n7740), .Q(\m04.YouGotIt ) );
  CFD1QXL \m01.YouGotIt_reg  ( .D(n5265), .CP(n7740), .Q(\m01.YouGotIt ) );
  CFD1QXL \m03.YouGotIt_reg  ( .D(n5255), .CP(n7740), .Q(\m03.YouGotIt ) );
  CFD1QX1 \m00.YouGotIt_reg  ( .D(n5225), .CP(\clock.sysClk ), .Q(
        \m00.YouGotIt ) );
  COR4X1 U5297 ( .A(n7185), .B(n7183), .C(n7553), .D(n7182), .Z(n6948) );
  COR4X1 U5298 ( .A(n7187), .B(n7186), .C(n7184), .D(n7180), .Z(n6947) );
  COR4X1 U5299 ( .A(n7532), .B(n7580), .C(n6789), .D(n6788), .Z(n5455) );
  COR8X1 U5300 ( .A(n7561), .B(\m01.addrM [45]), .C(\m01.addrM [46]), .D(
        \m01.addrM [47]), .E(\m01.addrM [41]), .F(\m01.addrM [42]), .G(
        \m01.addrM [43]), .H(\m01.addrM [44]), .Z(n5295) );
  COR4X1 U5301 ( .A(\m01.addrM [30]), .B(\m01.addrM [31]), .C(\m01.addrM [28]), 
        .D(\m01.addrM [29]), .Z(n5296) );
  COR4X1 U5302 ( .A(\m01.addrM [34]), .B(\m01.addrM [33]), .C(\m01.addrM [35]), 
        .D(n5296), .Z(n5297) );
  COR8X1 U5303 ( .A(\m01.addrM [37]), .B(\m01.addrM [38]), .C(\m01.addrM [39]), 
        .D(\m01.addrM [26]), .E(\m01.addrM [27]), .F(\m01.addrM [24]), .G(
        \m01.addrM [25]), .H(\m01.addrM [32]), .Z(n5298) );
  CNR4X1 U5304 ( .A(\m01.addrM [36]), .B(\m01.addrM [40]), .C(n5297), .D(n5298), .Z(n5299) );
  CND8X1 U5305 ( .A(\m01.addrM [17]), .B(\m01.addrM [20]), .C(\m01.addrM [19]), 
        .D(n5299), .E(\m01.addrM [21]), .F(\m01.addrM [23]), .G(
        \m01.addrM [22]), .H(\m01.addrM [18]), .Z(n5300) );
  CNR2X1 U5306 ( .A(n5295), .B(n5300), .Z(n7585) );
  CND3XL U5307 ( .A(n7531), .B(n6384), .C(n7515), .Z(n5301) );
  CND8X1 U5308 ( .A(n6558), .B(n6613), .C(n6601), .D(n6507), .E(n6325), .F(
        n7588), .G(n6503), .H(n7557), .Z(n5302) );
  CNR3XL U5309 ( .A(n6732), .B(n5301), .C(n5302), .Z(n5303) );
  CANR11X1 U5310 ( .A(n6664), .B(n6437), .C(n5303), .D(n7589), .Z(n6748) );
  COR8X1 U5311 ( .A(\m05.addrM [42]), .B(\m05.addrM [43]), .C(\m05.addrM [44]), 
        .D(\m05.addrM [45]), .E(\m05.addrM [38]), .F(\m05.addrM [39]), .G(
        \m05.addrM [40]), .H(\m05.addrM [41]), .Z(n5304) );
  CNR4X1 U5312 ( .A(\m05.addrM [33]), .B(\m05.addrM [30]), .C(\m05.addrM [27]), 
        .D(\m05.addrM [26]), .Z(n5305) );
  CAN4X1 U5313 ( .A(\m05.addrM [22]), .B(\m05.addrM [23]), .C(\m05.addrM [20]), 
        .D(\m05.addrM [17]), .Z(n5306) );
  CND4X1 U5314 ( .A(\m05.addrM [21]), .B(n5306), .C(\m05.addrM [18]), .D(
        \m05.addrM [19]), .Z(n5307) );
  CNR8X1 U5315 ( .A(n5307), .B(\m05.addrM [28]), .C(\m05.addrM [29]), .D(
        \m05.addrM [24]), .E(\m05.addrM [31]), .F(\m05.addrM [34]), .G(
        \m05.addrM [25]), .H(\m05.addrM [35]), .Z(n5308) );
  CND2X1 U5316 ( .A(n5305), .B(n5308), .Z(n5309) );
  COR8X1 U5317 ( .A(n5304), .B(n5309), .C(\m05.addrM [36]), .D(\m05.addrM [32]), .E(n6285), .F(\m05.addrM [46]), .G(\m05.addrM [47]), .H(\m05.addrM [37]), 
        .Z(n7589) );
  CIVX1 U5318 ( .A(n7300), .Z(n5310) );
  COR3X1 U5319 ( .A(\m03.addrM [2]), .B(\m03.addrM [0]), .C(n7299), .Z(n5311)
         );
  COND3X1 U5320 ( .A(n7318), .B(n7297), .C(n7298), .D(n5311), .Z(n5312) );
  CANR4CX1 U5321 ( .A(n7313), .B(n5310), .C(n7301), .D(n5312), .Z(n5313) );
  CND2X1 U5322 ( .A(\m03.addrM [14]), .B(\m03.addrM [13]), .Z(n5314) );
  CNR3XL U5323 ( .A(n7302), .B(n5313), .C(n5314), .Z(n5315) );
  CND3XL U5324 ( .A(\m03.addrM [15]), .B(\m03.addrM [16]), .C(n5315), .Z(n7484) );
  CND8X1 U5325 ( .A(n6677), .B(n7576), .C(n6332), .D(n6651), .E(n6392), .F(
        n6493), .G(n7514), .H(n6626), .Z(n5316) );
  CNR4XL U5326 ( .A(n7659), .B(n7667), .C(n6698), .D(n5316), .Z(n5317) );
  CAN4X1 U5327 ( .A(n6686), .B(n6579), .C(n6418), .D(n5317), .Z(n5318) );
  CNR2X1 U5328 ( .A(n7577), .B(n5318), .Z(n7679) );
  CAN3X1 U5329 ( .A(\m00.addrM [9]), .B(n5430), .C(n5371), .Z(n5376) );
  CIVX1 U5330 ( .A(n6849), .Z(n5319) );
  COND11X1 U5331 ( .A(n6483), .B(n6846), .C(n6828), .D(n6848), .Z(n5320) );
  COND1XL U5332 ( .A(\m04.addrM [5]), .B(n5320), .C(n6851), .Z(n5321) );
  CANR4CX1 U5333 ( .A(n6816), .B(n5319), .C(n5321), .D(n6854), .Z(n5322) );
  CAN2X1 U5334 ( .A(n6514), .B(n5322), .Z(n7243) );
  CND2X1 U5335 ( .A(n6634), .B(n6385), .Z(n5323) );
  COND1XL U5336 ( .A(\m03.addrM [0]), .B(n5323), .C(n7301), .Z(n5324) );
  CND2X1 U5337 ( .A(\m03.addrM [4]), .B(n6614), .Z(n5325) );
  CANR1XL U5338 ( .A(n6495), .B(n7296), .C(n7307), .Z(n5326) );
  COND4CX1 U5339 ( .A(n6633), .B(n5325), .C(n7298), .D(n5326), .Z(n5327) );
  CANR1XL U5340 ( .A(n6494), .B(n5324), .C(n5327), .Z(n5328) );
  CANR1XL U5341 ( .A(n7297), .B(n5328), .C(n6510), .Z(n5329) );
  CND2X1 U5342 ( .A(n7309), .B(n5329), .Z(n7436) );
  CAN4X1 U5343 ( .A(\m06.addrM [15]), .B(\m06.addrM [14]), .C(n6122), .D(n6093), .Z(n5330) );
  CND2IX1 U5344 ( .B(n6092), .A(\m06.addrM [3]), .Z(n5331) );
  COND1XL U5345 ( .A(n6149), .B(n6092), .C(n6127), .Z(n5332) );
  COND3X1 U5346 ( .A(n6156), .B(\m06.addrM [6]), .C(n6147), .D(n5332), .Z(
        n5333) );
  CANR11X1 U5347 ( .A(n6369), .B(n6138), .C(n6144), .D(n5333), .Z(n5334) );
  COND4CX1 U5348 ( .A(n6091), .B(n5331), .C(n6099), .D(n5334), .Z(n5335) );
  CND2X1 U5349 ( .A(n5330), .B(n5335), .Z(n7550) );
  CNR2IX1 U5350 ( .B(\m00.addrM [16]), .A(\m00.addrM [13]), .Z(n5361) );
  CIVX2 U5351 ( .A(\m00.addrM [14]), .Z(n5344) );
  CND2X1 U5352 ( .A(\m00.addrM [15]), .B(n5344), .Z(n5347) );
  CIVX2 U5353 ( .A(\m00.addrM [11]), .Z(n5378) );
  CNR3XL U5354 ( .A(\m00.addrM [12]), .B(n5347), .C(n5378), .Z(n5432) );
  CIVX2 U5355 ( .A(\m00.addrM [2]), .Z(n5397) );
  CND2X1 U5356 ( .A(\m00.addrM [4]), .B(\m00.addrM [3]), .Z(n5396) );
  CNR2X1 U5357 ( .A(n5397), .B(n5396), .Z(n5342) );
  CND2X1 U5358 ( .A(\m00.addrM [8]), .B(\m00.addrM [7]), .Z(n5390) );
  CIVX2 U5359 ( .A(n5390), .Z(n5365) );
  COND3X1 U5360 ( .A(\m00.addrM [5]), .B(n5342), .C(\m00.addrM [6]), .D(n5365), 
        .Z(n5339) );
  CNR2X1 U5361 ( .A(\m00.addrM [8]), .B(\m00.addrM [7]), .Z(n5399) );
  CIVX2 U5362 ( .A(\m00.addrM [8]), .Z(n5341) );
  CND2X1 U5363 ( .A(\m00.addrM [7]), .B(n5341), .Z(n5444) );
  CIVX2 U5364 ( .A(\m00.addrM [6]), .Z(n7563) );
  CNR2X1 U5365 ( .A(n5444), .B(n7563), .Z(n5385) );
  CIVX2 U5366 ( .A(\m00.addrM [5]), .Z(n5425) );
  CND2X1 U5367 ( .A(n5385), .B(n5425), .Z(n5422) );
  CNR3XL U5368 ( .A(\m00.addrM [0]), .B(\m00.addrM [1]), .C(n5422), .Z(n5337)
         );
  CANR4CX1 U5369 ( .A(\m00.addrM [5]), .B(n5342), .C(\m00.addrM [6]), .D(n5444), .Z(n5336) );
  COND11X1 U5370 ( .A(n5399), .B(n5337), .C(n5336), .D(\m00.addrM [9]), .Z(
        n5338) );
  CIVX2 U5371 ( .A(\m00.addrM [10]), .Z(n5430) );
  CANR4CX1 U5372 ( .A(\m00.addrM [9]), .B(n5339), .C(n5338), .D(n5430), .Z(
        n5340) );
  CND3XL U5373 ( .A(n5361), .B(n5432), .C(n5340), .Z(n6546) );
  CIVX2 U5374 ( .A(n6546), .Z(n6783) );
  CIVX2 U5375 ( .A(\m00.addrM [3]), .Z(n5381) );
  CND2X1 U5376 ( .A(n5397), .B(n5381), .Z(n5440) );
  CNR3XL U5377 ( .A(\m00.addrM [1]), .B(\m00.addrM [4]), .C(n5440), .Z(n5435)
         );
  CND2X1 U5378 ( .A(\m00.addrM [6]), .B(\m00.addrM [5]), .Z(n5429) );
  CNR2X1 U5379 ( .A(\m00.addrM [7]), .B(n5341), .Z(n5427) );
  CANR4CX1 U5380 ( .A(n5435), .B(n5429), .C(n5427), .D(n5385), .Z(n5346) );
  CNR2X1 U5381 ( .A(n5444), .B(n5425), .Z(n5343) );
  CNR2X1 U5382 ( .A(n5444), .B(n5425), .Z(n5384) );
  CIVX2 U5383 ( .A(\m00.addrM [1]), .Z(n5398) );
  CNR2X1 U5384 ( .A(n5398), .B(n5397), .Z(n5388) );
  CNR3XL U5385 ( .A(\m00.addrM [4]), .B(\m00.addrM [3]), .C(n5388), .Z(n5411)
         );
  CND2X1 U5386 ( .A(\m00.addrM [0]), .B(\m00.addrM [1]), .Z(n5382) );
  CNR2IX1 U5387 ( .B(n5342), .A(n5382), .Z(n5348) );
  CND3XL U5388 ( .A(\m00.addrM [0]), .B(\m00.addrM [2]), .C(n5398), .Z(n5352)
         );
  COND1XL U5389 ( .A(n5411), .B(n5348), .C(n5352), .Z(n5374) );
  CANR2X1 U5390 ( .A(\m00.addrM [4]), .B(n5343), .C(n5384), .D(n5374), .Z(
        n5345) );
  CAN2X1 U5391 ( .A(\m00.addrM [16]), .B(\m00.addrM [13]), .Z(n5431) );
  CIVX2 U5392 ( .A(\m00.addrM [15]), .Z(n5360) );
  CND3XL U5393 ( .A(n5431), .B(n5344), .C(n5360), .Z(n5443) );
  CNR2X1 U5394 ( .A(\m00.addrM [9]), .B(n5430), .Z(n5358) );
  CND3XL U5395 ( .A(\m00.addrM [12]), .B(\m00.addrM [11]), .C(n5358), .Z(n5408) );
  CANR3X1 U5396 ( .A(n5346), .B(n5345), .C(n5443), .D(n5408), .Z(n6782) );
  CANR2XL U5397 ( .A(n6783), .B(\s00.dataOut [0]), .C(n6782), .D(
        \s03.dataOut [0]), .Z(n5454) );
  CIVX2 U5398 ( .A(\m00.addrM [12]), .Z(n5379) );
  CNR2X1 U5399 ( .A(\m00.addrM [11]), .B(n5379), .Z(n5371) );
  CNR3XL U5400 ( .A(\m00.addrM [16]), .B(\m00.addrM [13]), .C(n5347), .Z(n5375) );
  CND3XL U5401 ( .A(\m00.addrM [6]), .B(n5427), .C(n5425), .Z(n5395) );
  COND3X1 U5402 ( .A(\m00.addrM [5]), .B(n5348), .C(n5427), .D(n7563), .Z(
        n5349) );
  COND4CX1 U5403 ( .A(\m00.addrM [4]), .B(n5440), .C(n5395), .D(n5349), .Z(
        n5350) );
  CAN4X1 U5404 ( .A(n5371), .B(n5358), .C(n5375), .D(n5350), .Z(n7580) );
  CND3XL U5405 ( .A(n5360), .B(\m00.addrM [14]), .C(n5431), .Z(n5416) );
  CIVX2 U5406 ( .A(n5416), .Z(n5359) );
  CNR2X1 U5407 ( .A(\m00.addrM [12]), .B(\m00.addrM [11]), .Z(n5357) );
  CIVX2 U5408 ( .A(n5388), .Z(n5351) );
  CIVX2 U5409 ( .A(\m00.addrM [4]), .Z(n5380) );
  CANR11X1 U5410 ( .A(n5352), .B(n5381), .C(n5351), .D(n5380), .Z(n5370) );
  CIVX2 U5411 ( .A(\m00.addrM [0]), .Z(n5403) );
  CNR2X1 U5412 ( .A(\m00.addrM [2]), .B(n5398), .Z(n5404) );
  CND3XL U5413 ( .A(\m00.addrM [4]), .B(n5404), .C(n5427), .Z(n5366) );
  CNR2IX1 U5414 ( .B(n5440), .A(n5380), .Z(n5353) );
  COND3X1 U5415 ( .A(\m00.addrM [5]), .B(n5353), .C(n7563), .D(n5427), .Z(
        n5368) );
  COND11X1 U5416 ( .A(n5403), .B(n5366), .C(\m00.addrM [6]), .D(n5368), .Z(
        n5354) );
  CIVX2 U5417 ( .A(n5354), .Z(n5355) );
  COND1XL U5418 ( .A(n5370), .B(n5395), .C(n5355), .Z(n5356) );
  CAN4X1 U5419 ( .A(n5359), .B(n5358), .C(n5357), .D(n5356), .Z(n6790) );
  CANR2X1 U5420 ( .A(\s04.dataOut [0]), .B(n7580), .C(\s10.dataOut [0]), .D(
        n6790), .Z(n5453) );
  CND3XL U5421 ( .A(\m00.addrM [14]), .B(n5361), .C(n5360), .Z(n5421) );
  CIVX2 U5422 ( .A(n5421), .Z(n5393) );
  CIVX2 U5423 ( .A(n5427), .Z(n5407) );
  CNR2X1 U5424 ( .A(n5429), .B(n5407), .Z(n5364) );
  CIVX2 U5425 ( .A(n5364), .Z(n5362) );
  COND2X1 U5426 ( .A(n5435), .B(n5395), .C(n5370), .D(n5362), .Z(n5363) );
  CND3XL U5427 ( .A(n5393), .B(n5376), .C(n5363), .Z(n5571) );
  CIVX2 U5428 ( .A(n5571), .Z(n7532) );
  CANR11X1 U5429 ( .A(\m00.addrM [1]), .B(\m00.addrM [2]), .C(\m00.addrM [3]), 
        .D(\m00.addrM [4]), .Z(n5420) );
  CANR4CX1 U5430 ( .A(n5429), .B(n5420), .C(n5365), .D(n5364), .Z(n5367) );
  CAN4X1 U5431 ( .A(n5368), .B(n5367), .C(n5366), .D(n5395), .Z(n5369) );
  CNR3X1 U5432 ( .A(n5369), .B(n5416), .C(n5408), .Z(n6784) );
  CANR2X1 U5433 ( .A(\s06.dataOut [0]), .B(n7532), .C(\s09.dataOut [0]), .D(
        n6784), .Z(n5452) );
  CND2X1 U5434 ( .A(n7563), .B(n5425), .Z(n5406) );
  COND1XL U5435 ( .A(n5370), .B(n5406), .C(n5399), .Z(n5373) );
  CNR2X1 U5436 ( .A(n5444), .B(n5406), .Z(n5387) );
  CND2X1 U5437 ( .A(n5411), .B(n5387), .Z(n5372) );
  CNR2X1 U5438 ( .A(\m00.addrM [10]), .B(\m00.addrM [9]), .Z(n5418) );
  CND2X1 U5439 ( .A(n5418), .B(n5371), .Z(n5442) );
  CANR3X1 U5440 ( .A(n5373), .B(n5372), .C(n5442), .D(n5416), .Z(n6797) );
  CNR2X1 U5441 ( .A(n5429), .B(n5390), .Z(n5377) );
  CAN4X1 U5442 ( .A(n5377), .B(n5376), .C(n5375), .D(n5374), .Z(n6789) );
  CND3XL U5443 ( .A(n5379), .B(n5378), .C(n5418), .Z(n5415) );
  CIVX2 U5444 ( .A(n5415), .Z(n5394) );
  COND4CX1 U5445 ( .A(n5397), .B(n5382), .C(n5381), .D(n5380), .Z(n5391) );
  CNR2X1 U5446 ( .A(n5444), .B(n5396), .Z(n5383) );
  COR4X1 U5447 ( .A(n5385), .B(n5384), .C(n5427), .D(n5383), .Z(n5386) );
  CANR11X1 U5448 ( .A(\m00.addrM [4]), .B(n5388), .C(n5387), .D(n5386), .Z(
        n5389) );
  COND11X1 U5449 ( .A(n5391), .B(n5390), .C(n5406), .D(n5389), .Z(n5392) );
  CND3XL U5450 ( .A(n5394), .B(n5393), .C(n5392), .Z(n6752) );
  CIVX2 U5451 ( .A(n6752), .Z(n6786) );
  CAOR2X2 U5452 ( .A(\s05.dataOut [0]), .B(n6789), .C(\s11.dataOut [0]), .D(
        n6786), .Z(n5450) );
  CIVX2 U5453 ( .A(\s07.dataOut [0]), .Z(n5448) );
  CIVX2 U5454 ( .A(n5395), .Z(n5405) );
  CANR1XL U5455 ( .A(n5398), .B(n5397), .C(n5396), .Z(n5424) );
  CND2X1 U5456 ( .A(n5427), .B(n5429), .Z(n5401) );
  CND2X1 U5457 ( .A(n5398), .B(n5397), .Z(n5400) );
  CNR2IX1 U5458 ( .B(n5399), .A(n5429), .Z(n5441) );
  COND4CX1 U5459 ( .A(\m00.addrM [3]), .B(n5400), .C(\m00.addrM [4]), .D(n5441), .Z(n5436) );
  COND4CX1 U5460 ( .A(n5424), .B(n5425), .C(n5401), .D(n5436), .Z(n5402) );
  CANR11X1 U5461 ( .A(n5405), .B(n5404), .C(n5403), .D(n5402), .Z(n5409) );
  CNR2X1 U5462 ( .A(n5407), .B(n5406), .Z(n5413) );
  CIVX2 U5463 ( .A(n5413), .Z(n5437) );
  CANR11X1 U5464 ( .A(n5409), .B(n5444), .C(n5437), .D(n5408), .Z(n5410) );
  CAN4X1 U5465 ( .A(\m00.addrM [14]), .B(\m00.addrM [15]), .C(n5431), .D(n5410), .Z(n6771) );
  CIVX2 U5466 ( .A(n6771), .Z(n7548) );
  CANR1XL U5467 ( .A(\m00.addrM [2]), .B(\m00.addrM [3]), .C(\m00.addrM [4]), 
        .Z(n5414) );
  CIVX2 U5468 ( .A(n5411), .Z(n5412) );
  CANR2X1 U5469 ( .A(n5414), .B(n5413), .C(n5441), .D(n5412), .Z(n5417) );
  CANR3X1 U5470 ( .A(n5417), .B(n5444), .C(n5416), .D(n5415), .Z(n6787) );
  CND3XL U5471 ( .A(\m00.addrM [12]), .B(\m00.addrM [11]), .C(n5418), .Z(n5419) );
  CNR4X1 U5472 ( .A(n5422), .B(n5421), .C(n5420), .D(n5419), .Z(n5423) );
  CNIVX1 U5473 ( .A(n5423), .Z(n6788) );
  CANR2XL U5474 ( .A(\s13.dataOut [0]), .B(n6787), .C(\s02.dataOut [0]), .D(
        n6788), .Z(n5447) );
  CIVX2 U5475 ( .A(n5424), .Z(n5428) );
  CANR3X1 U5476 ( .A(n5435), .B(n5425), .C(n5444), .D(n7563), .Z(n5426) );
  CANR4CX1 U5477 ( .A(n5429), .B(n5428), .C(n5427), .D(n5426), .Z(n5434) );
  CND4X1 U5478 ( .A(n5432), .B(\m00.addrM [9]), .C(n5431), .D(n5430), .Z(n5433) );
  CNR2X1 U5479 ( .A(n5434), .B(n5433), .Z(n6785) );
  CIVX2 U5480 ( .A(n5435), .Z(n5438) );
  COND11X1 U5481 ( .A(\m00.addrM [0]), .B(n5438), .C(n5437), .D(n5436), .Z(
        n5439) );
  CANR1XL U5482 ( .A(n5441), .B(n5440), .C(n5439), .Z(n5445) );
  CANR3X1 U5483 ( .A(n5445), .B(n5444), .C(n5443), .D(n5442), .Z(n6791) );
  CANR2XL U5484 ( .A(\s12.dataOut [0]), .B(n6785), .C(\s08.dataOut [0]), .D(
        n6791), .Z(n5446) );
  COND3X1 U5485 ( .A(n5448), .B(n7548), .C(n5447), .D(n5446), .Z(n5449) );
  CANR3XL U5486 ( .A(\s01.dataOut [0]), .B(n6797), .C(n5450), .D(n5449), .Z(
        n5451) );
  CND4X1 U5487 ( .A(n5454), .B(n5453), .C(n5452), .D(n5451), .Z(n5470) );
  CNR3XL U5488 ( .A(n6786), .B(n6784), .C(n6791), .Z(n5469) );
  CNR4XL U5489 ( .A(n6782), .B(n6797), .C(n6771), .D(n5455), .Z(n5456) );
  CIVX2 U5490 ( .A(n6785), .Z(n7522) );
  CIVX2 U5491 ( .A(n6787), .Z(n6506) );
  CAN4X1 U5492 ( .A(n5456), .B(n6546), .C(n7522), .D(n6506), .Z(n5468) );
  CIVX2 U5493 ( .A(n6790), .Z(n6774) );
  CAN4X1 U5494 ( .A(\m00.addrM [18]), .B(\m00.addrM [17]), .C(\m00.addrM [20]), 
        .D(\m00.addrM [19]), .Z(n5461) );
  CND3XL U5495 ( .A(\m00.addrM [21]), .B(\m00.addrM [22]), .C(\m00.addrM [23]), 
        .Z(n5457) );
  CNR2X1 U5496 ( .A(n5457), .B(\m00.addrM [39]), .Z(n5460) );
  CNR4X1 U5497 ( .A(\m00.addrM [44]), .B(\m00.addrM [45]), .C(\m00.addrM [46]), 
        .D(\m00.addrM [47]), .Z(n5459) );
  CNR4X1 U5498 ( .A(\m00.addrM [40]), .B(\m00.addrM [41]), .C(\m00.addrM [42]), 
        .D(\m00.addrM [43]), .Z(n5458) );
  CAN4X1 U5499 ( .A(n5461), .B(n5460), .C(n5459), .D(n5458), .Z(n5467) );
  CNR4X1 U5500 ( .A(\m00.addrM [27]), .B(\m00.addrM [28]), .C(\m00.addrM [29]), 
        .D(\m00.addrM [30]), .Z(n5465) );
  CIVXL U5501 ( .A(\m00.YouGotIt ), .Z(n7690) );
  CNR4X1 U5502 ( .A(\m00.addrM [25]), .B(\m00.addrM [24]), .C(\m00.addrM [26]), 
        .D(n7690), .Z(n5464) );
  CNR4X1 U5503 ( .A(\m00.addrM [35]), .B(\m00.addrM [36]), .C(\m00.addrM [37]), 
        .D(\m00.addrM [38]), .Z(n5463) );
  CNR4X1 U5504 ( .A(\m00.addrM [31]), .B(\m00.addrM [32]), .C(\m00.addrM [33]), 
        .D(\m00.addrM [34]), .Z(n5462) );
  CAN4X1 U5505 ( .A(n5465), .B(n5464), .C(n5463), .D(n5462), .Z(n5466) );
  CND2X1 U5506 ( .A(n5467), .B(n5466), .Z(n7549) );
  CANR11X1 U5507 ( .A(n5469), .B(n5468), .C(n6774), .D(n7549), .Z(n6802) );
  CMX2XL U5508 ( .A0(\m00.DinMast [0]), .A1(n5470), .S(n6802), .Z(n5026) );
  CANR2XL U5509 ( .A(n6783), .B(\s00.dataOut [1]), .C(\s01.dataOut [1]), .D(
        n6797), .Z(n5478) );
  CANR2XL U5510 ( .A(\s12.dataOut [1]), .B(n6785), .C(\s08.dataOut [1]), .D(
        n6791), .Z(n5477) );
  CANR2X1 U5511 ( .A(\s04.dataOut [1]), .B(n7580), .C(\s06.dataOut [1]), .D(
        n7532), .Z(n5476) );
  CAOR2XL U5512 ( .A(n6782), .B(\s03.dataOut [1]), .C(\s11.dataOut [1]), .D(
        n6786), .Z(n5474) );
  CIVX2 U5513 ( .A(\s07.dataOut [1]), .Z(n7343) );
  CANR2XL U5514 ( .A(\s13.dataOut [1]), .B(n6787), .C(\s02.dataOut [1]), .D(
        n6788), .Z(n5472) );
  CANR2X1 U5515 ( .A(\s10.dataOut [1]), .B(n6790), .C(\s09.dataOut [1]), .D(
        n6784), .Z(n5471) );
  COND3X1 U5516 ( .A(n7343), .B(n7548), .C(n5472), .D(n5471), .Z(n5473) );
  CANR3X1 U5517 ( .A(\s05.dataOut [1]), .B(n6789), .C(n5474), .D(n5473), .Z(
        n5475) );
  CND4X1 U5518 ( .A(n5478), .B(n5477), .C(n5476), .D(n5475), .Z(n5479) );
  CMX2XL U5519 ( .A0(\m00.DinMast [1]), .A1(n5479), .S(n6802), .Z(n5027) );
  CANR2XL U5520 ( .A(n6783), .B(\s00.dataOut [2]), .C(n6782), .D(
        \s03.dataOut [2]), .Z(n5487) );
  CANR2XL U5521 ( .A(\s07.dataOut [2]), .B(n6771), .C(\s08.dataOut [2]), .D(
        n6791), .Z(n5486) );
  CANR2X1 U5522 ( .A(\s12.dataOut [2]), .B(n6785), .C(\s04.dataOut [2]), .D(
        n7580), .Z(n5485) );
  CAOR2XL U5523 ( .A(\s13.dataOut [2]), .B(n6787), .C(\s11.dataOut [2]), .D(
        n6786), .Z(n5483) );
  CIVX2 U5524 ( .A(\s10.dataOut [2]), .Z(n6244) );
  CANR2XL U5525 ( .A(\s05.dataOut [2]), .B(n6789), .C(\s02.dataOut [2]), .D(
        n6788), .Z(n5481) );
  CANR2X1 U5526 ( .A(\s06.dataOut [2]), .B(n7532), .C(\s09.dataOut [2]), .D(
        n6784), .Z(n5480) );
  COND3X1 U5527 ( .A(n6244), .B(n6774), .C(n5481), .D(n5480), .Z(n5482) );
  CANR3XL U5528 ( .A(\s01.dataOut [2]), .B(n6797), .C(n5483), .D(n5482), .Z(
        n5484) );
  CND4X1 U5529 ( .A(n5487), .B(n5486), .C(n5485), .D(n5484), .Z(n5488) );
  CMX2XL U5530 ( .A0(\m00.DinMast [2]), .A1(n5488), .S(n6802), .Z(n5028) );
  CANR2XL U5531 ( .A(n6783), .B(\s00.dataOut [3]), .C(n6782), .D(
        \s03.dataOut [3]), .Z(n5497) );
  CANR2XL U5532 ( .A(\s08.dataOut [3]), .B(n6791), .C(\s09.dataOut [3]), .D(
        n6784), .Z(n5496) );
  CANR2X1 U5533 ( .A(\s12.dataOut [3]), .B(n6785), .C(\s10.dataOut [3]), .D(
        n6790), .Z(n5495) );
  CAOR2X2 U5534 ( .A(\s05.dataOut [3]), .B(n6789), .C(\s06.dataOut [3]), .D(
        n7532), .Z(n5493) );
  CIVX2 U5535 ( .A(\s11.dataOut [3]), .Z(n5491) );
  CANR2XL U5536 ( .A(\s02.dataOut [3]), .B(n6788), .C(\s13.dataOut [3]), .D(
        n6787), .Z(n5490) );
  CANR2X1 U5537 ( .A(\s07.dataOut [3]), .B(n6771), .C(\s04.dataOut [3]), .D(
        n7580), .Z(n5489) );
  COND3X1 U5538 ( .A(n5491), .B(n6752), .C(n5490), .D(n5489), .Z(n5492) );
  CANR3XL U5539 ( .A(\s01.dataOut [3]), .B(n6797), .C(n5493), .D(n5492), .Z(
        n5494) );
  CND4X1 U5540 ( .A(n5497), .B(n5496), .C(n5495), .D(n5494), .Z(n5498) );
  CMX2XL U5541 ( .A0(\m00.DinMast [3]), .A1(n5498), .S(n6802), .Z(n5029) );
  CANR2XL U5542 ( .A(n6783), .B(\s00.dataOut [4]), .C(\s01.dataOut [4]), .D(
        n6797), .Z(n5507) );
  CANR2X1 U5543 ( .A(\s04.dataOut [4]), .B(n7580), .C(\s10.dataOut [4]), .D(
        n6790), .Z(n5506) );
  CANR2XL U5544 ( .A(\s06.dataOut [4]), .B(n7532), .C(\s08.dataOut [4]), .D(
        n6791), .Z(n5505) );
  CAOR2X2 U5545 ( .A(\s05.dataOut [4]), .B(n6789), .C(\s12.dataOut [4]), .D(
        n6785), .Z(n5503) );
  CIVX2 U5546 ( .A(\s09.dataOut [4]), .Z(n5501) );
  CIVX2 U5547 ( .A(n6784), .Z(n5540) );
  CANR2XL U5548 ( .A(\s13.dataOut [4]), .B(n6787), .C(\s02.dataOut [4]), .D(
        n6788), .Z(n5500) );
  CANR2X1 U5549 ( .A(\s07.dataOut [4]), .B(n6771), .C(\s11.dataOut [4]), .D(
        n6786), .Z(n5499) );
  COND3X1 U5550 ( .A(n5501), .B(n5540), .C(n5500), .D(n5499), .Z(n5502) );
  CANR3XL U5551 ( .A(n6782), .B(\s03.dataOut [4]), .C(n5503), .D(n5502), .Z(
        n5504) );
  CND4X1 U5552 ( .A(n5507), .B(n5506), .C(n5505), .D(n5504), .Z(n5508) );
  CMX2XL U5553 ( .A0(\m00.DinMast [4]), .A1(n5508), .S(n6802), .Z(n5030) );
  CANR2XL U5554 ( .A(n6783), .B(\s00.dataOut [5]), .C(\s01.dataOut [5]), .D(
        n6797), .Z(n5516) );
  CANR2X1 U5555 ( .A(\s07.dataOut [5]), .B(n6771), .C(\s04.dataOut [5]), .D(
        n7580), .Z(n5515) );
  CANR2X1 U5556 ( .A(\s06.dataOut [5]), .B(n7532), .C(\s09.dataOut [5]), .D(
        n6784), .Z(n5514) );
  CAOR2XL U5557 ( .A(\s05.dataOut [5]), .B(n6789), .C(\s08.dataOut [5]), .D(
        n6791), .Z(n5512) );
  CIVX2 U5558 ( .A(\s11.dataOut [5]), .Z(n7384) );
  CANR2XL U5559 ( .A(\s13.dataOut [5]), .B(n6787), .C(\s02.dataOut [5]), .D(
        n6788), .Z(n5510) );
  CANR2X1 U5560 ( .A(\s12.dataOut [5]), .B(n6785), .C(\s10.dataOut [5]), .D(
        n6790), .Z(n5509) );
  COND3X1 U5561 ( .A(n7384), .B(n6752), .C(n5510), .D(n5509), .Z(n5511) );
  CANR3XL U5562 ( .A(n6782), .B(\s03.dataOut [5]), .C(n5512), .D(n5511), .Z(
        n5513) );
  CND4X1 U5563 ( .A(n5516), .B(n5515), .C(n5514), .D(n5513), .Z(n5517) );
  CMX2XL U5564 ( .A0(\m00.DinMast [5]), .A1(n5517), .S(n6802), .Z(n5031) );
  CANR2XL U5565 ( .A(n6783), .B(\s00.dataOut [6]), .C(n6782), .D(
        \s03.dataOut [6]), .Z(n5526) );
  CANR2X1 U5566 ( .A(\s07.dataOut [6]), .B(n6771), .C(\s11.dataOut [6]), .D(
        n6786), .Z(n5525) );
  CANR2X1 U5567 ( .A(\s06.dataOut [6]), .B(n7532), .C(\s04.dataOut [6]), .D(
        n7580), .Z(n5524) );
  CAOR2X2 U5568 ( .A(\s12.dataOut [6]), .B(n6785), .C(\s13.dataOut [6]), .D(
        n6787), .Z(n5522) );
  CIVX2 U5569 ( .A(\s09.dataOut [6]), .Z(n5520) );
  CANR2XL U5570 ( .A(\s05.dataOut [6]), .B(n6789), .C(\s02.dataOut [6]), .D(
        n6788), .Z(n5519) );
  CANR2XL U5571 ( .A(\s10.dataOut [6]), .B(n6790), .C(\s08.dataOut [6]), .D(
        n6791), .Z(n5518) );
  COND3X1 U5572 ( .A(n5520), .B(n5540), .C(n5519), .D(n5518), .Z(n5521) );
  CANR3XL U5573 ( .A(\s01.dataOut [6]), .B(n6797), .C(n5522), .D(n5521), .Z(
        n5523) );
  CND4X1 U5574 ( .A(n5526), .B(n5525), .C(n5524), .D(n5523), .Z(n5527) );
  CMX2XL U5575 ( .A0(\m00.DinMast [6]), .A1(n5527), .S(n6802), .Z(n5032) );
  CANR2XL U5576 ( .A(n6783), .B(\s00.dataOut [7]), .C(\s01.dataOut [7]), .D(
        n6797), .Z(n5536) );
  CANR2XL U5577 ( .A(\s08.dataOut [7]), .B(n6791), .C(\s11.dataOut [7]), .D(
        n6786), .Z(n5535) );
  CANR2X1 U5578 ( .A(\s06.dataOut [7]), .B(n7532), .C(\s07.dataOut [7]), .D(
        n6771), .Z(n5534) );
  CIVX2 U5579 ( .A(\s13.dataOut [7]), .Z(n6687) );
  CIVX2 U5580 ( .A(\s10.dataOut [7]), .Z(n6676) );
  COND2X1 U5581 ( .A(n6687), .B(n6506), .C(n6676), .D(n6774), .Z(n5532) );
  CIVX2 U5582 ( .A(\s09.dataOut [7]), .Z(n5530) );
  CANR2XL U5583 ( .A(\s05.dataOut [7]), .B(n6789), .C(\s02.dataOut [7]), .D(
        n6788), .Z(n5529) );
  CANR2X1 U5584 ( .A(\s04.dataOut [7]), .B(n7580), .C(\s12.dataOut [7]), .D(
        n6785), .Z(n5528) );
  COND3X1 U5585 ( .A(n5530), .B(n5540), .C(n5529), .D(n5528), .Z(n5531) );
  CANR3XL U5586 ( .A(n6782), .B(\s03.dataOut [7]), .C(n5532), .D(n5531), .Z(
        n5533) );
  CND4X1 U5587 ( .A(n5536), .B(n5535), .C(n5534), .D(n5533), .Z(n5537) );
  CMX2XL U5588 ( .A0(\m00.DinMast [7]), .A1(n5537), .S(n6802), .Z(n5033) );
  CANR2XL U5589 ( .A(n6783), .B(\s00.dataOut [8]), .C(\s01.dataOut [8]), .D(
        n6797), .Z(n5547) );
  CANR2X1 U5590 ( .A(\s06.dataOut [8]), .B(n7532), .C(\s11.dataOut [8]), .D(
        n6786), .Z(n5546) );
  CANR2X1 U5591 ( .A(\s04.dataOut [8]), .B(n7580), .C(\s10.dataOut [8]), .D(
        n6790), .Z(n5545) );
  CAOR2X2 U5592 ( .A(\s07.dataOut [8]), .B(n6771), .C(\s13.dataOut [8]), .D(
        n6787), .Z(n5543) );
  CIVX2 U5593 ( .A(\s09.dataOut [8]), .Z(n5541) );
  CANR2XL U5594 ( .A(\s05.dataOut [8]), .B(n6789), .C(\s02.dataOut [8]), .D(
        n6788), .Z(n5539) );
  CANR2XL U5595 ( .A(\s12.dataOut [8]), .B(n6785), .C(\s08.dataOut [8]), .D(
        n6791), .Z(n5538) );
  COND3X1 U5596 ( .A(n5541), .B(n5540), .C(n5539), .D(n5538), .Z(n5542) );
  CANR3XL U5597 ( .A(n6782), .B(\s03.dataOut [8]), .C(n5543), .D(n5542), .Z(
        n5544) );
  CND4X1 U5598 ( .A(n5547), .B(n5546), .C(n5545), .D(n5544), .Z(n5548) );
  CMX2XL U5599 ( .A0(\m00.DinMast [8]), .A1(n5548), .S(n6802), .Z(n5034) );
  CANR2XL U5600 ( .A(n6783), .B(\s00.dataOut [9]), .C(\s01.dataOut [9]), .D(
        n6797), .Z(n5557) );
  CANR2X1 U5601 ( .A(\s12.dataOut [9]), .B(n6785), .C(\s04.dataOut [9]), .D(
        n7580), .Z(n5556) );
  CANR2X1 U5602 ( .A(\s07.dataOut [9]), .B(n6771), .C(\s11.dataOut [9]), .D(
        n6786), .Z(n5555) );
  CAOR2X2 U5603 ( .A(\s05.dataOut [9]), .B(n6789), .C(\s09.dataOut [9]), .D(
        n6784), .Z(n5553) );
  CIVX2 U5604 ( .A(\s10.dataOut [9]), .Z(n5551) );
  CANR2XL U5605 ( .A(\s02.dataOut [9]), .B(n6788), .C(\s13.dataOut [9]), .D(
        n6787), .Z(n5550) );
  CANR2XL U5606 ( .A(\s06.dataOut [9]), .B(n7532), .C(\s08.dataOut [9]), .D(
        n6791), .Z(n5549) );
  COND3X1 U5607 ( .A(n5551), .B(n6774), .C(n5550), .D(n5549), .Z(n5552) );
  CANR3XL U5608 ( .A(n6782), .B(\s03.dataOut [9]), .C(n5553), .D(n5552), .Z(
        n5554) );
  CND4X1 U5609 ( .A(n5557), .B(n5556), .C(n5555), .D(n5554), .Z(n5558) );
  CMX2XL U5610 ( .A0(\m00.DinMast [9]), .A1(n5558), .S(n6802), .Z(n5035) );
  CANR2XL U5611 ( .A(n6783), .B(\s00.dataOut [10]), .C(\s01.dataOut [10]), .D(
        n6797), .Z(n5567) );
  CANR2X1 U5612 ( .A(\s07.dataOut [10]), .B(n6771), .C(\s12.dataOut [10]), .D(
        n6785), .Z(n5566) );
  CANR2X1 U5613 ( .A(\s06.dataOut [10]), .B(n7532), .C(\s11.dataOut [10]), .D(
        n6786), .Z(n5565) );
  CAOR2X2 U5614 ( .A(\s05.dataOut [10]), .B(n6789), .C(\s10.dataOut [10]), .D(
        n6790), .Z(n5563) );
  CIVX2 U5615 ( .A(\s04.dataOut [10]), .Z(n7448) );
  CIVX2 U5616 ( .A(n7580), .Z(n5561) );
  CANR2XL U5617 ( .A(\s02.dataOut [10]), .B(n6788), .C(\s13.dataOut [10]), .D(
        n6787), .Z(n5560) );
  CANR2XL U5618 ( .A(\s09.dataOut [10]), .B(n6784), .C(\s08.dataOut [10]), .D(
        n6791), .Z(n5559) );
  COND3X1 U5619 ( .A(n7448), .B(n5561), .C(n5560), .D(n5559), .Z(n5562) );
  CANR3XL U5620 ( .A(n6782), .B(\s03.dataOut [10]), .C(n5563), .D(n5562), .Z(
        n5564) );
  CND4X1 U5621 ( .A(n5567), .B(n5566), .C(n5565), .D(n5564), .Z(n5568) );
  CMX2XL U5622 ( .A0(\m00.DinMast [10]), .A1(n5568), .S(n6802), .Z(n5036) );
  CANR2X1 U5623 ( .A(n6783), .B(\s00.dataOut [11]), .C(\s01.dataOut [11]), .D(
        n6797), .Z(n5578) );
  CANR2XL U5624 ( .A(\s11.dataOut [11]), .B(n6786), .C(\s08.dataOut [11]), .D(
        n6791), .Z(n5577) );
  CANR2X1 U5625 ( .A(\s07.dataOut [11]), .B(n6771), .C(\s09.dataOut [11]), .D(
        n6784), .Z(n5576) );
  CAOR2X2 U5626 ( .A(\s05.dataOut [11]), .B(n6789), .C(\s10.dataOut [11]), .D(
        n6790), .Z(n5574) );
  CIVX2 U5627 ( .A(\s06.dataOut [11]), .Z(n5572) );
  CANR2XL U5628 ( .A(\s13.dataOut [11]), .B(n6787), .C(\s02.dataOut [11]), .D(
        n6788), .Z(n5570) );
  CANR2X1 U5629 ( .A(\s12.dataOut [11]), .B(n6785), .C(\s04.dataOut [11]), .D(
        n7580), .Z(n5569) );
  COND3X1 U5630 ( .A(n5572), .B(n5571), .C(n5570), .D(n5569), .Z(n5573) );
  CANR3XL U5631 ( .A(n6782), .B(\s03.dataOut [11]), .C(n5574), .D(n5573), .Z(
        n5575) );
  CND4X1 U5632 ( .A(n5578), .B(n5577), .C(n5576), .D(n5575), .Z(n5579) );
  CMX2XL U5633 ( .A0(\m00.DinMast [11]), .A1(n5579), .S(n6802), .Z(n5037) );
  CND2X1 U5634 ( .A(\m02.addrM [7]), .B(\m02.addrM [8]), .Z(n5689) );
  CIVX2 U5635 ( .A(\m02.addrM [2]), .Z(n5637) );
  CND2X1 U5636 ( .A(\m02.addrM [4]), .B(\m02.addrM [3]), .Z(n5634) );
  CNR2X1 U5637 ( .A(n5637), .B(n5634), .Z(n5605) );
  CIVX2 U5638 ( .A(\m02.addrM [10]), .Z(n5651) );
  CNR2X1 U5639 ( .A(\m02.addrM [9]), .B(n5651), .Z(n5622) );
  COND3X1 U5640 ( .A(\m02.addrM [5]), .B(n5605), .C(\m02.addrM [6]), .D(n5622), 
        .Z(n5584) );
  CIVX2 U5641 ( .A(\m02.addrM [7]), .Z(n7542) );
  CNR2X1 U5642 ( .A(n7542), .B(\m02.addrM [8]), .Z(n5683) );
  CIVX2 U5643 ( .A(n5683), .Z(n5639) );
  CANR4CX1 U5644 ( .A(\m02.addrM [5]), .B(n5605), .C(\m02.addrM [6]), .D(n5639), .Z(n5581) );
  CIVX2 U5645 ( .A(\m02.addrM [1]), .Z(n5585) );
  CND2X1 U5646 ( .A(\m02.addrM [2]), .B(n5585), .Z(n5610) );
  CIVX2 U5647 ( .A(\m02.addrM [6]), .Z(n7565) );
  CNR2X1 U5648 ( .A(n7565), .B(n5639), .Z(n5645) );
  CIVX2 U5649 ( .A(\m02.addrM [5]), .Z(n5621) );
  CND2X1 U5650 ( .A(n5645), .B(n5621), .Z(n5656) );
  COR2X1 U5651 ( .A(\m02.addrM [8]), .B(\m02.addrM [7]), .Z(n5666) );
  COND11X1 U5652 ( .A(\m02.addrM [0]), .B(n5610), .C(n5656), .D(n5666), .Z(
        n5580) );
  COND3X1 U5653 ( .A(n5581), .B(n5580), .C(\m02.addrM [10]), .D(\m02.addrM [9]), .Z(n5583) );
  CNR2X1 U5654 ( .A(\m02.addrM [13]), .B(\m02.addrM [14]), .Z(n5604) );
  CIVX2 U5655 ( .A(\m02.addrM [12]), .Z(n5600) );
  CAN4X1 U5656 ( .A(\m02.addrM [11]), .B(\m02.addrM [15]), .C(\m02.addrM [16]), 
        .D(n5600), .Z(n5653) );
  CND2X1 U5657 ( .A(n5604), .B(n5653), .Z(n5582) );
  CANR4CX1 U5658 ( .A(n5689), .B(n5584), .C(n5583), .D(n5582), .Z(n7265) );
  CNR2X1 U5659 ( .A(n5585), .B(n5637), .Z(n5663) );
  CNR2X1 U5660 ( .A(\m02.addrM [4]), .B(n5663), .Z(n5589) );
  CIVX2 U5661 ( .A(n5589), .Z(n5586) );
  CND2X1 U5662 ( .A(n5585), .B(n5637), .Z(n5635) );
  CND2X1 U5663 ( .A(\m02.addrM [3]), .B(n5635), .Z(n5587) );
  CNR2X1 U5664 ( .A(n5586), .B(n5587), .Z(n5698) );
  CNR2X1 U5665 ( .A(\m02.addrM [3]), .B(n5586), .Z(n5628) );
  CIVX2 U5666 ( .A(\m02.addrM [4]), .Z(n5619) );
  CND2X1 U5667 ( .A(n5619), .B(n5587), .Z(n5690) );
  CIVX2 U5668 ( .A(\m02.addrM [0]), .Z(n5674) );
  COND2X1 U5669 ( .A(n5628), .B(n5690), .C(n5674), .D(n5610), .Z(n5607) );
  CNR2X1 U5670 ( .A(n5639), .B(n5621), .Z(n5592) );
  CND2X1 U5671 ( .A(\m02.addrM [6]), .B(\m02.addrM [5]), .Z(n5606) );
  CND2X1 U5672 ( .A(\m02.addrM [8]), .B(n7542), .Z(n5692) );
  CNR2X1 U5673 ( .A(n5606), .B(n5692), .Z(n5682) );
  CNR2X1 U5674 ( .A(\m02.addrM [3]), .B(n5635), .Z(n5695) );
  CIVX2 U5675 ( .A(n5692), .Z(n5593) );
  CND2X1 U5676 ( .A(n5593), .B(n7565), .Z(n5677) );
  CNR2X1 U5677 ( .A(\m02.addrM [5]), .B(n5677), .Z(n5691) );
  CANR3X1 U5678 ( .A(n5682), .B(n5695), .C(n5645), .D(n5691), .Z(n5590) );
  CNR2X1 U5679 ( .A(\m02.addrM [6]), .B(\m02.addrM [5]), .Z(n5693) );
  CNR2X1 U5680 ( .A(n5693), .B(n5639), .Z(n5588) );
  CNR2X1 U5681 ( .A(n5588), .B(n5691), .Z(n5688) );
  CNR2X1 U5682 ( .A(\m02.addrM [4]), .B(\m02.addrM [3]), .Z(n5670) );
  CNR2X1 U5683 ( .A(n5589), .B(n5670), .Z(n5596) );
  CMXI2X1 U5684 ( .A0(n5590), .A1(n5688), .S(n5596), .Z(n5591) );
  CANR4CX1 U5685 ( .A(n5698), .B(n5607), .C(n5592), .D(n5591), .Z(n5594) );
  CNR2IX1 U5686 ( .B(n5606), .A(n5693), .Z(n5647) );
  CND2X1 U5687 ( .A(n5593), .B(n5647), .Z(n5646) );
  CIVX2 U5688 ( .A(\m02.addrM [16]), .Z(n5603) );
  CNR2X1 U5689 ( .A(\m02.addrM [15]), .B(n5603), .Z(n5609) );
  CIVX2 U5690 ( .A(\m02.addrM [13]), .Z(n5595) );
  CNR2X1 U5691 ( .A(\m02.addrM [14]), .B(n5595), .Z(n5652) );
  CND2X1 U5692 ( .A(n5609), .B(n5652), .Z(n5601) );
  CND3XL U5693 ( .A(\m02.addrM [11]), .B(\m02.addrM [12]), .C(n5622), .Z(n5700) );
  CANR3X1 U5694 ( .A(n5594), .B(n5646), .C(n5601), .D(n5700), .Z(n7264) );
  CANR2XL U5695 ( .A(n7265), .B(\s00.dataOut [0]), .C(n7264), .D(
        \s03.dataOut [0]), .Z(n5710) );
  CND3XL U5696 ( .A(\m02.addrM [14]), .B(n5609), .C(n5595), .Z(n5685) );
  CNR2X1 U5697 ( .A(\m02.addrM [9]), .B(\m02.addrM [10]), .Z(n5631) );
  CND4X1 U5698 ( .A(\m02.addrM [11]), .B(\m02.addrM [12]), .C(n5596), .D(n5631), .Z(n5597) );
  CNR3X1 U5699 ( .A(n5656), .B(n5685), .C(n5597), .Z(n7267) );
  CND2X1 U5700 ( .A(n5670), .B(n5637), .Z(n5598) );
  CNR2X1 U5701 ( .A(\m02.addrM [1]), .B(n5598), .Z(n5657) );
  CIVX2 U5702 ( .A(n5657), .Z(n5658) );
  CNR2X1 U5703 ( .A(\m02.addrM [0]), .B(n5658), .Z(n5599) );
  CNR2X1 U5704 ( .A(n5666), .B(n5606), .Z(n5636) );
  CANR2X1 U5705 ( .A(n5691), .B(n5599), .C(n5636), .D(n5598), .Z(n5602) );
  CNR2X1 U5706 ( .A(n5600), .B(\m02.addrM [11]), .Z(n5617) );
  CND2X1 U5707 ( .A(n5617), .B(n5631), .Z(n5671) );
  CANR3X1 U5708 ( .A(n5602), .B(n5639), .C(n5601), .D(n5671), .Z(n7266) );
  CANR2XL U5709 ( .A(\s02.dataOut [0]), .B(n7267), .C(\s08.dataOut [0]), .D(
        n7266), .Z(n5709) );
  CND3XL U5710 ( .A(\m02.addrM [9]), .B(n5617), .C(n5651), .Z(n5661) );
  CND3XL U5711 ( .A(\m02.addrM [15]), .B(n5604), .C(n5603), .Z(n5626) );
  CND3XL U5712 ( .A(\m02.addrM [0]), .B(\m02.addrM [1]), .C(n5605), .Z(n5618)
         );
  CNR2X1 U5713 ( .A(n5606), .B(n5689), .Z(n5699) );
  COND4CX1 U5714 ( .A(n5690), .B(n5618), .C(n5607), .D(n5699), .Z(n5608) );
  CNR3X1 U5715 ( .A(n5661), .B(n5626), .C(n5608), .Z(n7269) );
  CND3XL U5716 ( .A(\m02.addrM [13]), .B(\m02.addrM [14]), .C(n5609), .Z(n5701) );
  CNR2X1 U5717 ( .A(n5674), .B(n5610), .Z(n5611) );
  CND2X1 U5718 ( .A(\m02.addrM [4]), .B(n5611), .Z(n5612) );
  CND2X1 U5719 ( .A(n5634), .B(n5612), .Z(n5664) );
  CANR1XL U5720 ( .A(\m02.addrM [4]), .B(n5663), .C(n5664), .Z(n5660) );
  CNR2X1 U5721 ( .A(n5692), .B(\m02.addrM [5]), .Z(n5675) );
  CNR2IX1 U5722 ( .B(n5675), .A(n7565), .Z(n5659) );
  CANR3X1 U5723 ( .A(\m02.addrM [1]), .B(\m02.addrM [0]), .C(\m02.addrM [2]), 
        .D(\m02.addrM [3]), .Z(n5613) );
  CANR4CX1 U5724 ( .A(n5613), .B(n5619), .C(n5621), .D(n5677), .Z(n5614) );
  COND4CX1 U5725 ( .A(n5660), .B(n5659), .C(n5614), .D(n5622), .Z(n5615) );
  CNR4X1 U5726 ( .A(\m02.addrM [11]), .B(\m02.addrM [12]), .C(n5701), .D(n5615), .Z(n5616) );
  CNIVX1 U5727 ( .A(n5616), .Z(n7268) );
  CANR2XL U5728 ( .A(\s05.dataOut [0]), .B(n7269), .C(\s10.dataOut [0]), .D(
        n7268), .Z(n5708) );
  CIVX2 U5729 ( .A(n5617), .Z(n5627) );
  CIVX2 U5730 ( .A(n5618), .Z(n5624) );
  CNR2X1 U5731 ( .A(\m02.addrM [2]), .B(\m02.addrM [3]), .Z(n5620) );
  CNR2X1 U5732 ( .A(n5620), .B(n5619), .Z(n5665) );
  CANR1XL U5733 ( .A(n5665), .B(n5621), .C(n5646), .Z(n5623) );
  COND4CX1 U5734 ( .A(n5624), .B(n5691), .C(n5623), .D(n5622), .Z(n5625) );
  CNR3X1 U5735 ( .A(n5627), .B(n5626), .C(n5625), .Z(n7582) );
  CANR1XL U5736 ( .A(\m02.addrM [2]), .B(\m02.addrM [3]), .C(\m02.addrM [4]), 
        .Z(n5630) );
  CIVX2 U5737 ( .A(n5628), .Z(n5629) );
  CANR2X1 U5738 ( .A(n5691), .B(n5630), .C(n5636), .D(n5629), .Z(n5633) );
  CNR2X1 U5739 ( .A(\m02.addrM [11]), .B(\m02.addrM [12]), .Z(n5632) );
  CND2X1 U5740 ( .A(n5632), .B(n5631), .Z(n5686) );
  CANR3X1 U5741 ( .A(n5633), .B(n5639), .C(n5701), .D(n5686), .Z(n7270) );
  CANR2XL U5742 ( .A(\s04.dataOut [0]), .B(n7582), .C(\s13.dataOut [0]), .D(
        n7270), .Z(n5706) );
  CIVX2 U5743 ( .A(n5634), .Z(n5684) );
  CND2X1 U5744 ( .A(n5684), .B(n5635), .Z(n5650) );
  CANR2X1 U5745 ( .A(n5675), .B(n5650), .C(n5636), .D(n5690), .Z(n5640) );
  CND3XL U5746 ( .A(n5659), .B(n5674), .C(n5637), .Z(n5638) );
  CAN4X1 U5747 ( .A(n5640), .B(n5639), .C(n5677), .D(n5638), .Z(n5643) );
  CND2X1 U5748 ( .A(\m02.addrM [15]), .B(\m02.addrM [16]), .Z(n5642) );
  CND2X1 U5749 ( .A(\m02.addrM [13]), .B(\m02.addrM [14]), .Z(n5641) );
  CNR4X1 U5750 ( .A(n5643), .B(n5700), .C(n5642), .D(n5641), .Z(n5644) );
  CNIVX1 U5751 ( .A(n5644), .Z(n7552) );
  CIVX2 U5752 ( .A(n5645), .Z(n5648) );
  COND4CX1 U5753 ( .A(n5648), .B(n5677), .C(n5647), .D(n5646), .Z(n5649) );
  CANR1XL U5754 ( .A(n5682), .B(n5650), .C(n5649), .Z(n5655) );
  CND4X1 U5755 ( .A(\m02.addrM [9]), .B(n5653), .C(n5652), .D(n5651), .Z(n5654) );
  CANR4CX1 U5756 ( .A(n5657), .B(n5656), .C(n5655), .D(n5654), .Z(n7518) );
  CANR2XL U5757 ( .A(\s07.dataOut [0]), .B(n7552), .C(\s12.dataOut [0]), .D(
        n7518), .Z(n5705) );
  CANR2X1 U5758 ( .A(n5682), .B(n5660), .C(n5659), .D(n5658), .Z(n5662) );
  CNR3X1 U5759 ( .A(n5662), .B(n5685), .C(n5661), .Z(n7534) );
  CND2IX1 U5760 ( .B(n5663), .A(n5693), .Z(n5676) );
  CIVX2 U5761 ( .A(n5676), .Z(n5669) );
  CANR1XL U5762 ( .A(\m02.addrM [1]), .B(n5665), .C(n5664), .Z(n5667) );
  CANR1XL U5763 ( .A(n5693), .B(n5667), .C(n5666), .Z(n5668) );
  CANR11X1 U5764 ( .A(n5670), .B(n5683), .C(n5669), .D(n5668), .Z(n5672) );
  CNR3X1 U5765 ( .A(n5672), .B(n5671), .C(n5701), .Z(n7272) );
  CANR2X1 U5766 ( .A(\s06.dataOut [0]), .B(n7534), .C(\s01.dataOut [0]), .D(
        n7272), .Z(n5704) );
  CIVX2 U5767 ( .A(n5690), .Z(n5673) );
  CANR11X1 U5768 ( .A(\m02.addrM [1]), .B(n5698), .C(n5674), .D(n5673), .Z(
        n5680) );
  CND2IX1 U5769 ( .B(n5689), .A(n5693), .Z(n5679) );
  CANR11X1 U5770 ( .A(\m02.addrM [4]), .B(n5683), .C(n5676), .D(n5675), .Z(
        n5678) );
  COND3X1 U5771 ( .A(n5680), .B(n5679), .C(n5678), .D(n5677), .Z(n5681) );
  CANR3X1 U5772 ( .A(n5684), .B(n5683), .C(n5682), .D(n5681), .Z(n5687) );
  CANR3X1 U5773 ( .A(n5688), .B(n5687), .C(n5686), .D(n5685), .Z(n7273) );
  CANR11X1 U5774 ( .A(\m02.addrM [6]), .B(\m02.addrM [5]), .C(n5690), .D(n5689), .Z(n5697) );
  CND2X1 U5775 ( .A(\m02.addrM [4]), .B(n5691), .Z(n5694) );
  COND2X1 U5776 ( .A(n5695), .B(n5694), .C(n5693), .D(n5692), .Z(n5696) );
  CANR3X1 U5777 ( .A(n5699), .B(n5698), .C(n5697), .D(n5696), .Z(n5702) );
  CNR3X1 U5778 ( .A(n5702), .B(n5701), .C(n5700), .Z(n7271) );
  CANR2XL U5779 ( .A(\s11.dataOut [0]), .B(n7273), .C(\s09.dataOut [0]), .D(
        n7271), .Z(n5703) );
  CAN4X1 U5780 ( .A(n5706), .B(n5705), .C(n5704), .D(n5703), .Z(n5707) );
  CND4X1 U5781 ( .A(n5710), .B(n5709), .C(n5708), .D(n5707), .Z(n5728) );
  CNR3XL U5782 ( .A(n7269), .B(n7268), .C(n7267), .Z(n5727) );
  COR4XL U5783 ( .A(n7518), .B(n7552), .C(n7582), .D(n7266), .Z(n5712) );
  COR4XL U5784 ( .A(n7271), .B(n7534), .C(n7273), .D(n7272), .Z(n5711) );
  CNR4XL U5785 ( .A(n7265), .B(n7264), .C(n5712), .D(n5711), .Z(n5726) );
  CIVXL U5786 ( .A(n7270), .Z(n5725) );
  CNR3XL U5787 ( .A(\m02.addrM [25]), .B(\m02.addrM [26]), .C(\m02.addrM [24]), 
        .Z(n5713) );
  CND2X1 U5788 ( .A(\m02.addrM [18]), .B(n5713), .Z(n5723) );
  CND4X1 U5789 ( .A(\m02.addrM [22]), .B(\m02.addrM [21]), .C(\m02.addrM [17]), 
        .D(\m02.addrM [23]), .Z(n5722) );
  CNR4X1 U5790 ( .A(\m02.addrM [44]), .B(\m02.addrM [45]), .C(\m02.addrM [46]), 
        .D(\m02.addrM [47]), .Z(n5714) );
  CND3XL U5791 ( .A(\m02.addrM [20]), .B(\m02.addrM [19]), .C(n5714), .Z(n5720) );
  COR4X1 U5792 ( .A(\m02.addrM [31]), .B(\m02.addrM [32]), .C(\m02.addrM [33]), 
        .D(\m02.addrM [34]), .Z(n5718) );
  COR4X1 U5793 ( .A(\m02.addrM [27]), .B(\m02.addrM [28]), .C(\m02.addrM [29]), 
        .D(\m02.addrM [30]), .Z(n5717) );
  CNR2XL U5794 ( .A(\m00.YouGotIt ), .B(\m01.YouGotIt ), .Z(n5961) );
  CND2XL U5795 ( .A(\m02.YouGotIt ), .B(n5961), .Z(n7564) );
  COR4X1 U5796 ( .A(\m02.addrM [35]), .B(\m02.addrM [36]), .C(\m02.addrM [37]), 
        .D(\m02.addrM [38]), .Z(n5715) );
  COR4X1 U5797 ( .A(\m02.addrM [40]), .B(\m02.addrM [41]), .C(\m02.addrM [39]), 
        .D(n5715), .Z(n5716) );
  COR4X1 U5798 ( .A(n5718), .B(n5717), .C(n7564), .D(n5716), .Z(n5719) );
  COR4X1 U5799 ( .A(\m02.addrM [42]), .B(\m02.addrM [43]), .C(n5720), .D(n5719), .Z(n5721) );
  CNR3X1 U5800 ( .A(n5723), .B(n5722), .C(n5721), .Z(n7583) );
  CIVX2 U5801 ( .A(n7583), .Z(n5724) );
  CANR11X1 U5802 ( .A(n5727), .B(n5726), .C(n5725), .D(n5724), .Z(n7282) );
  CMX2XL U5803 ( .A0(\m02.DinMast [0]), .A1(n5728), .S(n7282), .Z(n4242) );
  CANR2XL U5804 ( .A(n7265), .B(\s00.dataOut [1]), .C(n7264), .D(
        \s03.dataOut [1]), .Z(n5736) );
  CANR2XL U5805 ( .A(\s10.dataOut [1]), .B(n7268), .C(\s02.dataOut [1]), .D(
        n7267), .Z(n5735) );
  CANR2X1 U5806 ( .A(\s05.dataOut [1]), .B(n7269), .C(\s04.dataOut [1]), .D(
        n7582), .Z(n5734) );
  CANR2XL U5807 ( .A(\s12.dataOut [1]), .B(n7518), .C(\s13.dataOut [1]), .D(
        n7270), .Z(n5732) );
  CANR2XL U5808 ( .A(\s06.dataOut [1]), .B(n7534), .C(\s08.dataOut [1]), .D(
        n7266), .Z(n5731) );
  CANR2XL U5809 ( .A(\s07.dataOut [1]), .B(n7552), .C(\s09.dataOut [1]), .D(
        n7271), .Z(n5730) );
  CANR2XL U5810 ( .A(\s11.dataOut [1]), .B(n7273), .C(\s01.dataOut [1]), .D(
        n7272), .Z(n5729) );
  CAN4X1 U5811 ( .A(n5732), .B(n5731), .C(n5730), .D(n5729), .Z(n5733) );
  CND4X1 U5812 ( .A(n5736), .B(n5735), .C(n5734), .D(n5733), .Z(n5737) );
  CMX2XL U5813 ( .A0(\m02.DinMast [1]), .A1(n5737), .S(n7282), .Z(n4243) );
  CANR2XL U5814 ( .A(n7265), .B(\s00.dataOut [2]), .C(n7264), .D(
        \s03.dataOut [2]), .Z(n5745) );
  CANR2XL U5815 ( .A(\s13.dataOut [2]), .B(n7270), .C(\s08.dataOut [2]), .D(
        n7266), .Z(n5744) );
  CANR2XL U5816 ( .A(\s02.dataOut [2]), .B(n7267), .C(\s10.dataOut [2]), .D(
        n7268), .Z(n5743) );
  CANR2XL U5817 ( .A(\s12.dataOut [2]), .B(n7518), .C(\s07.dataOut [2]), .D(
        n7552), .Z(n5741) );
  CANR2X1 U5818 ( .A(\s06.dataOut [2]), .B(n7534), .C(\s04.dataOut [2]), .D(
        n7582), .Z(n5740) );
  CANR2X1 U5819 ( .A(\s05.dataOut [2]), .B(n7269), .C(\s09.dataOut [2]), .D(
        n7271), .Z(n5739) );
  CANR2XL U5820 ( .A(\s11.dataOut [2]), .B(n7273), .C(\s01.dataOut [2]), .D(
        n7272), .Z(n5738) );
  CAN4X1 U5821 ( .A(n5741), .B(n5740), .C(n5739), .D(n5738), .Z(n5742) );
  CND4X1 U5822 ( .A(n5745), .B(n5744), .C(n5743), .D(n5742), .Z(n5746) );
  CMX2XL U5823 ( .A0(\m02.DinMast [2]), .A1(n5746), .S(n7282), .Z(n4244) );
  CANR2XL U5824 ( .A(n7265), .B(\s00.dataOut [3]), .C(n7264), .D(
        \s03.dataOut [3]), .Z(n5754) );
  CANR2X1 U5825 ( .A(\s06.dataOut [3]), .B(n7534), .C(\s02.dataOut [3]), .D(
        n7267), .Z(n5753) );
  CANR2XL U5826 ( .A(\s04.dataOut [3]), .B(n7582), .C(\s12.dataOut [3]), .D(
        n7518), .Z(n5752) );
  CANR2XL U5827 ( .A(\s05.dataOut [3]), .B(n7269), .C(\s08.dataOut [3]), .D(
        n7266), .Z(n5750) );
  CANR2XL U5828 ( .A(\s07.dataOut [3]), .B(n7552), .C(\s10.dataOut [3]), .D(
        n7268), .Z(n5749) );
  CANR2XL U5829 ( .A(\s13.dataOut [3]), .B(n7270), .C(\s11.dataOut [3]), .D(
        n7273), .Z(n5748) );
  CANR2X1 U5830 ( .A(\s01.dataOut [3]), .B(n7272), .C(\s09.dataOut [3]), .D(
        n7271), .Z(n5747) );
  CAN4X1 U5831 ( .A(n5750), .B(n5749), .C(n5748), .D(n5747), .Z(n5751) );
  CND4X1 U5832 ( .A(n5754), .B(n5753), .C(n5752), .D(n5751), .Z(n5755) );
  CMX2XL U5833 ( .A0(\m02.DinMast [3]), .A1(n5755), .S(n7282), .Z(n4245) );
  CANR2XL U5834 ( .A(n7265), .B(\s00.dataOut [4]), .C(n7264), .D(
        \s03.dataOut [4]), .Z(n5763) );
  CANR2XL U5835 ( .A(\s06.dataOut [4]), .B(n7534), .C(\s02.dataOut [4]), .D(
        n7267), .Z(n5762) );
  CANR2XL U5836 ( .A(\s13.dataOut [4]), .B(n7270), .C(\s07.dataOut [4]), .D(
        n7552), .Z(n5761) );
  CANR2XL U5837 ( .A(\s10.dataOut [4]), .B(n7268), .C(\s08.dataOut [4]), .D(
        n7266), .Z(n5759) );
  CANR2XL U5838 ( .A(\s05.dataOut [4]), .B(n7269), .C(\s12.dataOut [4]), .D(
        n7518), .Z(n5758) );
  CANR2XL U5839 ( .A(\s04.dataOut [4]), .B(n7582), .C(\s09.dataOut [4]), .D(
        n7271), .Z(n5757) );
  CANR2XL U5840 ( .A(\s11.dataOut [4]), .B(n7273), .C(\s01.dataOut [4]), .D(
        n7272), .Z(n5756) );
  CAN4X1 U5841 ( .A(n5759), .B(n5758), .C(n5757), .D(n5756), .Z(n5760) );
  CND4X1 U5842 ( .A(n5763), .B(n5762), .C(n5761), .D(n5760), .Z(n5764) );
  CMX2XL U5843 ( .A0(\m02.DinMast [4]), .A1(n5764), .S(n7282), .Z(n4246) );
  CANR2XL U5844 ( .A(n7265), .B(\s00.dataOut [5]), .C(n7264), .D(
        \s03.dataOut [5]), .Z(n5772) );
  CANR2XL U5845 ( .A(\s07.dataOut [5]), .B(n7552), .C(\s02.dataOut [5]), .D(
        n7267), .Z(n5771) );
  CANR2XL U5846 ( .A(\s06.dataOut [5]), .B(n7534), .C(\s13.dataOut [5]), .D(
        n7270), .Z(n5770) );
  CANR2XL U5847 ( .A(\s12.dataOut [5]), .B(n7518), .C(\s04.dataOut [5]), .D(
        n7582), .Z(n5768) );
  CANR2XL U5848 ( .A(\s05.dataOut [5]), .B(n7269), .C(\s08.dataOut [5]), .D(
        n7266), .Z(n5767) );
  CANR2XL U5849 ( .A(\s01.dataOut [5]), .B(n7272), .C(\s11.dataOut [5]), .D(
        n7273), .Z(n5766) );
  CANR2XL U5850 ( .A(\s09.dataOut [5]), .B(n7271), .C(\s10.dataOut [5]), .D(
        n7268), .Z(n5765) );
  CAN4X1 U5851 ( .A(n5768), .B(n5767), .C(n5766), .D(n5765), .Z(n5769) );
  CND4X1 U5852 ( .A(n5772), .B(n5771), .C(n5770), .D(n5769), .Z(n5773) );
  CMX2XL U5853 ( .A0(\m02.DinMast [5]), .A1(n5773), .S(n7282), .Z(n4247) );
  CANR2XL U5854 ( .A(n7265), .B(\s00.dataOut [6]), .C(n7264), .D(
        \s03.dataOut [6]), .Z(n5781) );
  CANR2XL U5855 ( .A(\s04.dataOut [6]), .B(n7582), .C(\s02.dataOut [6]), .D(
        n7267), .Z(n5780) );
  CANR2XL U5856 ( .A(\s12.dataOut [6]), .B(n7518), .C(\s13.dataOut [6]), .D(
        n7270), .Z(n5779) );
  CANR2XL U5857 ( .A(\s06.dataOut [6]), .B(n7534), .C(\s05.dataOut [6]), .D(
        n7269), .Z(n5777) );
  CANR2XL U5858 ( .A(\s07.dataOut [6]), .B(n7552), .C(\s08.dataOut [6]), .D(
        n7266), .Z(n5776) );
  CANR2X1 U5859 ( .A(\s09.dataOut [6]), .B(n7271), .C(\s01.dataOut [6]), .D(
        n7272), .Z(n5775) );
  CANR2XL U5860 ( .A(\s10.dataOut [6]), .B(n7268), .C(\s11.dataOut [6]), .D(
        n7273), .Z(n5774) );
  CAN4X1 U5861 ( .A(n5777), .B(n5776), .C(n5775), .D(n5774), .Z(n5778) );
  CND4X1 U5862 ( .A(n5781), .B(n5780), .C(n5779), .D(n5778), .Z(n5782) );
  CMX2XL U5863 ( .A0(\m02.DinMast [6]), .A1(n5782), .S(n7282), .Z(n4248) );
  CANR2XL U5864 ( .A(n7265), .B(\s00.dataOut [7]), .C(n7264), .D(
        \s03.dataOut [7]), .Z(n5790) );
  CANR2XL U5865 ( .A(\s02.dataOut [7]), .B(n7267), .C(\s10.dataOut [7]), .D(
        n7268), .Z(n5789) );
  CANR2XL U5866 ( .A(\s06.dataOut [7]), .B(n7534), .C(\s13.dataOut [7]), .D(
        n7270), .Z(n5788) );
  CANR2XL U5867 ( .A(\s12.dataOut [7]), .B(n7518), .C(\s08.dataOut [7]), .D(
        n7266), .Z(n5786) );
  CANR2X1 U5868 ( .A(\s04.dataOut [7]), .B(n7582), .C(\s05.dataOut [7]), .D(
        n7269), .Z(n5785) );
  CANR2XL U5869 ( .A(\s09.dataOut [7]), .B(n7271), .C(\s07.dataOut [7]), .D(
        n7552), .Z(n5784) );
  CANR2XL U5870 ( .A(\s01.dataOut [7]), .B(n7272), .C(\s11.dataOut [7]), .D(
        n7273), .Z(n5783) );
  CAN4X1 U5871 ( .A(n5786), .B(n5785), .C(n5784), .D(n5783), .Z(n5787) );
  CND4X1 U5872 ( .A(n5790), .B(n5789), .C(n5788), .D(n5787), .Z(n5791) );
  CMX2XL U5873 ( .A0(\m02.DinMast [7]), .A1(n5791), .S(n7282), .Z(n4249) );
  CANR2XL U5874 ( .A(n7265), .B(\s00.dataOut [8]), .C(n7264), .D(
        \s03.dataOut [8]), .Z(n5799) );
  CANR2XL U5875 ( .A(\s06.dataOut [8]), .B(n7534), .C(\s02.dataOut [8]), .D(
        n7267), .Z(n5798) );
  CANR2XL U5876 ( .A(\s04.dataOut [8]), .B(n7582), .C(\s13.dataOut [8]), .D(
        n7270), .Z(n5797) );
  CANR2XL U5877 ( .A(\s12.dataOut [8]), .B(n7518), .C(\s08.dataOut [8]), .D(
        n7266), .Z(n5795) );
  CANR2XL U5878 ( .A(\s07.dataOut [8]), .B(n7552), .C(\s05.dataOut [8]), .D(
        n7269), .Z(n5794) );
  CANR2XL U5879 ( .A(\s09.dataOut [8]), .B(n7271), .C(\s11.dataOut [8]), .D(
        n7273), .Z(n5793) );
  CANR2XL U5880 ( .A(\s01.dataOut [8]), .B(n7272), .C(\s10.dataOut [8]), .D(
        n7268), .Z(n5792) );
  CAN4X1 U5881 ( .A(n5795), .B(n5794), .C(n5793), .D(n5792), .Z(n5796) );
  CND4X1 U5882 ( .A(n5799), .B(n5798), .C(n5797), .D(n5796), .Z(n5800) );
  CMX2XL U5883 ( .A0(\m02.DinMast [8]), .A1(n5800), .S(n7282), .Z(n4250) );
  CANR2XL U5884 ( .A(n7265), .B(\s00.dataOut [9]), .C(n7264), .D(
        \s03.dataOut [9]), .Z(n5808) );
  CANR2XL U5885 ( .A(\s06.dataOut [9]), .B(n7534), .C(\s13.dataOut [9]), .D(
        n7270), .Z(n5807) );
  CANR2XL U5886 ( .A(\s07.dataOut [9]), .B(n7552), .C(\s02.dataOut [9]), .D(
        n7267), .Z(n5806) );
  CANR2X1 U5887 ( .A(\s04.dataOut [9]), .B(n7582), .C(\s05.dataOut [9]), .D(
        n7269), .Z(n5804) );
  CANR2XL U5888 ( .A(\s08.dataOut [9]), .B(n7266), .C(\s10.dataOut [9]), .D(
        n7268), .Z(n5803) );
  CANR2XL U5889 ( .A(\s12.dataOut [9]), .B(n7518), .C(\s09.dataOut [9]), .D(
        n7271), .Z(n5802) );
  CANR2XL U5890 ( .A(\s11.dataOut [9]), .B(n7273), .C(\s01.dataOut [9]), .D(
        n7272), .Z(n5801) );
  CAN4X1 U5891 ( .A(n5804), .B(n5803), .C(n5802), .D(n5801), .Z(n5805) );
  CND4X1 U5892 ( .A(n5808), .B(n5807), .C(n5806), .D(n5805), .Z(n5809) );
  CMX2XL U5893 ( .A0(\m02.DinMast [9]), .A1(n5809), .S(n7282), .Z(n4251) );
  CANR2XL U5894 ( .A(n7265), .B(\s00.dataOut [10]), .C(n7264), .D(
        \s03.dataOut [10]), .Z(n5817) );
  CANR2X1 U5895 ( .A(\s04.dataOut [10]), .B(n7582), .C(\s02.dataOut [10]), .D(
        n7267), .Z(n5816) );
  CANR2X1 U5896 ( .A(\s05.dataOut [10]), .B(n7269), .C(\s06.dataOut [10]), .D(
        n7534), .Z(n5815) );
  CANR2XL U5897 ( .A(\s13.dataOut [10]), .B(n7270), .C(\s10.dataOut [10]), .D(
        n7268), .Z(n5813) );
  CANR2XL U5898 ( .A(\s12.dataOut [10]), .B(n7518), .C(\s08.dataOut [10]), .D(
        n7266), .Z(n5812) );
  CANR2X1 U5899 ( .A(\s09.dataOut [10]), .B(n7271), .C(\s01.dataOut [10]), .D(
        n7272), .Z(n5811) );
  CANR2XL U5900 ( .A(\s07.dataOut [10]), .B(n7552), .C(\s11.dataOut [10]), .D(
        n7273), .Z(n5810) );
  CAN4X1 U5901 ( .A(n5813), .B(n5812), .C(n5811), .D(n5810), .Z(n5814) );
  CND4X1 U5902 ( .A(n5817), .B(n5816), .C(n5815), .D(n5814), .Z(n5818) );
  CMX2XL U5903 ( .A0(\m02.DinMast [10]), .A1(n5818), .S(n7282), .Z(n4252) );
  CANR2XL U5904 ( .A(n7265), .B(\s00.dataOut [11]), .C(n7264), .D(
        \s03.dataOut [11]), .Z(n5826) );
  CANR2XL U5905 ( .A(\s12.dataOut [11]), .B(n7518), .C(\s02.dataOut [11]), .D(
        n7267), .Z(n5825) );
  CANR2XL U5906 ( .A(\s06.dataOut [11]), .B(n7534), .C(\s08.dataOut [11]), .D(
        n7266), .Z(n5824) );
  CANR2XL U5907 ( .A(\s04.dataOut [11]), .B(n7582), .C(\s10.dataOut [11]), .D(
        n7268), .Z(n5822) );
  CANR2XL U5908 ( .A(\s05.dataOut [11]), .B(n7269), .C(\s07.dataOut [11]), .D(
        n7552), .Z(n5821) );
  CANR2XL U5909 ( .A(\s13.dataOut [11]), .B(n7270), .C(\s01.dataOut [11]), .D(
        n7272), .Z(n5820) );
  CANR2XL U5910 ( .A(\s11.dataOut [11]), .B(n7273), .C(\s09.dataOut [11]), .D(
        n7271), .Z(n5819) );
  CAN4X1 U5911 ( .A(n5822), .B(n5821), .C(n5820), .D(n5819), .Z(n5823) );
  CND4X1 U5912 ( .A(n5826), .B(n5825), .C(n5824), .D(n5823), .Z(n5827) );
  CMX2XL U5913 ( .A0(\m02.DinMast [11]), .A1(n5827), .S(n7282), .Z(n4253) );
  CNR2X1 U5914 ( .A(\m05.addrM [5]), .B(\m05.addrM [6]), .Z(n5849) );
  CNR2X1 U5915 ( .A(\m05.addrM [4]), .B(\m05.addrM [3]), .Z(n5832) );
  CIVX2 U5916 ( .A(\m05.addrM [4]), .Z(n5902) );
  CND2X1 U5917 ( .A(\m05.addrM [1]), .B(\m05.addrM [2]), .Z(n5845) );
  CND2X1 U5918 ( .A(n5902), .B(n5845), .Z(n5935) );
  CND2IX1 U5919 ( .B(n5832), .A(n5935), .Z(n5925) );
  CNR2X1 U5920 ( .A(\m05.addrM [0]), .B(\m05.addrM [1]), .Z(n5944) );
  CIVX2 U5921 ( .A(n5944), .Z(n5828) );
  CANR1XL U5922 ( .A(\m05.addrM [2]), .B(n5828), .C(\m05.addrM [3]), .Z(n5833)
         );
  CNR2X1 U5923 ( .A(\m05.addrM [4]), .B(n5833), .Z(n5887) );
  CND2X1 U5924 ( .A(\m05.addrM [5]), .B(n5887), .Z(n5829) );
  CIVX2 U5925 ( .A(\m05.addrM [7]), .Z(n5848) );
  CNR2X1 U5926 ( .A(\m05.addrM [8]), .B(n5848), .Z(n5942) );
  CIVX2 U5927 ( .A(n5942), .Z(n5871) );
  CANR4CX1 U5928 ( .A(n5849), .B(n5925), .C(n5829), .D(n5871), .Z(n5831) );
  CIVX2 U5929 ( .A(\m05.addrM [5]), .Z(n5931) );
  CIVX2 U5930 ( .A(\m05.addrM [6]), .Z(n5930) );
  CNR2X1 U5931 ( .A(n5931), .B(n5930), .Z(n5936) );
  CNR2X1 U5932 ( .A(\m05.addrM [2]), .B(\m05.addrM [3]), .Z(n5903) );
  CIVX2 U5933 ( .A(n5903), .Z(n5879) );
  CNR2X1 U5934 ( .A(\m05.addrM [4]), .B(n5879), .Z(n5950) );
  CIVX2 U5935 ( .A(\m05.addrM [1]), .Z(n5847) );
  CND2X1 U5936 ( .A(n5950), .B(n5847), .Z(n5896) );
  CND2X1 U5937 ( .A(\m05.addrM [8]), .B(n5848), .Z(n5928) );
  CNR2X1 U5938 ( .A(n5930), .B(n5871), .Z(n5913) );
  CIVX2 U5939 ( .A(n5849), .Z(n5834) );
  CNR2X1 U5940 ( .A(n5834), .B(n5928), .Z(n5943) );
  CNR2X1 U5941 ( .A(n5913), .B(n5943), .Z(n5839) );
  COND4CX1 U5942 ( .A(n5936), .B(n5896), .C(n5928), .D(n5839), .Z(n5830) );
  CIVXL U5943 ( .A(\m05.addrM [9]), .Z(n5857) );
  CND2X1 U5944 ( .A(\m05.addrM [10]), .B(n5857), .Z(n5911) );
  CND2X1 U5945 ( .A(\m05.addrM [12]), .B(\m05.addrM [11]), .Z(n5926) );
  CNR2X1 U5946 ( .A(n5911), .B(n5926), .Z(n5937) );
  CIVX2 U5947 ( .A(\m05.addrM [14]), .Z(n5882) );
  CND2X1 U5948 ( .A(\m05.addrM [16]), .B(n5882), .Z(n5858) );
  CIVXL U5949 ( .A(\m05.addrM [15]), .Z(n5881) );
  CND2X1 U5950 ( .A(\m05.addrM [13]), .B(n5881), .Z(n5835) );
  CNR2X1 U5951 ( .A(n5858), .B(n5835), .Z(n5946) );
  COND3X1 U5952 ( .A(n5831), .B(n5830), .C(n5937), .D(n5946), .Z(n6664) );
  CIVX2 U5953 ( .A(n6664), .Z(n6727) );
  CND2X1 U5954 ( .A(n5942), .B(n5849), .Z(n5838) );
  CND2X1 U5955 ( .A(n5832), .B(n5845), .Z(n5841) );
  CNR2X1 U5956 ( .A(n5902), .B(n5833), .Z(n5895) );
  CIVX2 U5957 ( .A(\m05.addrM [8]), .Z(n5917) );
  COND3X1 U5958 ( .A(n5895), .B(n5834), .C(n5848), .D(n5917), .Z(n5837) );
  CND2X1 U5959 ( .A(\m05.addrM [16]), .B(\m05.addrM [14]), .Z(n5870) );
  CNR2X1 U5960 ( .A(n5835), .B(n5870), .Z(n5940) );
  CIVX2 U5961 ( .A(\m05.addrM [11]), .Z(n5859) );
  CND2X1 U5962 ( .A(\m05.addrM [12]), .B(n5859), .Z(n5890) );
  CNR2X1 U5963 ( .A(\m05.addrM [9]), .B(\m05.addrM [10]), .Z(n5855) );
  CIVX2 U5964 ( .A(n5855), .Z(n5843) );
  CNR2X1 U5965 ( .A(n5890), .B(n5843), .Z(n5945) );
  CND2X1 U5966 ( .A(n5940), .B(n5945), .Z(n5836) );
  CANR4CX1 U5967 ( .A(n5838), .B(n5841), .C(n5837), .D(n5836), .Z(n6726) );
  CANR2XL U5968 ( .A(n6727), .B(\s03.dataOut [15]), .C(\s01.dataOut [15]), .D(
        n6726), .Z(n5958) );
  CIVX2 U5969 ( .A(n5936), .Z(n5894) );
  CNR2X1 U5970 ( .A(\m05.addrM [8]), .B(n5894), .Z(n5864) );
  CANR3X1 U5971 ( .A(\m05.addrM [2]), .B(\m05.addrM [3]), .C(\m05.addrM [4]), 
        .D(n5839), .Z(n5840) );
  CANR3X1 U5972 ( .A(n5864), .B(n5841), .C(n5942), .D(n5840), .Z(n5844) );
  CNR2X1 U5973 ( .A(\m05.addrM [12]), .B(\m05.addrM [11]), .Z(n5842) );
  CND2X1 U5974 ( .A(n5940), .B(n5842), .Z(n5910) );
  CNR3X1 U5975 ( .A(n5844), .B(n5843), .C(n5910), .Z(n6728) );
  CNR2X1 U5976 ( .A(n5849), .B(n5871), .Z(n5854) );
  CIVX2 U5977 ( .A(n5928), .Z(n5869) );
  CND2X1 U5978 ( .A(\m05.addrM [4]), .B(\m05.addrM [3]), .Z(n5874) );
  CND2IX1 U5979 ( .B(n5845), .A(\m05.addrM [4]), .Z(n5846) );
  CANR1XL U5980 ( .A(n5874), .B(n5846), .C(n5871), .Z(n5853) );
  CNR2X1 U5981 ( .A(n5847), .B(\m05.addrM [0]), .Z(n5868) );
  CIVX2 U5982 ( .A(n5868), .Z(n5851) );
  COND1XL U5983 ( .A(\m05.addrM [1]), .B(\m05.addrM [2]), .C(\m05.addrM [3]), 
        .Z(n5860) );
  CND2X1 U5984 ( .A(n5902), .B(n5860), .Z(n5934) );
  CNR2X1 U5985 ( .A(n5848), .B(n5917), .Z(n5932) );
  CND2X1 U5986 ( .A(n5849), .B(n5932), .Z(n5850) );
  CANR4CX1 U5987 ( .A(n5935), .B(n5851), .C(n5934), .D(n5850), .Z(n5852) );
  CNR4X1 U5988 ( .A(n5854), .B(n5869), .C(n5853), .D(n5852), .Z(n5856) );
  CNR3XL U5989 ( .A(\m05.addrM [13]), .B(\m05.addrM [15]), .C(n5870), .Z(n5898) );
  CND2X1 U5990 ( .A(n5898), .B(n5855), .Z(n5924) );
  CNR4X1 U5991 ( .A(\m05.addrM [12]), .B(\m05.addrM [11]), .C(n5856), .D(n5924), .Z(n5959) );
  CANR2XL U5992 ( .A(\s13.dataOut [15]), .B(n6728), .C(\s11.dataOut [15]), .D(
        n6733), .Z(n5957) );
  CNR2X1 U5993 ( .A(\m05.addrM [10]), .B(n5857), .Z(n5889) );
  CNR3XL U5994 ( .A(\m05.addrM [12]), .B(n5859), .C(n5858), .Z(n5923) );
  CNR2IX1 U5995 ( .B(\m05.addrM [13]), .A(n5881), .Z(n5863) );
  CNR2X1 U5996 ( .A(n5902), .B(n5860), .Z(n5866) );
  COND1XL U5997 ( .A(\m05.addrM [5]), .B(n5896), .C(n5913), .Z(n5861) );
  COND4CX1 U5998 ( .A(n5936), .B(n5866), .C(n5928), .D(n5861), .Z(n5862) );
  CAN4X1 U5999 ( .A(n5889), .B(n5923), .C(n5863), .D(n5862), .Z(n6734) );
  CND2X1 U6000 ( .A(n5869), .B(n5894), .Z(n5865) );
  CNR2X1 U6001 ( .A(n5930), .B(n5865), .Z(n5905) );
  CIVX2 U6002 ( .A(\m05.addrM [2]), .Z(n5875) );
  CIVX2 U6003 ( .A(n5934), .Z(n5885) );
  CIVX2 U6004 ( .A(n5864), .Z(n5949) );
  COND2X1 U6005 ( .A(n5885), .B(n5949), .C(n5866), .D(n5865), .Z(n5867) );
  CANR11X1 U6006 ( .A(n5905), .B(n5868), .C(n5875), .D(n5867), .Z(n5872) );
  CND2X1 U6007 ( .A(n5869), .B(n5930), .Z(n5876) );
  CANR11X1 U6008 ( .A(n5872), .B(n5871), .C(n5876), .D(n5870), .Z(n5873) );
  CAN4X1 U6009 ( .A(\m05.addrM [13]), .B(\m05.addrM [15]), .C(n5937), .D(n5873), .Z(n6729) );
  CANR2X1 U6010 ( .A(\s12.dataOut [15]), .B(n6734), .C(\s07.dataOut [15]), .D(
        n6729), .Z(n5956) );
  CNR2X1 U6011 ( .A(n5875), .B(n5874), .Z(n5914) );
  CND2X1 U6012 ( .A(\m05.addrM [0]), .B(\m05.addrM [1]), .Z(n5888) );
  CNR2IX1 U6013 ( .B(n5943), .A(n5888), .Z(n5904) );
  CIVX2 U6014 ( .A(n5905), .Z(n5878) );
  CIVX2 U6015 ( .A(n5876), .Z(n5908) );
  CND2X1 U6016 ( .A(\m05.addrM [5]), .B(n5908), .Z(n5877) );
  COND4CX1 U6017 ( .A(\m05.addrM [4]), .B(n5879), .C(n5878), .D(n5877), .Z(
        n5880) );
  CANR1XL U6018 ( .A(n5914), .B(n5904), .C(n5880), .Z(n5884) );
  CNR2X1 U6019 ( .A(\m05.addrM [13]), .B(n5881), .Z(n5922) );
  CIVX2 U6020 ( .A(\m05.addrM [16]), .Z(n5883) );
  CND3XL U6021 ( .A(n5922), .B(n5883), .C(n5882), .Z(n5891) );
  CNR4X1 U6022 ( .A(n5884), .B(n5890), .C(n5911), .D(n5891), .Z(n5960) );
  CNR2X1 U6023 ( .A(n5885), .B(n5914), .Z(n5886) );
  CANR3X1 U6024 ( .A(n5914), .B(n5888), .C(n5887), .D(n5886), .Z(n5893) );
  CND2IX1 U6025 ( .B(n5890), .A(n5889), .Z(n5899) );
  CND2X1 U6026 ( .A(n5936), .B(n5932), .Z(n5892) );
  CNR4X2 U6027 ( .A(n5893), .B(n5899), .C(n5892), .D(n5891), .Z(n6731) );
  CANR2XL U6028 ( .A(\s04.dataOut [15]), .B(n6735), .C(\s05.dataOut [15]), .D(
        n6731), .Z(n5954) );
  CNR2X1 U6029 ( .A(n5894), .B(n5928), .Z(n5897) );
  CIVX2 U6030 ( .A(n5895), .Z(n5906) );
  CANR2X1 U6031 ( .A(n5897), .B(n5906), .C(n5905), .D(n5896), .Z(n5901) );
  CIVX2 U6032 ( .A(n5898), .Z(n5900) );
  CNR3X1 U6033 ( .A(n5901), .B(n5900), .C(n5899), .Z(n6730) );
  CNR2X1 U6034 ( .A(n5903), .B(n5902), .Z(n5909) );
  CAOR2X2 U6035 ( .A(n5906), .B(n5905), .C(\m05.addrM [4]), .D(n5904), .Z(
        n5907) );
  CANR4CX1 U6036 ( .A(\m05.addrM [5]), .B(n5909), .C(n5908), .D(n5907), .Z(
        n5912) );
  CNR3X1 U6037 ( .A(n5912), .B(n5911), .C(n5910), .Z(n6732) );
  CANR2XL U6038 ( .A(\s06.dataOut [15]), .B(n6730), .C(\s10.dataOut [15]), .D(
        n6732), .Z(n5953) );
  CND2X1 U6039 ( .A(n5931), .B(n5913), .Z(n5927) );
  CIVX2 U6040 ( .A(n5927), .Z(n5915) );
  COND3XL U6041 ( .A(\m05.addrM [5]), .B(n5914), .C(\m05.addrM [6]), .D(
        \m05.addrM [7]), .Z(n5916) );
  CANR2X1 U6042 ( .A(n5944), .B(n5915), .C(n5917), .D(n5916), .Z(n5920) );
  CNR2X1 U6043 ( .A(n5917), .B(n5916), .Z(n5918) );
  COND1XL U6044 ( .A(n5918), .B(\m05.addrM [9]), .C(\m05.addrM [10]), .Z(n5919) );
  CANR1XL U6045 ( .A(\m05.addrM [9]), .B(n5920), .C(n5919), .Z(n5921) );
  CND3XL U6046 ( .A(n5923), .B(n5922), .C(n5921), .Z(n6558) );
  CIVX2 U6047 ( .A(n6558), .Z(n6737) );
  CNR4X2 U6048 ( .A(n5927), .B(n5926), .C(n5925), .D(n5924), .Z(n6739) );
  CANR2X1 U6049 ( .A(n6737), .B(\s00.dataOut [15]), .C(\s02.dataOut [15]), .D(
        n6739), .Z(n5952) );
  COND11XL U6050 ( .A(\m05.addrM [1]), .B(\m05.addrM [2]), .C(\m05.addrM [3]), 
        .D(\m05.addrM [4]), .Z(n5929) );
  CANR11X1 U6051 ( .A(n5931), .B(n5930), .C(n5929), .D(n5928), .Z(n5939) );
  CIVX2 U6052 ( .A(n5932), .Z(n5933) );
  CANR11X1 U6053 ( .A(n5936), .B(n5935), .C(n5934), .D(n5933), .Z(n5938) );
  COND1XL U6054 ( .A(n5939), .B(n5938), .C(n5937), .Z(n5941) );
  CND2IX1 U6055 ( .B(n5941), .A(n5940), .Z(n6437) );
  CIVX2 U6056 ( .A(n6437), .Z(n6738) );
  CANR11X1 U6057 ( .A(n5944), .B(n5950), .C(n5943), .D(n5942), .Z(n5948) );
  CND2X1 U6058 ( .A(n5946), .B(n5945), .Z(n5947) );
  CANR4CX1 U6059 ( .A(n5950), .B(n5949), .C(n5948), .D(n5947), .Z(n6736) );
  CANR2XL U6060 ( .A(\s09.dataOut [15]), .B(n6738), .C(\s08.dataOut [15]), .D(
        n6736), .Z(n5951) );
  CAN4X1 U6061 ( .A(n5954), .B(n5953), .C(n5952), .D(n5951), .Z(n5955) );
  CND4X1 U6062 ( .A(n5958), .B(n5957), .C(n5956), .D(n5955), .Z(n5962) );
  CIVX2 U6063 ( .A(n6730), .Z(n7531) );
  CIVX2 U6064 ( .A(n6734), .Z(n7515) );
  CIVX2 U6065 ( .A(n6736), .Z(n6384) );
  CIVX2 U6066 ( .A(n6729), .Z(n7557) );
  CIVDX1 U6067 ( .A(n5959), .Z0(n6503), .Z1(n6733) );
  CIVDX1 U6068 ( .A(n5960), .Z0(n7588), .Z1(n6735) );
  CIVX2 U6069 ( .A(n6731), .Z(n6325) );
  CIVXL U6070 ( .A(n6728), .Z(n6507) );
  CIVX2 U6071 ( .A(n6726), .Z(n6601) );
  CIVX2 U6072 ( .A(n6739), .Z(n6613) );
  CIVXL U6073 ( .A(\m02.YouGotIt ), .Z(n7699) );
  CND2X1 U6074 ( .A(n5961), .B(n7699), .Z(n6284) );
  CNR2XL U6075 ( .A(\m03.YouGotIt ), .B(n6284), .Z(n6286) );
  CND2IXL U6076 ( .B(\m04.YouGotIt ), .A(n6286), .Z(n6167) );
  CIVXL U6077 ( .A(\m05.YouGotIt ), .Z(n7694) );
  COR2X1 U6078 ( .A(n6167), .B(n7694), .Z(n6285) );
  CMX2XL U6079 ( .A0(\m05.DinMast [15]), .A1(n5962), .S(n6748), .Z(n4209) );
  CANR2XL U6080 ( .A(n6727), .B(\s03.dataOut [14]), .C(\s01.dataOut [14]), .D(
        n6726), .Z(n5970) );
  CANR2XL U6081 ( .A(\s05.dataOut [14]), .B(n6731), .C(\s08.dataOut [14]), .D(
        n6736), .Z(n5969) );
  CANR2X1 U6082 ( .A(\s12.dataOut [14]), .B(n6734), .C(\s10.dataOut [14]), .D(
        n6732), .Z(n5968) );
  CANR2X1 U6083 ( .A(\s07.dataOut [14]), .B(n6729), .C(\s06.dataOut [14]), .D(
        n6730), .Z(n5966) );
  CANR2XL U6084 ( .A(\s04.dataOut [14]), .B(n6735), .C(\s11.dataOut [14]), .D(
        n6733), .Z(n5965) );
  CANR2X1 U6085 ( .A(n6737), .B(\s00.dataOut [14]), .C(\s13.dataOut [14]), .D(
        n6728), .Z(n5964) );
  CANR2X1 U6086 ( .A(\s02.dataOut [14]), .B(n6739), .C(\s09.dataOut [14]), .D(
        n6738), .Z(n5963) );
  CAN4X1 U6087 ( .A(n5966), .B(n5965), .C(n5964), .D(n5963), .Z(n5967) );
  CND4X1 U6088 ( .A(n5970), .B(n5969), .C(n5968), .D(n5967), .Z(n5971) );
  CMX2XL U6089 ( .A0(\m05.DinMast [14]), .A1(n5971), .S(n6748), .Z(n4208) );
  CANR2XL U6090 ( .A(\s09.dataOut [13]), .B(n6738), .C(\s01.dataOut [13]), .D(
        n6726), .Z(n5979) );
  CANR2XL U6091 ( .A(\s07.dataOut [13]), .B(n6729), .C(\s11.dataOut [13]), .D(
        n6733), .Z(n5978) );
  CANR2X1 U6092 ( .A(\s12.dataOut [13]), .B(n6734), .C(\s13.dataOut [13]), .D(
        n6728), .Z(n5977) );
  CANR2X1 U6093 ( .A(\s05.dataOut [13]), .B(n6731), .C(\s06.dataOut [13]), .D(
        n6730), .Z(n5975) );
  CANR2XL U6094 ( .A(\s04.dataOut [13]), .B(n6735), .C(\s10.dataOut [13]), .D(
        n6732), .Z(n5974) );
  CANR2X1 U6095 ( .A(n6737), .B(\s00.dataOut [13]), .C(n6727), .D(
        \s03.dataOut [13]), .Z(n5973) );
  CANR2XL U6096 ( .A(\s02.dataOut [13]), .B(n6739), .C(\s08.dataOut [13]), .D(
        n6736), .Z(n5972) );
  CAN4X1 U6097 ( .A(n5975), .B(n5974), .C(n5973), .D(n5972), .Z(n5976) );
  CND4X1 U6098 ( .A(n5979), .B(n5978), .C(n5977), .D(n5976), .Z(n5980) );
  CMX2XL U6099 ( .A0(\m05.DinMast [13]), .A1(n5980), .S(n6748), .Z(n4207) );
  CANR2XL U6100 ( .A(n6727), .B(\s03.dataOut [12]), .C(\s01.dataOut [12]), .D(
        n6726), .Z(n5988) );
  CANR2XL U6101 ( .A(\s04.dataOut [12]), .B(n6735), .C(\s08.dataOut [12]), .D(
        n6736), .Z(n5987) );
  CANR2X1 U6102 ( .A(\s07.dataOut [12]), .B(n6729), .C(\s10.dataOut [12]), .D(
        n6732), .Z(n5986) );
  CANR2XL U6103 ( .A(\s05.dataOut [12]), .B(n6731), .C(\s11.dataOut [12]), .D(
        n6733), .Z(n5984) );
  CANR2XL U6104 ( .A(\s06.dataOut [12]), .B(n6730), .C(\s12.dataOut [12]), .D(
        n6734), .Z(n5983) );
  CANR2X1 U6105 ( .A(n6737), .B(\s00.dataOut [12]), .C(\s02.dataOut [12]), .D(
        n6739), .Z(n5982) );
  CANR2X1 U6106 ( .A(\s13.dataOut [12]), .B(n6728), .C(\s09.dataOut [12]), .D(
        n6738), .Z(n5981) );
  CAN4X1 U6107 ( .A(n5984), .B(n5983), .C(n5982), .D(n5981), .Z(n5985) );
  CND4X1 U6108 ( .A(n5988), .B(n5987), .C(n5986), .D(n5985), .Z(n5989) );
  CMX2XL U6109 ( .A0(\m05.DinMast [12]), .A1(n5989), .S(n6748), .Z(n4206) );
  CANR2XL U6110 ( .A(\s09.dataOut [11]), .B(n6738), .C(\s01.dataOut [11]), .D(
        n6726), .Z(n5997) );
  CANR2XL U6111 ( .A(\s07.dataOut [11]), .B(n6729), .C(\s08.dataOut [11]), .D(
        n6736), .Z(n5996) );
  CANR2XL U6112 ( .A(\s05.dataOut [11]), .B(n6731), .C(\s11.dataOut [11]), .D(
        n6733), .Z(n5995) );
  CANR2XL U6113 ( .A(\s12.dataOut [11]), .B(n6734), .C(\s04.dataOut [11]), .D(
        n6735), .Z(n5993) );
  CANR2XL U6114 ( .A(\s06.dataOut [11]), .B(n6730), .C(\s10.dataOut [11]), .D(
        n6732), .Z(n5992) );
  CANR2X1 U6115 ( .A(n6737), .B(\s00.dataOut [11]), .C(\s02.dataOut [11]), .D(
        n6739), .Z(n5991) );
  CANR2X1 U6116 ( .A(n6727), .B(\s03.dataOut [11]), .C(\s13.dataOut [11]), .D(
        n6728), .Z(n5990) );
  CAN4X1 U6117 ( .A(n5993), .B(n5992), .C(n5991), .D(n5990), .Z(n5994) );
  CND4X1 U6118 ( .A(n5997), .B(n5996), .C(n5995), .D(n5994), .Z(n5998) );
  CMX2XL U6119 ( .A0(\m05.DinMast [11]), .A1(n5998), .S(n6748), .Z(n4205) );
  CANR2XL U6120 ( .A(\s09.dataOut [10]), .B(n6738), .C(\s01.dataOut [10]), .D(
        n6726), .Z(n6006) );
  CANR2XL U6121 ( .A(\s07.dataOut [10]), .B(n6729), .C(\s11.dataOut [10]), .D(
        n6733), .Z(n6005) );
  CANR2XL U6122 ( .A(\s12.dataOut [10]), .B(n6734), .C(\s08.dataOut [10]), .D(
        n6736), .Z(n6004) );
  CANR2XL U6123 ( .A(\s04.dataOut [10]), .B(n6735), .C(\s10.dataOut [10]), .D(
        n6732), .Z(n6002) );
  CANR2X1 U6124 ( .A(\s05.dataOut [10]), .B(n6731), .C(\s06.dataOut [10]), .D(
        n6730), .Z(n6001) );
  CANR2X1 U6125 ( .A(n6737), .B(\s00.dataOut [10]), .C(\s02.dataOut [10]), .D(
        n6739), .Z(n6000) );
  CANR2X1 U6126 ( .A(n6727), .B(\s03.dataOut [10]), .C(\s13.dataOut [10]), .D(
        n6728), .Z(n5999) );
  CAN4X1 U6127 ( .A(n6002), .B(n6001), .C(n6000), .D(n5999), .Z(n6003) );
  CND4X1 U6128 ( .A(n6006), .B(n6005), .C(n6004), .D(n6003), .Z(n6007) );
  CMX2XL U6129 ( .A0(\m05.DinMast [10]), .A1(n6007), .S(n6748), .Z(n4204) );
  CANR2XL U6130 ( .A(\s01.dataOut [9]), .B(n6726), .C(\s09.dataOut [9]), .D(
        n6738), .Z(n6015) );
  CANR2XL U6131 ( .A(\s08.dataOut [9]), .B(n6736), .C(\s10.dataOut [9]), .D(
        n6732), .Z(n6014) );
  CANR2X1 U6132 ( .A(\s07.dataOut [9]), .B(n6729), .C(\s05.dataOut [9]), .D(
        n6731), .Z(n6013) );
  CANR2XL U6133 ( .A(\s06.dataOut [9]), .B(n6730), .C(\s11.dataOut [9]), .D(
        n6733), .Z(n6011) );
  CANR2XL U6134 ( .A(\s12.dataOut [9]), .B(n6734), .C(\s04.dataOut [9]), .D(
        n6735), .Z(n6010) );
  CANR2X1 U6135 ( .A(n6737), .B(\s00.dataOut [9]), .C(\s02.dataOut [9]), .D(
        n6739), .Z(n6009) );
  CANR2X1 U6136 ( .A(n6727), .B(\s03.dataOut [9]), .C(\s13.dataOut [9]), .D(
        n6728), .Z(n6008) );
  CAN4X1 U6137 ( .A(n6011), .B(n6010), .C(n6009), .D(n6008), .Z(n6012) );
  CND4X1 U6138 ( .A(n6015), .B(n6014), .C(n6013), .D(n6012), .Z(n6016) );
  CMX2XL U6139 ( .A0(\m05.DinMast [9]), .A1(n6016), .S(n6748), .Z(n4203) );
  CANR2X1 U6140 ( .A(n6727), .B(\s03.dataOut [8]), .C(\s09.dataOut [8]), .D(
        n6738), .Z(n6024) );
  CANR2XL U6141 ( .A(\s08.dataOut [8]), .B(n6736), .C(\s11.dataOut [8]), .D(
        n6733), .Z(n6023) );
  CANR2X1 U6142 ( .A(\s12.dataOut [8]), .B(n6734), .C(\s05.dataOut [8]), .D(
        n6731), .Z(n6022) );
  CANR2XL U6143 ( .A(\s06.dataOut [8]), .B(n6730), .C(\s04.dataOut [8]), .D(
        n6735), .Z(n6020) );
  CANR2XL U6144 ( .A(\s07.dataOut [8]), .B(n6729), .C(\s10.dataOut [8]), .D(
        n6732), .Z(n6019) );
  CANR2X1 U6145 ( .A(n6737), .B(\s00.dataOut [8]), .C(\s02.dataOut [8]), .D(
        n6739), .Z(n6018) );
  CANR2XL U6146 ( .A(\s13.dataOut [8]), .B(n6728), .C(\s01.dataOut [8]), .D(
        n6726), .Z(n6017) );
  CAN4X1 U6147 ( .A(n6020), .B(n6019), .C(n6018), .D(n6017), .Z(n6021) );
  CND4X1 U6148 ( .A(n6024), .B(n6023), .C(n6022), .D(n6021), .Z(n6025) );
  CMX2XL U6149 ( .A0(\m05.DinMast [8]), .A1(n6025), .S(n6748), .Z(n4202) );
  CANR2X1 U6150 ( .A(n6727), .B(\s03.dataOut [7]), .C(\s09.dataOut [7]), .D(
        n6738), .Z(n6033) );
  CANR2XL U6151 ( .A(\s04.dataOut [7]), .B(n6735), .C(\s08.dataOut [7]), .D(
        n6736), .Z(n6032) );
  CANR2XL U6152 ( .A(\s12.dataOut [7]), .B(n6734), .C(\s10.dataOut [7]), .D(
        n6732), .Z(n6031) );
  CANR2XL U6153 ( .A(\s05.dataOut [7]), .B(n6731), .C(\s11.dataOut [7]), .D(
        n6733), .Z(n6029) );
  CANR2XL U6154 ( .A(\s06.dataOut [7]), .B(n6730), .C(\s07.dataOut [7]), .D(
        n6729), .Z(n6028) );
  CANR2XL U6155 ( .A(n6737), .B(\s00.dataOut [7]), .C(\s01.dataOut [7]), .D(
        n6726), .Z(n6027) );
  CANR2XL U6156 ( .A(\s02.dataOut [7]), .B(n6739), .C(\s13.dataOut [7]), .D(
        n6728), .Z(n6026) );
  CAN4X1 U6157 ( .A(n6029), .B(n6028), .C(n6027), .D(n6026), .Z(n6030) );
  CND4X1 U6158 ( .A(n6033), .B(n6032), .C(n6031), .D(n6030), .Z(n6034) );
  CMX2XL U6159 ( .A0(\m05.DinMast [7]), .A1(n6034), .S(n6748), .Z(n4201) );
  CANR2XL U6160 ( .A(n6727), .B(\s03.dataOut [6]), .C(\s01.dataOut [6]), .D(
        n6726), .Z(n6042) );
  CANR2XL U6161 ( .A(\s04.dataOut [6]), .B(n6735), .C(\s13.dataOut [6]), .D(
        n6728), .Z(n6041) );
  CANR2XL U6162 ( .A(\s06.dataOut [6]), .B(n6730), .C(\s05.dataOut [6]), .D(
        n6731), .Z(n6040) );
  CANR2XL U6163 ( .A(\s10.dataOut [6]), .B(n6732), .C(\s11.dataOut [6]), .D(
        n6733), .Z(n6038) );
  CANR2X1 U6164 ( .A(\s12.dataOut [6]), .B(n6734), .C(\s07.dataOut [6]), .D(
        n6729), .Z(n6037) );
  CANR2X1 U6165 ( .A(n6737), .B(\s00.dataOut [6]), .C(\s02.dataOut [6]), .D(
        n6739), .Z(n6036) );
  CANR2XL U6166 ( .A(\s09.dataOut [6]), .B(n6738), .C(\s08.dataOut [6]), .D(
        n6736), .Z(n6035) );
  CAN4X1 U6167 ( .A(n6038), .B(n6037), .C(n6036), .D(n6035), .Z(n6039) );
  CND4X1 U6168 ( .A(n6042), .B(n6041), .C(n6040), .D(n6039), .Z(n6043) );
  CMX2XL U6169 ( .A0(\m05.DinMast [6]), .A1(n6043), .S(n6748), .Z(n4200) );
  CANR2XL U6170 ( .A(\s01.dataOut [5]), .B(n6726), .C(\s09.dataOut [5]), .D(
        n6738), .Z(n6051) );
  CANR2XL U6171 ( .A(\s07.dataOut [5]), .B(n6729), .C(\s13.dataOut [5]), .D(
        n6728), .Z(n6050) );
  CANR2XL U6172 ( .A(\s04.dataOut [5]), .B(n6735), .C(\s11.dataOut [5]), .D(
        n6733), .Z(n6049) );
  CANR2XL U6173 ( .A(\s06.dataOut [5]), .B(n6730), .C(\s10.dataOut [5]), .D(
        n6732), .Z(n6047) );
  CANR2X1 U6174 ( .A(\s05.dataOut [5]), .B(n6731), .C(\s12.dataOut [5]), .D(
        n6734), .Z(n6046) );
  CANR2X1 U6175 ( .A(n6737), .B(\s00.dataOut [5]), .C(n6727), .D(
        \s03.dataOut [5]), .Z(n6045) );
  CANR2XL U6176 ( .A(\s02.dataOut [5]), .B(n6739), .C(\s08.dataOut [5]), .D(
        n6736), .Z(n6044) );
  CAN4X1 U6177 ( .A(n6047), .B(n6046), .C(n6045), .D(n6044), .Z(n6048) );
  CND4X1 U6178 ( .A(n6051), .B(n6050), .C(n6049), .D(n6048), .Z(n6052) );
  CMX2XL U6179 ( .A0(\m05.DinMast [5]), .A1(n6052), .S(n6748), .Z(n4199) );
  CANR2X1 U6180 ( .A(n6727), .B(\s03.dataOut [4]), .C(\s09.dataOut [4]), .D(
        n6738), .Z(n6060) );
  CANR2XL U6181 ( .A(\s06.dataOut [4]), .B(n6730), .C(\s08.dataOut [4]), .D(
        n6736), .Z(n6059) );
  CANR2XL U6182 ( .A(\s12.dataOut [4]), .B(n6734), .C(\s11.dataOut [4]), .D(
        n6733), .Z(n6058) );
  CANR2XL U6183 ( .A(\s07.dataOut [4]), .B(n6729), .C(\s10.dataOut [4]), .D(
        n6732), .Z(n6056) );
  CANR2XL U6184 ( .A(\s04.dataOut [4]), .B(n6735), .C(\s05.dataOut [4]), .D(
        n6731), .Z(n6055) );
  CANR2X1 U6185 ( .A(n6737), .B(\s00.dataOut [4]), .C(\s02.dataOut [4]), .D(
        n6739), .Z(n6054) );
  CANR2XL U6186 ( .A(\s13.dataOut [4]), .B(n6728), .C(\s01.dataOut [4]), .D(
        n6726), .Z(n6053) );
  CAN4X1 U6187 ( .A(n6056), .B(n6055), .C(n6054), .D(n6053), .Z(n6057) );
  CND4X1 U6188 ( .A(n6060), .B(n6059), .C(n6058), .D(n6057), .Z(n6061) );
  CMX2XL U6189 ( .A0(\m05.DinMast [4]), .A1(n6061), .S(n6748), .Z(n4198) );
  CIVX2 U6190 ( .A(\s08.dataOut [14]), .Z(n6763) );
  CNR2X1 U6191 ( .A(\m06.addrM [4]), .B(\m06.addrM [3]), .Z(n6112) );
  CNR2X1 U6192 ( .A(\m06.addrM [2]), .B(\m06.addrM [1]), .Z(n6092) );
  CND2X1 U6193 ( .A(n6112), .B(n6092), .Z(n6137) );
  CIVXL U6194 ( .A(\m06.addrM [7]), .Z(n6082) );
  CND2X1 U6195 ( .A(\m06.addrM [8]), .B(n6082), .Z(n6156) );
  CIVXL U6196 ( .A(\m06.addrM [6]), .Z(n6076) );
  CIVX2 U6197 ( .A(\m06.addrM [5]), .Z(n6126) );
  CND2X1 U6198 ( .A(n6076), .B(n6126), .Z(n6068) );
  CNR2X1 U6199 ( .A(n6156), .B(n6068), .Z(n6121) );
  CIVX2 U6200 ( .A(n6121), .Z(n6129) );
  CNR3XL U6201 ( .A(\m06.addrM [0]), .B(n6137), .C(n6129), .Z(n6064) );
  CNR2X1 U6202 ( .A(\m06.addrM [2]), .B(\m06.addrM [3]), .Z(n6062) );
  CIVX2 U6203 ( .A(\m06.addrM [4]), .Z(n6091) );
  CNR2X1 U6204 ( .A(\m06.addrM [7]), .B(\m06.addrM [8]), .Z(n6085) );
  CNR2X1 U6205 ( .A(n6076), .B(n6126), .Z(n6119) );
  CND2X1 U6206 ( .A(n6085), .B(n6119), .Z(n6099) );
  CIVX2 U6207 ( .A(\m06.addrM [8]), .Z(n7612) );
  CND2X1 U6208 ( .A(\m06.addrM [7]), .B(n7612), .Z(n6147) );
  COND4CX1 U6209 ( .A(n6062), .B(n6091), .C(n6099), .D(n6147), .Z(n6063) );
  CND2X1 U6210 ( .A(\m06.addrM [16]), .B(\m06.addrM [13]), .Z(n6078) );
  CNR3XL U6211 ( .A(\m06.addrM [14]), .B(\m06.addrM [15]), .C(n6078), .Z(n6107) );
  CIVXL U6212 ( .A(\m06.addrM [10]), .Z(n6086) );
  CIVXL U6213 ( .A(\m06.addrM [9]), .Z(n6115) );
  CND2X1 U6214 ( .A(n6086), .B(n6115), .Z(n6103) );
  CIVX2 U6215 ( .A(\m06.addrM [11]), .Z(n6102) );
  CND2X1 U6216 ( .A(\m06.addrM [12]), .B(n6102), .Z(n6114) );
  CNR2X1 U6217 ( .A(n6103), .B(n6114), .Z(n6071) );
  COND3X1 U6218 ( .A(n6064), .B(n6063), .C(n6107), .D(n6071), .Z(n6392) );
  CND2X1 U6219 ( .A(\m06.addrM [10]), .B(n6115), .Z(n6134) );
  CNR3XL U6220 ( .A(\m06.addrM [5]), .B(n6076), .C(n6156), .Z(n6138) );
  COND1XL U6221 ( .A(\m06.addrM [2]), .B(\m06.addrM [3]), .C(\m06.addrM [4]), 
        .Z(n6128) );
  CIVX2 U6222 ( .A(\m06.addrM [2]), .Z(n6369) );
  CND2X1 U6223 ( .A(\m06.addrM [4]), .B(\m06.addrM [3]), .Z(n6149) );
  CNR2X1 U6224 ( .A(n6369), .B(n6149), .Z(n6083) );
  CND3XL U6225 ( .A(n6083), .B(\m06.addrM [0]), .C(\m06.addrM [1]), .Z(n6110)
         );
  CANR3X1 U6226 ( .A(n6126), .B(n6110), .C(\m06.addrM [6]), .D(n6156), .Z(
        n6065) );
  CIVX2 U6227 ( .A(\m06.addrM [14]), .Z(n6070) );
  CND2X1 U6228 ( .A(\m06.addrM [15]), .B(n6070), .Z(n6075) );
  CNR3XL U6229 ( .A(\m06.addrM [16]), .B(\m06.addrM [13]), .C(n6075), .Z(n6116) );
  COND4CX1 U6230 ( .A(n6138), .B(n6128), .C(n6065), .D(n6116), .Z(n6066) );
  CNR3X1 U6231 ( .A(n6134), .B(n6114), .C(n6066), .Z(n7656) );
  CND2X1 U6232 ( .A(\m06.addrM [2]), .B(\m06.addrM [1]), .Z(n6067) );
  CND2X1 U6233 ( .A(n6112), .B(n6067), .Z(n6111) );
  CIVX2 U6234 ( .A(n6068), .Z(n6152) );
  CND2IX1 U6235 ( .B(n6147), .A(n6152), .Z(n6074) );
  CIVX2 U6236 ( .A(\m06.addrM [0]), .Z(n6144) );
  CNR2X1 U6237 ( .A(n6369), .B(n6144), .Z(n6113) );
  CIVX2 U6238 ( .A(n6067), .Z(n6146) );
  COND11X1 U6239 ( .A(n6113), .B(\m06.addrM [3]), .C(n6146), .D(\m06.addrM [4]), .Z(n6139) );
  CIVX2 U6240 ( .A(n6139), .Z(n6069) );
  COND1XL U6241 ( .A(n6069), .B(n6068), .C(n6085), .Z(n6073) );
  CIVX2 U6242 ( .A(n6078), .Z(n6093) );
  CNR2X1 U6243 ( .A(\m06.addrM [15]), .B(n6070), .Z(n6094) );
  CND2X1 U6244 ( .A(n6093), .B(n6094), .Z(n6135) );
  CND2IX1 U6245 ( .B(n6135), .A(n6071), .Z(n6072) );
  CANR4CX1 U6246 ( .A(n6111), .B(n6074), .C(n6073), .D(n6072), .Z(n7658) );
  CANR2XL U6247 ( .A(\s04.dataOut [14]), .B(n7656), .C(\s01.dataOut [14]), .D(
        n7658), .Z(n6165) );
  CNR3XL U6248 ( .A(\m06.addrM [12]), .B(n6075), .C(n6102), .Z(n6090) );
  CIVX2 U6249 ( .A(n6137), .Z(n6080) );
  CNR2X1 U6250 ( .A(n6076), .B(n6147), .Z(n6109) );
  CND2X1 U6251 ( .A(n6109), .B(n6126), .Z(n6098) );
  CNR2IX1 U6252 ( .B(n6119), .A(n6156), .Z(n6140) );
  CMXI2X1 U6253 ( .A0(n6156), .A1(n6147), .S(n6119), .Z(n6077) );
  CANR4CX1 U6254 ( .A(n6092), .B(n6149), .C(n6140), .D(n6077), .Z(n6079) );
  CANR4CX1 U6255 ( .A(n6080), .B(n6098), .C(n6079), .D(n6078), .Z(n6081) );
  CAN4X1 U6256 ( .A(n6090), .B(\m06.addrM [9]), .C(n6081), .D(n6086), .Z(n7665) );
  CNR2IX1 U6257 ( .B(\m06.addrM [16]), .A(\m06.addrM [13]), .Z(n6095) );
  CNR2X1 U6258 ( .A(n6082), .B(n7612), .Z(n6153) );
  COND3X1 U6259 ( .A(\m06.addrM [5]), .B(n6083), .C(\m06.addrM [6]), .D(n6153), 
        .Z(n6088) );
  CNR2X1 U6260 ( .A(\m06.addrM [6]), .B(n6147), .Z(n6105) );
  CANR4CX1 U6261 ( .A(\m06.addrM [0]), .B(\m06.addrM [1]), .C(n6083), .D(n6098), .Z(n6084) );
  COND11X1 U6262 ( .A(n6105), .B(n6085), .C(n6084), .D(\m06.addrM [9]), .Z(
        n6087) );
  CANR4CX1 U6263 ( .A(\m06.addrM [9]), .B(n6088), .C(n6087), .D(n6086), .Z(
        n6089) );
  CND3XL U6264 ( .A(n6095), .B(n6090), .C(n6089), .Z(n6677) );
  CIVX2 U6265 ( .A(n6677), .Z(n7678) );
  CNR2X1 U6266 ( .A(n6119), .B(n6156), .Z(n6127) );
  CND2X1 U6267 ( .A(\m06.addrM [12]), .B(\m06.addrM [11]), .Z(n6096) );
  CNR2X1 U6268 ( .A(n6134), .B(n6096), .Z(n6122) );
  CIVX2 U6269 ( .A(n7550), .Z(n7667) );
  CAOR2X2 U6270 ( .A(n7678), .B(\s00.dataOut [14]), .C(\s07.dataOut [14]), .D(
        n7667), .Z(n6163) );
  CANR1XL U6271 ( .A(\m06.addrM [3]), .B(n6146), .C(\m06.addrM [4]), .Z(n6120)
         );
  CND2X1 U6272 ( .A(n6095), .B(n6094), .Z(n6155) );
  COR4X1 U6273 ( .A(n6120), .B(n6103), .C(n6096), .D(n6155), .Z(n6097) );
  CNR2X1 U6274 ( .A(n6098), .B(n6097), .Z(n7660) );
  CANR1XL U6275 ( .A(\m06.addrM [2]), .B(\m06.addrM [3]), .C(\m06.addrM [4]), 
        .Z(n6101) );
  CIVX2 U6276 ( .A(n6099), .Z(n6100) );
  CANR2X1 U6277 ( .A(n6101), .B(n6121), .C(n6100), .D(n6111), .Z(n6104) );
  CND2IX1 U6278 ( .B(\m06.addrM [12]), .A(n6102), .Z(n6133) );
  COR2X1 U6279 ( .A(n6103), .B(n6133), .Z(n6154) );
  CANR3X1 U6280 ( .A(n6104), .B(n6147), .C(n6135), .D(n6154), .Z(n7661) );
  CANR2X1 U6281 ( .A(\s02.dataOut [14]), .B(n7660), .C(\s13.dataOut [14]), .D(
        n7661), .Z(n6161) );
  COND3X1 U6282 ( .A(n6113), .B(n6111), .C(\m06.addrM [5]), .D(n6105), .Z(
        n6106) );
  COND4CX1 U6283 ( .A(n6119), .B(n6137), .C(n6156), .D(n6106), .Z(n6108) );
  COND3X1 U6284 ( .A(n6109), .B(n6108), .C(n6122), .D(n6107), .Z(n6651) );
  CIVX2 U6285 ( .A(n6651), .Z(n7663) );
  CANR2X1 U6286 ( .A(n6113), .B(n6112), .C(n6111), .D(n6110), .Z(n6118) );
  CNR3XL U6287 ( .A(\m06.addrM [10]), .B(n6115), .C(n6114), .Z(n6141) );
  CND4X1 U6288 ( .A(n6153), .B(n6119), .C(n6141), .D(n6116), .Z(n6117) );
  CNR2X1 U6289 ( .A(n6118), .B(n6117), .Z(n7657) );
  CANR2X1 U6290 ( .A(n7663), .B(\s03.dataOut [14]), .C(\s05.dataOut [14]), .D(
        n7657), .Z(n6160) );
  CND2IX1 U6291 ( .B(n6120), .A(n6119), .Z(n6124) );
  CND3XL U6292 ( .A(\m06.addrM [4]), .B(n6121), .C(\m06.addrM [1]), .Z(n6130)
         );
  COND4CX1 U6293 ( .A(n6152), .B(n6128), .C(n6156), .D(n6130), .Z(n6123) );
  COND4CX1 U6294 ( .A(n6153), .B(n6124), .C(n6123), .D(n6122), .Z(n6125) );
  CNR2X1 U6295 ( .A(n6135), .B(n6125), .Z(n7666) );
  CNR2IX1 U6296 ( .B(n6127), .A(n6126), .Z(n6132) );
  COND2X1 U6297 ( .A(n6144), .B(n6130), .C(n6129), .D(n6128), .Z(n6131) );
  CANR3X1 U6298 ( .A(n6138), .B(n6139), .C(n6132), .D(n6131), .Z(n6136) );
  CNR4X1 U6299 ( .A(n6136), .B(n6135), .C(n6134), .D(n6133), .Z(n6698) );
  CANR2XL U6300 ( .A(\s09.dataOut [14]), .B(n7666), .C(\s10.dataOut [14]), .D(
        n6698), .Z(n6159) );
  CANR2X1 U6301 ( .A(n6140), .B(n6139), .C(n6138), .D(n6137), .Z(n6143) );
  CIVX2 U6302 ( .A(n6141), .Z(n6142) );
  CNR3X1 U6303 ( .A(n6143), .B(n6155), .C(n6142), .Z(n7659) );
  CNR2IX1 U6304 ( .B(\m06.addrM [1]), .A(n6144), .Z(n6145) );
  CANR4CX1 U6305 ( .A(\m06.addrM [2]), .B(n6145), .C(\m06.addrM [3]), .D(
        \m06.addrM [4]), .Z(n6151) );
  CND2X1 U6306 ( .A(\m06.addrM [4]), .B(n6146), .Z(n6148) );
  CANR11X1 U6307 ( .A(n6152), .B(n6149), .C(n6148), .D(n6147), .Z(n6150) );
  CANR11X1 U6308 ( .A(n6153), .B(n6152), .C(n6151), .D(n6150), .Z(n6157) );
  CANR3X1 U6309 ( .A(n6157), .B(n6156), .C(n6155), .D(n6154), .Z(n7664) );
  CANR2XL U6310 ( .A(\s06.dataOut [14]), .B(n7659), .C(\s11.dataOut [14]), .D(
        n7664), .Z(n6158) );
  CND4X1 U6311 ( .A(n6161), .B(n6160), .C(n6159), .D(n6158), .Z(n6162) );
  CANR3X1 U6312 ( .A(\s12.dataOut [14]), .B(n7665), .C(n6163), .D(n6162), .Z(
        n6164) );
  COND3X1 U6313 ( .A(n6763), .B(n6392), .C(n6165), .D(n6164), .Z(n6178) );
  CIVX2 U6314 ( .A(n7657), .Z(n6332) );
  CIVX2 U6315 ( .A(n7656), .Z(n7576) );
  CIVX2 U6316 ( .A(n7660), .Z(n6626) );
  CIVX2 U6317 ( .A(n7665), .Z(n7514) );
  CIVX2 U6318 ( .A(n7664), .Z(n6493) );
  CIVX2 U6319 ( .A(n7658), .Z(n6579) );
  CIVXL U6320 ( .A(n7661), .Z(n6686) );
  CIVX2 U6321 ( .A(n7666), .Z(n6418) );
  CNR4XL U6322 ( .A(\m06.addrM [42]), .B(\m06.addrM [43]), .C(\m06.addrM [44]), 
        .D(\m06.addrM [45]), .Z(n6177) );
  CNR4XL U6323 ( .A(\m06.addrM [38]), .B(\m06.addrM [39]), .C(\m06.addrM [40]), 
        .D(\m06.addrM [41]), .Z(n6176) );
  CAN4X1 U6324 ( .A(\m06.addrM [20]), .B(\m06.addrM [19]), .C(\m06.addrM [23]), 
        .D(\m06.addrM [22]), .Z(n6166) );
  CND3XL U6325 ( .A(\m06.addrM [18]), .B(\m06.addrM [17]), .C(n6166), .Z(n6174) );
  CNR2XL U6326 ( .A(\m05.YouGotIt ), .B(n6167), .Z(n7618) );
  CND2XL U6327 ( .A(n7618), .B(\m06.YouGotIt ), .Z(n7613) );
  COR4X1 U6328 ( .A(\m06.addrM [26]), .B(\m06.addrM [27]), .C(\m06.addrM [28]), 
        .D(\m06.addrM [29]), .Z(n6172) );
  COR4X1 U6329 ( .A(\m06.addrM [30]), .B(\m06.addrM [31]), .C(\m06.addrM [32]), 
        .D(\m06.addrM [33]), .Z(n6171) );
  CNR4X1 U6330 ( .A(\m06.addrM [34]), .B(\m06.addrM [35]), .C(\m06.addrM [36]), 
        .D(\m06.addrM [37]), .Z(n6169) );
  CNR2X1 U6331 ( .A(\m06.addrM [24]), .B(\m06.addrM [25]), .Z(n6168) );
  CND3XL U6332 ( .A(\m06.addrM [21]), .B(n6169), .C(n6168), .Z(n6170) );
  COR4X1 U6333 ( .A(n7613), .B(n6172), .C(n6171), .D(n6170), .Z(n6173) );
  CNR4X1 U6334 ( .A(\m06.addrM [46]), .B(\m06.addrM [47]), .C(n6174), .D(n6173), .Z(n6175) );
  CND3X1 U6335 ( .A(n6177), .B(n6176), .C(n6175), .Z(n7577) );
  CMX2XL U6336 ( .A0(\m06.DinMast [14]), .A1(n6178), .S(n7679), .Z(n5200) );
  CIVX2 U6337 ( .A(\s07.dataOut [13]), .Z(n7485) );
  CANR2XL U6338 ( .A(\s11.dataOut [13]), .B(n7664), .C(\s01.dataOut [13]), .D(
        n7658), .Z(n6186) );
  CIVX2 U6339 ( .A(n6392), .Z(n7662) );
  CAOR2X2 U6340 ( .A(\s04.dataOut [13]), .B(n7656), .C(\s08.dataOut [13]), .D(
        n7662), .Z(n6184) );
  CANR2X1 U6341 ( .A(\s05.dataOut [13]), .B(n7657), .C(\s13.dataOut [13]), .D(
        n7661), .Z(n6182) );
  CANR2X1 U6342 ( .A(n7663), .B(\s03.dataOut [13]), .C(\s02.dataOut [13]), .D(
        n7660), .Z(n6181) );
  CANR2XL U6343 ( .A(\s09.dataOut [13]), .B(n7666), .C(\s10.dataOut [13]), .D(
        n6698), .Z(n6180) );
  CANR2X1 U6344 ( .A(\s12.dataOut [13]), .B(n7665), .C(\s06.dataOut [13]), .D(
        n7659), .Z(n6179) );
  CND4X1 U6345 ( .A(n6182), .B(n6181), .C(n6180), .D(n6179), .Z(n6183) );
  CANR3X1 U6346 ( .A(n7678), .B(\s00.dataOut [13]), .C(n6184), .D(n6183), .Z(
        n6185) );
  COND3X1 U6347 ( .A(n7485), .B(n7550), .C(n6186), .D(n6185), .Z(n6187) );
  CMX2XL U6348 ( .A0(\m06.DinMast [13]), .A1(n6187), .S(n7679), .Z(n5199) );
  CIVX2 U6349 ( .A(\s04.dataOut [12]), .Z(n7503) );
  CANR2XL U6350 ( .A(n7663), .B(\s03.dataOut [12]), .C(\s01.dataOut [12]), .D(
        n7658), .Z(n6195) );
  CAOR2X2 U6351 ( .A(n7678), .B(\s00.dataOut [12]), .C(\s07.dataOut [12]), .D(
        n7667), .Z(n6193) );
  CANR2X1 U6352 ( .A(\s05.dataOut [12]), .B(n7657), .C(\s13.dataOut [12]), .D(
        n7661), .Z(n6191) );
  CANR2X1 U6353 ( .A(\s02.dataOut [12]), .B(n7660), .C(\s08.dataOut [12]), .D(
        n7662), .Z(n6190) );
  CANR2XL U6354 ( .A(\s11.dataOut [12]), .B(n7664), .C(\s10.dataOut [12]), .D(
        n6698), .Z(n6189) );
  CANR2X1 U6355 ( .A(\s12.dataOut [12]), .B(n7665), .C(\s09.dataOut [12]), .D(
        n7666), .Z(n6188) );
  CND4X1 U6356 ( .A(n6191), .B(n6190), .C(n6189), .D(n6188), .Z(n6192) );
  CANR3XL U6357 ( .A(\s06.dataOut [12]), .B(n7659), .C(n6193), .D(n6192), .Z(
        n6194) );
  COND3X1 U6358 ( .A(n7503), .B(n7576), .C(n6195), .D(n6194), .Z(n6196) );
  CMX2XL U6359 ( .A0(\m06.DinMast [12]), .A1(n6196), .S(n7679), .Z(n5198) );
  CIVX2 U6360 ( .A(\s05.dataOut [11]), .Z(n6205) );
  CANR2XL U6361 ( .A(\s13.dataOut [11]), .B(n7661), .C(\s01.dataOut [11]), .D(
        n7658), .Z(n6204) );
  CAOR2X2 U6362 ( .A(n7678), .B(\s00.dataOut [11]), .C(\s09.dataOut [11]), .D(
        n7666), .Z(n6202) );
  CANR2X1 U6363 ( .A(n7663), .B(\s03.dataOut [11]), .C(\s02.dataOut [11]), .D(
        n7660), .Z(n6200) );
  CANR2X1 U6364 ( .A(\s04.dataOut [11]), .B(n7656), .C(\s08.dataOut [11]), .D(
        n7662), .Z(n6199) );
  CANR2XL U6365 ( .A(\s07.dataOut [11]), .B(n7667), .C(\s10.dataOut [11]), .D(
        n6698), .Z(n6198) );
  CANR2XL U6366 ( .A(\s12.dataOut [11]), .B(n7665), .C(\s11.dataOut [11]), .D(
        n7664), .Z(n6197) );
  CND4X1 U6367 ( .A(n6200), .B(n6199), .C(n6198), .D(n6197), .Z(n6201) );
  CANR3XL U6368 ( .A(\s06.dataOut [11]), .B(n7659), .C(n6202), .D(n6201), .Z(
        n6203) );
  COND3X1 U6369 ( .A(n6205), .B(n6332), .C(n6204), .D(n6203), .Z(n6206) );
  CMX2XL U6370 ( .A0(\m06.DinMast [11]), .A1(n6206), .S(n7679), .Z(n5197) );
  CIVX2 U6371 ( .A(\s07.dataOut [15]), .Z(n7438) );
  CANR2XL U6372 ( .A(\s10.dataOut [15]), .B(n6698), .C(\s01.dataOut [15]), .D(
        n7658), .Z(n6214) );
  CAOR2X2 U6373 ( .A(n7678), .B(\s00.dataOut [15]), .C(\s08.dataOut [15]), .D(
        n7662), .Z(n6212) );
  CANR2X1 U6374 ( .A(n7663), .B(\s03.dataOut [15]), .C(\s04.dataOut [15]), .D(
        n7656), .Z(n6210) );
  CANR2X1 U6375 ( .A(\s02.dataOut [15]), .B(n7660), .C(\s13.dataOut [15]), .D(
        n7661), .Z(n6209) );
  CANR2XL U6376 ( .A(\s06.dataOut [15]), .B(n7659), .C(\s12.dataOut [15]), .D(
        n7665), .Z(n6208) );
  CANR2XL U6377 ( .A(\s09.dataOut [15]), .B(n7666), .C(\s11.dataOut [15]), .D(
        n7664), .Z(n6207) );
  CND4X1 U6378 ( .A(n6210), .B(n6209), .C(n6208), .D(n6207), .Z(n6211) );
  CANR3X1 U6379 ( .A(\s05.dataOut [15]), .B(n7657), .C(n6212), .D(n6211), .Z(
        n6213) );
  COND3X1 U6380 ( .A(n7438), .B(n7550), .C(n6214), .D(n6213), .Z(n6215) );
  CMX2XL U6381 ( .A0(\m06.DinMast [15]), .A1(n6215), .S(n7679), .Z(n5201) );
  CIVX2 U6382 ( .A(\s00.dataOut [10]), .Z(n6224) );
  CANR2X1 U6383 ( .A(n7663), .B(\s03.dataOut [10]), .C(\s05.dataOut [10]), .D(
        n7657), .Z(n6223) );
  CAOR2XL U6384 ( .A(\s07.dataOut [10]), .B(n7667), .C(\s01.dataOut [10]), .D(
        n7658), .Z(n6221) );
  CANR2X1 U6385 ( .A(\s04.dataOut [10]), .B(n7656), .C(\s13.dataOut [10]), .D(
        n7661), .Z(n6219) );
  CANR2X1 U6386 ( .A(\s02.dataOut [10]), .B(n7660), .C(\s08.dataOut [10]), .D(
        n7662), .Z(n6218) );
  CANR2XL U6387 ( .A(\s06.dataOut [10]), .B(n7659), .C(\s11.dataOut [10]), .D(
        n7664), .Z(n6217) );
  CANR2XL U6388 ( .A(\s12.dataOut [10]), .B(n7665), .C(\s10.dataOut [10]), .D(
        n6698), .Z(n6216) );
  CND4X1 U6389 ( .A(n6219), .B(n6218), .C(n6217), .D(n6216), .Z(n6220) );
  CANR3X1 U6390 ( .A(\s09.dataOut [10]), .B(n7666), .C(n6221), .D(n6220), .Z(
        n6222) );
  COND3X1 U6391 ( .A(n6677), .B(n6224), .C(n6223), .D(n6222), .Z(n6225) );
  CMX2XL U6392 ( .A0(\m06.DinMast [10]), .A1(n6225), .S(n7679), .Z(n5196) );
  CIVX2 U6393 ( .A(\s05.dataOut [0]), .Z(n7326) );
  CANR2X1 U6394 ( .A(\s04.dataOut [0]), .B(n7656), .C(\s01.dataOut [0]), .D(
        n7658), .Z(n6233) );
  CAOR2X2 U6395 ( .A(\s07.dataOut [0]), .B(n7667), .C(\s09.dataOut [0]), .D(
        n7666), .Z(n6231) );
  CANR2X1 U6396 ( .A(\s02.dataOut [0]), .B(n7660), .C(\s08.dataOut [0]), .D(
        n7662), .Z(n6229) );
  CANR2XL U6397 ( .A(n7663), .B(\s03.dataOut [0]), .C(\s13.dataOut [0]), .D(
        n7661), .Z(n6228) );
  CANR2XL U6398 ( .A(\s06.dataOut [0]), .B(n7659), .C(\s10.dataOut [0]), .D(
        n6698), .Z(n6227) );
  CANR2XL U6399 ( .A(\s12.dataOut [0]), .B(n7665), .C(\s11.dataOut [0]), .D(
        n7664), .Z(n6226) );
  CND4X1 U6400 ( .A(n6229), .B(n6228), .C(n6227), .D(n6226), .Z(n6230) );
  CANR3X1 U6401 ( .A(n7678), .B(\s00.dataOut [0]), .C(n6231), .D(n6230), .Z(
        n6232) );
  COND3X1 U6402 ( .A(n7326), .B(n6332), .C(n6233), .D(n6232), .Z(n6234) );
  CMX2XL U6403 ( .A0(\m06.DinMast [0]), .A1(n6234), .S(n7679), .Z(n5186) );
  CIVX2 U6404 ( .A(\s03.dataOut [1]), .Z(n7340) );
  CANR2XL U6405 ( .A(n7678), .B(\s00.dataOut [1]), .C(\s13.dataOut [1]), .D(
        n7661), .Z(n6242) );
  CAOR2XL U6406 ( .A(\s10.dataOut [1]), .B(n6698), .C(\s01.dataOut [1]), .D(
        n7658), .Z(n6240) );
  CANR2X1 U6407 ( .A(\s04.dataOut [1]), .B(n7656), .C(\s02.dataOut [1]), .D(
        n7660), .Z(n6238) );
  CANR2X1 U6408 ( .A(\s05.dataOut [1]), .B(n7657), .C(\s08.dataOut [1]), .D(
        n7662), .Z(n6237) );
  CANR2XL U6409 ( .A(\s06.dataOut [1]), .B(n7659), .C(\s09.dataOut [1]), .D(
        n7666), .Z(n6236) );
  CANR2X1 U6410 ( .A(\s07.dataOut [1]), .B(n7667), .C(\s12.dataOut [1]), .D(
        n7665), .Z(n6235) );
  CND4X1 U6411 ( .A(n6238), .B(n6237), .C(n6236), .D(n6235), .Z(n6239) );
  CANR3XL U6412 ( .A(\s11.dataOut [1]), .B(n7664), .C(n6240), .D(n6239), .Z(
        n6241) );
  COND3X1 U6413 ( .A(n6651), .B(n7340), .C(n6242), .D(n6241), .Z(n6243) );
  CMX2XL U6414 ( .A0(\m06.DinMast [1]), .A1(n6243), .S(n7679), .Z(n5187) );
  CIVX2 U6415 ( .A(\s04.dataOut [2]), .Z(n6253) );
  CANR2XL U6416 ( .A(\s13.dataOut [2]), .B(n7661), .C(\s01.dataOut [2]), .D(
        n7658), .Z(n6252) );
  CIVX2 U6417 ( .A(\s00.dataOut [2]), .Z(n7353) );
  CIVXL U6418 ( .A(n6698), .Z(n7674) );
  COND2X1 U6419 ( .A(n6677), .B(n7353), .C(n6244), .D(n7674), .Z(n6250) );
  CANR2X1 U6420 ( .A(\s05.dataOut [2]), .B(n7657), .C(\s08.dataOut [2]), .D(
        n7662), .Z(n6248) );
  CANR2X1 U6421 ( .A(n7663), .B(\s03.dataOut [2]), .C(\s02.dataOut [2]), .D(
        n7660), .Z(n6247) );
  CANR2XL U6422 ( .A(\s06.dataOut [2]), .B(n7659), .C(\s07.dataOut [2]), .D(
        n7667), .Z(n6246) );
  CANR2XL U6423 ( .A(\s11.dataOut [2]), .B(n7664), .C(\s09.dataOut [2]), .D(
        n7666), .Z(n6245) );
  CND4X1 U6424 ( .A(n6248), .B(n6247), .C(n6246), .D(n6245), .Z(n6249) );
  CANR3X1 U6425 ( .A(\s12.dataOut [2]), .B(n7665), .C(n6250), .D(n6249), .Z(
        n6251) );
  COND3X1 U6426 ( .A(n6253), .B(n7576), .C(n6252), .D(n6251), .Z(n6254) );
  CMX2XL U6427 ( .A0(\m06.DinMast [2]), .A1(n6254), .S(n7679), .Z(n5188) );
  CIVX2 U6428 ( .A(\s05.dataOut [3]), .Z(n7363) );
  CANR2XL U6429 ( .A(n7663), .B(\s03.dataOut [3]), .C(\s01.dataOut [3]), .D(
        n7658), .Z(n6262) );
  CAOR2XL U6430 ( .A(\s12.dataOut [3]), .B(n7665), .C(\s11.dataOut [3]), .D(
        n7664), .Z(n6260) );
  CANR2X1 U6431 ( .A(\s02.dataOut [3]), .B(n7660), .C(\s08.dataOut [3]), .D(
        n7662), .Z(n6258) );
  CANR2XL U6432 ( .A(\s04.dataOut [3]), .B(n7656), .C(\s13.dataOut [3]), .D(
        n7661), .Z(n6257) );
  CANR2X1 U6433 ( .A(\s07.dataOut [3]), .B(n7667), .C(\s09.dataOut [3]), .D(
        n7666), .Z(n6256) );
  CANR2XL U6434 ( .A(\s06.dataOut [3]), .B(n7659), .C(\s10.dataOut [3]), .D(
        n6698), .Z(n6255) );
  CND4X1 U6435 ( .A(n6258), .B(n6257), .C(n6256), .D(n6255), .Z(n6259) );
  CANR3X1 U6436 ( .A(n7678), .B(\s00.dataOut [3]), .C(n6260), .D(n6259), .Z(
        n6261) );
  COND3X1 U6437 ( .A(n7363), .B(n6332), .C(n6262), .D(n6261), .Z(n6263) );
  CMX2XL U6438 ( .A0(\m06.DinMast [3]), .A1(n6263), .S(n7679), .Z(n5189) );
  CIVX2 U6439 ( .A(\s05.dataOut [4]), .Z(n6272) );
  CANR2XL U6440 ( .A(\s13.dataOut [4]), .B(n7661), .C(\s01.dataOut [4]), .D(
        n7658), .Z(n6271) );
  CAOR2XL U6441 ( .A(n7678), .B(\s00.dataOut [4]), .C(\s10.dataOut [4]), .D(
        n6698), .Z(n6269) );
  CANR2X1 U6442 ( .A(\s02.dataOut [4]), .B(n7660), .C(\s08.dataOut [4]), .D(
        n7662), .Z(n6267) );
  CANR2X1 U6443 ( .A(n7663), .B(\s03.dataOut [4]), .C(\s04.dataOut [4]), .D(
        n7656), .Z(n6266) );
  CANR2XL U6444 ( .A(\s06.dataOut [4]), .B(n7659), .C(\s12.dataOut [4]), .D(
        n7665), .Z(n6265) );
  CANR2XL U6445 ( .A(\s09.dataOut [4]), .B(n7666), .C(\s11.dataOut [4]), .D(
        n7664), .Z(n6264) );
  CND4X1 U6446 ( .A(n6267), .B(n6266), .C(n6265), .D(n6264), .Z(n6268) );
  CANR3X1 U6447 ( .A(\s07.dataOut [4]), .B(n7667), .C(n6269), .D(n6268), .Z(
        n6270) );
  COND3X1 U6448 ( .A(n6272), .B(n6332), .C(n6271), .D(n6270), .Z(n6273) );
  CMX2XL U6449 ( .A0(\m06.DinMast [4]), .A1(n6273), .S(n7679), .Z(n5190) );
  CIVX2 U6450 ( .A(\s04.dataOut [5]), .Z(n6282) );
  CANR2XL U6451 ( .A(\s13.dataOut [5]), .B(n7661), .C(\s01.dataOut [5]), .D(
        n7658), .Z(n6281) );
  CIVX2 U6452 ( .A(\s00.dataOut [5]), .Z(n7383) );
  CIVX2 U6453 ( .A(\s07.dataOut [5]), .Z(n7385) );
  COND2X1 U6454 ( .A(n6677), .B(n7383), .C(n7385), .D(n7550), .Z(n6279) );
  CANR2X1 U6455 ( .A(\s02.dataOut [5]), .B(n7660), .C(\s08.dataOut [5]), .D(
        n7662), .Z(n6277) );
  CANR2X1 U6456 ( .A(n7663), .B(\s03.dataOut [5]), .C(\s05.dataOut [5]), .D(
        n7657), .Z(n6276) );
  CANR2XL U6457 ( .A(\s10.dataOut [5]), .B(n6698), .C(\s11.dataOut [5]), .D(
        n7664), .Z(n6275) );
  CANR2XL U6458 ( .A(\s06.dataOut [5]), .B(n7659), .C(\s12.dataOut [5]), .D(
        n7665), .Z(n6274) );
  CND4X1 U6459 ( .A(n6277), .B(n6276), .C(n6275), .D(n6274), .Z(n6278) );
  CANR3X1 U6460 ( .A(\s09.dataOut [5]), .B(n7666), .C(n6279), .D(n6278), .Z(
        n6280) );
  COND3X1 U6461 ( .A(n6282), .B(n7576), .C(n6281), .D(n6280), .Z(n6283) );
  CMX2XL U6462 ( .A0(\m06.DinMast [5]), .A1(n6283), .S(n7679), .Z(n5191) );
  CND2XL U6463 ( .A(\m01.YouGotIt ), .B(n7690), .Z(n7561) );
  CIVX2 U6464 ( .A(n7561), .Z(n7642) );
  CANR2XL U6465 ( .A(\m00.YouGotIt ), .B(\m00.addrM [1]), .C(\m01.addrM [1]), 
        .D(n7642), .Z(n6290) );
  CND2IXL U6466 ( .B(n6284), .A(\m03.YouGotIt ), .Z(n7566) );
  CIVX2 U6467 ( .A(n7566), .Z(n7644) );
  CIVX2 U6468 ( .A(n7564), .Z(n7643) );
  CANR2X1 U6469 ( .A(\m03.addrM [1]), .B(n7644), .C(\m02.addrM [1]), .D(n7643), 
        .Z(n6289) );
  CIVX2 U6470 ( .A(n6285), .Z(n7641) );
  CIVX2 U6471 ( .A(n7613), .Z(n7640) );
  CANR2X1 U6472 ( .A(\m05.addrM [1]), .B(n7641), .C(n7640), .D(\m06.addrM [1]), 
        .Z(n6288) );
  CND2XL U6473 ( .A(\m04.YouGotIt ), .B(n6286), .Z(n7616) );
  CIVX2 U6474 ( .A(n7616), .Z(n7648) );
  CND2X1 U6475 ( .A(\m04.addrM [1]), .B(n7648), .Z(n6287) );
  CND4X1 U6476 ( .A(n6290), .B(n6289), .C(n6288), .D(n6287), .Z(n7687) );
  CNR4XL U6477 ( .A(\m03.addrM [34]), .B(\m03.addrM [35]), .C(\m03.addrM [36]), 
        .D(\m03.addrM [37]), .Z(n6301) );
  CNR4XL U6478 ( .A(\m03.addrM [30]), .B(\m03.addrM [31]), .C(\m03.addrM [32]), 
        .D(\m03.addrM [33]), .Z(n6300) );
  CAN4X1 U6479 ( .A(\m03.addrM [17]), .B(\m03.addrM [20]), .C(\m03.addrM [21]), 
        .D(\m03.addrM [19]), .Z(n6291) );
  CND3XL U6480 ( .A(\m03.addrM [23]), .B(\m03.addrM [18]), .C(n6291), .Z(n6298) );
  COR4X1 U6481 ( .A(\m03.addrM [42]), .B(\m03.addrM [43]), .C(\m03.addrM [44]), 
        .D(\m03.addrM [45]), .Z(n6296) );
  COR4X1 U6482 ( .A(\m03.addrM [38]), .B(\m03.addrM [39]), .C(\m03.addrM [40]), 
        .D(\m03.addrM [41]), .Z(n6295) );
  CNR4X1 U6483 ( .A(\m03.addrM [26]), .B(\m03.addrM [27]), .C(\m03.addrM [28]), 
        .D(\m03.addrM [29]), .Z(n6293) );
  CNR2X1 U6484 ( .A(\m03.addrM [24]), .B(\m03.addrM [25]), .Z(n6292) );
  CND3XL U6485 ( .A(\m03.addrM [22]), .B(n6293), .C(n6292), .Z(n6294) );
  COR4X1 U6486 ( .A(n6296), .B(n6295), .C(n7566), .D(n6294), .Z(n6297) );
  CNR4X1 U6487 ( .A(\m03.addrM [46]), .B(\m03.addrM [47]), .C(n6298), .D(n6297), .Z(n6299) );
  CND3XL U6488 ( .A(n6301), .B(n6300), .C(n6299), .Z(n7575) );
  CIVX2 U6489 ( .A(n7575), .Z(n7560) );
  CIVX2 U6490 ( .A(\m03.addrM [6]), .Z(n7567) );
  CND2X1 U6491 ( .A(\m03.addrM [7]), .B(\m03.addrM [8]), .Z(n6419) );
  CNR2X1 U6492 ( .A(n7567), .B(n6419), .Z(n6530) );
  CND2X1 U6493 ( .A(\m03.addrM [5]), .B(n6530), .Z(n6307) );
  CIVXL U6494 ( .A(\m03.addrM [10]), .Z(n6424) );
  CND2X1 U6495 ( .A(\m03.addrM [9]), .B(n6424), .Z(n7308) );
  CIVX2 U6496 ( .A(\m03.addrM [2]), .Z(n6385) );
  CIVX2 U6497 ( .A(\m03.addrM [1]), .Z(n7303) );
  CNR2X1 U6498 ( .A(n6385), .B(n7303), .Z(n6614) );
  CIVX2 U6499 ( .A(\m03.addrM [3]), .Z(n6635) );
  CIVX2 U6500 ( .A(\m03.addrM [4]), .Z(n6634) );
  CND2X1 U6501 ( .A(n6635), .B(n6634), .Z(n6302) );
  CNR2X1 U6502 ( .A(n6614), .B(n6302), .Z(n6585) );
  CND2X1 U6503 ( .A(\m03.addrM [2]), .B(\m03.addrM [0]), .Z(n6448) );
  CND2X1 U6504 ( .A(n6585), .B(n6448), .Z(n6638) );
  CNR2X1 U6505 ( .A(\m03.addrM [2]), .B(\m03.addrM [1]), .Z(n6636) );
  COND1XL U6506 ( .A(n6636), .B(n6635), .C(n6634), .Z(n7301) );
  CIVX2 U6507 ( .A(n7301), .Z(n6305) );
  CND2X1 U6508 ( .A(\m03.addrM [1]), .B(\m03.addrM [0]), .Z(n7289) );
  CIVX2 U6509 ( .A(n7289), .Z(n6449) );
  COND1XL U6510 ( .A(n6385), .B(n6634), .C(\m03.addrM [3]), .Z(n6303) );
  COND4CX1 U6511 ( .A(\m03.addrM [3]), .B(n6449), .C(n6634), .D(n6303), .Z(
        n6304) );
  CNR2X1 U6512 ( .A(\m03.addrM [13]), .B(\m03.addrM [14]), .Z(n6535) );
  CIVXL U6513 ( .A(\m03.addrM [12]), .Z(n6527) );
  CNR2X1 U6514 ( .A(\m03.addrM [11]), .B(n6527), .Z(n7310) );
  CIVXL U6515 ( .A(\m03.addrM [16]), .Z(n6388) );
  CAN4X1 U6516 ( .A(\m03.addrM [15]), .B(n6535), .C(n7310), .D(n6388), .Z(
        n7293) );
  COND4CX1 U6517 ( .A(n6638), .B(n6305), .C(n6304), .D(n7293), .Z(n6306) );
  CNR3X1 U6518 ( .A(n6307), .B(n7308), .C(n6306), .Z(n7497) );
  CNR4X1 U6519 ( .A(\m04.addrM [42]), .B(\m04.addrM [43]), .C(\m04.addrM [44]), 
        .D(\m04.addrM [45]), .Z(n6318) );
  CNR4X1 U6520 ( .A(\m04.addrM [38]), .B(\m04.addrM [39]), .C(\m04.addrM [40]), 
        .D(\m04.addrM [41]), .Z(n6317) );
  CAN4X1 U6521 ( .A(\m04.addrM [20]), .B(\m04.addrM [19]), .C(\m04.addrM [23]), 
        .D(\m04.addrM [22]), .Z(n6308) );
  CND3XL U6522 ( .A(\m04.addrM [18]), .B(\m04.addrM [17]), .C(n6308), .Z(n6315) );
  COR4X1 U6523 ( .A(\m04.addrM [26]), .B(\m04.addrM [27]), .C(\m04.addrM [28]), 
        .D(\m04.addrM [29]), .Z(n6313) );
  COR4X1 U6524 ( .A(\m04.addrM [30]), .B(\m04.addrM [31]), .C(\m04.addrM [32]), 
        .D(\m04.addrM [33]), .Z(n6312) );
  CNR4X1 U6525 ( .A(\m04.addrM [34]), .B(\m04.addrM [35]), .C(\m04.addrM [36]), 
        .D(\m04.addrM [37]), .Z(n6310) );
  CNR2X1 U6526 ( .A(\m04.addrM [24]), .B(\m04.addrM [25]), .Z(n6309) );
  CND3XL U6527 ( .A(\m04.addrM [21]), .B(n6310), .C(n6309), .Z(n6311) );
  COR4X1 U6528 ( .A(n7616), .B(n6313), .C(n6312), .D(n6311), .Z(n6314) );
  CNR4X1 U6529 ( .A(\m04.addrM [46]), .B(\m04.addrM [47]), .C(n6315), .D(n6314), .Z(n6316) );
  CND3X1 U6530 ( .A(n6318), .B(n6317), .C(n6316), .Z(n7539) );
  CIVX2 U6531 ( .A(\m04.addrM [5]), .Z(n6845) );
  CIVXL U6532 ( .A(\m04.addrM [8]), .Z(n7617) );
  CNR2IX1 U6533 ( .B(\m04.addrM [7]), .A(n7617), .Z(n6488) );
  CND2X1 U6534 ( .A(\m04.addrM [6]), .B(n6488), .Z(n6543) );
  CNR2X1 U6535 ( .A(n6845), .B(n6543), .Z(n6324) );
  CIVX2 U6536 ( .A(\m04.addrM [9]), .Z(n6805) );
  CIVX2 U6537 ( .A(\m04.addrM [11]), .Z(n6537) );
  CND2X1 U6538 ( .A(n6537), .B(\m04.addrM [12]), .Z(n6855) );
  CNR3XL U6539 ( .A(\m04.addrM [10]), .B(n6805), .C(n6855), .Z(n6821) );
  CIVX2 U6540 ( .A(\m04.addrM [13]), .Z(n6490) );
  CND2X1 U6541 ( .A(n6490), .B(\m04.addrM [15]), .Z(n6538) );
  CNR3XL U6542 ( .A(\m04.addrM [16]), .B(\m04.addrM [14]), .C(n6538), .Z(n6852) );
  CIVX2 U6543 ( .A(\m04.addrM [0]), .Z(n6846) );
  CIVX2 U6544 ( .A(\m04.addrM [1]), .Z(n6847) );
  CNR2X1 U6545 ( .A(n6846), .B(n6847), .Z(n6322) );
  CIVXL U6546 ( .A(\m04.addrM [2]), .Z(n6453) );
  CND2X1 U6547 ( .A(\m04.addrM [3]), .B(\m04.addrM [4]), .Z(n6826) );
  CNR2X1 U6548 ( .A(n6453), .B(n6826), .Z(n6830) );
  CIVX2 U6549 ( .A(n6830), .Z(n6321) );
  CNR2X1 U6550 ( .A(n6453), .B(n6846), .Z(n6319) );
  CNR2X1 U6551 ( .A(\m04.addrM [3]), .B(\m04.addrM [4]), .Z(n6378) );
  CNR2X1 U6552 ( .A(\m04.addrM [2]), .B(\m04.addrM [1]), .Z(n6827) );
  CIVX2 U6553 ( .A(\m04.addrM [4]), .Z(n6483) );
  CND2X1 U6554 ( .A(\m04.addrM [3]), .B(n6483), .Z(n6482) );
  CNR2X1 U6555 ( .A(n6827), .B(n6482), .Z(n6411) );
  CNR2X1 U6556 ( .A(\m04.addrM [4]), .B(n6411), .Z(n6480) );
  CND2X1 U6557 ( .A(\m04.addrM [2]), .B(\m04.addrM [1]), .Z(n6485) );
  CND2X1 U6558 ( .A(n6378), .B(n6485), .Z(n6592) );
  CANR2X1 U6559 ( .A(n6319), .B(n6378), .C(n6480), .D(n6592), .Z(n6645) );
  CIVX2 U6560 ( .A(\m04.addrM [3]), .Z(n6484) );
  COND1XL U6561 ( .A(n6453), .B(n6484), .C(n6483), .Z(n6619) );
  CNR2X1 U6562 ( .A(\m04.addrM [2]), .B(n6826), .Z(n6320) );
  CANR3X1 U6563 ( .A(n6826), .B(n6619), .C(n6411), .D(n6320), .Z(n6824) );
  COND3X1 U6564 ( .A(n6322), .B(n6321), .C(n6645), .D(n6824), .Z(n6323) );
  CAN4X1 U6565 ( .A(n6324), .B(n6821), .C(n6852), .D(n6323), .Z(n7237) );
  CIVX2 U6566 ( .A(n7237), .Z(n6866) );
  COND2X1 U6567 ( .A(n7589), .B(n6325), .C(n7539), .D(n6866), .Z(n6334) );
  CIVX2 U6568 ( .A(n7549), .Z(n7581) );
  CIVX2 U6569 ( .A(\m01.addrM [12]), .Z(n6555) );
  CNR2X1 U6570 ( .A(\m01.addrM [11]), .B(n6555), .Z(n6909) );
  CIVX2 U6571 ( .A(\m01.addrM [9]), .Z(n6892) );
  CNR2X1 U6572 ( .A(\m01.addrM [10]), .B(n6892), .Z(n6326) );
  CND2X1 U6573 ( .A(n6909), .B(n6326), .Z(n6901) );
  CNR2X1 U6574 ( .A(\m01.addrM [14]), .B(\m01.addrM [13]), .Z(n6327) );
  CIVX2 U6575 ( .A(\m01.addrM [16]), .Z(n6375) );
  CND3XL U6576 ( .A(n6327), .B(\m01.addrM [15]), .C(n6375), .Z(n6910) );
  CIVX2 U6577 ( .A(\m01.addrM [4]), .Z(n6605) );
  CIVX2 U6578 ( .A(\m01.addrM [3]), .Z(n6607) );
  CNR2X1 U6579 ( .A(n6605), .B(n6607), .Z(n6885) );
  CND2X1 U6580 ( .A(\m01.addrM [2]), .B(n6885), .Z(n6914) );
  CNR2X1 U6581 ( .A(\m01.addrM [0]), .B(n6914), .Z(n6549) );
  CIVX2 U6582 ( .A(\m01.addrM [2]), .Z(n6456) );
  CIVX2 U6583 ( .A(\m01.addrM [1]), .Z(n6905) );
  CND2X1 U6584 ( .A(n6905), .B(n6456), .Z(n6884) );
  CANR1XL U6585 ( .A(\m01.addrM [2]), .B(\m01.addrM [3]), .C(\m01.addrM [4]), 
        .Z(n6933) );
  CANR1XL U6586 ( .A(n6885), .B(n6884), .C(n6933), .Z(n6918) );
  CND2X1 U6587 ( .A(\m01.addrM [3]), .B(n6605), .Z(n6470) );
  CNR2IX1 U6588 ( .B(n6884), .A(n6470), .Z(n6427) );
  CANR3X1 U6589 ( .A(n6885), .B(n6456), .C(n6918), .D(n6427), .Z(n6917) );
  CNR2X1 U6590 ( .A(\m01.addrM [4]), .B(\m01.addrM [3]), .Z(n6373) );
  CND2X1 U6591 ( .A(\m01.addrM [1]), .B(\m01.addrM [2]), .Z(n6606) );
  CND2X1 U6592 ( .A(n6373), .B(n6606), .Z(n6570) );
  CANR1XL U6593 ( .A(\m01.addrM [3]), .B(n6884), .C(\m01.addrM [4]), .Z(n6473)
         );
  COND4CX1 U6594 ( .A(\m01.addrM [2]), .B(\m01.addrM [0]), .C(n6570), .D(n6473), .Z(n6653) );
  COND3X1 U6595 ( .A(\m01.addrM [1]), .B(n6914), .C(n6917), .D(n6653), .Z(
        n6328) );
  CND2X1 U6596 ( .A(\m01.addrM [5]), .B(\m01.addrM [6]), .Z(n6657) );
  CND2X1 U6597 ( .A(\m01.addrM [7]), .B(\m01.addrM [8]), .Z(n6471) );
  CNR2X1 U6598 ( .A(n6657), .B(n6471), .Z(n6428) );
  COND1XL U6599 ( .A(n6549), .B(n6328), .C(n6428), .Z(n6329) );
  CNR3X1 U6600 ( .A(n6901), .B(n6910), .C(n6329), .Z(n7179) );
  CANR2XL U6601 ( .A(n7581), .B(n6789), .C(n7585), .D(n7179), .Z(n6331) );
  CND2X1 U6602 ( .A(n7583), .B(n7269), .Z(n6330) );
  COND3X1 U6603 ( .A(n6332), .B(n7577), .C(n6331), .D(n6330), .Z(n6333) );
  CANR3X1 U6604 ( .A(n7560), .B(n7497), .C(n6334), .D(n6333), .Z(n7525) );
  CMX2X1 U6605 ( .A0(n7687), .A1(\s05.Adr [1]), .S(n7525), .Z(n4723) );
  CANR2XL U6606 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [15]), .C(n7642), .D(
        \m01.DoutM [15]), .Z(n6338) );
  CANR2X1 U6607 ( .A(n7644), .B(\m03.DoutM [15]), .C(n7643), .D(
        \m02.DoutM [15]), .Z(n6337) );
  CANR2X1 U6608 ( .A(n7641), .B(\m05.DoutM [15]), .C(n7640), .D(
        \m06.DoutM [15]), .Z(n6336) );
  CND2X1 U6609 ( .A(n7648), .B(\m04.DoutM [15]), .Z(n6335) );
  CND4X1 U6610 ( .A(n6338), .B(n6337), .C(n6336), .D(n6335), .Z(n7635) );
  CMX2X1 U6611 ( .A0(n7635), .A1(\s05.dbus_in [15]), .S(n7525), .Z(n4721) );
  CANR2XL U6612 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [14]), .C(n7642), .D(
        \m01.DoutM [14]), .Z(n6342) );
  CANR2X1 U6613 ( .A(n7644), .B(\m03.DoutM [14]), .C(n7643), .D(
        \m02.DoutM [14]), .Z(n6341) );
  CANR2X1 U6614 ( .A(n7641), .B(\m05.DoutM [14]), .C(n7640), .D(
        \m06.DoutM [14]), .Z(n6340) );
  CND2X1 U6615 ( .A(n7648), .B(\m04.DoutM [14]), .Z(n6339) );
  CND4X1 U6616 ( .A(n6342), .B(n6341), .C(n6340), .D(n6339), .Z(n7636) );
  CMX2X1 U6617 ( .A0(n7636), .A1(\s05.dbus_in [14]), .S(n7525), .Z(n4720) );
  CANR2XL U6618 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [11]), .C(n7642), .D(
        \m01.DoutM [11]), .Z(n6346) );
  CANR2X1 U6619 ( .A(n7644), .B(\m03.DoutM [11]), .C(n7643), .D(
        \m02.DoutM [11]), .Z(n6345) );
  CANR2X1 U6620 ( .A(n7641), .B(\m05.DoutM [11]), .C(n7640), .D(
        \m06.DoutM [11]), .Z(n6344) );
  CND2X1 U6621 ( .A(n7648), .B(\m04.DoutM [11]), .Z(n6343) );
  CND4X1 U6622 ( .A(n6346), .B(n6345), .C(n6344), .D(n6343), .Z(n7628) );
  CMX2X1 U6623 ( .A0(n7628), .A1(\s05.dbus_in [11]), .S(n7525), .Z(n4717) );
  CANR2XL U6624 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [7]), .C(n7642), .D(
        \m01.DoutM [7]), .Z(n6350) );
  CANR2X1 U6625 ( .A(n7644), .B(\m03.DoutM [7]), .C(n7643), .D(\m02.DoutM [7]), 
        .Z(n6349) );
  CANR2X1 U6626 ( .A(n7641), .B(\m05.DoutM [7]), .C(n7640), .D(\m06.DoutM [7]), 
        .Z(n6348) );
  CND2X1 U6627 ( .A(n7648), .B(\m04.DoutM [7]), .Z(n6347) );
  CND4X1 U6628 ( .A(n6350), .B(n6349), .C(n6348), .D(n6347), .Z(n7629) );
  CMX2X1 U6629 ( .A0(n7629), .A1(\s05.dbus_in [7]), .S(n7525), .Z(n4713) );
  CANR2XL U6630 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [5]), .C(n7642), .D(
        \m01.DoutM [5]), .Z(n6354) );
  CANR2X1 U6631 ( .A(n7644), .B(\m03.DoutM [5]), .C(n7643), .D(\m02.DoutM [5]), 
        .Z(n6353) );
  CANR2X1 U6632 ( .A(n7641), .B(\m05.DoutM [5]), .C(n7640), .D(\m06.DoutM [5]), 
        .Z(n6352) );
  CND2X1 U6633 ( .A(n7648), .B(\m04.DoutM [5]), .Z(n6351) );
  CND4X1 U6634 ( .A(n6354), .B(n6353), .C(n6352), .D(n6351), .Z(n7630) );
  CMX2X1 U6635 ( .A0(n7630), .A1(\s05.dbus_in [5]), .S(n7525), .Z(n4711) );
  CANR2XL U6636 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [4]), .C(n7642), .D(
        \m01.DoutM [4]), .Z(n6358) );
  CANR2X1 U6637 ( .A(n7644), .B(\m03.DoutM [4]), .C(n7643), .D(\m02.DoutM [4]), 
        .Z(n6357) );
  CANR2X1 U6638 ( .A(n7641), .B(\m05.DoutM [4]), .C(n7640), .D(\m06.DoutM [4]), 
        .Z(n6356) );
  CND2X1 U6639 ( .A(n7648), .B(\m04.DoutM [4]), .Z(n6355) );
  CND4X1 U6640 ( .A(n6358), .B(n6357), .C(n6356), .D(n6355), .Z(n7653) );
  CMX2X1 U6641 ( .A0(n7653), .A1(\s05.dbus_in [4]), .S(n7525), .Z(n4710) );
  CANR2XL U6642 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [2]), .C(n7642), .D(
        \m01.DoutM [2]), .Z(n6362) );
  CANR2X1 U6643 ( .A(n7644), .B(\m03.DoutM [2]), .C(n7643), .D(\m02.DoutM [2]), 
        .Z(n6361) );
  CANR2X1 U6644 ( .A(n7641), .B(\m05.DoutM [2]), .C(n7640), .D(\m06.DoutM [2]), 
        .Z(n6360) );
  CND2X1 U6645 ( .A(n7648), .B(\m04.DoutM [2]), .Z(n6359) );
  CND4X1 U6646 ( .A(n6362), .B(n6361), .C(n6360), .D(n6359), .Z(n7683) );
  CMX2X1 U6647 ( .A0(n7683), .A1(\s05.dbus_in [2]), .S(n7525), .Z(n4708) );
  CANR2XL U6648 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [0]), .C(n7642), .D(
        \m01.DoutM [0]), .Z(n6366) );
  CANR2X1 U6649 ( .A(n7644), .B(\m03.DoutM [0]), .C(n7643), .D(\m02.DoutM [0]), 
        .Z(n6365) );
  CANR2X1 U6650 ( .A(n7641), .B(\m05.DoutM [0]), .C(n7640), .D(\m06.DoutM [0]), 
        .Z(n6364) );
  CND2X1 U6651 ( .A(n7648), .B(\m04.DoutM [0]), .Z(n6363) );
  CND4X1 U6652 ( .A(n6366), .B(n6365), .C(n6364), .D(n6363), .Z(n7684) );
  CMX2X1 U6653 ( .A0(n7684), .A1(\s05.dbus_in [0]), .S(n7525), .Z(n4706) );
  CANR2XL U6654 ( .A(\m00.YouGotIt ), .B(\m00.addrM [2]), .C(\m01.addrM [2]), 
        .D(n7642), .Z(n6368) );
  CANR2X1 U6655 ( .A(\m03.addrM [2]), .B(n7644), .C(\m02.addrM [2]), .D(n7643), 
        .Z(n6367) );
  COND3X1 U6656 ( .A(n7613), .B(n6369), .C(n6368), .D(n6367), .Z(n6370) );
  CANR1XL U6657 ( .A(\m05.addrM [2]), .B(n7641), .C(n6370), .Z(n6371) );
  COND1X1 U6658 ( .A(n6453), .B(n7616), .C(n6371), .Z(n7621) );
  CIVX2 U6659 ( .A(\m01.addrM [8]), .Z(n6372) );
  CIVX2 U6660 ( .A(n6657), .Z(n6894) );
  CND2X1 U6661 ( .A(n6372), .B(n6894), .Z(n6915) );
  CIVX2 U6662 ( .A(n6915), .Z(n6925) );
  CND2X1 U6663 ( .A(n6373), .B(n6456), .Z(n6374) );
  CIVX2 U6664 ( .A(\m01.addrM [7]), .Z(n6547) );
  CNR2X1 U6665 ( .A(\m01.addrM [8]), .B(n6547), .Z(n6923) );
  CANR1XL U6666 ( .A(n6925), .B(n6374), .C(n6923), .Z(n6377) );
  CND2X1 U6667 ( .A(\m01.addrM [6]), .B(n6923), .Z(n6548) );
  CIVX2 U6668 ( .A(\m01.addrM [5]), .Z(n6882) );
  CND2X1 U6669 ( .A(\m01.addrM [8]), .B(n6547), .Z(n6883) );
  CIVX2 U6670 ( .A(n6883), .Z(n6895) );
  CND2X1 U6671 ( .A(n6882), .B(n6895), .Z(n6455) );
  CNR2X1 U6672 ( .A(n6455), .B(\m01.addrM [6]), .Z(n6519) );
  CIVX2 U6673 ( .A(n6519), .Z(n6919) );
  CND2X1 U6674 ( .A(n6548), .B(n6919), .Z(n6889) );
  CNR2X1 U6675 ( .A(n6455), .B(\m01.addrM [0]), .Z(n6916) );
  CNR2X1 U6676 ( .A(\m01.addrM [1]), .B(n6374), .Z(n6896) );
  CND3XL U6677 ( .A(n6889), .B(n6916), .C(n6896), .Z(n6376) );
  CNR2X1 U6678 ( .A(\m01.addrM [15]), .B(n6375), .Z(n6477) );
  CIVX2 U6679 ( .A(\m01.addrM [13]), .Z(n6476) );
  CNR2X1 U6680 ( .A(\m01.addrM [14]), .B(n6476), .Z(n6886) );
  CND2X1 U6681 ( .A(n6477), .B(n6886), .Z(n6659) );
  CNR2X1 U6682 ( .A(\m01.addrM [10]), .B(\m01.addrM [9]), .Z(n6604) );
  CND2X1 U6683 ( .A(n6909), .B(n6604), .Z(n6576) );
  CANR3X1 U6684 ( .A(n6377), .B(n6376), .C(n6659), .D(n6576), .Z(n7185) );
  CNR2X1 U6685 ( .A(\m04.addrM [9]), .B(\m04.addrM [10]), .Z(n6515) );
  CND2IX1 U6686 ( .B(n6855), .A(n6515), .Z(n6597) );
  CND2X1 U6687 ( .A(n6378), .B(n6827), .Z(n6817) );
  CIVX2 U6688 ( .A(n6817), .Z(n6809) );
  CNR2X1 U6689 ( .A(\m04.addrM [7]), .B(n7617), .Z(n6806) );
  CIVX2 U6690 ( .A(n6806), .Z(n6815) );
  CNR2X1 U6691 ( .A(\m04.addrM [6]), .B(n6815), .Z(n6851) );
  CND2X1 U6692 ( .A(n6851), .B(n6845), .Z(n6518) );
  CNR2X1 U6693 ( .A(\m04.addrM [0]), .B(n6518), .Z(n6381) );
  CNR2X1 U6694 ( .A(\m04.addrM [2]), .B(\m04.addrM [4]), .Z(n6379) );
  CND2X1 U6695 ( .A(\m04.addrM [5]), .B(\m04.addrM [6]), .Z(n6814) );
  CNR2X1 U6696 ( .A(\m04.addrM [7]), .B(\m04.addrM [8]), .Z(n6594) );
  CND2IX1 U6697 ( .B(n6814), .A(n6594), .Z(n6513) );
  CND2X1 U6698 ( .A(\m04.addrM [7]), .B(n7617), .Z(n6825) );
  COND4CX1 U6699 ( .A(n6379), .B(n6484), .C(n6513), .D(n6825), .Z(n6380) );
  CND2IX1 U6700 ( .B(\m04.addrM [14]), .A(\m04.addrM [16]), .Z(n6536) );
  CNR3XL U6701 ( .A(\m04.addrM [15]), .B(n6536), .C(n6490), .Z(n6650) );
  COND4CX1 U6702 ( .A(n6809), .B(n6381), .C(n6380), .D(n6650), .Z(n6382) );
  CNR2X1 U6703 ( .A(n6597), .B(n6382), .Z(n7242) );
  CIVX2 U6704 ( .A(n7242), .Z(n6383) );
  COND2X1 U6705 ( .A(n7589), .B(n6384), .C(n7539), .D(n6383), .Z(n6394) );
  CANR2XL U6706 ( .A(n7581), .B(n6791), .C(n7583), .D(n7266), .Z(n6391) );
  CIVX2 U6707 ( .A(\m03.addrM [7]), .Z(n7543) );
  CND2X1 U6708 ( .A(\m03.addrM [8]), .B(n7543), .Z(n7317) );
  COR2X1 U6709 ( .A(n7317), .B(\m03.addrM [6]), .Z(n6496) );
  CNR2X1 U6710 ( .A(\m03.addrM [5]), .B(n6496), .Z(n7284) );
  CNR2X1 U6711 ( .A(\m03.addrM [1]), .B(\m03.addrM [0]), .Z(n6529) );
  CND2X1 U6712 ( .A(n6385), .B(n6635), .Z(n6580) );
  CNR2X1 U6713 ( .A(\m03.addrM [4]), .B(n6580), .Z(n7304) );
  CIVX2 U6714 ( .A(n7304), .Z(n6387) );
  CNR2X1 U6715 ( .A(\m03.addrM [7]), .B(\m03.addrM [8]), .Z(n6587) );
  CIVXL U6716 ( .A(\m03.addrM [5]), .Z(n6633) );
  CNR2X1 U6717 ( .A(n7567), .B(n6633), .Z(n7319) );
  CND2X1 U6718 ( .A(n6587), .B(n7319), .Z(n7300) );
  CND2X1 U6719 ( .A(n6387), .B(n7300), .Z(n6386) );
  COND4CX1 U6720 ( .A(n7284), .B(n6529), .C(n6387), .D(n6386), .Z(n6389) );
  CNR2X1 U6721 ( .A(\m03.addrM [8]), .B(n7543), .Z(n6495) );
  CIVX2 U6722 ( .A(n6495), .Z(n6508) );
  CNR2X1 U6723 ( .A(\m03.addrM [15]), .B(n6388), .Z(n6500) );
  CIVX2 U6724 ( .A(\m03.addrM [13]), .Z(n6499) );
  CNR2X1 U6725 ( .A(\m03.addrM [14]), .B(n6499), .Z(n7323) );
  CND2X1 U6726 ( .A(n6500), .B(n7323), .Z(n6640) );
  CNR2X1 U6727 ( .A(\m03.addrM [9]), .B(\m03.addrM [10]), .Z(n6615) );
  CND2X1 U6728 ( .A(n6615), .B(n7310), .Z(n6588) );
  CANR3X1 U6729 ( .A(n6389), .B(n6508), .C(n6640), .D(n6588), .Z(n7496) );
  CND2X1 U6730 ( .A(n7560), .B(n7496), .Z(n6390) );
  COND3X1 U6731 ( .A(n6392), .B(n7577), .C(n6391), .D(n6390), .Z(n6393) );
  CANR3X1 U6732 ( .A(n7585), .B(n7185), .C(n6394), .D(n6393), .Z(n7573) );
  CMX2X1 U6733 ( .A0(n7621), .A1(\s08.Adr [2]), .S(n7573), .Z(n4532) );
  CANR2XL U6734 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [13]), .C(n7642), .D(
        \m01.DoutM [13]), .Z(n6398) );
  CANR2X1 U6735 ( .A(n7644), .B(\m03.DoutM [13]), .C(n7643), .D(
        \m02.DoutM [13]), .Z(n6397) );
  CANR2X1 U6736 ( .A(n7641), .B(\m05.DoutM [13]), .C(n7640), .D(
        \m06.DoutM [13]), .Z(n6396) );
  CND2X1 U6737 ( .A(n7648), .B(\m04.DoutM [13]), .Z(n6395) );
  CND4X1 U6738 ( .A(n6398), .B(n6397), .C(n6396), .D(n6395), .Z(n7627) );
  CMX2X1 U6739 ( .A0(n7627), .A1(\s08.dbus_in [13]), .S(n7573), .Z(n4527) );
  CMX2X1 U6740 ( .A0(n7628), .A1(\s08.dbus_in [11]), .S(n7573), .Z(n4525) );
  CANR2XL U6741 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [10]), .C(n7642), .D(
        \m01.DoutM [10]), .Z(n6402) );
  CANR2X1 U6742 ( .A(n7644), .B(\m03.DoutM [10]), .C(n7643), .D(
        \m02.DoutM [10]), .Z(n6401) );
  CANR2X1 U6743 ( .A(n7641), .B(\m05.DoutM [10]), .C(n7640), .D(
        \m06.DoutM [10]), .Z(n6400) );
  CND2X1 U6744 ( .A(n7648), .B(\m04.DoutM [10]), .Z(n6399) );
  CND4X1 U6745 ( .A(n6402), .B(n6401), .C(n6400), .D(n6399), .Z(n7626) );
  CMX2X1 U6746 ( .A0(n7626), .A1(\s08.dbus_in [10]), .S(n7573), .Z(n4524) );
  CMX2X1 U6747 ( .A0(n7629), .A1(\s08.dbus_in [7]), .S(n7573), .Z(n4521) );
  CMX2X1 U6748 ( .A0(n7630), .A1(\s08.dbus_in [5]), .S(n7573), .Z(n4519) );
  CANR2XL U6749 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [3]), .C(n7642), .D(
        \m01.DoutM [3]), .Z(n6406) );
  CANR2X1 U6750 ( .A(n7644), .B(\m03.DoutM [3]), .C(n7643), .D(\m02.DoutM [3]), 
        .Z(n6405) );
  CANR2X1 U6751 ( .A(n7641), .B(\m05.DoutM [3]), .C(n7640), .D(\m06.DoutM [3]), 
        .Z(n6404) );
  CND2X1 U6752 ( .A(n7648), .B(\m04.DoutM [3]), .Z(n6403) );
  CND4X1 U6753 ( .A(n6406), .B(n6405), .C(n6404), .D(n6403), .Z(n7631) );
  CMX2X1 U6754 ( .A0(n7631), .A1(\s08.dbus_in [3]), .S(n7573), .Z(n4517) );
  CANR2XL U6755 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [1]), .C(n7642), .D(
        \m01.DoutM [1]), .Z(n6410) );
  CANR2X1 U6756 ( .A(n7644), .B(\m03.DoutM [1]), .C(n7643), .D(\m02.DoutM [1]), 
        .Z(n6409) );
  CANR2X1 U6757 ( .A(n7641), .B(\m05.DoutM [1]), .C(n7640), .D(\m06.DoutM [1]), 
        .Z(n6408) );
  CND2X1 U6758 ( .A(n7648), .B(\m04.DoutM [1]), .Z(n6407) );
  CND4X1 U6759 ( .A(n6410), .B(n6409), .C(n6408), .D(n6407), .Z(n7632) );
  CMX2X1 U6760 ( .A0(n7632), .A1(\s08.dbus_in [1]), .S(n7573), .Z(n4515) );
  CND2X1 U6761 ( .A(\m04.addrM [16]), .B(\m04.addrM [14]), .Z(n6842) );
  CNR2X1 U6762 ( .A(\m04.addrM [15]), .B(n6842), .Z(n6491) );
  CND2X1 U6763 ( .A(\m04.addrM [13]), .B(n6491), .Z(n6596) );
  CND2X1 U6764 ( .A(n6411), .B(n6485), .Z(n6643) );
  CNR2X1 U6765 ( .A(\m04.addrM [5]), .B(\m04.addrM [6]), .Z(n6591) );
  CNR2X1 U6766 ( .A(n6591), .B(n6815), .Z(n6412) );
  CANR4CX1 U6767 ( .A(n6480), .B(n6814), .C(n6488), .D(n6412), .Z(n6413) );
  COND1XL U6768 ( .A(n6543), .B(n6643), .C(n6413), .Z(n6415) );
  CANR3X1 U6769 ( .A(n6827), .B(n6484), .C(n6483), .D(n6518), .Z(n6414) );
  CND2X1 U6770 ( .A(\m04.addrM [10]), .B(n6805), .Z(n6854) );
  CND2X1 U6771 ( .A(\m04.addrM [11]), .B(\m04.addrM [12]), .Z(n6621) );
  CNR2X1 U6772 ( .A(n6854), .B(n6621), .Z(n6839) );
  COND1XL U6773 ( .A(n6415), .B(n6414), .C(n6839), .Z(n6416) );
  CNR2X1 U6774 ( .A(n6596), .B(n6416), .Z(n7239) );
  CIVX2 U6775 ( .A(n7239), .Z(n6417) );
  COND2X1 U6776 ( .A(n7577), .B(n6418), .C(n7539), .D(n6417), .Z(n6439) );
  CNR2X1 U6777 ( .A(\m03.addrM [6]), .B(\m03.addrM [5]), .Z(n6583) );
  CNR2X1 U6778 ( .A(n7319), .B(n6583), .Z(n7285) );
  CNR2IX1 U6779 ( .B(n7319), .A(n7317), .Z(n7307) );
  CNR2IX1 U6780 ( .B(n6583), .A(n6419), .Z(n6494) );
  CANR3X1 U6781 ( .A(\m03.addrM [8]), .B(n7285), .C(n7307), .D(n6494), .Z(
        n6426) );
  CNR2X1 U6782 ( .A(n6614), .B(\m03.addrM [4]), .Z(n6423) );
  CIVX2 U6783 ( .A(n6636), .Z(n7295) );
  CNR2X1 U6784 ( .A(\m03.addrM [3]), .B(n7295), .Z(n6421) );
  CND2X1 U6785 ( .A(\m03.addrM [4]), .B(n7284), .Z(n6420) );
  COND2X1 U6786 ( .A(n6421), .B(n6420), .C(n7301), .D(n6419), .Z(n6422) );
  CANR1XL U6787 ( .A(n6423), .B(n6530), .C(n6422), .Z(n6425) );
  CND3XL U6788 ( .A(\m03.addrM [13]), .B(\m03.addrM [14]), .C(n6500), .Z(n6589) );
  CNR2X1 U6789 ( .A(\m03.addrM [9]), .B(n6424), .Z(n7294) );
  CND3XL U6790 ( .A(\m03.addrM [12]), .B(\m03.addrM [11]), .C(n7294), .Z(n7302) );
  CANR3X2 U6791 ( .A(n6426), .B(n6425), .C(n6589), .D(n7302), .Z(n7504) );
  CANR2X1 U6792 ( .A(n7560), .B(n7504), .C(n7581), .D(n6784), .Z(n6436) );
  CND2X1 U6793 ( .A(n6427), .B(n6606), .Z(n6652) );
  CIVX2 U6794 ( .A(n6428), .Z(n6432) );
  COND1XL U6795 ( .A(\m01.addrM [3]), .B(n6884), .C(\m01.addrM [4]), .Z(n6429)
         );
  COND2X1 U6796 ( .A(n6894), .B(n6471), .C(n6919), .D(n6429), .Z(n6430) );
  CANR4CX1 U6797 ( .A(\m01.addrM [5]), .B(\m01.addrM [6]), .C(n6895), .D(n6430), .Z(n6431) );
  COND1XL U6798 ( .A(n6652), .B(n6432), .C(n6431), .Z(n6433) );
  CANR11X1 U6799 ( .A(\m01.addrM [5]), .B(\m01.addrM [8]), .C(n6473), .D(n6433), .Z(n6434) );
  CND3XL U6800 ( .A(\m01.addrM [14]), .B(\m01.addrM [13]), .C(n6477), .Z(n6577) );
  CND2X1 U6801 ( .A(\m01.addrM [10]), .B(n6892), .Z(n6911) );
  CIVX2 U6802 ( .A(n6911), .Z(n6551) );
  CND3XL U6803 ( .A(n6551), .B(\m01.addrM [11]), .C(\m01.addrM [12]), .Z(n6936) );
  CNR3X1 U6804 ( .A(n6434), .B(n6577), .C(n6936), .Z(n7184) );
  CND2X1 U6805 ( .A(n7585), .B(n7184), .Z(n6435) );
  COND3X1 U6806 ( .A(n6437), .B(n7589), .C(n6436), .D(n6435), .Z(n6438) );
  CANR3X1 U6807 ( .A(n7583), .B(n7271), .C(n6439), .D(n6438), .Z(n7592) );
  CMX2X1 U6808 ( .A0(n7621), .A1(\s09.Adr [2]), .S(n7592), .Z(n4468) );
  CANR2XL U6809 ( .A(\m00.YouGotIt ), .B(\m00.addrM [0]), .C(\m01.addrM [0]), 
        .D(n7642), .Z(n6443) );
  CANR2X1 U6810 ( .A(\m03.addrM [0]), .B(n7644), .C(\m02.addrM [0]), .D(n7643), 
        .Z(n6442) );
  CANR2X1 U6811 ( .A(\m05.addrM [0]), .B(n7641), .C(n7640), .D(\m06.addrM [0]), 
        .Z(n6441) );
  CND2X1 U6812 ( .A(\m04.addrM [0]), .B(n7648), .Z(n6440) );
  CND4X1 U6813 ( .A(n6443), .B(n6442), .C(n6441), .D(n6440), .Z(n7625) );
  CMX2X1 U6814 ( .A0(n7625), .A1(\s09.Adr [0]), .S(n7592), .Z(n4466) );
  CMX2X1 U6815 ( .A0(n7635), .A1(\s09.dbus_in [15]), .S(n7592), .Z(n4465) );
  CANR2XL U6816 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [12]), .C(n7642), .D(
        \m01.DoutM [12]), .Z(n6447) );
  CANR2X1 U6817 ( .A(n7644), .B(\m03.DoutM [12]), .C(n7643), .D(
        \m02.DoutM [12]), .Z(n6446) );
  CANR2X1 U6818 ( .A(n7641), .B(\m05.DoutM [12]), .C(n7640), .D(
        \m06.DoutM [12]), .Z(n6445) );
  CND2X1 U6819 ( .A(n7648), .B(\m04.DoutM [12]), .Z(n6444) );
  CND4X1 U6820 ( .A(n6447), .B(n6446), .C(n6445), .D(n6444), .Z(n7637) );
  CMX2X1 U6821 ( .A0(n7637), .A1(\s09.dbus_in [12]), .S(n7592), .Z(n4462) );
  CMX2X1 U6822 ( .A0(n7626), .A1(\s09.dbus_in [10]), .S(n7592), .Z(n4460) );
  CMX2X1 U6823 ( .A0(n7629), .A1(\s09.dbus_in [7]), .S(n7592), .Z(n4457) );
  CMX2X1 U6824 ( .A0(n7630), .A1(\s09.dbus_in [5]), .S(n7592), .Z(n4455) );
  CMX2X1 U6825 ( .A0(n7631), .A1(\s09.dbus_in [3]), .S(n7592), .Z(n4453) );
  CMX2X1 U6826 ( .A0(n7632), .A1(\s09.dbus_in [1]), .S(n7592), .Z(n4451) );
  CNR2X1 U6827 ( .A(\m03.addrM [5]), .B(n7317), .Z(n6497) );
  CND2X1 U6828 ( .A(\m03.addrM [6]), .B(n6497), .Z(n7299) );
  CIVX2 U6829 ( .A(n7299), .Z(n7305) );
  CANR1XL U6830 ( .A(n6635), .B(n6448), .C(n6634), .Z(n6581) );
  CANR1XL U6831 ( .A(\m03.addrM [4]), .B(n6614), .C(n6581), .Z(n7306) );
  CNR2X1 U6832 ( .A(n6449), .B(n6580), .Z(n6450) );
  CANR4CX1 U6833 ( .A(n6450), .B(n6634), .C(n6633), .D(n6496), .Z(n6451) );
  COND4CX1 U6834 ( .A(n7305), .B(n7306), .C(n6451), .D(n7294), .Z(n6452) );
  CNR4X2 U6835 ( .A(\m03.addrM [12]), .B(\m03.addrM [11]), .C(n6589), .D(n6452), .Z(n7493) );
  CND2X1 U6836 ( .A(\m04.addrM [1]), .B(n6453), .Z(n6828) );
  COND1XL U6837 ( .A(\m04.addrM [2]), .B(\m04.addrM [3]), .C(\m04.addrM [4]), 
        .Z(n6848) );
  CND2X1 U6838 ( .A(n6806), .B(n6814), .Z(n6833) );
  CNR2IX1 U6839 ( .B(\m04.addrM [6]), .A(n6833), .Z(n6849) );
  COND1XL U6840 ( .A(\m04.addrM [0]), .B(\m04.addrM [1]), .C(\m04.addrM [2]), 
        .Z(n6539) );
  CANR1XL U6841 ( .A(n6539), .B(n6484), .C(n6483), .Z(n6816) );
  CNR3XL U6842 ( .A(\m04.addrM [11]), .B(\m04.addrM [12]), .C(n6596), .Z(n6514) );
  CIVXL U6843 ( .A(n7243), .Z(n6874) );
  COND2X1 U6844 ( .A(n7577), .B(n7674), .C(n7539), .D(n6874), .Z(n6465) );
  CIVX2 U6845 ( .A(n6732), .Z(n6463) );
  CANR2XL U6846 ( .A(n7581), .B(n6790), .C(n7583), .D(n7268), .Z(n6462) );
  CND2IX1 U6847 ( .B(n6606), .A(\m01.addrM [4]), .Z(n6468) );
  CND2X1 U6848 ( .A(\m01.addrM [0]), .B(\m01.addrM [2]), .Z(n6454) );
  CAOR1X1 U6849 ( .A(n6607), .B(n6454), .C(n6605), .Z(n6571) );
  CND2X1 U6850 ( .A(n6468), .B(n6571), .Z(n6899) );
  CND2IX1 U6851 ( .B(n6455), .A(\m01.addrM [6]), .Z(n6897) );
  CND2X1 U6852 ( .A(\m01.addrM [0]), .B(n6519), .Z(n6904) );
  CND2X1 U6853 ( .A(\m01.addrM [1]), .B(n6456), .Z(n6927) );
  COND1XL U6854 ( .A(\m01.addrM [2]), .B(\m01.addrM [3]), .C(\m01.addrM [4]), 
        .Z(n6907) );
  CIVX2 U6855 ( .A(\m01.addrM [6]), .Z(n7562) );
  CND2X1 U6856 ( .A(n6895), .B(n7562), .Z(n6929) );
  CAOR1X1 U6857 ( .A(n6882), .B(n6907), .C(n6929), .Z(n6457) );
  COND11X1 U6858 ( .A(n6605), .B(n6904), .C(n6927), .D(n6457), .Z(n6458) );
  CIVX2 U6859 ( .A(n6458), .Z(n6460) );
  COR4X1 U6860 ( .A(\m01.addrM [12]), .B(\m01.addrM [11]), .C(n6911), .D(n6577), .Z(n6459) );
  CANR4CX1 U6861 ( .A(n6899), .B(n6897), .C(n6460), .D(n6459), .Z(n7180) );
  CND2XL U6862 ( .A(n7585), .B(n7180), .Z(n6461) );
  COND3X1 U6863 ( .A(n6463), .B(n7589), .C(n6462), .D(n6461), .Z(n6464) );
  CANR3X1 U6864 ( .A(n7560), .B(n7493), .C(n6465), .D(n6464), .Z(n7593) );
  CMX2X1 U6865 ( .A0(n7621), .A1(\s10.Adr [2]), .S(n7593), .Z(n4404) );
  CMX2X1 U6866 ( .A0(n7687), .A1(\s10.Adr [1]), .S(n7593), .Z(n4403) );
  CMX2X1 U6867 ( .A0(n7636), .A1(\s10.dbus_in [14]), .S(n7593), .Z(n4400) );
  CMX2X1 U6868 ( .A0(n7637), .A1(\s10.dbus_in [12]), .S(n7593), .Z(n4398) );
  CMX2X1 U6869 ( .A0(n7628), .A1(\s10.dbus_in [11]), .S(n7593), .Z(n4397) );
  CMX2X1 U6870 ( .A0(n7629), .A1(\s10.dbus_in [7]), .S(n7593), .Z(n4393) );
  CMX2X1 U6871 ( .A0(n7630), .A1(\s10.dbus_in [5]), .S(n7593), .Z(n4391) );
  CMX2X1 U6872 ( .A0(n7631), .A1(\s10.dbus_in [3]), .S(n7593), .Z(n4389) );
  CMX2X1 U6873 ( .A0(n7632), .A1(\s10.dbus_in [1]), .S(n7593), .Z(n4387) );
  CND2X1 U6874 ( .A(n6923), .B(n7562), .Z(n6466) );
  CNR2X1 U6875 ( .A(n6882), .B(n6466), .Z(n6654) );
  CNR2X1 U6876 ( .A(n6466), .B(\m01.addrM [5]), .Z(n6574) );
  CIVX2 U6877 ( .A(n6574), .Z(n6467) );
  COND3X1 U6878 ( .A(n6468), .B(n6467), .C(n6548), .D(n6883), .Z(n6469) );
  CANR3X1 U6879 ( .A(n6923), .B(n6885), .C(n6654), .D(n6469), .Z(n6479) );
  CNR3XL U6880 ( .A(\m01.addrM [0]), .B(n6470), .C(n6927), .Z(n6474) );
  CIVX2 U6881 ( .A(n6471), .Z(n6472) );
  CNR2X1 U6882 ( .A(\m01.addrM [5]), .B(\m01.addrM [6]), .Z(n6658) );
  COND3X1 U6883 ( .A(n6474), .B(n6473), .C(n6472), .D(n6658), .Z(n6478) );
  CNR2X1 U6884 ( .A(\m01.addrM [11]), .B(\m01.addrM [12]), .Z(n6475) );
  CND2X1 U6885 ( .A(n6604), .B(n6475), .Z(n6520) );
  CND3XL U6886 ( .A(\m01.addrM [14]), .B(n6477), .C(n6476), .Z(n6902) );
  CANR3X1 U6887 ( .A(n6479), .B(n6478), .C(n6520), .D(n6902), .Z(n7187) );
  CIVX2 U6888 ( .A(n6480), .Z(n6481) );
  COND11X1 U6889 ( .A(\m04.addrM [0]), .B(n6482), .C(n6828), .D(n6481), .Z(
        n6487) );
  CANR3X1 U6890 ( .A(n6485), .B(n6484), .C(n6483), .D(n6825), .Z(n6486) );
  CANR11X1 U6891 ( .A(n6591), .B(n6488), .C(n6487), .D(n6486), .Z(n6489) );
  CND2X1 U6892 ( .A(\m04.addrM [6]), .B(n6836), .Z(n6808) );
  CND2X1 U6893 ( .A(\m04.addrM [5]), .B(n6836), .Z(n6642) );
  CAN4X1 U6894 ( .A(n6489), .B(n6808), .C(n6642), .D(n6815), .Z(n6492) );
  CAN2X1 U6895 ( .A(n6491), .B(n6490), .Z(n6820) );
  CND2X1 U6896 ( .A(n6515), .B(n6820), .Z(n6620) );
  CNR4X2 U6897 ( .A(\m04.addrM [11]), .B(\m04.addrM [12]), .C(n6492), .D(n6620), .Z(n7238) );
  CIVX2 U6898 ( .A(n7238), .Z(n6865) );
  COND2X1 U6899 ( .A(n7577), .B(n6493), .C(n7539), .D(n6865), .Z(n6505) );
  CND2X1 U6900 ( .A(n6495), .B(n7567), .Z(n7298) );
  CNR2X1 U6901 ( .A(n6635), .B(n6634), .Z(n7296) );
  CND2X1 U6902 ( .A(\m03.addrM [6]), .B(n6495), .Z(n6528) );
  CND2X1 U6903 ( .A(n6528), .B(n6496), .Z(n7313) );
  CNR2X1 U6904 ( .A(n6497), .B(n7313), .Z(n7297) );
  CNR2X1 U6905 ( .A(\m03.addrM [12]), .B(\m03.addrM [11]), .Z(n6498) );
  CND2X1 U6906 ( .A(n6615), .B(n6498), .Z(n6510) );
  CND3XL U6907 ( .A(\m03.addrM [14]), .B(n6500), .C(n6499), .Z(n6617) );
  CIVX2 U6908 ( .A(n6617), .Z(n7309) );
  CIVX2 U6909 ( .A(n7436), .Z(n7494) );
  CANR2XL U6910 ( .A(n7560), .B(n7494), .C(n7583), .D(n7273), .Z(n6502) );
  CND2X1 U6911 ( .A(n7581), .B(n6786), .Z(n6501) );
  COND3X1 U6912 ( .A(n6503), .B(n7589), .C(n6502), .D(n6501), .Z(n6504) );
  CANR3X1 U6913 ( .A(n7585), .B(n7187), .C(n6505), .D(n6504), .Z(n7594) );
  CMX2X1 U6914 ( .A0(n7621), .A1(\s11.Adr [2]), .S(n7594), .Z(n4340) );
  CMX2X1 U6915 ( .A0(n7625), .A1(\s11.Adr [0]), .S(n7594), .Z(n4338) );
  CMX2X1 U6916 ( .A0(n7627), .A1(\s11.dbus_in [13]), .S(n7594), .Z(n4335) );
  COND2X1 U6917 ( .A(n7589), .B(n6507), .C(n7549), .D(n6506), .Z(n6526) );
  COAN1X1 U6918 ( .A(n7300), .B(n6585), .C(n6508), .Z(n6512) );
  CANR1XL U6919 ( .A(\m03.addrM [2]), .B(\m03.addrM [3]), .C(\m03.addrM [4]), 
        .Z(n6509) );
  CND2X1 U6920 ( .A(n7284), .B(n6509), .Z(n6511) );
  CANR3X1 U6921 ( .A(n6512), .B(n6511), .C(n6510), .D(n6589), .Z(n7499) );
  CIVX2 U6922 ( .A(n7539), .Z(n7579) );
  CIVX2 U6923 ( .A(n6513), .Z(n6838) );
  CANR1XL U6924 ( .A(n6838), .B(n6592), .C(n6836), .Z(n6517) );
  CND2X1 U6925 ( .A(n6515), .B(n6514), .Z(n6516) );
  CANR4CX1 U6926 ( .A(n6619), .B(n6518), .C(n6517), .D(n6516), .Z(n7236) );
  CANR2XL U6927 ( .A(n7560), .B(n7499), .C(n7579), .D(n7236), .Z(n6524) );
  CANR2X1 U6928 ( .A(n6519), .B(n6933), .C(n6925), .D(n6570), .Z(n6522) );
  CIVX2 U6929 ( .A(n6923), .Z(n6521) );
  CANR3X1 U6930 ( .A(n6522), .B(n6521), .C(n6520), .D(n6577), .Z(n7183) );
  CND2X1 U6931 ( .A(n7585), .B(n7183), .Z(n6523) );
  COND3X1 U6932 ( .A(n6686), .B(n7577), .C(n6524), .D(n6523), .Z(n6525) );
  CANR3X1 U6933 ( .A(n7583), .B(n7270), .C(n6526), .D(n6525), .Z(n7595) );
  CMX2X1 U6934 ( .A0(n7621), .A1(\s13.Adr [2]), .S(n7595), .Z(n5124) );
  CMX2X1 U6935 ( .A0(n7625), .A1(\s13.Adr [0]), .S(n7595), .Z(n5122) );
  CMX2X1 U6936 ( .A0(n7627), .A1(\s13.dbus_in [13]), .S(n7595), .Z(n5119) );
  CMX2X1 U6937 ( .A0(n7628), .A1(\s13.dbus_in [11]), .S(n7595), .Z(n5117) );
  CMX2X1 U6938 ( .A0(n7626), .A1(\s13.dbus_in [10]), .S(n7595), .Z(n5116) );
  CMX2X1 U6939 ( .A0(n7629), .A1(\s13.dbus_in [7]), .S(n7595), .Z(n5113) );
  CMX2X1 U6940 ( .A0(n7630), .A1(\s13.dbus_in [5]), .S(n7595), .Z(n5111) );
  CMX2X1 U6941 ( .A0(n7631), .A1(\s13.dbus_in [3]), .S(n7595), .Z(n5109) );
  CMX2X1 U6942 ( .A0(n7632), .A1(\s13.dbus_in [1]), .S(n7595), .Z(n5107) );
  CAN4X1 U6943 ( .A(\m03.addrM [11]), .B(\m03.addrM [15]), .C(\m03.addrM [16]), 
        .D(n6527), .Z(n7322) );
  CND2X1 U6944 ( .A(\m03.addrM [2]), .B(n7296), .Z(n7290) );
  CNR2X1 U6945 ( .A(\m03.addrM [5]), .B(n6528), .Z(n7315) );
  CANR4CX1 U6946 ( .A(n6529), .B(n7290), .C(n7315), .D(n6587), .Z(n6533) );
  CIVX2 U6947 ( .A(n7290), .Z(n6531) );
  CANR4CX1 U6948 ( .A(\m03.addrM [5]), .B(n6531), .C(n6530), .D(\m03.addrM [9]), .Z(n6532) );
  CANR11X1 U6949 ( .A(\m03.addrM [9]), .B(n6533), .C(n7298), .D(n6532), .Z(
        n6534) );
  CND4X1 U6950 ( .A(n7322), .B(\m03.addrM [10]), .C(n6535), .D(n6534), .Z(
        n7471) );
  COND2X1 U6951 ( .A(n7577), .B(n6677), .C(n7471), .D(n7575), .Z(n6561) );
  CNR3XL U6952 ( .A(\m04.addrM [12]), .B(n6537), .C(n6536), .Z(n6812) );
  CIVX2 U6953 ( .A(n6538), .Z(n6545) );
  CNR2X1 U6954 ( .A(\m04.addrM [5]), .B(n6830), .Z(n6844) );
  CNR2X1 U6955 ( .A(n6539), .B(n6826), .Z(n6540) );
  CANR4CX1 U6956 ( .A(n6540), .B(\m04.addrM [5]), .C(\m04.addrM [6]), .D(n6825), .Z(n6541) );
  COND3X1 U6957 ( .A(n6594), .B(n6541), .C(\m04.addrM [9]), .D(\m04.addrM [10]), .Z(n6542) );
  COND11X1 U6958 ( .A(n6844), .B(n6854), .C(n6543), .D(n6542), .Z(n6544) );
  CND3XL U6959 ( .A(n6812), .B(n6545), .C(n6544), .Z(n6804) );
  COND2X1 U6960 ( .A(n7549), .B(n6546), .C(n6804), .D(n7539), .Z(n6560) );
  CANR3X1 U6961 ( .A(n6914), .B(n6882), .C(n7562), .D(n6547), .Z(n6552) );
  CNR2X1 U6962 ( .A(\m01.addrM [5]), .B(n6548), .Z(n6608) );
  CND2X1 U6963 ( .A(n6549), .B(n6608), .Z(n6550) );
  COND2X1 U6964 ( .A(\m01.addrM [8]), .B(n6552), .C(\m01.addrM [1]), .D(n6550), 
        .Z(n6554) );
  CAN3X2 U6965 ( .A(\m01.addrM [8]), .B(n6552), .C(n6551), .Z(n6553) );
  CANR11X1 U6966 ( .A(\m01.addrM [9]), .B(\m01.addrM [10]), .C(n6554), .D(
        n6553), .Z(n6556) );
  CND4X1 U6967 ( .A(\m01.addrM [11]), .B(\m01.addrM [16]), .C(\m01.addrM [15]), 
        .D(n6555), .Z(n6891) );
  CNR4X2 U6968 ( .A(\m01.addrM [14]), .B(\m01.addrM [13]), .C(n6556), .D(n6891), .Z(n7181) );
  CANR2XL U6969 ( .A(n7181), .B(n7585), .C(n7265), .D(n7583), .Z(n6557) );
  COND1XL U6970 ( .A(n6558), .B(n7589), .C(n6557), .Z(n6559) );
  CNR3XL U6971 ( .A(n6561), .B(n6560), .C(n6559), .Z(n7596) );
  CMX2X1 U6972 ( .A0(n7621), .A1(\s00.Adr [2]), .S(n7596), .Z(n5060) );
  CANR2XL U6973 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [8]), .C(n7642), .D(
        \m01.DoutM [8]), .Z(n6565) );
  CANR2X1 U6974 ( .A(n7644), .B(\m03.DoutM [8]), .C(n7643), .D(\m02.DoutM [8]), 
        .Z(n6564) );
  CANR2X1 U6975 ( .A(n7641), .B(\m05.DoutM [8]), .C(n7640), .D(\m06.DoutM [8]), 
        .Z(n6563) );
  CND2X1 U6976 ( .A(n7648), .B(\m04.DoutM [8]), .Z(n6562) );
  CND4X1 U6977 ( .A(n6565), .B(n6564), .C(n6563), .D(n6562), .Z(n7685) );
  CMX2X1 U6978 ( .A0(n7685), .A1(\s00.dbus_in [8]), .S(n7596), .Z(n5050) );
  CANR2XL U6979 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [6]), .C(n7642), .D(
        \m01.DoutM [6]), .Z(n6569) );
  CANR2X1 U6980 ( .A(n7644), .B(\m03.DoutM [6]), .C(n7643), .D(\m02.DoutM [6]), 
        .Z(n6568) );
  CANR2X1 U6981 ( .A(n7641), .B(\m05.DoutM [6]), .C(n7640), .D(\m06.DoutM [6]), 
        .Z(n6567) );
  CND2X1 U6982 ( .A(n7648), .B(\m04.DoutM [6]), .Z(n6566) );
  CND4X1 U6983 ( .A(n6569), .B(n6568), .C(n6567), .D(n6566), .Z(n7686) );
  CMX2X1 U6984 ( .A0(n7686), .A1(\s00.dbus_in [6]), .S(n7596), .Z(n5048) );
  CIVX2 U6985 ( .A(n6570), .Z(n6575) );
  CNR2X1 U6986 ( .A(\m01.addrM [7]), .B(\m01.addrM [8]), .Z(n6573) );
  COND3X1 U6987 ( .A(n6905), .B(n6907), .C(n6658), .D(n6571), .Z(n6572) );
  CANR2X1 U6988 ( .A(n6575), .B(n6574), .C(n6573), .D(n6572), .Z(n6578) );
  CNR3X1 U6989 ( .A(n6578), .B(n6577), .C(n6576), .Z(n7186) );
  CNR2X1 U6990 ( .A(n7577), .B(n6579), .Z(n6603) );
  CND2X1 U6991 ( .A(\m03.addrM [4]), .B(n6580), .Z(n7287) );
  CIVX2 U6992 ( .A(n6581), .Z(n6582) );
  COND3X1 U6993 ( .A(n7303), .B(n7287), .C(n6583), .D(n6582), .Z(n6586) );
  CNR2X1 U6994 ( .A(\m03.addrM [5]), .B(n7298), .Z(n6584) );
  CANR2X1 U6995 ( .A(n6587), .B(n6586), .C(n6585), .D(n6584), .Z(n6590) );
  CNR3X1 U6996 ( .A(n6590), .B(n6589), .C(n6588), .Z(n7507) );
  CANR2XL U6997 ( .A(n7560), .B(n7507), .C(n7581), .D(n6797), .Z(n6600) );
  CIVX2 U6998 ( .A(n6591), .Z(n6595) );
  CNR3XL U6999 ( .A(n6825), .B(n6595), .C(n6592), .Z(n6593) );
  CANR4CX1 U7000 ( .A(n6816), .B(n6595), .C(n6594), .D(n6593), .Z(n6598) );
  CNR3X1 U7001 ( .A(n6598), .B(n6597), .C(n6596), .Z(n7234) );
  CANR2XL U7002 ( .A(n7579), .B(n7234), .C(n7583), .D(n7272), .Z(n6599) );
  COND3X1 U7003 ( .A(n7589), .B(n6601), .C(n6600), .D(n6599), .Z(n6602) );
  CANR3X1 U7004 ( .A(n7186), .B(n7585), .C(n6603), .D(n6602), .Z(n7597) );
  CMX2X1 U7005 ( .A0(n7687), .A1(\s01.Adr [1]), .S(n7597), .Z(n4979) );
  CMX2X1 U7006 ( .A0(n7635), .A1(\s01.dbus_in [15]), .S(n7597), .Z(n4977) );
  CMX2X1 U7007 ( .A0(n7636), .A1(\s01.dbus_in [14]), .S(n7597), .Z(n4976) );
  CMX2X1 U7008 ( .A0(n7628), .A1(\s01.dbus_in [11]), .S(n7597), .Z(n4973) );
  CMX2X1 U7009 ( .A0(n7629), .A1(\s01.dbus_in [7]), .S(n7597), .Z(n4969) );
  CMX2X1 U7010 ( .A0(n7630), .A1(\s01.dbus_in [5]), .S(n7597), .Z(n4967) );
  CMX2X1 U7011 ( .A0(n7631), .A1(\s01.dbus_in [3]), .S(n7597), .Z(n4965) );
  CMX2X1 U7012 ( .A0(n7632), .A1(\s01.dbus_in [1]), .S(n7597), .Z(n4963) );
  CMX2X1 U7013 ( .A0(n7684), .A1(\s01.dbus_in [0]), .S(n7597), .Z(n4962) );
  CND2X1 U7014 ( .A(\m01.addrM [11]), .B(\m01.addrM [12]), .Z(n6611) );
  CIVX2 U7015 ( .A(n6604), .Z(n6610) );
  COND1XL U7016 ( .A(n6607), .B(n6606), .C(n6605), .Z(n6656) );
  CND2X1 U7017 ( .A(n6608), .B(n6656), .Z(n6609) );
  CNR4X1 U7018 ( .A(n6611), .B(n6902), .C(n6610), .D(n6609), .Z(n6612) );
  CNIVX1 U7019 ( .A(n6612), .Z(n7182) );
  CNR2X1 U7020 ( .A(n7589), .B(n6613), .Z(n6628) );
  CANR2XL U7021 ( .A(n7581), .B(n6788), .C(n7583), .D(n7267), .Z(n6625) );
  CANR1XL U7022 ( .A(\m03.addrM [3]), .B(n6614), .C(\m03.addrM [4]), .Z(n6618)
         );
  CND4X1 U7023 ( .A(\m03.addrM [12]), .B(\m03.addrM [11]), .C(n7315), .D(n6615), .Z(n6616) );
  CNR3X1 U7024 ( .A(n6618), .B(n6617), .C(n6616), .Z(n7498) );
  CND2IX1 U7025 ( .B(n6808), .A(n6845), .Z(n6622) );
  COND1XL U7026 ( .A(\m04.addrM [1]), .B(\m04.addrM [4]), .C(n6619), .Z(n6644)
         );
  CNR4X1 U7027 ( .A(n6622), .B(n6621), .C(n6644), .D(n6620), .Z(n6623) );
  CNIVX1 U7028 ( .A(n6623), .Z(n7241) );
  CANR2XL U7029 ( .A(n7560), .B(n7498), .C(n7579), .D(n7241), .Z(n6624) );
  COND3X1 U7030 ( .A(n7577), .B(n6626), .C(n6625), .D(n6624), .Z(n6627) );
  CANR3X1 U7031 ( .A(n7182), .B(n7585), .C(n6628), .D(n6627), .Z(n7598) );
  CMX2X1 U7032 ( .A0(n7687), .A1(\s02.Adr [1]), .S(n7598), .Z(n4915) );
  CMX2X1 U7033 ( .A0(n7625), .A1(\s02.Adr [0]), .S(n7598), .Z(n4914) );
  CMX2X1 U7034 ( .A0(n7636), .A1(\s02.dbus_in [14]), .S(n7598), .Z(n4912) );
  CMX2X1 U7035 ( .A0(n7637), .A1(\s02.dbus_in [12]), .S(n7598), .Z(n4910) );
  CMX2X1 U7036 ( .A0(n7626), .A1(\s02.dbus_in [10]), .S(n7598), .Z(n4908) );
  CANR2XL U7037 ( .A(\m00.YouGotIt ), .B(\m00.DoutM [9]), .C(n7642), .D(
        \m01.DoutM [9]), .Z(n6632) );
  CANR2X1 U7038 ( .A(n7644), .B(\m03.DoutM [9]), .C(n7643), .D(\m02.DoutM [9]), 
        .Z(n6631) );
  CANR2X1 U7039 ( .A(n7641), .B(\m05.DoutM [9]), .C(n7640), .D(\m06.DoutM [9]), 
        .Z(n6630) );
  CND2X1 U7040 ( .A(n7648), .B(\m04.DoutM [9]), .Z(n6629) );
  CND4X1 U7041 ( .A(n6632), .B(n6631), .C(n6630), .D(n6629), .Z(n7682) );
  CMX2X1 U7042 ( .A0(n7682), .A1(\s02.dbus_in [9]), .S(n7598), .Z(n4907) );
  CMX2X1 U7043 ( .A0(n7685), .A1(\s02.dbus_in [8]), .S(n7598), .Z(n4906) );
  CMX2X1 U7044 ( .A0(n7686), .A1(\s02.dbus_in [6]), .S(n7598), .Z(n4904) );
  CMX2X1 U7045 ( .A0(n7653), .A1(\s02.dbus_in [4]), .S(n7598), .Z(n4902) );
  CNR2X1 U7046 ( .A(n7298), .B(n6633), .Z(n6639) );
  CAN4X1 U7047 ( .A(n7307), .B(n6636), .C(n6635), .D(n6634), .Z(n6637) );
  CANR1XL U7048 ( .A(n6639), .B(n6638), .C(n6637), .Z(n6641) );
  CANR3X1 U7049 ( .A(n6641), .B(n7297), .C(n7302), .D(n6640), .Z(n7500) );
  CIVX2 U7050 ( .A(n6833), .Z(n6647) );
  CANR11X1 U7051 ( .A(n6645), .B(n6644), .C(n6643), .D(n6642), .Z(n6646) );
  CANR4CX1 U7052 ( .A(n6809), .B(n6647), .C(n6806), .D(n6646), .Z(n6648) );
  CND2X1 U7053 ( .A(n6808), .B(n6648), .Z(n6649) );
  CND3XL U7054 ( .A(n6650), .B(n6839), .C(n6649), .Z(n6823) );
  COND2X1 U7055 ( .A(n7577), .B(n6651), .C(n7539), .D(n6823), .Z(n6666) );
  CND2X1 U7056 ( .A(n6653), .B(n6652), .Z(n6655) );
  CANR4CX1 U7057 ( .A(n6656), .B(n6655), .C(n6654), .D(n6889), .Z(n6661) );
  CND2X1 U7058 ( .A(n6895), .B(n6657), .Z(n6921) );
  CNR2X1 U7059 ( .A(n6658), .B(n6921), .Z(n6932) );
  COND1XL U7060 ( .A(n6932), .B(n6896), .C(n6895), .Z(n6660) );
  CANR3X1 U7061 ( .A(n6661), .B(n6660), .C(n6659), .D(n6936), .Z(n7178) );
  CANR2X1 U7062 ( .A(n7585), .B(n7178), .C(n7583), .D(n7264), .Z(n6663) );
  CND2X1 U7063 ( .A(n7581), .B(n6782), .Z(n6662) );
  COND3X1 U7064 ( .A(n7589), .B(n6664), .C(n6663), .D(n6662), .Z(n6665) );
  CANR3X1 U7065 ( .A(n7560), .B(n7500), .C(n6666), .D(n6665), .Z(n7599) );
  CMX2X1 U7066 ( .A0(n7621), .A1(\s03.Adr [2]), .S(n7599), .Z(n4852) );
  CMX2X1 U7067 ( .A0(n7625), .A1(\s03.Adr [0]), .S(n7599), .Z(n4850) );
  CMX2X1 U7068 ( .A0(n7627), .A1(\s03.dbus_in [13]), .S(n7599), .Z(n4847) );
  CMX2X1 U7069 ( .A0(n7628), .A1(\s03.dbus_in [11]), .S(n7599), .Z(n4845) );
  CMX2X1 U7070 ( .A0(n7626), .A1(\s03.dbus_in [10]), .S(n7599), .Z(n4844) );
  CMX2X1 U7071 ( .A0(n7629), .A1(\s03.dbus_in [7]), .S(n7599), .Z(n4841) );
  CMX2X1 U7072 ( .A0(n7630), .A1(\s03.dbus_in [5]), .S(n7599), .Z(n4839) );
  CMX2X1 U7073 ( .A0(n7631), .A1(\s03.dbus_in [3]), .S(n7599), .Z(n4837) );
  CMX2X1 U7074 ( .A0(n7632), .A1(\s03.dbus_in [1]), .S(n7599), .Z(n4835) );
  CMX2X1 U7075 ( .A0(n7625), .A1(\s08.Adr [0]), .S(n7573), .Z(n4530) );
  CIVX2 U7076 ( .A(\s04.dataOut [9]), .Z(n7425) );
  CANR2X1 U7077 ( .A(n7678), .B(\s00.dataOut [9]), .C(\s08.dataOut [9]), .D(
        n7662), .Z(n6674) );
  CAOR2XL U7078 ( .A(\s01.dataOut [9]), .B(n7658), .C(\s09.dataOut [9]), .D(
        n7666), .Z(n6672) );
  CANR2XL U7079 ( .A(\s02.dataOut [9]), .B(n7660), .C(\s13.dataOut [9]), .D(
        n7661), .Z(n6670) );
  CANR2X1 U7080 ( .A(n7663), .B(\s03.dataOut [9]), .C(\s05.dataOut [9]), .D(
        n7657), .Z(n6669) );
  CANR2XL U7081 ( .A(\s07.dataOut [9]), .B(n7667), .C(\s10.dataOut [9]), .D(
        n6698), .Z(n6668) );
  CANR2X1 U7082 ( .A(\s12.dataOut [9]), .B(n7665), .C(\s06.dataOut [9]), .D(
        n7659), .Z(n6667) );
  CND4X1 U7083 ( .A(n6670), .B(n6669), .C(n6668), .D(n6667), .Z(n6671) );
  CANR3XL U7084 ( .A(\s11.dataOut [9]), .B(n7664), .C(n6672), .D(n6671), .Z(
        n6673) );
  COND3X1 U7085 ( .A(n7425), .B(n7576), .C(n6674), .D(n6673), .Z(n6675) );
  CMX2X1 U7086 ( .A0(\m06.DinMast [9]), .A1(n6675), .S(n7679), .Z(n5195) );
  CANR2XL U7087 ( .A(\s01.dataOut [7]), .B(n7658), .C(\s08.dataOut [7]), .D(
        n7662), .Z(n6685) );
  CIVX2 U7088 ( .A(\s00.dataOut [7]), .Z(n7405) );
  COND2X1 U7089 ( .A(n6677), .B(n7405), .C(n6676), .D(n7674), .Z(n6683) );
  CANR2X1 U7090 ( .A(n7663), .B(\s03.dataOut [7]), .C(\s02.dataOut [7]), .D(
        n7660), .Z(n6681) );
  CANR2X1 U7091 ( .A(\s04.dataOut [7]), .B(n7656), .C(\s05.dataOut [7]), .D(
        n7657), .Z(n6680) );
  CANR2X1 U7092 ( .A(\s09.dataOut [7]), .B(n7666), .C(\s07.dataOut [7]), .D(
        n7667), .Z(n6679) );
  CANR2X1 U7093 ( .A(\s06.dataOut [7]), .B(n7659), .C(\s11.dataOut [7]), .D(
        n7664), .Z(n6678) );
  CND4X1 U7094 ( .A(n6681), .B(n6680), .C(n6679), .D(n6678), .Z(n6682) );
  CANR3X1 U7095 ( .A(\s12.dataOut [7]), .B(n7665), .C(n6683), .D(n6682), .Z(
        n6684) );
  COND3X1 U7096 ( .A(n6687), .B(n6686), .C(n6685), .D(n6684), .Z(n6688) );
  CMX2X1 U7097 ( .A0(\m06.DinMast [7]), .A1(n6688), .S(n7679), .Z(n5193) );
  CANR2XL U7098 ( .A(\s01.dataOut [0]), .B(n6726), .C(\s09.dataOut [0]), .D(
        n6738), .Z(n6696) );
  CANR2XL U7099 ( .A(\s11.dataOut [0]), .B(n6733), .C(\s08.dataOut [0]), .D(
        n6736), .Z(n6695) );
  CANR2X1 U7100 ( .A(\s07.dataOut [0]), .B(n6729), .C(\s06.dataOut [0]), .D(
        n6730), .Z(n6694) );
  CANR2XL U7101 ( .A(\s05.dataOut [0]), .B(n6731), .C(\s04.dataOut [0]), .D(
        n6735), .Z(n6692) );
  CANR2X1 U7102 ( .A(\s12.dataOut [0]), .B(n6734), .C(\s10.dataOut [0]), .D(
        n6732), .Z(n6691) );
  CANR2X1 U7103 ( .A(\s13.dataOut [0]), .B(n6728), .C(\s02.dataOut [0]), .D(
        n6739), .Z(n6690) );
  CANR2X1 U7104 ( .A(n6737), .B(\s00.dataOut [0]), .C(n6727), .D(
        \s03.dataOut [0]), .Z(n6689) );
  CAN4X1 U7105 ( .A(n6692), .B(n6691), .C(n6690), .D(n6689), .Z(n6693) );
  CND4X1 U7106 ( .A(n6696), .B(n6695), .C(n6694), .D(n6693), .Z(n6697) );
  CMX2X1 U7107 ( .A0(\m05.DinMast [0]), .A1(n6697), .S(n6748), .Z(n4194) );
  CIVX2 U7108 ( .A(\s04.dataOut [6]), .Z(n7395) );
  CANR2XL U7109 ( .A(\s08.dataOut [6]), .B(n7662), .C(\s01.dataOut [6]), .D(
        n7658), .Z(n6706) );
  CAOR2X2 U7110 ( .A(\s09.dataOut [6]), .B(n7666), .C(\s10.dataOut [6]), .D(
        n6698), .Z(n6704) );
  CANR2XL U7111 ( .A(n7663), .B(\s03.dataOut [6]), .C(\s13.dataOut [6]), .D(
        n7661), .Z(n6702) );
  CANR2X1 U7112 ( .A(\s05.dataOut [6]), .B(n7657), .C(\s02.dataOut [6]), .D(
        n7660), .Z(n6701) );
  CANR2X1 U7113 ( .A(\s12.dataOut [6]), .B(n7665), .C(\s11.dataOut [6]), .D(
        n7664), .Z(n6700) );
  CANR2XL U7114 ( .A(\s06.dataOut [6]), .B(n7659), .C(\s07.dataOut [6]), .D(
        n7667), .Z(n6699) );
  CND4X1 U7115 ( .A(n6702), .B(n6701), .C(n6700), .D(n6699), .Z(n6703) );
  CANR3X1 U7116 ( .A(n7678), .B(\s00.dataOut [6]), .C(n6704), .D(n6703), .Z(
        n6705) );
  COND3X1 U7117 ( .A(n7395), .B(n7576), .C(n6706), .D(n6705), .Z(n6707) );
  CMX2X1 U7118 ( .A0(\m06.DinMast [6]), .A1(n6707), .S(n7679), .Z(n5192) );
  CANR2X1 U7119 ( .A(n6727), .B(\s03.dataOut [1]), .C(\s09.dataOut [1]), .D(
        n6738), .Z(n6715) );
  CANR2XL U7120 ( .A(\s12.dataOut [1]), .B(n6734), .C(\s04.dataOut [1]), .D(
        n6735), .Z(n6714) );
  CANR2XL U7121 ( .A(\s06.dataOut [1]), .B(n6730), .C(\s13.dataOut [1]), .D(
        n6728), .Z(n6713) );
  CANR2XL U7122 ( .A(\s05.dataOut [1]), .B(n6731), .C(\s11.dataOut [1]), .D(
        n6733), .Z(n6711) );
  CANR2XL U7123 ( .A(\s07.dataOut [1]), .B(n6729), .C(\s10.dataOut [1]), .D(
        n6732), .Z(n6710) );
  CANR2X1 U7124 ( .A(n6737), .B(\s00.dataOut [1]), .C(\s02.dataOut [1]), .D(
        n6739), .Z(n6709) );
  CANR2XL U7125 ( .A(\s08.dataOut [1]), .B(n6736), .C(\s01.dataOut [1]), .D(
        n6726), .Z(n6708) );
  CAN4X1 U7126 ( .A(n6711), .B(n6710), .C(n6709), .D(n6708), .Z(n6712) );
  CND4X1 U7127 ( .A(n6715), .B(n6714), .C(n6713), .D(n6712), .Z(n6716) );
  CMX2X1 U7128 ( .A0(\m05.DinMast [1]), .A1(n6716), .S(n6748), .Z(n4195) );
  CANR2X1 U7129 ( .A(n6727), .B(\s03.dataOut [2]), .C(\s01.dataOut [2]), .D(
        n6726), .Z(n6724) );
  CANR2X1 U7130 ( .A(\s07.dataOut [2]), .B(n6729), .C(\s08.dataOut [2]), .D(
        n6736), .Z(n6723) );
  CANR2XL U7131 ( .A(\s05.dataOut [2]), .B(n6731), .C(\s11.dataOut [2]), .D(
        n6733), .Z(n6722) );
  CANR2XL U7132 ( .A(\s04.dataOut [2]), .B(n6735), .C(\s10.dataOut [2]), .D(
        n6732), .Z(n6720) );
  CANR2X1 U7133 ( .A(\s06.dataOut [2]), .B(n6730), .C(\s12.dataOut [2]), .D(
        n6734), .Z(n6719) );
  CANR2XL U7134 ( .A(\s02.dataOut [2]), .B(n6739), .C(\s13.dataOut [2]), .D(
        n6728), .Z(n6718) );
  CANR2X1 U7135 ( .A(n6737), .B(\s00.dataOut [2]), .C(\s09.dataOut [2]), .D(
        n6738), .Z(n6717) );
  CAN4X1 U7136 ( .A(n6720), .B(n6719), .C(n6718), .D(n6717), .Z(n6721) );
  CND4X1 U7137 ( .A(n6724), .B(n6723), .C(n6722), .D(n6721), .Z(n6725) );
  CMX2X1 U7138 ( .A0(\m05.DinMast [2]), .A1(n6725), .S(n6748), .Z(n4196) );
  CANR2XL U7139 ( .A(n6727), .B(\s03.dataOut [3]), .C(\s01.dataOut [3]), .D(
        n6726), .Z(n6747) );
  CANR2XL U7140 ( .A(\s07.dataOut [3]), .B(n6729), .C(\s13.dataOut [3]), .D(
        n6728), .Z(n6746) );
  CANR2X1 U7141 ( .A(\s05.dataOut [3]), .B(n6731), .C(\s06.dataOut [3]), .D(
        n6730), .Z(n6745) );
  CANR2XL U7142 ( .A(\s11.dataOut [3]), .B(n6733), .C(\s10.dataOut [3]), .D(
        n6732), .Z(n6743) );
  CANR2XL U7143 ( .A(\s04.dataOut [3]), .B(n6735), .C(\s12.dataOut [3]), .D(
        n6734), .Z(n6742) );
  CANR2XL U7144 ( .A(n6737), .B(\s00.dataOut [3]), .C(\s08.dataOut [3]), .D(
        n6736), .Z(n6741) );
  CANR2X1 U7145 ( .A(\s02.dataOut [3]), .B(n6739), .C(\s09.dataOut [3]), .D(
        n6738), .Z(n6740) );
  CAN4X1 U7146 ( .A(n6743), .B(n6742), .C(n6741), .D(n6740), .Z(n6744) );
  CND4X1 U7147 ( .A(n6747), .B(n6746), .C(n6745), .D(n6744), .Z(n6749) );
  CMX2X1 U7148 ( .A0(\m05.DinMast [3]), .A1(n6749), .S(n6748), .Z(n4197) );
  CANR2X1 U7149 ( .A(n6783), .B(\s00.dataOut [15]), .C(n6782), .D(
        \s03.dataOut [15]), .Z(n6758) );
  CANR2X1 U7150 ( .A(\s12.dataOut [15]), .B(n6785), .C(\s10.dataOut [15]), .D(
        n6790), .Z(n6757) );
  CANR2X1 U7151 ( .A(\s04.dataOut [15]), .B(n7580), .C(\s07.dataOut [15]), .D(
        n6771), .Z(n6756) );
  CAOR2X2 U7152 ( .A(\s06.dataOut [15]), .B(n7532), .C(\s05.dataOut [15]), .D(
        n6789), .Z(n6754) );
  CIVX2 U7153 ( .A(\s11.dataOut [15]), .Z(n7437) );
  CANR2XL U7154 ( .A(\s02.dataOut [15]), .B(n6788), .C(\s13.dataOut [15]), .D(
        n6787), .Z(n6751) );
  CANR2XL U7155 ( .A(\s09.dataOut [15]), .B(n6784), .C(\s08.dataOut [15]), .D(
        n6791), .Z(n6750) );
  COND3X1 U7156 ( .A(n7437), .B(n6752), .C(n6751), .D(n6750), .Z(n6753) );
  CANR3XL U7157 ( .A(\s01.dataOut [15]), .B(n6797), .C(n6754), .D(n6753), .Z(
        n6755) );
  CND4X1 U7158 ( .A(n6758), .B(n6757), .C(n6756), .D(n6755), .Z(n6759) );
  CMX2X1 U7159 ( .A0(\m00.DinMast [15]), .A1(n6759), .S(n6802), .Z(n5041) );
  CANR2XL U7160 ( .A(n6783), .B(\s00.dataOut [14]), .C(n6782), .D(
        \s03.dataOut [14]), .Z(n6769) );
  CANR2X1 U7161 ( .A(\s12.dataOut [14]), .B(n6785), .C(\s10.dataOut [14]), .D(
        n6790), .Z(n6768) );
  CANR2X1 U7162 ( .A(\s09.dataOut [14]), .B(n6784), .C(\s11.dataOut [14]), .D(
        n6786), .Z(n6767) );
  CAOR2X2 U7163 ( .A(\s07.dataOut [14]), .B(n6771), .C(\s05.dataOut [14]), .D(
        n6789), .Z(n6765) );
  CIVXL U7164 ( .A(n6791), .Z(n6762) );
  CANR2XL U7165 ( .A(\s02.dataOut [14]), .B(n6788), .C(\s13.dataOut [14]), .D(
        n6787), .Z(n6761) );
  CANR2X1 U7166 ( .A(\s06.dataOut [14]), .B(n7532), .C(\s04.dataOut [14]), .D(
        n7580), .Z(n6760) );
  COND3X1 U7167 ( .A(n6763), .B(n6762), .C(n6761), .D(n6760), .Z(n6764) );
  CANR3XL U7168 ( .A(\s01.dataOut [14]), .B(n6797), .C(n6765), .D(n6764), .Z(
        n6766) );
  CND4X1 U7169 ( .A(n6769), .B(n6768), .C(n6767), .D(n6766), .Z(n6770) );
  CMX2X1 U7170 ( .A0(\m00.DinMast [14]), .A1(n6770), .S(n6802), .Z(n5040) );
  CANR2X1 U7171 ( .A(n6783), .B(\s00.dataOut [13]), .C(\s01.dataOut [13]), .D(
        n6797), .Z(n6780) );
  CANR2X1 U7172 ( .A(\s04.dataOut [13]), .B(n7580), .C(\s11.dataOut [13]), .D(
        n6786), .Z(n6779) );
  CANR2XL U7173 ( .A(\s06.dataOut [13]), .B(n7532), .C(\s08.dataOut [13]), .D(
        n6791), .Z(n6778) );
  CAOR2X2 U7174 ( .A(\s05.dataOut [13]), .B(n6789), .C(\s09.dataOut [13]), .D(
        n6784), .Z(n6776) );
  CIVX2 U7175 ( .A(\s10.dataOut [13]), .Z(n7483) );
  CANR2XL U7176 ( .A(\s02.dataOut [13]), .B(n6788), .C(\s13.dataOut [13]), .D(
        n6787), .Z(n6773) );
  CANR2X1 U7177 ( .A(\s07.dataOut [13]), .B(n6771), .C(\s12.dataOut [13]), .D(
        n6785), .Z(n6772) );
  COND3X1 U7178 ( .A(n7483), .B(n6774), .C(n6773), .D(n6772), .Z(n6775) );
  CANR3XL U7179 ( .A(n6782), .B(\s03.dataOut [13]), .C(n6776), .D(n6775), .Z(
        n6777) );
  CND4X1 U7180 ( .A(n6780), .B(n6779), .C(n6778), .D(n6777), .Z(n6781) );
  CMX2X1 U7181 ( .A0(\m00.DinMast [13]), .A1(n6781), .S(n6802), .Z(n5039) );
  CANR2XL U7182 ( .A(n6783), .B(\s00.dataOut [12]), .C(n6782), .D(
        \s03.dataOut [12]), .Z(n6801) );
  CANR2X1 U7183 ( .A(\s12.dataOut [12]), .B(n6785), .C(\s09.dataOut [12]), .D(
        n6784), .Z(n6800) );
  CANR2X1 U7184 ( .A(\s06.dataOut [12]), .B(n7532), .C(\s04.dataOut [12]), .D(
        n7580), .Z(n6799) );
  CAOR2XL U7185 ( .A(\s13.dataOut [12]), .B(n6787), .C(\s11.dataOut [12]), .D(
        n6786), .Z(n6796) );
  CIVX2 U7186 ( .A(\s07.dataOut [12]), .Z(n6794) );
  CANR2XL U7187 ( .A(\s05.dataOut [12]), .B(n6789), .C(\s02.dataOut [12]), .D(
        n6788), .Z(n6793) );
  CANR2XL U7188 ( .A(\s08.dataOut [12]), .B(n6791), .C(\s10.dataOut [12]), .D(
        n6790), .Z(n6792) );
  COND3X1 U7189 ( .A(n6794), .B(n7548), .C(n6793), .D(n6792), .Z(n6795) );
  CANR3XL U7190 ( .A(\s01.dataOut [12]), .B(n6797), .C(n6796), .D(n6795), .Z(
        n6798) );
  CND4X1 U7191 ( .A(n6801), .B(n6800), .C(n6799), .D(n6798), .Z(n6803) );
  CMX2X1 U7192 ( .A0(\m00.DinMast [12]), .A1(n6803), .S(n6802), .Z(n5038) );
  CIVX2 U7193 ( .A(n6804), .Z(n7235) );
  CANR2X1 U7194 ( .A(n7235), .B(\s00.dataOut [0]), .C(\s01.dataOut [0]), .D(
        n7234), .Z(n6864) );
  CND2X1 U7195 ( .A(\m04.addrM [15]), .B(\m04.addrM [13]), .Z(n6840) );
  CIVX2 U7196 ( .A(n6840), .Z(n6813) );
  CNR2X1 U7197 ( .A(\m04.addrM [10]), .B(n6805), .Z(n6811) );
  COND11X1 U7198 ( .A(n6827), .B(n6826), .C(n6814), .D(n6806), .Z(n6807) );
  COND4CX1 U7199 ( .A(n6809), .B(n6845), .C(n6808), .D(n6807), .Z(n6810) );
  CAN4X1 U7200 ( .A(n6813), .B(n6812), .C(n6811), .D(n6810), .Z(n7516) );
  CANR2X1 U7201 ( .A(\s05.dataOut [0]), .B(n7237), .C(\s12.dataOut [0]), .D(
        n7516), .Z(n6863) );
  CNR2X1 U7202 ( .A(n6815), .B(n6814), .Z(n6819) );
  CIVX2 U7203 ( .A(n6816), .Z(n6818) );
  CAOR2X2 U7204 ( .A(n6819), .B(n6818), .C(n6849), .D(n6817), .Z(n6822) );
  CND3XL U7205 ( .A(n6822), .B(n6821), .C(n6820), .Z(n7538) );
  CIVX2 U7206 ( .A(n7538), .Z(n7244) );
  CANR2XL U7207 ( .A(\s06.dataOut [0]), .B(n7244), .C(\s10.dataOut [0]), .D(
        n7243), .Z(n6862) );
  CIVX2 U7208 ( .A(n6823), .Z(n7240) );
  CIVX2 U7209 ( .A(n6824), .Z(n6837) );
  CIVX1 U7210 ( .A(n6825), .Z(n6836) );
  CNR2X1 U7211 ( .A(n6827), .B(n6826), .Z(n6834) );
  CIVX2 U7212 ( .A(n6828), .Z(n6829) );
  COND4CX1 U7213 ( .A(n6849), .B(n6846), .C(n6851), .D(n6829), .Z(n6832) );
  COND1XL U7214 ( .A(n6851), .B(n6838), .C(n6830), .Z(n6831) );
  COND3X1 U7215 ( .A(n6834), .B(n6833), .C(n6832), .D(n6831), .Z(n6835) );
  CANR3X1 U7216 ( .A(n6838), .B(n6837), .C(n6836), .D(n6835), .Z(n6843) );
  CIVX2 U7217 ( .A(n6839), .Z(n6841) );
  CNR4X2 U7218 ( .A(n6843), .B(n6842), .C(n6841), .D(n6840), .Z(n7554) );
  CANR2X1 U7219 ( .A(n7240), .B(\s03.dataOut [0]), .C(\s07.dataOut [0]), .D(
        n7554), .Z(n6860) );
  CANR2XL U7220 ( .A(\s13.dataOut [0]), .B(n7236), .C(\s08.dataOut [0]), .D(
        n7242), .Z(n6859) );
  CANR4CX1 U7221 ( .A(n6847), .B(n6846), .C(n6845), .D(n6844), .Z(n6850) );
  CANR2X1 U7222 ( .A(n6851), .B(n6850), .C(n6849), .D(n6848), .Z(n6856) );
  CIVX2 U7223 ( .A(n6852), .Z(n6853) );
  CNR4X2 U7224 ( .A(n6856), .B(n6855), .C(n6854), .D(n6853), .Z(n7578) );
  CANR2XL U7225 ( .A(\s04.dataOut [0]), .B(n7578), .C(\s02.dataOut [0]), .D(
        n7241), .Z(n6858) );
  CANR2X1 U7226 ( .A(\s11.dataOut [0]), .B(n7238), .C(\s09.dataOut [0]), .D(
        n7239), .Z(n6857) );
  CAN4X1 U7227 ( .A(n6860), .B(n6859), .C(n6858), .D(n6857), .Z(n6861) );
  CND4X1 U7228 ( .A(n6864), .B(n6863), .C(n6862), .D(n6861), .Z(n6871) );
  CNR4X1 U7229 ( .A(n7243), .B(n7244), .C(n7239), .D(n7516), .Z(n6870) );
  CNR4XL U7230 ( .A(n7236), .B(n7242), .C(n7578), .D(n7241), .Z(n6868) );
  CNR4XL U7231 ( .A(n7235), .B(n7240), .C(n7234), .D(n7554), .Z(n6867) );
  CAN4X1 U7232 ( .A(n6868), .B(n6867), .C(n6866), .D(n6865), .Z(n6869) );
  CANR1X2 U7233 ( .A(n6870), .B(n6869), .C(n7539), .Z(n7253) );
  CMX2X1 U7234 ( .A0(\m04.DinMast [0]), .A1(n6871), .S(n7253), .Z(n4210) );
  CANR2X1 U7235 ( .A(n7235), .B(\s00.dataOut [1]), .C(\s01.dataOut [1]), .D(
        n7234), .Z(n6880) );
  CANR2X1 U7236 ( .A(\s05.dataOut [1]), .B(n7237), .C(\s08.dataOut [1]), .D(
        n7242), .Z(n6879) );
  CANR2X1 U7237 ( .A(\s06.dataOut [1]), .B(n7244), .C(\s09.dataOut [1]), .D(
        n7239), .Z(n6878) );
  CAOR2XL U7238 ( .A(n7240), .B(\s03.dataOut [1]), .C(\s07.dataOut [1]), .D(
        n7554), .Z(n6876) );
  CIVX2 U7239 ( .A(\s10.dataOut [1]), .Z(n7342) );
  CANR2XL U7240 ( .A(\s12.dataOut [1]), .B(n7516), .C(\s02.dataOut [1]), .D(
        n7241), .Z(n6873) );
  CANR2XL U7241 ( .A(\s04.dataOut [1]), .B(n7578), .C(\s13.dataOut [1]), .D(
        n7236), .Z(n6872) );
  COND3X1 U7242 ( .A(n7342), .B(n6874), .C(n6873), .D(n6872), .Z(n6875) );
  CANR3X1 U7243 ( .A(\s11.dataOut [1]), .B(n7238), .C(n6876), .D(n6875), .Z(
        n6877) );
  CND4X1 U7244 ( .A(n6880), .B(n6879), .C(n6878), .D(n6877), .Z(n6881) );
  CMX2X1 U7245 ( .A0(\m04.DinMast [1]), .A1(n6881), .S(n7253), .Z(n4211) );
  CANR2XL U7246 ( .A(n7181), .B(\s00.dataOut [15]), .C(n7178), .D(
        \s03.dataOut [15]), .Z(n6946) );
  CND2X1 U7247 ( .A(n6896), .B(n6882), .Z(n6888) );
  CANR11X1 U7248 ( .A(n6885), .B(n6894), .C(n6884), .D(n6883), .Z(n6887) );
  COND4CX1 U7249 ( .A(n6889), .B(n6888), .C(n6887), .D(n6886), .Z(n6890) );
  CNR4X1 U7250 ( .A(\m01.addrM [10]), .B(n6892), .C(n6891), .D(n6890), .Z(
        n6893) );
  CNIVX1 U7251 ( .A(n6893), .Z(n7519) );
  CANR2XL U7252 ( .A(n7179), .B(\s05.dataOut [15]), .C(n7519), .D(
        \s12.dataOut [15]), .Z(n6945) );
  CND2X1 U7253 ( .A(n6895), .B(n6894), .Z(n6898) );
  COND2X1 U7254 ( .A(n6899), .B(n6898), .C(n6897), .D(n6896), .Z(n6900) );
  CIVX2 U7255 ( .A(n6900), .Z(n6903) );
  CNR3X1 U7256 ( .A(n6903), .B(n6902), .C(n6901), .Z(n7535) );
  CIVX2 U7257 ( .A(n6929), .Z(n6908) );
  CNR3XL U7258 ( .A(n6905), .B(n6914), .C(n6904), .Z(n6906) );
  CANR4CX1 U7259 ( .A(n6908), .B(n6907), .C(n6932), .D(n6906), .Z(n6913) );
  CIVX2 U7260 ( .A(n6909), .Z(n6912) );
  CNR4X2 U7261 ( .A(n6913), .B(n6912), .C(n6911), .D(n6910), .Z(n7584) );
  CANR2XL U7262 ( .A(n7535), .B(\s06.dataOut [15]), .C(n7584), .D(
        \s04.dataOut [15]), .Z(n6944) );
  CANR1XL U7263 ( .A(n6929), .B(n6915), .C(n6914), .Z(n6931) );
  CIVX2 U7264 ( .A(n6916), .Z(n6928) );
  CIVX2 U7265 ( .A(n6917), .Z(n6924) );
  CIVX2 U7266 ( .A(n6918), .Z(n6920) );
  COND1XL U7267 ( .A(n6921), .B(n6920), .C(n6919), .Z(n6922) );
  CANR3X1 U7268 ( .A(n6925), .B(n6924), .C(n6923), .D(n6922), .Z(n6926) );
  COND4CX1 U7269 ( .A(n6929), .B(n6928), .C(n6927), .D(n6926), .Z(n6930) );
  CANR3X1 U7270 ( .A(n6933), .B(n6932), .C(n6931), .D(n6930), .Z(n6937) );
  CND2X1 U7271 ( .A(\m01.addrM [16]), .B(\m01.addrM [15]), .Z(n6935) );
  CND2X1 U7272 ( .A(\m01.addrM [14]), .B(\m01.addrM [13]), .Z(n6934) );
  CNR4X1 U7273 ( .A(n6937), .B(n6936), .C(n6935), .D(n6934), .Z(n6938) );
  CNIVX1 U7274 ( .A(n6938), .Z(n7553) );
  CANR2XL U7275 ( .A(n7553), .B(\s07.dataOut [15]), .C(n7180), .D(
        \s10.dataOut [15]), .Z(n6942) );
  CANR2XL U7276 ( .A(n7183), .B(\s13.dataOut [15]), .C(n7182), .D(
        \s02.dataOut [15]), .Z(n6941) );
  CANR2XL U7277 ( .A(n7185), .B(\s08.dataOut [15]), .C(n7187), .D(
        \s11.dataOut [15]), .Z(n6940) );
  CANR2XL U7278 ( .A(n7186), .B(\s01.dataOut [15]), .C(n7184), .D(
        \s09.dataOut [15]), .Z(n6939) );
  CAN4X1 U7279 ( .A(n6942), .B(n6941), .C(n6940), .D(n6939), .Z(n6943) );
  CND4X1 U7280 ( .A(n6946), .B(n6945), .C(n6944), .D(n6943), .Z(n6952) );
  CNR4XL U7281 ( .A(n7535), .B(n7179), .C(n7584), .D(n7519), .Z(n6951) );
  CNR4XL U7282 ( .A(n7181), .B(n7178), .C(n6948), .D(n6947), .Z(n6950) );
  CIVX2 U7283 ( .A(n7585), .Z(n6949) );
  CANR1X2 U7284 ( .A(n6951), .B(n6950), .C(n6949), .Z(n7196) );
  CMX2X1 U7285 ( .A0(\m01.DinMast [15]), .A1(n6952), .S(n7196), .Z(n4273) );
  CANR2X1 U7286 ( .A(n7235), .B(\s00.dataOut [2]), .C(\s01.dataOut [2]), .D(
        n7234), .Z(n6960) );
  CANR2XL U7287 ( .A(\s13.dataOut [2]), .B(n7236), .C(\s11.dataOut [2]), .D(
        n7238), .Z(n6959) );
  CANR2XL U7288 ( .A(\s06.dataOut [2]), .B(n7244), .C(\s10.dataOut [2]), .D(
        n7243), .Z(n6958) );
  CANR2X1 U7289 ( .A(n7240), .B(\s03.dataOut [2]), .C(\s07.dataOut [2]), .D(
        n7554), .Z(n6956) );
  CANR2X1 U7290 ( .A(\s04.dataOut [2]), .B(n7578), .C(\s08.dataOut [2]), .D(
        n7242), .Z(n6955) );
  CANR2XL U7291 ( .A(\s12.dataOut [2]), .B(n7516), .C(\s02.dataOut [2]), .D(
        n7241), .Z(n6954) );
  CANR2X1 U7292 ( .A(\s05.dataOut [2]), .B(n7237), .C(\s09.dataOut [2]), .D(
        n7239), .Z(n6953) );
  CAN4X1 U7293 ( .A(n6956), .B(n6955), .C(n6954), .D(n6953), .Z(n6957) );
  CND4X1 U7294 ( .A(n6960), .B(n6959), .C(n6958), .D(n6957), .Z(n6961) );
  CMX2X1 U7295 ( .A0(\m04.DinMast [2]), .A1(n6961), .S(n7253), .Z(n4212) );
  CANR2XL U7296 ( .A(n7181), .B(\s00.dataOut [14]), .C(n7553), .D(
        \s07.dataOut [14]), .Z(n6969) );
  CANR2XL U7297 ( .A(n7535), .B(\s06.dataOut [14]), .C(n7584), .D(
        \s04.dataOut [14]), .Z(n6968) );
  CANR2XL U7298 ( .A(n7179), .B(\s05.dataOut [14]), .C(n7519), .D(
        \s12.dataOut [14]), .Z(n6967) );
  CANR2X1 U7299 ( .A(n7178), .B(\s03.dataOut [14]), .C(n7184), .D(
        \s09.dataOut [14]), .Z(n6965) );
  CANR2XL U7300 ( .A(n7183), .B(\s13.dataOut [14]), .C(n7182), .D(
        \s02.dataOut [14]), .Z(n6964) );
  CANR2XL U7301 ( .A(n7186), .B(\s01.dataOut [14]), .C(n7180), .D(
        \s10.dataOut [14]), .Z(n6963) );
  CANR2XL U7302 ( .A(n7185), .B(\s08.dataOut [14]), .C(n7187), .D(
        \s11.dataOut [14]), .Z(n6962) );
  CAN4X1 U7303 ( .A(n6965), .B(n6964), .C(n6963), .D(n6962), .Z(n6966) );
  CND4X1 U7304 ( .A(n6969), .B(n6968), .C(n6967), .D(n6966), .Z(n6970) );
  CMX2X1 U7305 ( .A0(\m01.DinMast [14]), .A1(n6970), .S(n7196), .Z(n4272) );
  CANR2X1 U7306 ( .A(n7235), .B(\s00.dataOut [3]), .C(\s01.dataOut [3]), .D(
        n7234), .Z(n6978) );
  CANR2X1 U7307 ( .A(\s08.dataOut [3]), .B(n7242), .C(\s09.dataOut [3]), .D(
        n7239), .Z(n6977) );
  CANR2XL U7308 ( .A(\s06.dataOut [3]), .B(n7244), .C(\s10.dataOut [3]), .D(
        n7243), .Z(n6976) );
  CANR2X1 U7309 ( .A(n7240), .B(\s03.dataOut [3]), .C(\s07.dataOut [3]), .D(
        n7554), .Z(n6974) );
  CANR2XL U7310 ( .A(\s02.dataOut [3]), .B(n7241), .C(\s13.dataOut [3]), .D(
        n7236), .Z(n6973) );
  CANR2X1 U7311 ( .A(\s04.dataOut [3]), .B(n7578), .C(\s12.dataOut [3]), .D(
        n7516), .Z(n6972) );
  CANR2X1 U7312 ( .A(\s05.dataOut [3]), .B(n7237), .C(\s11.dataOut [3]), .D(
        n7238), .Z(n6971) );
  CAN4X1 U7313 ( .A(n6974), .B(n6973), .C(n6972), .D(n6971), .Z(n6975) );
  CND4X1 U7314 ( .A(n6978), .B(n6977), .C(n6976), .D(n6975), .Z(n6979) );
  CMX2X1 U7315 ( .A0(\m04.DinMast [3]), .A1(n6979), .S(n7253), .Z(n4213) );
  CANR2XL U7316 ( .A(n7181), .B(\s00.dataOut [13]), .C(n7553), .D(
        \s07.dataOut [13]), .Z(n6987) );
  CANR2X1 U7317 ( .A(n7535), .B(\s06.dataOut [13]), .C(n7179), .D(
        \s05.dataOut [13]), .Z(n6986) );
  CANR2XL U7318 ( .A(n7584), .B(\s04.dataOut [13]), .C(n7519), .D(
        \s12.dataOut [13]), .Z(n6985) );
  CANR2XL U7319 ( .A(n7178), .B(\s03.dataOut [13]), .C(n7183), .D(
        \s13.dataOut [13]), .Z(n6983) );
  CANR2XL U7320 ( .A(n7182), .B(\s02.dataOut [13]), .C(n7187), .D(
        \s11.dataOut [13]), .Z(n6982) );
  CANR2XL U7321 ( .A(n7186), .B(\s01.dataOut [13]), .C(n7180), .D(
        \s10.dataOut [13]), .Z(n6981) );
  CANR2XL U7322 ( .A(n7185), .B(\s08.dataOut [13]), .C(n7184), .D(
        \s09.dataOut [13]), .Z(n6980) );
  CAN4X1 U7323 ( .A(n6983), .B(n6982), .C(n6981), .D(n6980), .Z(n6984) );
  CND4X1 U7324 ( .A(n6987), .B(n6986), .C(n6985), .D(n6984), .Z(n6988) );
  CMX2X1 U7325 ( .A0(\m01.DinMast [13]), .A1(n6988), .S(n7196), .Z(n4271) );
  CANR2XL U7326 ( .A(n7181), .B(\s00.dataOut [12]), .C(n7553), .D(
        \s07.dataOut [12]), .Z(n6996) );
  CANR2XL U7327 ( .A(n7179), .B(\s05.dataOut [12]), .C(n7584), .D(
        \s04.dataOut [12]), .Z(n6995) );
  CANR2XL U7328 ( .A(n7535), .B(\s06.dataOut [12]), .C(n7519), .D(
        \s12.dataOut [12]), .Z(n6994) );
  CANR2XL U7329 ( .A(n7178), .B(\s03.dataOut [12]), .C(n7187), .D(
        \s11.dataOut [12]), .Z(n6992) );
  CANR2XL U7330 ( .A(n7183), .B(\s13.dataOut [12]), .C(n7182), .D(
        \s02.dataOut [12]), .Z(n6991) );
  CANR2XL U7331 ( .A(n7185), .B(\s08.dataOut [12]), .C(n7180), .D(
        \s10.dataOut [12]), .Z(n6990) );
  CANR2XL U7332 ( .A(n7186), .B(\s01.dataOut [12]), .C(n7184), .D(
        \s09.dataOut [12]), .Z(n6989) );
  CAN4X1 U7333 ( .A(n6992), .B(n6991), .C(n6990), .D(n6989), .Z(n6993) );
  CND4X1 U7334 ( .A(n6996), .B(n6995), .C(n6994), .D(n6993), .Z(n6997) );
  CMX2X1 U7335 ( .A0(\m01.DinMast [12]), .A1(n6997), .S(n7196), .Z(n4270) );
  CANR2X1 U7336 ( .A(n7235), .B(\s00.dataOut [4]), .C(\s01.dataOut [4]), .D(
        n7234), .Z(n7005) );
  CANR2X1 U7337 ( .A(\s04.dataOut [4]), .B(n7578), .C(\s09.dataOut [4]), .D(
        n7239), .Z(n7004) );
  CANR2X1 U7338 ( .A(\s06.dataOut [4]), .B(n7244), .C(\s05.dataOut [4]), .D(
        n7237), .Z(n7003) );
  CANR2X1 U7339 ( .A(n7240), .B(\s03.dataOut [4]), .C(\s07.dataOut [4]), .D(
        n7554), .Z(n7001) );
  CANR2X1 U7340 ( .A(\s12.dataOut [4]), .B(n7516), .C(\s08.dataOut [4]), .D(
        n7242), .Z(n7000) );
  CANR2XL U7341 ( .A(\s13.dataOut [4]), .B(n7236), .C(\s02.dataOut [4]), .D(
        n7241), .Z(n6999) );
  CANR2XL U7342 ( .A(\s10.dataOut [4]), .B(n7243), .C(\s11.dataOut [4]), .D(
        n7238), .Z(n6998) );
  CAN4X1 U7343 ( .A(n7001), .B(n7000), .C(n6999), .D(n6998), .Z(n7002) );
  CND4X1 U7344 ( .A(n7005), .B(n7004), .C(n7003), .D(n7002), .Z(n7006) );
  CMX2X1 U7345 ( .A0(\m04.DinMast [4]), .A1(n7006), .S(n7253), .Z(n4214) );
  CANR2XL U7346 ( .A(n7181), .B(\s00.dataOut [11]), .C(n7178), .D(
        \s03.dataOut [11]), .Z(n7014) );
  CANR2XL U7347 ( .A(n7584), .B(\s04.dataOut [11]), .C(n7519), .D(
        \s12.dataOut [11]), .Z(n7013) );
  CANR2X1 U7348 ( .A(n7535), .B(\s06.dataOut [11]), .C(n7179), .D(
        \s05.dataOut [11]), .Z(n7012) );
  CANR2XL U7349 ( .A(n7553), .B(\s07.dataOut [11]), .C(n7182), .D(
        \s02.dataOut [11]), .Z(n7010) );
  CANR2XL U7350 ( .A(n7183), .B(\s13.dataOut [11]), .C(n7187), .D(
        \s11.dataOut [11]), .Z(n7009) );
  CANR2XL U7351 ( .A(n7186), .B(\s01.dataOut [11]), .C(n7184), .D(
        \s09.dataOut [11]), .Z(n7008) );
  CANR2XL U7352 ( .A(n7185), .B(\s08.dataOut [11]), .C(n7180), .D(
        \s10.dataOut [11]), .Z(n7007) );
  CAN4X1 U7353 ( .A(n7010), .B(n7009), .C(n7008), .D(n7007), .Z(n7011) );
  CND4X1 U7354 ( .A(n7014), .B(n7013), .C(n7012), .D(n7011), .Z(n7015) );
  CMX2X1 U7355 ( .A0(\m01.DinMast [11]), .A1(n7015), .S(n7196), .Z(n4269) );
  CANR2X1 U7356 ( .A(n7235), .B(\s00.dataOut [5]), .C(\s01.dataOut [5]), .D(
        n7234), .Z(n7023) );
  CANR2X1 U7357 ( .A(\s12.dataOut [5]), .B(n7516), .C(\s09.dataOut [5]), .D(
        n7239), .Z(n7022) );
  CANR2X1 U7358 ( .A(\s06.dataOut [5]), .B(n7244), .C(\s05.dataOut [5]), .D(
        n7237), .Z(n7021) );
  CANR2X1 U7359 ( .A(n7240), .B(\s03.dataOut [5]), .C(\s07.dataOut [5]), .D(
        n7554), .Z(n7019) );
  CANR2XL U7360 ( .A(\s13.dataOut [5]), .B(n7236), .C(\s08.dataOut [5]), .D(
        n7242), .Z(n7018) );
  CANR2XL U7361 ( .A(\s04.dataOut [5]), .B(n7578), .C(\s02.dataOut [5]), .D(
        n7241), .Z(n7017) );
  CANR2XL U7362 ( .A(\s10.dataOut [5]), .B(n7243), .C(\s11.dataOut [5]), .D(
        n7238), .Z(n7016) );
  CAN4X1 U7363 ( .A(n7019), .B(n7018), .C(n7017), .D(n7016), .Z(n7020) );
  CND4X1 U7364 ( .A(n7023), .B(n7022), .C(n7021), .D(n7020), .Z(n7024) );
  CMX2X1 U7365 ( .A0(\m04.DinMast [5]), .A1(n7024), .S(n7253), .Z(n4215) );
  CANR2XL U7366 ( .A(n7181), .B(\s00.dataOut [10]), .C(n7553), .D(
        \s07.dataOut [10]), .Z(n7032) );
  CANR2XL U7367 ( .A(n7535), .B(\s06.dataOut [10]), .C(n7519), .D(
        \s12.dataOut [10]), .Z(n7031) );
  CANR2XL U7368 ( .A(n7179), .B(\s05.dataOut [10]), .C(n7584), .D(
        \s04.dataOut [10]), .Z(n7030) );
  CANR2XL U7369 ( .A(n7178), .B(\s03.dataOut [10]), .C(n7183), .D(
        \s13.dataOut [10]), .Z(n7028) );
  CANR2XL U7370 ( .A(n7182), .B(\s02.dataOut [10]), .C(n7184), .D(
        \s09.dataOut [10]), .Z(n7027) );
  CANR2XL U7371 ( .A(n7185), .B(\s08.dataOut [10]), .C(n7180), .D(
        \s10.dataOut [10]), .Z(n7026) );
  CANR2XL U7372 ( .A(n7187), .B(\s11.dataOut [10]), .C(n7186), .D(
        \s01.dataOut [10]), .Z(n7025) );
  CAN4X1 U7373 ( .A(n7028), .B(n7027), .C(n7026), .D(n7025), .Z(n7029) );
  CND4X1 U7374 ( .A(n7032), .B(n7031), .C(n7030), .D(n7029), .Z(n7033) );
  CMX2X1 U7375 ( .A0(\m01.DinMast [10]), .A1(n7033), .S(n7196), .Z(n4268) );
  CANR2XL U7376 ( .A(n7235), .B(\s00.dataOut [6]), .C(\s01.dataOut [6]), .D(
        n7234), .Z(n7041) );
  CANR2X1 U7377 ( .A(\s12.dataOut [6]), .B(n7516), .C(\s09.dataOut [6]), .D(
        n7239), .Z(n7040) );
  CANR2XL U7378 ( .A(\s06.dataOut [6]), .B(n7244), .C(\s10.dataOut [6]), .D(
        n7243), .Z(n7039) );
  CANR2X1 U7379 ( .A(n7240), .B(\s03.dataOut [6]), .C(\s07.dataOut [6]), .D(
        n7554), .Z(n7037) );
  CANR2XL U7380 ( .A(\s02.dataOut [6]), .B(n7241), .C(\s08.dataOut [6]), .D(
        n7242), .Z(n7036) );
  CANR2X1 U7381 ( .A(\s04.dataOut [6]), .B(n7578), .C(\s13.dataOut [6]), .D(
        n7236), .Z(n7035) );
  CANR2X1 U7382 ( .A(\s05.dataOut [6]), .B(n7237), .C(\s11.dataOut [6]), .D(
        n7238), .Z(n7034) );
  CAN4X1 U7383 ( .A(n7037), .B(n7036), .C(n7035), .D(n7034), .Z(n7038) );
  CND4X1 U7384 ( .A(n7041), .B(n7040), .C(n7039), .D(n7038), .Z(n7042) );
  CMX2X1 U7385 ( .A0(\m04.DinMast [6]), .A1(n7042), .S(n7253), .Z(n4216) );
  CANR2XL U7386 ( .A(n7181), .B(\s00.dataOut [9]), .C(n7553), .D(
        \s07.dataOut [9]), .Z(n7050) );
  CANR2X1 U7387 ( .A(n7535), .B(\s06.dataOut [9]), .C(n7179), .D(
        \s05.dataOut [9]), .Z(n7049) );
  CANR2XL U7388 ( .A(n7584), .B(\s04.dataOut [9]), .C(n7519), .D(
        \s12.dataOut [9]), .Z(n7048) );
  CANR2XL U7389 ( .A(n7183), .B(\s13.dataOut [9]), .C(n7182), .D(
        \s02.dataOut [9]), .Z(n7046) );
  CANR2XL U7390 ( .A(n7178), .B(\s03.dataOut [9]), .C(n7187), .D(
        \s11.dataOut [9]), .Z(n7045) );
  CANR2XL U7391 ( .A(n7184), .B(\s09.dataOut [9]), .C(n7180), .D(
        \s10.dataOut [9]), .Z(n7044) );
  CANR2XL U7392 ( .A(n7185), .B(\s08.dataOut [9]), .C(n7186), .D(
        \s01.dataOut [9]), .Z(n7043) );
  CAN4X1 U7393 ( .A(n7046), .B(n7045), .C(n7044), .D(n7043), .Z(n7047) );
  CND4X1 U7394 ( .A(n7050), .B(n7049), .C(n7048), .D(n7047), .Z(n7051) );
  CMX2X1 U7395 ( .A0(\m01.DinMast [9]), .A1(n7051), .S(n7196), .Z(n4267) );
  CANR2XL U7396 ( .A(n7181), .B(\s00.dataOut [8]), .C(n7553), .D(
        \s07.dataOut [8]), .Z(n7059) );
  CANR2XL U7397 ( .A(n7535), .B(\s06.dataOut [8]), .C(n7584), .D(
        \s04.dataOut [8]), .Z(n7058) );
  CANR2XL U7398 ( .A(n7179), .B(\s05.dataOut [8]), .C(n7519), .D(
        \s12.dataOut [8]), .Z(n7057) );
  CANR2XL U7399 ( .A(n7178), .B(\s03.dataOut [8]), .C(n7185), .D(
        \s08.dataOut [8]), .Z(n7055) );
  CANR2XL U7400 ( .A(n7183), .B(\s13.dataOut [8]), .C(n7182), .D(
        \s02.dataOut [8]), .Z(n7054) );
  CANR2XL U7401 ( .A(n7187), .B(\s11.dataOut [8]), .C(n7180), .D(
        \s10.dataOut [8]), .Z(n7053) );
  CANR2XL U7402 ( .A(n7186), .B(\s01.dataOut [8]), .C(n7184), .D(
        \s09.dataOut [8]), .Z(n7052) );
  CAN4X1 U7403 ( .A(n7055), .B(n7054), .C(n7053), .D(n7052), .Z(n7056) );
  CND4X1 U7404 ( .A(n7059), .B(n7058), .C(n7057), .D(n7056), .Z(n7060) );
  CMX2X1 U7405 ( .A0(\m01.DinMast [8]), .A1(n7060), .S(n7196), .Z(n4266) );
  CANR2XL U7406 ( .A(n7235), .B(\s00.dataOut [7]), .C(\s01.dataOut [7]), .D(
        n7234), .Z(n7068) );
  CANR2XL U7407 ( .A(\s06.dataOut [7]), .B(n7244), .C(\s02.dataOut [7]), .D(
        n7241), .Z(n7067) );
  CANR2X1 U7408 ( .A(\s10.dataOut [7]), .B(n7243), .C(\s11.dataOut [7]), .D(
        n7238), .Z(n7066) );
  CANR2X1 U7409 ( .A(n7240), .B(\s03.dataOut [7]), .C(\s07.dataOut [7]), .D(
        n7554), .Z(n7064) );
  CANR2X1 U7410 ( .A(\s04.dataOut [7]), .B(n7578), .C(\s08.dataOut [7]), .D(
        n7242), .Z(n7063) );
  CANR2XL U7411 ( .A(\s12.dataOut [7]), .B(n7516), .C(\s13.dataOut [7]), .D(
        n7236), .Z(n7062) );
  CANR2X1 U7412 ( .A(\s05.dataOut [7]), .B(n7237), .C(\s09.dataOut [7]), .D(
        n7239), .Z(n7061) );
  CAN4X1 U7413 ( .A(n7064), .B(n7063), .C(n7062), .D(n7061), .Z(n7065) );
  CND4X1 U7414 ( .A(n7068), .B(n7067), .C(n7066), .D(n7065), .Z(n7069) );
  CMX2X1 U7415 ( .A0(\m04.DinMast [7]), .A1(n7069), .S(n7253), .Z(n4217) );
  CANR2XL U7416 ( .A(n7181), .B(\s00.dataOut [7]), .C(n7178), .D(
        \s03.dataOut [7]), .Z(n7077) );
  CANR2XL U7417 ( .A(n7535), .B(\s06.dataOut [7]), .C(n7519), .D(
        \s12.dataOut [7]), .Z(n7076) );
  CANR2XL U7418 ( .A(n7179), .B(\s05.dataOut [7]), .C(n7584), .D(
        \s04.dataOut [7]), .Z(n7075) );
  CANR2XL U7419 ( .A(n7183), .B(\s13.dataOut [7]), .C(n7553), .D(
        \s07.dataOut [7]), .Z(n7073) );
  CANR2XL U7420 ( .A(n7182), .B(\s02.dataOut [7]), .C(n7184), .D(
        \s09.dataOut [7]), .Z(n7072) );
  CANR2XL U7421 ( .A(n7187), .B(\s11.dataOut [7]), .C(n7180), .D(
        \s10.dataOut [7]), .Z(n7071) );
  CANR2XL U7422 ( .A(n7185), .B(\s08.dataOut [7]), .C(n7186), .D(
        \s01.dataOut [7]), .Z(n7070) );
  CAN4X1 U7423 ( .A(n7073), .B(n7072), .C(n7071), .D(n7070), .Z(n7074) );
  CND4X1 U7424 ( .A(n7077), .B(n7076), .C(n7075), .D(n7074), .Z(n7078) );
  CMX2X1 U7425 ( .A0(\m01.DinMast [7]), .A1(n7078), .S(n7196), .Z(n4265) );
  CANR2XL U7426 ( .A(n7235), .B(\s00.dataOut [8]), .C(\s01.dataOut [8]), .D(
        n7234), .Z(n7086) );
  CANR2XL U7427 ( .A(\s02.dataOut [8]), .B(n7241), .C(\s10.dataOut [8]), .D(
        n7243), .Z(n7085) );
  CANR2X1 U7428 ( .A(\s05.dataOut [8]), .B(n7237), .C(\s09.dataOut [8]), .D(
        n7239), .Z(n7084) );
  CANR2X1 U7429 ( .A(n7240), .B(\s03.dataOut [8]), .C(\s07.dataOut [8]), .D(
        n7554), .Z(n7082) );
  CANR2X1 U7430 ( .A(\s12.dataOut [8]), .B(n7516), .C(\s04.dataOut [8]), .D(
        n7578), .Z(n7081) );
  CANR2XL U7431 ( .A(\s13.dataOut [8]), .B(n7236), .C(\s08.dataOut [8]), .D(
        n7242), .Z(n7080) );
  CANR2X1 U7432 ( .A(\s06.dataOut [8]), .B(n7244), .C(\s11.dataOut [8]), .D(
        n7238), .Z(n7079) );
  CAN4X1 U7433 ( .A(n7082), .B(n7081), .C(n7080), .D(n7079), .Z(n7083) );
  CND4X1 U7434 ( .A(n7086), .B(n7085), .C(n7084), .D(n7083), .Z(n7087) );
  CMX2X1 U7435 ( .A0(\m04.DinMast [8]), .A1(n7087), .S(n7253), .Z(n4218) );
  CANR2XL U7436 ( .A(n7181), .B(\s00.dataOut [6]), .C(n7178), .D(
        \s03.dataOut [6]), .Z(n7095) );
  CANR2XL U7437 ( .A(n7179), .B(\s05.dataOut [6]), .C(n7584), .D(
        \s04.dataOut [6]), .Z(n7094) );
  CANR2XL U7438 ( .A(n7535), .B(\s06.dataOut [6]), .C(n7519), .D(
        \s12.dataOut [6]), .Z(n7093) );
  CANR2XL U7439 ( .A(n7183), .B(\s13.dataOut [6]), .C(n7182), .D(
        \s02.dataOut [6]), .Z(n7091) );
  CANR2XL U7440 ( .A(n7553), .B(\s07.dataOut [6]), .C(n7184), .D(
        \s09.dataOut [6]), .Z(n7090) );
  CANR2XL U7441 ( .A(n7187), .B(\s11.dataOut [6]), .C(n7186), .D(
        \s01.dataOut [6]), .Z(n7089) );
  CANR2XL U7442 ( .A(n7185), .B(\s08.dataOut [6]), .C(n7180), .D(
        \s10.dataOut [6]), .Z(n7088) );
  CAN4X1 U7443 ( .A(n7091), .B(n7090), .C(n7089), .D(n7088), .Z(n7092) );
  CND4X1 U7444 ( .A(n7095), .B(n7094), .C(n7093), .D(n7092), .Z(n7096) );
  CMX2X1 U7445 ( .A0(\m01.DinMast [6]), .A1(n7096), .S(n7196), .Z(n4264) );
  CANR2XL U7446 ( .A(n7235), .B(\s00.dataOut [9]), .C(\s01.dataOut [9]), .D(
        n7234), .Z(n7104) );
  CANR2XL U7447 ( .A(\s05.dataOut [9]), .B(n7237), .C(\s02.dataOut [9]), .D(
        n7241), .Z(n7103) );
  CANR2X1 U7448 ( .A(\s11.dataOut [9]), .B(n7238), .C(\s09.dataOut [9]), .D(
        n7239), .Z(n7102) );
  CANR2X1 U7449 ( .A(n7240), .B(\s03.dataOut [9]), .C(\s07.dataOut [9]), .D(
        n7554), .Z(n7100) );
  CANR2XL U7450 ( .A(\s13.dataOut [9]), .B(n7236), .C(\s08.dataOut [9]), .D(
        n7242), .Z(n7099) );
  CANR2X1 U7451 ( .A(\s12.dataOut [9]), .B(n7516), .C(\s04.dataOut [9]), .D(
        n7578), .Z(n7098) );
  CANR2XL U7452 ( .A(\s06.dataOut [9]), .B(n7244), .C(\s10.dataOut [9]), .D(
        n7243), .Z(n7097) );
  CAN4X1 U7453 ( .A(n7100), .B(n7099), .C(n7098), .D(n7097), .Z(n7101) );
  CND4X1 U7454 ( .A(n7104), .B(n7103), .C(n7102), .D(n7101), .Z(n7105) );
  CMX2X1 U7455 ( .A0(\m04.DinMast [9]), .A1(n7105), .S(n7253), .Z(n4219) );
  CANR2XL U7456 ( .A(n7178), .B(\s03.dataOut [5]), .C(n7553), .D(
        \s07.dataOut [5]), .Z(n7113) );
  CANR2XL U7457 ( .A(n7584), .B(\s04.dataOut [5]), .C(n7519), .D(
        \s12.dataOut [5]), .Z(n7112) );
  CANR2XL U7458 ( .A(n7535), .B(\s06.dataOut [5]), .C(n7179), .D(
        \s05.dataOut [5]), .Z(n7111) );
  CANR2XL U7459 ( .A(n7181), .B(\s00.dataOut [5]), .C(n7182), .D(
        \s02.dataOut [5]), .Z(n7109) );
  CANR2XL U7460 ( .A(n7183), .B(\s13.dataOut [5]), .C(n7186), .D(
        \s01.dataOut [5]), .Z(n7108) );
  CANR2XL U7461 ( .A(n7187), .B(\s11.dataOut [5]), .C(n7180), .D(
        \s10.dataOut [5]), .Z(n7107) );
  CANR2XL U7462 ( .A(n7185), .B(\s08.dataOut [5]), .C(n7184), .D(
        \s09.dataOut [5]), .Z(n7106) );
  CAN4X1 U7463 ( .A(n7109), .B(n7108), .C(n7107), .D(n7106), .Z(n7110) );
  CND4X1 U7464 ( .A(n7113), .B(n7112), .C(n7111), .D(n7110), .Z(n7114) );
  CMX2X1 U7465 ( .A0(\m01.DinMast [5]), .A1(n7114), .S(n7196), .Z(n4263) );
  CANR2XL U7466 ( .A(n7181), .B(\s00.dataOut [4]), .C(n7178), .D(
        \s03.dataOut [4]), .Z(n7122) );
  CANR2XL U7467 ( .A(n7179), .B(\s05.dataOut [4]), .C(n7519), .D(
        \s12.dataOut [4]), .Z(n7121) );
  CANR2X1 U7468 ( .A(n7535), .B(\s06.dataOut [4]), .C(n7584), .D(
        \s04.dataOut [4]), .Z(n7120) );
  CANR2XL U7469 ( .A(n7553), .B(\s07.dataOut [4]), .C(n7180), .D(
        \s10.dataOut [4]), .Z(n7118) );
  CANR2XL U7470 ( .A(n7183), .B(\s13.dataOut [4]), .C(n7182), .D(
        \s02.dataOut [4]), .Z(n7117) );
  CANR2XL U7471 ( .A(n7187), .B(\s11.dataOut [4]), .C(n7186), .D(
        \s01.dataOut [4]), .Z(n7116) );
  CANR2XL U7472 ( .A(n7185), .B(\s08.dataOut [4]), .C(n7184), .D(
        \s09.dataOut [4]), .Z(n7115) );
  CAN4X1 U7473 ( .A(n7118), .B(n7117), .C(n7116), .D(n7115), .Z(n7119) );
  CND4X1 U7474 ( .A(n7122), .B(n7121), .C(n7120), .D(n7119), .Z(n7123) );
  CMX2X1 U7475 ( .A0(\m01.DinMast [4]), .A1(n7123), .S(n7196), .Z(n4262) );
  CANR2XL U7476 ( .A(n7235), .B(\s00.dataOut [10]), .C(\s01.dataOut [10]), .D(
        n7234), .Z(n7131) );
  CANR2XL U7477 ( .A(\s02.dataOut [10]), .B(n7241), .C(\s10.dataOut [10]), .D(
        n7243), .Z(n7130) );
  CANR2X1 U7478 ( .A(\s09.dataOut [10]), .B(n7239), .C(\s11.dataOut [10]), .D(
        n7238), .Z(n7129) );
  CANR2X1 U7479 ( .A(n7240), .B(\s03.dataOut [10]), .C(\s07.dataOut [10]), .D(
        n7554), .Z(n7127) );
  CANR2X1 U7480 ( .A(\s04.dataOut [10]), .B(n7578), .C(\s08.dataOut [10]), .D(
        n7242), .Z(n7126) );
  CANR2XL U7481 ( .A(\s12.dataOut [10]), .B(n7516), .C(\s13.dataOut [10]), .D(
        n7236), .Z(n7125) );
  CANR2X1 U7482 ( .A(\s05.dataOut [10]), .B(n7237), .C(\s06.dataOut [10]), .D(
        n7244), .Z(n7124) );
  CAN4X1 U7483 ( .A(n7127), .B(n7126), .C(n7125), .D(n7124), .Z(n7128) );
  CND4X1 U7484 ( .A(n7131), .B(n7130), .C(n7129), .D(n7128), .Z(n7132) );
  CMX2X1 U7485 ( .A0(\m04.DinMast [10]), .A1(n7132), .S(n7253), .Z(n4220) );
  CANR2XL U7486 ( .A(n7181), .B(\s00.dataOut [3]), .C(n7553), .D(
        \s07.dataOut [3]), .Z(n7140) );
  CANR2XL U7487 ( .A(n7535), .B(\s06.dataOut [3]), .C(n7519), .D(
        \s12.dataOut [3]), .Z(n7139) );
  CANR2X1 U7488 ( .A(n7179), .B(\s05.dataOut [3]), .C(n7584), .D(
        \s04.dataOut [3]), .Z(n7138) );
  CANR2XL U7489 ( .A(n7183), .B(\s13.dataOut [3]), .C(n7182), .D(
        \s02.dataOut [3]), .Z(n7136) );
  CANR2XL U7490 ( .A(n7178), .B(\s03.dataOut [3]), .C(n7186), .D(
        \s01.dataOut [3]), .Z(n7135) );
  CANR2XL U7491 ( .A(n7184), .B(\s09.dataOut [3]), .C(n7180), .D(
        \s10.dataOut [3]), .Z(n7134) );
  CANR2XL U7492 ( .A(n7185), .B(\s08.dataOut [3]), .C(n7187), .D(
        \s11.dataOut [3]), .Z(n7133) );
  CAN4X1 U7493 ( .A(n7136), .B(n7135), .C(n7134), .D(n7133), .Z(n7137) );
  CND4X1 U7494 ( .A(n7140), .B(n7139), .C(n7138), .D(n7137), .Z(n7141) );
  CMX2X1 U7495 ( .A0(\m01.DinMast [3]), .A1(n7141), .S(n7196), .Z(n4261) );
  CANR2XL U7496 ( .A(n7235), .B(\s00.dataOut [11]), .C(\s01.dataOut [11]), .D(
        n7234), .Z(n7149) );
  CANR2X1 U7497 ( .A(\s06.dataOut [11]), .B(n7244), .C(\s04.dataOut [11]), .D(
        n7578), .Z(n7148) );
  CANR2X1 U7498 ( .A(\s05.dataOut [11]), .B(n7237), .C(\s10.dataOut [11]), .D(
        n7243), .Z(n7147) );
  CANR2X1 U7499 ( .A(n7240), .B(\s03.dataOut [11]), .C(\s07.dataOut [11]), .D(
        n7554), .Z(n7145) );
  CANR2XL U7500 ( .A(\s13.dataOut [11]), .B(n7236), .C(\s08.dataOut [11]), .D(
        n7242), .Z(n7144) );
  CANR2XL U7501 ( .A(\s12.dataOut [11]), .B(n7516), .C(\s02.dataOut [11]), .D(
        n7241), .Z(n7143) );
  CANR2X1 U7502 ( .A(\s11.dataOut [11]), .B(n7238), .C(\s09.dataOut [11]), .D(
        n7239), .Z(n7142) );
  CAN4X1 U7503 ( .A(n7145), .B(n7144), .C(n7143), .D(n7142), .Z(n7146) );
  CND4X1 U7504 ( .A(n7149), .B(n7148), .C(n7147), .D(n7146), .Z(n7150) );
  CMX2X1 U7505 ( .A0(\m04.DinMast [11]), .A1(n7150), .S(n7253), .Z(n4221) );
  CANR2XL U7506 ( .A(n7181), .B(\s00.dataOut [2]), .C(n7178), .D(
        \s03.dataOut [2]), .Z(n7158) );
  CANR2X1 U7507 ( .A(n7179), .B(\s05.dataOut [2]), .C(n7584), .D(
        \s04.dataOut [2]), .Z(n7157) );
  CANR2XL U7508 ( .A(n7535), .B(\s06.dataOut [2]), .C(n7519), .D(
        \s12.dataOut [2]), .Z(n7156) );
  CANR2XL U7509 ( .A(n7553), .B(\s07.dataOut [2]), .C(n7180), .D(
        \s10.dataOut [2]), .Z(n7154) );
  CANR2XL U7510 ( .A(n7183), .B(\s13.dataOut [2]), .C(n7182), .D(
        \s02.dataOut [2]), .Z(n7153) );
  CANR2XL U7511 ( .A(n7186), .B(\s01.dataOut [2]), .C(n7184), .D(
        \s09.dataOut [2]), .Z(n7152) );
  CANR2XL U7512 ( .A(n7185), .B(\s08.dataOut [2]), .C(n7187), .D(
        \s11.dataOut [2]), .Z(n7151) );
  CAN4X1 U7513 ( .A(n7154), .B(n7153), .C(n7152), .D(n7151), .Z(n7155) );
  CND4X1 U7514 ( .A(n7158), .B(n7157), .C(n7156), .D(n7155), .Z(n7159) );
  CMX2X1 U7515 ( .A0(\m01.DinMast [2]), .A1(n7159), .S(n7196), .Z(n4260) );
  CANR2XL U7516 ( .A(n7235), .B(\s00.dataOut [12]), .C(\s01.dataOut [12]), .D(
        n7234), .Z(n7167) );
  CANR2X1 U7517 ( .A(\s06.dataOut [12]), .B(n7244), .C(\s12.dataOut [12]), .D(
        n7516), .Z(n7166) );
  CANR2X1 U7518 ( .A(\s05.dataOut [12]), .B(n7237), .C(\s09.dataOut [12]), .D(
        n7239), .Z(n7165) );
  CANR2X1 U7519 ( .A(n7240), .B(\s03.dataOut [12]), .C(\s07.dataOut [12]), .D(
        n7554), .Z(n7163) );
  CANR2XL U7520 ( .A(\s13.dataOut [12]), .B(n7236), .C(\s08.dataOut [12]), .D(
        n7242), .Z(n7162) );
  CANR2XL U7521 ( .A(\s04.dataOut [12]), .B(n7578), .C(\s02.dataOut [12]), .D(
        n7241), .Z(n7161) );
  CANR2X1 U7522 ( .A(\s11.dataOut [12]), .B(n7238), .C(\s10.dataOut [12]), .D(
        n7243), .Z(n7160) );
  CAN4X1 U7523 ( .A(n7163), .B(n7162), .C(n7161), .D(n7160), .Z(n7164) );
  CND4X1 U7524 ( .A(n7167), .B(n7166), .C(n7165), .D(n7164), .Z(n7168) );
  CMX2X1 U7525 ( .A0(\m04.DinMast [12]), .A1(n7168), .S(n7253), .Z(n4222) );
  CANR2XL U7526 ( .A(n7178), .B(\s03.dataOut [1]), .C(n7553), .D(
        \s07.dataOut [1]), .Z(n7176) );
  CANR2X1 U7527 ( .A(n7535), .B(\s06.dataOut [1]), .C(n7584), .D(
        \s04.dataOut [1]), .Z(n7175) );
  CANR2XL U7528 ( .A(n7179), .B(\s05.dataOut [1]), .C(n7519), .D(
        \s12.dataOut [1]), .Z(n7174) );
  CANR2XL U7529 ( .A(n7181), .B(\s00.dataOut [1]), .C(n7182), .D(
        \s02.dataOut [1]), .Z(n7172) );
  CANR2XL U7530 ( .A(n7183), .B(\s13.dataOut [1]), .C(n7180), .D(
        \s10.dataOut [1]), .Z(n7171) );
  CANR2XL U7531 ( .A(n7185), .B(\s08.dataOut [1]), .C(n7186), .D(
        \s01.dataOut [1]), .Z(n7170) );
  CANR2XL U7532 ( .A(n7187), .B(\s11.dataOut [1]), .C(n7184), .D(
        \s09.dataOut [1]), .Z(n7169) );
  CAN4X1 U7533 ( .A(n7172), .B(n7171), .C(n7170), .D(n7169), .Z(n7173) );
  CND4X1 U7534 ( .A(n7176), .B(n7175), .C(n7174), .D(n7173), .Z(n7177) );
  CMX2X1 U7535 ( .A0(\m01.DinMast [1]), .A1(n7177), .S(n7196), .Z(n4259) );
  CANR2XL U7536 ( .A(n7178), .B(\s03.dataOut [0]), .C(n7553), .D(
        \s07.dataOut [0]), .Z(n7195) );
  CANR2XL U7537 ( .A(n7535), .B(\s06.dataOut [0]), .C(n7519), .D(
        \s12.dataOut [0]), .Z(n7194) );
  CANR2X1 U7538 ( .A(n7179), .B(\s05.dataOut [0]), .C(n7584), .D(
        \s04.dataOut [0]), .Z(n7193) );
  CANR2XL U7539 ( .A(n7181), .B(\s00.dataOut [0]), .C(n7180), .D(
        \s10.dataOut [0]), .Z(n7191) );
  CANR2XL U7540 ( .A(n7183), .B(\s13.dataOut [0]), .C(n7182), .D(
        \s02.dataOut [0]), .Z(n7190) );
  CANR2XL U7541 ( .A(n7185), .B(\s08.dataOut [0]), .C(n7184), .D(
        \s09.dataOut [0]), .Z(n7189) );
  CANR2XL U7542 ( .A(n7187), .B(\s11.dataOut [0]), .C(n7186), .D(
        \s01.dataOut [0]), .Z(n7188) );
  CAN4X1 U7543 ( .A(n7191), .B(n7190), .C(n7189), .D(n7188), .Z(n7192) );
  CND4X1 U7544 ( .A(n7195), .B(n7194), .C(n7193), .D(n7192), .Z(n7197) );
  CMX2X1 U7545 ( .A0(\m01.DinMast [0]), .A1(n7197), .S(n7196), .Z(n4258) );
  CANR2XL U7546 ( .A(n7235), .B(\s00.dataOut [13]), .C(\s01.dataOut [13]), .D(
        n7234), .Z(n7205) );
  CANR2X1 U7547 ( .A(\s05.dataOut [13]), .B(n7237), .C(\s08.dataOut [13]), .D(
        n7242), .Z(n7204) );
  CANR2X1 U7548 ( .A(\s11.dataOut [13]), .B(n7238), .C(\s10.dataOut [13]), .D(
        n7243), .Z(n7203) );
  CANR2X1 U7549 ( .A(n7240), .B(\s03.dataOut [13]), .C(\s07.dataOut [13]), .D(
        n7554), .Z(n7201) );
  CANR2XL U7550 ( .A(\s04.dataOut [13]), .B(n7578), .C(\s13.dataOut [13]), .D(
        n7236), .Z(n7200) );
  CANR2XL U7551 ( .A(\s12.dataOut [13]), .B(n7516), .C(\s02.dataOut [13]), .D(
        n7241), .Z(n7199) );
  CANR2X1 U7552 ( .A(\s06.dataOut [13]), .B(n7244), .C(\s09.dataOut [13]), .D(
        n7239), .Z(n7198) );
  CAN4X1 U7553 ( .A(n7201), .B(n7200), .C(n7199), .D(n7198), .Z(n7202) );
  CND4X1 U7554 ( .A(n7205), .B(n7204), .C(n7203), .D(n7202), .Z(n7206) );
  CMX2X1 U7555 ( .A0(\m04.DinMast [13]), .A1(n7206), .S(n7253), .Z(n4223) );
  CANR2XL U7556 ( .A(n7265), .B(\s00.dataOut [15]), .C(n7264), .D(
        \s03.dataOut [15]), .Z(n7214) );
  CANR2XL U7557 ( .A(\s12.dataOut [15]), .B(n7518), .C(\s02.dataOut [15]), .D(
        n7267), .Z(n7213) );
  CANR2XL U7558 ( .A(\s04.dataOut [15]), .B(n7582), .C(\s08.dataOut [15]), .D(
        n7266), .Z(n7212) );
  CANR2XL U7559 ( .A(\s05.dataOut [15]), .B(n7269), .C(\s13.dataOut [15]), .D(
        n7270), .Z(n7210) );
  CANR2XL U7560 ( .A(\s06.dataOut [15]), .B(n7534), .C(\s07.dataOut [15]), .D(
        n7552), .Z(n7209) );
  CANR2XL U7561 ( .A(\s10.dataOut [15]), .B(n7268), .C(\s01.dataOut [15]), .D(
        n7272), .Z(n7208) );
  CANR2XL U7562 ( .A(\s09.dataOut [15]), .B(n7271), .C(\s11.dataOut [15]), .D(
        n7273), .Z(n7207) );
  CAN4X1 U7563 ( .A(n7210), .B(n7209), .C(n7208), .D(n7207), .Z(n7211) );
  CND4X1 U7564 ( .A(n7214), .B(n7213), .C(n7212), .D(n7211), .Z(n7215) );
  CMX2X1 U7565 ( .A0(\m02.DinMast [15]), .A1(n7215), .S(n7282), .Z(n4257) );
  CANR2XL U7566 ( .A(n7235), .B(\s00.dataOut [14]), .C(\s01.dataOut [14]), .D(
        n7234), .Z(n7223) );
  CANR2X1 U7567 ( .A(\s06.dataOut [14]), .B(n7244), .C(\s08.dataOut [14]), .D(
        n7242), .Z(n7222) );
  CANR2X1 U7568 ( .A(\s09.dataOut [14]), .B(n7239), .C(\s11.dataOut [14]), .D(
        n7238), .Z(n7221) );
  CANR2X1 U7569 ( .A(n7240), .B(\s03.dataOut [14]), .C(\s07.dataOut [14]), .D(
        n7554), .Z(n7219) );
  CANR2XL U7570 ( .A(\s02.dataOut [14]), .B(n7241), .C(\s13.dataOut [14]), .D(
        n7236), .Z(n7218) );
  CANR2X1 U7571 ( .A(\s12.dataOut [14]), .B(n7516), .C(\s04.dataOut [14]), .D(
        n7578), .Z(n7217) );
  CANR2X1 U7572 ( .A(\s05.dataOut [14]), .B(n7237), .C(\s10.dataOut [14]), .D(
        n7243), .Z(n7216) );
  CAN4X1 U7573 ( .A(n7219), .B(n7218), .C(n7217), .D(n7216), .Z(n7220) );
  CND4X1 U7574 ( .A(n7223), .B(n7222), .C(n7221), .D(n7220), .Z(n7224) );
  CMX2X1 U7575 ( .A0(\m04.DinMast [14]), .A1(n7224), .S(n7253), .Z(n4224) );
  CANR2XL U7576 ( .A(n7265), .B(\s00.dataOut [14]), .C(n7264), .D(
        \s03.dataOut [14]), .Z(n7232) );
  CANR2XL U7577 ( .A(\s07.dataOut [14]), .B(n7552), .C(\s12.dataOut [14]), .D(
        n7518), .Z(n7231) );
  CANR2XL U7578 ( .A(\s02.dataOut [14]), .B(n7267), .C(\s13.dataOut [14]), .D(
        n7270), .Z(n7230) );
  CANR2XL U7579 ( .A(\s04.dataOut [14]), .B(n7582), .C(\s08.dataOut [14]), .D(
        n7266), .Z(n7228) );
  CANR2XL U7580 ( .A(\s06.dataOut [14]), .B(n7534), .C(\s10.dataOut [14]), .D(
        n7268), .Z(n7227) );
  CANR2XL U7581 ( .A(\s05.dataOut [14]), .B(n7269), .C(\s11.dataOut [14]), .D(
        n7273), .Z(n7226) );
  CANR2X1 U7582 ( .A(\s09.dataOut [14]), .B(n7271), .C(\s01.dataOut [14]), .D(
        n7272), .Z(n7225) );
  CAN4X1 U7583 ( .A(n7228), .B(n7227), .C(n7226), .D(n7225), .Z(n7229) );
  CND4X1 U7584 ( .A(n7232), .B(n7231), .C(n7230), .D(n7229), .Z(n7233) );
  CMX2X1 U7585 ( .A0(\m02.DinMast [14]), .A1(n7233), .S(n7282), .Z(n4256) );
  CANR2XL U7586 ( .A(n7235), .B(\s00.dataOut [15]), .C(\s01.dataOut [15]), .D(
        n7234), .Z(n7252) );
  CANR2XL U7587 ( .A(\s05.dataOut [15]), .B(n7237), .C(\s13.dataOut [15]), .D(
        n7236), .Z(n7251) );
  CANR2X1 U7588 ( .A(\s09.dataOut [15]), .B(n7239), .C(\s11.dataOut [15]), .D(
        n7238), .Z(n7250) );
  CANR2X1 U7589 ( .A(n7240), .B(\s03.dataOut [15]), .C(\s07.dataOut [15]), .D(
        n7554), .Z(n7248) );
  CANR2XL U7590 ( .A(\s04.dataOut [15]), .B(n7578), .C(\s02.dataOut [15]), .D(
        n7241), .Z(n7247) );
  CANR2X1 U7591 ( .A(\s12.dataOut [15]), .B(n7516), .C(\s08.dataOut [15]), .D(
        n7242), .Z(n7246) );
  CANR2X1 U7592 ( .A(\s06.dataOut [15]), .B(n7244), .C(\s10.dataOut [15]), .D(
        n7243), .Z(n7245) );
  CAN4X1 U7593 ( .A(n7248), .B(n7247), .C(n7246), .D(n7245), .Z(n7249) );
  CND4X1 U7594 ( .A(n7252), .B(n7251), .C(n7250), .D(n7249), .Z(n7254) );
  CMX2X1 U7595 ( .A0(\m04.DinMast [15]), .A1(n7254), .S(n7253), .Z(n4225) );
  CANR2XL U7596 ( .A(n7265), .B(\s00.dataOut [13]), .C(n7264), .D(
        \s03.dataOut [13]), .Z(n7262) );
  CANR2XL U7597 ( .A(\s13.dataOut [13]), .B(n7270), .C(\s10.dataOut [13]), .D(
        n7268), .Z(n7261) );
  CANR2XL U7598 ( .A(\s12.dataOut [13]), .B(n7518), .C(\s02.dataOut [13]), .D(
        n7267), .Z(n7260) );
  CANR2XL U7599 ( .A(\s05.dataOut [13]), .B(n7269), .C(\s08.dataOut [13]), .D(
        n7266), .Z(n7258) );
  CANR2XL U7600 ( .A(\s04.dataOut [13]), .B(n7582), .C(\s06.dataOut [13]), .D(
        n7534), .Z(n7257) );
  CANR2XL U7601 ( .A(\s07.dataOut [13]), .B(n7552), .C(\s09.dataOut [13]), .D(
        n7271), .Z(n7256) );
  CANR2XL U7602 ( .A(\s11.dataOut [13]), .B(n7273), .C(\s01.dataOut [13]), .D(
        n7272), .Z(n7255) );
  CAN4X1 U7603 ( .A(n7258), .B(n7257), .C(n7256), .D(n7255), .Z(n7259) );
  CND4X1 U7604 ( .A(n7262), .B(n7261), .C(n7260), .D(n7259), .Z(n7263) );
  CMX2X1 U7605 ( .A0(\m02.DinMast [13]), .A1(n7263), .S(n7282), .Z(n4255) );
  CANR2XL U7606 ( .A(n7265), .B(\s00.dataOut [12]), .C(n7264), .D(
        \s03.dataOut [12]), .Z(n7281) );
  CANR2XL U7607 ( .A(\s02.dataOut [12]), .B(n7267), .C(\s08.dataOut [12]), .D(
        n7266), .Z(n7280) );
  CANR2XL U7608 ( .A(\s05.dataOut [12]), .B(n7269), .C(\s10.dataOut [12]), .D(
        n7268), .Z(n7279) );
  CANR2XL U7609 ( .A(\s12.dataOut [12]), .B(n7518), .C(\s04.dataOut [12]), .D(
        n7582), .Z(n7277) );
  CANR2XL U7610 ( .A(\s06.dataOut [12]), .B(n7534), .C(\s13.dataOut [12]), .D(
        n7270), .Z(n7276) );
  CANR2XL U7611 ( .A(\s07.dataOut [12]), .B(n7552), .C(\s09.dataOut [12]), .D(
        n7271), .Z(n7275) );
  CANR2XL U7612 ( .A(\s11.dataOut [12]), .B(n7273), .C(\s01.dataOut [12]), .D(
        n7272), .Z(n7274) );
  CAN4X1 U7613 ( .A(n7277), .B(n7276), .C(n7275), .D(n7274), .Z(n7278) );
  CND4X1 U7614 ( .A(n7281), .B(n7280), .C(n7279), .D(n7278), .Z(n7283) );
  CMX2X1 U7615 ( .A0(\m02.DinMast [12]), .A1(n7283), .S(n7282), .Z(n4254) );
  CANR2XL U7616 ( .A(\s01.dataOut [0]), .B(n7507), .C(\s09.dataOut [0]), .D(
        n7504), .Z(n7332) );
  CANR2XL U7617 ( .A(n7500), .B(\s03.dataOut [0]), .C(\s13.dataOut [0]), .D(
        n7499), .Z(n7331) );
  CIVX2 U7618 ( .A(n7471), .Z(n7495) );
  CIVX2 U7619 ( .A(n7284), .Z(n7291) );
  CIVX2 U7620 ( .A(n7285), .Z(n7312) );
  CNR2X1 U7621 ( .A(n7317), .B(n7312), .Z(n7286) );
  COND1XL U7622 ( .A(\m03.addrM [5]), .B(n7287), .C(n7286), .Z(n7288) );
  COND11X1 U7623 ( .A(n7291), .B(n7290), .C(n7289), .D(n7288), .Z(n7292) );
  CND3XL U7624 ( .A(n7294), .B(n7293), .C(n7292), .Z(n7574) );
  CIVX2 U7625 ( .A(n7574), .Z(n7467) );
  CANR2X1 U7626 ( .A(n7495), .B(\s00.dataOut [0]), .C(\s04.dataOut [0]), .D(
        n7467), .Z(n7330) );
  CAN2X1 U7627 ( .A(n7296), .B(n7295), .Z(n7318) );
  CIVX2 U7628 ( .A(n7484), .Z(n7559) );
  CIVX2 U7629 ( .A(n7497), .Z(n7458) );
  CANR2XL U7630 ( .A(\s02.dataOut [0]), .B(n7498), .C(\s08.dataOut [0]), .D(
        n7496), .Z(n7325) );
  CND2X1 U7631 ( .A(n7304), .B(n7303), .Z(n7314) );
  CAOR2X2 U7632 ( .A(n7307), .B(n7306), .C(n7305), .D(n7314), .Z(n7311) );
  CIVX2 U7633 ( .A(n7308), .Z(n7321) );
  CAN4X1 U7634 ( .A(n7311), .B(n7321), .C(n7310), .D(n7309), .Z(n7533) );
  CANR2X1 U7635 ( .A(n7315), .B(n7314), .C(n7313), .D(n7312), .Z(n7316) );
  COND4CX1 U7636 ( .A(n7319), .B(n7318), .C(n7317), .D(n7316), .Z(n7320) );
  CAN4X1 U7637 ( .A(n7323), .B(n7322), .C(n7321), .D(n7320), .Z(n7517) );
  CANR2X1 U7638 ( .A(\s06.dataOut [0]), .B(n7533), .C(\s12.dataOut [0]), .D(
        n7517), .Z(n7324) );
  COND3X1 U7639 ( .A(n7326), .B(n7458), .C(n7325), .D(n7324), .Z(n7328) );
  CAOR2X2 U7640 ( .A(\s10.dataOut [0]), .B(n7493), .C(\s11.dataOut [0]), .D(
        n7494), .Z(n7327) );
  CANR3X1 U7641 ( .A(\s07.dataOut [0]), .B(n7559), .C(n7328), .D(n7327), .Z(
        n7329) );
  CND4X1 U7642 ( .A(n7332), .B(n7331), .C(n7330), .D(n7329), .Z(n7337) );
  CNR3XL U7643 ( .A(n7500), .B(n7496), .C(n7517), .Z(n7336) );
  COR4XL U7644 ( .A(n7495), .B(n7497), .C(n7499), .D(n7498), .Z(n7333) );
  COR4XL U7645 ( .A(n7507), .B(n7493), .C(n7533), .D(n7333), .Z(n7334) );
  CNR4XL U7646 ( .A(n7494), .B(n7504), .C(n7559), .D(n7334), .Z(n7335) );
  CANR11X2 U7647 ( .A(n7336), .B(n7335), .C(n7574), .D(n7575), .Z(n7512) );
  CMX2X1 U7648 ( .A0(\m03.DinMast [0]), .A1(n7337), .S(n7512), .Z(n4226) );
  CANR2X1 U7649 ( .A(\s11.dataOut [1]), .B(n7494), .C(\s09.dataOut [1]), .D(
        n7504), .Z(n7349) );
  CANR2XL U7650 ( .A(\s05.dataOut [1]), .B(n7497), .C(\s08.dataOut [1]), .D(
        n7496), .Z(n7348) );
  CANR2X1 U7651 ( .A(n7495), .B(\s00.dataOut [1]), .C(\s04.dataOut [1]), .D(
        n7467), .Z(n7347) );
  CIVXL U7652 ( .A(n7500), .Z(n7341) );
  CANR2XL U7653 ( .A(\s13.dataOut [1]), .B(n7499), .C(\s02.dataOut [1]), .D(
        n7498), .Z(n7339) );
  CANR2X1 U7654 ( .A(\s12.dataOut [1]), .B(n7517), .C(\s06.dataOut [1]), .D(
        n7533), .Z(n7338) );
  COND3X1 U7655 ( .A(n7341), .B(n7340), .C(n7339), .D(n7338), .Z(n7345) );
  CIVX2 U7656 ( .A(n7493), .Z(n7482) );
  COND2X1 U7657 ( .A(n7343), .B(n7484), .C(n7342), .D(n7482), .Z(n7344) );
  CANR3X1 U7658 ( .A(\s01.dataOut [1]), .B(n7507), .C(n7345), .D(n7344), .Z(
        n7346) );
  CND4X1 U7659 ( .A(n7349), .B(n7348), .C(n7347), .D(n7346), .Z(n7350) );
  CMX2X1 U7660 ( .A0(\m03.DinMast [1]), .A1(n7350), .S(n7512), .Z(n4227) );
  CANR2X1 U7661 ( .A(\s11.dataOut [2]), .B(n7494), .C(\s09.dataOut [2]), .D(
        n7504), .Z(n7359) );
  CANR2XL U7662 ( .A(n7500), .B(\s03.dataOut [2]), .C(\s08.dataOut [2]), .D(
        n7496), .Z(n7358) );
  CANR2X1 U7663 ( .A(\s12.dataOut [2]), .B(n7517), .C(\s05.dataOut [2]), .D(
        n7497), .Z(n7357) );
  CANR2XL U7664 ( .A(\s02.dataOut [2]), .B(n7498), .C(\s13.dataOut [2]), .D(
        n7499), .Z(n7352) );
  CANR2X1 U7665 ( .A(\s06.dataOut [2]), .B(n7533), .C(\s04.dataOut [2]), .D(
        n7467), .Z(n7351) );
  COND3X1 U7666 ( .A(n7471), .B(n7353), .C(n7352), .D(n7351), .Z(n7355) );
  CAOR2X2 U7667 ( .A(\s10.dataOut [2]), .B(n7493), .C(\s07.dataOut [2]), .D(
        n7559), .Z(n7354) );
  CANR3XL U7668 ( .A(\s01.dataOut [2]), .B(n7507), .C(n7355), .D(n7354), .Z(
        n7356) );
  CND4X1 U7669 ( .A(n7359), .B(n7358), .C(n7357), .D(n7356), .Z(n7360) );
  CMX2X1 U7670 ( .A0(\m03.DinMast [2]), .A1(n7360), .S(n7512), .Z(n4228) );
  CANR2XL U7671 ( .A(\s01.dataOut [3]), .B(n7507), .C(\s10.dataOut [3]), .D(
        n7493), .Z(n7369) );
  CANR2XL U7672 ( .A(\s06.dataOut [3]), .B(n7533), .C(\s08.dataOut [3]), .D(
        n7496), .Z(n7368) );
  CANR2XL U7673 ( .A(n7495), .B(\s00.dataOut [3]), .C(n7500), .D(
        \s03.dataOut [3]), .Z(n7367) );
  CANR2XL U7674 ( .A(\s02.dataOut [3]), .B(n7498), .C(\s13.dataOut [3]), .D(
        n7499), .Z(n7362) );
  CANR2X1 U7675 ( .A(\s04.dataOut [3]), .B(n7467), .C(\s12.dataOut [3]), .D(
        n7517), .Z(n7361) );
  COND3X1 U7676 ( .A(n7363), .B(n7458), .C(n7362), .D(n7361), .Z(n7365) );
  CAOR2X2 U7677 ( .A(\s11.dataOut [3]), .B(n7494), .C(\s09.dataOut [3]), .D(
        n7504), .Z(n7364) );
  CANR3X1 U7678 ( .A(\s07.dataOut [3]), .B(n7559), .C(n7365), .D(n7364), .Z(
        n7366) );
  CND4X1 U7679 ( .A(n7369), .B(n7368), .C(n7367), .D(n7366), .Z(n7370) );
  CMX2X1 U7680 ( .A0(\m03.DinMast [3]), .A1(n7370), .S(n7512), .Z(n4229) );
  CANR2X1 U7681 ( .A(\s11.dataOut [4]), .B(n7494), .C(\s01.dataOut [4]), .D(
        n7507), .Z(n7379) );
  CANR2XL U7682 ( .A(\s12.dataOut [4]), .B(n7517), .C(\s08.dataOut [4]), .D(
        n7496), .Z(n7378) );
  CANR2XL U7683 ( .A(n7500), .B(\s03.dataOut [4]), .C(\s06.dataOut [4]), .D(
        n7533), .Z(n7377) );
  CIVX2 U7684 ( .A(\s00.dataOut [4]), .Z(n7373) );
  CANR2XL U7685 ( .A(\s13.dataOut [4]), .B(n7499), .C(\s02.dataOut [4]), .D(
        n7498), .Z(n7372) );
  CANR2X1 U7686 ( .A(\s04.dataOut [4]), .B(n7467), .C(\s05.dataOut [4]), .D(
        n7497), .Z(n7371) );
  COND3X1 U7687 ( .A(n7471), .B(n7373), .C(n7372), .D(n7371), .Z(n7375) );
  CAOR2X2 U7688 ( .A(\s10.dataOut [4]), .B(n7493), .C(\s09.dataOut [4]), .D(
        n7504), .Z(n7374) );
  CANR3X1 U7689 ( .A(\s07.dataOut [4]), .B(n7559), .C(n7375), .D(n7374), .Z(
        n7376) );
  CND4X1 U7690 ( .A(n7379), .B(n7378), .C(n7377), .D(n7376), .Z(n7380) );
  CMX2X1 U7691 ( .A0(\m03.DinMast [4]), .A1(n7380), .S(n7512), .Z(n4230) );
  CANR2XL U7692 ( .A(\s09.dataOut [5]), .B(n7504), .C(\s10.dataOut [5]), .D(
        n7493), .Z(n7391) );
  CANR2X1 U7693 ( .A(\s12.dataOut [5]), .B(n7517), .C(\s13.dataOut [5]), .D(
        n7499), .Z(n7390) );
  CANR2XL U7694 ( .A(n7500), .B(\s03.dataOut [5]), .C(\s05.dataOut [5]), .D(
        n7497), .Z(n7389) );
  CANR2XL U7695 ( .A(\s02.dataOut [5]), .B(n7498), .C(\s08.dataOut [5]), .D(
        n7496), .Z(n7382) );
  CANR2X1 U7696 ( .A(\s06.dataOut [5]), .B(n7533), .C(\s04.dataOut [5]), .D(
        n7467), .Z(n7381) );
  COND3X1 U7697 ( .A(n7471), .B(n7383), .C(n7382), .D(n7381), .Z(n7387) );
  COND2X1 U7698 ( .A(n7385), .B(n7484), .C(n7384), .D(n7436), .Z(n7386) );
  CANR3XL U7699 ( .A(\s01.dataOut [5]), .B(n7507), .C(n7387), .D(n7386), .Z(
        n7388) );
  CND4X1 U7700 ( .A(n7391), .B(n7390), .C(n7389), .D(n7388), .Z(n7392) );
  CMX2X1 U7701 ( .A0(\m03.DinMast [5]), .A1(n7392), .S(n7512), .Z(n4231) );
  CANR2X1 U7702 ( .A(\s11.dataOut [6]), .B(n7494), .C(\s01.dataOut [6]), .D(
        n7507), .Z(n7401) );
  CANR2XL U7703 ( .A(n7500), .B(\s03.dataOut [6]), .C(\s08.dataOut [6]), .D(
        n7496), .Z(n7400) );
  CANR2X1 U7704 ( .A(n7495), .B(\s00.dataOut [6]), .C(\s05.dataOut [6]), .D(
        n7497), .Z(n7399) );
  CANR2XL U7705 ( .A(\s02.dataOut [6]), .B(n7498), .C(\s13.dataOut [6]), .D(
        n7499), .Z(n7394) );
  CANR2X1 U7706 ( .A(\s12.dataOut [6]), .B(n7517), .C(\s06.dataOut [6]), .D(
        n7533), .Z(n7393) );
  COND3X1 U7707 ( .A(n7395), .B(n7574), .C(n7394), .D(n7393), .Z(n7397) );
  CAOR2X2 U7708 ( .A(\s07.dataOut [6]), .B(n7559), .C(\s10.dataOut [6]), .D(
        n7493), .Z(n7396) );
  CANR3X1 U7709 ( .A(\s09.dataOut [6]), .B(n7504), .C(n7397), .D(n7396), .Z(
        n7398) );
  CND4X1 U7710 ( .A(n7401), .B(n7400), .C(n7399), .D(n7398), .Z(n7402) );
  CMX2X1 U7711 ( .A0(\m03.DinMast [6]), .A1(n7402), .S(n7512), .Z(n4232) );
  CANR2X1 U7712 ( .A(\s01.dataOut [7]), .B(n7507), .C(\s11.dataOut [7]), .D(
        n7494), .Z(n7411) );
  CANR2XL U7713 ( .A(n7500), .B(\s03.dataOut [7]), .C(\s13.dataOut [7]), .D(
        n7499), .Z(n7410) );
  CANR2X1 U7714 ( .A(\s04.dataOut [7]), .B(n7467), .C(\s06.dataOut [7]), .D(
        n7533), .Z(n7409) );
  CANR2XL U7715 ( .A(\s02.dataOut [7]), .B(n7498), .C(\s08.dataOut [7]), .D(
        n7496), .Z(n7404) );
  CANR2X1 U7716 ( .A(\s05.dataOut [7]), .B(n7497), .C(\s12.dataOut [7]), .D(
        n7517), .Z(n7403) );
  COND3X1 U7717 ( .A(n7471), .B(n7405), .C(n7404), .D(n7403), .Z(n7407) );
  CAOR2X2 U7718 ( .A(\s07.dataOut [7]), .B(n7559), .C(\s10.dataOut [7]), .D(
        n7493), .Z(n7406) );
  CANR3X1 U7719 ( .A(\s09.dataOut [7]), .B(n7504), .C(n7407), .D(n7406), .Z(
        n7408) );
  CND4X1 U7720 ( .A(n7411), .B(n7410), .C(n7409), .D(n7408), .Z(n7412) );
  CMX2X1 U7721 ( .A0(\m03.DinMast [7]), .A1(n7412), .S(n7512), .Z(n4233) );
  CANR2X1 U7722 ( .A(\s09.dataOut [8]), .B(n7504), .C(\s11.dataOut [8]), .D(
        n7494), .Z(n7421) );
  CANR2XL U7723 ( .A(\s12.dataOut [8]), .B(n7517), .C(\s08.dataOut [8]), .D(
        n7496), .Z(n7420) );
  CANR2X1 U7724 ( .A(n7495), .B(\s00.dataOut [8]), .C(\s04.dataOut [8]), .D(
        n7467), .Z(n7419) );
  CIVX2 U7725 ( .A(\s05.dataOut [8]), .Z(n7415) );
  CANR2XL U7726 ( .A(\s13.dataOut [8]), .B(n7499), .C(\s02.dataOut [8]), .D(
        n7498), .Z(n7414) );
  CANR2XL U7727 ( .A(n7500), .B(\s03.dataOut [8]), .C(\s06.dataOut [8]), .D(
        n7533), .Z(n7413) );
  COND3X1 U7728 ( .A(n7415), .B(n7458), .C(n7414), .D(n7413), .Z(n7417) );
  CAOR2X2 U7729 ( .A(\s07.dataOut [8]), .B(n7559), .C(\s10.dataOut [8]), .D(
        n7493), .Z(n7416) );
  CANR3XL U7730 ( .A(\s01.dataOut [8]), .B(n7507), .C(n7417), .D(n7416), .Z(
        n7418) );
  CND4X1 U7731 ( .A(n7421), .B(n7420), .C(n7419), .D(n7418), .Z(n7422) );
  CMX2X1 U7732 ( .A0(\m03.DinMast [8]), .A1(n7422), .S(n7512), .Z(n4234) );
  CANR2X1 U7733 ( .A(\s11.dataOut [9]), .B(n7494), .C(\s09.dataOut [9]), .D(
        n7504), .Z(n7431) );
  CANR2XL U7734 ( .A(\s06.dataOut [9]), .B(n7533), .C(\s08.dataOut [9]), .D(
        n7496), .Z(n7430) );
  CANR2X1 U7735 ( .A(n7495), .B(\s00.dataOut [9]), .C(\s05.dataOut [9]), .D(
        n7497), .Z(n7429) );
  CANR2XL U7736 ( .A(\s02.dataOut [9]), .B(n7498), .C(\s13.dataOut [9]), .D(
        n7499), .Z(n7424) );
  CANR2XL U7737 ( .A(n7500), .B(\s03.dataOut [9]), .C(\s12.dataOut [9]), .D(
        n7517), .Z(n7423) );
  COND3X1 U7738 ( .A(n7425), .B(n7574), .C(n7424), .D(n7423), .Z(n7427) );
  CAOR2X2 U7739 ( .A(\s07.dataOut [9]), .B(n7559), .C(\s10.dataOut [9]), .D(
        n7493), .Z(n7426) );
  CANR3XL U7740 ( .A(\s01.dataOut [9]), .B(n7507), .C(n7427), .D(n7426), .Z(
        n7428) );
  CND4X1 U7741 ( .A(n7431), .B(n7430), .C(n7429), .D(n7428), .Z(n7432) );
  CMX2X1 U7742 ( .A0(\m03.DinMast [9]), .A1(n7432), .S(n7512), .Z(n4235) );
  CANR2X1 U7743 ( .A(\s10.dataOut [15]), .B(n7493), .C(\s09.dataOut [15]), .D(
        n7504), .Z(n7444) );
  CANR2X1 U7744 ( .A(\s05.dataOut [15]), .B(n7497), .C(\s13.dataOut [15]), .D(
        n7499), .Z(n7443) );
  CANR2X1 U7745 ( .A(n7495), .B(\s00.dataOut [15]), .C(\s06.dataOut [15]), .D(
        n7533), .Z(n7442) );
  CIVX2 U7746 ( .A(\s04.dataOut [15]), .Z(n7435) );
  CANR2XL U7747 ( .A(\s02.dataOut [15]), .B(n7498), .C(\s08.dataOut [15]), .D(
        n7496), .Z(n7434) );
  CANR2XL U7748 ( .A(n7500), .B(\s03.dataOut [15]), .C(\s12.dataOut [15]), .D(
        n7517), .Z(n7433) );
  COND3X1 U7749 ( .A(n7435), .B(n7574), .C(n7434), .D(n7433), .Z(n7440) );
  COND2X1 U7750 ( .A(n7438), .B(n7484), .C(n7437), .D(n7436), .Z(n7439) );
  CANR3XL U7751 ( .A(\s01.dataOut [15]), .B(n7507), .C(n7440), .D(n7439), .Z(
        n7441) );
  CND4X1 U7752 ( .A(n7444), .B(n7443), .C(n7442), .D(n7441), .Z(n7445) );
  CMX2X1 U7753 ( .A0(\m03.DinMast [15]), .A1(n7445), .S(n7512), .Z(n4241) );
  CANR2XL U7754 ( .A(\s09.dataOut [10]), .B(n7504), .C(\s10.dataOut [10]), .D(
        n7493), .Z(n7454) );
  CANR2XL U7755 ( .A(n7495), .B(\s00.dataOut [10]), .C(\s08.dataOut [10]), .D(
        n7496), .Z(n7453) );
  CANR2X1 U7756 ( .A(\s05.dataOut [10]), .B(n7497), .C(\s06.dataOut [10]), .D(
        n7533), .Z(n7452) );
  CANR2XL U7757 ( .A(\s02.dataOut [10]), .B(n7498), .C(\s13.dataOut [10]), .D(
        n7499), .Z(n7447) );
  CANR2XL U7758 ( .A(n7500), .B(\s03.dataOut [10]), .C(\s12.dataOut [10]), .D(
        n7517), .Z(n7446) );
  COND3X1 U7759 ( .A(n7448), .B(n7574), .C(n7447), .D(n7446), .Z(n7450) );
  CAOR2X2 U7760 ( .A(\s07.dataOut [10]), .B(n7559), .C(\s11.dataOut [10]), .D(
        n7494), .Z(n7449) );
  CANR3XL U7761 ( .A(\s01.dataOut [10]), .B(n7507), .C(n7450), .D(n7449), .Z(
        n7451) );
  CND4X1 U7762 ( .A(n7454), .B(n7453), .C(n7452), .D(n7451), .Z(n7455) );
  CMX2X1 U7763 ( .A0(\m03.DinMast [10]), .A1(n7455), .S(n7512), .Z(n4236) );
  CANR2X1 U7764 ( .A(\s11.dataOut [14]), .B(n7494), .C(\s01.dataOut [14]), .D(
        n7507), .Z(n7465) );
  CANR2XL U7765 ( .A(\s06.dataOut [14]), .B(n7533), .C(\s13.dataOut [14]), .D(
        n7499), .Z(n7464) );
  CANR2XL U7766 ( .A(n7500), .B(\s03.dataOut [14]), .C(\s04.dataOut [14]), .D(
        n7467), .Z(n7463) );
  CIVX2 U7767 ( .A(\s05.dataOut [14]), .Z(n7459) );
  CANR2XL U7768 ( .A(\s02.dataOut [14]), .B(n7498), .C(\s08.dataOut [14]), .D(
        n7496), .Z(n7457) );
  CANR2X1 U7769 ( .A(n7495), .B(\s00.dataOut [14]), .C(\s12.dataOut [14]), .D(
        n7517), .Z(n7456) );
  COND3X1 U7770 ( .A(n7459), .B(n7458), .C(n7457), .D(n7456), .Z(n7461) );
  CAOR2X2 U7771 ( .A(\s07.dataOut [14]), .B(n7559), .C(\s10.dataOut [14]), .D(
        n7493), .Z(n7460) );
  CANR3X1 U7772 ( .A(\s09.dataOut [14]), .B(n7504), .C(n7461), .D(n7460), .Z(
        n7462) );
  CND4X1 U7773 ( .A(n7465), .B(n7464), .C(n7463), .D(n7462), .Z(n7466) );
  CMX2X1 U7774 ( .A0(\m03.DinMast [14]), .A1(n7466), .S(n7512), .Z(n4240) );
  CANR2X1 U7775 ( .A(\s11.dataOut [11]), .B(n7494), .C(\s10.dataOut [11]), .D(
        n7493), .Z(n7477) );
  CANR2XL U7776 ( .A(n7500), .B(\s03.dataOut [11]), .C(\s08.dataOut [11]), .D(
        n7496), .Z(n7476) );
  CANR2X1 U7777 ( .A(\s05.dataOut [11]), .B(n7497), .C(\s12.dataOut [11]), .D(
        n7517), .Z(n7475) );
  CIVX2 U7778 ( .A(\s00.dataOut [11]), .Z(n7470) );
  CANR2XL U7779 ( .A(\s13.dataOut [11]), .B(n7499), .C(\s02.dataOut [11]), .D(
        n7498), .Z(n7469) );
  CANR2X1 U7780 ( .A(\s06.dataOut [11]), .B(n7533), .C(\s04.dataOut [11]), .D(
        n7467), .Z(n7468) );
  COND3X1 U7781 ( .A(n7471), .B(n7470), .C(n7469), .D(n7468), .Z(n7473) );
  CAOR2X2 U7782 ( .A(\s07.dataOut [11]), .B(n7559), .C(\s09.dataOut [11]), .D(
        n7504), .Z(n7472) );
  CANR3XL U7783 ( .A(\s01.dataOut [11]), .B(n7507), .C(n7473), .D(n7472), .Z(
        n7474) );
  CND4X1 U7784 ( .A(n7477), .B(n7476), .C(n7475), .D(n7474), .Z(n7478) );
  CMX2X1 U7785 ( .A0(\m03.DinMast [11]), .A1(n7478), .S(n7512), .Z(n4237) );
  CANR2X1 U7786 ( .A(\s11.dataOut [13]), .B(n7494), .C(\s01.dataOut [13]), .D(
        n7507), .Z(n7491) );
  CANR2XL U7787 ( .A(n7495), .B(\s00.dataOut [13]), .C(n7500), .D(
        \s03.dataOut [13]), .Z(n7490) );
  CANR2XL U7788 ( .A(\s12.dataOut [13]), .B(n7517), .C(\s13.dataOut [13]), .D(
        n7499), .Z(n7489) );
  CIVX2 U7789 ( .A(\s04.dataOut [13]), .Z(n7481) );
  CANR2XL U7790 ( .A(\s02.dataOut [13]), .B(n7498), .C(\s08.dataOut [13]), .D(
        n7496), .Z(n7480) );
  CANR2X1 U7791 ( .A(\s05.dataOut [13]), .B(n7497), .C(\s06.dataOut [13]), .D(
        n7533), .Z(n7479) );
  COND3X1 U7792 ( .A(n7481), .B(n7574), .C(n7480), .D(n7479), .Z(n7487) );
  COND2X1 U7793 ( .A(n7485), .B(n7484), .C(n7483), .D(n7482), .Z(n7486) );
  CANR3X1 U7794 ( .A(\s09.dataOut [13]), .B(n7504), .C(n7487), .D(n7486), .Z(
        n7488) );
  CND4X1 U7795 ( .A(n7491), .B(n7490), .C(n7489), .D(n7488), .Z(n7492) );
  CMX2X1 U7796 ( .A0(\m03.DinMast [13]), .A1(n7492), .S(n7512), .Z(n4239) );
  CANR2X1 U7797 ( .A(\s11.dataOut [12]), .B(n7494), .C(\s10.dataOut [12]), .D(
        n7493), .Z(n7511) );
  CANR2X1 U7798 ( .A(n7495), .B(\s00.dataOut [12]), .C(\s12.dataOut [12]), .D(
        n7517), .Z(n7510) );
  CANR2XL U7799 ( .A(\s05.dataOut [12]), .B(n7497), .C(\s08.dataOut [12]), .D(
        n7496), .Z(n7509) );
  CANR2XL U7800 ( .A(\s13.dataOut [12]), .B(n7499), .C(\s02.dataOut [12]), .D(
        n7498), .Z(n7502) );
  CANR2XL U7801 ( .A(n7500), .B(\s03.dataOut [12]), .C(\s06.dataOut [12]), .D(
        n7533), .Z(n7501) );
  COND3X1 U7802 ( .A(n7503), .B(n7574), .C(n7502), .D(n7501), .Z(n7506) );
  CAOR2X2 U7803 ( .A(\s07.dataOut [12]), .B(n7559), .C(\s09.dataOut [12]), .D(
        n7504), .Z(n7505) );
  CANR3XL U7804 ( .A(\s01.dataOut [12]), .B(n7507), .C(n7506), .D(n7505), .Z(
        n7508) );
  CND4X1 U7805 ( .A(n7511), .B(n7510), .C(n7509), .D(n7508), .Z(n7513) );
  CMX2X1 U7806 ( .A0(\m03.DinMast [12]), .A1(n7513), .S(n7512), .Z(n4238) );
  CMX2X1 U7807 ( .A0(n7628), .A1(\s11.dbus_in [11]), .S(n7594), .Z(n4333) );
  CMX2X1 U7808 ( .A0(n7632), .A1(\s11.dbus_in [1]), .S(n7594), .Z(n4323) );
  CMX2X1 U7809 ( .A0(n7629), .A1(\s11.dbus_in [7]), .S(n7594), .Z(n4329) );
  CMX2X1 U7810 ( .A0(n7631), .A1(\s11.dbus_in [3]), .S(n7594), .Z(n4325) );
  CMX2X1 U7811 ( .A0(n7626), .A1(\s11.dbus_in [10]), .S(n7594), .Z(n4332) );
  CMX2X1 U7812 ( .A0(n7630), .A1(\s11.dbus_in [5]), .S(n7594), .Z(n4327) );
  COND2X1 U7813 ( .A(n7589), .B(n7515), .C(n7577), .D(n7514), .Z(n7524) );
  CANR2X1 U7814 ( .A(n7560), .B(n7517), .C(n7579), .D(n7516), .Z(n7521) );
  CANR2XL U7815 ( .A(n7585), .B(n7519), .C(n7583), .D(n7518), .Z(n7520) );
  COND3X1 U7816 ( .A(n7549), .B(n7522), .C(n7521), .D(n7520), .Z(n7523) );
  CNR2X1 U7817 ( .A(n7524), .B(n7523), .Z(n7622) );
  CMX2X1 U7818 ( .A0(n7636), .A1(\s12.dbus_in [14]), .S(n7622), .Z(n5184) );
  CNIVX1 U7819 ( .A(n7525), .Z(n7710) );
  CMX2X1 U7820 ( .A0(n7621), .A1(\s05.Adr [2]), .S(n7710), .Z(n4724) );
  CANR2XL U7821 ( .A(\m00.YouGotIt ), .B(\m00.addrM [4]), .C(\m01.addrM [4]), 
        .D(n7642), .Z(n7529) );
  CANR2X1 U7822 ( .A(\m03.addrM [4]), .B(n7644), .C(\m02.addrM [4]), .D(n7643), 
        .Z(n7528) );
  CANR2X1 U7823 ( .A(\m05.addrM [4]), .B(n7641), .C(n7640), .D(\m06.addrM [4]), 
        .Z(n7527) );
  CND2X1 U7824 ( .A(\m04.addrM [4]), .B(n7648), .Z(n7526) );
  CND4X1 U7825 ( .A(n7529), .B(n7528), .C(n7527), .D(n7526), .Z(n7634) );
  CIVX2 U7826 ( .A(n7659), .Z(n7530) );
  COND2X1 U7827 ( .A(n7589), .B(n7531), .C(n7577), .D(n7530), .Z(n7541) );
  CANR2X1 U7828 ( .A(n7560), .B(n7533), .C(n7581), .D(n7532), .Z(n7537) );
  CANR2X1 U7829 ( .A(n7585), .B(n7535), .C(n7583), .D(n7534), .Z(n7536) );
  COND3X1 U7830 ( .A(n7539), .B(n7538), .C(n7537), .D(n7536), .Z(n7540) );
  CNR2X1 U7831 ( .A(n7541), .B(n7540), .Z(n7623) );
  CMX2X1 U7832 ( .A0(n7634), .A1(\s06.Adr [4]), .S(n7623), .Z(n4662) );
  CMX2X1 U7833 ( .A0(n7621), .A1(\s06.Adr [2]), .S(n7623), .Z(n4660) );
  CMX2X1 U7834 ( .A0(n7687), .A1(\s06.Adr [1]), .S(n7623), .Z(n4659) );
  CMX2X1 U7835 ( .A0(n7625), .A1(\s06.Adr [0]), .S(n7623), .Z(n4658) );
  CMX2X1 U7836 ( .A0(n7627), .A1(\s06.dbus_in [13]), .S(n7623), .Z(n4655) );
  CMX2X1 U7837 ( .A0(n7628), .A1(\s06.dbus_in [11]), .S(n7623), .Z(n4653) );
  CMX2X1 U7838 ( .A0(n7626), .A1(\s06.dbus_in [10]), .S(n7623), .Z(n4652) );
  CMX2X1 U7839 ( .A0(n7629), .A1(\s06.dbus_in [7]), .S(n7623), .Z(n4649) );
  CMX2X1 U7840 ( .A0(n7630), .A1(\s06.dbus_in [5]), .S(n7623), .Z(n4647) );
  CMX2X1 U7841 ( .A0(n7631), .A1(\s06.dbus_in [3]), .S(n7623), .Z(n4645) );
  CMX2X1 U7842 ( .A0(n7684), .A1(\s06.dbus_in [0]), .S(n7623), .Z(n4642) );
  CAOR2XL U7843 ( .A(\m00.YouGotIt ), .B(\m00.addrM [7]), .C(\m01.addrM [7]), 
        .D(n7642), .Z(n7545) );
  COND2X1 U7844 ( .A(n7543), .B(n7566), .C(n7542), .D(n7564), .Z(n7544) );
  CANR3X1 U7845 ( .A(n7640), .B(\m06.addrM [7]), .C(n7545), .D(n7544), .Z(
        n7547) );
  CANR2X1 U7846 ( .A(\m05.addrM [7]), .B(n7641), .C(\m04.addrM [7]), .D(n7648), 
        .Z(n7546) );
  CND2X1 U7847 ( .A(n7547), .B(n7546), .Z(n7624) );
  COND2X1 U7848 ( .A(n7577), .B(n7550), .C(n7549), .D(n7548), .Z(n7551) );
  CANR1XL U7849 ( .A(n7583), .B(n7552), .C(n7551), .Z(n7556) );
  CANR2XL U7850 ( .A(n7579), .B(n7554), .C(n7585), .D(n7553), .Z(n7555) );
  COND3X1 U7851 ( .A(n7589), .B(n7557), .C(n7556), .D(n7555), .Z(n7558) );
  CANR1XL U7852 ( .A(n7560), .B(n7559), .C(n7558), .Z(n7572) );
  CNIVX1 U7853 ( .A(n7572), .Z(n7714) );
  CMX2X1 U7854 ( .A0(n7624), .A1(\s07.Adr [7]), .S(n7714), .Z(n4601) );
  COND2X1 U7855 ( .A(n7690), .B(n7563), .C(n7562), .D(n7561), .Z(n7569) );
  COND2X1 U7856 ( .A(n7567), .B(n7566), .C(n7565), .D(n7564), .Z(n7568) );
  CANR3X1 U7857 ( .A(n7640), .B(\m06.addrM [6]), .C(n7569), .D(n7568), .Z(
        n7571) );
  CANR2X1 U7858 ( .A(\m05.addrM [6]), .B(n7641), .C(\m04.addrM [6]), .D(n7648), 
        .Z(n7570) );
  CND2X1 U7859 ( .A(n7571), .B(n7570), .Z(n7609) );
  CMX2X1 U7860 ( .A0(n7609), .A1(\s07.Adr [6]), .S(n7714), .Z(n4600) );
  CMX2X1 U7861 ( .A0(n7621), .A1(\s07.Adr [2]), .S(n7572), .Z(n4596) );
  CMX2X1 U7862 ( .A0(n7629), .A1(\s07.dbus_in [7]), .S(n7572), .Z(n4585) );
  CMX2X1 U7863 ( .A0(n7630), .A1(\s07.dbus_in [5]), .S(n7572), .Z(n4583) );
  CMX2X1 U7864 ( .A0(n7631), .A1(\s07.dbus_in [3]), .S(n7572), .Z(n4581) );
  CNIVX1 U7865 ( .A(n7573), .Z(n7716) );
  CMX2X1 U7866 ( .A0(n7624), .A1(\s08.Adr [7]), .S(n7716), .Z(n4537) );
  CMX2X1 U7867 ( .A0(n7609), .A1(\s08.Adr [6]), .S(n7716), .Z(n4536) );
  COND2X1 U7868 ( .A(n7577), .B(n7576), .C(n7575), .D(n7574), .Z(n7591) );
  CANR2X1 U7869 ( .A(n7581), .B(n7580), .C(n7579), .D(n7578), .Z(n7587) );
  CANR2X1 U7870 ( .A(n7585), .B(n7584), .C(n7583), .D(n7582), .Z(n7586) );
  COND3X1 U7871 ( .A(n7589), .B(n7588), .C(n7587), .D(n7586), .Z(n7590) );
  CNR2X1 U7872 ( .A(n7591), .B(n7590), .Z(n7608) );
  CMX2X1 U7873 ( .A0(n7632), .A1(\s04.dbus_in [1]), .S(n7608), .Z(n4771) );
  CNIVX1 U7874 ( .A(n7592), .Z(n7718) );
  CMX2X1 U7875 ( .A0(n7609), .A1(\s09.Adr [6]), .S(n7718), .Z(n4472) );
  CMX2X1 U7876 ( .A0(n7682), .A1(\s09.dbus_in [9]), .S(n7718), .Z(n4459) );
  CMX2X1 U7877 ( .A0(n7683), .A1(\s09.dbus_in [2]), .S(n7718), .Z(n4452) );
  CNIVX1 U7878 ( .A(n7593), .Z(n7720) );
  CMX2X1 U7879 ( .A0(n7609), .A1(\s10.Adr [6]), .S(n7720), .Z(n4408) );
  CNIVX1 U7880 ( .A(n7594), .Z(n7722) );
  CMX2X1 U7881 ( .A0(n7624), .A1(\s11.Adr [7]), .S(n7722), .Z(n4345) );
  CMX2X1 U7882 ( .A0(n7609), .A1(\s11.Adr [6]), .S(n7722), .Z(n4344) );
  CMX2X1 U7883 ( .A0(n7637), .A1(\s12.dbus_in [12]), .S(n7622), .Z(n5182) );
  CMX2X1 U7884 ( .A0(n7626), .A1(\s12.dbus_in [10]), .S(n7622), .Z(n5180) );
  CMX2X1 U7885 ( .A0(n7685), .A1(\s12.dbus_in [8]), .S(n7622), .Z(n5178) );
  CMX2X1 U7886 ( .A0(n7686), .A1(\s12.dbus_in [6]), .S(n7622), .Z(n5176) );
  CMX2X1 U7887 ( .A0(n7631), .A1(\s12.dbus_in [3]), .S(n7622), .Z(n5173) );
  CMX2X1 U7888 ( .A0(n7632), .A1(\s12.dbus_in [1]), .S(n7622), .Z(n5171) );
  CNIVX1 U7889 ( .A(n7595), .Z(n7700) );
  CMX2X1 U7890 ( .A0(n7624), .A1(\s13.Adr [7]), .S(n7700), .Z(n5129) );
  CMX2X1 U7891 ( .A0(n7609), .A1(\s13.Adr [6]), .S(n7700), .Z(n5128) );
  CNIVX1 U7892 ( .A(n7596), .Z(n7702) );
  CMX2X1 U7893 ( .A0(n7624), .A1(\s00.Adr [7]), .S(n7702), .Z(n5065) );
  CMX2X1 U7894 ( .A0(n7609), .A1(\s00.Adr [6]), .S(n7702), .Z(n5064) );
  CNIVX1 U7895 ( .A(n7597), .Z(n7704) );
  CMX2X1 U7896 ( .A0(n7609), .A1(\s01.Adr [6]), .S(n7704), .Z(n4984) );
  CMX2X1 U7897 ( .A0(n7621), .A1(\s01.Adr [2]), .S(n7704), .Z(n4980) );
  CMX2X1 U7898 ( .A0(n7682), .A1(\s01.dbus_in [9]), .S(n7704), .Z(n4971) );
  CMX2X1 U7899 ( .A0(n7683), .A1(\s01.dbus_in [2]), .S(n7704), .Z(n4964) );
  CNIVX1 U7900 ( .A(n7598), .Z(n7638) );
  CMX2X1 U7901 ( .A0(n7621), .A1(\s02.Adr [2]), .S(n7638), .Z(n4916) );
  CNIVX1 U7902 ( .A(n7599), .Z(n7706) );
  CMX2X1 U7903 ( .A0(n7624), .A1(\s03.Adr [7]), .S(n7706), .Z(n4857) );
  CMX2X1 U7904 ( .A0(n7609), .A1(\s03.Adr [6]), .S(n7706), .Z(n4856) );
  CNIVX1 U7905 ( .A(n7608), .Z(n7708) );
  CMX2X1 U7906 ( .A0(n7609), .A1(\s04.Adr [6]), .S(n7708), .Z(n4792) );
  CANR2XL U7907 ( .A(\m00.YouGotIt ), .B(\m00.addrM [5]), .C(\m01.addrM [5]), 
        .D(n7642), .Z(n7603) );
  CANR2X1 U7908 ( .A(\m03.addrM [5]), .B(n7644), .C(\m02.addrM [5]), .D(n7643), 
        .Z(n7602) );
  CANR2X1 U7909 ( .A(\m05.addrM [5]), .B(n7641), .C(n7640), .D(\m06.addrM [5]), 
        .Z(n7601) );
  CND2X1 U7910 ( .A(\m04.addrM [5]), .B(n7648), .Z(n7600) );
  CND4X1 U7911 ( .A(n7603), .B(n7602), .C(n7601), .D(n7600), .Z(n7654) );
  CMX2X1 U7912 ( .A0(n7654), .A1(\s04.Adr [5]), .S(n7608), .Z(n4791) );
  CANR2XL U7913 ( .A(\m00.YouGotIt ), .B(\m00.addrM [3]), .C(\m01.addrM [3]), 
        .D(n7642), .Z(n7607) );
  CANR2X1 U7914 ( .A(\m03.addrM [3]), .B(n7644), .C(\m02.addrM [3]), .D(n7643), 
        .Z(n7606) );
  CANR2X1 U7915 ( .A(\m05.addrM [3]), .B(n7641), .C(n7640), .D(\m06.addrM [3]), 
        .Z(n7605) );
  CND2X1 U7916 ( .A(\m04.addrM [3]), .B(n7648), .Z(n7604) );
  CND4X1 U7917 ( .A(n7607), .B(n7606), .C(n7605), .D(n7604), .Z(n7655) );
  CMX2X1 U7918 ( .A0(n7655), .A1(\s04.Adr [3]), .S(n7608), .Z(n4789) );
  CMX2X1 U7919 ( .A0(n7621), .A1(\s04.Adr [2]), .S(n7708), .Z(n4788) );
  CMX2X1 U7920 ( .A0(n7687), .A1(\s04.Adr [1]), .S(n7608), .Z(n4787) );
  CMX2X1 U7921 ( .A0(n7625), .A1(\s04.Adr [0]), .S(n7608), .Z(n4786) );
  CMX2X1 U7922 ( .A0(n7627), .A1(\s04.dbus_in [13]), .S(n7608), .Z(n4783) );
  CMX2X1 U7923 ( .A0(n7628), .A1(\s04.dbus_in [11]), .S(n7608), .Z(n4781) );
  CMX2X1 U7924 ( .A0(n7626), .A1(\s04.dbus_in [10]), .S(n7608), .Z(n4780) );
  CMX2X1 U7925 ( .A0(n7629), .A1(\s04.dbus_in [7]), .S(n7608), .Z(n4777) );
  CMX2X1 U7926 ( .A0(n7630), .A1(\s04.dbus_in [5]), .S(n7608), .Z(n4775) );
  CMX2X1 U7927 ( .A0(n7631), .A1(\s04.dbus_in [3]), .S(n7608), .Z(n4773) );
  CMX2X1 U7928 ( .A0(n7609), .A1(\s12.Adr [6]), .S(n7622), .Z(n4280) );
  CANR2XL U7929 ( .A(\m00.YouGotIt ), .B(\m00.addrM [8]), .C(\m01.addrM [8]), 
        .D(n7642), .Z(n7611) );
  CANR2X1 U7930 ( .A(\m03.addrM [8]), .B(n7644), .C(\m02.addrM [8]), .D(n7643), 
        .Z(n7610) );
  COND3X1 U7931 ( .A(n7613), .B(n7612), .C(n7611), .D(n7610), .Z(n7614) );
  CANR1XL U7932 ( .A(\m05.addrM [8]), .B(n7641), .C(n7614), .Z(n7615) );
  COND1XL U7933 ( .A(n7617), .B(n7616), .C(n7615), .Z(n7633) );
  CMX2X1 U7934 ( .A0(n7633), .A1(\s12.Adr [8]), .S(n7622), .Z(n4282) );
  CMX2X1 U7935 ( .A0(n7625), .A1(\s12.Adr [0]), .S(n7622), .Z(n4274) );
  CNIVX1 U7936 ( .A(n7622), .Z(n7724) );
  CMX2X1 U7937 ( .A0(n7624), .A1(\s12.Adr [7]), .S(n7724), .Z(n4281) );
  CIVXL U7938 ( .A(\m06.YouGotIt ), .Z(n7620) );
  CND2X1 U7939 ( .A(n7618), .B(n7620), .Z(n7689) );
  CNR2X1 U7940 ( .A(\m00.need ), .B(n7689), .Z(n7695) );
  CND2IX1 U7941 ( .B(\m04.need ), .A(n7695), .Z(n7693) );
  CNR2X1 U7942 ( .A(\m05.need ), .B(n7693), .Z(n7691) );
  CNR2IX1 U7943 ( .B(n7691), .A(\m03.need ), .Z(n7652) );
  CNR2IX1 U7944 ( .B(n7652), .A(\m01.need ), .Z(n7697) );
  CND2X1 U7945 ( .A(n7697), .B(\m06.need ), .Z(n7619) );
  COND2XL U7946 ( .A(\clock.rst ), .B(n7620), .C(\m02.need ), .D(n7619), .Z(
        n5285) );
  CMX2X1 U7947 ( .A0(n7621), .A1(\s12.Adr [2]), .S(n7622), .Z(n4276) );
  CMX2X1 U7948 ( .A0(n7634), .A1(\s12.Adr [4]), .S(n7622), .Z(n4278) );
  CNIVXL U7949 ( .A(\clock.sysClk ), .Z(n7737) );
  CNIVXL U7950 ( .A(\clock.sysClk ), .Z(n7745) );
  CNIVXL U7951 ( .A(\clock.sysClk ), .Z(n7744) );
  CNIVXL U7952 ( .A(\clock.sysClk ), .Z(n7743) );
  CNIVXL U7953 ( .A(\clock.sysClk ), .Z(n7742) );
  CNIVXL U7954 ( .A(\clock.sysClk ), .Z(n7735) );
  CNIVXL U7955 ( .A(\clock.sysClk ), .Z(n7726) );
  CNIVXL U7956 ( .A(\clock.sysClk ), .Z(n7730) );
  CNIVXL U7957 ( .A(\clock.sysClk ), .Z(n7729) );
  CNIVXL U7958 ( .A(\clock.sysClk ), .Z(n7728) );
  CNIVXL U7959 ( .A(\clock.sysClk ), .Z(n7727) );
  CNIVXL U7960 ( .A(\clock.sysClk ), .Z(n7734) );
  CNIVXL U7961 ( .A(\clock.sysClk ), .Z(n7732) );
  CNIVXL U7962 ( .A(\clock.sysClk ), .Z(n7731) );
  CNIVXL U7963 ( .A(\clock.sysClk ), .Z(n7736) );
  CMX2X1 U7964 ( .A0(n7684), .A1(\s04.dbus_in [0]), .S(n7708), .Z(n4770) );
  CMX2X1 U7965 ( .A0(n7634), .A1(\s05.Adr [4]), .S(n7710), .Z(n4726) );
  CMX2X1 U7966 ( .A0(n7655), .A1(\s05.Adr [3]), .S(n7710), .Z(n4725) );
  CMX2X1 U7967 ( .A0(n7625), .A1(\s05.Adr [0]), .S(n7710), .Z(n4722) );
  CMX2X1 U7968 ( .A0(n7627), .A1(\s05.dbus_in [13]), .S(n7710), .Z(n4719) );
  CMX2X1 U7969 ( .A0(n7637), .A1(\s05.dbus_in [12]), .S(n7710), .Z(n4718) );
  CMX2X1 U7970 ( .A0(n7626), .A1(\s05.dbus_in [10]), .S(n7710), .Z(n4716) );
  CMX2X1 U7971 ( .A0(n7682), .A1(\s05.dbus_in [9]), .S(n7710), .Z(n4715) );
  CMX2X1 U7972 ( .A0(n7685), .A1(\s05.dbus_in [8]), .S(n7710), .Z(n4714) );
  CMX2X1 U7973 ( .A0(n7686), .A1(\s05.dbus_in [6]), .S(n7710), .Z(n4712) );
  CMX2X1 U7974 ( .A0(n7631), .A1(\s05.dbus_in [3]), .S(n7710), .Z(n4709) );
  CMX2X1 U7975 ( .A0(n7632), .A1(\s05.dbus_in [1]), .S(n7710), .Z(n4707) );
  CNIVX1 U7976 ( .A(n7623), .Z(n7712) );
  CMX2X1 U7977 ( .A0(n7654), .A1(\s06.Adr [5]), .S(n7712), .Z(n4663) );
  CMX2X1 U7978 ( .A0(n7655), .A1(\s06.Adr [3]), .S(n7712), .Z(n4661) );
  CMX2X1 U7979 ( .A0(n7635), .A1(\s06.dbus_in [15]), .S(n7712), .Z(n4657) );
  CMX2X1 U7980 ( .A0(n7636), .A1(\s06.dbus_in [14]), .S(n7712), .Z(n4656) );
  CMX2X1 U7981 ( .A0(n7637), .A1(\s06.dbus_in [12]), .S(n7712), .Z(n4654) );
  CMX2X1 U7982 ( .A0(n7682), .A1(\s06.dbus_in [9]), .S(n7712), .Z(n4651) );
  CMX2X1 U7983 ( .A0(n7685), .A1(\s06.dbus_in [8]), .S(n7712), .Z(n4650) );
  CMX2X1 U7984 ( .A0(n7686), .A1(\s06.dbus_in [6]), .S(n7712), .Z(n4648) );
  CMX2X1 U7985 ( .A0(n7653), .A1(\s06.dbus_in [4]), .S(n7712), .Z(n4646) );
  CMX2X1 U7986 ( .A0(n7683), .A1(\s06.dbus_in [2]), .S(n7712), .Z(n4644) );
  CMX2X1 U7987 ( .A0(n7632), .A1(\s06.dbus_in [1]), .S(n7712), .Z(n4643) );
  CMX2X1 U7988 ( .A0(n7633), .A1(\s07.Adr [8]), .S(n7714), .Z(n4602) );
  CMX2X1 U7989 ( .A0(n7654), .A1(\s07.Adr [5]), .S(n7714), .Z(n4599) );
  CMX2X1 U7990 ( .A0(n7634), .A1(\s07.Adr [4]), .S(n7714), .Z(n4598) );
  CMX2X1 U7991 ( .A0(n7655), .A1(\s07.Adr [3]), .S(n7714), .Z(n4597) );
  CMX2X1 U7992 ( .A0(n7687), .A1(\s07.Adr [1]), .S(n7714), .Z(n4595) );
  CMX2X1 U7993 ( .A0(n7625), .A1(\s07.Adr [0]), .S(n7714), .Z(n4594) );
  CMX2X1 U7994 ( .A0(n7635), .A1(\s07.dbus_in [15]), .S(n7714), .Z(n4593) );
  CMX2X1 U7995 ( .A0(n7636), .A1(\s07.dbus_in [14]), .S(n7714), .Z(n4592) );
  CMX2X1 U7996 ( .A0(n7627), .A1(\s07.dbus_in [13]), .S(n7714), .Z(n4591) );
  CMX2X1 U7997 ( .A0(n7637), .A1(\s07.dbus_in [12]), .S(n7714), .Z(n4590) );
  CMX2X1 U7998 ( .A0(n7628), .A1(\s07.dbus_in [11]), .S(n7714), .Z(n4589) );
  CMX2X1 U7999 ( .A0(n7626), .A1(\s07.dbus_in [10]), .S(n7714), .Z(n4588) );
  CMX2X1 U8000 ( .A0(n7682), .A1(\s07.dbus_in [9]), .S(n7714), .Z(n4587) );
  CMX2X1 U8001 ( .A0(n7685), .A1(\s07.dbus_in [8]), .S(n7714), .Z(n4586) );
  CMX2X1 U8002 ( .A0(n7686), .A1(\s07.dbus_in [6]), .S(n7714), .Z(n4584) );
  CMX2X1 U8003 ( .A0(n7653), .A1(\s07.dbus_in [4]), .S(n7714), .Z(n4582) );
  CMX2X1 U8004 ( .A0(n7683), .A1(\s07.dbus_in [2]), .S(n7714), .Z(n4580) );
  CMX2X1 U8005 ( .A0(n7632), .A1(\s07.dbus_in [1]), .S(n7714), .Z(n4579) );
  CMX2X1 U8006 ( .A0(n7684), .A1(\s07.dbus_in [0]), .S(n7714), .Z(n4578) );
  CMX2X1 U8007 ( .A0(n7633), .A1(\s08.Adr [8]), .S(n7716), .Z(n4538) );
  CMX2X1 U8008 ( .A0(n7654), .A1(\s08.Adr [5]), .S(n7716), .Z(n4535) );
  CMX2X1 U8009 ( .A0(n7634), .A1(\s08.Adr [4]), .S(n7716), .Z(n4534) );
  CMX2X1 U8010 ( .A0(n7655), .A1(\s08.Adr [3]), .S(n7716), .Z(n4533) );
  CMX2X1 U8011 ( .A0(n7687), .A1(\s08.Adr [1]), .S(n7716), .Z(n4531) );
  CMX2X1 U8012 ( .A0(n7635), .A1(\s12.dbus_in [15]), .S(n7724), .Z(n5185) );
  CMX2X1 U8013 ( .A0(n7635), .A1(\s08.dbus_in [15]), .S(n7716), .Z(n4529) );
  CMX2X1 U8014 ( .A0(n7636), .A1(\s08.dbus_in [14]), .S(n7716), .Z(n4528) );
  CMX2X1 U8015 ( .A0(n7637), .A1(\s08.dbus_in [12]), .S(n7716), .Z(n4526) );
  CMX2X1 U8016 ( .A0(n7682), .A1(\s08.dbus_in [9]), .S(n7716), .Z(n4523) );
  CMX2X1 U8017 ( .A0(n7685), .A1(\s08.dbus_in [8]), .S(n7716), .Z(n4522) );
  CMX2X1 U8018 ( .A0(n7686), .A1(\s08.dbus_in [6]), .S(n7716), .Z(n4520) );
  CMX2X1 U8019 ( .A0(n7653), .A1(\s08.dbus_in [4]), .S(n7716), .Z(n4518) );
  CMX2X1 U8020 ( .A0(n7683), .A1(\s08.dbus_in [2]), .S(n7716), .Z(n4516) );
  CMX2X1 U8021 ( .A0(n7684), .A1(\s08.dbus_in [0]), .S(n7716), .Z(n4514) );
  CMX2X1 U8022 ( .A0(n7624), .A1(\s09.Adr [7]), .S(n7718), .Z(n4473) );
  CMX2X1 U8023 ( .A0(n7654), .A1(\s09.Adr [5]), .S(n7718), .Z(n4471) );
  CMX2X1 U8024 ( .A0(n7634), .A1(\s09.Adr [4]), .S(n7718), .Z(n4470) );
  CMX2X1 U8025 ( .A0(n7655), .A1(\s09.Adr [3]), .S(n7718), .Z(n4469) );
  CMX2X1 U8026 ( .A0(n7687), .A1(\s09.Adr [1]), .S(n7718), .Z(n4467) );
  CMX2X1 U8027 ( .A0(n7636), .A1(\s09.dbus_in [14]), .S(n7718), .Z(n4464) );
  CMX2X1 U8028 ( .A0(n7627), .A1(\s09.dbus_in [13]), .S(n7718), .Z(n4463) );
  CMX2X1 U8029 ( .A0(n7628), .A1(\s09.dbus_in [11]), .S(n7718), .Z(n4461) );
  CMX2X1 U8030 ( .A0(n7685), .A1(\s09.dbus_in [8]), .S(n7718), .Z(n4458) );
  CMX2X1 U8031 ( .A0(n7686), .A1(\s09.dbus_in [6]), .S(n7718), .Z(n4456) );
  CMX2X1 U8032 ( .A0(n7653), .A1(\s09.dbus_in [4]), .S(n7718), .Z(n4454) );
  CMX2X1 U8033 ( .A0(n7684), .A1(\s09.dbus_in [0]), .S(n7718), .Z(n4450) );
  CMX2X1 U8034 ( .A0(n7654), .A1(\s10.Adr [5]), .S(n7720), .Z(n4407) );
  CMX2X1 U8035 ( .A0(n7634), .A1(\s10.Adr [4]), .S(n7720), .Z(n4406) );
  CMX2X1 U8036 ( .A0(n7655), .A1(\s10.Adr [3]), .S(n7720), .Z(n4405) );
  CMX2X1 U8037 ( .A0(n7625), .A1(\s10.Adr [0]), .S(n7720), .Z(n4402) );
  CMX2X1 U8038 ( .A0(n7635), .A1(\s10.dbus_in [15]), .S(n7720), .Z(n4401) );
  CMX2X1 U8039 ( .A0(n7627), .A1(\s10.dbus_in [13]), .S(n7720), .Z(n4399) );
  CMX2X1 U8040 ( .A0(n7626), .A1(\s10.dbus_in [10]), .S(n7720), .Z(n4396) );
  CMX2X1 U8041 ( .A0(n7682), .A1(\s10.dbus_in [9]), .S(n7720), .Z(n4395) );
  CMX2X1 U8042 ( .A0(n7685), .A1(\s10.dbus_in [8]), .S(n7720), .Z(n4394) );
  CMX2X1 U8043 ( .A0(n7686), .A1(\s10.dbus_in [6]), .S(n7720), .Z(n4392) );
  CMX2X1 U8044 ( .A0(n7653), .A1(\s10.dbus_in [4]), .S(n7720), .Z(n4390) );
  CMX2X1 U8045 ( .A0(n7683), .A1(\s10.dbus_in [2]), .S(n7720), .Z(n4388) );
  CMX2X1 U8046 ( .A0(n7684), .A1(\s10.dbus_in [0]), .S(n7720), .Z(n4386) );
  CMX2X1 U8047 ( .A0(n7633), .A1(\s11.Adr [8]), .S(n7722), .Z(n4346) );
  CMX2X1 U8048 ( .A0(n7654), .A1(\s11.Adr [5]), .S(n7722), .Z(n4343) );
  CMX2X1 U8049 ( .A0(n7634), .A1(\s11.Adr [4]), .S(n7722), .Z(n4342) );
  CMX2X1 U8050 ( .A0(n7655), .A1(\s11.Adr [3]), .S(n7722), .Z(n4341) );
  CMX2X1 U8051 ( .A0(n7687), .A1(\s11.Adr [1]), .S(n7722), .Z(n4339) );
  CMX2X1 U8052 ( .A0(n7635), .A1(\s11.dbus_in [15]), .S(n7722), .Z(n4337) );
  CMX2X1 U8053 ( .A0(n7636), .A1(\s11.dbus_in [14]), .S(n7722), .Z(n4336) );
  CMX2X1 U8054 ( .A0(n7683), .A1(\s04.dbus_in [2]), .S(n7708), .Z(n4772) );
  CMX2X1 U8055 ( .A0(n7628), .A1(\s12.dbus_in [11]), .S(n7724), .Z(n5181) );
  CMX2X1 U8056 ( .A0(n7682), .A1(\s12.dbus_in [9]), .S(n7724), .Z(n5179) );
  CMX2X1 U8057 ( .A0(n7629), .A1(\s12.dbus_in [7]), .S(n7724), .Z(n5177) );
  CMX2X1 U8058 ( .A0(n7630), .A1(\s12.dbus_in [5]), .S(n7724), .Z(n5175) );
  CMX2X1 U8059 ( .A0(n7653), .A1(\s12.dbus_in [4]), .S(n7724), .Z(n5174) );
  CMX2X1 U8060 ( .A0(n7683), .A1(\s12.dbus_in [2]), .S(n7724), .Z(n5172) );
  CMX2X1 U8061 ( .A0(n7684), .A1(\s12.dbus_in [0]), .S(n7724), .Z(n5170) );
  CMX2X1 U8062 ( .A0(n7633), .A1(\s13.Adr [8]), .S(n7700), .Z(n5130) );
  CMX2X1 U8063 ( .A0(n7654), .A1(\s13.Adr [5]), .S(n7700), .Z(n5127) );
  CMX2X1 U8064 ( .A0(n7634), .A1(\s13.Adr [4]), .S(n7700), .Z(n5126) );
  CMX2X1 U8065 ( .A0(n7655), .A1(\s13.Adr [3]), .S(n7700), .Z(n5125) );
  CMX2X1 U8066 ( .A0(n7687), .A1(\s13.Adr [1]), .S(n7700), .Z(n5123) );
  CMX2X1 U8067 ( .A0(n7635), .A1(\s13.dbus_in [15]), .S(n7700), .Z(n5121) );
  CMX2X1 U8068 ( .A0(n7636), .A1(\s13.dbus_in [14]), .S(n7700), .Z(n5120) );
  CMX2X1 U8069 ( .A0(n7637), .A1(\s13.dbus_in [12]), .S(n7700), .Z(n5118) );
  CMX2X1 U8070 ( .A0(n7682), .A1(\s13.dbus_in [9]), .S(n7700), .Z(n5115) );
  CMX2X1 U8071 ( .A0(n7685), .A1(\s13.dbus_in [8]), .S(n7700), .Z(n5114) );
  CMX2X1 U8072 ( .A0(n7686), .A1(\s13.dbus_in [6]), .S(n7700), .Z(n5112) );
  CMX2X1 U8073 ( .A0(n7653), .A1(\s13.dbus_in [4]), .S(n7700), .Z(n5110) );
  CMX2X1 U8074 ( .A0(n7683), .A1(\s13.dbus_in [2]), .S(n7700), .Z(n5108) );
  CMX2X1 U8075 ( .A0(n7684), .A1(\s13.dbus_in [0]), .S(n7700), .Z(n5106) );
  CMX2X1 U8076 ( .A0(n7633), .A1(\s00.Adr [8]), .S(n7702), .Z(n5066) );
  CMX2X1 U8077 ( .A0(n7654), .A1(\s00.Adr [5]), .S(n7702), .Z(n5063) );
  CMX2X1 U8078 ( .A0(n7634), .A1(\s00.Adr [4]), .S(n7702), .Z(n5062) );
  CMX2X1 U8079 ( .A0(n7655), .A1(\s00.Adr [3]), .S(n7702), .Z(n5061) );
  CMX2X1 U8080 ( .A0(n7687), .A1(\s00.Adr [1]), .S(n7702), .Z(n5059) );
  CMX2X1 U8081 ( .A0(n7625), .A1(\s00.Adr [0]), .S(n7702), .Z(n5058) );
  CMX2X1 U8082 ( .A0(n7635), .A1(\s00.dbus_in [15]), .S(n7702), .Z(n5057) );
  CMX2X1 U8083 ( .A0(n7636), .A1(\s00.dbus_in [14]), .S(n7702), .Z(n5056) );
  CMX2X1 U8084 ( .A0(n7627), .A1(\s00.dbus_in [13]), .S(n7702), .Z(n5055) );
  CMX2X1 U8085 ( .A0(n7637), .A1(\s00.dbus_in [12]), .S(n7702), .Z(n5054) );
  CMX2X1 U8086 ( .A0(n7628), .A1(\s00.dbus_in [11]), .S(n7702), .Z(n5053) );
  CMX2X1 U8087 ( .A0(n7626), .A1(\s00.dbus_in [10]), .S(n7702), .Z(n5052) );
  CMX2X1 U8088 ( .A0(n7682), .A1(\s00.dbus_in [9]), .S(n7702), .Z(n5051) );
  CMX2X1 U8089 ( .A0(n7629), .A1(\s00.dbus_in [7]), .S(n7702), .Z(n5049) );
  CMX2X1 U8090 ( .A0(n7630), .A1(\s00.dbus_in [5]), .S(n7702), .Z(n5047) );
  CMX2X1 U8091 ( .A0(n7653), .A1(\s00.dbus_in [4]), .S(n7702), .Z(n5046) );
  CMX2X1 U8092 ( .A0(n7631), .A1(\s00.dbus_in [3]), .S(n7702), .Z(n5045) );
  CMX2X1 U8093 ( .A0(n7683), .A1(\s00.dbus_in [2]), .S(n7702), .Z(n5044) );
  CMX2X1 U8094 ( .A0(n7632), .A1(\s00.dbus_in [1]), .S(n7702), .Z(n5043) );
  CMX2X1 U8095 ( .A0(n7684), .A1(\s00.dbus_in [0]), .S(n7702), .Z(n5042) );
  CMX2X1 U8096 ( .A0(n7624), .A1(\s01.Adr [7]), .S(n7704), .Z(n4985) );
  CMX2X1 U8097 ( .A0(n7654), .A1(\s01.Adr [5]), .S(n7704), .Z(n4983) );
  CMX2X1 U8098 ( .A0(n7634), .A1(\s01.Adr [4]), .S(n7704), .Z(n4982) );
  CMX2X1 U8099 ( .A0(n7655), .A1(\s01.Adr [3]), .S(n7704), .Z(n4981) );
  CMX2X1 U8100 ( .A0(n7625), .A1(\s01.Adr [0]), .S(n7704), .Z(n4978) );
  CMX2X1 U8101 ( .A0(n7627), .A1(\s01.dbus_in [13]), .S(n7704), .Z(n4975) );
  CMX2X1 U8102 ( .A0(n7637), .A1(\s01.dbus_in [12]), .S(n7704), .Z(n4974) );
  CMX2X1 U8103 ( .A0(n7626), .A1(\s01.dbus_in [10]), .S(n7704), .Z(n4972) );
  CMX2X1 U8104 ( .A0(n7627), .A1(\s12.dbus_in [13]), .S(n7724), .Z(n5183) );
  CMX2X1 U8105 ( .A0(n7685), .A1(\s01.dbus_in [8]), .S(n7704), .Z(n4970) );
  CMX2X1 U8106 ( .A0(n7686), .A1(\s01.dbus_in [6]), .S(n7704), .Z(n4968) );
  CMX2X1 U8107 ( .A0(n7653), .A1(\s01.dbus_in [4]), .S(n7704), .Z(n4966) );
  CMX2X1 U8108 ( .A0(n7634), .A1(\s02.Adr [4]), .S(n7638), .Z(n4918) );
  CMX2X1 U8109 ( .A0(n7655), .A1(\s02.Adr [3]), .S(n7638), .Z(n4917) );
  CMX2X1 U8110 ( .A0(n7635), .A1(\s02.dbus_in [15]), .S(n7638), .Z(n4913) );
  CMX2X1 U8111 ( .A0(n7627), .A1(\s02.dbus_in [13]), .S(n7638), .Z(n4911) );
  CMX2X1 U8112 ( .A0(n7628), .A1(\s02.dbus_in [11]), .S(n7638), .Z(n4909) );
  CMX2X1 U8113 ( .A0(n7629), .A1(\s02.dbus_in [7]), .S(n7638), .Z(n4905) );
  CMX2X1 U8114 ( .A0(n7630), .A1(\s02.dbus_in [5]), .S(n7638), .Z(n4903) );
  CMX2X1 U8115 ( .A0(n7631), .A1(\s02.dbus_in [3]), .S(n7638), .Z(n4901) );
  CMX2X1 U8116 ( .A0(n7683), .A1(\s02.dbus_in [2]), .S(n7638), .Z(n4900) );
  CMX2X1 U8117 ( .A0(n7632), .A1(\s02.dbus_in [1]), .S(n7638), .Z(n4899) );
  CMX2X1 U8118 ( .A0(n7684), .A1(\s02.dbus_in [0]), .S(n7638), .Z(n4898) );
  CMX2X1 U8119 ( .A0(n7633), .A1(\s03.Adr [8]), .S(n7706), .Z(n4858) );
  CMX2X1 U8120 ( .A0(n7654), .A1(\s03.Adr [5]), .S(n7706), .Z(n4855) );
  CMX2X1 U8121 ( .A0(n7634), .A1(\s03.Adr [4]), .S(n7706), .Z(n4854) );
  CMX2X1 U8122 ( .A0(n7655), .A1(\s03.Adr [3]), .S(n7706), .Z(n4853) );
  CMX2X1 U8123 ( .A0(n7687), .A1(\s03.Adr [1]), .S(n7706), .Z(n4851) );
  CMX2X1 U8124 ( .A0(n7635), .A1(\s03.dbus_in [15]), .S(n7706), .Z(n4849) );
  CMX2X1 U8125 ( .A0(n7636), .A1(\s03.dbus_in [14]), .S(n7706), .Z(n4848) );
  CMX2X1 U8126 ( .A0(n7637), .A1(\s03.dbus_in [12]), .S(n7706), .Z(n4846) );
  CMX2X1 U8127 ( .A0(n7682), .A1(\s03.dbus_in [9]), .S(n7706), .Z(n4843) );
  CMX2X1 U8128 ( .A0(n7685), .A1(\s03.dbus_in [8]), .S(n7706), .Z(n4842) );
  CMX2X1 U8129 ( .A0(n7686), .A1(\s03.dbus_in [6]), .S(n7706), .Z(n4840) );
  CMX2X1 U8130 ( .A0(n7653), .A1(\s03.dbus_in [4]), .S(n7706), .Z(n4838) );
  CMX2X1 U8131 ( .A0(n7683), .A1(\s03.dbus_in [2]), .S(n7706), .Z(n4836) );
  CMX2X1 U8132 ( .A0(n7684), .A1(\s03.dbus_in [0]), .S(n7706), .Z(n4834) );
  CMX2X1 U8133 ( .A0(n7634), .A1(\s04.Adr [4]), .S(n7708), .Z(n4790) );
  CMX2X1 U8134 ( .A0(n7635), .A1(\s04.dbus_in [15]), .S(n7708), .Z(n4785) );
  CMX2X1 U8135 ( .A0(n7636), .A1(\s04.dbus_in [14]), .S(n7708), .Z(n4784) );
  CMX2X1 U8136 ( .A0(n7637), .A1(\s04.dbus_in [12]), .S(n7708), .Z(n4782) );
  CMX2X1 U8137 ( .A0(n7682), .A1(\s04.dbus_in [9]), .S(n7708), .Z(n4779) );
  CMX2X1 U8138 ( .A0(n7685), .A1(\s04.dbus_in [8]), .S(n7708), .Z(n4778) );
  CMX2X1 U8139 ( .A0(n7686), .A1(\s04.dbus_in [6]), .S(n7708), .Z(n4776) );
  CMX2X1 U8140 ( .A0(n7653), .A1(\s04.dbus_in [4]), .S(n7708), .Z(n4774) );
  CMX2X1 U8141 ( .A0(n7637), .A1(\s11.dbus_in [12]), .S(n7722), .Z(n4334) );
  CIVXL U8142 ( .A(\clock.rst ), .Z(n7696) );
  CND2X1 U8143 ( .A(\s02.tarActive ), .B(n7696), .Z(n7639) );
  CND2X1 U8144 ( .A(n7639), .B(n7638), .Z(n5212) );
  CANR2X1 U8145 ( .A(\m05.addrM [9]), .B(n7641), .C(n7640), .D(\m06.addrM [9]), 
        .Z(n7651) );
  CANR2XL U8146 ( .A(\m00.YouGotIt ), .B(\m00.addrM [9]), .C(\m01.addrM [9]), 
        .D(n7642), .Z(n7646) );
  CANR2X1 U8147 ( .A(\m03.addrM [9]), .B(n7644), .C(\m02.addrM [9]), .D(n7643), 
        .Z(n7645) );
  CND2X1 U8148 ( .A(n7646), .B(n7645), .Z(n7647) );
  CANR1XL U8149 ( .A(n7648), .B(\m04.addrM [9]), .C(n7647), .Z(n7650) );
  CND2X1 U8150 ( .A(n7702), .B(\s00.Adr [9]), .Z(n7649) );
  COND4CX1 U8151 ( .A(n7651), .B(n7650), .C(n7702), .D(n7649), .Z(n5067) );
  CAOR2XL U8152 ( .A(n7696), .B(\m01.YouGotIt ), .C(n7652), .D(\m01.need ), 
        .Z(n5265) );
  CMX2X1 U8153 ( .A0(n7653), .A1(\s11.dbus_in [4]), .S(n7722), .Z(n4326) );
  CMX2X1 U8154 ( .A0(n7654), .A1(\s12.Adr [5]), .S(n7724), .Z(n4279) );
  CMX2X1 U8155 ( .A0(n7655), .A1(\s12.Adr [3]), .S(n7724), .Z(n4277) );
  CIVX2 U8156 ( .A(\m06.DinMast [8]), .Z(n7681) );
  CAOR2X2 U8157 ( .A(\s05.dataOut [8]), .B(n7657), .C(\s04.dataOut [8]), .D(
        n7656), .Z(n7677) );
  CIVX2 U8158 ( .A(\s10.dataOut [8]), .Z(n7675) );
  CANR2XL U8159 ( .A(\s06.dataOut [8]), .B(n7659), .C(\s01.dataOut [8]), .D(
        n7658), .Z(n7673) );
  CANR2X1 U8160 ( .A(\s13.dataOut [8]), .B(n7661), .C(\s02.dataOut [8]), .D(
        n7660), .Z(n7671) );
  CANR2X1 U8161 ( .A(n7663), .B(\s03.dataOut [8]), .C(\s08.dataOut [8]), .D(
        n7662), .Z(n7670) );
  CANR2XL U8162 ( .A(\s12.dataOut [8]), .B(n7665), .C(\s11.dataOut [8]), .D(
        n7664), .Z(n7669) );
  CANR2X1 U8163 ( .A(\s07.dataOut [8]), .B(n7667), .C(\s09.dataOut [8]), .D(
        n7666), .Z(n7668) );
  CAN4X1 U8164 ( .A(n7671), .B(n7670), .C(n7669), .D(n7668), .Z(n7672) );
  COND3X1 U8165 ( .A(n7675), .B(n7674), .C(n7673), .D(n7672), .Z(n7676) );
  CANR3X1 U8166 ( .A(n7678), .B(\s00.dataOut [8]), .C(n7677), .D(n7676), .Z(
        n7680) );
  CMXI2X1 U8167 ( .A0(n7681), .A1(n7680), .S(n7679), .Z(n5194) );
  CMX2X1 U8168 ( .A0(n7682), .A1(\s11.dbus_in [9]), .S(n7722), .Z(n4331) );
  CMX2X1 U8169 ( .A0(n7683), .A1(\s11.dbus_in [2]), .S(n7722), .Z(n4324) );
  CMX2X1 U8170 ( .A0(n7684), .A1(\s11.dbus_in [0]), .S(n7722), .Z(n4322) );
  CMX2X1 U8171 ( .A0(n7685), .A1(\s11.dbus_in [8]), .S(n7722), .Z(n4330) );
  CMX2X1 U8172 ( .A0(n7686), .A1(\s11.dbus_in [6]), .S(n7722), .Z(n4328) );
  CMX2X1 U8173 ( .A0(n7687), .A1(\s12.Adr [1]), .S(n7724), .Z(n4275) );
  CNIVXL U8174 ( .A(\clock.sysClk ), .Z(n7741) );
  CNIVXL U8175 ( .A(\clock.sysClk ), .Z(n7746) );
  CNIVXL U8176 ( .A(\clock.sysClk ), .Z(n7739) );
  CNIVX1 U8177 ( .A(n7734), .Z(n7740) );
  CIVX2 U8178 ( .A(\m00.need ), .Z(n7688) );
  COND2XL U8179 ( .A(\clock.rst ), .B(n7690), .C(n7689), .D(n7688), .Z(n5225)
         );
  CAOR2XL U8180 ( .A(\m03.YouGotIt ), .B(n7696), .C(\m03.need ), .D(n7691), 
        .Z(n5255) );
  CIVX2 U8181 ( .A(\m05.need ), .Z(n7692) );
  COND2XL U8182 ( .A(\clock.rst ), .B(n7694), .C(n7693), .D(n7692), .Z(n5245)
         );
  CAOR2XL U8183 ( .A(\m04.YouGotIt ), .B(n7696), .C(n7695), .D(\m04.need ), 
        .Z(n5235) );
  CNIVXL U8184 ( .A(\clock.sysClk ), .Z(n7738) );
  CNIVXL U8185 ( .A(\clock.sysClk ), .Z(n7733) );
  CND2X1 U8748 ( .A(n7697), .B(\m02.need ), .Z(n7698) );
  COND1XL U8749 ( .A(n7699), .B(\clock.rst ), .C(n7698), .Z(n5275) );
  CIVX2 U8750 ( .A(\s13.tarActive ), .Z(n7701) );
  COND1XL U8751 ( .A(\clock.rst ), .B(n7701), .C(n7700), .Z(n5224) );
  CIVX2 U8752 ( .A(\s00.tarActive ), .Z(n7703) );
  COND1XL U8753 ( .A(\clock.rst ), .B(n7703), .C(n7702), .Z(n5214) );
  CIVX2 U8754 ( .A(\s01.tarActive ), .Z(n7705) );
  COND1XL U8755 ( .A(\clock.rst ), .B(n7705), .C(n7704), .Z(n5213) );
  CIVX2 U8756 ( .A(\s03.tarActive ), .Z(n7707) );
  COND1XL U8757 ( .A(\clock.rst ), .B(n7707), .C(n7706), .Z(n5211) );
  CIVX2 U8758 ( .A(\s04.tarActive ), .Z(n7709) );
  COND1XL U8759 ( .A(\clock.rst ), .B(n7709), .C(n7708), .Z(n5210) );
  CIVX2 U8760 ( .A(\s05.tarActive ), .Z(n7711) );
  COND1XL U8761 ( .A(\clock.rst ), .B(n7711), .C(n7710), .Z(n5209) );
  CIVX2 U8762 ( .A(\s06.tarActive ), .Z(n7713) );
  COND1XL U8763 ( .A(\clock.rst ), .B(n7713), .C(n7712), .Z(n5208) );
  CIVX2 U8764 ( .A(\s07.tarActive ), .Z(n7715) );
  COND1XL U8765 ( .A(\clock.rst ), .B(n7715), .C(n7714), .Z(n5207) );
  CIVX2 U8766 ( .A(\s08.tarActive ), .Z(n7717) );
  COND1XL U8767 ( .A(\clock.rst ), .B(n7717), .C(n7716), .Z(n5206) );
  CIVX2 U8768 ( .A(\s09.tarActive ), .Z(n7719) );
  COND1XL U8769 ( .A(\clock.rst ), .B(n7719), .C(n7718), .Z(n5205) );
  CIVX2 U8770 ( .A(\s10.tarActive ), .Z(n7721) );
  COND1XL U8771 ( .A(\clock.rst ), .B(n7721), .C(n7720), .Z(n5204) );
  CIVX2 U8772 ( .A(\s11.tarActive ), .Z(n7723) );
  COND1XL U8773 ( .A(\clock.rst ), .B(n7723), .C(n7722), .Z(n5203) );
  CIVX2 U8774 ( .A(\s12.tarActive ), .Z(n7725) );
  COND1XL U8775 ( .A(\clock.rst ), .B(n7725), .C(n7724), .Z(n5202) );
endmodule

