
module gpr ( clk, RegWrite, rd_addr1, rd_addr2, wr_addr, wr_data, rd_data2, 
        \rd_data1[31]_BAR , \rd_data1[30] , \rd_data1[29] , \rd_data1[28] , 
        \rd_data1[27] , \rd_data1[26] , \rd_data1[25] , \rd_data1[24] , 
        \rd_data1[23] , \rd_data1[22] , \rd_data1[21] , \rd_data1[20] , 
        \rd_data1[19] , \rd_data1[17] , \rd_data1[16] , \rd_data1[15] , 
        \rd_data1[14] , \rd_data1[13] , \rd_data1[12] , \rd_data1[11] , 
        \rd_data1[10] , \rd_data1[9] , \rd_data1[8] , \rd_data1[7] , 
        \rd_data1[6] , \rd_data1[5] , \rd_data1[4] , \rd_data1[3] , 
        \rd_data1[2] , \rd_data1[1] , \rd_data1[0] , \rd_data1[18]_BAR  );
  input [4:0] rd_addr1;
  input [4:0] rd_addr2;
  input [4:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_data2;
  input clk, RegWrite;
  output \rd_data1[31]_BAR , \rd_data1[30] , \rd_data1[29] , \rd_data1[28] ,
         \rd_data1[27] , \rd_data1[26] , \rd_data1[25] , \rd_data1[24] ,
         \rd_data1[23] , \rd_data1[22] , \rd_data1[21] , \rd_data1[20] ,
         \rd_data1[19] , \rd_data1[17] , \rd_data1[16] , \rd_data1[15] ,
         \rd_data1[14] , \rd_data1[13] , \rd_data1[12] , \rd_data1[11] ,
         \rd_data1[10] , \rd_data1[9] , \rd_data1[8] , \rd_data1[7] ,
         \rd_data1[6] , \rd_data1[5] , \rd_data1[4] , \rd_data1[3] ,
         \rd_data1[2] , \rd_data1[1] , \rd_data1[0] , \rd_data1[18]_BAR ;
  wire   \gpr[1][31] , \gpr[1][30] , \gpr[1][29] , \gpr[1][28] , \gpr[1][27] ,
         \gpr[1][26] , \gpr[1][25] , \gpr[1][24] , \gpr[1][23] , \gpr[1][22] ,
         \gpr[1][21] , \gpr[1][20] , \gpr[1][19] , \gpr[1][18] , \gpr[1][17] ,
         \gpr[1][16] , \gpr[1][15] , \gpr[1][14] , \gpr[1][13] , \gpr[1][12] ,
         \gpr[1][11] , \gpr[1][10] , \gpr[1][9] , \gpr[1][8] , \gpr[1][7] ,
         \gpr[1][6] , \gpr[1][5] , \gpr[1][4] , \gpr[1][3] , \gpr[1][2] ,
         \gpr[1][1] , \gpr[1][0] , \gpr[2][31] , \gpr[2][30] , \gpr[2][29] ,
         \gpr[2][28] , \gpr[2][27] , \gpr[2][26] , \gpr[2][25] , \gpr[2][24] ,
         \gpr[2][23] , \gpr[2][22] , \gpr[2][21] , \gpr[2][20] , \gpr[2][19] ,
         \gpr[2][18] , \gpr[2][17] , \gpr[2][16] , \gpr[2][15] , \gpr[2][14] ,
         \gpr[2][13] , \gpr[2][12] , \gpr[2][11] , \gpr[2][10] , \gpr[2][9] ,
         \gpr[2][8] , \gpr[2][7] , \gpr[2][6] , \gpr[2][5] , \gpr[2][4] ,
         \gpr[2][3] , \gpr[2][2] , \gpr[2][1] , \gpr[2][0] , \gpr[3][31] ,
         \gpr[3][30] , \gpr[3][29] , \gpr[3][28] , \gpr[3][27] , \gpr[3][26] ,
         \gpr[3][25] , \gpr[3][24] , \gpr[3][23] , \gpr[3][22] , \gpr[3][21] ,
         \gpr[3][20] , \gpr[3][19] , \gpr[3][18] , \gpr[3][17] , \gpr[3][16] ,
         \gpr[3][15] , \gpr[3][14] , \gpr[3][13] , \gpr[3][12] , \gpr[3][11] ,
         \gpr[3][10] , \gpr[3][9] , \gpr[3][8] , \gpr[3][7] , \gpr[3][6] ,
         \gpr[3][5] , \gpr[3][4] , \gpr[3][3] , \gpr[3][2] , \gpr[3][1] ,
         \gpr[3][0] , \gpr[4][31] , \gpr[4][30] , \gpr[4][29] , \gpr[4][28] ,
         \gpr[4][27] , \gpr[4][26] , \gpr[4][25] , \gpr[4][24] , \gpr[4][23] ,
         \gpr[4][22] , \gpr[4][21] , \gpr[4][20] , \gpr[4][19] , \gpr[4][18] ,
         \gpr[4][17] , \gpr[4][16] , \gpr[4][15] , \gpr[4][14] , \gpr[4][13] ,
         \gpr[4][12] , \gpr[4][11] , \gpr[4][10] , \gpr[4][9] , \gpr[4][8] ,
         \gpr[4][7] , \gpr[4][6] , \gpr[4][5] , \gpr[4][4] , \gpr[4][3] ,
         \gpr[4][2] , \gpr[4][1] , \gpr[4][0] , \gpr[5][31] , \gpr[5][30] ,
         \gpr[5][29] , \gpr[5][28] , \gpr[5][27] , \gpr[5][26] , \gpr[5][25] ,
         \gpr[5][24] , \gpr[5][23] , \gpr[5][22] , \gpr[5][21] , \gpr[5][20] ,
         \gpr[5][19] , \gpr[5][18] , \gpr[5][17] , \gpr[5][16] , \gpr[5][15] ,
         \gpr[5][14] , \gpr[5][13] , \gpr[5][12] , \gpr[5][11] , \gpr[5][10] ,
         \gpr[5][9] , \gpr[5][8] , \gpr[5][7] , \gpr[5][6] , \gpr[5][5] ,
         \gpr[5][4] , \gpr[5][3] , \gpr[5][2] , \gpr[5][1] , \gpr[5][0] ,
         \gpr[6][31] , \gpr[6][30] , \gpr[6][29] , \gpr[6][28] , \gpr[6][27] ,
         \gpr[6][26] , \gpr[6][25] , \gpr[6][24] , \gpr[6][23] , \gpr[6][22] ,
         \gpr[6][21] , \gpr[6][20] , \gpr[6][19] , \gpr[6][18] , \gpr[6][17] ,
         \gpr[6][16] , \gpr[6][15] , \gpr[6][14] , \gpr[6][13] , \gpr[6][12] ,
         \gpr[6][11] , \gpr[6][10] , \gpr[6][9] , \gpr[6][8] , \gpr[6][7] ,
         \gpr[6][6] , \gpr[6][5] , \gpr[6][4] , \gpr[6][3] , \gpr[6][2] ,
         \gpr[6][1] , \gpr[6][0] , \gpr[7][31] , \gpr[7][30] , \gpr[7][29] ,
         \gpr[7][28] , \gpr[7][27] , \gpr[7][26] , \gpr[7][25] , \gpr[7][24] ,
         \gpr[7][23] , \gpr[7][22] , \gpr[7][21] , \gpr[7][20] , \gpr[7][19] ,
         \gpr[7][18] , \gpr[7][17] , \gpr[7][16] , \gpr[7][15] , \gpr[7][14] ,
         \gpr[7][13] , \gpr[7][12] , \gpr[7][11] , \gpr[7][10] , \gpr[7][9] ,
         \gpr[7][8] , \gpr[7][7] , \gpr[7][6] , \gpr[7][5] , \gpr[7][4] ,
         \gpr[7][3] , \gpr[7][2] , \gpr[7][1] , \gpr[7][0] , \gpr[8][31] ,
         \gpr[8][30] , \gpr[8][29] , \gpr[8][28] , \gpr[8][27] , \gpr[8][26] ,
         \gpr[8][25] , \gpr[8][24] , \gpr[8][23] , \gpr[8][22] , \gpr[8][21] ,
         \gpr[8][20] , \gpr[8][19] , \gpr[8][18] , \gpr[8][17] , \gpr[8][16] ,
         \gpr[8][15] , \gpr[8][14] , \gpr[8][13] , \gpr[8][12] , \gpr[8][11] ,
         \gpr[8][10] , \gpr[8][9] , \gpr[8][8] , \gpr[8][7] , \gpr[8][6] ,
         \gpr[8][5] , \gpr[8][4] , \gpr[8][3] , \gpr[8][2] , \gpr[8][1] ,
         \gpr[8][0] , \gpr[9][31] , \gpr[9][30] , \gpr[9][29] , \gpr[9][28] ,
         \gpr[9][27] , \gpr[9][26] , \gpr[9][25] , \gpr[9][24] , \gpr[9][23] ,
         \gpr[9][22] , \gpr[9][21] , \gpr[9][20] , \gpr[9][19] , \gpr[9][18] ,
         \gpr[9][17] , \gpr[9][16] , \gpr[9][15] , \gpr[9][14] , \gpr[9][13] ,
         \gpr[9][12] , \gpr[9][11] , \gpr[9][10] , \gpr[9][9] , \gpr[9][8] ,
         \gpr[9][7] , \gpr[9][6] , \gpr[9][5] , \gpr[9][4] , \gpr[9][3] ,
         \gpr[9][2] , \gpr[9][1] , \gpr[9][0] , \gpr[10][31] , \gpr[10][30] ,
         \gpr[10][29] , \gpr[10][28] , \gpr[10][27] , \gpr[10][26] ,
         \gpr[10][25] , \gpr[10][24] , \gpr[10][23] , \gpr[10][22] ,
         \gpr[10][21] , \gpr[10][20] , \gpr[10][19] , \gpr[10][18] ,
         \gpr[10][17] , \gpr[10][16] , \gpr[10][15] , \gpr[10][14] ,
         \gpr[10][13] , \gpr[10][12] , \gpr[10][11] , \gpr[10][10] ,
         \gpr[10][9] , \gpr[10][8] , \gpr[10][7] , \gpr[10][6] , \gpr[10][5] ,
         \gpr[10][4] , \gpr[10][3] , \gpr[10][2] , \gpr[10][1] , \gpr[10][0] ,
         \gpr[11][31] , \gpr[11][30] , \gpr[11][29] , \gpr[11][28] ,
         \gpr[11][27] , \gpr[11][26] , \gpr[11][25] , \gpr[11][24] ,
         \gpr[11][23] , \gpr[11][22] , \gpr[11][21] , \gpr[11][20] ,
         \gpr[11][19] , \gpr[11][18] , \gpr[11][17] , \gpr[11][16] ,
         \gpr[11][15] , \gpr[11][14] , \gpr[11][13] , \gpr[11][12] ,
         \gpr[11][11] , \gpr[11][10] , \gpr[11][9] , \gpr[11][8] ,
         \gpr[11][7] , \gpr[11][6] , \gpr[11][5] , \gpr[11][4] , \gpr[11][3] ,
         \gpr[11][2] , \gpr[11][1] , \gpr[11][0] , \gpr[12][31] ,
         \gpr[12][30] , \gpr[12][29] , \gpr[12][28] , \gpr[12][27] ,
         \gpr[12][26] , \gpr[12][25] , \gpr[12][24] , \gpr[12][23] ,
         \gpr[12][22] , \gpr[12][21] , \gpr[12][20] , \gpr[12][19] ,
         \gpr[12][18] , \gpr[12][17] , \gpr[12][16] , \gpr[12][15] ,
         \gpr[12][14] , \gpr[12][13] , \gpr[12][12] , \gpr[12][11] ,
         \gpr[12][10] , \gpr[12][9] , \gpr[12][8] , \gpr[12][7] , \gpr[12][6] ,
         \gpr[12][5] , \gpr[12][4] , \gpr[12][3] , \gpr[12][2] , \gpr[12][1] ,
         \gpr[12][0] , \gpr[13][31] , \gpr[13][30] , \gpr[13][29] ,
         \gpr[13][28] , \gpr[13][27] , \gpr[13][26] , \gpr[13][25] ,
         \gpr[13][24] , \gpr[13][23] , \gpr[13][22] , \gpr[13][21] ,
         \gpr[13][20] , \gpr[13][19] , \gpr[13][18] , \gpr[13][17] ,
         \gpr[13][16] , \gpr[13][15] , \gpr[13][14] , \gpr[13][13] ,
         \gpr[13][12] , \gpr[13][11] , \gpr[13][10] , \gpr[13][9] ,
         \gpr[13][8] , \gpr[13][7] , \gpr[13][6] , \gpr[13][5] , \gpr[13][4] ,
         \gpr[13][3] , \gpr[13][2] , \gpr[13][1] , \gpr[13][0] , \gpr[14][31] ,
         \gpr[14][30] , \gpr[14][29] , \gpr[14][28] , \gpr[14][27] ,
         \gpr[14][26] , \gpr[14][25] , \gpr[14][24] , \gpr[14][23] ,
         \gpr[14][22] , \gpr[14][21] , \gpr[14][20] , \gpr[14][19] ,
         \gpr[14][18] , \gpr[14][17] , \gpr[14][16] , \gpr[14][15] ,
         \gpr[14][14] , \gpr[14][13] , \gpr[14][12] , \gpr[14][11] ,
         \gpr[14][10] , \gpr[14][9] , \gpr[14][8] , \gpr[14][7] , \gpr[14][6] ,
         \gpr[14][5] , \gpr[14][4] , \gpr[14][3] , \gpr[14][2] , \gpr[14][1] ,
         \gpr[14][0] , \gpr[15][31] , \gpr[15][30] , \gpr[15][29] ,
         \gpr[15][28] , \gpr[15][27] , \gpr[15][26] , \gpr[15][25] ,
         \gpr[15][24] , \gpr[15][23] , \gpr[15][22] , \gpr[15][21] ,
         \gpr[15][20] , \gpr[15][19] , \gpr[15][18] , \gpr[15][17] ,
         \gpr[15][16] , \gpr[15][15] , \gpr[15][14] , \gpr[15][13] ,
         \gpr[15][12] , \gpr[15][11] , \gpr[15][10] , \gpr[15][9] ,
         \gpr[15][8] , \gpr[15][7] , \gpr[15][6] , \gpr[15][5] , \gpr[15][4] ,
         \gpr[15][3] , \gpr[15][2] , \gpr[15][1] , \gpr[15][0] , \gpr[16][31] ,
         \gpr[16][30] , \gpr[16][29] , \gpr[16][28] , \gpr[16][27] ,
         \gpr[16][26] , \gpr[16][25] , \gpr[16][24] , \gpr[16][23] ,
         \gpr[16][22] , \gpr[16][21] , \gpr[16][20] , \gpr[16][19] ,
         \gpr[16][18] , \gpr[16][17] , \gpr[16][16] , \gpr[16][15] ,
         \gpr[16][14] , \gpr[16][13] , \gpr[16][12] , \gpr[16][11] ,
         \gpr[16][10] , \gpr[16][9] , \gpr[16][8] , \gpr[16][7] , \gpr[16][6] ,
         \gpr[16][5] , \gpr[16][4] , \gpr[16][3] , \gpr[16][2] , \gpr[16][1] ,
         \gpr[16][0] , \gpr[17][31] , \gpr[17][30] , \gpr[17][29] ,
         \gpr[17][28] , \gpr[17][27] , \gpr[17][26] , \gpr[17][25] ,
         \gpr[17][24] , \gpr[17][23] , \gpr[17][22] , \gpr[17][21] ,
         \gpr[17][20] , \gpr[17][19] , \gpr[17][18] , \gpr[17][17] ,
         \gpr[17][16] , \gpr[17][15] , \gpr[17][14] , \gpr[17][13] ,
         \gpr[17][12] , \gpr[17][11] , \gpr[17][10] , \gpr[17][9] ,
         \gpr[17][8] , \gpr[17][7] , \gpr[17][6] , \gpr[17][5] , \gpr[17][4] ,
         \gpr[17][3] , \gpr[17][2] , \gpr[17][1] , \gpr[17][0] , \gpr[18][31] ,
         \gpr[18][30] , \gpr[18][29] , \gpr[18][28] , \gpr[18][27] ,
         \gpr[18][26] , \gpr[18][25] , \gpr[18][24] , \gpr[18][23] ,
         \gpr[18][22] , \gpr[18][21] , \gpr[18][20] , \gpr[18][19] ,
         \gpr[18][18] , \gpr[18][17] , \gpr[18][16] , \gpr[18][15] ,
         \gpr[18][14] , \gpr[18][13] , \gpr[18][12] , \gpr[18][11] ,
         \gpr[18][10] , \gpr[18][9] , \gpr[18][8] , \gpr[18][7] , \gpr[18][6] ,
         \gpr[18][5] , \gpr[18][4] , \gpr[18][3] , \gpr[18][2] , \gpr[18][1] ,
         \gpr[18][0] , \gpr[19][31] , \gpr[19][30] , \gpr[19][29] ,
         \gpr[19][28] , \gpr[19][27] , \gpr[19][26] , \gpr[19][25] ,
         \gpr[19][24] , \gpr[19][23] , \gpr[19][22] , \gpr[19][21] ,
         \gpr[19][20] , \gpr[19][19] , \gpr[19][18] , \gpr[19][17] ,
         \gpr[19][16] , \gpr[19][15] , \gpr[19][14] , \gpr[19][13] ,
         \gpr[19][12] , \gpr[19][11] , \gpr[19][10] , \gpr[19][9] ,
         \gpr[19][8] , \gpr[19][7] , \gpr[19][6] , \gpr[19][5] , \gpr[19][4] ,
         \gpr[19][3] , \gpr[19][2] , \gpr[19][1] , \gpr[19][0] , \gpr[20][31] ,
         \gpr[20][30] , \gpr[20][29] , \gpr[20][28] , \gpr[20][27] ,
         \gpr[20][26] , \gpr[20][25] , \gpr[20][24] , \gpr[20][23] ,
         \gpr[20][22] , \gpr[20][21] , \gpr[20][20] , \gpr[20][19] ,
         \gpr[20][18] , \gpr[20][17] , \gpr[20][16] , \gpr[20][15] ,
         \gpr[20][14] , \gpr[20][13] , \gpr[20][12] , \gpr[20][11] ,
         \gpr[20][10] , \gpr[20][9] , \gpr[20][8] , \gpr[20][7] , \gpr[20][6] ,
         \gpr[20][5] , \gpr[20][4] , \gpr[20][3] , \gpr[20][2] , \gpr[20][1] ,
         \gpr[20][0] , \gpr[21][31] , \gpr[21][30] , \gpr[21][29] ,
         \gpr[21][28] , \gpr[21][27] , \gpr[21][26] , \gpr[21][25] ,
         \gpr[21][24] , \gpr[21][23] , \gpr[21][22] , \gpr[21][21] ,
         \gpr[21][20] , \gpr[21][19] , \gpr[21][18] , \gpr[21][17] ,
         \gpr[21][16] , \gpr[21][15] , \gpr[21][14] , \gpr[21][13] ,
         \gpr[21][12] , \gpr[21][11] , \gpr[21][10] , \gpr[21][9] ,
         \gpr[21][8] , \gpr[21][7] , \gpr[21][6] , \gpr[21][5] , \gpr[21][4] ,
         \gpr[21][3] , \gpr[21][2] , \gpr[21][1] , \gpr[21][0] , \gpr[22][31] ,
         \gpr[22][30] , \gpr[22][29] , \gpr[22][28] , \gpr[22][27] ,
         \gpr[22][26] , \gpr[22][25] , \gpr[22][24] , \gpr[22][23] ,
         \gpr[22][22] , \gpr[22][21] , \gpr[22][20] , \gpr[22][19] ,
         \gpr[22][18] , \gpr[22][17] , \gpr[22][16] , \gpr[22][15] ,
         \gpr[22][14] , \gpr[22][13] , \gpr[22][12] , \gpr[22][11] ,
         \gpr[22][10] , \gpr[22][9] , \gpr[22][8] , \gpr[22][7] , \gpr[22][6] ,
         \gpr[22][5] , \gpr[22][4] , \gpr[22][3] , \gpr[22][2] , \gpr[22][1] ,
         \gpr[22][0] , \gpr[23][31] , \gpr[23][30] , \gpr[23][29] ,
         \gpr[23][28] , \gpr[23][27] , \gpr[23][26] , \gpr[23][25] ,
         \gpr[23][24] , \gpr[23][23] , \gpr[23][22] , \gpr[23][21] ,
         \gpr[23][20] , \gpr[23][19] , \gpr[23][18] , \gpr[23][17] ,
         \gpr[23][16] , \gpr[23][15] , \gpr[23][14] , \gpr[23][13] ,
         \gpr[23][12] , \gpr[23][11] , \gpr[23][10] , \gpr[23][9] ,
         \gpr[23][8] , \gpr[23][7] , \gpr[23][6] , \gpr[23][5] , \gpr[23][4] ,
         \gpr[23][3] , \gpr[23][2] , \gpr[23][1] , \gpr[23][0] , \gpr[24][31] ,
         \gpr[24][30] , \gpr[24][29] , \gpr[24][28] , \gpr[24][27] ,
         \gpr[24][26] , \gpr[24][25] , \gpr[24][24] , \gpr[24][23] ,
         \gpr[24][22] , \gpr[24][21] , \gpr[24][20] , \gpr[24][19] ,
         \gpr[24][18] , \gpr[24][17] , \gpr[24][16] , \gpr[24][15] ,
         \gpr[24][14] , \gpr[24][13] , \gpr[24][12] , \gpr[24][11] ,
         \gpr[24][10] , \gpr[24][9] , \gpr[24][8] , \gpr[24][7] , \gpr[24][6] ,
         \gpr[24][5] , \gpr[24][4] , \gpr[24][3] , \gpr[24][2] , \gpr[24][1] ,
         \gpr[24][0] , \gpr[25][31] , \gpr[25][30] , \gpr[25][29] ,
         \gpr[25][28] , \gpr[25][27] , \gpr[25][26] , \gpr[25][25] ,
         \gpr[25][24] , \gpr[25][23] , \gpr[25][22] , \gpr[25][21] ,
         \gpr[25][20] , \gpr[25][19] , \gpr[25][18] , \gpr[25][17] ,
         \gpr[25][16] , \gpr[25][15] , \gpr[25][14] , \gpr[25][13] ,
         \gpr[25][12] , \gpr[25][11] , \gpr[25][10] , \gpr[25][9] ,
         \gpr[25][8] , \gpr[25][7] , \gpr[25][6] , \gpr[25][5] , \gpr[25][4] ,
         \gpr[25][3] , \gpr[25][2] , \gpr[25][1] , \gpr[25][0] , \gpr[26][31] ,
         \gpr[26][30] , \gpr[26][29] , \gpr[26][28] , \gpr[26][27] ,
         \gpr[26][26] , \gpr[26][25] , \gpr[26][24] , \gpr[26][23] ,
         \gpr[26][22] , \gpr[26][21] , \gpr[26][20] , \gpr[26][19] ,
         \gpr[26][18] , \gpr[26][17] , \gpr[26][16] , \gpr[26][15] ,
         \gpr[26][14] , \gpr[26][13] , \gpr[26][12] , \gpr[26][11] ,
         \gpr[26][10] , \gpr[26][9] , \gpr[26][8] , \gpr[26][7] , \gpr[26][6] ,
         \gpr[26][5] , \gpr[26][4] , \gpr[26][3] , \gpr[26][2] , \gpr[26][1] ,
         \gpr[26][0] , \gpr[27][31] , \gpr[27][30] , \gpr[27][29] ,
         \gpr[27][28] , \gpr[27][27] , \gpr[27][26] , \gpr[27][25] ,
         \gpr[27][24] , \gpr[27][23] , \gpr[27][22] , \gpr[27][21] ,
         \gpr[27][20] , \gpr[27][19] , \gpr[27][18] , \gpr[27][17] ,
         \gpr[27][16] , \gpr[27][15] , \gpr[27][14] , \gpr[27][13] ,
         \gpr[27][12] , \gpr[27][11] , \gpr[27][10] , \gpr[27][9] ,
         \gpr[27][8] , \gpr[27][7] , \gpr[27][6] , \gpr[27][5] , \gpr[27][4] ,
         \gpr[27][3] , \gpr[27][2] , \gpr[27][1] , \gpr[27][0] , \gpr[28][31] ,
         \gpr[28][30] , \gpr[28][29] , \gpr[28][28] , \gpr[28][27] ,
         \gpr[28][26] , \gpr[28][25] , \gpr[28][24] , \gpr[28][23] ,
         \gpr[28][22] , \gpr[28][21] , \gpr[28][20] , \gpr[28][19] ,
         \gpr[28][17] , \gpr[28][16] , \gpr[28][15] , \gpr[28][14] ,
         \gpr[28][13] , \gpr[28][12] , \gpr[28][11] , \gpr[28][10] ,
         \gpr[28][9] , \gpr[28][8] , \gpr[28][7] , \gpr[28][6] , \gpr[28][5] ,
         \gpr[28][4] , \gpr[28][3] , \gpr[28][2] , \gpr[28][1] , \gpr[28][0] ,
         \gpr[29][31] , \gpr[29][30] , \gpr[29][29] , \gpr[29][28] ,
         \gpr[29][27] , \gpr[29][26] , \gpr[29][25] , \gpr[29][24] ,
         \gpr[29][23] , \gpr[29][22] , \gpr[29][21] , \gpr[29][20] ,
         \gpr[29][19] , \gpr[29][18] , \gpr[29][17] , \gpr[29][16] ,
         \gpr[29][15] , \gpr[29][14] , \gpr[29][13] , \gpr[29][12] ,
         \gpr[29][11] , \gpr[29][10] , \gpr[29][9] , \gpr[29][8] ,
         \gpr[29][7] , \gpr[29][6] , \gpr[29][5] , \gpr[29][4] , \gpr[29][3] ,
         \gpr[29][2] , \gpr[29][1] , \gpr[29][0] , \gpr[30][30] ,
         \gpr[30][28] , \gpr[30][27] , \gpr[30][26] , \gpr[30][25] ,
         \gpr[30][24] , \gpr[30][23] , \gpr[30][22] , \gpr[30][21] ,
         \gpr[30][20] , \gpr[30][19] , \gpr[30][18] , \gpr[30][17] ,
         \gpr[30][16] , \gpr[30][15] , \gpr[30][14] , \gpr[30][13] ,
         \gpr[30][12] , \gpr[30][11] , \gpr[30][10] , \gpr[30][9] ,
         \gpr[30][8] , \gpr[30][7] , \gpr[30][6] , \gpr[30][5] , \gpr[30][4] ,
         \gpr[30][3] , \gpr[30][2] , \gpr[30][1] , \gpr[30][0] , \gpr[31][31] ,
         \gpr[31][30] , \gpr[31][29] , \gpr[31][28] , \gpr[31][27] ,
         \gpr[31][26] , \gpr[31][25] , \gpr[31][24] , \gpr[31][23] ,
         \gpr[31][22] , \gpr[31][21] , \gpr[31][20] , \gpr[31][19] ,
         \gpr[31][18] , \gpr[31][17] , \gpr[31][16] , \gpr[31][15] ,
         \gpr[31][14] , \gpr[31][13] , \gpr[31][12] , \gpr[31][11] ,
         \gpr[31][10] , \gpr[31][9] , \gpr[31][8] , \gpr[31][7] , \gpr[31][6] ,
         \gpr[31][5] , \gpr[31][4] , \gpr[31][3] , \gpr[31][2] , \gpr[31][1] ,
         \gpr[31][0] , n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724;
  wire   [31:0] rd_data1;

  FD1 \gpr_reg[1][31]  ( .D(n3346), .CP(clk), .Q(\gpr[1][31] ), .QN(n5667) );
  FD1 \gpr_reg[1][30]  ( .D(n3345), .CP(clk), .Q(\gpr[1][30] ), .QN(n5642) );
  FD1 \gpr_reg[1][29]  ( .D(n3344), .CP(clk), .Q(\gpr[1][29] ), .QN(n5614) );
  FD1 \gpr_reg[1][28]  ( .D(n3343), .CP(clk), .Q(\gpr[1][28] ), .QN(n5591) );
  FD1 \gpr_reg[1][26]  ( .D(n3341), .CP(clk), .Q(\gpr[1][26] ), .QN(n5540) );
  FD1 \gpr_reg[1][25]  ( .D(n3340), .CP(clk), .Q(\gpr[1][25] ), .QN(n5509) );
  FD1 \gpr_reg[1][24]  ( .D(n3339), .CP(clk), .Q(\gpr[1][24] ), .QN(n5492) );
  FD1 \gpr_reg[1][23]  ( .D(n3338), .CP(clk), .Q(\gpr[1][23] ), .QN(n5465) );
  FD1 \gpr_reg[1][21]  ( .D(n3336), .CP(clk), .Q(\gpr[1][21] ), .QN(n5421) );
  FD1 \gpr_reg[1][20]  ( .D(n3335), .CP(clk), .Q(\gpr[1][20] ), .QN(n5395) );
  FD1 \gpr_reg[1][19]  ( .D(n3334), .CP(clk), .Q(\gpr[1][19] ), .QN(n5369) );
  FD1 \gpr_reg[1][18]  ( .D(n3333), .CP(clk), .Q(\gpr[1][18] ), .QN(n311) );
  FD1 \gpr_reg[1][17]  ( .D(n3332), .CP(clk), .Q(\gpr[1][17] ), .QN(n5312) );
  FD1 \gpr_reg[1][16]  ( .D(n3331), .CP(clk), .Q(\gpr[1][16] ), .QN(n5303) );
  FD1 \gpr_reg[1][15]  ( .D(n3330), .CP(clk), .Q(\gpr[1][15] ), .QN(n5276) );
  FD1 \gpr_reg[1][14]  ( .D(n3329), .CP(clk), .Q(\gpr[1][14] ), .QN(n5250) );
  FD1 \gpr_reg[1][13]  ( .D(n3328), .CP(clk), .Q(\gpr[1][13] ), .QN(n5223) );
  FD1 \gpr_reg[1][10]  ( .D(n3325), .CP(clk), .Q(\gpr[1][10] ), .QN(n5153) );
  FD1 \gpr_reg[1][9]  ( .D(n3324), .CP(clk), .Q(\gpr[1][9] ), .QN(n5124) );
  FD1 \gpr_reg[1][8]  ( .D(n3323), .CP(clk), .Q(\gpr[1][8] ), .QN(n5097) );
  FD1 \gpr_reg[1][7]  ( .D(n3322), .CP(clk), .Q(\gpr[1][7] ), .QN(n5070) );
  FD1 \gpr_reg[1][6]  ( .D(n3321), .CP(clk), .Q(\gpr[1][6] ), .QN(n5045) );
  FD1 \gpr_reg[1][5]  ( .D(n3320), .CP(clk), .Q(\gpr[1][5] ), .QN(n5017) );
  FD1 \gpr_reg[1][3]  ( .D(n3318), .CP(clk), .Q(\gpr[1][3] ), .QN(n4972) );
  FD1 \gpr_reg[1][2]  ( .D(n3317), .CP(clk), .Q(\gpr[1][2] ), .QN(n4947) );
  FD1 \gpr_reg[1][1]  ( .D(n3316), .CP(clk), .Q(\gpr[1][1] ), .QN(n4920) );
  FD1 \gpr_reg[2][31]  ( .D(n3314), .CP(clk), .Q(\gpr[2][31] ), .QN(n5663) );
  FD1 \gpr_reg[2][30]  ( .D(n3313), .CP(clk), .Q(\gpr[2][30] ), .QN(n5638) );
  FD1 \gpr_reg[2][29]  ( .D(n3312), .CP(clk), .Q(\gpr[2][29] ), .QN(n5610) );
  FD1 \gpr_reg[2][28]  ( .D(n3311), .CP(clk), .Q(\gpr[2][28] ), .QN(n5587) );
  FD1 \gpr_reg[2][27]  ( .D(n3310), .CP(clk), .Q(\gpr[2][27] ), .QN(n5564) );
  FD1 \gpr_reg[2][26]  ( .D(n3309), .CP(clk), .Q(\gpr[2][26] ), .QN(n5536) );
  FD1 \gpr_reg[2][25]  ( .D(n3308), .CP(clk), .Q(\gpr[2][25] ), .QN(n5508) );
  FD1 \gpr_reg[2][24]  ( .D(n3307), .CP(clk), .Q(\gpr[2][24] ), .QN(n5488) );
  FD1 \gpr_reg[2][23]  ( .D(n3306), .CP(clk), .Q(\gpr[2][23] ), .QN(n5461) );
  FD1 \gpr_reg[2][22]  ( .D(n3305), .CP(clk), .Q(\gpr[2][22] ), .QN(n5442) );
  FD1 \gpr_reg[2][21]  ( .D(n3304), .CP(clk), .Q(\gpr[2][21] ), .QN(n5417) );
  FD1 \gpr_reg[2][20]  ( .D(n3303), .CP(clk), .Q(\gpr[2][20] ), .QN(n5391) );
  FD1 \gpr_reg[2][19]  ( .D(n3302), .CP(clk), .Q(\gpr[2][19] ), .QN(n5365) );
  FD1 \gpr_reg[2][18]  ( .D(n3301), .CP(clk), .Q(\gpr[2][18] ), .QN(n5344) );
  FD1 \gpr_reg[2][17]  ( .D(n3300), .CP(clk), .Q(\gpr[2][17] ), .QN(n5318) );
  FD1 \gpr_reg[2][16]  ( .D(n3299), .CP(clk), .Q(\gpr[2][16] ), .QN(n5299) );
  FD1 \gpr_reg[2][15]  ( .D(n3298), .CP(clk), .Q(\gpr[2][15] ), .QN(n5272) );
  FD1 \gpr_reg[2][14]  ( .D(n3297), .CP(clk), .Q(\gpr[2][14] ), .QN(n5246) );
  FD1 \gpr_reg[2][13]  ( .D(n3296), .CP(clk), .Q(\gpr[2][13] ), .QN(n5219) );
  FD1 \gpr_reg[2][12]  ( .D(n3295), .CP(clk), .Q(\gpr[2][12] ), .QN(n5197) );
  FD1 \gpr_reg[2][11]  ( .D(n3294), .CP(clk), .Q(\gpr[2][11] ), .QN(n5176) );
  FD1 \gpr_reg[2][10]  ( .D(n3293), .CP(clk), .Q(\gpr[2][10] ), .QN(n5149) );
  FD1 \gpr_reg[2][9]  ( .D(n3292), .CP(clk), .Q(\gpr[2][9] ), .QN(n5120) );
  FD1 \gpr_reg[2][8]  ( .D(n3291), .CP(clk), .Q(\gpr[2][8] ), .QN(n5093) );
  FD1 \gpr_reg[2][7]  ( .D(n3290), .CP(clk), .Q(\gpr[2][7] ), .QN(n5066) );
  FD1 \gpr_reg[2][6]  ( .D(n3289), .CP(clk), .Q(\gpr[2][6] ), .QN(n5041) );
  FD1 \gpr_reg[2][5]  ( .D(n3288), .CP(clk), .Q(\gpr[2][5] ), .QN(n5013) );
  FD1 \gpr_reg[2][4]  ( .D(n3287), .CP(clk), .Q(\gpr[2][4] ), .QN(n4992) );
  FD1 \gpr_reg[2][3]  ( .D(n3286), .CP(clk), .Q(\gpr[2][3] ), .QN(n4968) );
  FD1 \gpr_reg[2][2]  ( .D(n3285), .CP(clk), .Q(\gpr[2][2] ), .QN(n4943) );
  FD1 \gpr_reg[2][1]  ( .D(n3284), .CP(clk), .Q(\gpr[2][1] ), .QN(n4914) );
  FD1 \gpr_reg[2][0]  ( .D(n3283), .CP(clk), .Q(\gpr[2][0] ), .QN(n4899) );
  FD1 \gpr_reg[3][31]  ( .D(n3282), .CP(clk), .Q(\gpr[3][31] ), .QN(n5668) );
  FD1 \gpr_reg[3][30]  ( .D(n3281), .CP(clk), .Q(\gpr[3][30] ), .QN(n5643) );
  FD1 \gpr_reg[3][29]  ( .D(n3280), .CP(clk), .Q(\gpr[3][29] ), .QN(n5615) );
  FD1 \gpr_reg[3][28]  ( .D(n3279), .CP(clk), .Q(\gpr[3][28] ), .QN(n5592) );
  FD1 \gpr_reg[3][26]  ( .D(n3277), .CP(clk), .Q(\gpr[3][26] ), .QN(n5541) );
  FD1 \gpr_reg[3][25]  ( .D(n3276), .CP(clk), .Q(\gpr[3][25] ), .QN(n5510) );
  FD1 \gpr_reg[3][24]  ( .D(n3275), .CP(clk), .Q(\gpr[3][24] ), .QN(n5493) );
  FD1 \gpr_reg[3][23]  ( .D(n3274), .CP(clk), .Q(\gpr[3][23] ), .QN(n5466) );
  FD1 \gpr_reg[3][21]  ( .D(n3272), .CP(clk), .Q(\gpr[3][21] ), .QN(n5422) );
  FD1 \gpr_reg[3][20]  ( .D(n3271), .CP(clk), .Q(\gpr[3][20] ), .QN(n5396) );
  FD1 \gpr_reg[3][19]  ( .D(n3270), .CP(clk), .Q(\gpr[3][19] ), .QN(n5370) );
  FD1 \gpr_reg[3][18]  ( .D(n3269), .CP(clk), .Q(\gpr[3][18] ), .QN(n5346) );
  FD1 \gpr_reg[3][17]  ( .D(n3268), .CP(clk), .Q(\gpr[3][17] ), .QN(n5313) );
  FD1 \gpr_reg[3][16]  ( .D(n3267), .CP(clk), .Q(\gpr[3][16] ), .QN(n5304) );
  FD1 \gpr_reg[3][15]  ( .D(n3266), .CP(clk), .Q(\gpr[3][15] ), .QN(n5277) );
  FD1 \gpr_reg[3][14]  ( .D(n3265), .CP(clk), .Q(\gpr[3][14] ), .QN(n5251) );
  FD1 \gpr_reg[3][13]  ( .D(n3264), .CP(clk), .Q(\gpr[3][13] ), .QN(n5224) );
  FD1 \gpr_reg[3][10]  ( .D(n3261), .CP(clk), .Q(\gpr[3][10] ), .QN(n5154) );
  FD1 \gpr_reg[3][9]  ( .D(n3260), .CP(clk), .Q(\gpr[3][9] ), .QN(n5125) );
  FD1 \gpr_reg[3][8]  ( .D(n3259), .CP(clk), .Q(\gpr[3][8] ), .QN(n5098) );
  FD1 \gpr_reg[3][7]  ( .D(n3258), .CP(clk), .Q(\gpr[3][7] ), .QN(n5071) );
  FD1 \gpr_reg[3][6]  ( .D(n3257), .CP(clk), .Q(\gpr[3][6] ), .QN(n5046) );
  FD1 \gpr_reg[3][5]  ( .D(n3256), .CP(clk), .Q(\gpr[3][5] ), .QN(n5018) );
  FD1 \gpr_reg[3][3]  ( .D(n3254), .CP(clk), .Q(\gpr[3][3] ), .QN(n4973) );
  FD1 \gpr_reg[3][2]  ( .D(n3253), .CP(clk), .Q(\gpr[3][2] ), .QN(n4948) );
  FD1 \gpr_reg[3][1]  ( .D(n3252), .CP(clk), .Q(\gpr[3][1] ), .QN(n4915) );
  FD1 \gpr_reg[4][31]  ( .D(n3250), .CP(clk), .Q(\gpr[4][31] ), .QN(n5662) );
  FD1 \gpr_reg[4][30]  ( .D(n3249), .CP(clk), .Q(\gpr[4][30] ), .QN(n5637) );
  FD1 \gpr_reg[4][29]  ( .D(n3248), .CP(clk), .Q(\gpr[4][29] ), .QN(n5609) );
  FD1 \gpr_reg[4][28]  ( .D(n3247), .CP(clk), .Q(\gpr[4][28] ), .QN(n5586) );
  FD1 \gpr_reg[4][27]  ( .D(n3246), .CP(clk), .Q(\gpr[4][27] ), .QN(n5563) );
  FD1 \gpr_reg[4][26]  ( .D(n3245), .CP(clk), .Q(\gpr[4][26] ) );
  FD1 \gpr_reg[4][25]  ( .D(n3244), .CP(clk), .Q(\gpr[4][25] ), .QN(n5507) );
  FD1 \gpr_reg[4][24]  ( .D(n3243), .CP(clk), .Q(\gpr[4][24] ), .QN(n5487) );
  FD1 \gpr_reg[4][23]  ( .D(n3242), .CP(clk), .Q(\gpr[4][23] ), .QN(n5460) );
  FD1 \gpr_reg[4][22]  ( .D(n3241), .CP(clk), .Q(\gpr[4][22] ), .QN(n5441) );
  FD1 \gpr_reg[4][21]  ( .D(n3240), .CP(clk), .Q(\gpr[4][21] ), .QN(n5416) );
  FD1 \gpr_reg[4][20]  ( .D(n3239), .CP(clk), .Q(\gpr[4][20] ), .QN(n5390) );
  FD1 \gpr_reg[4][19]  ( .D(n3238), .CP(clk), .Q(\gpr[4][19] ), .QN(n5364) );
  FD1 \gpr_reg[4][17]  ( .D(n3236), .CP(clk), .Q(\gpr[4][17] ), .QN(n5311) );
  FD1 \gpr_reg[4][16]  ( .D(n3235), .CP(clk), .Q(\gpr[4][16] ), .QN(n5298) );
  FD1 \gpr_reg[4][15]  ( .D(n3234), .CP(clk), .Q(\gpr[4][15] ), .QN(n5271) );
  FD1 \gpr_reg[4][14]  ( .D(n3233), .CP(clk), .Q(\gpr[4][14] ), .QN(n5245) );
  FD1 \gpr_reg[4][13]  ( .D(n3232), .CP(clk), .Q(\gpr[4][13] ), .QN(n5218) );
  FD1 \gpr_reg[4][12]  ( .D(n3231), .CP(clk), .Q(\gpr[4][12] ), .QN(n5196) );
  FD1 \gpr_reg[4][11]  ( .D(n3230), .CP(clk), .Q(\gpr[4][11] ), .QN(n5175) );
  FD1 \gpr_reg[4][10]  ( .D(n3229), .CP(clk), .Q(\gpr[4][10] ), .QN(n5148) );
  FD1 \gpr_reg[4][9]  ( .D(n3228), .CP(clk), .Q(\gpr[4][9] ), .QN(n5119) );
  FD1 \gpr_reg[4][8]  ( .D(n3227), .CP(clk), .Q(\gpr[4][8] ), .QN(n5092) );
  FD1 \gpr_reg[4][7]  ( .D(n3226), .CP(clk), .Q(\gpr[4][7] ), .QN(n5065) );
  FD1 \gpr_reg[4][6]  ( .D(n3225), .CP(clk), .Q(\gpr[4][6] ), .QN(n5040) );
  FD1 \gpr_reg[4][5]  ( .D(n3224), .CP(clk), .Q(\gpr[4][5] ), .QN(n5012) );
  FD1 \gpr_reg[4][4]  ( .D(n3223), .CP(clk), .Q(\gpr[4][4] ), .QN(n4991) );
  FD1 \gpr_reg[4][3]  ( .D(n3222), .CP(clk), .Q(\gpr[4][3] ), .QN(n4967) );
  FD1 \gpr_reg[4][1]  ( .D(n3220), .CP(clk), .Q(\gpr[4][1] ), .QN(n4913) );
  FD1 \gpr_reg[4][0]  ( .D(n3219), .CP(clk), .Q(\gpr[4][0] ), .QN(n4898) );
  FD1 \gpr_reg[5][31]  ( .D(n3218), .CP(clk), .Q(\gpr[5][31] ), .QN(n5666) );
  FD1 \gpr_reg[5][30]  ( .D(n3217), .CP(clk), .Q(\gpr[5][30] ), .QN(n5641) );
  FD1 \gpr_reg[5][29]  ( .D(n3216), .CP(clk), .Q(\gpr[5][29] ), .QN(n5613) );
  FD1 \gpr_reg[5][28]  ( .D(n3215), .CP(clk), .Q(\gpr[5][28] ), .QN(n5590) );
  FD1 \gpr_reg[5][27]  ( .D(n3214), .CP(clk), .Q(\gpr[5][27] ) );
  FD1 \gpr_reg[5][26]  ( .D(n3213), .CP(clk), .Q(\gpr[5][26] ), .QN(n5539) );
  FD1 \gpr_reg[5][25]  ( .D(n3212), .CP(clk), .Q(\gpr[5][25] ), .QN(n5502) );
  FD1 \gpr_reg[5][24]  ( .D(n3211), .CP(clk), .Q(\gpr[5][24] ), .QN(n5491) );
  FD1 \gpr_reg[5][23]  ( .D(n3210), .CP(clk), .Q(\gpr[5][23] ), .QN(n5464) );
  FD1 \gpr_reg[5][21]  ( .D(n3208), .CP(clk), .Q(\gpr[5][21] ), .QN(n5420) );
  FD1 \gpr_reg[5][20]  ( .D(n3207), .CP(clk), .Q(\gpr[5][20] ), .QN(n5394) );
  FD1 \gpr_reg[5][19]  ( .D(n3206), .CP(clk), .Q(\gpr[5][19] ), .QN(n5368) );
  FD1 \gpr_reg[5][17]  ( .D(n3204), .CP(clk), .Q(\gpr[5][17] ), .QN(n5321) );
  FD1 \gpr_reg[5][16]  ( .D(n3203), .CP(clk), .Q(\gpr[5][16] ), .QN(n5302) );
  FD1 \gpr_reg[5][15]  ( .D(n3202), .CP(clk), .Q(\gpr[5][15] ), .QN(n5275) );
  FD1 \gpr_reg[5][14]  ( .D(n3201), .CP(clk), .Q(\gpr[5][14] ), .QN(n5249) );
  FD1 \gpr_reg[5][13]  ( .D(n3200), .CP(clk), .Q(\gpr[5][13] ), .QN(n5222) );
  FD1 \gpr_reg[5][10]  ( .D(n3197), .CP(clk), .Q(\gpr[5][10] ), .QN(n5152) );
  FD1 \gpr_reg[5][9]  ( .D(n3196), .CP(clk), .Q(\gpr[5][9] ), .QN(n5123) );
  FD1 \gpr_reg[5][8]  ( .D(n3195), .CP(clk), .Q(\gpr[5][8] ), .QN(n5096) );
  FD1 \gpr_reg[5][7]  ( .D(n3194), .CP(clk), .Q(\gpr[5][7] ), .QN(n5069) );
  FD1 \gpr_reg[5][6]  ( .D(n3193), .CP(clk), .Q(\gpr[5][6] ), .QN(n5044) );
  FD1 \gpr_reg[5][5]  ( .D(n3192), .CP(clk), .Q(\gpr[5][5] ), .QN(n5016) );
  FD1 \gpr_reg[5][3]  ( .D(n3190), .CP(clk), .Q(\gpr[5][3] ), .QN(n4971) );
  FD1 \gpr_reg[5][2]  ( .D(n3189), .CP(clk), .Q(\gpr[5][2] ), .QN(n4946) );
  FD1 \gpr_reg[6][31]  ( .D(n3186), .CP(clk), .Q(\gpr[6][31] ), .QN(n5665) );
  FD1 \gpr_reg[6][30]  ( .D(n3185), .CP(clk), .Q(\gpr[6][30] ), .QN(n5640) );
  FD1 \gpr_reg[6][29]  ( .D(n3184), .CP(clk), .Q(\gpr[6][29] ), .QN(n5612) );
  FD1 \gpr_reg[6][28]  ( .D(n3183), .CP(clk), .Q(\gpr[6][28] ), .QN(n5589) );
  FD1 \gpr_reg[6][26]  ( .D(n3181), .CP(clk), .Q(\gpr[6][26] ), .QN(n5538) );
  FD1 \gpr_reg[6][25]  ( .D(n3180), .CP(clk), .Q(\gpr[6][25] ), .QN(n5501) );
  FD1 \gpr_reg[6][24]  ( .D(n3179), .CP(clk), .Q(\gpr[6][24] ), .QN(n5490) );
  FD1 \gpr_reg[6][23]  ( .D(n3178), .CP(clk), .Q(\gpr[6][23] ), .QN(n5463) );
  FD1 \gpr_reg[6][21]  ( .D(n3176), .CP(clk), .Q(\gpr[6][21] ), .QN(n5419) );
  FD1 \gpr_reg[6][20]  ( .D(n3175), .CP(clk), .Q(\gpr[6][20] ), .QN(n5393) );
  FD1 \gpr_reg[6][19]  ( .D(n3174), .CP(clk), .Q(\gpr[6][19] ), .QN(n5367) );
  FD1 \gpr_reg[6][18]  ( .D(n3173), .CP(clk), .Q(\gpr[6][18] ), .QN(n310) );
  FD1 \gpr_reg[6][17]  ( .D(n3172), .CP(clk), .Q(\gpr[6][17] ), .QN(n5320) );
  FD1 \gpr_reg[6][16]  ( .D(n3171), .CP(clk), .Q(\gpr[6][16] ), .QN(n5301) );
  FD1 \gpr_reg[6][15]  ( .D(n3170), .CP(clk), .Q(\gpr[6][15] ), .QN(n5274) );
  FD1 \gpr_reg[6][14]  ( .D(n3169), .CP(clk), .Q(\gpr[6][14] ), .QN(n5248) );
  FD1 \gpr_reg[6][13]  ( .D(n3168), .CP(clk), .Q(\gpr[6][13] ), .QN(n5221) );
  FD1 \gpr_reg[6][10]  ( .D(n3165), .CP(clk), .Q(\gpr[6][10] ), .QN(n5151) );
  FD1 \gpr_reg[6][9]  ( .D(n3164), .CP(clk), .Q(\gpr[6][9] ), .QN(n5122) );
  FD1 \gpr_reg[6][8]  ( .D(n3163), .CP(clk), .Q(\gpr[6][8] ), .QN(n5095) );
  FD1 \gpr_reg[6][7]  ( .D(n3162), .CP(clk), .Q(\gpr[6][7] ), .QN(n5068) );
  FD1 \gpr_reg[6][6]  ( .D(n3161), .CP(clk), .Q(\gpr[6][6] ), .QN(n5043) );
  FD1 \gpr_reg[6][5]  ( .D(n3160), .CP(clk), .Q(\gpr[6][5] ), .QN(n5015) );
  FD1 \gpr_reg[6][3]  ( .D(n3158), .CP(clk), .Q(\gpr[6][3] ), .QN(n4970) );
  FD1 \gpr_reg[6][2]  ( .D(n3157), .CP(clk), .Q(\gpr[6][2] ), .QN(n4945) );
  FD1 \gpr_reg[6][1]  ( .D(n3156), .CP(clk), .Q(\gpr[6][1] ), .QN(n4919) );
  FD1 \gpr_reg[6][0]  ( .D(n3155), .CP(clk), .Q(\gpr[6][0] ), .QN(n4901) );
  FD1 \gpr_reg[7][31]  ( .D(n3154), .CP(clk), .Q(\gpr[7][31] ), .QN(n5664) );
  FD1 \gpr_reg[7][30]  ( .D(n3153), .CP(clk), .Q(\gpr[7][30] ), .QN(n5639) );
  FD1 \gpr_reg[7][29]  ( .D(n3152), .CP(clk), .Q(\gpr[7][29] ), .QN(n5611) );
  FD1 \gpr_reg[7][28]  ( .D(n3151), .CP(clk), .Q(\gpr[7][28] ), .QN(n5588) );
  FD1 \gpr_reg[7][27]  ( .D(n3150), .CP(clk), .Q(\gpr[7][27] ), .QN(n5565) );
  FD1 \gpr_reg[7][26]  ( .D(n3149), .CP(clk), .Q(\gpr[7][26] ), .QN(n5537) );
  FD1 \gpr_reg[7][25]  ( .D(n3148), .CP(clk), .Q(\gpr[7][25] ), .QN(n5500) );
  FD1 \gpr_reg[7][24]  ( .D(n3147), .CP(clk), .Q(\gpr[7][24] ), .QN(n5489) );
  FD1 \gpr_reg[7][23]  ( .D(n3146), .CP(clk), .Q(\gpr[7][23] ), .QN(n5462) );
  FD1 \gpr_reg[7][21]  ( .D(n3144), .CP(clk), .Q(\gpr[7][21] ), .QN(n5418) );
  FD1 \gpr_reg[7][20]  ( .D(n3143), .CP(clk), .Q(\gpr[7][20] ), .QN(n5392) );
  FD1 \gpr_reg[7][19]  ( .D(n3142), .CP(clk), .Q(\gpr[7][19] ), .QN(n5366) );
  FD1 \gpr_reg[7][18]  ( .D(n3141), .CP(clk), .Q(\gpr[7][18] ), .QN(n5345) );
  FD1 \gpr_reg[7][17]  ( .D(n3140), .CP(clk), .Q(\gpr[7][17] ), .QN(n5319) );
  FD1 \gpr_reg[7][16]  ( .D(n3139), .CP(clk), .Q(\gpr[7][16] ), .QN(n5300) );
  FD1 \gpr_reg[7][15]  ( .D(n3138), .CP(clk), .Q(\gpr[7][15] ), .QN(n5273) );
  FD1 \gpr_reg[7][14]  ( .D(n3137), .CP(clk), .Q(\gpr[7][14] ), .QN(n5247) );
  FD1 \gpr_reg[7][13]  ( .D(n3136), .CP(clk), .Q(\gpr[7][13] ), .QN(n5220) );
  FD1 \gpr_reg[7][11]  ( .D(n3134), .CP(clk), .Q(\gpr[7][11] ), .QN(n5177) );
  FD1 \gpr_reg[7][10]  ( .D(n3133), .CP(clk), .Q(\gpr[7][10] ), .QN(n5150) );
  FD1 \gpr_reg[7][9]  ( .D(n3132), .CP(clk), .Q(\gpr[7][9] ), .QN(n5121) );
  FD1 \gpr_reg[7][8]  ( .D(n3131), .CP(clk), .Q(\gpr[7][8] ), .QN(n5094) );
  FD1 \gpr_reg[7][7]  ( .D(n3130), .CP(clk), .Q(\gpr[7][7] ), .QN(n5067) );
  FD1 \gpr_reg[7][6]  ( .D(n3129), .CP(clk), .Q(\gpr[7][6] ), .QN(n5042) );
  FD1 \gpr_reg[7][5]  ( .D(n3128), .CP(clk), .Q(\gpr[7][5] ), .QN(n5014) );
  FD1 \gpr_reg[7][3]  ( .D(n3126), .CP(clk), .Q(\gpr[7][3] ), .QN(n4969) );
  FD1 \gpr_reg[7][2]  ( .D(n3125), .CP(clk), .Q(\gpr[7][2] ), .QN(n4944) );
  FD1 \gpr_reg[7][1]  ( .D(n3124), .CP(clk), .Q(\gpr[7][1] ), .QN(n4837) );
  FD1 \gpr_reg[7][0]  ( .D(n3123), .CP(clk), .Q(\gpr[7][0] ), .QN(n4900) );
  FD1 \gpr_reg[8][31]  ( .D(n3122), .CP(clk), .Q(\gpr[8][31] ), .QN(n5657) );
  FD1 \gpr_reg[8][30]  ( .D(n3121), .CP(clk), .Q(\gpr[8][30] ), .QN(n5632) );
  FD1 \gpr_reg[8][29]  ( .D(n3120), .CP(clk), .Q(\gpr[8][29] ), .QN(n5604) );
  FD1 \gpr_reg[8][28]  ( .D(n3119), .CP(clk), .Q(\gpr[8][28] ), .QN(n5581) );
  FD1 \gpr_reg[8][27]  ( .D(n3118), .CP(clk), .Q(\gpr[8][27] ), .QN(n5557) );
  FD1 \gpr_reg[8][26]  ( .D(n3117), .CP(clk), .Q(\gpr[8][26] ), .QN(n5530) );
  FD1 \gpr_reg[8][25]  ( .D(n3116), .CP(clk), .Q(\gpr[8][25] ), .QN(n315) );
  FD1 \gpr_reg[8][24]  ( .D(n3115), .CP(clk), .Q(\gpr[8][24] ), .QN(n5482) );
  FD1 \gpr_reg[8][23]  ( .D(n3114), .CP(clk), .Q(\gpr[8][23] ), .QN(n5455) );
  FD1 \gpr_reg[8][22]  ( .D(n3113), .CP(clk), .Q(\gpr[8][22] ), .QN(n5438) );
  FD1 \gpr_reg[8][21]  ( .D(n3112), .CP(clk), .Q(\gpr[8][21] ), .QN(n5411) );
  FD1 \gpr_reg[8][20]  ( .D(n3111), .CP(clk), .Q(\gpr[8][20] ), .QN(n5724) );
  FD1 \gpr_reg[8][19]  ( .D(n3110), .CP(clk), .Q(\gpr[8][19] ), .QN(n5359) );
  FD1 \gpr_reg[8][18]  ( .D(n3109), .CP(clk), .Q(\gpr[8][18] ), .QN(n5341) );
  FD1 \gpr_reg[8][17]  ( .D(n3108), .CP(clk), .Q(\gpr[8][17] ), .QN(n5315) );
  FD1 \gpr_reg[8][16]  ( .D(n3107), .CP(clk), .Q(\gpr[8][16] ), .QN(n5293) );
  FD1 \gpr_reg[8][15]  ( .D(n3106), .CP(clk), .Q(\gpr[8][15] ), .QN(n5266) );
  FD1 \gpr_reg[8][14]  ( .D(n3105), .CP(clk), .Q(\gpr[8][14] ), .QN(n5240) );
  FD1 \gpr_reg[8][13]  ( .D(n3104), .CP(clk), .Q(\gpr[8][13] ), .QN(n5213) );
  FD1 \gpr_reg[8][12]  ( .D(n3103), .CP(clk), .Q(\gpr[8][12] ), .QN(n5193) );
  FD1 \gpr_reg[8][11]  ( .D(n3102), .CP(clk), .Q(\gpr[8][11] ), .QN(n5169) );
  FD1 \gpr_reg[8][10]  ( .D(n3101), .CP(clk), .Q(\gpr[8][10] ), .QN(n5143) );
  FD1 \gpr_reg[8][9]  ( .D(n3100), .CP(clk), .Q(\gpr[8][9] ), .QN(n5114) );
  FD1 \gpr_reg[8][8]  ( .D(n3099), .CP(clk), .Q(\gpr[8][8] ), .QN(n5087) );
  FD1 \gpr_reg[8][7]  ( .D(n3098), .CP(clk), .Q(\gpr[8][7] ), .QN(n5060) );
  FD1 \gpr_reg[8][6]  ( .D(n3097), .CP(clk), .Q(\gpr[8][6] ), .QN(n5035) );
  FD1 \gpr_reg[8][5]  ( .D(n3096), .CP(clk), .Q(\gpr[8][5] ), .QN(n5007) );
  FD1 \gpr_reg[8][4]  ( .D(n3095), .CP(clk), .Q(\gpr[8][4] ), .QN(n4989) );
  FD1 \gpr_reg[8][3]  ( .D(n3094), .CP(clk), .Q(\gpr[8][3] ), .QN(n4962) );
  FD1 \gpr_reg[8][2]  ( .D(n3093), .CP(clk), .Q(\gpr[8][2] ), .QN(n4938) );
  FD1 \gpr_reg[8][0]  ( .D(n3091), .CP(clk), .Q(\gpr[8][0] ), .QN(n4904) );
  FD1 \gpr_reg[9][31]  ( .D(n3090), .CP(clk), .Q(\gpr[9][31] ), .QN(n5659) );
  FD1 \gpr_reg[9][30]  ( .D(n3089), .CP(clk), .Q(\gpr[9][30] ), .QN(n5634) );
  FD1 \gpr_reg[9][29]  ( .D(n3088), .CP(clk), .Q(\gpr[9][29] ), .QN(n5606) );
  FD1 \gpr_reg[9][28]  ( .D(n3087), .CP(clk), .Q(\gpr[9][28] ), .QN(n5583) );
  FD1 \gpr_reg[9][27]  ( .D(n3086), .CP(clk), .Q(\gpr[9][27] ), .QN(n5559) );
  FD1 \gpr_reg[9][26]  ( .D(n3085), .CP(clk), .Q(\gpr[9][26] ), .QN(n5532) );
  FD1 \gpr_reg[9][25]  ( .D(n3084), .CP(clk), .Q(\gpr[9][25] ), .QN(n5505) );
  FD1 \gpr_reg[9][24]  ( .D(n3083), .CP(clk), .Q(\gpr[9][24] ), .QN(n5484) );
  FD1 \gpr_reg[9][23]  ( .D(n3082), .CP(clk), .Q(\gpr[9][23] ), .QN(n5457) );
  FD1 \gpr_reg[9][21]  ( .D(n3080), .CP(clk), .Q(\gpr[9][21] ), .QN(n5413) );
  FD1 \gpr_reg[9][20]  ( .D(n3079), .CP(clk), .Q(\gpr[9][20] ), .QN(n5387) );
  FD1 \gpr_reg[9][19]  ( .D(n3078), .CP(clk), .Q(\gpr[9][19] ), .QN(n5361) );
  FD1 \gpr_reg[9][18]  ( .D(n3077), .CP(clk), .Q(\gpr[9][18] ), .QN(n308) );
  FD1 \gpr_reg[9][17]  ( .D(n3076), .CP(clk), .Q(\gpr[9][17] ), .QN(n5317) );
  FD1 \gpr_reg[9][16]  ( .D(n3075), .CP(clk), .Q(\gpr[9][16] ), .QN(n5295) );
  FD1 \gpr_reg[9][15]  ( .D(n3074), .CP(clk), .Q(\gpr[9][15] ), .QN(n5268) );
  FD1 \gpr_reg[9][14]  ( .D(n3073), .CP(clk), .Q(\gpr[9][14] ), .QN(n5242) );
  FD1 \gpr_reg[9][13]  ( .D(n3072), .CP(clk), .Q(\gpr[9][13] ), .QN(n5215) );
  FD1 \gpr_reg[9][11]  ( .D(n3070), .CP(clk), .Q(\gpr[9][11] ), .QN(n5171) );
  FD1 \gpr_reg[9][10]  ( .D(n3069), .CP(clk), .Q(\gpr[9][10] ), .QN(n5145) );
  FD1 \gpr_reg[9][9]  ( .D(n3068), .CP(clk), .Q(\gpr[9][9] ), .QN(n5116) );
  FD1 \gpr_reg[9][8]  ( .D(n3067), .CP(clk), .Q(\gpr[9][8] ), .QN(n5089) );
  FD1 \gpr_reg[9][7]  ( .D(n3066), .CP(clk), .Q(\gpr[9][7] ), .QN(n5062) );
  FD1 \gpr_reg[9][6]  ( .D(n3065), .CP(clk), .Q(\gpr[9][6] ), .QN(n5037) );
  FD1 \gpr_reg[9][5]  ( .D(n3064), .CP(clk), .Q(\gpr[9][5] ), .QN(n5009) );
  FD1 \gpr_reg[9][3]  ( .D(n3062), .CP(clk), .Q(\gpr[9][3] ), .QN(n4964) );
  FD1 \gpr_reg[9][2]  ( .D(n3061), .CP(clk), .Q(\gpr[9][2] ), .QN(n4940) );
  FD1 \gpr_reg[9][1]  ( .D(n3060), .CP(clk), .Q(\gpr[9][1] ), .QN(n4918) );
  FD1 \gpr_reg[9][0]  ( .D(n3059), .CP(clk), .Q(\gpr[9][0] ), .QN(n4906) );
  FD1 \gpr_reg[10][31]  ( .D(n3058), .CP(clk), .Q(\gpr[10][31] ), .QN(n5660)
         );
  FD1 \gpr_reg[10][30]  ( .D(n3057), .CP(clk), .Q(\gpr[10][30] ), .QN(n5636)
         );
  FD1 \gpr_reg[10][29]  ( .D(n3056), .CP(clk), .Q(\gpr[10][29] ), .QN(n5607)
         );
  FD1 \gpr_reg[10][28]  ( .D(n3055), .CP(clk), .Q(\gpr[10][28] ), .QN(n5584)
         );
  FD1 \gpr_reg[10][27]  ( .D(n3054), .CP(clk), .Q(\gpr[10][27] ), .QN(n5561)
         );
  FD1 \gpr_reg[10][26]  ( .D(n3053), .CP(clk), .Q(\gpr[10][26] ), .QN(n5534)
         );
  FD1 \gpr_reg[10][25]  ( .D(n3052), .CP(clk), .Q(\gpr[10][25] ), .QN(n4799)
         );
  FD1 \gpr_reg[10][24]  ( .D(n3051), .CP(clk), .Q(\gpr[10][24] ), .QN(n5485)
         );
  FD1 \gpr_reg[10][23]  ( .D(n3050), .CP(clk), .Q(\gpr[10][23] ), .QN(n5458)
         );
  FD1 \gpr_reg[10][22]  ( .D(n3049), .CP(clk), .Q(\gpr[10][22] ), .QN(n5439)
         );
  FD1 \gpr_reg[10][21]  ( .D(n3048), .CP(clk), .Q(\gpr[10][21] ), .QN(n5414)
         );
  FD1 \gpr_reg[10][20]  ( .D(n3047), .CP(clk), .Q(\gpr[10][20] ), .QN(n5388)
         );
  FD1 \gpr_reg[10][19]  ( .D(n3046), .CP(clk), .Q(\gpr[10][19] ), .QN(n5362)
         );
  FD1 \gpr_reg[10][18]  ( .D(n3045), .CP(clk), .Q(\gpr[10][18] ), .QN(n309) );
  FD1 \gpr_reg[10][17]  ( .D(n3044), .CP(clk), .Q(\gpr[10][17] ), .QN(n4839)
         );
  FD1 \gpr_reg[10][16]  ( .D(n3043), .CP(clk), .Q(\gpr[10][16] ), .QN(n5296)
         );
  FD1 \gpr_reg[10][15]  ( .D(n3042), .CP(clk), .Q(\gpr[10][15] ), .QN(n5269)
         );
  FD1 \gpr_reg[10][14]  ( .D(n3041), .CP(clk), .Q(\gpr[10][14] ), .QN(n5243)
         );
  FD1 \gpr_reg[10][13]  ( .D(n3040), .CP(clk), .Q(\gpr[10][13] ), .QN(n5216)
         );
  FD1 \gpr_reg[10][12]  ( .D(n3039), .CP(clk), .Q(\gpr[10][12] ), .QN(n5194)
         );
  FD1 \gpr_reg[10][11]  ( .D(n3038), .CP(clk), .Q(\gpr[10][11] ), .QN(n5173)
         );
  FD1 \gpr_reg[10][10]  ( .D(n3037), .CP(clk), .Q(\gpr[10][10] ), .QN(n5147)
         );
  FD1 \gpr_reg[10][9]  ( .D(n3036), .CP(clk), .Q(\gpr[10][9] ), .QN(n5117) );
  FD1 \gpr_reg[10][8]  ( .D(n3035), .CP(clk), .Q(\gpr[10][8] ), .QN(n5090) );
  FD1 \gpr_reg[10][7]  ( .D(n3034), .CP(clk), .Q(\gpr[10][7] ), .QN(n5063) );
  FD1 \gpr_reg[10][6]  ( .D(n3033), .CP(clk), .Q(\gpr[10][6] ), .QN(n5039) );
  FD1 \gpr_reg[10][5]  ( .D(n3032), .CP(clk), .Q(\gpr[10][5] ), .QN(n5010) );
  FD1 \gpr_reg[10][4]  ( .D(n3031), .CP(clk), .Q(\gpr[10][4] ), .QN(n4990) );
  FD1 \gpr_reg[10][3]  ( .D(n3030), .CP(clk), .Q(\gpr[10][3] ), .QN(n4965) );
  FD1 \gpr_reg[10][2]  ( .D(n3029), .CP(clk), .Q(\gpr[10][2] ), .QN(n4941) );
  FD1 \gpr_reg[10][1]  ( .D(n3028), .CP(clk), .Q(\gpr[10][1] ), .QN(n4838) );
  FD1 \gpr_reg[10][0]  ( .D(n3027), .CP(clk), .Q(\gpr[10][0] ), .QN(n298) );
  FD1 \gpr_reg[11][31]  ( .D(n3026), .CP(clk), .Q(\gpr[11][31] ), .QN(n5658)
         );
  FD1 \gpr_reg[11][30]  ( .D(n3025), .CP(clk), .Q(\gpr[11][30] ), .QN(n5633)
         );
  FD1 \gpr_reg[11][29]  ( .D(n3024), .CP(clk), .Q(\gpr[11][29] ), .QN(n5605)
         );
  FD1 \gpr_reg[11][28]  ( .D(n3023), .CP(clk), .Q(\gpr[11][28] ), .QN(n5582)
         );
  FD1 \gpr_reg[11][27]  ( .D(n3022), .CP(clk), .Q(\gpr[11][27] ), .QN(n5558)
         );
  FD1 \gpr_reg[11][26]  ( .D(n3021), .CP(clk), .Q(\gpr[11][26] ), .QN(n5531)
         );
  FD1 \gpr_reg[11][25]  ( .D(n3020), .CP(clk), .Q(\gpr[11][25] ), .QN(n5504)
         );
  FD1 \gpr_reg[11][24]  ( .D(n3019), .CP(clk), .Q(\gpr[11][24] ), .QN(n5483)
         );
  FD1 \gpr_reg[11][23]  ( .D(n3018), .CP(clk), .Q(\gpr[11][23] ), .QN(n5456)
         );
  FD1 \gpr_reg[11][21]  ( .D(n3016), .CP(clk), .Q(\gpr[11][21] ), .QN(n5412)
         );
  FD1 \gpr_reg[11][20]  ( .D(n3015), .CP(clk), .Q(\gpr[11][20] ), .QN(n5386)
         );
  FD1 \gpr_reg[11][19]  ( .D(n3014), .CP(clk), .Q(\gpr[11][19] ), .QN(n5360)
         );
  FD1 \gpr_reg[11][18]  ( .D(n3013), .CP(clk), .Q(\gpr[11][18] ), .QN(n307) );
  FD1 \gpr_reg[11][17]  ( .D(n3012), .CP(clk), .Q(\gpr[11][17] ), .QN(n5316)
         );
  FD1 \gpr_reg[11][16]  ( .D(n3011), .CP(clk), .Q(\gpr[11][16] ), .QN(n5294)
         );
  FD1 \gpr_reg[11][15]  ( .D(n3010), .CP(clk), .Q(\gpr[11][15] ), .QN(n5267)
         );
  FD1 \gpr_reg[11][14]  ( .D(n3009), .CP(clk), .Q(\gpr[11][14] ), .QN(n5241)
         );
  FD1 \gpr_reg[11][13]  ( .D(n3008), .CP(clk), .Q(\gpr[11][13] ), .QN(n5214)
         );
  FD1 \gpr_reg[11][11]  ( .D(n3006), .CP(clk), .Q(\gpr[11][11] ), .QN(n5170)
         );
  FD1 \gpr_reg[11][10]  ( .D(n3005), .CP(clk), .Q(\gpr[11][10] ), .QN(n5144)
         );
  FD1 \gpr_reg[11][9]  ( .D(n3004), .CP(clk), .Q(\gpr[11][9] ), .QN(n5115) );
  FD1 \gpr_reg[11][8]  ( .D(n3003), .CP(clk), .Q(\gpr[11][8] ), .QN(n5088) );
  FD1 \gpr_reg[11][7]  ( .D(n3002), .CP(clk), .Q(\gpr[11][7] ), .QN(n5061) );
  FD1 \gpr_reg[11][6]  ( .D(n3001), .CP(clk), .Q(\gpr[11][6] ), .QN(n5036) );
  FD1 \gpr_reg[11][5]  ( .D(n3000), .CP(clk), .Q(\gpr[11][5] ), .QN(n5008) );
  FD1 \gpr_reg[11][3]  ( .D(n2998), .CP(clk), .Q(\gpr[11][3] ), .QN(n4963) );
  FD1 \gpr_reg[11][2]  ( .D(n2997), .CP(clk), .Q(\gpr[11][2] ), .QN(n4939) );
  FD1 \gpr_reg[11][1]  ( .D(n2996), .CP(clk), .Q(\gpr[11][1] ), .QN(n4917) );
  FD1 \gpr_reg[11][0]  ( .D(n2995), .CP(clk), .Q(\gpr[11][0] ), .QN(n4905) );
  FD1 \gpr_reg[12][31]  ( .D(n2994), .CP(clk), .Q(\gpr[12][31] ), .QN(n5656)
         );
  FD1 \gpr_reg[12][30]  ( .D(n2993), .CP(clk), .Q(\gpr[12][30] ), .QN(n5631)
         );
  FD1 \gpr_reg[12][29]  ( .D(n2992), .CP(clk), .Q(\gpr[12][29] ), .QN(n5603)
         );
  FD1 \gpr_reg[12][28]  ( .D(n2991), .CP(clk), .Q(\gpr[12][28] ), .QN(n5580)
         );
  FD1 \gpr_reg[12][27]  ( .D(n2990), .CP(clk), .Q(\gpr[12][27] ), .QN(n5556)
         );
  FD1 \gpr_reg[12][25]  ( .D(n2988), .CP(clk), .Q(\gpr[12][25] ), .QN(n5503)
         );
  FD1 \gpr_reg[12][24]  ( .D(n2987), .CP(clk), .Q(\gpr[12][24] ), .QN(n5481)
         );
  FD1 \gpr_reg[12][23]  ( .D(n2986), .CP(clk), .Q(\gpr[12][23] ), .QN(n5454)
         );
  FD1 \gpr_reg[12][22]  ( .D(n2985), .CP(clk), .Q(\gpr[12][22] ), .QN(n5437)
         );
  FD1 \gpr_reg[12][21]  ( .D(n2984), .CP(clk), .Q(\gpr[12][21] ), .QN(n5410)
         );
  FD1 \gpr_reg[12][20]  ( .D(n2983), .CP(clk), .Q(\gpr[12][20] ), .QN(n5385)
         );
  FD1 \gpr_reg[12][19]  ( .D(n2982), .CP(clk), .Q(\gpr[12][19] ), .QN(n5358)
         );
  FD1 \gpr_reg[12][18]  ( .D(n2981), .CP(clk), .Q(\gpr[12][18] ), .QN(n306) );
  FD1 \gpr_reg[12][17]  ( .D(n2980), .CP(clk), .Q(\gpr[12][17] ), .QN(n5314)
         );
  FD1 \gpr_reg[12][16]  ( .D(n2979), .CP(clk), .Q(\gpr[12][16] ), .QN(n5292)
         );
  FD1 \gpr_reg[12][15]  ( .D(n2978), .CP(clk), .Q(\gpr[12][15] ), .QN(n5265)
         );
  FD1 \gpr_reg[12][14]  ( .D(n2977), .CP(clk), .Q(\gpr[12][14] ), .QN(n5239)
         );
  FD1 \gpr_reg[12][13]  ( .D(n2976), .CP(clk), .Q(\gpr[12][13] ), .QN(n5212)
         );
  FD1 \gpr_reg[12][12]  ( .D(n2975), .CP(clk), .Q(\gpr[12][12] ), .QN(n5192)
         );
  FD1 \gpr_reg[12][11]  ( .D(n2974), .CP(clk), .Q(\gpr[12][11] ), .QN(n5168)
         );
  FD1 \gpr_reg[12][10]  ( .D(n2973), .CP(clk), .Q(\gpr[12][10] ), .QN(n5142)
         );
  FD1 \gpr_reg[12][9]  ( .D(n2972), .CP(clk), .Q(\gpr[12][9] ), .QN(n5113) );
  FD1 \gpr_reg[12][8]  ( .D(n2971), .CP(clk), .Q(\gpr[12][8] ), .QN(n5086) );
  FD1 \gpr_reg[12][7]  ( .D(n2970), .CP(clk), .Q(\gpr[12][7] ), .QN(n5059) );
  FD1 \gpr_reg[12][6]  ( .D(n2969), .CP(clk), .Q(\gpr[12][6] ), .QN(n5034) );
  FD1 \gpr_reg[12][5]  ( .D(n2968), .CP(clk), .Q(\gpr[12][5] ), .QN(n5006) );
  FD1 \gpr_reg[12][4]  ( .D(n2967), .CP(clk), .Q(\gpr[12][4] ), .QN(n4988) );
  FD1 \gpr_reg[12][3]  ( .D(n2966), .CP(clk), .Q(\gpr[12][3] ), .QN(n4961) );
  FD1 \gpr_reg[12][1]  ( .D(n2964), .CP(clk), .Q(\gpr[12][1] ), .QN(n4916) );
  FD1 \gpr_reg[12][0]  ( .D(n2963), .CP(clk), .Q(\gpr[12][0] ), .QN(n4903) );
  FD1 \gpr_reg[13][31]  ( .D(n2962), .CP(clk), .Q(\gpr[13][31] ), .QN(n4804)
         );
  FD1 \gpr_reg[13][30]  ( .D(n2961), .CP(clk), .Q(\gpr[13][30] ), .QN(n5629)
         );
  FD1 \gpr_reg[13][29]  ( .D(n2960), .CP(clk), .Q(\gpr[13][29] ), .QN(n4803)
         );
  FD1 \gpr_reg[13][28]  ( .D(n2959), .CP(clk), .Q(\gpr[13][28] ), .QN(n4802)
         );
  FD1 \gpr_reg[13][27]  ( .D(n2958), .CP(clk), .Q(\gpr[13][27] ), .QN(n4801)
         );
  FD1 \gpr_reg[13][26]  ( .D(n2957), .CP(clk), .Q(\gpr[13][26] ), .QN(n4800)
         );
  FD1 \gpr_reg[13][25]  ( .D(n2956), .CP(clk), .Q(\gpr[13][25] ), .QN(n4798)
         );
  FD1 \gpr_reg[13][24]  ( .D(n2955), .CP(clk), .Q(\gpr[13][24] ), .QN(n4769)
         );
  FD1 \gpr_reg[13][23]  ( .D(n2954), .CP(clk), .Q(\gpr[13][23] ), .QN(n4795)
         );
  FD1 \gpr_reg[13][22]  ( .D(n2953), .CP(clk), .Q(\gpr[13][22] ), .QN(n4794)
         );
  FD1 \gpr_reg[13][21]  ( .D(n2952), .CP(clk), .Q(\gpr[13][21] ), .QN(n4793)
         );
  FD1 \gpr_reg[13][20]  ( .D(n2951), .CP(clk), .Q(\gpr[13][20] ), .QN(n4768)
         );
  FD1 \gpr_reg[13][19]  ( .D(n2950), .CP(clk), .Q(\gpr[13][19] ), .QN(n4792)
         );
  FD1 \gpr_reg[13][18]  ( .D(n2949), .CP(clk), .Q(\gpr[13][18] ), .QN(n4791)
         );
  FD1 \gpr_reg[13][17]  ( .D(n2948), .CP(clk), .Q(\gpr[13][17] ), .QN(n4790)
         );
  FD1 \gpr_reg[13][16]  ( .D(n2947), .CP(clk), .Q(\gpr[13][16] ), .QN(n4767)
         );
  FD1 \gpr_reg[13][15]  ( .D(n2946), .CP(clk), .Q(\gpr[13][15] ), .QN(n4787)
         );
  FD1 \gpr_reg[13][14]  ( .D(n2945), .CP(clk), .Q(\gpr[13][14] ), .QN(n4766)
         );
  FD1 \gpr_reg[13][13]  ( .D(n2944), .CP(clk), .Q(\gpr[13][13] ), .QN(n4786)
         );
  FD1 \gpr_reg[13][12]  ( .D(n2943), .CP(clk), .Q(\gpr[13][12] ), .QN(n4785)
         );
  FD1 \gpr_reg[13][11]  ( .D(n2942), .CP(clk), .Q(\gpr[13][11] ), .QN(n4784)
         );
  FD1 \gpr_reg[13][10]  ( .D(n2941), .CP(clk), .Q(\gpr[13][10] ), .QN(n5140)
         );
  FD1 \gpr_reg[13][9]  ( .D(n2940), .CP(clk), .Q(\gpr[13][9] ), .QN(n4783) );
  FD1 \gpr_reg[13][8]  ( .D(n2939), .CP(clk), .Q(\gpr[13][8] ), .QN(n4765) );
  FD1 \gpr_reg[13][7]  ( .D(n2938), .CP(clk), .Q(\gpr[13][7] ), .QN(n4782) );
  FD1 \gpr_reg[13][6]  ( .D(n2937), .CP(clk), .Q(\gpr[13][6] ), .QN(n5032) );
  FD1 \gpr_reg[13][5]  ( .D(n2936), .CP(clk), .Q(\gpr[13][5] ), .QN(n4781) );
  FD1 \gpr_reg[13][3]  ( .D(n2934), .CP(clk), .Q(\gpr[13][3] ), .QN(n4780) );
  FD1 \gpr_reg[13][2]  ( .D(n2933), .CP(clk), .Q(\gpr[13][2] ), .QN(n4778) );
  FD1 \gpr_reg[13][1]  ( .D(n2932), .CP(clk), .Q(\gpr[13][1] ), .QN(n4911) );
  FD1 \gpr_reg[13][0]  ( .D(n2931), .CP(clk), .Q(\gpr[13][0] ), .QN(n4777) );
  FD1 \gpr_reg[14][31]  ( .D(n2930), .CP(clk), .Q(\gpr[14][31] ), .QN(n4826)
         );
  FD1 \gpr_reg[14][30]  ( .D(n2929), .CP(clk), .Q(\gpr[14][30] ), .QN(n5635)
         );
  FD1 \gpr_reg[14][29]  ( .D(n2928), .CP(clk), .Q(\gpr[14][29] ), .QN(n4825)
         );
  FD1 \gpr_reg[14][28]  ( .D(n2927), .CP(clk), .Q(\gpr[14][28] ), .QN(n4824)
         );
  FD1 \gpr_reg[14][27]  ( .D(n2926), .CP(clk), .Q(\gpr[14][27] ), .QN(n5560)
         );
  FD1 \gpr_reg[14][26]  ( .D(n2925), .CP(clk), .Q(\gpr[14][26] ), .QN(n5533)
         );
  FD1 \gpr_reg[14][25]  ( .D(n2924), .CP(clk), .Q(\gpr[14][25] ), .QN(n5506)
         );
  FD1 \gpr_reg[14][24]  ( .D(n2923), .CP(clk), .Q(\gpr[14][24] ), .QN(n4775)
         );
  FD1 \gpr_reg[14][23]  ( .D(n2922), .CP(clk), .Q(\gpr[14][23] ), .QN(n4823)
         );
  FD1 \gpr_reg[14][22]  ( .D(n2921), .CP(clk), .Q(\gpr[14][22] ), .QN(n4822)
         );
  FD1 \gpr_reg[14][21]  ( .D(n2920), .CP(clk), .Q(\gpr[14][21] ), .QN(n4821)
         );
  FD1 \gpr_reg[14][20]  ( .D(n2919), .CP(clk), .Q(\gpr[14][20] ), .QN(n4774)
         );
  FD1 \gpr_reg[14][19]  ( .D(n2918), .CP(clk), .Q(\gpr[14][19] ), .QN(n4820)
         );
  FD1 \gpr_reg[14][18]  ( .D(n2917), .CP(clk), .Q(\gpr[14][18] ), .QN(n5342)
         );
  FD1 \gpr_reg[14][16]  ( .D(n2915), .CP(clk), .Q(\gpr[14][16] ), .QN(n4773)
         );
  FD1 \gpr_reg[14][15]  ( .D(n2914), .CP(clk), .Q(\gpr[14][15] ), .QN(n4819)
         );
  FD1 \gpr_reg[14][14]  ( .D(n2913), .CP(clk), .Q(\gpr[14][14] ), .QN(n4772)
         );
  FD1 \gpr_reg[14][13]  ( .D(n2912), .CP(clk), .Q(\gpr[14][13] ), .QN(n4818)
         );
  FD1 \gpr_reg[14][12]  ( .D(n2911), .CP(clk), .Q(\gpr[14][12] ), .QN(n4817)
         );
  FD1 \gpr_reg[14][11]  ( .D(n2910), .CP(clk), .Q(\gpr[14][11] ), .QN(n5172)
         );
  FD1 \gpr_reg[14][10]  ( .D(n2909), .CP(clk), .Q(\gpr[14][10] ), .QN(n5146)
         );
  FD1 \gpr_reg[14][9]  ( .D(n2908), .CP(clk), .Q(\gpr[14][9] ), .QN(n4816) );
  FD1 \gpr_reg[14][8]  ( .D(n2907), .CP(clk), .Q(\gpr[14][8] ), .QN(n4771) );
  FD1 \gpr_reg[14][7]  ( .D(n2906), .CP(clk), .Q(\gpr[14][7] ), .QN(n4815) );
  FD1 \gpr_reg[14][6]  ( .D(n2905), .CP(clk), .Q(\gpr[14][6] ), .QN(n5038) );
  FD1 \gpr_reg[14][5]  ( .D(n2904), .CP(clk), .Q(\gpr[14][5] ), .QN(n4814) );
  FD1 \gpr_reg[14][3]  ( .D(n2902), .CP(clk), .Q(\gpr[14][3] ), .QN(n4813) );
  FD1 \gpr_reg[14][2]  ( .D(n2901), .CP(clk), .Q(\gpr[14][2] ), .QN(n4812) );
  FD1 \gpr_reg[14][0]  ( .D(n2899), .CP(clk), .Q(\gpr[14][0] ), .QN(n4907) );
  FD1 \gpr_reg[15][31]  ( .D(n2898), .CP(clk), .Q(\gpr[15][31] ), .QN(n5661)
         );
  FD1 \gpr_reg[15][30]  ( .D(n2897), .CP(clk), .Q(\gpr[15][30] ), .QN(n5630)
         );
  FD1 \gpr_reg[15][29]  ( .D(n2896), .CP(clk), .Q(\gpr[15][29] ), .QN(n5608)
         );
  FD1 \gpr_reg[15][28]  ( .D(n2895), .CP(clk), .Q(\gpr[15][28] ), .QN(n5585)
         );
  FD1 \gpr_reg[15][27]  ( .D(n2894), .CP(clk), .Q(\gpr[15][27] ), .QN(n5562)
         );
  FD1 \gpr_reg[15][26]  ( .D(n2893), .CP(clk), .Q(\gpr[15][26] ), .QN(n5535)
         );
  FD1 \gpr_reg[15][25]  ( .D(n2892), .CP(clk), .Q(\gpr[15][25] ), .QN(n5499)
         );
  FD1 \gpr_reg[15][24]  ( .D(n2891), .CP(clk), .Q(\gpr[15][24] ), .QN(n5486)
         );
  FD1 \gpr_reg[15][23]  ( .D(n2890), .CP(clk), .Q(\gpr[15][23] ), .QN(n5459)
         );
  FD1 \gpr_reg[15][22]  ( .D(n2889), .CP(clk), .Q(\gpr[15][22] ), .QN(n5440)
         );
  FD1 \gpr_reg[15][21]  ( .D(n2888), .CP(clk), .Q(\gpr[15][21] ), .QN(n5415)
         );
  FD1 \gpr_reg[15][20]  ( .D(n2887), .CP(clk), .Q(\gpr[15][20] ), .QN(n5389)
         );
  FD1 \gpr_reg[15][19]  ( .D(n2886), .CP(clk), .Q(\gpr[15][19] ), .QN(n5363)
         );
  FD1 \gpr_reg[15][18]  ( .D(n2885), .CP(clk), .Q(\gpr[15][18] ), .QN(n5343)
         );
  FD1 \gpr_reg[15][17]  ( .D(n2884), .CP(clk), .Q(\gpr[15][17] ), .QN(n5310)
         );
  FD1 \gpr_reg[15][16]  ( .D(n2883), .CP(clk), .Q(\gpr[15][16] ), .QN(n5297)
         );
  FD1 \gpr_reg[15][15]  ( .D(n2882), .CP(clk), .Q(\gpr[15][15] ), .QN(n5270)
         );
  FD1 \gpr_reg[15][14]  ( .D(n2881), .CP(clk), .Q(\gpr[15][14] ), .QN(n5244)
         );
  FD1 \gpr_reg[15][13]  ( .D(n2880), .CP(clk), .Q(\gpr[15][13] ), .QN(n5217)
         );
  FD1 \gpr_reg[15][12]  ( .D(n2879), .CP(clk), .Q(\gpr[15][12] ), .QN(n5195)
         );
  FD1 \gpr_reg[15][11]  ( .D(n2878), .CP(clk), .Q(\gpr[15][11] ), .QN(n5174)
         );
  FD1 \gpr_reg[15][10]  ( .D(n2877), .CP(clk), .Q(\gpr[15][10] ), .QN(n5141)
         );
  FD1 \gpr_reg[15][9]  ( .D(n2876), .CP(clk), .Q(\gpr[15][9] ), .QN(n5118) );
  FD1 \gpr_reg[15][8]  ( .D(n2875), .CP(clk), .Q(\gpr[15][8] ), .QN(n5091) );
  FD1 \gpr_reg[15][7]  ( .D(n2874), .CP(clk), .Q(\gpr[15][7] ), .QN(n5064) );
  FD1 \gpr_reg[15][6]  ( .D(n2873), .CP(clk), .Q(\gpr[15][6] ), .QN(n5033) );
  FD1 \gpr_reg[15][5]  ( .D(n2872), .CP(clk), .Q(\gpr[15][5] ), .QN(n5011) );
  FD1 \gpr_reg[15][3]  ( .D(n2870), .CP(clk), .Q(\gpr[15][3] ), .QN(n4966) );
  FD1 \gpr_reg[15][2]  ( .D(n2869), .CP(clk), .Q(\gpr[15][2] ), .QN(n4942) );
  FD1 \gpr_reg[15][1]  ( .D(n2868), .CP(clk), .Q(\gpr[15][1] ), .QN(n4912) );
  FD1 \gpr_reg[15][0]  ( .D(n2867), .CP(clk), .Q(\gpr[15][0] ), .QN(n4902) );
  FD1 \gpr_reg[16][31]  ( .D(n2866), .CP(clk), .Q(\gpr[16][31] ), .QN(n5648)
         );
  FD1 \gpr_reg[16][29]  ( .D(n2864), .CP(clk), .Q(\gpr[16][29] ), .QN(n5594)
         );
  FD1 \gpr_reg[16][28]  ( .D(n2863), .CP(clk), .Q(\gpr[16][28] ), .QN(n5575)
         );
  FD1 \gpr_reg[16][27]  ( .D(n2862), .CP(clk), .Q(\gpr[16][27] ), .QN(n5543)
         );
  FD1 \gpr_reg[16][26]  ( .D(n2861), .CP(clk), .Q(\gpr[16][26] ), .QN(n5524)
         );
  FD1 \gpr_reg[16][25]  ( .D(n2860), .CP(clk), .Q(\gpr[16][25] ), .QN(n5513)
         );
  FD1 \gpr_reg[16][24]  ( .D(n2859), .CP(clk), .Q(\gpr[16][24] ), .QN(n5479)
         );
  FD1 \gpr_reg[16][23]  ( .D(n2858), .CP(clk), .Q(\gpr[16][23] ), .QN(n5450)
         );
  FD1 \gpr_reg[16][22]  ( .D(n2857), .CP(clk), .Q(\gpr[16][22] ), .QN(n5428)
         );
  FD1 \gpr_reg[16][21]  ( .D(n2856), .CP(clk), .Q(\gpr[16][21] ), .QN(n5408)
         );
  FD1 \gpr_reg[16][20]  ( .D(n2855), .CP(clk), .Q(\gpr[16][20] ), .QN(n5379)
         );
  FD1 \gpr_reg[16][19]  ( .D(n2854), .CP(clk), .Q(\gpr[16][19] ), .QN(n5348)
         );
  FD1 \gpr_reg[16][18]  ( .D(n2853), .CP(clk), .Q(\gpr[16][18] ), .QN(n5339)
         );
  FD1 \gpr_reg[16][17]  ( .D(n2852), .CP(clk), .Q(\gpr[16][17] ), .QN(n5324)
         );
  FD1 \gpr_reg[16][16]  ( .D(n2851), .CP(clk), .Q(\gpr[16][16] ), .QN(n5290)
         );
  FD1 \gpr_reg[16][14]  ( .D(n2849), .CP(clk), .Q(\gpr[16][14] ), .QN(n5234)
         );
  FD1 \gpr_reg[16][13]  ( .D(n2848), .CP(clk), .Q(\gpr[16][13] ), .QN(n5207)
         );
  FD1 \gpr_reg[16][12]  ( .D(n2847), .CP(clk), .Q(\gpr[16][12] ), .QN(n5187)
         );
  FD1 \gpr_reg[16][11]  ( .D(n2846), .CP(clk), .Q(\gpr[16][11] ), .QN(n5157)
         );
  FD1 \gpr_reg[16][10]  ( .D(n2845), .CP(clk), .Q(\gpr[16][10] ), .QN(n5138)
         );
  FD1 \gpr_reg[16][9]  ( .D(n2844), .CP(clk), .Q(\gpr[16][9] ), .QN(n5108) );
  FD1 \gpr_reg[16][8]  ( .D(n2843), .CP(clk), .Q(\gpr[16][8] ), .QN(n5077) );
  FD1 \gpr_reg[16][7]  ( .D(n2842), .CP(clk), .Q(\gpr[16][7] ), .QN(n5057) );
  FD1 \gpr_reg[16][6]  ( .D(n2841), .CP(clk), .Q(\gpr[16][6] ), .QN(n301) );
  FD1 \gpr_reg[16][5]  ( .D(n2840), .CP(clk), .Q(\gpr[16][5] ), .QN(n4994) );
  FD1 \gpr_reg[16][4]  ( .D(n2839), .CP(clk), .Q(\gpr[16][4] ), .QN(n4984) );
  FD1 \gpr_reg[16][3]  ( .D(n2838), .CP(clk), .Q(\gpr[16][3] ), .QN(n4957) );
  FD1 \gpr_reg[16][2]  ( .D(n2837), .CP(clk), .Q(\gpr[16][2] ), .QN(n4936) );
  FD1 \gpr_reg[16][0]  ( .D(n2835), .CP(clk), .Q(\gpr[16][0] ), .QN(n4895) );
  FD1 \gpr_reg[17][31]  ( .D(n2834), .CP(clk), .Q(\gpr[17][31] ), .QN(n5646)
         );
  FD1 \gpr_reg[17][30]  ( .D(n2833), .CP(clk), .Q(\gpr[17][30] ), .QN(n5626)
         );
  FD1 \gpr_reg[17][29]  ( .D(n2832), .CP(clk), .Q(\gpr[17][29] ), .QN(n5597)
         );
  FD1 \gpr_reg[17][28]  ( .D(n2831), .CP(clk), .Q(\gpr[17][28] ), .QN(n5578)
         );
  FD1 \gpr_reg[17][27]  ( .D(n2830), .CP(clk), .Q(\gpr[17][27] ), .QN(n5544)
         );
  FD1 \gpr_reg[17][26]  ( .D(n2829), .CP(clk), .Q(\gpr[17][26] ), .QN(n5525)
         );
  FD1 \gpr_reg[17][25]  ( .D(n2828), .CP(clk), .Q(\gpr[17][25] ), .QN(n5515)
         );
  FD1 \gpr_reg[17][24]  ( .D(n2827), .CP(clk), .Q(\gpr[17][24] ), .QN(n5476)
         );
  FD1 \gpr_reg[17][23]  ( .D(n2826), .CP(clk), .Q(\gpr[17][23] ), .QN(n5452)
         );
  FD1 \gpr_reg[17][22]  ( .D(n2825), .CP(clk), .Q(\gpr[17][22] ), .QN(n5429)
         );
  FD1 \gpr_reg[17][21]  ( .D(n2824), .CP(clk), .Q(\gpr[17][21] ), .QN(n5405)
         );
  FD1 \gpr_reg[17][20]  ( .D(n2823), .CP(clk), .Q(\gpr[17][20] ), .QN(n5380)
         );
  FD1 \gpr_reg[17][19]  ( .D(n2822), .CP(clk), .Q(\gpr[17][19] ), .QN(n5351)
         );
  FD1 \gpr_reg[17][18]  ( .D(n2821), .CP(clk), .Q(\gpr[17][18] ), .QN(n5340)
         );
  FD1 \gpr_reg[17][17]  ( .D(n2820), .CP(clk), .Q(\gpr[17][17] ), .QN(n5326)
         );
  FD1 \gpr_reg[17][16]  ( .D(n2819), .CP(clk), .Q(\gpr[17][16] ), .QN(n5287)
         );
  FD1 \gpr_reg[17][15]  ( .D(n2818), .CP(clk), .Q(\gpr[17][15] ), .QN(n5255)
         );
  FD1 \gpr_reg[17][14]  ( .D(n2817), .CP(clk), .Q(\gpr[17][14] ), .QN(n5235)
         );
  FD1 \gpr_reg[17][13]  ( .D(n2816), .CP(clk), .Q(\gpr[17][13] ), .QN(n5210)
         );
  FD1 \gpr_reg[17][12]  ( .D(n2815), .CP(clk), .Q(\gpr[17][12] ), .QN(n5190)
         );
  FD1 \gpr_reg[17][11]  ( .D(n2814), .CP(clk), .Q(\gpr[17][11] ), .QN(n5160)
         );
  FD1 \gpr_reg[17][10]  ( .D(n2813), .CP(clk), .Q(\gpr[17][10] ), .QN(n5135)
         );
  FD1 \gpr_reg[17][9]  ( .D(n2812), .CP(clk), .Q(\gpr[17][9] ), .QN(n5109) );
  FD1 \gpr_reg[17][8]  ( .D(n2811), .CP(clk), .Q(\gpr[17][8] ), .QN(n5075) );
  FD1 \gpr_reg[17][7]  ( .D(n2810), .CP(clk), .Q(\gpr[17][7] ), .QN(n5055) );
  FD1 \gpr_reg[17][6]  ( .D(n2809), .CP(clk), .Q(\gpr[17][6] ), .QN(n5023) );
  FD1 \gpr_reg[17][5]  ( .D(n2808), .CP(clk), .Q(\gpr[17][5] ), .QN(n4997) );
  FD1 \gpr_reg[17][4]  ( .D(n2807), .CP(clk), .Q(\gpr[17][4] ), .QN(n4986) );
  FD1 \gpr_reg[17][3]  ( .D(n2806), .CP(clk), .Q(\gpr[17][3] ), .QN(n4959) );
  FD1 \gpr_reg[17][2]  ( .D(n2805), .CP(clk), .Q(\gpr[17][2] ), .QN(n4934) );
  FD1 \gpr_reg[17][0]  ( .D(n2803), .CP(clk), .Q(\gpr[17][0] ), .QN(n4897) );
  FD1 \gpr_reg[18][31]  ( .D(n2802), .CP(clk), .Q(\gpr[18][31] ), .QN(n5647)
         );
  FD1 \gpr_reg[18][30]  ( .D(n2801), .CP(clk), .Q(\gpr[18][30] ), .QN(n5627)
         );
  FD1 \gpr_reg[18][29]  ( .D(n2800), .CP(clk), .Q(\gpr[18][29] ), .QN(n5596)
         );
  FD1 \gpr_reg[18][28]  ( .D(n2799), .CP(clk), .Q(\gpr[18][28] ), .QN(n5577)
         );
  FD1 \gpr_reg[18][27]  ( .D(n2798), .CP(clk), .Q(\gpr[18][27] ), .QN(n5546)
         );
  FD1 \gpr_reg[18][26]  ( .D(n2797), .CP(clk), .Q(\gpr[18][26] ), .QN(n5527)
         );
  FD1 \gpr_reg[18][25]  ( .D(n2796), .CP(clk), .Q(\gpr[18][25] ), .QN(n4796)
         );
  FD1 \gpr_reg[18][24]  ( .D(n2795), .CP(clk), .Q(\gpr[18][24] ), .QN(n5478)
         );
  FD1 \gpr_reg[18][23]  ( .D(n2794), .CP(clk), .Q(\gpr[18][23] ), .QN(n5451)
         );
  FD1 \gpr_reg[18][22]  ( .D(n2793), .CP(clk), .Q(\gpr[18][22] ), .QN(n5427)
         );
  FD1 \gpr_reg[18][21]  ( .D(n2792), .CP(clk), .Q(\gpr[18][21] ), .QN(n5407)
         );
  FD1 \gpr_reg[18][20]  ( .D(n2791), .CP(clk), .Q(\gpr[18][20] ), .QN(n5382)
         );
  FD1 \gpr_reg[18][19]  ( .D(n2790), .CP(clk), .Q(\gpr[18][19] ), .QN(n5350)
         );
  FD1 \gpr_reg[18][18]  ( .D(n2789), .CP(clk), .Q(\gpr[18][18] ), .QN(n5338)
         );
  FD1 \gpr_reg[18][17]  ( .D(n2788), .CP(clk), .Q(\gpr[18][17] ), .QN(n4788)
         );
  FD1 \gpr_reg[18][16]  ( .D(n2787), .CP(clk), .Q(\gpr[18][16] ), .QN(n5289)
         );
  FD1 \gpr_reg[18][15]  ( .D(n2786), .CP(clk), .Q(\gpr[18][15] ), .QN(n5256)
         );
  FD1 \gpr_reg[18][14]  ( .D(n2785), .CP(clk), .Q(\gpr[18][14] ), .QN(n5237)
         );
  FD1 \gpr_reg[18][13]  ( .D(n2784), .CP(clk), .Q(\gpr[18][13] ), .QN(n5209)
         );
  FD1 \gpr_reg[18][12]  ( .D(n2783), .CP(clk), .Q(\gpr[18][12] ), .QN(n5189)
         );
  FD1 \gpr_reg[18][11]  ( .D(n2782), .CP(clk), .Q(\gpr[18][11] ), .QN(n5159)
         );
  FD1 \gpr_reg[18][10]  ( .D(n2781), .CP(clk), .Q(\gpr[18][10] ), .QN(n5137)
         );
  FD1 \gpr_reg[18][9]  ( .D(n2780), .CP(clk), .Q(\gpr[18][9] ), .QN(n5110) );
  FD1 \gpr_reg[18][8]  ( .D(n2779), .CP(clk), .Q(\gpr[18][8] ), .QN(n5076) );
  FD1 \gpr_reg[18][7]  ( .D(n2778), .CP(clk), .Q(\gpr[18][7] ), .QN(n5056) );
  FD1 \gpr_reg[18][6]  ( .D(n2777), .CP(clk), .Q(\gpr[18][6] ), .QN(n5022) );
  FD1 \gpr_reg[18][5]  ( .D(n2776), .CP(clk), .Q(\gpr[18][5] ), .QN(n4996) );
  FD1 \gpr_reg[18][4]  ( .D(n2775), .CP(clk), .Q(\gpr[18][4] ), .QN(n4985) );
  FD1 \gpr_reg[18][3]  ( .D(n2774), .CP(clk), .Q(\gpr[18][3] ), .QN(n299) );
  FD1 \gpr_reg[18][2]  ( .D(n2773), .CP(clk), .Q(\gpr[18][2] ), .QN(n4935) );
  FD1 \gpr_reg[18][1]  ( .D(n2772), .CP(clk), .Q(\gpr[18][1] ), .QN(n4836) );
  FD1 \gpr_reg[18][0]  ( .D(n2771), .CP(clk), .Q(\gpr[18][0] ), .QN(n4892) );
  FD1 \gpr_reg[19][31]  ( .D(n2770), .CP(clk), .Q(\gpr[19][31] ), .QN(n5645)
         );
  FD1 \gpr_reg[19][30]  ( .D(n2769), .CP(clk), .Q(\gpr[19][30] ), .QN(n5625)
         );
  FD1 \gpr_reg[19][29]  ( .D(n2768), .CP(clk), .Q(\gpr[19][29] ), .QN(n5595)
         );
  FD1 \gpr_reg[19][28]  ( .D(n2767), .CP(clk), .Q(\gpr[19][28] ), .QN(n5579)
         );
  FD1 \gpr_reg[19][27]  ( .D(n2766), .CP(clk), .Q(\gpr[19][27] ), .QN(n5547)
         );
  FD1 \gpr_reg[19][26]  ( .D(n2765), .CP(clk), .Q(\gpr[19][26] ), .QN(n5528)
         );
  FD1 \gpr_reg[19][25]  ( .D(n2764), .CP(clk), .Q(\gpr[19][25] ), .QN(n5514)
         );
  FD1 \gpr_reg[19][24]  ( .D(n2763), .CP(clk), .Q(\gpr[19][24] ), .QN(n5475)
         );
  FD1 \gpr_reg[19][23]  ( .D(n2762), .CP(clk), .Q(\gpr[19][23] ), .QN(n5453)
         );
  FD1 \gpr_reg[19][22]  ( .D(n2761), .CP(clk), .Q(\gpr[19][22] ), .QN(n5426)
         );
  FD1 \gpr_reg[19][21]  ( .D(n2760), .CP(clk), .Q(\gpr[19][21] ), .QN(n5404)
         );
  FD1 \gpr_reg[19][20]  ( .D(n2759), .CP(clk), .Q(\gpr[19][20] ), .QN(n5383)
         );
  FD1 \gpr_reg[19][19]  ( .D(n2758), .CP(clk), .Q(\gpr[19][19] ), .QN(n5349)
         );
  FD1 \gpr_reg[19][18]  ( .D(n2757), .CP(clk), .Q(\gpr[19][18] ), .QN(n5337)
         );
  FD1 \gpr_reg[19][17]  ( .D(n2756), .CP(clk), .Q(\gpr[19][17] ), .QN(n5325)
         );
  FD1 \gpr_reg[19][16]  ( .D(n2755), .CP(clk), .Q(\gpr[19][16] ), .QN(n5286)
         );
  FD1 \gpr_reg[19][15]  ( .D(n2754), .CP(clk), .Q(\gpr[19][15] ), .QN(n5254)
         );
  FD1 \gpr_reg[19][14]  ( .D(n2753), .CP(clk), .Q(\gpr[19][14] ), .QN(n5238)
         );
  FD1 \gpr_reg[19][13]  ( .D(n2752), .CP(clk), .Q(\gpr[19][13] ), .QN(n5211)
         );
  FD1 \gpr_reg[19][12]  ( .D(n2751), .CP(clk), .Q(\gpr[19][12] ), .QN(n5188)
         );
  FD1 \gpr_reg[19][11]  ( .D(n2750), .CP(clk), .Q(\gpr[19][11] ), .QN(n5158)
         );
  FD1 \gpr_reg[19][10]  ( .D(n2749), .CP(clk), .Q(\gpr[19][10] ), .QN(n5139)
         );
  FD1 \gpr_reg[19][9]  ( .D(n2748), .CP(clk), .Q(\gpr[19][9] ), .QN(n5111) );
  FD1 \gpr_reg[19][8]  ( .D(n2747), .CP(clk), .Q(\gpr[19][8] ), .QN(n5074) );
  FD1 \gpr_reg[19][7]  ( .D(n2746), .CP(clk), .Q(\gpr[19][7] ), .QN(n5054) );
  FD1 \gpr_reg[19][6]  ( .D(n2745), .CP(clk), .Q(\gpr[19][6] ), .QN(n5024) );
  FD1 \gpr_reg[19][5]  ( .D(n2744), .CP(clk), .Q(\gpr[19][5] ), .QN(n4995) );
  FD1 \gpr_reg[19][4]  ( .D(n2743), .CP(clk), .Q(\gpr[19][4] ), .QN(n4987) );
  FD1 \gpr_reg[19][3]  ( .D(n2742), .CP(clk), .Q(\gpr[19][3] ), .QN(n4958) );
  FD1 \gpr_reg[19][2]  ( .D(n2741), .CP(clk), .Q(\gpr[19][2] ), .QN(n4933) );
  FD1 \gpr_reg[19][1]  ( .D(n2740), .CP(clk), .Q(\gpr[19][1] ), .QN(n4909) );
  FD1 \gpr_reg[19][0]  ( .D(n2739), .CP(clk), .Q(\gpr[19][0] ), .QN(n4896) );
  FD1 \gpr_reg[20][31]  ( .D(n2738), .CP(clk), .Q(\gpr[20][31] ), .QN(n317) );
  FD1 \gpr_reg[20][30]  ( .D(n2737), .CP(clk), .Q(\gpr[20][30] ), .QN(n5628)
         );
  FD1 \gpr_reg[20][28]  ( .D(n2735), .CP(clk), .Q(\gpr[20][28] ), .QN(n5574)
         );
  FD1 \gpr_reg[20][27]  ( .D(n2734), .CP(clk), .Q(\gpr[20][27] ), .QN(n4877)
         );
  FD1 \gpr_reg[20][26]  ( .D(n2733), .CP(clk), .Q(\gpr[20][26] ), .QN(n5523)
         );
  FD1 \gpr_reg[20][25]  ( .D(n2732), .CP(clk), .Q(\gpr[20][25] ), .QN(n316) );
  FD1 \gpr_reg[20][24]  ( .D(n2731), .CP(clk), .Q(\gpr[20][24] ), .QN(n5474)
         );
  FD1 \gpr_reg[20][23]  ( .D(n2730), .CP(clk), .Q(\gpr[20][23] ) );
  FD1 \gpr_reg[20][22]  ( .D(n2729), .CP(clk), .Q(\gpr[20][22] ), .QN(n5425)
         );
  FD1 \gpr_reg[20][21]  ( .D(n2728), .CP(clk), .Q(\gpr[20][21] ), .QN(n4868)
         );
  FD1 \gpr_reg[20][20]  ( .D(n2727), .CP(clk), .Q(\gpr[20][20] ), .QN(n5378)
         );
  FD1 \gpr_reg[20][19]  ( .D(n2726), .CP(clk), .Q(\gpr[20][19] ), .QN(n312) );
  FD1 \gpr_reg[20][18]  ( .D(n2725), .CP(clk), .Q(\gpr[20][18] ), .QN(n5336)
         );
  FD1 \gpr_reg[20][17]  ( .D(n2724), .CP(clk), .Q(\gpr[20][17] ), .QN(n305) );
  FD1 \gpr_reg[20][16]  ( .D(n2723), .CP(clk), .Q(\gpr[20][16] ), .QN(n5285)
         );
  FD1 \gpr_reg[20][15]  ( .D(n2722), .CP(clk), .Q(\gpr[20][15] ), .QN(n5257)
         );
  FD1 \gpr_reg[20][14]  ( .D(n2721), .CP(clk), .Q(\gpr[20][14] ), .QN(n5233)
         );
  FD1 \gpr_reg[20][13]  ( .D(n2720), .CP(clk), .Q(\gpr[20][13] ), .QN(n5206)
         );
  FD1 \gpr_reg[20][12]  ( .D(n2719), .CP(clk), .Q(\gpr[20][12] ), .QN(n5186)
         );
  FD1 \gpr_reg[20][11]  ( .D(n2718), .CP(clk), .Q(\gpr[20][11] ), .QN(n5161)
         );
  FD1 \gpr_reg[20][10]  ( .D(n2717), .CP(clk), .Q(\gpr[20][10] ), .QN(n5134)
         );
  FD1 \gpr_reg[20][9]  ( .D(n2716), .CP(clk), .Q(\gpr[20][9] ), .QN(n5112) );
  FD1 \gpr_reg[20][8]  ( .D(n2715), .CP(clk), .Q(\gpr[20][8] ), .QN(n5073) );
  FD1 \gpr_reg[20][7]  ( .D(n2714), .CP(clk), .Q(\gpr[20][7] ), .QN(n303) );
  FD1 \gpr_reg[20][6]  ( .D(n2713), .CP(clk), .Q(\gpr[20][6] ), .QN(n5021) );
  FD1 \gpr_reg[20][5]  ( .D(n2712), .CP(clk), .Q(\gpr[20][5] ), .QN(n300) );
  FD1 \gpr_reg[20][4]  ( .D(n2711), .CP(clk), .Q(\gpr[20][4] ), .QN(n4983) );
  FD1 \gpr_reg[20][3]  ( .D(n2710), .CP(clk), .Q(\gpr[20][3] ), .QN(n4956) );
  FD1 \gpr_reg[20][2]  ( .D(n2709), .CP(clk), .Q(\gpr[20][2] ), .QN(n4937) );
  FD1 \gpr_reg[20][1]  ( .D(n2708), .CP(clk), .Q(\gpr[20][1] ), .QN(n4908) );
  FD1 \gpr_reg[20][0]  ( .D(n2707), .CP(clk), .Q(\gpr[20][0] ), .QN(n4891) );
  FD1 \gpr_reg[21][31]  ( .D(n2706), .CP(clk), .Q(\gpr[21][31] ), .QN(n5644)
         );
  FD1 \gpr_reg[21][30]  ( .D(n2705), .CP(clk), .Q(\gpr[21][30] ), .QN(n5624)
         );
  FD1 \gpr_reg[21][29]  ( .D(n2704), .CP(clk), .Q(\gpr[21][29] ), .QN(n5593)
         );
  FD1 \gpr_reg[21][28]  ( .D(n2703), .CP(clk), .Q(\gpr[21][28] ), .QN(n5573)
         );
  FD1 \gpr_reg[21][27]  ( .D(n2702), .CP(clk), .Q(\gpr[21][27] ), .QN(n5542)
         );
  FD1 \gpr_reg[21][26]  ( .D(n2701), .CP(clk), .Q(\gpr[21][26] ), .QN(n4876)
         );
  FD1 \gpr_reg[21][25]  ( .D(n2700), .CP(clk), .Q(\gpr[21][25] ), .QN(n5512)
         );
  FD1 \gpr_reg[21][24]  ( .D(n2699), .CP(clk), .Q(\gpr[21][24] ), .QN(n4776)
         );
  FD1 \gpr_reg[21][23]  ( .D(n2698), .CP(clk), .Q(\gpr[21][23] ), .QN(n5449)
         );
  FD1 \gpr_reg[21][22]  ( .D(n2697), .CP(clk), .Q(\gpr[21][22] ), .QN(n5424)
         );
  FD1 \gpr_reg[21][21]  ( .D(n2696), .CP(clk), .Q(\gpr[21][21] ), .QN(n5403)
         );
  FD1 \gpr_reg[21][20]  ( .D(n2695), .CP(clk), .Q(\gpr[21][20] ), .QN(n4832)
         );
  FD1 \gpr_reg[21][19]  ( .D(n2694), .CP(clk), .Q(\gpr[21][19] ), .QN(n5347)
         );
  FD1 \gpr_reg[21][18]  ( .D(n2693), .CP(clk), .Q(\gpr[21][18] ), .QN(n5335)
         );
  FD1 \gpr_reg[21][17]  ( .D(n2692), .CP(clk), .Q(\gpr[21][17] ), .QN(n5323)
         );
  FD1 \gpr_reg[21][16]  ( .D(n2691), .CP(clk), .Q(\gpr[21][16] ), .QN(n4807)
         );
  FD1 \gpr_reg[21][15]  ( .D(n2690), .CP(clk), .Q(\gpr[21][15] ), .QN(n5253)
         );
  FD1 \gpr_reg[21][14]  ( .D(n2689), .CP(clk), .Q(\gpr[21][14] ), .QN(n5232)
         );
  FD1 \gpr_reg[21][13]  ( .D(n2688), .CP(clk), .Q(\gpr[21][13] ), .QN(n5205)
         );
  FD1 \gpr_reg[21][12]  ( .D(n2687), .CP(clk), .Q(\gpr[21][12] ), .QN(n5185)
         );
  FD1 \gpr_reg[21][11]  ( .D(n2686), .CP(clk), .Q(\gpr[21][11] ), .QN(n5156)
         );
  FD1 \gpr_reg[21][10]  ( .D(n2685), .CP(clk), .Q(\gpr[21][10] ), .QN(n5133)
         );
  FD1 \gpr_reg[21][9]  ( .D(n2684), .CP(clk), .Q(\gpr[21][9] ), .QN(n5107) );
  FD1 \gpr_reg[21][8]  ( .D(n2683), .CP(clk), .Q(\gpr[21][8] ), .QN(n5072) );
  FD1 \gpr_reg[21][7]  ( .D(n2682), .CP(clk), .Q(\gpr[21][7] ), .QN(n5053) );
  FD1 \gpr_reg[21][6]  ( .D(n2681), .CP(clk), .Q(\gpr[21][6] ), .QN(n5020) );
  FD1 \gpr_reg[21][5]  ( .D(n2680), .CP(clk), .Q(\gpr[21][5] ), .QN(n4993) );
  FD1 \gpr_reg[21][4]  ( .D(n2679), .CP(clk), .Q(\gpr[21][4] ), .QN(n4982) );
  FD1 \gpr_reg[21][3]  ( .D(n2678), .CP(clk), .Q(\gpr[21][3] ), .QN(n4955) );
  FD1 \gpr_reg[21][2]  ( .D(n2677), .CP(clk), .Q(\gpr[21][2] ), .QN(n4932) );
  FD1 \gpr_reg[21][1]  ( .D(n2676), .CP(clk), .Q(\gpr[21][1] ), .QN(n4841) );
  FD1 \gpr_reg[21][0]  ( .D(n2675), .CP(clk), .Q(\gpr[21][0] ), .QN(n4894) );
  FD1 \gpr_reg[22][31]  ( .D(n2674), .CP(clk), .Q(\gpr[22][31] ), .QN(n4883)
         );
  FD1 \gpr_reg[22][30]  ( .D(n2673), .CP(clk), .Q(\gpr[22][30] ), .QN(n4882)
         );
  FD1 \gpr_reg[22][29]  ( .D(n2672), .CP(clk), .Q(\gpr[22][29] ), .QN(n4880)
         );
  FD1 \gpr_reg[22][28]  ( .D(n2671), .CP(clk), .Q(\gpr[22][28] ), .QN(n5576)
         );
  FD1 \gpr_reg[22][27]  ( .D(n2670), .CP(clk), .Q(\gpr[22][27] ), .QN(n5545)
         );
  FD1 \gpr_reg[22][26]  ( .D(n2669), .CP(clk), .Q(\gpr[22][26] ), .QN(n5526)
         );
  FD1 \gpr_reg[22][25]  ( .D(n2668), .CP(clk), .Q(\gpr[22][25] ), .QN(n4875)
         );
  FD1 \gpr_reg[22][24]  ( .D(n2667), .CP(clk), .Q(\gpr[22][24] ), .QN(n5477)
         );
  FD1 \gpr_reg[22][23]  ( .D(n2666), .CP(clk), .Q(\gpr[22][23] ), .QN(n4872)
         );
  FD1 \gpr_reg[22][22]  ( .D(n2665), .CP(clk), .Q(\gpr[22][22] ), .QN(n4870)
         );
  FD1 \gpr_reg[22][21]  ( .D(n2664), .CP(clk), .Q(\gpr[22][21] ), .QN(n5406)
         );
  FD1 \gpr_reg[22][20]  ( .D(n2663), .CP(clk), .Q(\gpr[22][20] ), .QN(n5381)
         );
  FD1 \gpr_reg[22][19]  ( .D(n2662), .CP(clk), .Q(\gpr[22][19] ), .QN(n4867)
         );
  FD1 \gpr_reg[22][18]  ( .D(n2661), .CP(clk), .Q(\gpr[22][18] ), .QN(n4865)
         );
  FD1 \gpr_reg[22][17]  ( .D(n2660), .CP(clk), .Q(\gpr[22][17] ), .QN(n4863)
         );
  FD1 \gpr_reg[22][16]  ( .D(n2659), .CP(clk), .Q(\gpr[22][16] ), .QN(n5288)
         );
  FD1 \gpr_reg[22][15]  ( .D(n2658), .CP(clk), .Q(\gpr[22][15] ), .QN(n4862)
         );
  FD1 \gpr_reg[22][14]  ( .D(n2657), .CP(clk), .Q(\gpr[22][14] ), .QN(n5236)
         );
  FD1 \gpr_reg[22][13]  ( .D(n2656), .CP(clk), .Q(\gpr[22][13] ), .QN(n5208)
         );
  FD1 \gpr_reg[22][12]  ( .D(n2655), .CP(clk), .Q(\gpr[22][12] ), .QN(n4856)
         );
  FD1 \gpr_reg[22][11]  ( .D(n2654), .CP(clk), .Q(\gpr[22][11] ), .QN(n4854)
         );
  FD1 \gpr_reg[22][10]  ( .D(n2653), .CP(clk), .Q(\gpr[22][10] ), .QN(n5136)
         );
  FD1 \gpr_reg[22][9]  ( .D(n2652), .CP(clk), .Q(\gpr[22][9] ), .QN(n4852) );
  FD1 \gpr_reg[22][8]  ( .D(n2651), .CP(clk), .Q(\gpr[22][8] ), .QN(n4850) );
  FD1 \gpr_reg[22][7]  ( .D(n2650), .CP(clk), .Q(\gpr[22][7] ), .QN(n4848) );
  FD1 \gpr_reg[22][6]  ( .D(n2649), .CP(clk), .Q(\gpr[22][6] ), .QN(n4846) );
  FD1 \gpr_reg[22][5]  ( .D(n2648), .CP(clk), .Q(\gpr[22][5] ), .QN(n4844) );
  FD1 \gpr_reg[22][4]  ( .D(n2647), .CP(clk), .Q(\gpr[22][4] ), .QN(n4805) );
  FD1 \gpr_reg[22][3]  ( .D(n2646), .CP(clk), .Q(\gpr[22][3] ), .QN(n4764) );
  FD1 \gpr_reg[22][2]  ( .D(n2645), .CP(clk), .Q(\gpr[22][2] ), .QN(n4763) );
  FD1 \gpr_reg[22][0]  ( .D(n2643), .CP(clk), .Q(\gpr[22][0] ), .QN(n4762) );
  FD1 \gpr_reg[23][31]  ( .D(n2642), .CP(clk), .Q(\gpr[23][31] ), .QN(n5649)
         );
  FD1 \gpr_reg[23][30]  ( .D(n2641), .CP(clk), .Q(\gpr[23][30] ), .QN(n5623)
         );
  FD1 \gpr_reg[23][29]  ( .D(n2640), .CP(clk), .Q(\gpr[23][29] ), .QN(n5598)
         );
  FD1 \gpr_reg[23][28]  ( .D(n2639), .CP(clk), .Q(\gpr[23][28] ), .QN(n4879)
         );
  FD1 \gpr_reg[23][27]  ( .D(n2638), .CP(clk), .Q(\gpr[23][27] ), .QN(n5548)
         );
  FD1 \gpr_reg[23][26]  ( .D(n2637), .CP(clk), .Q(\gpr[23][26] ), .QN(n5529)
         );
  FD1 \gpr_reg[23][25]  ( .D(n2636), .CP(clk), .Q(\gpr[23][25] ), .QN(n5511)
         );
  FD1 \gpr_reg[23][24]  ( .D(n2635), .CP(clk), .Q(\gpr[23][24] ), .QN(n5480)
         );
  FD1 \gpr_reg[23][23]  ( .D(n2634), .CP(clk), .Q(\gpr[23][23] ), .QN(n5448)
         );
  FD1 \gpr_reg[23][22]  ( .D(n2633), .CP(clk), .Q(\gpr[23][22] ), .QN(n5423)
         );
  FD1 \gpr_reg[23][21]  ( .D(n2632), .CP(clk), .Q(\gpr[23][21] ), .QN(n5409)
         );
  FD1 \gpr_reg[23][20]  ( .D(n2631), .CP(clk), .Q(\gpr[23][20] ), .QN(n5384)
         );
  FD1 \gpr_reg[23][19]  ( .D(n2630), .CP(clk), .Q(\gpr[23][19] ), .QN(n5352)
         );
  FD1 \gpr_reg[23][18]  ( .D(n2629), .CP(clk), .Q(\gpr[23][18] ), .QN(n5334)
         );
  FD1 \gpr_reg[23][17]  ( .D(n2628), .CP(clk), .Q(\gpr[23][17] ), .QN(n5322)
         );
  FD1 \gpr_reg[23][16]  ( .D(n2627), .CP(clk), .Q(\gpr[23][16] ), .QN(n5291)
         );
  FD1 \gpr_reg[23][15]  ( .D(n2626), .CP(clk), .Q(\gpr[23][15] ), .QN(n5252)
         );
  FD1 \gpr_reg[23][14]  ( .D(n2625), .CP(clk), .Q(\gpr[23][14] ), .QN(n4860)
         );
  FD1 \gpr_reg[23][13]  ( .D(n2624), .CP(clk), .Q(\gpr[23][13] ), .QN(n4858)
         );
  FD1 \gpr_reg[23][12]  ( .D(n2623), .CP(clk), .Q(\gpr[23][12] ), .QN(n5191)
         );
  FD1 \gpr_reg[23][11]  ( .D(n2622), .CP(clk), .Q(\gpr[23][11] ), .QN(n5155)
         );
  FD1 \gpr_reg[23][10]  ( .D(n2621), .CP(clk), .Q(\gpr[23][10] ), .QN(n4853)
         );
  FD1 \gpr_reg[23][9]  ( .D(n2620), .CP(clk), .Q(\gpr[23][9] ), .QN(n5106) );
  FD1 \gpr_reg[23][8]  ( .D(n2619), .CP(clk), .Q(\gpr[23][8] ), .QN(n5078) );
  FD1 \gpr_reg[23][7]  ( .D(n2618), .CP(clk), .Q(\gpr[23][7] ), .QN(n5058) );
  FD1 \gpr_reg[23][6]  ( .D(n2617), .CP(clk), .Q(\gpr[23][6] ), .QN(n5019) );
  FD1 \gpr_reg[23][5]  ( .D(n2616), .CP(clk), .Q(\gpr[23][5] ), .QN(n4998) );
  FD1 \gpr_reg[23][4]  ( .D(n2615), .CP(clk), .Q(\gpr[23][4] ), .QN(n4981) );
  FD1 \gpr_reg[23][3]  ( .D(n2614), .CP(clk), .Q(\gpr[23][3] ), .QN(n4960) );
  FD1 \gpr_reg[23][2]  ( .D(n2613), .CP(clk), .Q(\gpr[23][2] ), .QN(n4931) );
  FD1 \gpr_reg[23][1]  ( .D(n2612), .CP(clk), .Q(\gpr[23][1] ), .QN(n4910) );
  FD1 \gpr_reg[23][0]  ( .D(n2611), .CP(clk), .Q(\gpr[23][0] ), .QN(n4893) );
  FD1 \gpr_reg[24][31]  ( .D(n2610), .CP(clk), .Q(\gpr[24][31] ), .QN(n5651)
         );
  FD1 \gpr_reg[24][30]  ( .D(n2609), .CP(clk), .Q(\gpr[24][30] ), .QN(n5617)
         );
  FD1 \gpr_reg[24][29]  ( .D(n2608), .CP(clk), .Q(\gpr[24][29] ), .QN(n5600)
         );
  FD1 \gpr_reg[24][28]  ( .D(n2607), .CP(clk), .Q(\gpr[24][28] ), .QN(n5569)
         );
  FD1 \gpr_reg[24][27]  ( .D(n2606), .CP(clk), .Q(\gpr[24][27] ), .QN(n5550)
         );
  FD1 \gpr_reg[24][26]  ( .D(n2605), .CP(clk), .Q(\gpr[24][26] ), .QN(n5519)
         );
  FD1 \gpr_reg[24][25]  ( .D(n2604), .CP(clk), .Q(\gpr[24][25] ), .QN(n5497)
         );
  FD1 \gpr_reg[24][24]  ( .D(n2603), .CP(clk), .Q(\gpr[24][24] ), .QN(n5469)
         );
  FD1 \gpr_reg[24][22]  ( .D(n2601), .CP(clk), .Q(\gpr[24][22] ), .QN(n5432)
         );
  FD1 \gpr_reg[24][21]  ( .D(n2600), .CP(clk), .Q(\gpr[24][21] ), .QN(n5398)
         );
  FD1 \gpr_reg[24][20]  ( .D(n2599), .CP(clk), .Q(\gpr[24][20] ), .QN(n5371)
         );
  FD1 \gpr_reg[24][18]  ( .D(n2597), .CP(clk), .Q(\gpr[24][18] ), .QN(n5328)
         );
  FD1 \gpr_reg[24][17]  ( .D(n2596), .CP(clk), .Q(\gpr[24][17] ), .QN(n5308)
         );
  FD1 \gpr_reg[24][16]  ( .D(n2595), .CP(clk), .Q(\gpr[24][16] ), .QN(n5279)
         );
  FD1 \gpr_reg[24][15]  ( .D(n2594), .CP(clk), .Q(\gpr[24][15] ), .QN(n5260)
         );
  FD1 \gpr_reg[24][14]  ( .D(n2593), .CP(clk), .Q(\gpr[24][14] ), .QN(n5226)
         );
  FD1 \gpr_reg[24][13]  ( .D(n2592), .CP(clk), .Q(\gpr[24][13] ), .QN(n5200)
         );
  FD1 \gpr_reg[24][12]  ( .D(n2591), .CP(clk), .Q(\gpr[24][12] ), .QN(n5183)
         );
  FD1 \gpr_reg[24][11]  ( .D(n2590), .CP(clk), .Q(\gpr[24][11] ), .QN(n5163)
         );
  FD1 \gpr_reg[24][10]  ( .D(n2589), .CP(clk), .Q(\gpr[24][10] ), .QN(n5128)
         );
  FD1 \gpr_reg[24][9]  ( .D(n2588), .CP(clk), .Q(\gpr[24][9] ), .QN(n5101) );
  FD1 \gpr_reg[24][8]  ( .D(n2587), .CP(clk), .Q(\gpr[24][8] ), .QN(n5080) );
  FD1 \gpr_reg[24][7]  ( .D(n2586), .CP(clk), .Q(\gpr[24][7] ), .QN(n5049) );
  FD1 \gpr_reg[24][6]  ( .D(n2585), .CP(clk), .Q(\gpr[24][6] ), .QN(n5027) );
  FD1 \gpr_reg[24][5]  ( .D(n2584), .CP(clk), .Q(\gpr[24][5] ), .QN(n5000) );
  FD1 \gpr_reg[24][4]  ( .D(n2583), .CP(clk), .Q(\gpr[24][4] ), .QN(n4979) );
  FD1 \gpr_reg[24][3]  ( .D(n2582), .CP(clk), .Q(\gpr[24][3] ), .QN(n4951) );
  FD1 \gpr_reg[24][2]  ( .D(n2581), .CP(clk), .Q(\gpr[24][2] ), .QN(n4926) );
  FD1 \gpr_reg[24][1]  ( .D(n2580), .CP(clk), .Q(\gpr[24][1] ), .QN(n4922) );
  FD1 \gpr_reg[24][0]  ( .D(n2579), .CP(clk), .Q(\gpr[24][0] ), .QN(n4888) );
  FD1 \gpr_reg[25][31]  ( .D(n2578), .CP(clk), .Q(\gpr[25][31] ), .QN(n5653)
         );
  FD1 \gpr_reg[25][30]  ( .D(n2577), .CP(clk), .Q(\gpr[25][30] ), .QN(n5619)
         );
  FD1 \gpr_reg[25][28]  ( .D(n2575), .CP(clk), .Q(\gpr[25][28] ), .QN(n5571)
         );
  FD1 \gpr_reg[25][27]  ( .D(n2574), .CP(clk), .Q(\gpr[25][27] ), .QN(n5552)
         );
  FD1 \gpr_reg[25][26]  ( .D(n2573), .CP(clk), .Q(\gpr[25][26] ), .QN(n5521)
         );
  FD1 \gpr_reg[25][25]  ( .D(n2572), .CP(clk), .Q(\gpr[25][25] ), .QN(n5498)
         );
  FD1 \gpr_reg[25][24]  ( .D(n2571), .CP(clk), .Q(\gpr[25][24] ), .QN(n5473)
         );
  FD1 \gpr_reg[25][23]  ( .D(n2570), .CP(clk), .Q(\gpr[25][23] ), .QN(n5447)
         );
  FD1 \gpr_reg[25][22]  ( .D(n2569), .CP(clk), .Q(\gpr[25][22] ), .QN(n5435)
         );
  FD1 \gpr_reg[25][21]  ( .D(n2568), .CP(clk), .Q(\gpr[25][21] ), .QN(n5401)
         );
  FD1 \gpr_reg[25][20]  ( .D(n2567), .CP(clk), .Q(\gpr[25][20] ), .QN(n5373)
         );
  FD1 \gpr_reg[25][19]  ( .D(n2566), .CP(clk), .Q(\gpr[25][19] ), .QN(n5355)
         );
  FD1 \gpr_reg[25][18]  ( .D(n2565), .CP(clk), .Q(\gpr[25][18] ), .QN(n5330)
         );
  FD1 \gpr_reg[25][17]  ( .D(n2564), .CP(clk), .Q(\gpr[25][17] ), .QN(n5309)
         );
  FD1 \gpr_reg[25][16]  ( .D(n2563), .CP(clk), .Q(\gpr[25][16] ), .QN(n5283)
         );
  FD1 \gpr_reg[25][15]  ( .D(n2562), .CP(clk), .Q(\gpr[25][15] ), .QN(n5263)
         );
  FD1 \gpr_reg[25][14]  ( .D(n2561), .CP(clk), .Q(\gpr[25][14] ), .QN(n5227)
         );
  FD1 \gpr_reg[25][13]  ( .D(n2560), .CP(clk), .Q(\gpr[25][13] ), .QN(n5201)
         );
  FD1 \gpr_reg[25][12]  ( .D(n2559), .CP(clk), .Q(\gpr[25][12] ), .QN(n5181)
         );
  FD1 \gpr_reg[25][11]  ( .D(n2558), .CP(clk), .Q(\gpr[25][11] ), .QN(n5166)
         );
  FD1 \gpr_reg[25][10]  ( .D(n2557), .CP(clk), .Q(\gpr[25][10] ), .QN(n5129)
         );
  FD1 \gpr_reg[25][9]  ( .D(n2556), .CP(clk), .Q(\gpr[25][9] ), .QN(n5102) );
  FD1 \gpr_reg[25][8]  ( .D(n2555), .CP(clk), .Q(\gpr[25][8] ), .QN(n5084) );
  FD1 \gpr_reg[25][7]  ( .D(n2554), .CP(clk), .Q(\gpr[25][7] ), .QN(n5052) );
  FD1 \gpr_reg[25][6]  ( .D(n2553), .CP(clk), .Q(\gpr[25][6] ), .QN(n5028) );
  FD1 \gpr_reg[25][5]  ( .D(n2552), .CP(clk), .Q(\gpr[25][5] ), .QN(n5001) );
  FD1 \gpr_reg[25][4]  ( .D(n2551), .CP(clk), .Q(\gpr[25][4] ), .QN(n4980) );
  FD1 \gpr_reg[25][3]  ( .D(n2550), .CP(clk), .Q(\gpr[25][3] ), .QN(n4953) );
  FD1 \gpr_reg[25][2]  ( .D(n2549), .CP(clk), .Q(\gpr[25][2] ), .QN(n4929) );
  FD1 \gpr_reg[25][0]  ( .D(n2547), .CP(clk), .Q(\gpr[25][0] ), .QN(n4890) );
  FD1 \gpr_reg[26][31]  ( .D(n2546), .CP(clk), .Q(\gpr[26][31] ), .QN(n5654)
         );
  FD1 \gpr_reg[26][30]  ( .D(n2545), .CP(clk), .Q(\gpr[26][30] ), .QN(n5620)
         );
  FD1 \gpr_reg[26][29]  ( .D(n2544), .CP(clk), .Q(\gpr[26][29] ), .QN(n5601)
         );
  FD1 \gpr_reg[26][28]  ( .D(n2543), .CP(clk), .Q(\gpr[26][28] ), .QN(n5570)
         );
  FD1 \gpr_reg[26][27]  ( .D(n2542), .CP(clk), .Q(\gpr[26][27] ), .QN(n5554)
         );
  FD1 \gpr_reg[26][26]  ( .D(n2541), .CP(clk), .Q(\gpr[26][26] ), .QN(n5520)
         );
  FD1 \gpr_reg[26][25]  ( .D(n2540), .CP(clk), .Q(\gpr[26][25] ), .QN(n4797)
         );
  FD1 \gpr_reg[26][24]  ( .D(n2539), .CP(clk), .Q(\gpr[26][24] ), .QN(n5472)
         );
  FD1 \gpr_reg[26][23]  ( .D(n2538), .CP(clk), .Q(\gpr[26][23] ), .QN(n5446)
         );
  FD1 \gpr_reg[26][22]  ( .D(n2537), .CP(clk), .Q(\gpr[26][22] ), .QN(n5434)
         );
  FD1 \gpr_reg[26][21]  ( .D(n2536), .CP(clk), .Q(\gpr[26][21] ), .QN(n5400)
         );
  FD1 \gpr_reg[26][20]  ( .D(n2535), .CP(clk), .Q(\gpr[26][20] ), .QN(n5375)
         );
  FD1 \gpr_reg[26][19]  ( .D(n2534), .CP(clk), .Q(\gpr[26][19] ), .QN(n5356)
         );
  FD1 \gpr_reg[26][18]  ( .D(n2533), .CP(clk), .Q(\gpr[26][18] ), .QN(n5332)
         );
  FD1 \gpr_reg[26][17]  ( .D(n2532), .CP(clk), .Q(\gpr[26][17] ), .QN(n4789)
         );
  FD1 \gpr_reg[26][16]  ( .D(n2531), .CP(clk), .Q(\gpr[26][16] ), .QN(n5282)
         );
  FD1 \gpr_reg[26][15]  ( .D(n2530), .CP(clk), .Q(\gpr[26][15] ), .QN(n5262)
         );
  FD1 \gpr_reg[26][14]  ( .D(n2529), .CP(clk), .Q(\gpr[26][14] ), .QN(n5229)
         );
  FD1 \gpr_reg[26][13]  ( .D(n2528), .CP(clk), .Q(\gpr[26][13] ), .QN(n5202)
         );
  FD1 \gpr_reg[26][12]  ( .D(n2527), .CP(clk), .Q(\gpr[26][12] ), .QN(n5182)
         );
  FD1 \gpr_reg[26][11]  ( .D(n2526), .CP(clk), .Q(\gpr[26][11] ), .QN(n5165)
         );
  FD1 \gpr_reg[26][10]  ( .D(n2525), .CP(clk), .Q(\gpr[26][10] ), .QN(n5131)
         );
  FD1 \gpr_reg[26][9]  ( .D(n2524), .CP(clk), .Q(\gpr[26][9] ), .QN(n5103) );
  FD1 \gpr_reg[26][8]  ( .D(n2523), .CP(clk), .Q(\gpr[26][8] ), .QN(n5083) );
  FD1 \gpr_reg[26][7]  ( .D(n2522), .CP(clk), .Q(\gpr[26][7] ), .QN(n5051) );
  FD1 \gpr_reg[26][6]  ( .D(n2521), .CP(clk), .Q(\gpr[26][6] ), .QN(n5029) );
  FD1 \gpr_reg[26][5]  ( .D(n2520), .CP(clk), .Q(\gpr[26][5] ), .QN(n5003) );
  FD1 \gpr_reg[26][4]  ( .D(n2519), .CP(clk), .Q(\gpr[26][4] ), .QN(n4978) );
  FD1 \gpr_reg[26][3]  ( .D(n2518), .CP(clk), .Q(\gpr[26][3] ), .QN(n4779) );
  FD1 \gpr_reg[26][2]  ( .D(n2517), .CP(clk), .Q(\gpr[26][2] ), .QN(n4928) );
  FD1 \gpr_reg[26][1]  ( .D(n2516), .CP(clk), .Q(\gpr[26][1] ), .QN(n4835) );
  FD1 \gpr_reg[26][0]  ( .D(n2515), .CP(clk), .Q(\gpr[26][0] ), .QN(n4885) );
  FD1 \gpr_reg[27][31]  ( .D(n2514), .CP(clk), .Q(\gpr[27][31] ), .QN(n5652)
         );
  FD1 \gpr_reg[27][30]  ( .D(n2513), .CP(clk), .Q(\gpr[27][30] ), .QN(n5618)
         );
  FD1 \gpr_reg[27][28]  ( .D(n2511), .CP(clk), .Q(\gpr[27][28] ), .QN(n5572)
         );
  FD1 \gpr_reg[27][27]  ( .D(n2510), .CP(clk), .Q(\gpr[27][27] ), .QN(n5551)
         );
  FD1 \gpr_reg[27][26]  ( .D(n2509), .CP(clk), .Q(\gpr[27][26] ), .QN(n5522)
         );
  FD1 \gpr_reg[27][25]  ( .D(n2508), .CP(clk), .Q(\gpr[27][25] ), .QN(n5494)
         );
  FD1 \gpr_reg[27][24]  ( .D(n2507), .CP(clk), .Q(\gpr[27][24] ), .QN(n5470)
         );
  FD1 \gpr_reg[27][23]  ( .D(n2506), .CP(clk), .Q(\gpr[27][23] ), .QN(n5445)
         );
  FD1 \gpr_reg[27][22]  ( .D(n2505), .CP(clk), .Q(\gpr[27][22] ), .QN(n5433)
         );
  FD1 \gpr_reg[27][21]  ( .D(n2504), .CP(clk), .Q(\gpr[27][21] ), .QN(n5399)
         );
  FD1 \gpr_reg[27][20]  ( .D(n2503), .CP(clk), .Q(\gpr[27][20] ), .QN(n5372)
         );
  FD1 \gpr_reg[27][19]  ( .D(n2502), .CP(clk), .Q(\gpr[27][19] ), .QN(n5354)
         );
  FD1 \gpr_reg[27][18]  ( .D(n2501), .CP(clk), .Q(\gpr[27][18] ), .QN(n5329)
         );
  FD1 \gpr_reg[27][17]  ( .D(n2500), .CP(clk), .Q(\gpr[27][17] ), .QN(n5305)
         );
  FD1 \gpr_reg[27][16]  ( .D(n2499), .CP(clk), .Q(\gpr[27][16] ), .QN(n5280)
         );
  FD1 \gpr_reg[27][15]  ( .D(n2498), .CP(clk), .Q(\gpr[27][15] ), .QN(n5261)
         );
  FD1 \gpr_reg[27][14]  ( .D(n2497), .CP(clk), .Q(\gpr[27][14] ), .QN(n5230)
         );
  FD1 \gpr_reg[27][13]  ( .D(n2496), .CP(clk), .Q(\gpr[27][13] ), .QN(n5203)
         );
  FD1 \gpr_reg[27][12]  ( .D(n2495), .CP(clk), .Q(\gpr[27][12] ), .QN(n5180)
         );
  FD1 \gpr_reg[27][11]  ( .D(n2494), .CP(clk), .Q(\gpr[27][11] ), .QN(n5164)
         );
  FD1 \gpr_reg[27][10]  ( .D(n2493), .CP(clk), .Q(\gpr[27][10] ), .QN(n5132)
         );
  FD1 \gpr_reg[27][9]  ( .D(n2492), .CP(clk), .Q(\gpr[27][9] ), .QN(n5104) );
  FD1 \gpr_reg[27][8]  ( .D(n2491), .CP(clk), .Q(\gpr[27][8] ), .QN(n5081) );
  FD1 \gpr_reg[27][7]  ( .D(n2490), .CP(clk), .Q(\gpr[27][7] ), .QN(n5050) );
  FD1 \gpr_reg[27][6]  ( .D(n2489), .CP(clk), .Q(\gpr[27][6] ), .QN(n5030) );
  FD1 \gpr_reg[27][5]  ( .D(n2488), .CP(clk), .Q(\gpr[27][5] ), .QN(n5004) );
  FD1 \gpr_reg[27][4]  ( .D(n2487), .CP(clk), .Q(\gpr[27][4] ), .QN(n4977) );
  FD1 \gpr_reg[27][3]  ( .D(n2486), .CP(clk), .Q(\gpr[27][3] ), .QN(n4952) );
  FD1 \gpr_reg[27][2]  ( .D(n2485), .CP(clk), .Q(\gpr[27][2] ), .QN(n4927) );
  FD1 \gpr_reg[27][0]  ( .D(n2483), .CP(clk), .Q(\gpr[27][0] ), .QN(n4889) );
  FD1 \gpr_reg[28][31]  ( .D(n2482), .CP(clk), .Q(\gpr[28][31] ), .QN(n318) );
  FD1 \gpr_reg[28][30]  ( .D(n2481), .CP(clk), .Q(\gpr[28][30] ), .QN(n5621)
         );
  FD1 \gpr_reg[28][28]  ( .D(n2479), .CP(clk), .Q(\gpr[28][28] ), .QN(n5568)
         );
  FD1 \gpr_reg[28][27]  ( .D(n2478), .CP(clk), .Q(\gpr[28][27] ), .QN(n5555)
         );
  FD1 \gpr_reg[28][26]  ( .D(n2477), .CP(clk), .Q(\gpr[28][26] ), .QN(n5518)
         );
  FD1 \gpr_reg[28][25]  ( .D(n2476), .CP(clk), .Q(\gpr[28][25] ), .QN(n314) );
  FD1 \gpr_reg[28][24]  ( .D(n2475), .CP(clk), .Q(\gpr[28][24] ), .QN(n5468)
         );
  FD1 \gpr_reg[28][23]  ( .D(n2474), .CP(clk), .Q(\gpr[28][23] ) );
  FD1 \gpr_reg[28][22]  ( .D(n2473), .CP(clk), .Q(\gpr[28][22] ), .QN(n5431)
         );
  FD1 \gpr_reg[28][20]  ( .D(n2471), .CP(clk), .Q(\gpr[28][20] ), .QN(n5376)
         );
  FD1 \gpr_reg[28][19]  ( .D(n2470), .CP(clk), .Q(\gpr[28][19] ), .QN(n313) );
  FD1 \gpr_reg[28][18]  ( .D(n2469), .CP(clk), .QN(n4770) );
  FD1 \gpr_reg[28][17]  ( .D(n2468), .CP(clk), .Q(\gpr[28][17] ), .QN(n304) );
  FD1 \gpr_reg[28][16]  ( .D(n2467), .CP(clk), .Q(\gpr[28][16] ), .QN(n5284)
         );
  FD1 \gpr_reg[28][15]  ( .D(n2466), .CP(clk), .Q(\gpr[28][15] ), .QN(n5264)
         );
  FD1 \gpr_reg[28][14]  ( .D(n2465), .CP(clk), .Q(\gpr[28][14] ), .QN(n5225)
         );
  FD1 \gpr_reg[28][13]  ( .D(n2464), .CP(clk), .Q(\gpr[28][13] ), .QN(n5204)
         );
  FD1 \gpr_reg[28][12]  ( .D(n2463), .CP(clk), .Q(\gpr[28][12] ), .QN(n5179)
         );
  FD1 \gpr_reg[28][11]  ( .D(n2462), .CP(clk), .Q(\gpr[28][11] ) );
  FD1 \gpr_reg[28][10]  ( .D(n2461), .CP(clk), .Q(\gpr[28][10] ), .QN(n5127)
         );
  FD1 \gpr_reg[28][9]  ( .D(n2460), .CP(clk), .Q(\gpr[28][9] ), .QN(n5105) );
  FD1 \gpr_reg[28][8]  ( .D(n2459), .CP(clk), .Q(\gpr[28][8] ), .QN(n5079) );
  FD1 \gpr_reg[28][7]  ( .D(n2458), .CP(clk), .Q(\gpr[28][7] ), .QN(n302) );
  FD1 \gpr_reg[28][6]  ( .D(n2457), .CP(clk), .Q(\gpr[28][6] ), .QN(n5031) );
  FD1 \gpr_reg[28][5]  ( .D(n2456), .CP(clk), .Q(\gpr[28][5] ), .QN(n4845) );
  FD1 \gpr_reg[28][4]  ( .D(n2455), .CP(clk), .Q(\gpr[28][4] ), .QN(n4976) );
  FD1 \gpr_reg[28][3]  ( .D(n2454), .CP(clk), .Q(\gpr[28][3] ), .QN(n4950) );
  FD1 \gpr_reg[28][2]  ( .D(n2453), .CP(clk), .Q(\gpr[28][2] ), .QN(n4925) );
  FD1 \gpr_reg[28][1]  ( .D(n2452), .CP(clk), .Q(\gpr[28][1] ), .QN(n4921) );
  FD1 \gpr_reg[28][0]  ( .D(n2451), .CP(clk), .Q(\gpr[28][0] ), .QN(n4887) );
  FD1 \gpr_reg[29][31]  ( .D(n2450), .CP(clk), .Q(\gpr[29][31] ), .QN(n5650)
         );
  FD1 \gpr_reg[29][30]  ( .D(n2449), .CP(clk), .Q(\gpr[29][30] ), .QN(n5622)
         );
  FD1 \gpr_reg[29][29]  ( .D(n2448), .CP(clk), .Q(\gpr[29][29] ), .QN(n5599)
         );
  FD1 \gpr_reg[29][28]  ( .D(n2447), .CP(clk), .Q(\gpr[29][28] ), .QN(n5567)
         );
  FD1 \gpr_reg[29][27]  ( .D(n2446), .CP(clk), .Q(\gpr[29][27] ), .QN(n4834)
         );
  FD1 \gpr_reg[29][26]  ( .D(n2445), .CP(clk), .Q(\gpr[29][26] ), .QN(n5517)
         );
  FD1 \gpr_reg[29][25]  ( .D(n2444), .CP(clk), .Q(\gpr[29][25] ), .QN(n5496)
         );
  FD1 \gpr_reg[29][24]  ( .D(n2443), .CP(clk), .Q(\gpr[29][24] ), .QN(n5467)
         );
  FD1 \gpr_reg[29][23]  ( .D(n2442), .CP(clk), .Q(\gpr[29][23] ), .QN(n5444)
         );
  FD1 \gpr_reg[29][22]  ( .D(n2441), .CP(clk), .Q(\gpr[29][22] ), .QN(n5430)
         );
  FD1 \gpr_reg[29][21]  ( .D(n2440), .CP(clk), .Q(\gpr[29][21] ), .QN(n5397)
         );
  FD1 \gpr_reg[29][20]  ( .D(n2439), .CP(clk), .Q(\gpr[29][20] ), .QN(n4833)
         );
  FD1 \gpr_reg[29][19]  ( .D(n2438), .CP(clk), .Q(\gpr[29][19] ), .QN(n5353)
         );
  FD1 \gpr_reg[29][18]  ( .D(n2437), .CP(clk), .Q(\gpr[29][18] ), .QN(n5327)
         );
  FD1 \gpr_reg[29][17]  ( .D(n2436), .CP(clk), .Q(\gpr[29][17] ), .QN(n5307)
         );
  FD1 \gpr_reg[29][16]  ( .D(n2435), .CP(clk), .Q(\gpr[29][16] ), .QN(n4831)
         );
  FD1 \gpr_reg[29][15]  ( .D(n2434), .CP(clk), .Q(\gpr[29][15] ), .QN(n5259)
         );
  FD1 \gpr_reg[29][14]  ( .D(n2433), .CP(clk), .Q(\gpr[29][14] ), .QN(n4830)
         );
  FD1 \gpr_reg[29][13]  ( .D(n2432), .CP(clk), .Q(\gpr[29][13] ), .QN(n5199)
         );
  FD1 \gpr_reg[29][12]  ( .D(n2431), .CP(clk), .Q(\gpr[29][12] ), .QN(n5178)
         );
  FD1 \gpr_reg[29][11]  ( .D(n2430), .CP(clk), .Q(\gpr[29][11] ), .QN(n5162)
         );
  FD1 \gpr_reg[29][10]  ( .D(n2429), .CP(clk), .Q(\gpr[29][10] ), .QN(n4829)
         );
  FD1 \gpr_reg[29][9]  ( .D(n2428), .CP(clk), .Q(\gpr[29][9] ), .QN(n5100) );
  FD1 \gpr_reg[29][8]  ( .D(n2427), .CP(clk), .Q(\gpr[29][8] ), .QN(n4828) );
  FD1 \gpr_reg[29][7]  ( .D(n2426), .CP(clk), .Q(\gpr[29][7] ), .QN(n5048) );
  FD1 \gpr_reg[29][6]  ( .D(n2425), .CP(clk), .Q(\gpr[29][6] ), .QN(n5026) );
  FD1 \gpr_reg[29][5]  ( .D(n2424), .CP(clk), .Q(\gpr[29][5] ), .QN(n4999) );
  FD1 \gpr_reg[29][4]  ( .D(n2423), .CP(clk), .Q(\gpr[29][4] ), .QN(n4975) );
  FD1 \gpr_reg[29][3]  ( .D(n2422), .CP(clk), .Q(\gpr[29][3] ), .QN(n4949) );
  FD1 \gpr_reg[29][2]  ( .D(n2421), .CP(clk), .Q(\gpr[29][2] ), .QN(n4924) );
  FD1 \gpr_reg[29][1]  ( .D(n2420), .CP(clk), .Q(\gpr[29][1] ), .QN(n4827) );
  FD1 \gpr_reg[29][0]  ( .D(n2419), .CP(clk), .Q(\gpr[29][0] ), .QN(n4886) );
  FD1 \gpr_reg[30][31]  ( .D(n2418), .CP(clk), .QN(n4811) );
  FD1 \gpr_reg[30][30]  ( .D(n2417), .CP(clk), .Q(\gpr[30][30] ), .QN(n4881)
         );
  FD1 \gpr_reg[30][29]  ( .D(n2416), .CP(clk), .QN(n4810) );
  FD1 \gpr_reg[30][28]  ( .D(n2415), .CP(clk), .Q(\gpr[30][28] ), .QN(n4878)
         );
  FD1 \gpr_reg[30][27]  ( .D(n2414), .CP(clk), .Q(\gpr[30][27] ), .QN(n5553)
         );
  FD1 \gpr_reg[30][26]  ( .D(n2413), .CP(clk), .Q(\gpr[30][26] ), .QN(n4809)
         );
  FD1 \gpr_reg[30][25]  ( .D(n2412), .CP(clk), .Q(\gpr[30][25] ), .QN(n4874)
         );
  FD1 \gpr_reg[30][24]  ( .D(n2411), .CP(clk), .Q(\gpr[30][24] ), .QN(n5471)
         );
  FD1 \gpr_reg[30][23]  ( .D(n2410), .CP(clk), .Q(\gpr[30][23] ), .QN(n4873)
         );
  FD1 \gpr_reg[30][22]  ( .D(n2409), .CP(clk), .Q(\gpr[30][22] ), .QN(n4871)
         );
  FD1 \gpr_reg[30][21]  ( .D(n2408), .CP(clk), .Q(\gpr[30][21] ), .QN(n4869)
         );
  FD1 \gpr_reg[30][20]  ( .D(n2407), .CP(clk), .Q(\gpr[30][20] ), .QN(n5374)
         );
  FD1 \gpr_reg[30][19]  ( .D(n2406), .CP(clk), .Q(\gpr[30][19] ), .QN(n4866)
         );
  FD1 \gpr_reg[30][18]  ( .D(n2405), .CP(clk), .Q(\gpr[30][18] ), .QN(n5331)
         );
  FD1 \gpr_reg[30][17]  ( .D(n2404), .CP(clk), .Q(\gpr[30][17] ), .QN(n4864)
         );
  FD1 \gpr_reg[30][16]  ( .D(n2403), .CP(clk), .Q(\gpr[30][16] ), .QN(n5281)
         );
  FD1 \gpr_reg[30][15]  ( .D(n2402), .CP(clk), .Q(\gpr[30][15] ), .QN(n4861)
         );
  FD1 \gpr_reg[30][14]  ( .D(n2401), .CP(clk), .Q(\gpr[30][14] ), .QN(n5228)
         );
  FD1 \gpr_reg[30][13]  ( .D(n2400), .CP(clk), .Q(\gpr[30][13] ), .QN(n4859)
         );
  FD1 \gpr_reg[30][12]  ( .D(n2399), .CP(clk), .Q(\gpr[30][12] ), .QN(n4857)
         );
  FD1 \gpr_reg[30][11]  ( .D(n2398), .CP(clk), .Q(\gpr[30][11] ), .QN(n4855)
         );
  FD1 \gpr_reg[30][10]  ( .D(n2397), .CP(clk), .Q(\gpr[30][10] ), .QN(n5130)
         );
  FD1 \gpr_reg[30][9]  ( .D(n2396), .CP(clk), .Q(\gpr[30][9] ), .QN(n4851) );
  FD1 \gpr_reg[30][8]  ( .D(n2395), .CP(clk), .Q(\gpr[30][8] ), .QN(n5082) );
  FD1 \gpr_reg[30][7]  ( .D(n2394), .CP(clk), .Q(\gpr[30][7] ), .QN(n4849) );
  FD1 \gpr_reg[30][6]  ( .D(n2393), .CP(clk), .Q(\gpr[30][6] ), .QN(n4847) );
  FD1 \gpr_reg[30][5]  ( .D(n2392), .CP(clk), .Q(\gpr[30][5] ), .QN(n5002) );
  FD1 \gpr_reg[30][4]  ( .D(n2391), .CP(clk), .Q(\gpr[30][4] ), .QN(n4806) );
  FD1 \gpr_reg[30][3]  ( .D(n2390), .CP(clk), .Q(\gpr[30][3] ), .QN(n4843) );
  FD1 \gpr_reg[30][2]  ( .D(n2389), .CP(clk), .Q(\gpr[30][2] ), .QN(n4842) );
  FD1 \gpr_reg[30][1]  ( .D(n2388), .CP(clk), .Q(\gpr[30][1] ), .QN(n4923) );
  FD1 \gpr_reg[30][0]  ( .D(n2387), .CP(clk), .Q(\gpr[30][0] ), .QN(n4884) );
  FD1 \gpr_reg[31][31]  ( .D(n2386), .CP(clk), .Q(\gpr[31][31] ), .QN(n5655)
         );
  FD1 \gpr_reg[31][30]  ( .D(n2385), .CP(clk), .Q(\gpr[31][30] ), .QN(n5616)
         );
  FD1 \gpr_reg[31][29]  ( .D(n2384), .CP(clk), .Q(\gpr[31][29] ), .QN(n5602)
         );
  FD1 \gpr_reg[31][28]  ( .D(n2383), .CP(clk), .Q(\gpr[31][28] ), .QN(n5566)
         );
  FD1 \gpr_reg[31][27]  ( .D(n2382), .CP(clk), .Q(\gpr[31][27] ), .QN(n5549)
         );
  FD1 \gpr_reg[31][26]  ( .D(n2381), .CP(clk), .Q(\gpr[31][26] ), .QN(n5516)
         );
  FD1 \gpr_reg[31][25]  ( .D(n2380), .CP(clk), .Q(\gpr[31][25] ), .QN(n5495)
         );
  FD1 \gpr_reg[31][24]  ( .D(n2379), .CP(clk), .Q(\gpr[31][24] ), .QN(n4808)
         );
  FD1 \gpr_reg[31][23]  ( .D(n2378), .CP(clk), .Q(\gpr[31][23] ), .QN(n5443)
         );
  FD1 \gpr_reg[31][22]  ( .D(n2377), .CP(clk), .Q(\gpr[31][22] ), .QN(n5436)
         );
  FD1 \gpr_reg[31][21]  ( .D(n2376), .CP(clk), .Q(\gpr[31][21] ), .QN(n5402)
         );
  FD1 \gpr_reg[31][20]  ( .D(n2375), .CP(clk), .Q(\gpr[31][20] ), .QN(n5377)
         );
  FD1 \gpr_reg[31][19]  ( .D(n2374), .CP(clk), .Q(\gpr[31][19] ), .QN(n5357)
         );
  FD1 \gpr_reg[31][18]  ( .D(n2373), .CP(clk), .Q(\gpr[31][18] ), .QN(n5333)
         );
  FD1 \gpr_reg[31][17]  ( .D(n2372), .CP(clk), .Q(\gpr[31][17] ), .QN(n5306)
         );
  FD1 \gpr_reg[31][16]  ( .D(n2371), .CP(clk), .Q(\gpr[31][16] ), .QN(n5278)
         );
  FD1 \gpr_reg[31][15]  ( .D(n2370), .CP(clk), .Q(\gpr[31][15] ), .QN(n5258)
         );
  FD1 \gpr_reg[31][14]  ( .D(n2369), .CP(clk), .Q(\gpr[31][14] ), .QN(n5231)
         );
  FD1 \gpr_reg[31][13]  ( .D(n2368), .CP(clk), .Q(\gpr[31][13] ), .QN(n5198)
         );
  FD1 \gpr_reg[31][12]  ( .D(n2367), .CP(clk), .Q(\gpr[31][12] ), .QN(n5184)
         );
  FD1 \gpr_reg[31][11]  ( .D(n2366), .CP(clk), .Q(\gpr[31][11] ), .QN(n5167)
         );
  FD1 \gpr_reg[31][10]  ( .D(n2365), .CP(clk), .Q(\gpr[31][10] ), .QN(n5126)
         );
  FD1 \gpr_reg[31][9]  ( .D(n2364), .CP(clk), .Q(\gpr[31][9] ), .QN(n5099) );
  FD1 \gpr_reg[31][8]  ( .D(n2363), .CP(clk), .Q(\gpr[31][8] ), .QN(n5085) );
  FD1 \gpr_reg[31][7]  ( .D(n2362), .CP(clk), .Q(\gpr[31][7] ), .QN(n5047) );
  FD1 \gpr_reg[31][6]  ( .D(n2361), .CP(clk), .Q(\gpr[31][6] ), .QN(n5025) );
  FD1 \gpr_reg[31][5]  ( .D(n2360), .CP(clk), .Q(\gpr[31][5] ), .QN(n5005) );
  FD1 \gpr_reg[31][4]  ( .D(n2359), .CP(clk), .Q(\gpr[31][4] ), .QN(n4974) );
  FD1 \gpr_reg[31][3]  ( .D(n2358), .CP(clk), .Q(\gpr[31][3] ), .QN(n4954) );
  FD1 \gpr_reg[31][2]  ( .D(n2357), .CP(clk), .Q(\gpr[31][2] ), .QN(n4930) );
  FD1 \gpr_reg[31][0]  ( .D(n2355), .CP(clk), .Q(\gpr[31][0] ), .QN(n4840) );
  FD1 \gpr_reg[12][2]  ( .D(n2965), .CP(clk), .Q(\gpr[12][2] ), .QN(n5680) );
  FD1 \gpr_reg[4][2]  ( .D(n3221), .CP(clk), .Q(\gpr[4][2] ), .QN(n5681) );
  FD1 \gpr_reg[5][0]  ( .D(n3187), .CP(clk), .Q(\gpr[5][0] ), .QN(n5669) );
  FD1 \gpr_reg[3][0]  ( .D(n3251), .CP(clk), .Q(\gpr[3][0] ), .QN(n5671) );
  FD1 \gpr_reg[1][0]  ( .D(n3315), .CP(clk), .Q(\gpr[1][0] ), .QN(n5670) );
  FD1 \gpr_reg[31][1]  ( .D(n2356), .CP(clk), .Q(\gpr[31][1] ), .QN(n5677) );
  FD1 \gpr_reg[27][1]  ( .D(n2484), .CP(clk), .Q(\gpr[27][1] ), .QN(n5678) );
  FD1 \gpr_reg[25][1]  ( .D(n2548), .CP(clk), .Q(\gpr[25][1] ), .QN(n5679) );
  FD1 \gpr_reg[22][1]  ( .D(n2644), .CP(clk), .Q(\gpr[22][1] ), .QN(n5674) );
  FD1 \gpr_reg[17][1]  ( .D(n2804), .CP(clk), .Q(\gpr[17][1] ), .QN(n5673) );
  FD1 \gpr_reg[16][1]  ( .D(n2836), .CP(clk), .Q(\gpr[16][1] ), .QN(n5672) );
  FD1 \gpr_reg[15][4]  ( .D(n2871), .CP(clk), .Q(\gpr[15][4] ), .QN(n5683) );
  FD1 \gpr_reg[14][4]  ( .D(n2903), .CP(clk), .Q(\gpr[14][4] ), .QN(n5686) );
  FD1 \gpr_reg[14][1]  ( .D(n2900), .CP(clk), .Q(\gpr[14][1] ), .QN(n4760) );
  FD1 \gpr_reg[13][4]  ( .D(n2935), .CP(clk), .Q(\gpr[13][4] ), .QN(n5682) );
  FD1 \gpr_reg[11][22]  ( .D(n3017), .CP(clk), .Q(\gpr[11][22] ), .QN(n5707)
         );
  FD1 \gpr_reg[11][12]  ( .D(n3007), .CP(clk), .Q(\gpr[11][12] ), .QN(n5695)
         );
  FD1 \gpr_reg[11][4]  ( .D(n2999), .CP(clk), .Q(\gpr[11][4] ), .QN(n5684) );
  FD1 \gpr_reg[9][22]  ( .D(n3081), .CP(clk), .Q(\gpr[9][22] ), .QN(n5708) );
  FD1 \gpr_reg[9][12]  ( .D(n3071), .CP(clk), .Q(\gpr[9][12] ), .QN(n5696) );
  FD1 \gpr_reg[9][4]  ( .D(n3063), .CP(clk), .Q(\gpr[9][4] ), .QN(n5685) );
  FD1 \gpr_reg[8][1]  ( .D(n3092), .CP(clk), .Q(\gpr[8][1] ), .QN(n5675) );
  FD1 \gpr_reg[7][22]  ( .D(n3145), .CP(clk), .Q(\gpr[7][22] ), .QN(n5709) );
  FD1 \gpr_reg[7][12]  ( .D(n3135), .CP(clk), .Q(\gpr[7][12] ), .QN(n5697) );
  FD1 \gpr_reg[7][4]  ( .D(n3127), .CP(clk), .Q(\gpr[7][4] ), .QN(n5687) );
  FD1 \gpr_reg[6][22]  ( .D(n3177), .CP(clk), .Q(\gpr[6][22] ), .QN(n5710) );
  FD1 \gpr_reg[6][12]  ( .D(n3167), .CP(clk), .Q(\gpr[6][12] ), .QN(n5698) );
  FD1 \gpr_reg[6][4]  ( .D(n3159), .CP(clk), .Q(\gpr[6][4] ), .QN(n5688) );
  FD1 \gpr_reg[5][22]  ( .D(n3209), .CP(clk), .Q(\gpr[5][22] ), .QN(n5711) );
  FD1 \gpr_reg[5][12]  ( .D(n3199), .CP(clk), .Q(\gpr[5][12] ), .QN(n5699) );
  FD1 \gpr_reg[5][4]  ( .D(n3191), .CP(clk), .Q(\gpr[5][4] ), .QN(n5689) );
  FD1 \gpr_reg[5][1]  ( .D(n3188), .CP(clk), .Q(\gpr[5][1] ), .QN(n5676) );
  FD1 \gpr_reg[3][22]  ( .D(n3273), .CP(clk), .Q(\gpr[3][22] ), .QN(n5713) );
  FD1 \gpr_reg[3][12]  ( .D(n3263), .CP(clk), .Q(\gpr[3][12] ), .QN(n5701) );
  FD1 \gpr_reg[3][4]  ( .D(n3255), .CP(clk), .Q(\gpr[3][4] ), .QN(n5691) );
  FD1 \gpr_reg[1][22]  ( .D(n3337), .CP(clk), .Q(\gpr[1][22] ), .QN(n5712) );
  FD1 \gpr_reg[1][12]  ( .D(n3327), .CP(clk), .Q(\gpr[1][12] ), .QN(n5700) );
  FD1 \gpr_reg[1][4]  ( .D(n3319), .CP(clk), .Q(\gpr[1][4] ), .QN(n5690) );
  FD1 \gpr_reg[16][15]  ( .D(n2850), .CP(clk), .Q(\gpr[16][15] ), .QN(n5702)
         );
  FD1 \gpr_reg[24][23]  ( .D(n2602), .CP(clk), .Q(\gpr[24][23] ), .QN(n5714)
         );
  FD1 \gpr_reg[24][19]  ( .D(n2598), .CP(clk), .Q(\gpr[24][19] ), .QN(n5705)
         );
  FD1 \gpr_reg[16][30]  ( .D(n2865), .CP(clk), .Q(\gpr[16][30] ), .QN(n5723)
         );
  FD1 \gpr_reg[14][17]  ( .D(n2916), .CP(clk), .Q(\gpr[14][17] ), .QN(n5703)
         );
  FD1 \gpr_reg[6][27]  ( .D(n3182), .CP(clk), .Q(\gpr[6][27] ), .QN(n5716) );
  FD1 \gpr_reg[3][27]  ( .D(n3278), .CP(clk), .Q(\gpr[3][27] ), .QN(n5718) );
  FD1 \gpr_reg[1][27]  ( .D(n3342), .CP(clk), .Q(\gpr[1][27] ), .QN(n5717) );
  FD1 \gpr_reg[12][26]  ( .D(n2989), .CP(clk), .Q(\gpr[12][26] ), .QN(n5715)
         );
  FD1 \gpr_reg[28][29]  ( .D(n2480), .CP(clk), .Q(\gpr[28][29] ), .QN(n5720)
         );
  FD1 \gpr_reg[25][29]  ( .D(n2576), .CP(clk), .Q(\gpr[25][29] ), .QN(n5721)
         );
  FD1 \gpr_reg[20][29]  ( .D(n2736), .CP(clk), .Q(\gpr[20][29] ), .QN(n5719)
         );
  FD1 \gpr_reg[6][11]  ( .D(n3166), .CP(clk), .Q(\gpr[6][11] ), .QN(n5692) );
  FD1 \gpr_reg[3][11]  ( .D(n3262), .CP(clk), .Q(\gpr[3][11] ), .QN(n5694) );
  FD1 \gpr_reg[1][11]  ( .D(n3326), .CP(clk), .Q(\gpr[1][11] ), .QN(n5693) );
  FD1 \gpr_reg[28][21]  ( .D(n2472), .CP(clk), .Q(\gpr[28][21] ), .QN(n5706)
         );
  FD1 \gpr_reg[5][11]  ( .D(n3198), .CP(clk), .Q(\gpr[5][11] ), .QN(n4761) );
  FD1 \gpr_reg[27][29]  ( .D(n2512), .CP(clk), .Q(\gpr[27][29] ), .QN(n5722)
         );
  FD1 \gpr_reg[4][18]  ( .D(n3237), .CP(clk), .Q(\gpr[4][18] ), .QN(n5704) );
  FD1 \gpr_reg[5][18]  ( .D(n3205), .CP(clk), .Q(\gpr[5][18] ), .QN(n4759) );
  AN2I U4 ( .A(n2), .B(n1), .Z(n2264) );
  IVI U5 ( .A(n2263), .Z(n1) );
  AN2I U6 ( .A(n2262), .B(n3), .Z(n2) );
  NR2I U7 ( .A(n2261), .B(n4), .Z(n3) );
  ND2I U8 ( .A(n2260), .B(n259), .Z(n4) );
  ND2I U9 ( .A(n7), .B(n5), .Z(n1710) );
  NR2I U10 ( .A(n1708), .B(n6), .Z(n5) );
  ND2I U11 ( .A(n172), .B(n1706), .Z(n6) );
  NR2I U12 ( .A(n12), .B(n8), .Z(n7) );
  ND2I U13 ( .A(n1707), .B(n9), .Z(n8) );
  AN2I U14 ( .A(n11), .B(n10), .Z(n9) );
  ND2I U15 ( .A(\gpr[24][21] ), .B(n1598), .Z(n10) );
  IVI U16 ( .A(n1063), .Z(n1598) );
  ND2I U17 ( .A(\gpr[25][21] ), .B(n1466), .Z(n11) );
  IVI U18 ( .A(n1275), .Z(n1466) );
  IVI U19 ( .A(n279), .Z(n12) );
  ND2I U20 ( .A(\gpr[2][28] ), .B(n13), .Z(n2321) );
  IVI U21 ( .A(n1148), .Z(n13) );
  ND2I U22 ( .A(n685), .B(n378), .Z(n1148) );
  NR2I U23 ( .A(n18), .B(n14), .Z(n2336) );
  ND2I U24 ( .A(n2304), .B(n15), .Z(n14) );
  AN2I U25 ( .A(n2305), .B(n16), .Z(n15) );
  IVI U26 ( .A(n17), .Z(n16) );
  ND2I U27 ( .A(n2309), .B(n2314), .Z(n17) );
  ND2I U28 ( .A(n20), .B(n19), .Z(n18) );
  ND2I U29 ( .A(n2303), .B(\gpr[4][28] ), .Z(n19) );
  IVI U30 ( .A(n21), .Z(n20) );
  ND2I U31 ( .A(n2316), .B(n22), .Z(n21) );
  AN2I U32 ( .A(n2310), .B(n2313), .Z(n22) );
  ND2I U33 ( .A(n4700), .B(n23), .Z(n4717) );
  IVI U34 ( .A(n24), .Z(n23) );
  ND2I U35 ( .A(n4698), .B(n25), .Z(n24) );
  AN2I U36 ( .A(n4699), .B(n26), .Z(n25) );
  AN2I U37 ( .A(n28), .B(n27), .Z(n26) );
  ND2I U38 ( .A(\gpr[31][25] ), .B(n2275), .Z(n27) );
  IVI U39 ( .A(n940), .Z(n2275) );
  ND2I U40 ( .A(\gpr[24][25] ), .B(n4686), .Z(n28) );
  IVI U41 ( .A(n1553), .Z(n4686) );
  AN2I U42 ( .A(n32), .B(n29), .Z(\rd_data1[26] ) );
  ND2I U43 ( .A(n31), .B(n30), .Z(n29) );
  NR2I U44 ( .A(n40), .B(n43), .Z(n30) );
  NR2I U45 ( .A(n39), .B(n1039), .Z(n31) );
  IVI U46 ( .A(n33), .Z(n32) );
  ND2I U47 ( .A(n35), .B(n34), .Z(n33) );
  ND2I U48 ( .A(n44), .B(n1017), .Z(n34) );
  ND2I U49 ( .A(n48), .B(n36), .Z(n35) );
  NR2I U50 ( .A(n38), .B(n37), .Z(n36) );
  ND2I U51 ( .A(n45), .B(n46), .Z(n37) );
  IVI U52 ( .A(n1005), .Z(n38) );
  ND2I U53 ( .A(n41), .B(n1026), .Z(n39) );
  IVI U54 ( .A(n1037), .Z(n40) );
  IVI U55 ( .A(n42), .Z(n41) );
  ND2I U56 ( .A(n1038), .B(n1020), .Z(n42) );
  ND4P U57 ( .A(n1019), .B(n1027), .C(n1018), .D(n498), .Z(n43) );
  AN2I U58 ( .A(n1015), .B(n1016), .Z(n44) );
  IVI U59 ( .A(n996), .Z(n45) );
  AN2I U60 ( .A(n1002), .B(n47), .Z(n46) );
  IVI U61 ( .A(n997), .Z(n47) );
  IVI U62 ( .A(n49), .Z(n48) );
  ND2I U63 ( .A(n1004), .B(n1003), .Z(n49) );
  IVI U64 ( .A(n50), .Z(n59) );
  ND2I U65 ( .A(n2301), .B(n51), .Z(n50) );
  IVI U66 ( .A(n52), .Z(n51) );
  ND2I U67 ( .A(n53), .B(n2293), .Z(n52) );
  IVI U68 ( .A(n54), .Z(n53) );
  ND2I U69 ( .A(n60), .B(n61), .Z(n54) );
  ND2I U70 ( .A(n58), .B(n55), .Z(n2302) );
  ND2I U71 ( .A(n2288), .B(n56), .Z(n55) );
  IVI U72 ( .A(n57), .Z(n56) );
  ND2I U73 ( .A(n260), .B(n2287), .Z(n57) );
  ND2I U74 ( .A(n62), .B(n59), .Z(n58) );
  ND2I U75 ( .A(\gpr[18][28] ), .B(n4702), .Z(n60) );
  ND2I U76 ( .A(\gpr[16][28] ), .B(n2296), .Z(n61) );
  AN2I U77 ( .A(n2294), .B(n63), .Z(n62) );
  IVI U78 ( .A(n2295), .Z(n63) );
  ND4P U79 ( .A(n908), .B(n907), .C(n498), .D(n64), .Z(n915) );
  ND2I U80 ( .A(n4719), .B(\gpr[1][22] ), .Z(n64) );
  ND2I U81 ( .A(n68), .B(n65), .Z(n70) );
  NR2I U82 ( .A(n67), .B(n66), .Z(n65) );
  ND2I U83 ( .A(n2123), .B(n71), .Z(n66) );
  ND2I U84 ( .A(n2121), .B(n80), .Z(n67) );
  IVI U85 ( .A(n69), .Z(n68) );
  ND2I U86 ( .A(n254), .B(n2139), .Z(n69) );
  ND2I U87 ( .A(n73), .B(n70), .Z(n74) );
  IVI U88 ( .A(n72), .Z(n71) );
  ND2I U89 ( .A(n2122), .B(n2124), .Z(n72) );
  AN2I U90 ( .A(n75), .B(n78), .Z(n73) );
  IVI U91 ( .A(n74), .Z(rd_data1[3]) );
  ND2I U92 ( .A(n2106), .B(n76), .Z(n75) );
  IVI U93 ( .A(n77), .Z(n76) );
  ND2I U94 ( .A(n2105), .B(n2107), .Z(n77) );
  ND2I U95 ( .A(n2089), .B(n79), .Z(n78) );
  NR2I U96 ( .A(n2088), .B(n2087), .Z(n79) );
  IVI U97 ( .A(n2140), .Z(n80) );
  IVI U98 ( .A(n81), .Z(rd_data1[5]) );
  AO3P U99 ( .A(n83), .B(n82), .C(n91), .D(n94), .Z(n81) );
  ND2I U100 ( .A(n86), .B(n84), .Z(n82) );
  ND2I U101 ( .A(n1628), .B(n90), .Z(n83) );
  IVI U102 ( .A(n85), .Z(n84) );
  ND2I U103 ( .A(n88), .B(n1627), .Z(n85) );
  NR2I U104 ( .A(n1614), .B(n87), .Z(n86) );
  ND2I U105 ( .A(n224), .B(n1613), .Z(n87) );
  IVI U106 ( .A(n89), .Z(n88) );
  ND2I U107 ( .A(n1611), .B(n1612), .Z(n89) );
  IVI U108 ( .A(n1617), .Z(n90) );
  ND2I U109 ( .A(n1605), .B(n92), .Z(n91) );
  IVI U110 ( .A(n93), .Z(n92) );
  ND2I U111 ( .A(n1603), .B(n1604), .Z(n93) );
  ND2I U112 ( .A(n1590), .B(n95), .Z(n94) );
  NR2I U113 ( .A(n1589), .B(n1588), .Z(n95) );
  B4IP U114 ( .A(rd_addr2[0]), .Z(n725) );
  ND2I U115 ( .A(n97), .B(n96), .Z(n722) );
  IVI U116 ( .A(n4442), .Z(n96) );
  IVI U117 ( .A(n3538), .Z(n97) );
  ND2I U118 ( .A(n724), .B(n98), .Z(n3538) );
  NR2I U119 ( .A(rd_addr2[0]), .B(n99), .Z(n98) );
  IVI U120 ( .A(rd_addr2[1]), .Z(n99) );
  ND2I U121 ( .A(n656), .B(n100), .Z(n119) );
  AN2I U122 ( .A(n657), .B(n658), .Z(n100) );
  ND4P U123 ( .A(n733), .B(n732), .C(n731), .D(n730), .Z(n741) );
  IVI U124 ( .A(n1915), .Z(n101) );
  IVI U125 ( .A(n1915), .Z(n102) );
  AO6P U126 ( .A(n105), .B(\gpr[6][4] ), .C(n178), .Z(n266) );
  ND4P U127 ( .A(n2086), .B(n2085), .C(n2084), .D(n2083), .Z(n2087) );
  ND2I U128 ( .A(n1077), .B(n2307), .Z(n103) );
  B4I U129 ( .A(n2297), .Z(n2215) );
  AN2I U130 ( .A(n1075), .B(n1204), .Z(n104) );
  AN2I U131 ( .A(n1075), .B(n1204), .Z(n105) );
  IVI U132 ( .A(n556), .Z(n106) );
  ND2I U133 ( .A(n110), .B(n107), .Z(n112) );
  NR2I U134 ( .A(n109), .B(n108), .Z(n107) );
  ND2I U135 ( .A(n233), .B(n683), .Z(n108) );
  ND2I U136 ( .A(n695), .B(n114), .Z(n109) );
  IVI U137 ( .A(n111), .Z(n110) );
  ND2I U138 ( .A(n696), .B(n113), .Z(n111) );
  ND2I U139 ( .A(n115), .B(n112), .Z(\rd_data1[31]_BAR ) );
  IVI U140 ( .A(n684), .Z(n113) );
  IVI U141 ( .A(n699), .Z(n114) );
  AN2I U142 ( .A(n119), .B(n116), .Z(n115) );
  ND2I U143 ( .A(n671), .B(n117), .Z(n116) );
  IVI U144 ( .A(n118), .Z(n117) );
  ND2I U145 ( .A(n669), .B(n670), .Z(n118) );
  ND2I U146 ( .A(n1319), .B(n120), .Z(n1327) );
  AN2I U147 ( .A(n122), .B(n121), .Z(n120) );
  ND2I U148 ( .A(n1983), .B(\gpr[10][2] ), .Z(n121) );
  IVI U149 ( .A(n123), .Z(n122) );
  ND2I U150 ( .A(n124), .B(n1318), .Z(n123) );
  IVI U151 ( .A(n1915), .Z(n1983) );
  ND2I U152 ( .A(\gpr[12][2] ), .B(n2132), .Z(n124) );
  ND4P U153 ( .A(n498), .B(n568), .C(n567), .D(n566), .Z(n569) );
  B5IP U154 ( .A(n594), .Z(n2094) );
  IVI U155 ( .A(n1136), .Z(n1268) );
  AO3 U156 ( .A(n2022), .B(n4841), .C(n2094), .D(n2021), .Z(n2023) );
  IVI U157 ( .A(n850), .Z(n2108) );
  AO3 U158 ( .A(n1007), .B(n4876), .C(n2094), .D(n1006), .Z(n1008) );
  AO3 U159 ( .A(n2022), .B(n4807), .C(n2094), .D(n819), .Z(n820) );
  AO2 U160 ( .A(n4704), .B(\gpr[23][8] ), .C(n1402), .D(\gpr[16][8] ), .Z(
        n1364) );
  ND4 U161 ( .A(n1236), .B(n1235), .C(n1234), .D(n1233), .Z(n1237) );
  ND4 U162 ( .A(n210), .B(n1544), .C(n1543), .D(n1542), .Z(n1581) );
  AO2 U163 ( .A(n4659), .B(\gpr[2][1] ), .C(n4657), .D(\gpr[3][1] ), .Z(n125)
         );
  AN4P U164 ( .A(n125), .B(n3422), .C(n3421), .D(n3432), .Z(n126) );
  ND4 U165 ( .A(n3413), .B(n3412), .C(n3411), .D(n3410), .Z(n127) );
  ND4 U166 ( .A(n3407), .B(n3406), .C(n3405), .D(n3404), .Z(n128) );
  ND2 U167 ( .A(n127), .B(n128), .Z(n129) );
  AO6P U168 ( .A(n126), .B(n3431), .C(n129), .Z(rd_data2[1]) );
  ND2I U169 ( .A(n4209), .B(\gpr[23][2] ), .Z(n130) );
  ND2I U170 ( .A(n130), .B(n4628), .Z(n131) );
  AO6 U171 ( .A(n4497), .B(\gpr[16][2] ), .C(n131), .Z(n3440) );
  ND2 U172 ( .A(\gpr[24][10] ), .B(n4637), .Z(n132) );
  ND2 U173 ( .A(\gpr[25][10] ), .B(n4001), .Z(n133) );
  ND2 U174 ( .A(n132), .B(n133), .Z(n134) );
  NR2I U175 ( .A(n802), .B(n134), .Z(n803) );
  ND2I U176 ( .A(n4548), .B(\gpr[23][15] ), .Z(n135) );
  ND2I U177 ( .A(n135), .B(n4628), .Z(n136) );
  AO6 U178 ( .A(n4432), .B(\gpr[16][15] ), .C(n136), .Z(n3939) );
  AO2 U179 ( .A(\gpr[17][30] ), .B(n4636), .C(n4623), .D(\gpr[19][30] ), .Z(
        n4552) );
  AO2 U180 ( .A(\gpr[26][28] ), .B(n4622), .C(n4623), .D(\gpr[27][28] ), .Z(
        n4454) );
  ND2I U181 ( .A(n4548), .B(\gpr[23][30] ), .Z(n137) );
  ND2I U182 ( .A(n137), .B(n4628), .Z(n138) );
  AO6 U183 ( .A(n4549), .B(\gpr[16][30] ), .C(n138), .Z(n4550) );
  AO2 U184 ( .A(n4623), .B(\gpr[19][31] ), .C(\gpr[18][31] ), .D(n4622), .Z(
        n4634) );
  ND2 U185 ( .A(n4543), .B(\gpr[31][30] ), .Z(n139) );
  ND2I U186 ( .A(n139), .B(n4641), .Z(n140) );
  AO6 U187 ( .A(n4624), .B(\gpr[28][30] ), .C(n140), .Z(n4544) );
  AO2 U188 ( .A(n4624), .B(\gpr[28][28] ), .C(\gpr[24][28] ), .D(n4450), .Z(
        n141) );
  ND4P U189 ( .A(n141), .B(n4456), .C(n4455), .D(n4454), .Z(n4463) );
  ND2 U190 ( .A(n4251), .B(\gpr[31][10] ), .Z(n142) );
  ND2I U191 ( .A(n142), .B(n4641), .Z(n143) );
  AO6 U192 ( .A(n4501), .B(\gpr[27][10] ), .C(n143), .Z(n804) );
  AO2 U193 ( .A(n4623), .B(\gpr[27][30] ), .C(\gpr[25][30] ), .D(n4636), .Z(
        n4546) );
  ND2I U194 ( .A(n4624), .B(\gpr[28][25] ), .Z(n144) );
  ND3P U195 ( .A(n4340), .B(n4341), .C(n144), .Z(n145) );
  AO1P U196 ( .A(\gpr[30][25] ), .B(n4431), .C(n4344), .D(n145), .Z(n146) );
  AO2 U197 ( .A(\gpr[24][25] ), .B(n4637), .C(\gpr[25][25] ), .D(n4636), .Z(
        n147) );
  ND2I U198 ( .A(n146), .B(n147), .Z(n4345) );
  AO3 U199 ( .A(n4687), .B(n4844), .C(n1582), .D(n2094), .Z(n1589) );
  ND2 U200 ( .A(n4650), .B(n4801), .Z(n148) );
  AO3 U201 ( .A(\gpr[15][27] ), .B(n4639), .C(n4652), .D(n148), .Z(n149) );
  ND2I U202 ( .A(n149), .B(n4561), .Z(n150) );
  AO6 U203 ( .A(n4524), .B(\gpr[6][27] ), .C(n150), .Z(n4446) );
  ND2I U204 ( .A(n2157), .B(\gpr[29][18] ), .Z(n151) );
  ND3P U205 ( .A(n534), .B(n533), .C(n151), .Z(n535) );
  ND2I U206 ( .A(n2020), .B(\gpr[22][21] ), .Z(n152) );
  ND2 U207 ( .A(n152), .B(n2094), .Z(n153) );
  AO6 U208 ( .A(n2204), .B(\gpr[20][21] ), .C(n153), .Z(n277) );
  AO2 U209 ( .A(n4636), .B(\gpr[17][28] ), .C(n4457), .D(\gpr[23][28] ), .Z(
        n154) );
  ND4 U210 ( .A(n4628), .B(n293), .C(n4461), .D(n154), .Z(n4462) );
  AO2 U211 ( .A(n4623), .B(\gpr[27][27] ), .C(\gpr[25][27] ), .D(n4636), .Z(
        n4423) );
  ND4P U212 ( .A(n4309), .B(n4310), .C(n4311), .D(n4312), .Z(n155) );
  AO3 U213 ( .A(n4775), .B(n3446), .C(n4561), .D(n4307), .Z(n156) );
  NR2I U214 ( .A(n155), .B(n156), .Z(n4329) );
  ND2I U215 ( .A(n4548), .B(\gpr[31][23] ), .Z(n157) );
  ND2I U216 ( .A(n157), .B(n4453), .Z(n158) );
  AO6 U217 ( .A(n4497), .B(\gpr[24][23] ), .C(n158), .Z(n4247) );
  AO4 U218 ( .A(n484), .B(n4985), .C(n1507), .D(n4984), .Z(n597) );
  NR2I U219 ( .A(n4776), .B(n2006), .Z(n159) );
  NR2 U220 ( .A(n5477), .B(n1546), .Z(n160) );
  NR2I U221 ( .A(n159), .B(n160), .Z(n161) );
  ND2I U222 ( .A(n2094), .B(n161), .Z(n1547) );
  IVI U223 ( .A(wr_data[17]), .Z(n4000) );
  AO2 U224 ( .A(n4268), .B(\gpr[10][4] ), .C(n4659), .D(\gpr[2][4] ), .Z(n162)
         );
  AO2 U225 ( .A(n4666), .B(\gpr[4][4] ), .C(n3558), .D(\gpr[9][4] ), .Z(n163)
         );
  ND2I U226 ( .A(n162), .B(n163), .Z(n3559) );
  ND4P U227 ( .A(n3455), .B(n3456), .C(n3457), .D(n3458), .Z(n164) );
  ND4 U228 ( .A(n3459), .B(n3460), .C(n3461), .D(n3462), .Z(n165) );
  NR2I U229 ( .A(n164), .B(n165), .Z(n3463) );
  ND2I U230 ( .A(n4209), .B(\gpr[23][22] ), .Z(n166) );
  ND2I U231 ( .A(n166), .B(n4628), .Z(n167) );
  AO6 U232 ( .A(n4497), .B(\gpr[16][22] ), .C(n167), .Z(n4210) );
  ND4P U233 ( .A(n4154), .B(n4155), .C(n4156), .D(n4157), .Z(n168) );
  AO3 U234 ( .A(n4774), .B(n4150), .C(n4561), .D(n4152), .Z(n169) );
  NR2I U235 ( .A(n168), .B(n169), .Z(n4168) );
  AO2 U236 ( .A(n4333), .B(\gpr[31][18] ), .C(n4090), .D(\gpr[29][18] ), .Z(
        n170) );
  AO2 U237 ( .A(n4635), .B(\gpr[27][18] ), .C(n4214), .D(\gpr[26][18] ), .Z(
        n171) );
  ND4P U238 ( .A(n4058), .B(n4059), .C(n170), .D(n171), .Z(n4069) );
  EO1 U239 ( .A(n1367), .B(\gpr[14][20] ), .C(n5724), .D(n1136), .Z(n1137) );
  ND2I U240 ( .A(n2207), .B(\gpr[26][21] ), .Z(n172) );
  ND3 U241 ( .A(n2292), .B(n2307), .C(\gpr[13][26] ), .Z(n1020) );
  ND2I U242 ( .A(\gpr[18][7] ), .B(n2077), .Z(n173) );
  ND2I U243 ( .A(\gpr[16][7] ), .B(n1598), .Z(n174) );
  ND2I U244 ( .A(n173), .B(n174), .Z(n175) );
  NR3P U245 ( .A(n1062), .B(n1061), .C(n175), .Z(n1064) );
  ND2I U246 ( .A(\gpr[7][4] ), .B(n2061), .Z(n176) );
  ND2I U247 ( .A(\gpr[11][4] ), .B(n4739), .Z(n177) );
  ND2I U248 ( .A(n176), .B(n177), .Z(n178) );
  IVI U249 ( .A(wr_data[29]), .Z(n4486) );
  ND2 U250 ( .A(n226), .B(n2194), .Z(n179) );
  ND4P U251 ( .A(n2195), .B(n2196), .C(n2198), .D(n2199), .Z(n180) );
  NR2I U252 ( .A(n179), .B(n180), .Z(n2200) );
  AO2 U253 ( .A(n4623), .B(\gpr[19][29] ), .C(\gpr[20][29] ), .D(n4624), .Z(
        n4495) );
  AO2 U254 ( .A(n4474), .B(\gpr[9][28] ), .C(\gpr[8][28] ), .D(n4570), .Z(n181) );
  AO2 U255 ( .A(\gpr[10][28] ), .B(n4473), .C(\gpr[2][28] ), .D(n4659), .Z(
        n182) );
  ND2I U256 ( .A(n181), .B(n182), .Z(n4481) );
  ND2I U257 ( .A(n4457), .B(\gpr[31][27] ), .Z(n183) );
  ND2I U258 ( .A(n183), .B(n4453), .Z(n184) );
  AO6 U259 ( .A(n4498), .B(\gpr[28][27] ), .C(n184), .Z(n4421) );
  ND2I U260 ( .A(n4625), .B(\gpr[22][21] ), .Z(n185) );
  ND2I U261 ( .A(n185), .B(n4628), .Z(n186) );
  AO6 U262 ( .A(n4549), .B(\gpr[16][21] ), .C(n186), .Z(n4178) );
  ND2 U263 ( .A(n4184), .B(n4791), .Z(n187) );
  AO3 U264 ( .A(\gpr[15][18] ), .B(n4090), .C(n4652), .D(n187), .Z(n188) );
  ND2I U265 ( .A(n188), .B(n4561), .Z(n189) );
  AO6 U266 ( .A(n4475), .B(\gpr[6][18] ), .C(n189), .Z(n4086) );
  ND3 U267 ( .A(RegWrite), .B(n3348), .C(wr_addr[3]), .Z(n3356) );
  AO2 U268 ( .A(\gpr[6][0] ), .B(n105), .C(n1523), .D(\gpr[15][0] ), .Z(n190)
         );
  AO2 U269 ( .A(\gpr[7][0] ), .B(n4747), .C(\gpr[14][0] ), .D(n4748), .Z(n191)
         );
  ND2I U270 ( .A(n190), .B(n191), .Z(n360) );
  ND2I U271 ( .A(n2233), .B(\gpr[24][29] ), .Z(n192) );
  ND2I U272 ( .A(\gpr[26][29] ), .B(n2077), .Z(n193) );
  ND2I U273 ( .A(n192), .B(n193), .Z(n2234) );
  ND3 U274 ( .A(n2157), .B(n2037), .C(\gpr[5][1] ), .Z(n2039) );
  AO3 U275 ( .A(n2092), .B(n4805), .C(n2094), .D(n595), .Z(n194) );
  NR2I U276 ( .A(n597), .B(n194), .Z(n598) );
  IVI U277 ( .A(wr_data[4]), .Z(n3537) );
  AO2 U278 ( .A(n4572), .B(\gpr[15][4] ), .C(\gpr[12][4] ), .D(n4573), .Z(n195) );
  AO2 U279 ( .A(n4571), .B(\gpr[11][4] ), .C(\gpr[8][4] ), .D(n3960), .Z(n196)
         );
  ND2I U280 ( .A(n195), .B(n196), .Z(n3568) );
  ND4P U281 ( .A(n4159), .B(n4160), .C(n4161), .D(n4162), .Z(n197) );
  ND4 U282 ( .A(n4163), .B(n4164), .C(n4165), .D(n4166), .Z(n198) );
  NR2I U283 ( .A(n197), .B(n198), .Z(n4167) );
  ND2I U284 ( .A(\gpr[30][19] ), .B(n4625), .Z(n199) );
  ND2I U285 ( .A(n199), .B(n4453), .Z(n200) );
  AO6 U286 ( .A(n4357), .B(\gpr[24][19] ), .C(n200), .Z(n4098) );
  AO2 U287 ( .A(n4475), .B(\gpr[6][17] ), .C(\gpr[7][17] ), .D(n4675), .Z(n201) );
  AO2 U288 ( .A(n4666), .B(\gpr[4][17] ), .C(\gpr[1][17] ), .D(n4556), .Z(n202) );
  ND2I U289 ( .A(n201), .B(n202), .Z(n4023) );
  ND2I U290 ( .A(\gpr[23][9] ), .B(n4209), .Z(n203) );
  ND2I U291 ( .A(n203), .B(n4628), .Z(n204) );
  AO6 U292 ( .A(n4623), .B(\gpr[19][9] ), .C(n204), .Z(n3743) );
  ND2 U293 ( .A(\gpr[23][10] ), .B(n3864), .Z(n205) );
  ND3 U294 ( .A(n805), .B(n4628), .C(n205), .Z(n234) );
  ND3 U295 ( .A(wr_addr[1]), .B(n2344), .C(wr_addr[0]), .Z(n3353) );
  AO2 U296 ( .A(n1583), .B(\gpr[16][14] ), .C(\gpr[19][14] ), .D(n4703), .Z(
        n1233) );
  ND3 U297 ( .A(n2307), .B(n206), .C(\gpr[9][11] ), .Z(n1796) );
  AO2 U298 ( .A(\gpr[26][11] ), .B(n4726), .C(n2292), .D(\gpr[29][11] ), .Z(
        n1774) );
  AO2 U299 ( .A(\gpr[7][24] ), .B(n2306), .C(\gpr[6][24] ), .D(n105), .Z(n1544) );
  AO2 U300 ( .A(n4666), .B(\gpr[4][0] ), .C(\gpr[7][0] ), .D(n4675), .Z(n3392)
         );
  EO1 U301 ( .A(n4604), .B(n4246), .C(\gpr[28][23] ), .D(n4604), .Z(n2474) );
  EO1 U302 ( .A(n4591), .B(n4246), .C(\gpr[20][23] ), .D(n4591), .Z(n2730) );
  EO1 U303 ( .A(n4607), .B(n4129), .C(\gpr[8][20] ), .D(n4607), .Z(n3111) );
  EO1 U304 ( .A(n4618), .B(n4412), .C(\gpr[5][27] ), .D(n4618), .Z(n3214) );
  EO1 U305 ( .A(n4614), .B(n4371), .C(\gpr[4][26] ), .D(n4614), .Z(n3245) );
  IVI U306 ( .A(n659), .Z(n206) );
  IVDA U307 ( .A(n1546), .Y(n207), .Z(n2050) );
  AN2I U308 ( .A(n485), .B(n264), .Z(n209) );
  AN2I U309 ( .A(n244), .B(n1526), .Z(n210) );
  AN2I U310 ( .A(n1210), .B(n1209), .Z(n211) );
  AN4P U311 ( .A(n2174), .B(n1431), .C(n1430), .D(n1429), .Z(n212) );
  AN2I U312 ( .A(n1609), .B(n2174), .Z(n213) );
  AN2I U313 ( .A(n1640), .B(n1639), .Z(n214) );
  AN2I U314 ( .A(n1780), .B(n2174), .Z(n215) );
  AN2I U315 ( .A(n1819), .B(n282), .Z(n216) );
  AN2I U316 ( .A(n1971), .B(n2174), .Z(n217) );
  AN2I U317 ( .A(n2134), .B(n2174), .Z(n218) );
  AN2I U318 ( .A(n487), .B(n486), .Z(n221) );
  AN2I U319 ( .A(n505), .B(n504), .Z(n222) );
  AN2I U320 ( .A(n1537), .B(n1536), .Z(n223) );
  AN2I U321 ( .A(n213), .B(n1610), .Z(n224) );
  AN2I U322 ( .A(n1861), .B(n1860), .Z(n225) );
  AN2I U323 ( .A(n2193), .B(n2192), .Z(n226) );
  AN2I U324 ( .A(n386), .B(n385), .Z(n227) );
  ND2I U325 ( .A(n396), .B(n395), .Z(n228) );
  AN2I U326 ( .A(n433), .B(n432), .Z(n229) );
  AN2I U327 ( .A(n454), .B(n453), .Z(n230) );
  AN2I U328 ( .A(n555), .B(n554), .Z(n231) );
  AN2I U329 ( .A(n638), .B(n637), .Z(n232) );
  AN2I U330 ( .A(n679), .B(n678), .Z(n233) );
  AN2I U331 ( .A(n4723), .B(\gpr[5][30] ), .Z(n235) );
  AN2I U332 ( .A(n1070), .B(n1069), .Z(n236) );
  AN2I U333 ( .A(n1203), .B(n1202), .Z(n237) );
  AN2I U334 ( .A(n1223), .B(n1222), .Z(n238) );
  AN2I U335 ( .A(n1314), .B(n1313), .Z(n239) );
  AN2I U336 ( .A(n1444), .B(n1443), .Z(n240) );
  AN2I U337 ( .A(n1428), .B(n1427), .Z(n241) );
  AN2I U338 ( .A(n1473), .B(n1472), .Z(n242) );
  AN2I U339 ( .A(n1485), .B(n1484), .Z(n243) );
  AN2I U340 ( .A(n1522), .B(n1521), .Z(n244) );
  ND2I U341 ( .A(n1555), .B(n1554), .Z(n245) );
  AN2I U342 ( .A(n1636), .B(n1635), .Z(n246) );
  AN2I U343 ( .A(n1646), .B(n1645), .Z(n247) );
  AN2I U344 ( .A(\gpr[4][21] ), .B(n4732), .Z(n248) );
  AN2I U345 ( .A(n1711), .B(n1710), .Z(n249) );
  AN2I U346 ( .A(n1805), .B(n1804), .Z(n250) );
  AN2I U347 ( .A(n1845), .B(n1844), .Z(n251) );
  AN2I U348 ( .A(n4723), .B(\gpr[5][9] ), .Z(n252) );
  AN2I U349 ( .A(\gpr[15][3] ), .B(n2312), .Z(n253) );
  AN2I U350 ( .A(n2131), .B(n2130), .Z(n254) );
  AN2I U351 ( .A(n2152), .B(n2151), .Z(n255) );
  AN2I U352 ( .A(n2166), .B(n2165), .Z(n256) );
  AN2I U353 ( .A(n2230), .B(n2229), .Z(n257) );
  AN2I U354 ( .A(n2303), .B(\gpr[4][29] ), .Z(n258) );
  AN2I U355 ( .A(n2258), .B(n2257), .Z(n259) );
  AN2I U356 ( .A(n2286), .B(n2285), .Z(n260) );
  B4IP U357 ( .A(n779), .Z(n4652) );
  B4IP U358 ( .A(n3414), .Z(n4675) );
  B2I U359 ( .A(n4473), .Z2(n3679) );
  AN2I U360 ( .A(n4690), .B(n350), .Z(n261) );
  AN2I U361 ( .A(n1498), .B(n2174), .Z(n262) );
  AN2I U362 ( .A(\gpr[14][12] ), .B(n2252), .Z(n263) );
  OR2P U363 ( .A(n2092), .B(n4873), .Z(n264) );
  AN2I U364 ( .A(n622), .B(n498), .Z(n265) );
  AN2I U365 ( .A(n859), .B(n858), .Z(n267) );
  AN2I U366 ( .A(n498), .B(n966), .Z(n268) );
  AN2I U367 ( .A(n1021), .B(n2292), .Z(n269) );
  AN2I U368 ( .A(n1078), .B(n2174), .Z(n270) );
  AN2I U369 ( .A(n2252), .B(\gpr[14][7] ), .Z(n271) );
  OR2P U370 ( .A(n1889), .B(n4861), .Z(n272) );
  AN2I U371 ( .A(n4690), .B(n1196), .Z(n273) );
  AN2I U372 ( .A(n1386), .B(n1385), .Z(n274) );
  AN2I U373 ( .A(n1420), .B(n1419), .Z(n275) );
  AN2I U374 ( .A(n1649), .B(n1648), .Z(n276) );
  OR2P U375 ( .A(n1889), .B(n4869), .Z(n278) );
  AN2I U376 ( .A(n4690), .B(n1709), .Z(n279) );
  AN2I U377 ( .A(n1990), .B(\gpr[14][11] ), .Z(n280) );
  OR2P U378 ( .A(n1810), .B(n4866), .Z(n281) );
  AN2I U379 ( .A(n4690), .B(n1818), .Z(n282) );
  OR2P U380 ( .A(n1889), .B(n4859), .Z(n283) );
  AN2I U381 ( .A(n4690), .B(n1901), .Z(n284) );
  AN2I U382 ( .A(n1905), .B(n2174), .Z(n285) );
  OR2P U383 ( .A(n1765), .B(n4851), .Z(n286) );
  AN2I U384 ( .A(n4690), .B(n1950), .Z(n287) );
  AN2I U385 ( .A(\gpr[19][17] ), .B(n4703), .Z(n288) );
  AN2I U386 ( .A(n4690), .B(n2154), .Z(n289) );
  OR2P U387 ( .A(n2159), .B(n4864), .Z(n290) );
  OR2P U388 ( .A(n1889), .B(n4810), .Z(n291) );
  AN2I U389 ( .A(\gpr[15][29] ), .B(n2312), .Z(n292) );
  AN2I U390 ( .A(n4460), .B(n4459), .Z(n293) );
  B2IP U391 ( .A(n702), .Z1(n294), .Z2(n295) );
  AN2I U392 ( .A(n2037), .B(\gpr[5][11] ), .Z(n296) );
  AN2I U393 ( .A(n4725), .B(\gpr[10][25] ), .Z(n297) );
  AN2I U394 ( .A(rd_addr1[2]), .B(rd_addr1[1]), .Z(n357) );
  IVI U395 ( .A(rd_addr1[0]), .Z(n356) );
  ND2I U396 ( .A(n357), .B(n356), .Z(n525) );
  IVI U397 ( .A(n525), .Z(n1204) );
  IVI U398 ( .A(n1204), .Z(n1810) );
  NR2I U399 ( .A(n1810), .B(n4762), .Z(n321) );
  IVI U400 ( .A(rd_addr1[3]), .Z(n685) );
  ND2I U401 ( .A(rd_addr1[4]), .B(n685), .Z(n594) );
  IVI U402 ( .A(n594), .Z(n4709) );
  NR2I U403 ( .A(rd_addr1[2]), .B(rd_addr1[1]), .Z(n333) );
  ND2I U404 ( .A(n333), .B(rd_addr1[0]), .Z(n383) );
  IVI U405 ( .A(n383), .Z(n601) );
  IVI U406 ( .A(n601), .Z(n1252) );
  ND2I U407 ( .A(n1938), .B(\gpr[17][0] ), .Z(n319) );
  ND2I U408 ( .A(n4709), .B(n319), .Z(n320) );
  NR2I U409 ( .A(n321), .B(n320), .Z(n339) );
  IVI U410 ( .A(rd_addr1[1]), .Z(n322) );
  AN2I U411 ( .A(rd_addr1[2]), .B(n322), .Z(n361) );
  ND2I U412 ( .A(rd_addr1[0]), .B(n361), .Z(n1545) );
  ND2I U413 ( .A(\gpr[21][0] ), .B(n2292), .Z(n325) );
  NR2I U414 ( .A(rd_addr1[0]), .B(rd_addr1[2]), .Z(n323) );
  AN2I U415 ( .A(rd_addr1[1]), .B(n323), .Z(n378) );
  IVI U416 ( .A(n378), .Z(n596) );
  B4I U417 ( .A(n596), .Z(n2077) );
  ND2I U418 ( .A(\gpr[18][0] ), .B(n2077), .Z(n324) );
  AN2I U419 ( .A(n325), .B(n324), .Z(n328) );
  ND2I U420 ( .A(n361), .B(n356), .Z(n326) );
  B4IP U421 ( .A(n326), .Z(n1631) );
  ND2I U422 ( .A(\gpr[20][0] ), .B(n2204), .Z(n327) );
  ND2I U423 ( .A(n328), .B(n327), .Z(n337) );
  AN2I U424 ( .A(n357), .B(rd_addr1[0]), .Z(n576) );
  IVI U425 ( .A(n576), .Z(n940) );
  B5IP U426 ( .A(n940), .Z(n4704) );
  ND2I U427 ( .A(\gpr[23][0] ), .B(n4704), .Z(n332) );
  IVI U428 ( .A(rd_addr1[2]), .Z(n330) );
  AN2I U429 ( .A(rd_addr1[1]), .B(rd_addr1[0]), .Z(n329) );
  ND2I U430 ( .A(n330), .B(n329), .Z(n362) );
  IVI U431 ( .A(n362), .Z(n503) );
  IVI U432 ( .A(n503), .Z(n467) );
  B5IP U433 ( .A(n467), .Z(n2284) );
  ND2I U434 ( .A(\gpr[19][0] ), .B(n2284), .Z(n331) );
  AN2I U435 ( .A(n332), .B(n331), .Z(n335) );
  ND2I U436 ( .A(n333), .B(n356), .Z(n1136) );
  IVI U437 ( .A(n1268), .Z(n1363) );
  IVI U438 ( .A(n1363), .Z(n2004) );
  ND2I U439 ( .A(\gpr[16][0] ), .B(n2004), .Z(n334) );
  ND2I U440 ( .A(n335), .B(n334), .Z(n336) );
  NR2I U441 ( .A(n337), .B(n336), .Z(n338) );
  ND2I U442 ( .A(n339), .B(n338), .Z(n355) );
  ND2I U443 ( .A(\gpr[29][0] ), .B(n4701), .Z(n340) );
  IVI U444 ( .A(n340), .Z(n344) );
  IVI U445 ( .A(n378), .Z(n484) );
  B4IP U446 ( .A(n596), .Z(n4702) );
  ND2I U447 ( .A(\gpr[26][0] ), .B(n2077), .Z(n342) );
  IVI U448 ( .A(n1268), .Z(n934) );
  IVI U449 ( .A(n934), .Z(n1205) );
  ND2I U450 ( .A(\gpr[24][0] ), .B(n1205), .Z(n341) );
  ND2I U451 ( .A(n342), .B(n341), .Z(n343) );
  NR2I U452 ( .A(n344), .B(n343), .Z(n353) );
  ND2I U453 ( .A(n2158), .B(\gpr[28][0] ), .Z(n346) );
  ND2I U454 ( .A(n357), .B(n356), .Z(n1546) );
  ND2I U455 ( .A(\gpr[30][0] ), .B(n862), .Z(n345) );
  AN2I U456 ( .A(n346), .B(n345), .Z(n352) );
  IVI U457 ( .A(n576), .Z(n2297) );
  NR2I U458 ( .A(n2297), .B(n4840), .Z(n347) );
  IVI U459 ( .A(n347), .Z(n349) );
  ND2I U460 ( .A(\gpr[25][0] ), .B(n1824), .Z(n348) );
  AN2I U461 ( .A(n349), .B(n348), .Z(n351) );
  ND2I U462 ( .A(rd_addr1[4]), .B(n4725), .Z(n401) );
  IVI U463 ( .A(n401), .Z(n4690) );
  IVI U464 ( .A(n362), .Z(n4688) );
  ND2I U465 ( .A(n4688), .B(\gpr[27][0] ), .Z(n350) );
  ND4P U466 ( .A(n353), .B(n352), .C(n351), .D(n261), .Z(n354) );
  AN2I U467 ( .A(n355), .B(n354), .Z(n392) );
  ND2I U468 ( .A(n576), .B(n4725), .Z(n1432) );
  IVI U469 ( .A(n1432), .Z(n1523) );
  ND2I U470 ( .A(n576), .B(n685), .Z(n2173) );
  IVI U471 ( .A(n2173), .Z(n4747) );
  ND2I U472 ( .A(n357), .B(n356), .Z(n492) );
  IVI U473 ( .A(n492), .Z(n862) );
  ND2I U474 ( .A(n4725), .B(n862), .Z(n1606) );
  ND2I U475 ( .A(n1631), .B(n685), .Z(n850) );
  B2IP U476 ( .A(n2108), .Z2(n4732) );
  ND2I U477 ( .A(n4732), .B(\gpr[4][0] ), .Z(n358) );
  IVI U478 ( .A(n358), .Z(n359) );
  NR2I U479 ( .A(n360), .B(n359), .Z(n390) );
  B2IP U480 ( .A(rd_addr1[3]), .Z1(n2037), .Z2(n4725) );
  ND2I U481 ( .A(rd_addr1[0]), .B(n361), .Z(n1469) );
  ND2I U482 ( .A(n2037), .B(n1752), .Z(n562) );
  B4IP U483 ( .A(n562), .Z(n4723) );
  ND2I U484 ( .A(n4723), .B(\gpr[5][0] ), .Z(n369) );
  IVI U485 ( .A(n362), .Z(n1077) );
  ND2I U486 ( .A(n685), .B(n1077), .Z(n1434) );
  ND2I U487 ( .A(n2110), .B(\gpr[3][0] ), .Z(n367) );
  ND2I U488 ( .A(n4725), .B(n1631), .Z(n556) );
  IVI U489 ( .A(n556), .Z(n2132) );
  ND2I U490 ( .A(n2132), .B(\gpr[12][0] ), .Z(n364) );
  B2IP U491 ( .A(rd_addr1[3]), .Z1(n1075), .Z2(n2307) );
  ND2I U492 ( .A(n1077), .B(n2307), .Z(n1308) );
  IVI U493 ( .A(n1308), .Z(n1970) );
  ND2I U494 ( .A(n1970), .B(\gpr[11][0] ), .Z(n363) );
  ND2I U495 ( .A(n364), .B(n363), .Z(n365) );
  IVI U496 ( .A(n365), .Z(n366) );
  AN2I U497 ( .A(n367), .B(n366), .Z(n368) );
  ND2I U498 ( .A(n369), .B(n368), .Z(n377) );
  IVI U499 ( .A(n601), .Z(n659) );
  IVI U500 ( .A(n659), .Z(n370) );
  ND2I U501 ( .A(n2307), .B(n370), .Z(n1320) );
  IVI U502 ( .A(n1320), .Z(n2125) );
  ND2I U503 ( .A(n2125), .B(\gpr[9][0] ), .Z(n375) );
  IVI U504 ( .A(n1136), .Z(n2048) );
  AN2I U505 ( .A(n4725), .B(n2048), .Z(n672) );
  IVI U506 ( .A(n672), .Z(n2239) );
  IVI U507 ( .A(n2239), .Z(n4738) );
  ND2I U508 ( .A(n4738), .B(\gpr[8][0] ), .Z(n372) );
  IVI U509 ( .A(n484), .Z(n1535) );
  ND2I U510 ( .A(n4725), .B(n1535), .Z(n1915) );
  ND2I U511 ( .A(n1983), .B(\gpr[10][0] ), .Z(n371) );
  ND2I U512 ( .A(n372), .B(n371), .Z(n373) );
  IVI U513 ( .A(n373), .Z(n374) );
  ND2I U514 ( .A(n375), .B(n374), .Z(n376) );
  NR2I U515 ( .A(n377), .B(n376), .Z(n387) );
  ND2I U516 ( .A(n1752), .B(n2307), .Z(n1083) );
  IVI U517 ( .A(n1083), .Z(n2188) );
  ND2I U518 ( .A(\gpr[13][0] ), .B(n2188), .Z(n381) );
  IVI U519 ( .A(n1148), .Z(n2115) );
  ND2I U520 ( .A(n2115), .B(\gpr[2][0] ), .Z(n379) );
  IVI U521 ( .A(rd_addr1[4]), .Z(n2174) );
  AN2I U522 ( .A(n379), .B(n2174), .Z(n380) );
  ND2I U523 ( .A(n381), .B(n380), .Z(n382) );
  IVI U524 ( .A(n382), .Z(n386) );
  IVI U525 ( .A(n383), .Z(n384) );
  AN2I U526 ( .A(n384), .B(n685), .Z(n2320) );
  B2IP U527 ( .A(n2320), .Z2(n4719) );
  ND2I U528 ( .A(\gpr[1][0] ), .B(n4719), .Z(n385) );
  ND2I U529 ( .A(n387), .B(n227), .Z(n388) );
  IVI U530 ( .A(n388), .Z(n389) );
  ND2I U531 ( .A(n390), .B(n389), .Z(n391) );
  ND2I U532 ( .A(n392), .B(n391), .Z(n393) );
  IVI U533 ( .A(n393), .Z(rd_data1[0]) );
  IVI U534 ( .A(n1252), .Z(n2276) );
  ND2I U535 ( .A(\gpr[25][12] ), .B(n2276), .Z(n396) );
  IVI U536 ( .A(n503), .Z(n394) );
  B4IP U537 ( .A(n394), .Z(n4703) );
  ND2I U538 ( .A(\gpr[27][12] ), .B(n4703), .Z(n395) );
  IVI U539 ( .A(n576), .Z(n397) );
  B4IP U540 ( .A(n397), .Z(n2100) );
  ND2I U541 ( .A(n2100), .B(\gpr[31][12] ), .Z(n399) );
  IVI U542 ( .A(n1631), .Z(n413) );
  ND2I U543 ( .A(\gpr[28][12] ), .B(n2204), .Z(n398) );
  ND2I U544 ( .A(n399), .B(n398), .Z(n400) );
  NR2I U545 ( .A(n228), .B(n400), .Z(n409) );
  IVI U546 ( .A(n1204), .Z(n1889) );
  NR2I U547 ( .A(n1889), .B(n4857), .Z(n404) );
  IVI U548 ( .A(n401), .Z(n2079) );
  IVI U549 ( .A(n1268), .Z(n1507) );
  IVI U550 ( .A(n1507), .Z(n878) );
  ND2I U551 ( .A(n878), .B(\gpr[24][12] ), .Z(n402) );
  ND2I U552 ( .A(n2079), .B(n402), .Z(n403) );
  NR2I U553 ( .A(n404), .B(n403), .Z(n406) );
  B4I U554 ( .A(n484), .Z(n4726) );
  AO2P U555 ( .A(n4726), .B(\gpr[26][12] ), .C(n4701), .D(\gpr[29][12] ), .Z(
        n405) );
  ND2I U556 ( .A(n406), .B(n405), .Z(n407) );
  IVI U557 ( .A(n407), .Z(n408) );
  ND2I U558 ( .A(n409), .B(n408), .Z(n429) );
  IVI U559 ( .A(n1546), .Z(n1367) );
  IVI U560 ( .A(n1367), .Z(n1765) );
  NR2I U561 ( .A(n1765), .B(n4856), .Z(n412) );
  IVI U562 ( .A(n934), .Z(n2147) );
  ND2I U563 ( .A(n2147), .B(\gpr[16][12] ), .Z(n410) );
  ND2I U564 ( .A(n4709), .B(n410), .Z(n411) );
  NR2I U565 ( .A(n412), .B(n411), .Z(n427) );
  ND2I U566 ( .A(\gpr[23][12] ), .B(n2100), .Z(n415) );
  B5IP U567 ( .A(n413), .Z(n4694) );
  ND2I U568 ( .A(\gpr[20][12] ), .B(n4694), .Z(n414) );
  ND2I U569 ( .A(n415), .B(n414), .Z(n416) );
  IVI U570 ( .A(n416), .Z(n424) );
  ND2I U571 ( .A(\gpr[19][12] ), .B(n4703), .Z(n418) );
  ND2I U572 ( .A(n2292), .B(\gpr[21][12] ), .Z(n417) );
  ND2I U573 ( .A(n418), .B(n417), .Z(n422) );
  ND2I U574 ( .A(\gpr[17][12] ), .B(n206), .Z(n420) );
  ND2I U575 ( .A(\gpr[18][12] ), .B(n4726), .Z(n419) );
  ND2I U576 ( .A(n420), .B(n419), .Z(n421) );
  NR2I U577 ( .A(n422), .B(n421), .Z(n423) );
  ND2I U578 ( .A(n424), .B(n423), .Z(n425) );
  IVI U579 ( .A(n425), .Z(n426) );
  ND2I U580 ( .A(n427), .B(n426), .Z(n428) );
  ND2I U581 ( .A(n429), .B(n428), .Z(n430) );
  IVI U582 ( .A(n430), .Z(n461) );
  IVI U583 ( .A(n1083), .Z(n4718) );
  ND2I U584 ( .A(\gpr[13][12] ), .B(n4718), .Z(n434) );
  ND2I U585 ( .A(n2108), .B(\gpr[4][12] ), .Z(n433) );
  ND2I U586 ( .A(n2247), .B(\gpr[7][12] ), .Z(n431) );
  AN2I U587 ( .A(n431), .B(n2174), .Z(n432) );
  ND2I U588 ( .A(n434), .B(n229), .Z(n435) );
  IVI U589 ( .A(n1606), .Z(n2252) );
  NR2I U590 ( .A(n435), .B(n263), .Z(n445) );
  IVI U591 ( .A(n1915), .Z(n1797) );
  ND2I U592 ( .A(n101), .B(\gpr[10][12] ), .Z(n442) );
  IVI U593 ( .A(n672), .Z(n619) );
  IVI U594 ( .A(n619), .Z(n2197) );
  ND2I U595 ( .A(n2197), .B(\gpr[8][12] ), .Z(n439) );
  IVI U596 ( .A(n103), .Z(n1669) );
  ND2I U597 ( .A(n1669), .B(\gpr[11][12] ), .Z(n437) );
  IVI U598 ( .A(n1148), .Z(n1670) );
  ND2I U599 ( .A(n1670), .B(\gpr[2][12] ), .Z(n436) );
  AN2I U600 ( .A(n437), .B(n436), .Z(n438) );
  ND2I U601 ( .A(n439), .B(n438), .Z(n440) );
  IVI U602 ( .A(n440), .Z(n441) );
  ND2I U603 ( .A(n442), .B(n441), .Z(n443) );
  IVI U604 ( .A(n443), .Z(n444) );
  ND2I U605 ( .A(n445), .B(n444), .Z(n446) );
  IVI U606 ( .A(n446), .Z(n459) );
  ND2I U607 ( .A(\gpr[9][12] ), .B(n2125), .Z(n450) );
  IVI U608 ( .A(n556), .Z(n4740) );
  ND2I U609 ( .A(n2317), .B(\gpr[12][12] ), .Z(n448) );
  IVI U610 ( .A(n1432), .Z(n1846) );
  ND2I U611 ( .A(\gpr[15][12] ), .B(n1846), .Z(n447) );
  AN2I U612 ( .A(n448), .B(n447), .Z(n449) );
  ND2I U613 ( .A(n450), .B(n449), .Z(n457) );
  ND2I U614 ( .A(n4719), .B(\gpr[1][12] ), .Z(n455) );
  ND2I U615 ( .A(n105), .B(\gpr[6][12] ), .Z(n454) );
  IVI U616 ( .A(n1434), .Z(n909) );
  ND2I U617 ( .A(n2110), .B(\gpr[3][12] ), .Z(n452) );
  AN2I U618 ( .A(n1752), .B(n2037), .Z(n1520) );
  ND2I U619 ( .A(n1520), .B(\gpr[5][12] ), .Z(n451) );
  AN2I U620 ( .A(n452), .B(n451), .Z(n453) );
  ND2I U621 ( .A(n455), .B(n230), .Z(n456) );
  NR2I U622 ( .A(n457), .B(n456), .Z(n458) );
  ND2I U623 ( .A(n459), .B(n458), .Z(n460) );
  AN2I U624 ( .A(n461), .B(n460), .Z(rd_data1[12]) );
  IVI U625 ( .A(n492), .Z(n600) );
  IVI U626 ( .A(n600), .Z(n4707) );
  NR2I U627 ( .A(n4707), .B(n4872), .Z(n464) );
  IVI U628 ( .A(n1252), .Z(n1360) );
  ND2I U629 ( .A(n1360), .B(\gpr[17][23] ), .Z(n462) );
  ND2I U630 ( .A(n4709), .B(n462), .Z(n463) );
  NR2I U631 ( .A(n464), .B(n463), .Z(n478) );
  ND2I U632 ( .A(\gpr[20][23] ), .B(n2204), .Z(n466) );
  ND2I U633 ( .A(\gpr[21][23] ), .B(n2268), .Z(n465) );
  AN2I U634 ( .A(n466), .B(n465), .Z(n475) );
  B4I U635 ( .A(n467), .Z(n2216) );
  ND2I U636 ( .A(n2216), .B(\gpr[19][23] ), .Z(n469) );
  ND2I U637 ( .A(n4726), .B(\gpr[18][23] ), .Z(n468) );
  ND2I U638 ( .A(n469), .B(n468), .Z(n473) );
  ND2I U639 ( .A(\gpr[16][23] ), .B(n1762), .Z(n471) );
  ND2I U640 ( .A(n4704), .B(\gpr[23][23] ), .Z(n470) );
  ND2I U641 ( .A(n471), .B(n470), .Z(n472) );
  NR2I U642 ( .A(n473), .B(n472), .Z(n474) );
  ND2I U643 ( .A(n475), .B(n474), .Z(n476) );
  IVI U644 ( .A(n476), .Z(n477) );
  ND2I U645 ( .A(n478), .B(n477), .Z(n491) );
  IVI U646 ( .A(n601), .Z(n1275) );
  AO2 U647 ( .A(n2157), .B(\gpr[29][23] ), .C(n2276), .D(\gpr[25][23] ), .Z(
        n489) );
  ND2I U648 ( .A(n2147), .B(\gpr[24][23] ), .Z(n479) );
  ND2I U649 ( .A(n4690), .B(n479), .Z(n480) );
  IVI U650 ( .A(n480), .Z(n482) );
  ND2I U651 ( .A(n2216), .B(\gpr[27][23] ), .Z(n481) );
  ND2I U652 ( .A(n482), .B(n481), .Z(n483) );
  IVI U653 ( .A(n483), .Z(n488) );
  B4I U654 ( .A(n484), .Z(n2207) );
  ND2I U655 ( .A(\gpr[26][23] ), .B(n2207), .Z(n485) );
  IVI U656 ( .A(n600), .Z(n2092) );
  ND2I U657 ( .A(\gpr[28][23] ), .B(n2158), .Z(n487) );
  ND2I U658 ( .A(n2215), .B(\gpr[31][23] ), .Z(n486) );
  ND4P U659 ( .A(n489), .B(n488), .C(n209), .D(n221), .Z(n490) );
  AN2I U660 ( .A(n491), .B(n490), .Z(n523) );
  ND2I U661 ( .A(\gpr[15][23] ), .B(n1523), .Z(n497) );
  OR2P U662 ( .A(n2307), .B(n492), .Z(n493) );
  B4IP U663 ( .A(n493), .Z(n4746) );
  ND2I U664 ( .A(n4746), .B(\gpr[6][23] ), .Z(n496) );
  ND2I U665 ( .A(n1791), .B(\gpr[7][23] ), .Z(n495) );
  IVI U666 ( .A(n1606), .Z(n1990) );
  ND2I U667 ( .A(n1990), .B(\gpr[14][23] ), .Z(n494) );
  ND4 U668 ( .A(n497), .B(n496), .C(n495), .D(n494), .Z(n510) );
  ND2I U669 ( .A(n1307), .B(\gpr[8][23] ), .Z(n508) );
  IVI U670 ( .A(n1148), .Z(n1618) );
  ND2I U671 ( .A(n2189), .B(\gpr[2][23] ), .Z(n502) );
  IVI U672 ( .A(n1308), .Z(n2255) );
  ND2I U673 ( .A(n2255), .B(\gpr[11][23] ), .Z(n499) );
  IVI U674 ( .A(rd_addr1[4]), .Z(n498) );
  ND2I U675 ( .A(n499), .B(n498), .Z(n500) );
  IVI U676 ( .A(n500), .Z(n501) );
  AN2I U677 ( .A(n502), .B(n501), .Z(n507) );
  ND2I U678 ( .A(n4740), .B(\gpr[12][23] ), .Z(n505) );
  ND2I U679 ( .A(n503), .B(n685), .Z(n1499) );
  IVI U680 ( .A(n1499), .Z(n1346) );
  ND2I U681 ( .A(n1089), .B(\gpr[3][23] ), .Z(n504) );
  ND2I U682 ( .A(n2125), .B(\gpr[9][23] ), .Z(n506) );
  ND4P U683 ( .A(n508), .B(n507), .C(n222), .D(n506), .Z(n509) );
  NR2I U684 ( .A(n510), .B(n509), .Z(n521) );
  ND2I U685 ( .A(n4732), .B(\gpr[4][23] ), .Z(n515) );
  ND2I U686 ( .A(\gpr[13][23] ), .B(n4718), .Z(n512) );
  ND2I U687 ( .A(n4723), .B(\gpr[5][23] ), .Z(n511) );
  ND2I U688 ( .A(n512), .B(n511), .Z(n513) );
  IVI U689 ( .A(n513), .Z(n514) );
  ND2I U690 ( .A(n515), .B(n514), .Z(n519) );
  ND2I U691 ( .A(\gpr[1][23] ), .B(n4719), .Z(n517) );
  IVI U692 ( .A(n1915), .Z(n2328) );
  ND2I U693 ( .A(n2328), .B(\gpr[10][23] ), .Z(n516) );
  ND2I U694 ( .A(n517), .B(n516), .Z(n518) );
  NR2I U695 ( .A(n519), .B(n518), .Z(n520) );
  ND2I U696 ( .A(n521), .B(n520), .Z(n522) );
  ND2I U697 ( .A(n523), .B(n522), .Z(n524) );
  IVI U698 ( .A(n524), .Z(rd_data1[23]) );
  IVI U699 ( .A(n525), .Z(n2020) );
  ND2I U700 ( .A(n2020), .B(\gpr[30][18] ), .Z(n526) );
  AO3 U701 ( .A(n1633), .B(n4770), .C(n2079), .D(n526), .Z(n527) );
  IVI U702 ( .A(n527), .Z(n538) );
  ND2I U703 ( .A(\gpr[31][18] ), .B(n4704), .Z(n532) );
  ND2I U704 ( .A(\gpr[26][18] ), .B(n4702), .Z(n529) );
  ND2I U705 ( .A(\gpr[24][18] ), .B(n2233), .Z(n528) );
  ND2I U706 ( .A(n529), .B(n528), .Z(n530) );
  IVI U707 ( .A(n530), .Z(n531) );
  ND2I U708 ( .A(n532), .B(n531), .Z(n536) );
  ND2I U709 ( .A(\gpr[27][18] ), .B(n4703), .Z(n534) );
  IVI U710 ( .A(n1252), .Z(n2146) );
  ND2I U711 ( .A(\gpr[25][18] ), .B(n2146), .Z(n533) );
  NR2I U712 ( .A(n536), .B(n535), .Z(n537) );
  ND2I U713 ( .A(n538), .B(n537), .Z(n553) );
  NR2I U714 ( .A(n1810), .B(n4865), .Z(n541) );
  ND2I U715 ( .A(n1824), .B(\gpr[17][18] ), .Z(n539) );
  ND2I U716 ( .A(n4709), .B(n539), .Z(n540) );
  NR2I U717 ( .A(n541), .B(n540), .Z(n551) );
  ND2I U718 ( .A(\gpr[21][18] ), .B(n2157), .Z(n543) );
  ND2I U719 ( .A(\gpr[20][18] ), .B(n2204), .Z(n542) );
  ND2I U720 ( .A(n543), .B(n542), .Z(n549) );
  ND2I U721 ( .A(\gpr[16][18] ), .B(n2233), .Z(n547) );
  ND2I U722 ( .A(\gpr[23][18] ), .B(n2275), .Z(n546) );
  ND2I U723 ( .A(\gpr[19][18] ), .B(n4703), .Z(n545) );
  ND2I U724 ( .A(\gpr[18][18] ), .B(n4702), .Z(n544) );
  ND4P U725 ( .A(n547), .B(n546), .C(n545), .D(n544), .Z(n548) );
  NR2I U726 ( .A(n549), .B(n548), .Z(n550) );
  ND2I U727 ( .A(n551), .B(n550), .Z(n552) );
  AN2I U728 ( .A(n553), .B(n552), .Z(n586) );
  IVI U729 ( .A(n103), .Z(n4739) );
  ND2I U730 ( .A(n4739), .B(\gpr[11][18] ), .Z(n555) );
  ND2I U731 ( .A(n909), .B(\gpr[3][18] ), .Z(n554) );
  IVI U732 ( .A(n556), .Z(n2317) );
  ND2I U733 ( .A(n4740), .B(\gpr[12][18] ), .Z(n557) );
  ND2I U734 ( .A(n231), .B(n557), .Z(n558) );
  IVI U735 ( .A(n558), .Z(n560) );
  ND2I U736 ( .A(n102), .B(\gpr[10][18] ), .Z(n559) );
  ND2I U737 ( .A(n560), .B(n559), .Z(n561) );
  IVI U738 ( .A(n561), .Z(n572) );
  ND2I U739 ( .A(n2315), .B(\gpr[8][18] ), .Z(n564) );
  OR2I U740 ( .A(n562), .B(n4759), .Z(n563) );
  ND2I U741 ( .A(n564), .B(n563), .Z(n570) );
  AN2I U742 ( .A(n2307), .B(\gpr[13][18] ), .Z(n565) );
  ND2I U743 ( .A(n2268), .B(n565), .Z(n568) );
  ND2I U744 ( .A(\gpr[1][18] ), .B(n2320), .Z(n567) );
  IVI U745 ( .A(n1148), .Z(n1246) );
  ND2I U746 ( .A(n1246), .B(\gpr[2][18] ), .Z(n566) );
  NR2I U747 ( .A(n570), .B(n569), .Z(n571) );
  ND2I U748 ( .A(n572), .B(n571), .Z(n573) );
  IVI U749 ( .A(n573), .Z(n584) );
  ND2I U750 ( .A(n2125), .B(\gpr[9][18] ), .Z(n575) );
  ND2I U751 ( .A(\gpr[4][18] ), .B(n2303), .Z(n574) );
  ND2I U752 ( .A(n575), .B(n574), .Z(n582) );
  ND2I U753 ( .A(\gpr[6][18] ), .B(n4746), .Z(n580) );
  IVI U754 ( .A(n1432), .Z(n4745) );
  ND2I U755 ( .A(\gpr[15][18] ), .B(n4745), .Z(n579) );
  ND2I U756 ( .A(n576), .B(n685), .Z(n1446) );
  ND2I U757 ( .A(n2114), .B(\gpr[7][18] ), .Z(n578) );
  IVI U758 ( .A(n1606), .Z(n2311) );
  ND2I U759 ( .A(n2311), .B(\gpr[14][18] ), .Z(n577) );
  ND4P U760 ( .A(n580), .B(n579), .C(n578), .D(n577), .Z(n581) );
  NR2I U761 ( .A(n582), .B(n581), .Z(n583) );
  ND2I U762 ( .A(n584), .B(n583), .Z(n585) );
  ND2I U763 ( .A(n586), .B(n585), .Z(\rd_data1[18]_BAR ) );
  ND2I U764 ( .A(\gpr[19][4] ), .B(n2284), .Z(n589) );
  ND2I U765 ( .A(\gpr[21][4] ), .B(n2292), .Z(n588) );
  ND2I U766 ( .A(n589), .B(n588), .Z(n593) );
  ND2I U767 ( .A(\gpr[20][4] ), .B(n2158), .Z(n591) );
  ND2I U768 ( .A(\gpr[23][4] ), .B(n2100), .Z(n590) );
  ND2I U769 ( .A(n591), .B(n590), .Z(n592) );
  NR2I U770 ( .A(n593), .B(n592), .Z(n599) );
  ND2I U771 ( .A(n1938), .B(\gpr[17][4] ), .Z(n595) );
  ND2I U772 ( .A(n599), .B(n598), .Z(n618) );
  IVI U773 ( .A(n600), .Z(n4687) );
  NR2I U774 ( .A(n4687), .B(n4806), .Z(n604) );
  IVI U775 ( .A(n1275), .Z(n1952) );
  ND2I U776 ( .A(n1952), .B(\gpr[25][4] ), .Z(n602) );
  ND2I U777 ( .A(n4690), .B(n602), .Z(n603) );
  NR2I U778 ( .A(n604), .B(n603), .Z(n616) );
  ND2I U779 ( .A(\gpr[29][4] ), .B(n2268), .Z(n606) );
  ND2I U780 ( .A(\gpr[26][4] ), .B(n2077), .Z(n605) );
  AN2I U781 ( .A(n606), .B(n605), .Z(n608) );
  ND2I U782 ( .A(\gpr[28][4] ), .B(n2204), .Z(n607) );
  ND2I U783 ( .A(n608), .B(n607), .Z(n614) );
  ND2I U784 ( .A(n2100), .B(\gpr[31][4] ), .Z(n610) );
  ND2I U785 ( .A(n2284), .B(\gpr[27][4] ), .Z(n609) );
  AN2I U786 ( .A(n610), .B(n609), .Z(n612) );
  ND2I U787 ( .A(\gpr[24][4] ), .B(n1402), .Z(n611) );
  ND2I U788 ( .A(n612), .B(n611), .Z(n613) );
  NR2I U789 ( .A(n614), .B(n613), .Z(n615) );
  ND2I U790 ( .A(n616), .B(n615), .Z(n617) );
  AN2I U791 ( .A(n618), .B(n617), .Z(n645) );
  ND2I U792 ( .A(\gpr[1][4] ), .B(n4719), .Z(n621) );
  IVI U793 ( .A(n619), .Z(n1725) );
  ND2I U794 ( .A(\gpr[8][4] ), .B(n1725), .Z(n620) );
  ND2I U795 ( .A(n621), .B(n620), .Z(n626) );
  IVI U796 ( .A(n1446), .Z(n2061) );
  IVI U797 ( .A(n1148), .Z(n2189) );
  ND2I U798 ( .A(n1246), .B(\gpr[2][4] ), .Z(n622) );
  ND2I U799 ( .A(n2317), .B(\gpr[12][4] ), .Z(n623) );
  AN2I U800 ( .A(n265), .B(n623), .Z(n624) );
  ND2I U801 ( .A(n266), .B(n624), .Z(n625) );
  NR2I U802 ( .A(n626), .B(n625), .Z(n643) );
  ND2I U803 ( .A(\gpr[14][4] ), .B(n4748), .Z(n628) );
  ND2I U804 ( .A(n2125), .B(\gpr[9][4] ), .Z(n627) );
  ND2I U805 ( .A(n628), .B(n627), .Z(n641) );
  ND2I U806 ( .A(n1523), .B(\gpr[15][4] ), .Z(n630) );
  ND2I U807 ( .A(n101), .B(\gpr[10][4] ), .Z(n629) );
  AN2I U808 ( .A(n630), .B(n629), .Z(n639) );
  ND2I U809 ( .A(n1528), .B(\gpr[4][4] ), .Z(n632) );
  ND2I U810 ( .A(n1520), .B(\gpr[5][4] ), .Z(n631) );
  ND2I U811 ( .A(n632), .B(n631), .Z(n633) );
  IVI U812 ( .A(n633), .Z(n638) );
  IVI U813 ( .A(n1083), .Z(n2259) );
  ND2I U814 ( .A(n2259), .B(\gpr[13][4] ), .Z(n635) );
  ND2I U815 ( .A(n2110), .B(\gpr[3][4] ), .Z(n634) );
  ND2I U816 ( .A(n635), .B(n634), .Z(n636) );
  IVI U817 ( .A(n636), .Z(n637) );
  ND2I U818 ( .A(n639), .B(n232), .Z(n640) );
  NR2I U819 ( .A(n641), .B(n640), .Z(n642) );
  ND2I U820 ( .A(n643), .B(n642), .Z(n644) );
  ND2I U821 ( .A(n645), .B(n644), .Z(n646) );
  IVI U822 ( .A(n646), .Z(rd_data1[4]) );
  AO2 U823 ( .A(n2207), .B(\gpr[26][31] ), .C(n2268), .D(\gpr[29][31] ), .Z(
        n658) );
  NR2I U824 ( .A(n2092), .B(n4811), .Z(n649) );
  ND2I U825 ( .A(n1824), .B(\gpr[25][31] ), .Z(n647) );
  ND2I U826 ( .A(n2079), .B(n647), .Z(n648) );
  NR2I U827 ( .A(n649), .B(n648), .Z(n657) );
  ND2I U828 ( .A(\gpr[31][31] ), .B(n4704), .Z(n651) );
  ND2I U829 ( .A(\gpr[27][31] ), .B(n2216), .Z(n650) );
  ND2I U830 ( .A(n651), .B(n650), .Z(n655) );
  ND2I U831 ( .A(\gpr[28][31] ), .B(n2099), .Z(n653) );
  ND2I U832 ( .A(\gpr[24][31] ), .B(n878), .Z(n652) );
  ND2I U833 ( .A(n653), .B(n652), .Z(n654) );
  NR2I U834 ( .A(n655), .B(n654), .Z(n656) );
  IVI U835 ( .A(n659), .Z(n2047) );
  AO2 U836 ( .A(n1598), .B(\gpr[16][31] ), .C(n2047), .D(\gpr[17][31] ), .Z(
        n671) );
  NR2I U837 ( .A(n4687), .B(n4883), .Z(n662) );
  ND2I U838 ( .A(n2207), .B(\gpr[18][31] ), .Z(n660) );
  ND2I U839 ( .A(n2094), .B(n660), .Z(n661) );
  NR2I U840 ( .A(n662), .B(n661), .Z(n670) );
  ND2I U841 ( .A(n2216), .B(\gpr[19][31] ), .Z(n664) );
  ND2I U842 ( .A(\gpr[21][31] ), .B(n2292), .Z(n663) );
  ND2I U843 ( .A(n664), .B(n663), .Z(n668) );
  ND2I U844 ( .A(n2099), .B(\gpr[20][31] ), .Z(n666) );
  ND2I U845 ( .A(\gpr[23][31] ), .B(n2100), .Z(n665) );
  ND2I U846 ( .A(n666), .B(n665), .Z(n667) );
  NR2I U847 ( .A(n668), .B(n667), .Z(n669) );
  IVI U848 ( .A(n672), .Z(n1977) );
  IVI U849 ( .A(n1977), .Z(n1307) );
  ND2I U850 ( .A(n1307), .B(\gpr[8][31] ), .Z(n674) );
  ND2I U851 ( .A(\gpr[1][31] ), .B(n4719), .Z(n673) );
  ND2I U852 ( .A(n674), .B(n673), .Z(n684) );
  ND2I U853 ( .A(\gpr[13][31] ), .B(n2259), .Z(n679) );
  ND2I U854 ( .A(n104), .B(\gpr[6][31] ), .Z(n676) );
  ND2I U855 ( .A(\gpr[15][31] ), .B(n1523), .Z(n675) );
  ND2I U856 ( .A(n676), .B(n675), .Z(n677) );
  IVI U857 ( .A(n677), .Z(n678) );
  ND2I U858 ( .A(\gpr[5][31] ), .B(n4723), .Z(n681) );
  ND2I U859 ( .A(\gpr[10][31] ), .B(n102), .Z(n680) );
  ND2I U860 ( .A(n681), .B(n680), .Z(n682) );
  IVI U861 ( .A(n682), .Z(n683) );
  ND2I U862 ( .A(n1077), .B(n685), .Z(n1022) );
  IVI U863 ( .A(n1022), .Z(n1859) );
  ND2I U864 ( .A(n1859), .B(\gpr[3][31] ), .Z(n688) );
  ND2I U865 ( .A(n2306), .B(\gpr[7][31] ), .Z(n686) );
  AN2I U866 ( .A(n686), .B(n2174), .Z(n687) );
  ND2I U867 ( .A(n688), .B(n687), .Z(n694) );
  ND2I U868 ( .A(n106), .B(\gpr[12][31] ), .Z(n692) );
  ND2I U869 ( .A(n4739), .B(\gpr[11][31] ), .Z(n690) );
  ND2I U870 ( .A(n1246), .B(\gpr[2][31] ), .Z(n689) );
  AN2I U871 ( .A(n690), .B(n689), .Z(n691) );
  ND2I U872 ( .A(n692), .B(n691), .Z(n693) );
  NR2I U873 ( .A(n694), .B(n693), .Z(n696) );
  ND2I U874 ( .A(\gpr[4][31] ), .B(n4732), .Z(n695) );
  ND2I U875 ( .A(n2125), .B(\gpr[9][31] ), .Z(n698) );
  ND2I U876 ( .A(n1990), .B(\gpr[14][31] ), .Z(n697) );
  ND2I U877 ( .A(n698), .B(n697), .Z(n699) );
  ND2I U878 ( .A(rd_addr2[2]), .B(rd_addr2[1]), .Z(n734) );
  IVI U879 ( .A(n734), .Z(n701) );
  AN2I U880 ( .A(n725), .B(n701), .Z(n4500) );
  IVI U881 ( .A(n4500), .Z(n735) );
  B5IP U882 ( .A(n735), .Z(n4625) );
  ND2I U883 ( .A(n4625), .B(n4442), .Z(n3953) );
  IVI U884 ( .A(n3953), .Z(n3873) );
  IVI U885 ( .A(rd_addr2[4]), .Z(n702) );
  IVI U886 ( .A(n294), .Z(n4561) );
  IVI U887 ( .A(rd_addr2[1]), .Z(n707) );
  ND2I U888 ( .A(rd_addr2[2]), .B(n707), .Z(n711) );
  NR2I U889 ( .A(n725), .B(n711), .Z(n3365) );
  AN2I U890 ( .A(rd_addr2[2]), .B(rd_addr2[0]), .Z(n703) );
  ND2I U891 ( .A(n4442), .B(n703), .Z(n779) );
  IVI U892 ( .A(n707), .Z(n4223) );
  IVI U893 ( .A(n4223), .Z(n4184) );
  ND2I U894 ( .A(n4767), .B(n4184), .Z(n704) );
  AO3 U895 ( .A(\gpr[15][16] ), .B(n4090), .C(n4652), .D(n704), .Z(n705) );
  AO3 U896 ( .A(n4773), .B(n3953), .C(n4561), .D(n705), .Z(n721) );
  ND2I U897 ( .A(rd_addr2[0]), .B(n724), .Z(n706) );
  IVI U898 ( .A(n706), .Z(n708) );
  ND2I U899 ( .A(n708), .B(n4223), .Z(n4054) );
  IVI U900 ( .A(n4054), .Z(n709) );
  B2IP U901 ( .A(rd_addr2[3]), .Z1(n3428), .Z2(n4442) );
  AN2I U902 ( .A(n709), .B(n3428), .Z(n710) );
  B4IP U903 ( .A(n710), .Z(n767) );
  B4IP U904 ( .A(n767), .Z(n4557) );
  ND2I U905 ( .A(\gpr[3][16] ), .B(n4557), .Z(n719) );
  NR2I U906 ( .A(n725), .B(n711), .Z(n4104) );
  ND2I U907 ( .A(n4104), .B(n3428), .Z(n712) );
  B5IP U908 ( .A(n712), .Z(n4658) );
  ND2I U909 ( .A(\gpr[5][16] ), .B(n4658), .Z(n718) );
  NR2I U910 ( .A(rd_addr2[2]), .B(rd_addr2[1]), .Z(n723) );
  ND2I U911 ( .A(rd_addr2[0]), .B(n3428), .Z(n713) );
  IVI U912 ( .A(n713), .Z(n714) );
  ND2I U913 ( .A(n723), .B(n714), .Z(n766) );
  IVI U914 ( .A(n766), .Z(n4556) );
  ND2I U915 ( .A(\gpr[1][16] ), .B(n4556), .Z(n717) );
  AN2I U916 ( .A(rd_addr2[2]), .B(n725), .Z(n715) );
  IVI U917 ( .A(n4223), .Z(n726) );
  ND2I U918 ( .A(n715), .B(n726), .Z(n3401) );
  IVI U919 ( .A(n3401), .Z(n4138) );
  ND2I U920 ( .A(n4138), .B(n3428), .Z(n772) );
  IVI U921 ( .A(n772), .Z(n4153) );
  ND2I U922 ( .A(\gpr[4][16] ), .B(n4153), .Z(n716) );
  ND4 U923 ( .A(n719), .B(n718), .C(n717), .D(n716), .Z(n720) );
  NR2I U924 ( .A(n721), .B(n720), .Z(n743) );
  IVI U925 ( .A(rd_addr2[2]), .Z(n724) );
  B4IP U926 ( .A(n722), .Z(n4659) );
  ND2I U927 ( .A(\gpr[2][16] ), .B(n4659), .Z(n733) );
  ND2I U928 ( .A(n4442), .B(n3703), .Z(n771) );
  IVI U929 ( .A(n771), .Z(n4313) );
  ND2I U930 ( .A(\gpr[10][16] ), .B(n4313), .Z(n732) );
  ND2I U931 ( .A(n723), .B(rd_addr2[0]), .Z(n745) );
  IVI U932 ( .A(n745), .Z(n4490) );
  ND2I U933 ( .A(n4442), .B(n4490), .Z(n3598) );
  IVI U934 ( .A(n3598), .Z(n3558) );
  ND2I U935 ( .A(\gpr[9][16] ), .B(n3558), .Z(n731) );
  AN2I U936 ( .A(n725), .B(n724), .Z(n727) );
  ND2I U937 ( .A(n727), .B(n726), .Z(n3485) );
  IVI U938 ( .A(n3485), .Z(n728) );
  ND2I U939 ( .A(n728), .B(n4442), .Z(n729) );
  IVI U940 ( .A(n729), .Z(n3680) );
  IVI U941 ( .A(n3680), .Z(n3561) );
  IVI U942 ( .A(n3561), .Z(n3599) );
  ND2I U943 ( .A(\gpr[8][16] ), .B(n3599), .Z(n730) );
  ND2I U944 ( .A(n4442), .B(n709), .Z(n3513) );
  IVI U945 ( .A(n3513), .Z(n4320) );
  ND2I U946 ( .A(\gpr[11][16] ), .B(n4320), .Z(n739) );
  ND2I U947 ( .A(n4138), .B(n4442), .Z(n3514) );
  IVI U948 ( .A(n3514), .Z(n4321) );
  ND2I U949 ( .A(\gpr[12][16] ), .B(n4321), .Z(n738) );
  AN2I U950 ( .A(n701), .B(rd_addr2[0]), .Z(n3539) );
  ND2I U951 ( .A(n3539), .B(n3428), .Z(n3414) );
  ND2I U952 ( .A(\gpr[7][16] ), .B(n4675), .Z(n737) );
  IVI U953 ( .A(n735), .Z(n4489) );
  ND2I U954 ( .A(n4489), .B(n3428), .Z(n3562) );
  IVI U955 ( .A(n3562), .Z(n4524) );
  ND2I U956 ( .A(\gpr[6][16] ), .B(n4524), .Z(n736) );
  ND4 U957 ( .A(n739), .B(n738), .C(n737), .D(n736), .Z(n740) );
  NR2I U958 ( .A(n741), .B(n740), .Z(n742) );
  ND2I U959 ( .A(n743), .B(n742), .Z(n765) );
  IVI U960 ( .A(n4054), .Z(n744) );
  B2I U961 ( .A(n744), .Z2(n4009) );
  AO2 U962 ( .A(\gpr[18][16] ), .B(n3703), .C(\gpr[19][16] ), .D(n4009), .Z(
        n753) );
  IVI U963 ( .A(n745), .Z(n4286) );
  IVI U964 ( .A(n4286), .Z(n3400) );
  IVI U965 ( .A(n3400), .Z(n4296) );
  IVDAP U966 ( .A(n3401), .Y(n219), .Z(n796) );
  AO2 U967 ( .A(\gpr[17][16] ), .B(n4296), .C(\gpr[20][16] ), .D(n220), .Z(
        n752) );
  IVI U968 ( .A(n3539), .Z(n4130) );
  AO2 U969 ( .A(\gpr[23][16] ), .B(n4342), .C(\gpr[21][16] ), .D(n4090), .Z(
        n751) );
  AN2I U970 ( .A(\gpr[22][16] ), .B(n4625), .Z(n749) );
  ND2I U971 ( .A(rd_addr2[4]), .B(n3428), .Z(n746) );
  B5IP U972 ( .A(n746), .Z(n4628) );
  IVI U973 ( .A(n3485), .Z(n4637) );
  ND2I U974 ( .A(\gpr[16][16] ), .B(n4637), .Z(n747) );
  ND2I U975 ( .A(n4628), .B(n747), .Z(n748) );
  NR2I U976 ( .A(n749), .B(n748), .Z(n750) );
  ND4 U977 ( .A(n753), .B(n752), .C(n751), .D(n750), .Z(n762) );
  IVI U978 ( .A(n3538), .Z(n4214) );
  AO2 U979 ( .A(\gpr[26][16] ), .B(n4214), .C(\gpr[28][16] ), .D(n219), .Z(
        n760) );
  IVI U980 ( .A(n3485), .Z(n4450) );
  AO2 U981 ( .A(\gpr[24][16] ), .B(n4450), .C(\gpr[27][16] ), .D(n4009), .Z(
        n759) );
  IVI U982 ( .A(n4500), .Z(n3367) );
  B4IP U983 ( .A(n3367), .Z(n4431) );
  AO2 U984 ( .A(\gpr[30][16] ), .B(n4431), .C(\gpr[29][16] ), .D(n4090), .Z(
        n758) );
  AN2I U985 ( .A(n4442), .B(rd_addr2[4]), .Z(n792) );
  IVI U986 ( .A(n754), .Z(n4453) );
  IVI U987 ( .A(n4130), .Z(n4499) );
  ND2I U988 ( .A(\gpr[31][16] ), .B(n4499), .Z(n756) );
  ND2I U989 ( .A(\gpr[25][16] ), .B(n4490), .Z(n755) );
  AN3 U990 ( .A(n4453), .B(n756), .C(n755), .Z(n757) );
  ND4 U991 ( .A(n760), .B(n759), .C(n758), .D(n757), .Z(n761) );
  ND2I U992 ( .A(n762), .B(n761), .Z(n763) );
  IVI U993 ( .A(n763), .Z(n764) );
  AN2I U994 ( .A(n765), .B(n764), .Z(rd_data2[16]) );
  B5IP U995 ( .A(n766), .Z(n4656) );
  ND2I U996 ( .A(\gpr[1][10] ), .B(n4656), .Z(n770) );
  B4IP U997 ( .A(n767), .Z(n4657) );
  ND2I U998 ( .A(\gpr[3][10] ), .B(n4657), .Z(n769) );
  ND2I U999 ( .A(\gpr[5][10] ), .B(n4658), .Z(n768) );
  ND4 U1000 ( .A(n295), .B(n770), .C(n769), .D(n768), .Z(n778) );
  ND2I U1001 ( .A(\gpr[2][10] ), .B(n4659), .Z(n776) );
  IVI U1002 ( .A(n771), .Z(n4268) );
  ND2I U1003 ( .A(\gpr[10][10] ), .B(n4268), .Z(n775) );
  IVI U1004 ( .A(n772), .Z(n4308) );
  ND2I U1005 ( .A(\gpr[4][10] ), .B(n4153), .Z(n774) );
  ND2I U1006 ( .A(\gpr[9][10] ), .B(n3558), .Z(n773) );
  ND4 U1007 ( .A(n776), .B(n775), .C(n774), .D(n773), .Z(n777) );
  NR2I U1008 ( .A(n778), .B(n777), .Z(n791) );
  IVI U1009 ( .A(n3680), .Z(n3508) );
  ND2I U1010 ( .A(\gpr[8][10] ), .B(n3720), .Z(n783) );
  IVI U1011 ( .A(n3513), .Z(n4667) );
  ND2I U1012 ( .A(\gpr[11][10] ), .B(n4667), .Z(n782) );
  AN2I U1013 ( .A(rd_addr2[1]), .B(n4652), .Z(n4572) );
  ND2I U1014 ( .A(\gpr[15][10] ), .B(n4572), .Z(n781) );
  IVI U1015 ( .A(n3514), .Z(n4673) );
  ND2I U1016 ( .A(\gpr[12][10] ), .B(n4673), .Z(n780) );
  ND4 U1017 ( .A(n783), .B(n782), .C(n781), .D(n780), .Z(n789) );
  IVI U1018 ( .A(n3562), .Z(n4674) );
  ND2I U1019 ( .A(\gpr[6][10] ), .B(n4674), .Z(n787) );
  IVI U1020 ( .A(n4223), .Z(n3833) );
  AN2I U1021 ( .A(n4652), .B(n3833), .Z(n4578) );
  ND2I U1022 ( .A(\gpr[13][10] ), .B(n4578), .Z(n786) );
  ND2I U1023 ( .A(\gpr[7][10] ), .B(n4675), .Z(n785) );
  ND2I U1024 ( .A(n4625), .B(n4442), .Z(n4150) );
  IVI U1025 ( .A(n4150), .Z(n4579) );
  ND2I U1026 ( .A(\gpr[14][10] ), .B(n4579), .Z(n784) );
  ND4 U1027 ( .A(n787), .B(n786), .C(n785), .D(n784), .Z(n788) );
  NR2I U1028 ( .A(n789), .B(n788), .Z(n790) );
  ND2I U1029 ( .A(n791), .B(n790), .Z(n818) );
  IVI U1030 ( .A(n3539), .Z(n3778) );
  IVI U1031 ( .A(n3778), .Z(n4251) );
  B2I U1032 ( .A(n792), .Z1(n754), .Z2(n4641) );
  B2I U1033 ( .A(n709), .Z2(n4501) );
  IVI U1034 ( .A(n3400), .Z(n4001) );
  ND2I U1035 ( .A(n4214), .B(\gpr[26][10] ), .Z(n794) );
  B2IP U1036 ( .A(n3365), .Z2(n4090) );
  IVI U1037 ( .A(n3366), .Z(n4097) );
  ND2I U1038 ( .A(\gpr[29][10] ), .B(n4097), .Z(n793) );
  ND2I U1039 ( .A(n794), .B(n793), .Z(n795) );
  IVI U1040 ( .A(n795), .Z(n801) );
  ND2I U1041 ( .A(n4431), .B(\gpr[30][10] ), .Z(n798) );
  B5IP U1042 ( .A(n796), .Z(n4498) );
  ND2I U1043 ( .A(n4498), .B(\gpr[28][10] ), .Z(n797) );
  ND2I U1044 ( .A(n798), .B(n797), .Z(n799) );
  IVI U1045 ( .A(n799), .Z(n800) );
  ND2I U1046 ( .A(n801), .B(n800), .Z(n802) );
  ND2I U1047 ( .A(n804), .B(n803), .Z(n815) );
  IVI U1048 ( .A(n3538), .Z(n4293) );
  AO2 U1049 ( .A(\gpr[19][10] ), .B(n4009), .C(\gpr[18][10] ), .D(n4293), .Z(
        n813) );
  AO2 U1050 ( .A(\gpr[21][10] ), .B(n4090), .C(\gpr[22][10] ), .D(n4431), .Z(
        n811) );
  IVI U1051 ( .A(n3778), .Z(n3864) );
  ND2I U1052 ( .A(\gpr[16][10] ), .B(n4450), .Z(n805) );
  ND2I U1053 ( .A(n4001), .B(\gpr[17][10] ), .Z(n808) );
  B2I U1054 ( .A(n3401), .Z1(n220), .Z2(n806) );
  B5IP U1055 ( .A(n806), .Z(n4624) );
  ND2I U1056 ( .A(\gpr[20][10] ), .B(n4624), .Z(n807) );
  ND2I U1057 ( .A(n808), .B(n807), .Z(n809) );
  NR2I U1058 ( .A(n234), .B(n809), .Z(n810) );
  AN2I U1059 ( .A(n811), .B(n810), .Z(n812) );
  ND2I U1060 ( .A(n813), .B(n812), .Z(n814) );
  ND2I U1061 ( .A(n815), .B(n814), .Z(n816) );
  IVI U1062 ( .A(n816), .Z(n817) );
  AN2I U1063 ( .A(n818), .B(n817), .Z(rd_data2[10]) );
  ND2I U1064 ( .A(n2020), .B(\gpr[22][16] ), .Z(n819) );
  IVI U1065 ( .A(n820), .Z(n831) );
  ND2I U1066 ( .A(\gpr[18][16] ), .B(n2207), .Z(n822) );
  IVI U1067 ( .A(n1275), .Z(n1938) );
  ND2I U1068 ( .A(\gpr[17][16] ), .B(n1938), .Z(n821) );
  AN2I U1069 ( .A(n822), .B(n821), .Z(n830) );
  ND2I U1070 ( .A(\gpr[23][16] ), .B(n2215), .Z(n824) );
  ND2I U1071 ( .A(\gpr[19][16] ), .B(n4703), .Z(n823) );
  AN2I U1072 ( .A(n824), .B(n823), .Z(n829) );
  ND2I U1073 ( .A(\gpr[20][16] ), .B(n4694), .Z(n826) );
  IVI U1074 ( .A(n1268), .Z(n1553) );
  ND2I U1075 ( .A(\gpr[16][16] ), .B(n4686), .Z(n825) );
  ND2I U1076 ( .A(n826), .B(n825), .Z(n827) );
  IVI U1077 ( .A(n827), .Z(n828) );
  ND4P U1078 ( .A(n831), .B(n830), .C(n829), .D(n828), .Z(n848) );
  B3IP U1079 ( .A(n1545), .Z1(n2292), .Z2(n1007) );
  ND2I U1080 ( .A(n2020), .B(\gpr[30][16] ), .Z(n832) );
  AO3 U1081 ( .A(n1007), .B(n4831), .C(n4690), .D(n832), .Z(n833) );
  IVI U1082 ( .A(n833), .Z(n846) );
  ND2I U1083 ( .A(n2215), .B(\gpr[31][16] ), .Z(n835) );
  ND2I U1084 ( .A(\gpr[27][16] ), .B(n4703), .Z(n834) );
  ND2I U1085 ( .A(n835), .B(n834), .Z(n844) );
  IVI U1086 ( .A(n1275), .Z(n1383) );
  ND2I U1087 ( .A(\gpr[25][16] ), .B(n1383), .Z(n837) );
  ND2I U1088 ( .A(\gpr[24][16] ), .B(n1762), .Z(n836) );
  AN2I U1089 ( .A(n837), .B(n836), .Z(n842) );
  B2IP U1090 ( .A(n1631), .Z1(n838), .Z2(n2204) );
  IVI U1091 ( .A(n838), .Z(n1424) );
  ND2I U1092 ( .A(n1424), .B(\gpr[28][16] ), .Z(n840) );
  ND2I U1093 ( .A(\gpr[26][16] ), .B(n2207), .Z(n839) );
  AN2I U1094 ( .A(n840), .B(n839), .Z(n841) );
  ND2I U1095 ( .A(n842), .B(n841), .Z(n843) );
  NR2I U1096 ( .A(n844), .B(n843), .Z(n845) );
  ND2I U1097 ( .A(n846), .B(n845), .Z(n847) );
  ND2I U1098 ( .A(n848), .B(n847), .Z(n849) );
  IVI U1099 ( .A(n849), .Z(n876) );
  AO2 U1100 ( .A(\gpr[15][16] ), .B(n1846), .C(n105), .D(\gpr[6][16] ), .Z(
        n874) );
  IVI U1101 ( .A(n850), .Z(n1528) );
  ND2I U1102 ( .A(n1528), .B(\gpr[4][16] ), .Z(n851) );
  ND2I U1103 ( .A(n498), .B(n851), .Z(n855) );
  ND2I U1104 ( .A(\gpr[13][16] ), .B(n2188), .Z(n853) );
  IVI U1105 ( .A(n1499), .Z(n4724) );
  ND2I U1106 ( .A(n4724), .B(\gpr[3][16] ), .Z(n852) );
  ND2I U1107 ( .A(n853), .B(n852), .Z(n854) );
  NR2I U1108 ( .A(n855), .B(n854), .Z(n873) );
  B2I U1109 ( .A(n2320), .Z2(n1240) );
  ND2I U1110 ( .A(\gpr[1][16] ), .B(n1240), .Z(n857) );
  IVI U1111 ( .A(n1148), .Z(n2256) );
  ND2I U1112 ( .A(\gpr[2][16] ), .B(n2256), .Z(n856) );
  AN2I U1113 ( .A(n857), .B(n856), .Z(n860) );
  IVI U1114 ( .A(n2173), .Z(n2306) );
  ND2I U1115 ( .A(\gpr[7][16] ), .B(n2306), .Z(n859) );
  ND2I U1116 ( .A(\gpr[5][16] ), .B(n1520), .Z(n858) );
  ND2I U1117 ( .A(n860), .B(n267), .Z(n861) );
  IVI U1118 ( .A(n861), .Z(n872) );
  AO2 U1119 ( .A(n4702), .B(\gpr[10][16] ), .C(n1360), .D(\gpr[9][16] ), .Z(
        n869) );
  ND2I U1120 ( .A(n2204), .B(\gpr[12][16] ), .Z(n866) );
  ND2I U1121 ( .A(n4688), .B(\gpr[11][16] ), .Z(n864) );
  AO2 U1122 ( .A(n862), .B(\gpr[14][16] ), .C(n2048), .D(\gpr[8][16] ), .Z(
        n863) );
  AN2I U1123 ( .A(n864), .B(n863), .Z(n865) );
  ND2I U1124 ( .A(n866), .B(n865), .Z(n867) );
  IVI U1125 ( .A(n867), .Z(n868) );
  ND2I U1126 ( .A(n869), .B(n868), .Z(n870) );
  ND2I U1127 ( .A(n2307), .B(n870), .Z(n871) );
  ND4P U1128 ( .A(n874), .B(n873), .C(n872), .D(n871), .Z(n875) );
  ND2I U1129 ( .A(n876), .B(n875), .Z(n877) );
  IVI U1130 ( .A(n877), .Z(rd_data1[16]) );
  NR2I U1131 ( .A(n1765), .B(n4870), .Z(n881) );
  ND2I U1132 ( .A(n878), .B(\gpr[16][22] ), .Z(n879) );
  ND2I U1133 ( .A(n4709), .B(n879), .Z(n880) );
  NR2I U1134 ( .A(n881), .B(n880), .Z(n891) );
  ND2I U1135 ( .A(\gpr[17][22] ), .B(n2146), .Z(n883) );
  ND2I U1136 ( .A(\gpr[21][22] ), .B(n4701), .Z(n882) );
  ND2I U1137 ( .A(n883), .B(n882), .Z(n889) );
  ND2I U1138 ( .A(\gpr[19][22] ), .B(n2284), .Z(n887) );
  ND2I U1139 ( .A(\gpr[18][22] ), .B(n2207), .Z(n886) );
  ND2I U1140 ( .A(\gpr[20][22] ), .B(n4694), .Z(n885) );
  ND2I U1141 ( .A(\gpr[23][22] ), .B(n4704), .Z(n884) );
  ND4P U1142 ( .A(n887), .B(n886), .C(n885), .D(n884), .Z(n888) );
  NR2I U1143 ( .A(n889), .B(n888), .Z(n890) );
  ND2I U1144 ( .A(n891), .B(n890), .Z(n906) );
  AO2 U1145 ( .A(n2207), .B(\gpr[26][22] ), .C(n2157), .D(\gpr[29][22] ), .Z(
        n904) );
  NR2I U1146 ( .A(n1889), .B(n4871), .Z(n894) );
  ND2I U1147 ( .A(n1205), .B(\gpr[24][22] ), .Z(n892) );
  ND2I U1148 ( .A(n4690), .B(n892), .Z(n893) );
  NR2I U1149 ( .A(n894), .B(n893), .Z(n902) );
  ND2I U1150 ( .A(n4704), .B(\gpr[31][22] ), .Z(n896) );
  ND2I U1151 ( .A(n2284), .B(\gpr[27][22] ), .Z(n895) );
  ND2I U1152 ( .A(n896), .B(n895), .Z(n900) );
  ND2I U1153 ( .A(n2204), .B(\gpr[28][22] ), .Z(n898) );
  ND2I U1154 ( .A(\gpr[25][22] ), .B(n2146), .Z(n897) );
  ND2I U1155 ( .A(n898), .B(n897), .Z(n899) );
  NR2I U1156 ( .A(n900), .B(n899), .Z(n901) );
  AN2I U1157 ( .A(n902), .B(n901), .Z(n903) );
  ND2I U1158 ( .A(n904), .B(n903), .Z(n905) );
  AN2I U1159 ( .A(n906), .B(n905), .Z(n932) );
  ND2I U1160 ( .A(\gpr[13][22] ), .B(n2259), .Z(n908) );
  ND2I U1161 ( .A(n1670), .B(\gpr[2][22] ), .Z(n907) );
  ND2I U1162 ( .A(n4723), .B(\gpr[5][22] ), .Z(n913) );
  ND2I U1163 ( .A(n1528), .B(\gpr[4][22] ), .Z(n912) );
  ND2I U1164 ( .A(n909), .B(\gpr[3][22] ), .Z(n911) );
  ND2I U1165 ( .A(n1797), .B(\gpr[10][22] ), .Z(n910) );
  ND4 U1166 ( .A(n913), .B(n912), .C(n911), .D(n910), .Z(n914) );
  NR2I U1167 ( .A(n915), .B(n914), .Z(n930) );
  ND2I U1168 ( .A(\gpr[15][22] ), .B(n4745), .Z(n919) );
  ND2I U1169 ( .A(n4746), .B(\gpr[6][22] ), .Z(n918) );
  ND2I U1170 ( .A(n1791), .B(\gpr[7][22] ), .Z(n917) );
  ND2I U1171 ( .A(n2252), .B(\gpr[14][22] ), .Z(n916) );
  ND4 U1172 ( .A(n919), .B(n918), .C(n917), .D(n916), .Z(n928) );
  ND2I U1173 ( .A(n2125), .B(\gpr[9][22] ), .Z(n926) );
  ND2I U1174 ( .A(n2197), .B(\gpr[8][22] ), .Z(n924) );
  ND2I U1175 ( .A(n106), .B(\gpr[12][22] ), .Z(n921) );
  ND2I U1176 ( .A(n1970), .B(\gpr[11][22] ), .Z(n920) );
  ND2I U1177 ( .A(n921), .B(n920), .Z(n922) );
  IVI U1178 ( .A(n922), .Z(n923) );
  AN2I U1179 ( .A(n924), .B(n923), .Z(n925) );
  ND2I U1180 ( .A(n926), .B(n925), .Z(n927) );
  NR2I U1181 ( .A(n928), .B(n927), .Z(n929) );
  ND2I U1182 ( .A(n930), .B(n929), .Z(n931) );
  ND2I U1183 ( .A(n932), .B(n931), .Z(n933) );
  IVI U1184 ( .A(n933), .Z(rd_data1[22]) );
  IVI U1185 ( .A(n934), .Z(n2296) );
  AO2 U1186 ( .A(n2296), .B(\gpr[24][30] ), .C(n4688), .D(\gpr[27][30] ), .Z(
        n948) );
  NR2I U1187 ( .A(n1889), .B(n4881), .Z(n937) );
  ND2I U1188 ( .A(n206), .B(\gpr[25][30] ), .Z(n935) );
  ND2I U1189 ( .A(n4690), .B(n935), .Z(n936) );
  NR2I U1190 ( .A(n937), .B(n936), .Z(n946) );
  ND2I U1191 ( .A(\gpr[29][30] ), .B(n2292), .Z(n939) );
  ND2I U1192 ( .A(\gpr[26][30] ), .B(n2077), .Z(n938) );
  ND2I U1193 ( .A(n939), .B(n938), .Z(n944) );
  ND2I U1194 ( .A(\gpr[28][30] ), .B(n2099), .Z(n942) );
  ND2I U1195 ( .A(\gpr[31][30] ), .B(n4704), .Z(n941) );
  ND2I U1196 ( .A(n942), .B(n941), .Z(n943) );
  NR2I U1197 ( .A(n944), .B(n943), .Z(n945) );
  AN2I U1198 ( .A(n946), .B(n945), .Z(n947) );
  ND2I U1199 ( .A(n948), .B(n947), .Z(n964) );
  AO2 U1200 ( .A(n4702), .B(\gpr[18][30] ), .C(n1647), .D(\gpr[17][30] ), .Z(
        n952) );
  ND2I U1201 ( .A(\gpr[19][30] ), .B(n4688), .Z(n950) );
  ND2I U1202 ( .A(\gpr[23][30] ), .B(n4704), .Z(n949) );
  AN2I U1203 ( .A(n950), .B(n949), .Z(n951) );
  AN2I U1204 ( .A(n952), .B(n951), .Z(n962) );
  NR2I U1205 ( .A(n4707), .B(n4882), .Z(n955) );
  IVI U1206 ( .A(n1268), .Z(n1063) );
  IVI U1207 ( .A(n1063), .Z(n2017) );
  ND2I U1208 ( .A(\gpr[16][30] ), .B(n2017), .Z(n953) );
  ND2I U1209 ( .A(n4709), .B(n953), .Z(n954) );
  NR2I U1210 ( .A(n955), .B(n954), .Z(n959) );
  ND2I U1211 ( .A(n2158), .B(\gpr[20][30] ), .Z(n957) );
  ND2I U1212 ( .A(\gpr[21][30] ), .B(n2292), .Z(n956) );
  AN2I U1213 ( .A(n957), .B(n956), .Z(n958) );
  ND2I U1214 ( .A(n959), .B(n958), .Z(n960) );
  IVI U1215 ( .A(n960), .Z(n961) );
  ND2I U1216 ( .A(n962), .B(n961), .Z(n963) );
  AN2I U1217 ( .A(n964), .B(n963), .Z(n994) );
  ND2I U1218 ( .A(n4719), .B(\gpr[1][30] ), .Z(n965) );
  IVI U1219 ( .A(n965), .Z(n969) );
  ND2I U1220 ( .A(n2259), .B(\gpr[13][30] ), .Z(n967) );
  ND2I U1221 ( .A(n1669), .B(\gpr[11][30] ), .Z(n966) );
  ND2I U1222 ( .A(n967), .B(n268), .Z(n968) );
  NR2I U1223 ( .A(n969), .B(n968), .Z(n979) );
  ND2I U1224 ( .A(\gpr[10][30] ), .B(n101), .Z(n976) );
  ND2I U1225 ( .A(n106), .B(\gpr[12][30] ), .Z(n973) );
  ND2I U1226 ( .A(n1618), .B(\gpr[2][30] ), .Z(n971) );
  IVI U1227 ( .A(n1022), .Z(n2040) );
  ND2I U1228 ( .A(n2040), .B(\gpr[3][30] ), .Z(n970) );
  AN2I U1229 ( .A(n971), .B(n970), .Z(n972) );
  ND2I U1230 ( .A(n973), .B(n972), .Z(n974) );
  IVI U1231 ( .A(n974), .Z(n975) );
  ND2I U1232 ( .A(n976), .B(n975), .Z(n977) );
  NR2I U1233 ( .A(n235), .B(n977), .Z(n978) );
  AN2I U1234 ( .A(n979), .B(n978), .Z(n992) );
  ND2I U1235 ( .A(n1846), .B(\gpr[15][30] ), .Z(n983) );
  ND2I U1236 ( .A(n4746), .B(\gpr[6][30] ), .Z(n982) );
  ND2I U1237 ( .A(n1791), .B(\gpr[7][30] ), .Z(n981) );
  ND2I U1238 ( .A(n2252), .B(\gpr[14][30] ), .Z(n980) );
  ND4 U1239 ( .A(n983), .B(n982), .C(n981), .D(n980), .Z(n990) );
  ND2I U1240 ( .A(\gpr[4][30] ), .B(n2303), .Z(n988) );
  ND2I U1241 ( .A(n2129), .B(\gpr[8][30] ), .Z(n985) );
  IVI U1242 ( .A(n1320), .Z(n4737) );
  ND2I U1243 ( .A(\gpr[9][30] ), .B(n4737), .Z(n984) );
  ND2I U1244 ( .A(n985), .B(n984), .Z(n986) );
  IVI U1245 ( .A(n986), .Z(n987) );
  ND2I U1246 ( .A(n988), .B(n987), .Z(n989) );
  NR2I U1247 ( .A(n990), .B(n989), .Z(n991) );
  ND2I U1248 ( .A(n992), .B(n991), .Z(n993) );
  AN2I U1249 ( .A(n994), .B(n993), .Z(rd_data1[30]) );
  NR2I U1250 ( .A(n4707), .B(n4809), .Z(n997) );
  IVI U1251 ( .A(n1363), .Z(n1583) );
  ND2I U1252 ( .A(n1583), .B(\gpr[24][26] ), .Z(n995) );
  ND2I U1253 ( .A(n2079), .B(n995), .Z(n996) );
  ND2I U1254 ( .A(\gpr[25][26] ), .B(n206), .Z(n999) );
  ND2I U1255 ( .A(\gpr[29][26] ), .B(n2157), .Z(n998) );
  AN2I U1256 ( .A(n999), .B(n998), .Z(n1005) );
  ND2I U1257 ( .A(\gpr[31][26] ), .B(n2275), .Z(n1001) );
  ND2I U1258 ( .A(\gpr[26][26] ), .B(n4702), .Z(n1000) );
  AN2I U1259 ( .A(n1001), .B(n1000), .Z(n1003) );
  ND2I U1260 ( .A(\gpr[27][26] ), .B(n2284), .Z(n1002) );
  ND2I U1261 ( .A(\gpr[28][26] ), .B(n1424), .Z(n1004) );
  IVI U1262 ( .A(n1275), .Z(n1824) );
  AO2 U1263 ( .A(n1402), .B(\gpr[16][26] ), .C(n1824), .D(\gpr[17][26] ), .Z(
        n1017) );
  ND2I U1264 ( .A(n2020), .B(\gpr[22][26] ), .Z(n1006) );
  IVI U1265 ( .A(n1008), .Z(n1016) );
  ND2I U1266 ( .A(n4704), .B(\gpr[23][26] ), .Z(n1010) );
  ND2I U1267 ( .A(n2207), .B(\gpr[18][26] ), .Z(n1009) );
  ND2I U1268 ( .A(n1010), .B(n1009), .Z(n1014) );
  ND2I U1269 ( .A(\gpr[20][26] ), .B(n2099), .Z(n1012) );
  ND2I U1270 ( .A(n2284), .B(\gpr[19][26] ), .Z(n1011) );
  ND2I U1271 ( .A(n1012), .B(n1011), .Z(n1013) );
  NR2I U1272 ( .A(n1014), .B(n1013), .Z(n1015) );
  ND2I U1273 ( .A(\gpr[1][26] ), .B(n4719), .Z(n1019) );
  ND2I U1274 ( .A(n2115), .B(\gpr[2][26] ), .Z(n1018) );
  ND2I U1275 ( .A(n102), .B(\gpr[10][26] ), .Z(n1027) );
  AN2I U1276 ( .A(n2037), .B(\gpr[5][26] ), .Z(n1021) );
  IVI U1277 ( .A(n1022), .Z(n1089) );
  ND2I U1278 ( .A(n1089), .B(\gpr[3][26] ), .Z(n1024) );
  ND2I U1279 ( .A(n1528), .B(\gpr[4][26] ), .Z(n1023) );
  ND2I U1280 ( .A(n1024), .B(n1023), .Z(n1025) );
  NR2I U1281 ( .A(n269), .B(n1025), .Z(n1026) );
  ND2I U1282 ( .A(\gpr[15][26] ), .B(n1846), .Z(n1031) );
  ND2I U1283 ( .A(n4746), .B(\gpr[6][26] ), .Z(n1030) );
  ND2I U1284 ( .A(n4747), .B(\gpr[7][26] ), .Z(n1029) );
  ND2I U1285 ( .A(n2252), .B(\gpr[14][26] ), .Z(n1028) );
  ND4 U1286 ( .A(n1031), .B(n1030), .C(n1029), .D(n1028), .Z(n1039) );
  ND2I U1287 ( .A(n2125), .B(\gpr[9][26] ), .Z(n1038) );
  ND2I U1288 ( .A(n2129), .B(\gpr[8][26] ), .Z(n1036) );
  ND2I U1289 ( .A(n2317), .B(\gpr[12][26] ), .Z(n1033) );
  ND2I U1290 ( .A(n2255), .B(\gpr[11][26] ), .Z(n1032) );
  ND2I U1291 ( .A(n1033), .B(n1032), .Z(n1034) );
  IVI U1292 ( .A(n1034), .Z(n1035) );
  AN2I U1293 ( .A(n1036), .B(n1035), .Z(n1037) );
  AO2 U1294 ( .A(n4726), .B(\gpr[26][7] ), .C(n2268), .D(\gpr[29][7] ), .Z(
        n1053) );
  ND2I U1295 ( .A(n4703), .B(\gpr[27][7] ), .Z(n1041) );
  ND2I U1296 ( .A(\gpr[24][7] ), .B(n2017), .Z(n1040) );
  ND2I U1297 ( .A(n1041), .B(n1040), .Z(n1045) );
  ND2I U1298 ( .A(n2100), .B(\gpr[31][7] ), .Z(n1043) );
  ND2I U1299 ( .A(\gpr[28][7] ), .B(n4694), .Z(n1042) );
  ND2I U1300 ( .A(n1043), .B(n1042), .Z(n1044) );
  NR2I U1301 ( .A(n1045), .B(n1044), .Z(n1050) );
  NR2I U1302 ( .A(n1810), .B(n4849), .Z(n1048) );
  ND2I U1303 ( .A(n1466), .B(\gpr[25][7] ), .Z(n1046) );
  ND2I U1304 ( .A(n4690), .B(n1046), .Z(n1047) );
  NR2I U1305 ( .A(n1048), .B(n1047), .Z(n1049) );
  ND2I U1306 ( .A(n1050), .B(n1049), .Z(n1051) );
  IVI U1307 ( .A(n1051), .Z(n1052) );
  ND2I U1308 ( .A(n1053), .B(n1052), .Z(n1067) );
  ND2I U1309 ( .A(\gpr[21][7] ), .B(n4701), .Z(n1055) );
  ND2I U1310 ( .A(\gpr[19][7] ), .B(n4703), .Z(n1054) );
  ND2I U1311 ( .A(n1055), .B(n1054), .Z(n1059) );
  ND2I U1312 ( .A(\gpr[23][7] ), .B(n2100), .Z(n1057) );
  ND2I U1313 ( .A(\gpr[20][7] ), .B(n2158), .Z(n1056) );
  ND2I U1314 ( .A(n1057), .B(n1056), .Z(n1058) );
  NR2I U1315 ( .A(n1059), .B(n1058), .Z(n1065) );
  NR2I U1316 ( .A(n1810), .B(n4848), .Z(n1062) );
  ND2I U1317 ( .A(n1938), .B(\gpr[17][7] ), .Z(n1060) );
  ND2I U1318 ( .A(n2094), .B(n1060), .Z(n1061) );
  ND2I U1319 ( .A(n1065), .B(n1064), .Z(n1066) );
  ND2I U1320 ( .A(n1067), .B(n1066), .Z(n1068) );
  IVI U1321 ( .A(n1068), .Z(n1104) );
  ND2I U1322 ( .A(\gpr[1][7] ), .B(n4719), .Z(n1071) );
  ND2I U1323 ( .A(n1307), .B(\gpr[8][7] ), .Z(n1070) );
  ND2I U1324 ( .A(n2328), .B(\gpr[10][7] ), .Z(n1069) );
  ND2I U1325 ( .A(n1071), .B(n236), .Z(n1074) );
  ND2I U1326 ( .A(n2303), .B(\gpr[4][7] ), .Z(n1072) );
  IVI U1327 ( .A(n1072), .Z(n1073) );
  NR2I U1328 ( .A(n1074), .B(n1073), .Z(n1102) );
  ND2I U1329 ( .A(\gpr[9][7] ), .B(n2125), .Z(n1082) );
  ND2I U1330 ( .A(n2317), .B(\gpr[12][7] ), .Z(n1079) );
  NR2I U1331 ( .A(n1075), .B(n5061), .Z(n1076) );
  ND2I U1332 ( .A(n1077), .B(n1076), .Z(n1078) );
  ND2I U1333 ( .A(n1079), .B(n270), .Z(n1080) );
  NR2I U1334 ( .A(n1080), .B(n271), .Z(n1081) );
  ND2I U1335 ( .A(n1082), .B(n1081), .Z(n1100) );
  ND2I U1336 ( .A(n104), .B(\gpr[6][7] ), .Z(n1085) );
  IVI U1337 ( .A(n1083), .Z(n2058) );
  ND2I U1338 ( .A(\gpr[13][7] ), .B(n2058), .Z(n1084) );
  ND2I U1339 ( .A(n1085), .B(n1084), .Z(n1088) );
  ND2I U1340 ( .A(\gpr[15][7] ), .B(n4745), .Z(n1086) );
  IVI U1341 ( .A(n1086), .Z(n1087) );
  NR2I U1342 ( .A(n1088), .B(n1087), .Z(n1098) );
  ND2I U1343 ( .A(n1089), .B(\gpr[3][7] ), .Z(n1093) );
  ND2I U1344 ( .A(n2061), .B(\gpr[7][7] ), .Z(n1091) );
  ND2I U1345 ( .A(n1727), .B(\gpr[2][7] ), .Z(n1090) );
  AN2I U1346 ( .A(n1091), .B(n1090), .Z(n1092) );
  ND2I U1347 ( .A(n1093), .B(n1092), .Z(n1096) );
  ND2I U1348 ( .A(\gpr[5][7] ), .B(n4723), .Z(n1094) );
  IVI U1349 ( .A(n1094), .Z(n1095) );
  NR2I U1350 ( .A(n1096), .B(n1095), .Z(n1097) );
  ND2I U1351 ( .A(n1098), .B(n1097), .Z(n1099) );
  NR2I U1352 ( .A(n1100), .B(n1099), .Z(n1101) );
  ND2I U1353 ( .A(n1102), .B(n1101), .Z(n1103) );
  AN2I U1354 ( .A(n1104), .B(n1103), .Z(rd_data1[7]) );
  IVI U1355 ( .A(n1553), .Z(n1762) );
  AO2 U1356 ( .A(n1762), .B(\gpr[16][20] ), .C(n1466), .D(\gpr[17][20] ), .Z(
        n1113) );
  B3IP U1357 ( .A(n1545), .Z1(n2157), .Z2(n4693) );
  ND2I U1358 ( .A(n2020), .B(\gpr[22][20] ), .Z(n1105) );
  AO3 U1359 ( .A(n4693), .B(n4832), .C(n2094), .D(n1105), .Z(n1111) );
  ND2I U1360 ( .A(\gpr[19][20] ), .B(n4703), .Z(n1109) );
  ND2I U1361 ( .A(\gpr[18][20] ), .B(n4702), .Z(n1108) );
  ND2I U1362 ( .A(\gpr[20][20] ), .B(n2099), .Z(n1107) );
  ND2I U1363 ( .A(\gpr[23][20] ), .B(n2275), .Z(n1106) );
  ND4P U1364 ( .A(n1109), .B(n1108), .C(n1107), .D(n1106), .Z(n1110) );
  NR2I U1365 ( .A(n1111), .B(n1110), .Z(n1112) );
  ND2I U1366 ( .A(n1113), .B(n1112), .Z(n1131) );
  ND2I U1367 ( .A(\gpr[26][20] ), .B(n2207), .Z(n1115) );
  ND2I U1368 ( .A(\gpr[27][20] ), .B(n2216), .Z(n1114) );
  ND2I U1369 ( .A(n1115), .B(n1114), .Z(n1125) );
  ND2I U1370 ( .A(\gpr[28][20] ), .B(n2158), .Z(n1123) );
  IVI U1371 ( .A(n1136), .Z(n2233) );
  ND2I U1372 ( .A(\gpr[24][20] ), .B(n2233), .Z(n1117) );
  ND2I U1373 ( .A(\gpr[25][20] ), .B(n2276), .Z(n1116) );
  ND2I U1374 ( .A(n1117), .B(n1116), .Z(n1118) );
  IVI U1375 ( .A(n1118), .Z(n1120) );
  ND2I U1376 ( .A(\gpr[30][20] ), .B(n207), .Z(n1119) );
  ND2I U1377 ( .A(n1120), .B(n1119), .Z(n1121) );
  IVI U1378 ( .A(n1121), .Z(n1122) );
  ND2I U1379 ( .A(n1123), .B(n1122), .Z(n1124) );
  NR2I U1380 ( .A(n1125), .B(n1124), .Z(n1129) );
  B3IP U1381 ( .A(n1469), .Z1(n2268), .Z2(n2022) );
  ND2I U1382 ( .A(n4704), .B(\gpr[31][20] ), .Z(n1126) );
  AO3 U1383 ( .A(n2022), .B(n4833), .C(n4690), .D(n1126), .Z(n1127) );
  IVI U1384 ( .A(n1127), .Z(n1128) );
  ND2I U1385 ( .A(n1129), .B(n1128), .Z(n1130) );
  AN2I U1386 ( .A(n1131), .B(n1130), .Z(n1159) );
  ND2I U1387 ( .A(\gpr[1][20] ), .B(n4719), .Z(n1133) );
  IVDAP U1388 ( .A(n1528), .Z(n1168) );
  ND2I U1389 ( .A(n1168), .B(\gpr[4][20] ), .Z(n1132) );
  ND2I U1390 ( .A(n1133), .B(n1132), .Z(n1147) );
  IVI U1391 ( .A(n1446), .Z(n2114) );
  AO2 U1392 ( .A(n104), .B(\gpr[6][20] ), .C(n2114), .D(\gpr[7][20] ), .Z(
        n1145) );
  IVI U1393 ( .A(n1252), .Z(n1647) );
  ND2I U1394 ( .A(\gpr[9][20] ), .B(n1647), .Z(n1135) );
  ND2I U1395 ( .A(\gpr[10][20] ), .B(n4702), .Z(n1134) );
  ND2I U1396 ( .A(n1135), .B(n1134), .Z(n1140) );
  ND2I U1397 ( .A(n4688), .B(\gpr[11][20] ), .Z(n1138) );
  ND2I U1398 ( .A(n1138), .B(n1137), .Z(n1139) );
  NR2I U1399 ( .A(n1140), .B(n1139), .Z(n1142) );
  ND2I U1400 ( .A(\gpr[12][20] ), .B(n2204), .Z(n1141) );
  ND2I U1401 ( .A(n1142), .B(n1141), .Z(n1143) );
  ND2I U1402 ( .A(n4725), .B(n1143), .Z(n1144) );
  ND2I U1403 ( .A(n1145), .B(n1144), .Z(n1146) );
  NR2I U1404 ( .A(n1147), .B(n1146), .Z(n1157) );
  AO2 U1405 ( .A(\gpr[15][20] ), .B(n1523), .C(n4724), .D(\gpr[3][20] ), .Z(
        n1154) );
  AO2 U1406 ( .A(n1246), .B(\gpr[2][20] ), .C(n1520), .D(\gpr[5][20] ), .Z(
        n1152) );
  ND2I U1407 ( .A(\gpr[13][20] ), .B(n2058), .Z(n1149) );
  ND2I U1408 ( .A(n2174), .B(n1149), .Z(n1150) );
  IVI U1409 ( .A(n1150), .Z(n1151) );
  AN2I U1410 ( .A(n1152), .B(n1151), .Z(n1153) );
  ND2I U1411 ( .A(n1154), .B(n1153), .Z(n1155) );
  IVI U1412 ( .A(n1155), .Z(n1156) );
  ND2I U1413 ( .A(n1157), .B(n1156), .Z(n1158) );
  AN2I U1414 ( .A(n1159), .B(n1158), .Z(rd_data1[20]) );
  ND2I U1415 ( .A(n4723), .B(\gpr[5][15] ), .Z(n1164) );
  ND2I U1416 ( .A(n909), .B(\gpr[3][15] ), .Z(n1163) );
  ND2I U1417 ( .A(n2115), .B(\gpr[2][15] ), .Z(n1160) );
  AN2I U1418 ( .A(n1160), .B(n2174), .Z(n1162) );
  ND2I U1419 ( .A(\gpr[10][15] ), .B(n102), .Z(n1161) );
  ND4P U1420 ( .A(n1164), .B(n1163), .C(n1162), .D(n1161), .Z(n1172) );
  ND2I U1421 ( .A(\gpr[13][15] ), .B(n4718), .Z(n1166) );
  ND2I U1422 ( .A(n4719), .B(\gpr[1][15] ), .Z(n1165) );
  ND2I U1423 ( .A(n1166), .B(n1165), .Z(n1167) );
  IVI U1424 ( .A(n1167), .Z(n1170) );
  ND2I U1425 ( .A(\gpr[4][15] ), .B(n1168), .Z(n1169) );
  ND2I U1426 ( .A(n1170), .B(n1169), .Z(n1171) );
  NR2I U1427 ( .A(n1172), .B(n1171), .Z(n1184) );
  ND2I U1428 ( .A(n4737), .B(\gpr[9][15] ), .Z(n1176) );
  ND2I U1429 ( .A(n1725), .B(\gpr[8][15] ), .Z(n1175) );
  ND2I U1430 ( .A(n1669), .B(\gpr[11][15] ), .Z(n1174) );
  ND2I U1431 ( .A(n2317), .B(\gpr[12][15] ), .Z(n1173) );
  ND4 U1432 ( .A(n1176), .B(n1175), .C(n1174), .D(n1173), .Z(n1182) );
  IVI U1433 ( .A(n1432), .Z(n2172) );
  ND2I U1434 ( .A(\gpr[15][15] ), .B(n2172), .Z(n1180) );
  ND2I U1435 ( .A(n4746), .B(\gpr[6][15] ), .Z(n1179) );
  IVI U1436 ( .A(n1446), .Z(n1791) );
  ND2I U1437 ( .A(n1791), .B(\gpr[7][15] ), .Z(n1178) );
  ND2I U1438 ( .A(n1990), .B(\gpr[14][15] ), .Z(n1177) );
  ND4 U1439 ( .A(n1180), .B(n1179), .C(n1178), .D(n1177), .Z(n1181) );
  NR2I U1440 ( .A(n1182), .B(n1181), .Z(n1183) );
  ND2I U1441 ( .A(n1184), .B(n1183), .Z(n1215) );
  ND2I U1442 ( .A(\gpr[26][15] ), .B(n2207), .Z(n1185) );
  ND2I U1443 ( .A(n272), .B(n1185), .Z(n1187) );
  AN2I U1444 ( .A(\gpr[24][15] ), .B(n1402), .Z(n1186) );
  NR2I U1445 ( .A(n1187), .B(n1186), .Z(n1195) );
  ND2I U1446 ( .A(\gpr[29][15] ), .B(n2268), .Z(n1189) );
  ND2I U1447 ( .A(\gpr[27][15] ), .B(n4703), .Z(n1188) );
  ND2I U1448 ( .A(n1189), .B(n1188), .Z(n1193) );
  ND2I U1449 ( .A(\gpr[31][15] ), .B(n2100), .Z(n1191) );
  ND2I U1450 ( .A(\gpr[28][15] ), .B(n2158), .Z(n1190) );
  ND2I U1451 ( .A(n1191), .B(n1190), .Z(n1192) );
  NR2I U1452 ( .A(n1193), .B(n1192), .Z(n1194) );
  AN2I U1453 ( .A(n1195), .B(n1194), .Z(n1197) );
  ND2I U1454 ( .A(n1952), .B(\gpr[25][15] ), .Z(n1196) );
  ND2I U1455 ( .A(n1197), .B(n273), .Z(n1212) );
  ND2I U1456 ( .A(\gpr[20][15] ), .B(n1424), .Z(n1203) );
  ND2I U1457 ( .A(n4703), .B(\gpr[19][15] ), .Z(n1199) );
  ND2I U1458 ( .A(n2268), .B(\gpr[21][15] ), .Z(n1198) );
  ND2I U1459 ( .A(n1199), .B(n1198), .Z(n1201) );
  AN2I U1460 ( .A(n2100), .B(\gpr[23][15] ), .Z(n1200) );
  NR2I U1461 ( .A(n1201), .B(n1200), .Z(n1202) );
  IVI U1462 ( .A(n1204), .Z(n2159) );
  NR2I U1463 ( .A(n2159), .B(n4862), .Z(n1208) );
  ND2I U1464 ( .A(n1205), .B(\gpr[16][15] ), .Z(n1206) );
  ND2I U1465 ( .A(n4709), .B(n1206), .Z(n1207) );
  NR2I U1466 ( .A(n1208), .B(n1207), .Z(n1210) );
  IVI U1467 ( .A(n1275), .Z(n2231) );
  AO2 U1468 ( .A(n4726), .B(\gpr[18][15] ), .C(n2231), .D(\gpr[17][15] ), .Z(
        n1209) );
  ND2I U1469 ( .A(n237), .B(n211), .Z(n1211) );
  ND2I U1470 ( .A(n1212), .B(n1211), .Z(n1213) );
  IVI U1471 ( .A(n1213), .Z(n1214) );
  AN2I U1472 ( .A(n1215), .B(n1214), .Z(rd_data1[15]) );
  ND2I U1473 ( .A(\gpr[27][14] ), .B(n4703), .Z(n1217) );
  ND2I U1474 ( .A(\gpr[26][14] ), .B(n4726), .Z(n1216) );
  ND2I U1475 ( .A(n1217), .B(n1216), .Z(n1221) );
  ND2I U1476 ( .A(\gpr[28][14] ), .B(n2204), .Z(n1219) );
  ND2I U1477 ( .A(\gpr[31][14] ), .B(n2100), .Z(n1218) );
  ND2I U1478 ( .A(n1219), .B(n1218), .Z(n1220) );
  NR2I U1479 ( .A(n1221), .B(n1220), .Z(n1223) );
  AO2 U1480 ( .A(n2233), .B(\gpr[24][14] ), .C(n1466), .D(\gpr[25][14] ), .Z(
        n1222) );
  ND2I U1481 ( .A(n2020), .B(\gpr[30][14] ), .Z(n1224) );
  AO3 U1482 ( .A(n2022), .B(n4830), .C(n4690), .D(n1224), .Z(n1225) );
  IVI U1483 ( .A(n1225), .Z(n1226) );
  ND2I U1484 ( .A(n238), .B(n1226), .Z(n1238) );
  NR2I U1485 ( .A(n2297), .B(n4860), .Z(n1229) );
  ND2I U1486 ( .A(n2077), .B(\gpr[18][14] ), .Z(n1227) );
  ND2I U1487 ( .A(n4709), .B(n1227), .Z(n1228) );
  NR2I U1488 ( .A(n1229), .B(n1228), .Z(n1236) );
  AO2 U1489 ( .A(n4701), .B(\gpr[21][14] ), .C(n1360), .D(\gpr[17][14] ), .Z(
        n1235) );
  B2IP U1490 ( .A(n1631), .Z1(n1230), .Z2(n2158) );
  IVI U1491 ( .A(n1230), .Z(n2291) );
  ND2I U1492 ( .A(n2291), .B(\gpr[20][14] ), .Z(n1232) );
  ND2I U1493 ( .A(\gpr[22][14] ), .B(n2020), .Z(n1231) );
  AN2I U1494 ( .A(n1232), .B(n1231), .Z(n1234) );
  ND2I U1495 ( .A(n1238), .B(n1237), .Z(n1239) );
  IVI U1496 ( .A(n1239), .Z(n1267) );
  AO2 U1497 ( .A(n2061), .B(\gpr[7][14] ), .C(n2040), .D(\gpr[3][14] ), .Z(
        n1245) );
  ND2I U1498 ( .A(\gpr[4][14] ), .B(n1528), .Z(n1242) );
  ND2I U1499 ( .A(\gpr[1][14] ), .B(n1240), .Z(n1241) );
  ND2I U1500 ( .A(n1242), .B(n1241), .Z(n1243) );
  IVI U1501 ( .A(n1243), .Z(n1244) );
  AN2I U1502 ( .A(n1245), .B(n1244), .Z(n1265) );
  AO2 U1503 ( .A(\gpr[15][14] ), .B(n1523), .C(n104), .D(\gpr[6][14] ), .Z(
        n1264) );
  ND2I U1504 ( .A(n2189), .B(\gpr[2][14] ), .Z(n1247) );
  ND2I U1505 ( .A(n498), .B(n1247), .Z(n1251) );
  ND2I U1506 ( .A(\gpr[13][14] ), .B(n2259), .Z(n1249) );
  ND2I U1507 ( .A(n1520), .B(\gpr[5][14] ), .Z(n1248) );
  ND2I U1508 ( .A(n1249), .B(n1248), .Z(n1250) );
  NR2I U1509 ( .A(n1251), .B(n1250), .Z(n1263) );
  AO2 U1510 ( .A(n2077), .B(\gpr[10][14] ), .C(n1824), .D(\gpr[9][14] ), .Z(
        n1260) );
  ND2I U1511 ( .A(\gpr[8][14] ), .B(n2017), .Z(n1254) );
  ND2I U1512 ( .A(n207), .B(\gpr[14][14] ), .Z(n1253) );
  ND2I U1513 ( .A(n1254), .B(n1253), .Z(n1258) );
  ND2I U1514 ( .A(n4694), .B(\gpr[12][14] ), .Z(n1256) );
  ND2I U1515 ( .A(n4688), .B(\gpr[11][14] ), .Z(n1255) );
  ND2I U1516 ( .A(n1256), .B(n1255), .Z(n1257) );
  NR2I U1517 ( .A(n1258), .B(n1257), .Z(n1259) );
  ND2I U1518 ( .A(n1260), .B(n1259), .Z(n1261) );
  ND2I U1519 ( .A(n4725), .B(n1261), .Z(n1262) );
  ND4P U1520 ( .A(n1265), .B(n1264), .C(n1263), .D(n1262), .Z(n1266) );
  AN2I U1521 ( .A(n1267), .B(n1266), .Z(rd_data1[14]) );
  IVI U1522 ( .A(n1268), .Z(n1384) );
  IVI U1523 ( .A(n1384), .Z(n2155) );
  ND2I U1524 ( .A(n2155), .B(\gpr[16][2] ), .Z(n1270) );
  ND2I U1525 ( .A(n2204), .B(\gpr[20][2] ), .Z(n1269) );
  ND2I U1526 ( .A(n1270), .B(n1269), .Z(n1274) );
  ND2I U1527 ( .A(\gpr[21][2] ), .B(n4701), .Z(n1272) );
  ND2I U1528 ( .A(\gpr[18][2] ), .B(n2077), .Z(n1271) );
  ND2I U1529 ( .A(n1272), .B(n1271), .Z(n1273) );
  NR2I U1530 ( .A(n1274), .B(n1273), .Z(n1285) );
  NR2I U1531 ( .A(n2159), .B(n4763), .Z(n1278) );
  IVI U1532 ( .A(n1275), .Z(n1595) );
  ND2I U1533 ( .A(n1595), .B(\gpr[17][2] ), .Z(n1276) );
  ND2I U1534 ( .A(n2094), .B(n1276), .Z(n1277) );
  NR2I U1535 ( .A(n1278), .B(n1277), .Z(n1283) );
  ND2I U1536 ( .A(n2100), .B(\gpr[23][2] ), .Z(n1280) );
  ND2I U1537 ( .A(n2284), .B(\gpr[19][2] ), .Z(n1279) );
  ND2I U1538 ( .A(n1280), .B(n1279), .Z(n1281) );
  IVI U1539 ( .A(n1281), .Z(n1282) );
  AN2I U1540 ( .A(n1283), .B(n1282), .Z(n1284) );
  ND2I U1541 ( .A(n1285), .B(n1284), .Z(n1301) );
  ND2I U1542 ( .A(\gpr[31][2] ), .B(n2100), .Z(n1287) );
  ND2I U1543 ( .A(\gpr[27][2] ), .B(n2284), .Z(n1286) );
  ND2I U1544 ( .A(n1287), .B(n1286), .Z(n1291) );
  ND2I U1545 ( .A(\gpr[28][2] ), .B(n2158), .Z(n1289) );
  ND2I U1546 ( .A(\gpr[24][2] ), .B(n2155), .Z(n1288) );
  ND2I U1547 ( .A(n1289), .B(n1288), .Z(n1290) );
  NR2I U1548 ( .A(n1291), .B(n1290), .Z(n1299) );
  NR2I U1549 ( .A(n2159), .B(n4842), .Z(n1294) );
  ND2I U1550 ( .A(n1938), .B(\gpr[25][2] ), .Z(n1292) );
  ND2I U1551 ( .A(n2079), .B(n1292), .Z(n1293) );
  NR2I U1552 ( .A(n1294), .B(n1293), .Z(n1296) );
  AO2P U1553 ( .A(n4702), .B(\gpr[26][2] ), .C(n2268), .D(\gpr[29][2] ), .Z(
        n1295) );
  ND2I U1554 ( .A(n1296), .B(n1295), .Z(n1297) );
  IVI U1555 ( .A(n1297), .Z(n1298) );
  ND2I U1556 ( .A(n1299), .B(n1298), .Z(n1300) );
  ND2I U1557 ( .A(n1301), .B(n1300), .Z(n1302) );
  IVI U1558 ( .A(n1302), .Z(n1331) );
  ND2I U1559 ( .A(\gpr[15][2] ), .B(n2172), .Z(n1306) );
  ND2I U1560 ( .A(n104), .B(\gpr[6][2] ), .Z(n1305) );
  ND2I U1561 ( .A(n1791), .B(\gpr[7][2] ), .Z(n1304) );
  IVI U1562 ( .A(n1606), .Z(n2126) );
  ND2I U1563 ( .A(n2126), .B(\gpr[14][2] ), .Z(n1303) );
  ND4 U1564 ( .A(n1306), .B(n1305), .C(n1304), .D(n1303), .Z(n1317) );
  ND2I U1565 ( .A(n1307), .B(\gpr[8][2] ), .Z(n1315) );
  ND2I U1566 ( .A(\gpr[13][2] ), .B(n2188), .Z(n1314) );
  ND2I U1567 ( .A(n2256), .B(\gpr[2][2] ), .Z(n1312) );
  IVI U1568 ( .A(n1308), .Z(n2133) );
  ND2I U1569 ( .A(n2133), .B(\gpr[11][2] ), .Z(n1309) );
  ND2I U1570 ( .A(n2174), .B(n1309), .Z(n1310) );
  IVI U1571 ( .A(n1310), .Z(n1311) );
  AN2I U1572 ( .A(n1312), .B(n1311), .Z(n1313) );
  ND2I U1573 ( .A(n1315), .B(n239), .Z(n1316) );
  NR2I U1574 ( .A(n1317), .B(n1316), .Z(n1329) );
  ND2I U1575 ( .A(\gpr[1][2] ), .B(n4719), .Z(n1319) );
  ND2I U1576 ( .A(n1859), .B(\gpr[3][2] ), .Z(n1318) );
  ND2I U1577 ( .A(n2303), .B(\gpr[4][2] ), .Z(n1325) );
  OR2I U1578 ( .A(n1320), .B(n4940), .Z(n1322) );
  ND2I U1579 ( .A(\gpr[5][2] ), .B(n4723), .Z(n1321) );
  ND2I U1580 ( .A(n1322), .B(n1321), .Z(n1323) );
  IVI U1581 ( .A(n1323), .Z(n1324) );
  ND2I U1582 ( .A(n1325), .B(n1324), .Z(n1326) );
  NR2I U1583 ( .A(n1327), .B(n1326), .Z(n1328) );
  ND2I U1584 ( .A(n1329), .B(n1328), .Z(n1330) );
  AN2I U1585 ( .A(n1331), .B(n1330), .Z(rd_data1[2]) );
  ND2I U1586 ( .A(\gpr[4][8] ), .B(n1528), .Z(n1339) );
  ND2I U1587 ( .A(n1727), .B(\gpr[2][8] ), .Z(n1332) );
  ND2I U1588 ( .A(n498), .B(n1332), .Z(n1337) );
  ND2I U1589 ( .A(\gpr[1][8] ), .B(n2320), .Z(n1335) );
  AN2I U1590 ( .A(n2307), .B(\gpr[13][8] ), .Z(n1333) );
  ND2I U1591 ( .A(n4701), .B(n1333), .Z(n1334) );
  ND2I U1592 ( .A(n1335), .B(n1334), .Z(n1336) );
  NR2I U1593 ( .A(n1337), .B(n1336), .Z(n1338) );
  ND2I U1594 ( .A(n1339), .B(n1338), .Z(n1345) );
  ND2I U1595 ( .A(n104), .B(\gpr[6][8] ), .Z(n1343) );
  ND2I U1596 ( .A(n1791), .B(\gpr[7][8] ), .Z(n1341) );
  ND2I U1597 ( .A(\gpr[5][8] ), .B(n1520), .Z(n1340) );
  AN2I U1598 ( .A(n1341), .B(n1340), .Z(n1342) );
  ND2I U1599 ( .A(n1343), .B(n1342), .Z(n1344) );
  NR2I U1600 ( .A(n1345), .B(n1344), .Z(n1348) );
  AO2 U1601 ( .A(\gpr[15][8] ), .B(n4745), .C(n1346), .D(\gpr[3][8] ), .Z(
        n1347) );
  AN2I U1602 ( .A(n1348), .B(n1347), .Z(n1359) );
  AO2 U1603 ( .A(n4726), .B(\gpr[10][8] ), .C(n2231), .D(\gpr[9][8] ), .Z(
        n1356) );
  ND2I U1604 ( .A(\gpr[8][8] ), .B(n1205), .Z(n1350) );
  ND2I U1605 ( .A(\gpr[14][8] ), .B(n862), .Z(n1349) );
  ND2I U1606 ( .A(n1350), .B(n1349), .Z(n1354) );
  ND2I U1607 ( .A(n4688), .B(\gpr[11][8] ), .Z(n1352) );
  ND2I U1608 ( .A(n2158), .B(\gpr[12][8] ), .Z(n1351) );
  ND2I U1609 ( .A(n1352), .B(n1351), .Z(n1353) );
  NR2I U1610 ( .A(n1354), .B(n1353), .Z(n1355) );
  ND2I U1611 ( .A(n1356), .B(n1355), .Z(n1357) );
  ND2I U1612 ( .A(rd_addr1[3]), .B(n1357), .Z(n1358) );
  ND2I U1613 ( .A(n1359), .B(n1358), .Z(n1395) );
  ND2I U1614 ( .A(\gpr[20][8] ), .B(n2158), .Z(n1362) );
  ND2I U1615 ( .A(\gpr[17][8] ), .B(n1360), .Z(n1361) );
  AN2I U1616 ( .A(n1362), .B(n1361), .Z(n1365) );
  IVI U1617 ( .A(n1363), .Z(n1402) );
  ND2I U1618 ( .A(n1365), .B(n1364), .Z(n1366) );
  IVI U1619 ( .A(n1366), .Z(n1375) );
  AO2 U1620 ( .A(n2157), .B(\gpr[21][8] ), .C(n4703), .D(\gpr[19][8] ), .Z(
        n1372) );
  NR2I U1621 ( .A(n1765), .B(n4850), .Z(n1370) );
  ND2I U1622 ( .A(n2207), .B(\gpr[18][8] ), .Z(n1368) );
  ND2I U1623 ( .A(n2094), .B(n1368), .Z(n1369) );
  NR2I U1624 ( .A(n1370), .B(n1369), .Z(n1371) );
  ND2I U1625 ( .A(n1372), .B(n1371), .Z(n1373) );
  IVI U1626 ( .A(n1373), .Z(n1374) );
  ND2I U1627 ( .A(n1375), .B(n1374), .Z(n1392) );
  AO2 U1628 ( .A(n4726), .B(\gpr[26][8] ), .C(n4703), .D(\gpr[27][8] ), .Z(
        n1379) );
  ND2I U1629 ( .A(n2020), .B(\gpr[30][8] ), .Z(n1376) );
  AO3 U1630 ( .A(n4693), .B(n4828), .C(n2079), .D(n1376), .Z(n1377) );
  IVI U1631 ( .A(n1377), .Z(n1378) );
  ND2I U1632 ( .A(n1379), .B(n1378), .Z(n1380) );
  IVI U1633 ( .A(n1380), .Z(n1390) );
  ND2I U1634 ( .A(\gpr[28][8] ), .B(n2204), .Z(n1382) );
  ND2I U1635 ( .A(\gpr[31][8] ), .B(n2100), .Z(n1381) );
  AN2I U1636 ( .A(n1382), .B(n1381), .Z(n1387) );
  ND2I U1637 ( .A(\gpr[25][8] ), .B(n1383), .Z(n1386) );
  IVI U1638 ( .A(n1384), .Z(n2271) );
  ND2I U1639 ( .A(\gpr[24][8] ), .B(n2271), .Z(n1385) );
  ND2I U1640 ( .A(n1387), .B(n274), .Z(n1388) );
  IVI U1641 ( .A(n1388), .Z(n1389) );
  ND2I U1642 ( .A(n1390), .B(n1389), .Z(n1391) );
  ND2I U1643 ( .A(n1392), .B(n1391), .Z(n1393) );
  IVI U1644 ( .A(n1393), .Z(n1394) );
  ND2I U1645 ( .A(n1395), .B(n1394), .Z(n1396) );
  IVI U1646 ( .A(n1396), .Z(rd_data1[8]) );
  AO2 U1647 ( .A(n2077), .B(\gpr[26][6] ), .C(n2157), .D(\gpr[29][6] ), .Z(
        n1410) );
  NR2I U1648 ( .A(n1810), .B(n4847), .Z(n1399) );
  ND2I U1649 ( .A(n1595), .B(\gpr[25][6] ), .Z(n1397) );
  ND2I U1650 ( .A(n4690), .B(n1397), .Z(n1398) );
  NR2I U1651 ( .A(n1399), .B(n1398), .Z(n1408) );
  ND2I U1652 ( .A(n2100), .B(\gpr[31][6] ), .Z(n1401) );
  ND2I U1653 ( .A(n2284), .B(\gpr[27][6] ), .Z(n1400) );
  ND2I U1654 ( .A(n1401), .B(n1400), .Z(n1406) );
  ND2I U1655 ( .A(\gpr[28][6] ), .B(n2099), .Z(n1404) );
  ND2I U1656 ( .A(\gpr[24][6] ), .B(n1402), .Z(n1403) );
  ND2I U1657 ( .A(n1404), .B(n1403), .Z(n1405) );
  NR2I U1658 ( .A(n1406), .B(n1405), .Z(n1407) );
  AN2I U1659 ( .A(n1408), .B(n1407), .Z(n1409) );
  ND2I U1660 ( .A(n1410), .B(n1409), .Z(n1428) );
  ND2I U1661 ( .A(n2292), .B(\gpr[21][6] ), .Z(n1415) );
  ND2I U1662 ( .A(\gpr[18][6] ), .B(n2077), .Z(n1412) );
  ND2I U1663 ( .A(\gpr[23][6] ), .B(n2100), .Z(n1411) );
  ND2I U1664 ( .A(n1412), .B(n1411), .Z(n1413) );
  IVI U1665 ( .A(n1413), .Z(n1414) );
  ND2I U1666 ( .A(n1415), .B(n1414), .Z(n1423) );
  NR2I U1667 ( .A(n4687), .B(n4846), .Z(n1418) );
  ND2I U1668 ( .A(n2004), .B(\gpr[16][6] ), .Z(n1416) );
  ND2I U1669 ( .A(n2094), .B(n1416), .Z(n1417) );
  NR2I U1670 ( .A(n1418), .B(n1417), .Z(n1421) );
  ND2I U1671 ( .A(\gpr[17][6] ), .B(n1952), .Z(n1420) );
  ND2I U1672 ( .A(\gpr[19][6] ), .B(n2284), .Z(n1419) );
  ND2I U1673 ( .A(n1421), .B(n275), .Z(n1422) );
  NR2I U1674 ( .A(n1423), .B(n1422), .Z(n1426) );
  ND2I U1675 ( .A(n1424), .B(\gpr[20][6] ), .Z(n1425) );
  ND2I U1676 ( .A(n1426), .B(n1425), .Z(n1427) );
  ND2I U1677 ( .A(n4718), .B(\gpr[13][6] ), .Z(n1431) );
  ND2I U1678 ( .A(\gpr[1][6] ), .B(n4719), .Z(n1430) );
  IVI U1679 ( .A(n1148), .Z(n1727) );
  ND2I U1680 ( .A(n1727), .B(\gpr[2][6] ), .Z(n1429) );
  ND2I U1681 ( .A(n4732), .B(\gpr[4][6] ), .Z(n1442) );
  IVI U1682 ( .A(n1432), .Z(n2312) );
  ND2I U1683 ( .A(n2312), .B(\gpr[15][6] ), .Z(n1433) );
  IVI U1684 ( .A(n1433), .Z(n1438) );
  IVI U1685 ( .A(n1434), .Z(n2110) );
  ND2I U1686 ( .A(n2110), .B(\gpr[3][6] ), .Z(n1436) );
  ND2I U1687 ( .A(n2132), .B(\gpr[12][6] ), .Z(n1435) );
  ND2I U1688 ( .A(n1436), .B(n1435), .Z(n1437) );
  NR2I U1689 ( .A(n1438), .B(n1437), .Z(n1440) );
  ND2I U1690 ( .A(n1797), .B(\gpr[10][6] ), .Z(n1439) );
  AN2I U1691 ( .A(n1440), .B(n1439), .Z(n1441) );
  ND2I U1692 ( .A(n1442), .B(n1441), .Z(n1457) );
  ND2I U1693 ( .A(n4737), .B(\gpr[9][6] ), .Z(n1444) );
  ND2I U1694 ( .A(n2126), .B(\gpr[14][6] ), .Z(n1443) );
  ND2I U1695 ( .A(n4738), .B(\gpr[8][6] ), .Z(n1445) );
  IVI U1696 ( .A(n1445), .Z(n1454) );
  ND2I U1697 ( .A(n2133), .B(\gpr[11][6] ), .Z(n1448) );
  OR2I U1698 ( .A(n1446), .B(n5042), .Z(n1447) );
  AN2I U1699 ( .A(n1448), .B(n1447), .Z(n1450) );
  ND2I U1700 ( .A(n104), .B(\gpr[6][6] ), .Z(n1449) );
  AN2I U1701 ( .A(n1450), .B(n1449), .Z(n1452) );
  ND2I U1702 ( .A(n4723), .B(\gpr[5][6] ), .Z(n1451) );
  ND2I U1703 ( .A(n1452), .B(n1451), .Z(n1453) );
  NR2I U1704 ( .A(n1454), .B(n1453), .Z(n1455) );
  ND2I U1705 ( .A(n240), .B(n1455), .Z(n1456) );
  NR2I U1706 ( .A(n1457), .B(n1456), .Z(n1458) );
  ND2I U1707 ( .A(n212), .B(n1458), .Z(n1459) );
  AN2I U1708 ( .A(n241), .B(n1459), .Z(rd_data1[6]) );
  ND2I U1709 ( .A(\gpr[27][10] ), .B(n4703), .Z(n1461) );
  ND2I U1710 ( .A(\gpr[26][10] ), .B(n4726), .Z(n1460) );
  ND2I U1711 ( .A(n1461), .B(n1460), .Z(n1465) );
  ND2I U1712 ( .A(\gpr[28][10] ), .B(n2099), .Z(n1463) );
  ND2I U1713 ( .A(\gpr[31][10] ), .B(n2100), .Z(n1462) );
  ND2I U1714 ( .A(n1463), .B(n1462), .Z(n1464) );
  NR2I U1715 ( .A(n1465), .B(n1464), .Z(n1474) );
  ND2I U1716 ( .A(\gpr[25][10] ), .B(n1466), .Z(n1468) );
  ND2I U1717 ( .A(\gpr[24][10] ), .B(n2017), .Z(n1467) );
  AN2I U1718 ( .A(n1468), .B(n1467), .Z(n1473) );
  B3IP U1719 ( .A(n1469), .Z1(n1752), .Z2(n1651) );
  ND2I U1720 ( .A(n2020), .B(\gpr[30][10] ), .Z(n1470) );
  AO3 U1721 ( .A(n1651), .B(n4829), .C(n2079), .D(n1470), .Z(n1471) );
  IVI U1722 ( .A(n1471), .Z(n1472) );
  ND2I U1723 ( .A(n1474), .B(n242), .Z(n1488) );
  ND2I U1724 ( .A(\gpr[16][10] ), .B(n1598), .Z(n1476) );
  ND2I U1725 ( .A(\gpr[22][10] ), .B(n207), .Z(n1475) );
  ND2I U1726 ( .A(n1476), .B(n1475), .Z(n1480) );
  ND2I U1727 ( .A(\gpr[20][10] ), .B(n2099), .Z(n1478) );
  ND2I U1728 ( .A(\gpr[19][10] ), .B(n4703), .Z(n1477) );
  ND2I U1729 ( .A(n1478), .B(n1477), .Z(n1479) );
  NR2I U1730 ( .A(n1480), .B(n1479), .Z(n1486) );
  NR2I U1731 ( .A(n2297), .B(n4853), .Z(n1483) );
  ND2I U1732 ( .A(n4702), .B(\gpr[18][10] ), .Z(n1481) );
  ND2I U1733 ( .A(n2094), .B(n1481), .Z(n1482) );
  NR2I U1734 ( .A(n1483), .B(n1482), .Z(n1485) );
  AO2P U1735 ( .A(n2268), .B(\gpr[21][10] ), .C(n1952), .D(\gpr[17][10] ), .Z(
        n1484) );
  ND2I U1736 ( .A(n1486), .B(n243), .Z(n1487) );
  AN2I U1737 ( .A(n1488), .B(n1487), .Z(n1519) );
  ND2I U1738 ( .A(n1528), .B(\gpr[4][10] ), .Z(n1491) );
  AN2I U1739 ( .A(n2307), .B(\gpr[13][10] ), .Z(n1489) );
  ND2I U1740 ( .A(n2268), .B(n1489), .Z(n1490) );
  ND2I U1741 ( .A(n1491), .B(n1490), .Z(n1495) );
  ND2I U1742 ( .A(n105), .B(\gpr[6][10] ), .Z(n1493) );
  ND2I U1743 ( .A(n4723), .B(\gpr[5][10] ), .Z(n1492) );
  ND2I U1744 ( .A(n1493), .B(n1492), .Z(n1494) );
  NR2I U1745 ( .A(n1495), .B(n1494), .Z(n1505) );
  ND2I U1746 ( .A(n2114), .B(\gpr[7][10] ), .Z(n1497) );
  ND2I U1747 ( .A(\gpr[2][10] ), .B(n1727), .Z(n1496) );
  AN2I U1748 ( .A(n1497), .B(n1496), .Z(n1502) );
  ND2I U1749 ( .A(n1846), .B(\gpr[15][10] ), .Z(n1501) );
  ND2I U1750 ( .A(\gpr[1][10] ), .B(n2320), .Z(n1498) );
  ND2I U1751 ( .A(\gpr[3][10] ), .B(n1089), .Z(n1500) );
  ND4P U1752 ( .A(n1502), .B(n1501), .C(n262), .D(n1500), .Z(n1503) );
  IVI U1753 ( .A(n1503), .Z(n1504) );
  ND2I U1754 ( .A(n1505), .B(n1504), .Z(n1506) );
  IVI U1755 ( .A(n1506), .Z(n1517) );
  AO2 U1756 ( .A(n2077), .B(\gpr[10][10] ), .C(n1647), .D(\gpr[9][10] ), .Z(
        n1514) );
  ND2I U1757 ( .A(n2291), .B(\gpr[12][10] ), .Z(n1511) );
  ND2I U1758 ( .A(\gpr[14][10] ), .B(n862), .Z(n1510) );
  ND2I U1759 ( .A(n4688), .B(\gpr[11][10] ), .Z(n1509) );
  ND2I U1760 ( .A(\gpr[8][10] ), .B(n2155), .Z(n1508) );
  ND4P U1761 ( .A(n1511), .B(n1510), .C(n1509), .D(n1508), .Z(n1512) );
  IVI U1762 ( .A(n1512), .Z(n1513) );
  ND2I U1763 ( .A(n1514), .B(n1513), .Z(n1515) );
  ND2I U1764 ( .A(n1515), .B(n2307), .Z(n1516) );
  ND2I U1765 ( .A(n1517), .B(n1516), .Z(n1518) );
  AN2I U1766 ( .A(n1519), .B(n1518), .Z(rd_data1[10]) );
  ND2I U1767 ( .A(\gpr[1][24] ), .B(n2320), .Z(n1522) );
  ND2I U1768 ( .A(\gpr[5][24] ), .B(n1520), .Z(n1521) );
  ND2I U1769 ( .A(n1089), .B(\gpr[3][24] ), .Z(n1525) );
  ND2I U1770 ( .A(n1523), .B(\gpr[15][24] ), .Z(n1524) );
  AN2I U1771 ( .A(n1525), .B(n1524), .Z(n1526) );
  ND2I U1772 ( .A(n2115), .B(\gpr[2][24] ), .Z(n1527) );
  ND2I U1773 ( .A(n2174), .B(n1527), .Z(n1532) );
  ND2I U1774 ( .A(n1528), .B(\gpr[4][24] ), .Z(n1530) );
  ND2I U1775 ( .A(\gpr[13][24] ), .B(n2058), .Z(n1529) );
  ND2I U1776 ( .A(n1530), .B(n1529), .Z(n1531) );
  NR2I U1777 ( .A(n1532), .B(n1531), .Z(n1543) );
  ND2I U1778 ( .A(n4694), .B(\gpr[12][24] ), .Z(n1540) );
  ND2I U1779 ( .A(n4688), .B(\gpr[11][24] ), .Z(n1534) );
  ND2I U1780 ( .A(\gpr[9][24] ), .B(n2276), .Z(n1533) );
  AN2I U1781 ( .A(n1534), .B(n1533), .Z(n1539) );
  ND2I U1782 ( .A(\gpr[8][24] ), .B(n2271), .Z(n1538) );
  ND2I U1783 ( .A(n600), .B(\gpr[14][24] ), .Z(n1537) );
  ND2I U1784 ( .A(\gpr[10][24] ), .B(n1535), .Z(n1536) );
  ND4P U1785 ( .A(n1540), .B(n1539), .C(n1538), .D(n223), .Z(n1541) );
  ND2I U1786 ( .A(n2307), .B(n1541), .Z(n1542) );
  B3IP U1787 ( .A(n1545), .Z1(n4701), .Z2(n2006) );
  IVI U1788 ( .A(n1547), .Z(n1552) );
  ND2I U1789 ( .A(\gpr[23][24] ), .B(n4704), .Z(n1549) );
  ND2I U1790 ( .A(\gpr[18][24] ), .B(n2207), .Z(n1548) );
  ND2I U1791 ( .A(n1549), .B(n1548), .Z(n1550) );
  IVI U1792 ( .A(n1550), .Z(n1551) );
  AN2I U1793 ( .A(n1552), .B(n1551), .Z(n1560) );
  ND2I U1794 ( .A(\gpr[17][24] ), .B(n1383), .Z(n1555) );
  ND2I U1795 ( .A(\gpr[16][24] ), .B(n2271), .Z(n1554) );
  ND2I U1796 ( .A(\gpr[19][24] ), .B(n2284), .Z(n1557) );
  ND2I U1797 ( .A(\gpr[20][24] ), .B(n4694), .Z(n1556) );
  ND2I U1798 ( .A(n1557), .B(n1556), .Z(n1558) );
  NR2I U1799 ( .A(n245), .B(n1558), .Z(n1559) );
  ND2I U1800 ( .A(n1560), .B(n1559), .Z(n1579) );
  ND2I U1801 ( .A(\gpr[27][24] ), .B(n2284), .Z(n1562) );
  ND2I U1802 ( .A(\gpr[30][24] ), .B(n600), .Z(n1561) );
  ND2I U1803 ( .A(n1562), .B(n1561), .Z(n1569) );
  ND2I U1804 ( .A(\gpr[25][24] ), .B(n2047), .Z(n1564) );
  ND2I U1805 ( .A(\gpr[29][24] ), .B(n2268), .Z(n1563) );
  AN2I U1806 ( .A(n1564), .B(n1563), .Z(n1567) );
  NR2I U1807 ( .A(n2297), .B(n4808), .Z(n1565) );
  IVI U1808 ( .A(n1565), .Z(n1566) );
  ND2I U1809 ( .A(n1567), .B(n1566), .Z(n1568) );
  NR2I U1810 ( .A(n1569), .B(n1568), .Z(n1577) );
  ND2I U1811 ( .A(\gpr[28][24] ), .B(n2158), .Z(n1571) );
  ND2I U1812 ( .A(\gpr[24][24] ), .B(n1762), .Z(n1570) );
  AN2I U1813 ( .A(n1571), .B(n1570), .Z(n1575) );
  ND2I U1814 ( .A(n2207), .B(\gpr[26][24] ), .Z(n1572) );
  ND2I U1815 ( .A(n4690), .B(n1572), .Z(n1573) );
  IVI U1816 ( .A(n1573), .Z(n1574) );
  AN2I U1817 ( .A(n1575), .B(n1574), .Z(n1576) );
  ND2I U1818 ( .A(n1577), .B(n1576), .Z(n1578) );
  AN2I U1819 ( .A(n1579), .B(n1578), .Z(n1580) );
  AN2I U1820 ( .A(n1581), .B(n1580), .Z(rd_data1[24]) );
  AO2 U1821 ( .A(n2077), .B(\gpr[18][5] ), .C(n2268), .D(\gpr[21][5] ), .Z(
        n1590) );
  ND2I U1822 ( .A(n1595), .B(\gpr[17][5] ), .Z(n1582) );
  ND2I U1823 ( .A(\gpr[20][5] ), .B(n4694), .Z(n1587) );
  ND2I U1824 ( .A(\gpr[16][5] ), .B(n1583), .Z(n1586) );
  ND2I U1825 ( .A(\gpr[23][5] ), .B(n2100), .Z(n1585) );
  ND2I U1826 ( .A(\gpr[19][5] ), .B(n2216), .Z(n1584) );
  ND4P U1827 ( .A(n1587), .B(n1586), .C(n1585), .D(n1584), .Z(n1588) );
  AO2 U1828 ( .A(n2077), .B(\gpr[26][5] ), .C(n2157), .D(\gpr[29][5] ), .Z(
        n1605) );
  ND2I U1829 ( .A(n2020), .B(\gpr[30][5] ), .Z(n1591) );
  AN2I U1830 ( .A(n2079), .B(n1591), .Z(n1593) );
  ND2I U1831 ( .A(n2204), .B(\gpr[28][5] ), .Z(n1592) );
  ND2I U1832 ( .A(n1593), .B(n1592), .Z(n1594) );
  IVI U1833 ( .A(n1594), .Z(n1604) );
  ND2I U1834 ( .A(n2216), .B(\gpr[27][5] ), .Z(n1597) );
  ND2I U1835 ( .A(\gpr[25][5] ), .B(n1595), .Z(n1596) );
  ND2I U1836 ( .A(n1597), .B(n1596), .Z(n1602) );
  ND2I U1837 ( .A(\gpr[24][5] ), .B(n1598), .Z(n1600) );
  ND2I U1838 ( .A(n2100), .B(\gpr[31][5] ), .Z(n1599) );
  ND2I U1839 ( .A(n1600), .B(n1599), .Z(n1601) );
  NR2I U1840 ( .A(n1602), .B(n1601), .Z(n1603) );
  ND2I U1841 ( .A(n2125), .B(\gpr[9][5] ), .Z(n1608) );
  IVI U1842 ( .A(n1606), .Z(n4748) );
  ND2I U1843 ( .A(n4748), .B(\gpr[14][5] ), .Z(n1607) );
  ND2I U1844 ( .A(n1608), .B(n1607), .Z(n1614) );
  ND2I U1845 ( .A(n4723), .B(\gpr[5][5] ), .Z(n1613) );
  ND2I U1846 ( .A(n102), .B(\gpr[10][5] ), .Z(n1612) );
  ND2I U1847 ( .A(\gpr[15][5] ), .B(n2172), .Z(n1611) );
  ND2I U1848 ( .A(n1669), .B(\gpr[11][5] ), .Z(n1609) );
  ND2I U1849 ( .A(n106), .B(\gpr[12][5] ), .Z(n1610) );
  ND2I U1850 ( .A(n1725), .B(\gpr[8][5] ), .Z(n1616) );
  ND2I U1851 ( .A(\gpr[1][5] ), .B(n4719), .Z(n1615) );
  ND2I U1852 ( .A(n1616), .B(n1615), .Z(n1617) );
  ND2I U1853 ( .A(n4724), .B(\gpr[3][5] ), .Z(n1622) );
  ND2I U1854 ( .A(n4747), .B(\gpr[7][5] ), .Z(n1620) );
  ND2I U1855 ( .A(n1618), .B(\gpr[2][5] ), .Z(n1619) );
  AN2I U1856 ( .A(n1620), .B(n1619), .Z(n1621) );
  ND2I U1857 ( .A(n1622), .B(n1621), .Z(n1626) );
  ND2I U1858 ( .A(n104), .B(\gpr[6][5] ), .Z(n1624) );
  ND2I U1859 ( .A(\gpr[13][5] ), .B(n4718), .Z(n1623) );
  ND2I U1860 ( .A(n1624), .B(n1623), .Z(n1625) );
  NR2I U1861 ( .A(n1626), .B(n1625), .Z(n1628) );
  ND2I U1862 ( .A(n4732), .B(\gpr[4][5] ), .Z(n1627) );
  ND2I U1863 ( .A(\gpr[16][27] ), .B(n4686), .Z(n1630) );
  ND2I U1864 ( .A(\gpr[23][27] ), .B(n2215), .Z(n1629) );
  AN2I U1865 ( .A(n1630), .B(n1629), .Z(n1636) );
  B2IP U1866 ( .A(n1631), .Z1(n1633), .Z2(n2099) );
  ND2I U1867 ( .A(n2020), .B(\gpr[22][27] ), .Z(n1632) );
  AO3 U1868 ( .A(n1633), .B(n4877), .C(n2094), .D(n1632), .Z(n1634) );
  IVI U1869 ( .A(n1634), .Z(n1635) );
  ND2I U1870 ( .A(\gpr[19][27] ), .B(n2216), .Z(n1638) );
  ND2I U1871 ( .A(\gpr[17][27] ), .B(n1466), .Z(n1637) );
  AN2I U1872 ( .A(n1638), .B(n1637), .Z(n1640) );
  AO2 U1873 ( .A(n4702), .B(\gpr[18][27] ), .C(n2157), .D(\gpr[21][27] ), .Z(
        n1639) );
  ND2I U1874 ( .A(n246), .B(n214), .Z(n1656) );
  ND2I U1875 ( .A(\gpr[28][27] ), .B(n2291), .Z(n1642) );
  ND2I U1876 ( .A(\gpr[30][27] ), .B(n600), .Z(n1641) );
  AN2I U1877 ( .A(n1642), .B(n1641), .Z(n1646) );
  ND2I U1878 ( .A(n2216), .B(\gpr[27][27] ), .Z(n1644) );
  ND2I U1879 ( .A(\gpr[26][27] ), .B(n4726), .Z(n1643) );
  AN2I U1880 ( .A(n1644), .B(n1643), .Z(n1645) );
  ND2I U1881 ( .A(\gpr[25][27] ), .B(n1647), .Z(n1649) );
  ND2I U1882 ( .A(\gpr[24][27] ), .B(n2017), .Z(n1648) );
  ND2I U1883 ( .A(n2275), .B(\gpr[31][27] ), .Z(n1650) );
  AO3 U1884 ( .A(n1651), .B(n4834), .C(n2079), .D(n1650), .Z(n1652) );
  IVI U1885 ( .A(n1652), .Z(n1653) );
  AN2I U1886 ( .A(n276), .B(n1653), .Z(n1654) );
  ND2I U1887 ( .A(n247), .B(n1654), .Z(n1655) );
  AN2I U1888 ( .A(n1656), .B(n1655), .Z(n1692) );
  ND2I U1889 ( .A(n2328), .B(\gpr[10][27] ), .Z(n1662) );
  ND2I U1890 ( .A(n1791), .B(\gpr[7][27] ), .Z(n1659) );
  ND2I U1891 ( .A(\gpr[3][27] ), .B(n1346), .Z(n1658) );
  ND2I U1892 ( .A(n1846), .B(\gpr[15][27] ), .Z(n1657) );
  ND4P U1893 ( .A(n1659), .B(n498), .C(n1658), .D(n1657), .Z(n1660) );
  IVI U1894 ( .A(n1660), .Z(n1661) );
  AN2I U1895 ( .A(n1662), .B(n1661), .Z(n1667) );
  ND2I U1896 ( .A(n4723), .B(\gpr[5][27] ), .Z(n1664) );
  ND2I U1897 ( .A(\gpr[4][27] ), .B(n2303), .Z(n1663) );
  ND2I U1898 ( .A(n1664), .B(n1663), .Z(n1665) );
  IVI U1899 ( .A(n1665), .Z(n1666) );
  ND2I U1900 ( .A(n1667), .B(n1666), .Z(n1668) );
  IVI U1901 ( .A(n1668), .Z(n1690) );
  ND2I U1902 ( .A(n4740), .B(\gpr[12][27] ), .Z(n1674) );
  ND2I U1903 ( .A(n1669), .B(\gpr[11][27] ), .Z(n1672) );
  ND2I U1904 ( .A(n1670), .B(\gpr[2][27] ), .Z(n1671) );
  AN2I U1905 ( .A(n1672), .B(n1671), .Z(n1673) );
  ND2I U1906 ( .A(n1674), .B(n1673), .Z(n1675) );
  IVI U1907 ( .A(n1675), .Z(n1677) );
  ND2I U1908 ( .A(\gpr[13][27] ), .B(n4718), .Z(n1676) );
  ND2I U1909 ( .A(n1677), .B(n1676), .Z(n1681) );
  ND2I U1910 ( .A(n4737), .B(\gpr[9][27] ), .Z(n1679) );
  ND2I U1911 ( .A(\gpr[1][27] ), .B(n4719), .Z(n1678) );
  ND2I U1912 ( .A(n1679), .B(n1678), .Z(n1680) );
  NR2I U1913 ( .A(n1681), .B(n1680), .Z(n1688) );
  ND2I U1914 ( .A(n4738), .B(\gpr[8][27] ), .Z(n1685) );
  ND2I U1915 ( .A(n2126), .B(\gpr[14][27] ), .Z(n1683) );
  ND2I U1916 ( .A(n4746), .B(\gpr[6][27] ), .Z(n1682) );
  AN2I U1917 ( .A(n1683), .B(n1682), .Z(n1684) );
  ND2I U1918 ( .A(n1685), .B(n1684), .Z(n1686) );
  IVI U1919 ( .A(n1686), .Z(n1687) );
  AN2I U1920 ( .A(n1688), .B(n1687), .Z(n1689) );
  ND2I U1921 ( .A(n1690), .B(n1689), .Z(n1691) );
  AN2I U1922 ( .A(n1692), .B(n1691), .Z(rd_data1[27]) );
  ND2I U1923 ( .A(\gpr[17][21] ), .B(n206), .Z(n1694) );
  ND2I U1924 ( .A(n2292), .B(\gpr[21][21] ), .Z(n1693) );
  ND2I U1925 ( .A(n1694), .B(n1693), .Z(n1695) );
  IVI U1926 ( .A(n1695), .Z(n1697) );
  ND2I U1927 ( .A(\gpr[23][21] ), .B(n2215), .Z(n1696) );
  ND2I U1928 ( .A(n1697), .B(n1696), .Z(n1703) );
  ND2I U1929 ( .A(\gpr[18][21] ), .B(n2207), .Z(n1699) );
  ND2I U1930 ( .A(\gpr[19][21] ), .B(n4703), .Z(n1698) );
  AN2I U1931 ( .A(n1699), .B(n1698), .Z(n1701) );
  ND2I U1932 ( .A(\gpr[16][21] ), .B(n2233), .Z(n1700) );
  ND2I U1933 ( .A(n1701), .B(n1700), .Z(n1702) );
  NR2I U1934 ( .A(n1703), .B(n1702), .Z(n1704) );
  ND2I U1935 ( .A(n277), .B(n1704), .Z(n1711) );
  ND2I U1936 ( .A(n2215), .B(\gpr[31][21] ), .Z(n1705) );
  ND2I U1937 ( .A(n1705), .B(n278), .Z(n1708) );
  ND2I U1938 ( .A(\gpr[29][21] ), .B(n2292), .Z(n1707) );
  ND2I U1939 ( .A(\gpr[28][21] ), .B(n2158), .Z(n1706) );
  ND2I U1940 ( .A(n4688), .B(\gpr[27][21] ), .Z(n1709) );
  ND2I U1941 ( .A(n4723), .B(\gpr[5][21] ), .Z(n1715) );
  ND2I U1942 ( .A(\gpr[13][21] ), .B(n2259), .Z(n1714) );
  ND2I U1943 ( .A(n4740), .B(\gpr[12][21] ), .Z(n1713) );
  ND2I U1944 ( .A(n1970), .B(\gpr[11][21] ), .Z(n1712) );
  ND4P U1945 ( .A(n1715), .B(n1714), .C(n1713), .D(n1712), .Z(n1716) );
  NR2I U1946 ( .A(n1716), .B(n248), .Z(n1740) );
  ND2I U1947 ( .A(\gpr[15][21] ), .B(n2172), .Z(n1720) );
  ND2I U1948 ( .A(n4746), .B(\gpr[6][21] ), .Z(n1719) );
  ND2I U1949 ( .A(n2061), .B(\gpr[7][21] ), .Z(n1718) );
  ND2I U1950 ( .A(n4748), .B(\gpr[14][21] ), .Z(n1717) );
  ND4 U1951 ( .A(n1720), .B(n1719), .C(n1718), .D(n1717), .Z(n1724) );
  ND2I U1952 ( .A(\gpr[1][21] ), .B(n4719), .Z(n1722) );
  ND2I U1953 ( .A(n2328), .B(\gpr[10][21] ), .Z(n1721) );
  ND2I U1954 ( .A(n1722), .B(n1721), .Z(n1723) );
  NR2I U1955 ( .A(n1724), .B(n1723), .Z(n1737) );
  ND2I U1956 ( .A(\gpr[9][21] ), .B(n2125), .Z(n1735) );
  ND2I U1957 ( .A(n1725), .B(\gpr[8][21] ), .Z(n1732) );
  ND2I U1958 ( .A(n4724), .B(\gpr[3][21] ), .Z(n1726) );
  AN2I U1959 ( .A(n498), .B(n1726), .Z(n1729) );
  ND2I U1960 ( .A(\gpr[2][21] ), .B(n1727), .Z(n1728) );
  ND2I U1961 ( .A(n1729), .B(n1728), .Z(n1730) );
  IVI U1962 ( .A(n1730), .Z(n1731) );
  ND2I U1963 ( .A(n1732), .B(n1731), .Z(n1733) );
  IVI U1964 ( .A(n1733), .Z(n1734) );
  AN2I U1965 ( .A(n1735), .B(n1734), .Z(n1736) );
  ND2I U1966 ( .A(n1737), .B(n1736), .Z(n1738) );
  IVI U1967 ( .A(n1738), .Z(n1739) );
  ND2I U1968 ( .A(n1740), .B(n1739), .Z(n1741) );
  ND2I U1969 ( .A(n249), .B(n1741), .Z(n1742) );
  IVI U1970 ( .A(n1742), .Z(rd_data1[21]) );
  NR2I U1971 ( .A(n1765), .B(n4854), .Z(n1745) );
  ND2I U1972 ( .A(n1583), .B(\gpr[16][11] ), .Z(n1743) );
  ND2I U1973 ( .A(n2094), .B(n1743), .Z(n1744) );
  NR2I U1974 ( .A(n1745), .B(n1744), .Z(n1759) );
  ND2I U1975 ( .A(\gpr[19][11] ), .B(n4703), .Z(n1747) );
  ND2I U1976 ( .A(\gpr[18][11] ), .B(n4726), .Z(n1746) );
  ND2I U1977 ( .A(n1747), .B(n1746), .Z(n1751) );
  ND2I U1978 ( .A(\gpr[20][11] ), .B(n2204), .Z(n1749) );
  ND2I U1979 ( .A(\gpr[23][11] ), .B(n2100), .Z(n1748) );
  ND2I U1980 ( .A(n1749), .B(n1748), .Z(n1750) );
  NR2I U1981 ( .A(n1751), .B(n1750), .Z(n1756) );
  ND2I U1982 ( .A(\gpr[17][11] ), .B(n2276), .Z(n1754) );
  ND2I U1983 ( .A(\gpr[21][11] ), .B(n2268), .Z(n1753) );
  AN2I U1984 ( .A(n1754), .B(n1753), .Z(n1755) );
  ND2I U1985 ( .A(n1756), .B(n1755), .Z(n1757) );
  IVI U1986 ( .A(n1757), .Z(n1758) );
  ND2I U1987 ( .A(n1759), .B(n1758), .Z(n1776) );
  ND2I U1988 ( .A(n2100), .B(\gpr[31][11] ), .Z(n1761) );
  ND2I U1989 ( .A(n4703), .B(\gpr[27][11] ), .Z(n1760) );
  AN2I U1990 ( .A(n1761), .B(n1760), .Z(n1764) );
  ND2I U1991 ( .A(\gpr[24][11] ), .B(n1762), .Z(n1763) );
  ND2I U1992 ( .A(n1764), .B(n1763), .Z(n1772) );
  NR2I U1993 ( .A(n1765), .B(n4855), .Z(n1768) );
  ND2I U1994 ( .A(n1383), .B(\gpr[25][11] ), .Z(n1766) );
  ND2I U1995 ( .A(n2079), .B(n1766), .Z(n1767) );
  NR2I U1996 ( .A(n1768), .B(n1767), .Z(n1770) );
  ND2I U1997 ( .A(n2204), .B(\gpr[28][11] ), .Z(n1769) );
  ND2I U1998 ( .A(n1770), .B(n1769), .Z(n1771) );
  NR2I U1999 ( .A(n1772), .B(n1771), .Z(n1773) );
  ND2I U2000 ( .A(n1774), .B(n1773), .Z(n1775) );
  AN2I U2001 ( .A(n1776), .B(n1775), .Z(n1808) );
  ND2I U2002 ( .A(n2129), .B(\gpr[8][11] ), .Z(n1778) );
  ND2I U2003 ( .A(\gpr[1][11] ), .B(n4719), .Z(n1777) );
  ND2I U2004 ( .A(n1778), .B(n1777), .Z(n1779) );
  ND2I U2005 ( .A(n4740), .B(\gpr[12][11] ), .Z(n1781) );
  ND2I U2006 ( .A(n1970), .B(\gpr[11][11] ), .Z(n1780) );
  ND2I U2007 ( .A(n1781), .B(n215), .Z(n1787) );
  ND2I U2008 ( .A(\gpr[13][11] ), .B(n2188), .Z(n1785) );
  ND2I U2009 ( .A(n2189), .B(\gpr[2][11] ), .Z(n1783) );
  ND2I U2010 ( .A(n2110), .B(\gpr[3][11] ), .Z(n1782) );
  AN2I U2011 ( .A(n1783), .B(n1782), .Z(n1784) );
  ND2I U2012 ( .A(n1785), .B(n1784), .Z(n1786) );
  NR2I U2013 ( .A(n1787), .B(n1786), .Z(n1789) );
  ND2I U2014 ( .A(\gpr[4][11] ), .B(n4732), .Z(n1788) );
  ND2I U2015 ( .A(n1789), .B(n1788), .Z(n1790) );
  NR2I U2016 ( .A(n1779), .B(n1790), .Z(n1806) );
  ND2I U2017 ( .A(n1791), .B(\gpr[7][11] ), .Z(n1793) );
  ND2I U2018 ( .A(n104), .B(\gpr[6][11] ), .Z(n1792) );
  ND2I U2019 ( .A(n1793), .B(n1792), .Z(n1794) );
  NR2I U2020 ( .A(n1794), .B(n280), .Z(n1795) );
  AN2I U2021 ( .A(n1796), .B(n1795), .Z(n1805) );
  ND2I U2022 ( .A(\gpr[10][11] ), .B(n101), .Z(n1802) );
  ND2I U2023 ( .A(n2157), .B(n296), .Z(n1799) );
  ND2I U2024 ( .A(\gpr[15][11] ), .B(n2172), .Z(n1798) );
  ND2I U2025 ( .A(n1799), .B(n1798), .Z(n1800) );
  IVI U2026 ( .A(n1800), .Z(n1801) );
  ND2I U2027 ( .A(n1802), .B(n1801), .Z(n1803) );
  IVI U2028 ( .A(n1803), .Z(n1804) );
  ND2I U2029 ( .A(n1806), .B(n250), .Z(n1807) );
  ND2I U2030 ( .A(n1808), .B(n1807), .Z(n1809) );
  IVI U2031 ( .A(n1809), .Z(rd_data1[11]) );
  ND2I U2032 ( .A(\gpr[28][19] ), .B(n2204), .Z(n1811) );
  ND2I U2033 ( .A(n1811), .B(n281), .Z(n1817) );
  ND2I U2034 ( .A(\gpr[31][19] ), .B(n4704), .Z(n1813) );
  ND2I U2035 ( .A(\gpr[27][19] ), .B(n4703), .Z(n1812) );
  AN2I U2036 ( .A(n1813), .B(n1812), .Z(n1815) );
  ND2I U2037 ( .A(\gpr[24][19] ), .B(n2233), .Z(n1814) );
  ND2I U2038 ( .A(n1815), .B(n1814), .Z(n1816) );
  NR2I U2039 ( .A(n1817), .B(n1816), .Z(n1820) );
  AO2 U2040 ( .A(n4702), .B(\gpr[26][19] ), .C(n2268), .D(\gpr[29][19] ), .Z(
        n1819) );
  ND2I U2041 ( .A(n2231), .B(\gpr[25][19] ), .Z(n1818) );
  ND2I U2042 ( .A(n1820), .B(n216), .Z(n1838) );
  NR2I U2043 ( .A(n2159), .B(n4867), .Z(n1823) );
  ND2I U2044 ( .A(n2155), .B(\gpr[16][19] ), .Z(n1821) );
  ND2I U2045 ( .A(n4709), .B(n1821), .Z(n1822) );
  NR2I U2046 ( .A(n1823), .B(n1822), .Z(n1836) );
  AO2 U2047 ( .A(n4702), .B(\gpr[18][19] ), .C(n1824), .D(\gpr[17][19] ), .Z(
        n1833) );
  ND2I U2048 ( .A(\gpr[20][19] ), .B(n2099), .Z(n1826) );
  ND2I U2049 ( .A(\gpr[21][19] ), .B(n2157), .Z(n1825) );
  AN2I U2050 ( .A(n1826), .B(n1825), .Z(n1830) );
  ND2I U2051 ( .A(\gpr[19][19] ), .B(n4703), .Z(n1828) );
  ND2I U2052 ( .A(n4704), .B(\gpr[23][19] ), .Z(n1827) );
  AN2I U2053 ( .A(n1828), .B(n1827), .Z(n1829) );
  ND2I U2054 ( .A(n1830), .B(n1829), .Z(n1831) );
  IVI U2055 ( .A(n1831), .Z(n1832) );
  ND2I U2056 ( .A(n1833), .B(n1832), .Z(n1834) );
  IVI U2057 ( .A(n1834), .Z(n1835) );
  ND2I U2058 ( .A(n1836), .B(n1835), .Z(n1837) );
  AN2I U2059 ( .A(n1838), .B(n1837), .Z(n1872) );
  ND2I U2060 ( .A(n2311), .B(\gpr[14][19] ), .Z(n1840) );
  ND2I U2061 ( .A(n4746), .B(\gpr[6][19] ), .Z(n1839) );
  ND2I U2062 ( .A(n1840), .B(n1839), .Z(n1843) );
  ND2I U2063 ( .A(n4723), .B(\gpr[5][19] ), .Z(n1841) );
  IVI U2064 ( .A(n1841), .Z(n1842) );
  NR2I U2065 ( .A(n1843), .B(n1842), .Z(n1857) );
  ND2I U2066 ( .A(\gpr[2][19] ), .B(n2189), .Z(n1845) );
  ND2I U2067 ( .A(\gpr[11][19] ), .B(n1970), .Z(n1844) );
  ND2I U2068 ( .A(\gpr[15][19] ), .B(n1846), .Z(n1850) );
  ND2I U2069 ( .A(n4747), .B(\gpr[7][19] ), .Z(n1847) );
  ND2I U2070 ( .A(n1847), .B(n498), .Z(n1848) );
  IVI U2071 ( .A(n1848), .Z(n1849) );
  AN2I U2072 ( .A(n1850), .B(n1849), .Z(n1851) );
  ND2I U2073 ( .A(n251), .B(n1851), .Z(n1852) );
  IVI U2074 ( .A(n1852), .Z(n1854) );
  ND2I U2075 ( .A(\gpr[4][19] ), .B(n2303), .Z(n1853) );
  ND2I U2076 ( .A(n1854), .B(n1853), .Z(n1855) );
  IVI U2077 ( .A(n1855), .Z(n1856) );
  ND2I U2078 ( .A(n1857), .B(n1856), .Z(n1858) );
  IVI U2079 ( .A(n1858), .Z(n1870) );
  ND2I U2080 ( .A(n2328), .B(\gpr[10][19] ), .Z(n1864) );
  ND2I U2081 ( .A(n4737), .B(\gpr[9][19] ), .Z(n1863) );
  ND2I U2082 ( .A(\gpr[13][19] ), .B(n2188), .Z(n1862) );
  ND2I U2083 ( .A(n4740), .B(\gpr[12][19] ), .Z(n1861) );
  ND2I U2084 ( .A(n1859), .B(\gpr[3][19] ), .Z(n1860) );
  ND4P U2085 ( .A(n1864), .B(n1863), .C(n1862), .D(n225), .Z(n1868) );
  ND2I U2086 ( .A(n2315), .B(\gpr[8][19] ), .Z(n1866) );
  ND2I U2087 ( .A(\gpr[1][19] ), .B(n4719), .Z(n1865) );
  ND2I U2088 ( .A(n1866), .B(n1865), .Z(n1867) );
  NR2I U2089 ( .A(n1868), .B(n1867), .Z(n1869) );
  ND2I U2090 ( .A(n1870), .B(n1869), .Z(n1871) );
  AN2I U2091 ( .A(n1872), .B(n1871), .Z(rd_data1[19]) );
  NR2I U2092 ( .A(n2297), .B(n4858), .Z(n1875) );
  ND2I U2093 ( .A(n1360), .B(\gpr[17][13] ), .Z(n1873) );
  ND2I U2094 ( .A(n4709), .B(n1873), .Z(n1874) );
  NR2I U2095 ( .A(n1875), .B(n1874), .Z(n1887) );
  AO2 U2096 ( .A(n4702), .B(\gpr[18][13] ), .C(n2233), .D(\gpr[16][13] ), .Z(
        n1884) );
  ND2I U2097 ( .A(\gpr[20][13] ), .B(n2099), .Z(n1877) );
  ND2I U2098 ( .A(\gpr[22][13] ), .B(n207), .Z(n1876) );
  AN2I U2099 ( .A(n1877), .B(n1876), .Z(n1881) );
  ND2I U2100 ( .A(\gpr[19][13] ), .B(n4703), .Z(n1879) );
  ND2I U2101 ( .A(\gpr[21][13] ), .B(n2268), .Z(n1878) );
  AN2I U2102 ( .A(n1879), .B(n1878), .Z(n1880) );
  ND2I U2103 ( .A(n1881), .B(n1880), .Z(n1882) );
  IVI U2104 ( .A(n1882), .Z(n1883) );
  ND2I U2105 ( .A(n1884), .B(n1883), .Z(n1885) );
  IVI U2106 ( .A(n1885), .Z(n1886) );
  ND2I U2107 ( .A(n1887), .B(n1886), .Z(n1904) );
  ND2I U2108 ( .A(n4726), .B(\gpr[26][13] ), .Z(n1888) );
  IVI U2109 ( .A(n1888), .Z(n1892) );
  ND2I U2110 ( .A(\gpr[24][13] ), .B(n1205), .Z(n1890) );
  ND2I U2111 ( .A(n283), .B(n1890), .Z(n1891) );
  NR2I U2112 ( .A(n1892), .B(n1891), .Z(n1900) );
  ND2I U2113 ( .A(\gpr[29][13] ), .B(n4701), .Z(n1894) );
  ND2I U2114 ( .A(n4703), .B(\gpr[27][13] ), .Z(n1893) );
  ND2I U2115 ( .A(n1894), .B(n1893), .Z(n1898) );
  ND2I U2116 ( .A(\gpr[31][13] ), .B(n2100), .Z(n1896) );
  ND2I U2117 ( .A(\gpr[28][13] ), .B(n2099), .Z(n1895) );
  ND2I U2118 ( .A(n1896), .B(n1895), .Z(n1897) );
  NR2I U2119 ( .A(n1898), .B(n1897), .Z(n1899) );
  AN2I U2120 ( .A(n1900), .B(n1899), .Z(n1902) );
  ND2I U2121 ( .A(\gpr[25][13] ), .B(n206), .Z(n1901) );
  ND2I U2122 ( .A(n1902), .B(n284), .Z(n1903) );
  AN2I U2123 ( .A(n1904), .B(n1903), .Z(n1937) );
  ND2I U2124 ( .A(n4740), .B(\gpr[12][13] ), .Z(n1906) );
  ND2I U2125 ( .A(n2255), .B(\gpr[11][13] ), .Z(n1905) );
  ND2I U2126 ( .A(n1906), .B(n285), .Z(n1912) );
  ND2I U2127 ( .A(\gpr[13][13] ), .B(n2188), .Z(n1910) );
  ND2I U2128 ( .A(n2189), .B(\gpr[2][13] ), .Z(n1908) );
  ND2I U2129 ( .A(n2110), .B(\gpr[3][13] ), .Z(n1907) );
  AN2I U2130 ( .A(n1908), .B(n1907), .Z(n1909) );
  ND2I U2131 ( .A(n1910), .B(n1909), .Z(n1911) );
  NR2I U2132 ( .A(n1912), .B(n1911), .Z(n1920) );
  ND2I U2133 ( .A(n2125), .B(\gpr[9][13] ), .Z(n1918) );
  ND2I U2134 ( .A(n104), .B(\gpr[6][13] ), .Z(n1914) );
  ND2I U2135 ( .A(n2306), .B(\gpr[7][13] ), .Z(n1913) );
  AO3P U2136 ( .A(n1915), .B(n5216), .C(n1914), .D(n1913), .Z(n1916) );
  IVI U2137 ( .A(n1916), .Z(n1917) );
  AN2I U2138 ( .A(n1918), .B(n1917), .Z(n1919) );
  ND2I U2139 ( .A(n1920), .B(n1919), .Z(n1921) );
  IVI U2140 ( .A(n1921), .Z(n1935) );
  ND2I U2141 ( .A(\gpr[15][13] ), .B(n4745), .Z(n1923) );
  ND2I U2142 ( .A(\gpr[5][13] ), .B(n4723), .Z(n1922) );
  ND2I U2143 ( .A(n1923), .B(n1922), .Z(n1924) );
  IVI U2144 ( .A(n1924), .Z(n1926) );
  ND2I U2145 ( .A(\gpr[14][13] ), .B(n1990), .Z(n1925) );
  ND2I U2146 ( .A(n1926), .B(n1925), .Z(n1933) );
  ND2I U2147 ( .A(n4732), .B(\gpr[4][13] ), .Z(n1931) );
  ND2I U2148 ( .A(n1307), .B(\gpr[8][13] ), .Z(n1928) );
  ND2I U2149 ( .A(\gpr[1][13] ), .B(n4719), .Z(n1927) );
  ND2I U2150 ( .A(n1928), .B(n1927), .Z(n1929) );
  IVI U2151 ( .A(n1929), .Z(n1930) );
  ND2I U2152 ( .A(n1931), .B(n1930), .Z(n1932) );
  NR2I U2153 ( .A(n1933), .B(n1932), .Z(n1934) );
  ND2I U2154 ( .A(n1935), .B(n1934), .Z(n1936) );
  AN2I U2155 ( .A(n1937), .B(n1936), .Z(rd_data1[13]) );
  AO2 U2156 ( .A(n4726), .B(\gpr[26][9] ), .C(n1938), .D(\gpr[25][9] ), .Z(
        n1948) );
  ND2I U2157 ( .A(\gpr[28][9] ), .B(n2204), .Z(n1940) );
  ND2I U2158 ( .A(\gpr[31][9] ), .B(n2100), .Z(n1939) );
  ND2I U2159 ( .A(n1940), .B(n1939), .Z(n1946) );
  ND2I U2160 ( .A(\gpr[27][9] ), .B(n2284), .Z(n1944) );
  ND2I U2161 ( .A(\gpr[29][9] ), .B(n2268), .Z(n1941) );
  ND2I U2162 ( .A(n1941), .B(n286), .Z(n1942) );
  IVI U2163 ( .A(n1942), .Z(n1943) );
  ND2I U2164 ( .A(n1944), .B(n1943), .Z(n1945) );
  NR2I U2165 ( .A(n1946), .B(n1945), .Z(n1947) );
  ND2I U2166 ( .A(n1948), .B(n1947), .Z(n1949) );
  IVI U2167 ( .A(n1949), .Z(n1951) );
  ND2I U2168 ( .A(n2147), .B(\gpr[24][9] ), .Z(n1950) );
  ND2I U2169 ( .A(n1951), .B(n287), .Z(n1968) );
  AO2 U2170 ( .A(n4701), .B(\gpr[21][9] ), .C(n1952), .D(\gpr[17][9] ), .Z(
        n1966) );
  NR2I U2171 ( .A(n1889), .B(n4852), .Z(n1955) );
  ND2I U2172 ( .A(n4686), .B(\gpr[16][9] ), .Z(n1953) );
  ND2I U2173 ( .A(n2094), .B(n1953), .Z(n1954) );
  NR2I U2174 ( .A(n1955), .B(n1954), .Z(n1963) );
  ND2I U2175 ( .A(n4703), .B(\gpr[19][9] ), .Z(n1957) );
  ND2I U2176 ( .A(\gpr[18][9] ), .B(n4726), .Z(n1956) );
  ND2I U2177 ( .A(n1957), .B(n1956), .Z(n1961) );
  ND2I U2178 ( .A(n2158), .B(\gpr[20][9] ), .Z(n1959) );
  ND2I U2179 ( .A(n2100), .B(\gpr[23][9] ), .Z(n1958) );
  ND2I U2180 ( .A(n1959), .B(n1958), .Z(n1960) );
  NR2I U2181 ( .A(n1961), .B(n1960), .Z(n1962) );
  ND2I U2182 ( .A(n1963), .B(n1962), .Z(n1964) );
  IVI U2183 ( .A(n1964), .Z(n1965) );
  ND2I U2184 ( .A(n1966), .B(n1965), .Z(n1967) );
  ND2I U2185 ( .A(n1968), .B(n1967), .Z(n1969) );
  IVI U2186 ( .A(n1969), .Z(n2003) );
  ND2I U2187 ( .A(\gpr[9][9] ), .B(n4737), .Z(n1975) );
  ND2I U2188 ( .A(n106), .B(\gpr[12][9] ), .Z(n1972) );
  ND2I U2189 ( .A(n1970), .B(\gpr[11][9] ), .Z(n1971) );
  ND2I U2190 ( .A(n1972), .B(n217), .Z(n1973) );
  IVI U2191 ( .A(n1973), .Z(n1974) );
  ND2I U2192 ( .A(n1975), .B(n1974), .Z(n1976) );
  NR2I U2193 ( .A(n252), .B(n1976), .Z(n1982) );
  IVI U2194 ( .A(n1977), .Z(n2129) );
  ND2I U2195 ( .A(n2129), .B(\gpr[8][9] ), .Z(n1979) );
  ND2I U2196 ( .A(\gpr[1][9] ), .B(n4719), .Z(n1978) );
  ND2I U2197 ( .A(n1979), .B(n1978), .Z(n1980) );
  IVI U2198 ( .A(n1980), .Z(n1981) );
  AN2I U2199 ( .A(n1982), .B(n1981), .Z(n2001) );
  ND2I U2200 ( .A(n1797), .B(\gpr[10][9] ), .Z(n1984) );
  ND2I U2201 ( .A(\gpr[13][9] ), .B(n4718), .Z(n1988) );
  ND2I U2202 ( .A(n2115), .B(\gpr[2][9] ), .Z(n1986) );
  ND2I U2203 ( .A(n2110), .B(\gpr[3][9] ), .Z(n1985) );
  AN2I U2204 ( .A(n1986), .B(n1985), .Z(n1987) );
  AN2I U2205 ( .A(n1988), .B(n1987), .Z(n1989) );
  ND2I U2206 ( .A(n1984), .B(n1989), .Z(n1999) );
  ND2I U2207 ( .A(\gpr[4][9] ), .B(n2303), .Z(n1997) );
  ND2I U2208 ( .A(n105), .B(\gpr[6][9] ), .Z(n1994) );
  ND2I U2209 ( .A(\gpr[15][9] ), .B(n4745), .Z(n1993) );
  ND2I U2210 ( .A(n2114), .B(\gpr[7][9] ), .Z(n1992) );
  ND2I U2211 ( .A(n1990), .B(\gpr[14][9] ), .Z(n1991) );
  ND4P U2212 ( .A(n1994), .B(n1993), .C(n1992), .D(n1991), .Z(n1995) );
  IVI U2213 ( .A(n1995), .Z(n1996) );
  ND2I U2214 ( .A(n1997), .B(n1996), .Z(n1998) );
  NR2I U2215 ( .A(n1999), .B(n1998), .Z(n2000) );
  ND2I U2216 ( .A(n2001), .B(n2000), .Z(n2002) );
  AN2I U2217 ( .A(n2003), .B(n2002), .Z(rd_data1[9]) );
  AO2 U2218 ( .A(n2004), .B(\gpr[24][1] ), .C(n2146), .D(\gpr[25][1] ), .Z(
        n2016) );
  ND2I U2219 ( .A(n2020), .B(\gpr[30][1] ), .Z(n2005) );
  AO3 U2220 ( .A(n2006), .B(n4827), .C(n2079), .D(n2005), .Z(n2007) );
  IVI U2221 ( .A(n2007), .Z(n2015) );
  ND2I U2222 ( .A(\gpr[31][1] ), .B(n2100), .Z(n2008) );
  IVI U2223 ( .A(n2008), .Z(n2012) );
  ND2I U2224 ( .A(\gpr[26][1] ), .B(n2077), .Z(n2010) );
  ND2I U2225 ( .A(n2216), .B(\gpr[27][1] ), .Z(n2009) );
  ND2I U2226 ( .A(n2010), .B(n2009), .Z(n2011) );
  NR2I U2227 ( .A(n2012), .B(n2011), .Z(n2014) );
  ND2I U2228 ( .A(\gpr[28][1] ), .B(n2158), .Z(n2013) );
  ND4P U2229 ( .A(n2016), .B(n2015), .C(n2014), .D(n2013), .Z(n2035) );
  ND2I U2230 ( .A(\gpr[16][1] ), .B(n2017), .Z(n2019) );
  ND2I U2231 ( .A(\gpr[18][1] ), .B(n2077), .Z(n2018) );
  AN2I U2232 ( .A(n2019), .B(n2018), .Z(n2033) );
  ND2I U2233 ( .A(n2020), .B(\gpr[22][1] ), .Z(n2021) );
  IVI U2234 ( .A(n2023), .Z(n2031) );
  ND2I U2235 ( .A(n2216), .B(\gpr[19][1] ), .Z(n2025) );
  ND2I U2236 ( .A(\gpr[17][1] ), .B(n2047), .Z(n2024) );
  ND2I U2237 ( .A(n2025), .B(n2024), .Z(n2029) );
  ND2I U2238 ( .A(\gpr[20][1] ), .B(n2158), .Z(n2027) );
  ND2I U2239 ( .A(n2100), .B(\gpr[23][1] ), .Z(n2026) );
  ND2I U2240 ( .A(n2027), .B(n2026), .Z(n2028) );
  NR2I U2241 ( .A(n2029), .B(n2028), .Z(n2030) );
  AN2I U2242 ( .A(n2031), .B(n2030), .Z(n2032) );
  ND2I U2243 ( .A(n2033), .B(n2032), .Z(n2034) );
  ND2I U2244 ( .A(n2035), .B(n2034), .Z(n2036) );
  IVI U2245 ( .A(n2036), .Z(n2076) );
  ND2I U2246 ( .A(\gpr[1][1] ), .B(n4719), .Z(n2046) );
  ND2I U2247 ( .A(\gpr[2][1] ), .B(n1246), .Z(n2038) );
  ND2I U2248 ( .A(n2039), .B(n2038), .Z(n2044) );
  ND2I U2249 ( .A(\gpr[3][1] ), .B(n2040), .Z(n2042) );
  ND2I U2250 ( .A(\gpr[15][1] ), .B(n2172), .Z(n2041) );
  ND2I U2251 ( .A(n2042), .B(n2041), .Z(n2043) );
  NR2I U2252 ( .A(n2044), .B(n2043), .Z(n2045) );
  AN2I U2253 ( .A(n2046), .B(n2045), .Z(n2074) );
  AO2 U2254 ( .A(n4726), .B(\gpr[10][1] ), .C(n2047), .D(\gpr[9][1] ), .Z(
        n2056) );
  ND2I U2255 ( .A(\gpr[8][1] ), .B(n2048), .Z(n2049) );
  AO7 U2256 ( .A(n2050), .B(n4760), .C(n2049), .Z(n2054) );
  ND2I U2257 ( .A(n4694), .B(\gpr[12][1] ), .Z(n2052) );
  ND2I U2258 ( .A(n4688), .B(\gpr[11][1] ), .Z(n2051) );
  ND2I U2259 ( .A(n2052), .B(n2051), .Z(n2053) );
  NR2I U2260 ( .A(n2054), .B(n2053), .Z(n2055) );
  ND2I U2261 ( .A(n2056), .B(n2055), .Z(n2057) );
  ND2I U2262 ( .A(n2307), .B(n2057), .Z(n2071) );
  ND2I U2263 ( .A(\gpr[4][1] ), .B(n2303), .Z(n2068) );
  ND2I U2264 ( .A(n2058), .B(\gpr[13][1] ), .Z(n2059) );
  ND2I U2265 ( .A(n2174), .B(n2059), .Z(n2060) );
  IVI U2266 ( .A(n2060), .Z(n2065) );
  ND2I U2267 ( .A(\gpr[7][1] ), .B(n2061), .Z(n2063) );
  ND2I U2268 ( .A(\gpr[6][1] ), .B(n105), .Z(n2062) );
  AN2I U2269 ( .A(n2063), .B(n2062), .Z(n2064) );
  ND2I U2270 ( .A(n2065), .B(n2064), .Z(n2066) );
  IVI U2271 ( .A(n2066), .Z(n2067) );
  ND2I U2272 ( .A(n2068), .B(n2067), .Z(n2069) );
  IVI U2273 ( .A(n2069), .Z(n2070) );
  ND2I U2274 ( .A(n2071), .B(n2070), .Z(n2072) );
  IVI U2275 ( .A(n2072), .Z(n2073) );
  ND2I U2276 ( .A(n2074), .B(n2073), .Z(n2075) );
  AN2I U2277 ( .A(n2076), .B(n2075), .Z(rd_data1[1]) );
  AO2 U2278 ( .A(n2077), .B(\gpr[26][3] ), .C(n1647), .D(\gpr[25][3] ), .Z(
        n2089) );
  NR2I U2279 ( .A(n2092), .B(n4843), .Z(n2081) );
  ND2I U2280 ( .A(n2296), .B(\gpr[24][3] ), .Z(n2078) );
  ND2I U2281 ( .A(n2079), .B(n2078), .Z(n2080) );
  NR2I U2282 ( .A(n2081), .B(n2080), .Z(n2082) );
  IVI U2283 ( .A(n2082), .Z(n2088) );
  ND2I U2284 ( .A(\gpr[28][3] ), .B(n4694), .Z(n2086) );
  ND2I U2285 ( .A(\gpr[31][3] ), .B(n2100), .Z(n2085) );
  ND2I U2286 ( .A(\gpr[27][3] ), .B(n2216), .Z(n2084) );
  ND2I U2287 ( .A(\gpr[29][3] ), .B(n2292), .Z(n2083) );
  ND2I U2288 ( .A(\gpr[17][3] ), .B(n1383), .Z(n2091) );
  ND2I U2289 ( .A(\gpr[16][3] ), .B(n1583), .Z(n2090) );
  AN2I U2290 ( .A(n2091), .B(n2090), .Z(n2107) );
  NR2I U2291 ( .A(n2092), .B(n4764), .Z(n2096) );
  ND2I U2292 ( .A(n2077), .B(\gpr[18][3] ), .Z(n2093) );
  ND2I U2293 ( .A(n2094), .B(n2093), .Z(n2095) );
  NR2I U2294 ( .A(n2096), .B(n2095), .Z(n2106) );
  ND2I U2295 ( .A(n2216), .B(\gpr[19][3] ), .Z(n2098) );
  ND2I U2296 ( .A(n2292), .B(\gpr[21][3] ), .Z(n2097) );
  ND2I U2297 ( .A(n2098), .B(n2097), .Z(n2104) );
  ND2I U2298 ( .A(\gpr[20][3] ), .B(n2099), .Z(n2102) );
  ND2I U2299 ( .A(n2100), .B(\gpr[23][3] ), .Z(n2101) );
  ND2I U2300 ( .A(n2102), .B(n2101), .Z(n2103) );
  NR2I U2301 ( .A(n2104), .B(n2103), .Z(n2105) );
  ND2I U2302 ( .A(\gpr[1][3] ), .B(n4719), .Z(n2124) );
  B3IP U2303 ( .A(n2108), .Z1(n2109), .Z2(n2303) );
  OR2I U2304 ( .A(n2109), .B(n4967), .Z(n2123) );
  ND2I U2305 ( .A(\gpr[13][3] ), .B(n2188), .Z(n2112) );
  ND2I U2306 ( .A(n2110), .B(\gpr[3][3] ), .Z(n2111) );
  ND2I U2307 ( .A(n2112), .B(n2111), .Z(n2113) );
  IVI U2308 ( .A(n2113), .Z(n2122) );
  ND2I U2309 ( .A(n105), .B(\gpr[6][3] ), .Z(n2119) );
  ND2I U2310 ( .A(n2114), .B(\gpr[7][3] ), .Z(n2117) );
  ND2I U2311 ( .A(n2115), .B(\gpr[2][3] ), .Z(n2116) );
  AN2I U2312 ( .A(n2117), .B(n2116), .Z(n2118) );
  ND2I U2313 ( .A(n2119), .B(n2118), .Z(n2120) );
  IVI U2314 ( .A(n2120), .Z(n2121) );
  ND2I U2315 ( .A(n2125), .B(\gpr[9][3] ), .Z(n2128) );
  ND2I U2316 ( .A(n2126), .B(\gpr[14][3] ), .Z(n2127) );
  ND2I U2317 ( .A(n2128), .B(n2127), .Z(n2140) );
  ND2I U2318 ( .A(n2129), .B(\gpr[8][3] ), .Z(n2131) );
  ND2I U2319 ( .A(n1797), .B(\gpr[10][3] ), .Z(n2130) );
  ND2I U2320 ( .A(\gpr[5][3] ), .B(n4723), .Z(n2138) );
  ND2I U2321 ( .A(n2132), .B(\gpr[12][3] ), .Z(n2135) );
  ND2I U2322 ( .A(n2133), .B(\gpr[11][3] ), .Z(n2134) );
  ND2I U2323 ( .A(n2135), .B(n218), .Z(n2136) );
  NR2I U2324 ( .A(n253), .B(n2136), .Z(n2137) );
  AN2I U2325 ( .A(n2138), .B(n2137), .Z(n2139) );
  ND2I U2326 ( .A(\gpr[20][17] ), .B(n2204), .Z(n2145) );
  ND2I U2327 ( .A(\gpr[21][17] ), .B(n2268), .Z(n2142) );
  ND2I U2328 ( .A(\gpr[23][17] ), .B(n4704), .Z(n2141) );
  ND2I U2329 ( .A(n2142), .B(n2141), .Z(n2143) );
  NR2I U2330 ( .A(n288), .B(n2143), .Z(n2144) );
  AN2I U2331 ( .A(n2145), .B(n2144), .Z(n2153) );
  AO2 U2332 ( .A(n4702), .B(\gpr[18][17] ), .C(n2146), .D(\gpr[17][17] ), .Z(
        n2152) );
  NR2I U2333 ( .A(n2159), .B(n4863), .Z(n2150) );
  ND2I U2334 ( .A(n2147), .B(\gpr[16][17] ), .Z(n2148) );
  ND2I U2335 ( .A(n4709), .B(n2148), .Z(n2149) );
  NR2I U2336 ( .A(n2150), .B(n2149), .Z(n2151) );
  ND2I U2337 ( .A(n2153), .B(n255), .Z(n2169) );
  ND2I U2338 ( .A(n4688), .B(\gpr[27][17] ), .Z(n2154) );
  AO2 U2339 ( .A(n2155), .B(\gpr[24][17] ), .C(n2231), .D(\gpr[25][17] ), .Z(
        n2156) );
  AN2I U2340 ( .A(n289), .B(n2156), .Z(n2167) );
  AO2 U2341 ( .A(n4702), .B(\gpr[26][17] ), .C(n2157), .D(\gpr[29][17] ), .Z(
        n2166) );
  ND2I U2342 ( .A(\gpr[28][17] ), .B(n2158), .Z(n2163) );
  ND2I U2343 ( .A(\gpr[31][17] ), .B(n4704), .Z(n2160) );
  ND2I U2344 ( .A(n290), .B(n2160), .Z(n2161) );
  IVI U2345 ( .A(n2161), .Z(n2162) );
  ND2I U2346 ( .A(n2163), .B(n2162), .Z(n2164) );
  IVI U2347 ( .A(n2164), .Z(n2165) );
  ND2I U2348 ( .A(n2167), .B(n256), .Z(n2168) );
  AN2I U2349 ( .A(n2169), .B(n2168), .Z(n2203) );
  ND2I U2350 ( .A(n2311), .B(\gpr[14][17] ), .Z(n2171) );
  ND2I U2351 ( .A(n4746), .B(\gpr[6][17] ), .Z(n2170) );
  ND2I U2352 ( .A(n2171), .B(n2170), .Z(n2187) );
  ND2I U2353 ( .A(n4732), .B(\gpr[4][17] ), .Z(n2185) );
  ND2I U2354 ( .A(n4723), .B(\gpr[5][17] ), .Z(n2182) );
  ND2I U2355 ( .A(\gpr[15][17] ), .B(n2172), .Z(n2180) );
  IVI U2356 ( .A(n2173), .Z(n2247) );
  ND2I U2357 ( .A(n2247), .B(\gpr[7][17] ), .Z(n2175) );
  AN2I U2358 ( .A(n2175), .B(n2174), .Z(n2177) );
  ND2I U2359 ( .A(n909), .B(\gpr[3][17] ), .Z(n2176) );
  ND2I U2360 ( .A(n2177), .B(n2176), .Z(n2178) );
  IVI U2361 ( .A(n2178), .Z(n2179) );
  AN2I U2362 ( .A(n2180), .B(n2179), .Z(n2181) );
  ND2I U2363 ( .A(n2182), .B(n2181), .Z(n2183) );
  IVI U2364 ( .A(n2183), .Z(n2184) );
  ND2I U2365 ( .A(n2185), .B(n2184), .Z(n2186) );
  NR2I U2366 ( .A(n2187), .B(n2186), .Z(n2201) );
  ND2I U2367 ( .A(n2328), .B(\gpr[10][17] ), .Z(n2196) );
  ND2I U2368 ( .A(n4737), .B(\gpr[9][17] ), .Z(n2195) );
  ND2I U2369 ( .A(\gpr[13][17] ), .B(n2188), .Z(n2194) );
  ND2I U2370 ( .A(n2317), .B(\gpr[12][17] ), .Z(n2193) );
  ND2I U2371 ( .A(n2255), .B(\gpr[11][17] ), .Z(n2191) );
  ND2I U2372 ( .A(n1618), .B(\gpr[2][17] ), .Z(n2190) );
  AN2I U2373 ( .A(n2191), .B(n2190), .Z(n2192) );
  ND2I U2374 ( .A(n2197), .B(\gpr[8][17] ), .Z(n2199) );
  ND2I U2375 ( .A(\gpr[1][17] ), .B(n4719), .Z(n2198) );
  ND2I U2376 ( .A(n2201), .B(n2200), .Z(n2202) );
  AN2I U2377 ( .A(n2203), .B(n2202), .Z(rd_data1[17]) );
  ND2I U2378 ( .A(\gpr[20][29] ), .B(n2158), .Z(n2206) );
  ND2I U2379 ( .A(\gpr[16][29] ), .B(n1598), .Z(n2205) );
  ND2I U2380 ( .A(n2206), .B(n2205), .Z(n2211) );
  ND2I U2381 ( .A(\gpr[21][29] ), .B(n2292), .Z(n2209) );
  ND2I U2382 ( .A(\gpr[18][29] ), .B(n2207), .Z(n2208) );
  ND2I U2383 ( .A(n2209), .B(n2208), .Z(n2210) );
  NR2I U2384 ( .A(n2211), .B(n2210), .Z(n2223) );
  NR2I U2385 ( .A(n1765), .B(n4880), .Z(n2214) );
  ND2I U2386 ( .A(n2047), .B(\gpr[17][29] ), .Z(n2212) );
  ND2I U2387 ( .A(n4709), .B(n2212), .Z(n2213) );
  NR2I U2388 ( .A(n2214), .B(n2213), .Z(n2221) );
  ND2I U2389 ( .A(\gpr[23][29] ), .B(n2215), .Z(n2218) );
  ND2I U2390 ( .A(\gpr[19][29] ), .B(n2216), .Z(n2217) );
  ND2I U2391 ( .A(n2218), .B(n2217), .Z(n2219) );
  IVI U2392 ( .A(n2219), .Z(n2220) );
  AN2I U2393 ( .A(n2221), .B(n2220), .Z(n2222) );
  ND2I U2394 ( .A(n2223), .B(n2222), .Z(n2238) );
  ND2I U2395 ( .A(\gpr[28][29] ), .B(n2158), .Z(n2230) );
  ND2I U2396 ( .A(\gpr[27][29] ), .B(n4688), .Z(n2224) );
  ND2I U2397 ( .A(n291), .B(n2224), .Z(n2228) );
  ND2I U2398 ( .A(\gpr[31][29] ), .B(n2215), .Z(n2226) );
  ND2I U2399 ( .A(\gpr[29][29] ), .B(n4701), .Z(n2225) );
  ND2I U2400 ( .A(n2226), .B(n2225), .Z(n2227) );
  NR2I U2401 ( .A(n2228), .B(n2227), .Z(n2229) );
  ND2I U2402 ( .A(n2231), .B(\gpr[25][29] ), .Z(n2232) );
  ND2I U2403 ( .A(n4690), .B(n2232), .Z(n2235) );
  NR2I U2404 ( .A(n2235), .B(n2234), .Z(n2236) );
  ND2I U2405 ( .A(n257), .B(n2236), .Z(n2237) );
  AN2I U2406 ( .A(n2238), .B(n2237), .Z(n2267) );
  ND2I U2407 ( .A(n2317), .B(\gpr[12][29] ), .Z(n2243) );
  ND2I U2408 ( .A(n4723), .B(\gpr[5][29] ), .Z(n2242) );
  IVI U2409 ( .A(n2239), .Z(n2315) );
  ND2I U2410 ( .A(n2315), .B(\gpr[8][29] ), .Z(n2241) );
  ND2I U2411 ( .A(\gpr[9][29] ), .B(n4737), .Z(n2240) );
  ND4P U2412 ( .A(n2243), .B(n2242), .C(n2241), .D(n2240), .Z(n2244) );
  NR2I U2413 ( .A(n258), .B(n2244), .Z(n2265) );
  ND2I U2414 ( .A(\gpr[1][29] ), .B(n4719), .Z(n2246) );
  ND2I U2415 ( .A(n1797), .B(\gpr[10][29] ), .Z(n2245) );
  ND2I U2416 ( .A(n2246), .B(n2245), .Z(n2263) );
  ND2I U2417 ( .A(n1089), .B(\gpr[3][29] ), .Z(n2250) );
  ND2I U2418 ( .A(n2247), .B(\gpr[7][29] ), .Z(n2248) );
  AN2I U2419 ( .A(n2248), .B(n498), .Z(n2249) );
  ND2I U2420 ( .A(n2250), .B(n2249), .Z(n2251) );
  NR2I U2421 ( .A(n292), .B(n2251), .Z(n2262) );
  ND2I U2422 ( .A(n2252), .B(\gpr[14][29] ), .Z(n2254) );
  ND2I U2423 ( .A(n4746), .B(\gpr[6][29] ), .Z(n2253) );
  ND2I U2424 ( .A(n2254), .B(n2253), .Z(n2261) );
  ND2I U2425 ( .A(n2255), .B(\gpr[11][29] ), .Z(n2258) );
  ND2I U2426 ( .A(n2256), .B(\gpr[2][29] ), .Z(n2257) );
  ND2I U2427 ( .A(\gpr[13][29] ), .B(n2259), .Z(n2260) );
  ND2I U2428 ( .A(n2265), .B(n2264), .Z(n2266) );
  AN2I U2429 ( .A(n2267), .B(n2266), .Z(rd_data1[29]) );
  ND2I U2430 ( .A(\gpr[28][28] ), .B(n4694), .Z(n2270) );
  ND2I U2431 ( .A(n2268), .B(\gpr[29][28] ), .Z(n2269) );
  ND2I U2432 ( .A(n2270), .B(n2269), .Z(n2274) );
  ND2I U2433 ( .A(\gpr[24][28] ), .B(n2271), .Z(n2272) );
  ND2I U2434 ( .A(n4690), .B(n2272), .Z(n2273) );
  NR2I U2435 ( .A(n2274), .B(n2273), .Z(n2288) );
  ND2I U2436 ( .A(\gpr[31][28] ), .B(n4704), .Z(n2281) );
  ND2I U2437 ( .A(\gpr[25][28] ), .B(n2276), .Z(n2278) );
  ND2I U2438 ( .A(n4702), .B(\gpr[26][28] ), .Z(n2277) );
  ND2I U2439 ( .A(n2278), .B(n2277), .Z(n2279) );
  IVI U2440 ( .A(n2279), .Z(n2280) );
  ND2I U2441 ( .A(n2281), .B(n2280), .Z(n2282) );
  IVI U2442 ( .A(n2282), .Z(n2287) );
  NR2I U2443 ( .A(n4707), .B(n4878), .Z(n2283) );
  IVI U2444 ( .A(n2283), .Z(n2286) );
  ND2I U2445 ( .A(n2284), .B(\gpr[27][28] ), .Z(n2285) );
  ND2I U2446 ( .A(\gpr[22][28] ), .B(n207), .Z(n2290) );
  ND2I U2447 ( .A(\gpr[19][28] ), .B(n4688), .Z(n2289) );
  ND2I U2448 ( .A(n2290), .B(n2289), .Z(n2295) );
  ND2I U2449 ( .A(\gpr[20][28] ), .B(n2291), .Z(n2294) );
  ND2I U2450 ( .A(\gpr[21][28] ), .B(n2292), .Z(n2293) );
  NR2I U2451 ( .A(n2297), .B(n4879), .Z(n2300) );
  ND2I U2452 ( .A(n206), .B(\gpr[17][28] ), .Z(n2298) );
  ND2I U2453 ( .A(n4709), .B(n2298), .Z(n2299) );
  NR2I U2454 ( .A(n2300), .B(n2299), .Z(n2301) );
  IVI U2455 ( .A(n2302), .Z(n2338) );
  ND2I U2456 ( .A(\gpr[6][28] ), .B(n4746), .Z(n2305) );
  ND2I U2457 ( .A(n4723), .B(\gpr[5][28] ), .Z(n2304) );
  ND2I U2458 ( .A(n2306), .B(\gpr[7][28] ), .Z(n2310) );
  AN2I U2459 ( .A(n2307), .B(\gpr[13][28] ), .Z(n2308) );
  ND2I U2460 ( .A(n4701), .B(n2308), .Z(n2309) );
  ND2I U2461 ( .A(n2311), .B(\gpr[14][28] ), .Z(n2314) );
  ND2I U2462 ( .A(n2312), .B(\gpr[15][28] ), .Z(n2313) );
  ND2I U2463 ( .A(\gpr[8][28] ), .B(n2315), .Z(n2316) );
  ND2I U2464 ( .A(n106), .B(\gpr[12][28] ), .Z(n2327) );
  ND2I U2465 ( .A(n4739), .B(\gpr[11][28] ), .Z(n2319) );
  ND2I U2466 ( .A(n1859), .B(\gpr[3][28] ), .Z(n2318) );
  ND2I U2467 ( .A(n2319), .B(n2318), .Z(n2325) );
  ND2I U2468 ( .A(\gpr[1][28] ), .B(n2320), .Z(n2323) );
  AN2I U2469 ( .A(n2321), .B(n498), .Z(n2322) );
  ND2I U2470 ( .A(n2323), .B(n2322), .Z(n2324) );
  NR2I U2471 ( .A(n2325), .B(n2324), .Z(n2326) );
  AN2I U2472 ( .A(n2327), .B(n2326), .Z(n2333) );
  ND2I U2473 ( .A(n4737), .B(\gpr[9][28] ), .Z(n2330) );
  ND2I U2474 ( .A(n101), .B(\gpr[10][28] ), .Z(n2329) );
  ND2I U2475 ( .A(n2330), .B(n2329), .Z(n2331) );
  IVI U2476 ( .A(n2331), .Z(n2332) );
  ND2I U2477 ( .A(n2333), .B(n2332), .Z(n2334) );
  IVI U2478 ( .A(n2334), .Z(n2335) );
  ND2I U2479 ( .A(n2336), .B(n2335), .Z(n2337) );
  AN2I U2480 ( .A(n2338), .B(n2337), .Z(rd_data1[28]) );
  B5IP U2481 ( .A(wr_data[0]), .Z(n3358) );
  AN2I U2482 ( .A(wr_addr[2]), .B(wr_addr[1]), .Z(n2341) );
  IVI U2483 ( .A(wr_addr[0]), .Z(n2339) );
  ND2I U2484 ( .A(n2341), .B(n2339), .Z(n3355) );
  AN2I U2485 ( .A(wr_addr[4]), .B(RegWrite), .Z(n2348) );
  ND2I U2486 ( .A(wr_addr[3]), .B(n2348), .Z(n2346) );
  OR2P U2487 ( .A(n3355), .B(n2346), .Z(n3772) );
  B4I U2488 ( .A(n3772), .Z(n3976) );
  MUX21L U2489 ( .A(n4884), .B(n3358), .S(n3976), .Z(n2387) );
  IVI U2490 ( .A(wr_addr[1]), .Z(n2342) );
  NR2I U2491 ( .A(wr_addr[0]), .B(n2342), .Z(n2340) );
  IVI U2492 ( .A(wr_addr[2]), .Z(n2344) );
  ND2I U2493 ( .A(n2340), .B(n2344), .Z(n3357) );
  OR2P U2494 ( .A(n3357), .B(n2346), .Z(n3773) );
  B4I U2495 ( .A(n3773), .Z(n3977) );
  MUX21L U2496 ( .A(n4885), .B(n3358), .S(n3977), .Z(n2515) );
  ND2I U2497 ( .A(wr_addr[0]), .B(n2341), .Z(n3349) );
  OR2P U2498 ( .A(n3349), .B(n2346), .Z(n3771) );
  B4I U2499 ( .A(n3771), .Z(n3975) );
  MUX21L U2500 ( .A(n4840), .B(n3358), .S(n3975), .Z(n2355) );
  AN2I U2501 ( .A(wr_addr[0]), .B(n2342), .Z(n2345) );
  ND2I U2502 ( .A(wr_addr[2]), .B(n2345), .Z(n3350) );
  NR2I U2503 ( .A(n3350), .B(n2346), .Z(n4036) );
  IVI U2504 ( .A(n3525), .Z(n3467) );
  MUX21L U2505 ( .A(n4886), .B(n3358), .S(n3467), .Z(n2419) );
  NR2I U2506 ( .A(wr_addr[0]), .B(wr_addr[1]), .Z(n2343) );
  ND2I U2507 ( .A(wr_addr[2]), .B(n2343), .Z(n3351) );
  OR2P U2508 ( .A(n3351), .B(n2346), .Z(n4038) );
  IVI U2509 ( .A(n4038), .Z(n3468) );
  MUX21L U2510 ( .A(n4887), .B(n3358), .S(n3468), .Z(n2451) );
  ND2I U2511 ( .A(n2343), .B(n2344), .Z(n3352) );
  OR2P U2512 ( .A(n3352), .B(n2346), .Z(n4037) );
  IVI U2513 ( .A(n4037), .Z(n3469) );
  MUX21L U2514 ( .A(n4888), .B(n3358), .S(n3469), .Z(n2579) );
  OR2P U2515 ( .A(n3353), .B(n2346), .Z(n3526) );
  IVI U2516 ( .A(n3526), .Z(n4535) );
  MUX21L U2517 ( .A(n4889), .B(n3358), .S(n4535), .Z(n2483) );
  ND2I U2518 ( .A(n2345), .B(n2344), .Z(n3354) );
  NR2I U2519 ( .A(n3354), .B(n2346), .Z(n3398) );
  B5IP U2520 ( .A(n2347), .Z(n3983) );
  MUX21L U2521 ( .A(n4890), .B(n3358), .S(n3983), .Z(n2547) );
  IVI U2522 ( .A(wr_addr[3]), .Z(n2352) );
  ND2I U2523 ( .A(n2348), .B(n2352), .Z(n2351) );
  OR2P U2524 ( .A(n3351), .B(n2351), .Z(n4039) );
  IVI U2525 ( .A(n4039), .Z(n3470) );
  MUX21L U2526 ( .A(n4891), .B(n3358), .S(n3470), .Z(n2707) );
  OR2P U2527 ( .A(n3357), .B(n2351), .Z(n3774) );
  B4I U2528 ( .A(n3774), .Z(n3978) );
  MUX21L U2529 ( .A(n4892), .B(n3358), .S(n3978), .Z(n2771) );
  OR2P U2530 ( .A(n3349), .B(n2351), .Z(n3527) );
  B4I U2531 ( .A(n3527), .Z(n4536) );
  MUX21L U2532 ( .A(n4893), .B(n3358), .S(n4536), .Z(n2611) );
  NR2I U2533 ( .A(n3350), .B(n2351), .Z(n3396) );
  B5IP U2534 ( .A(n2349), .Z(n3996) );
  MUX21L U2535 ( .A(n4894), .B(n3358), .S(n3996), .Z(n2675) );
  OR2P U2536 ( .A(n3352), .B(n2351), .Z(n4040) );
  IVI U2537 ( .A(n4040), .Z(n3471) );
  MUX21L U2538 ( .A(n4895), .B(n3358), .S(n3471), .Z(n2835) );
  OR2P U2539 ( .A(n3353), .B(n2351), .Z(n3530) );
  IVI U2540 ( .A(n3530), .Z(n4537) );
  MUX21L U2541 ( .A(n4896), .B(n3358), .S(n4537), .Z(n2739) );
  NR2I U2542 ( .A(n3354), .B(n2351), .Z(n3397) );
  B5IP U2543 ( .A(n2350), .Z(n3999) );
  MUX21L U2544 ( .A(n4897), .B(n3358), .S(n3999), .Z(n2803) );
  NR2I U2545 ( .A(n3355), .B(n2351), .Z(n3528) );
  MUX21L U2546 ( .A(n4762), .B(n3358), .S(n4538), .Z(n2643) );
  AN2I U2547 ( .A(RegWrite), .B(n2352), .Z(n2353) );
  IVI U2548 ( .A(wr_addr[4]), .Z(n3348) );
  ND2I U2549 ( .A(n2353), .B(n3348), .Z(n2354) );
  OR2P U2550 ( .A(n3351), .B(n2354), .Z(n4048) );
  IVI U2551 ( .A(n4048), .Z(n3479) );
  MUX21L U2552 ( .A(n4898), .B(n3358), .S(n3479), .Z(n3219) );
  OR2P U2553 ( .A(n2354), .B(n3357), .Z(n3534) );
  B4I U2554 ( .A(n3534), .Z(n4540) );
  MUX21L U2555 ( .A(n4899), .B(n3358), .S(n4540), .Z(n3283) );
  OR2P U2556 ( .A(n2354), .B(n3349), .Z(n4049) );
  IVI U2557 ( .A(n4049), .Z(n3480) );
  MUX21L U2558 ( .A(n4900), .B(n3358), .S(n3480), .Z(n3123) );
  OR2P U2559 ( .A(n2354), .B(n3355), .Z(n4050) );
  IVI U2560 ( .A(n4050), .Z(n3481) );
  MUX21L U2561 ( .A(n4901), .B(n3358), .S(n3481), .Z(n3155) );
  NR2I U2562 ( .A(n2354), .B(n3350), .Z(n4051) );
  IVI U2563 ( .A(n3535), .Z(n3482) );
  MUX21L U2564 ( .A(n5669), .B(n3358), .S(n3482), .Z(n3187) );
  NR2I U2565 ( .A(n2354), .B(n3354), .Z(n4052) );
  IVI U2566 ( .A(n3536), .Z(n3483) );
  MUX21L U2567 ( .A(n5670), .B(n3358), .S(n3483), .Z(n3315) );
  OR2P U2568 ( .A(n2354), .B(n3353), .Z(n3347) );
  B4IP U2569 ( .A(n3347), .Z(n4620) );
  MUX21L U2570 ( .A(n5671), .B(n3358), .S(n4620), .Z(n3251) );
  OR2P U2571 ( .A(n3356), .B(n3349), .Z(n4046) );
  IVI U2572 ( .A(n4046), .Z(n3477) );
  MUX21L U2573 ( .A(n4902), .B(n3358), .S(n3477), .Z(n2867) );
  NR2I U2574 ( .A(n3356), .B(n3350), .Z(n4047) );
  IVI U2575 ( .A(n3531), .Z(n3478) );
  MUX21L U2576 ( .A(n4777), .B(n3358), .S(n3478), .Z(n2931) );
  OR2P U2577 ( .A(n3351), .B(n3356), .Z(n4041) );
  IVI U2578 ( .A(n4041), .Z(n3472) );
  MUX21L U2579 ( .A(n4903), .B(n3358), .S(n3472), .Z(n2963) );
  OR2P U2580 ( .A(n3356), .B(n3352), .Z(n4042) );
  IVI U2581 ( .A(n4042), .Z(n3473) );
  MUX21L U2582 ( .A(n4904), .B(n3358), .S(n3473), .Z(n3091) );
  OR2P U2583 ( .A(n3356), .B(n3353), .Z(n3532) );
  IVI U2584 ( .A(n3532), .Z(n4539) );
  MUX21L U2585 ( .A(n4905), .B(n3358), .S(n4539), .Z(n2995) );
  NR2I U2586 ( .A(n3356), .B(n3354), .Z(n4043) );
  IVI U2587 ( .A(n3533), .Z(n3474) );
  MUX21L U2588 ( .A(n4906), .B(n3358), .S(n3474), .Z(n3059) );
  OR2P U2589 ( .A(n3356), .B(n3355), .Z(n4044) );
  IVI U2590 ( .A(n4044), .Z(n3475) );
  MUX21L U2591 ( .A(n4907), .B(n3358), .S(n3475), .Z(n2899) );
  OR2P U2592 ( .A(n3357), .B(n3356), .Z(n4045) );
  IVI U2593 ( .A(n4045), .Z(n3476) );
  MUX21L U2594 ( .A(n298), .B(n3358), .S(n3476), .Z(n3027) );
  AO2 U2595 ( .A(\gpr[25][0] ), .B(n4001), .C(\gpr[28][0] ), .D(n4498), .Z(
        n3364) );
  IVI U2596 ( .A(n3485), .Z(n4357) );
  AO2 U2597 ( .A(\gpr[29][0] ), .B(n4090), .C(\gpr[24][0] ), .D(n4357), .Z(
        n3363) );
  IVI U2598 ( .A(n4356), .Z(n4487) );
  IVI U2599 ( .A(n3539), .Z(n3897) );
  IVI U2600 ( .A(n3897), .Z(n4457) );
  AO2 U2601 ( .A(\gpr[26][0] ), .B(n4487), .C(\gpr[31][0] ), .D(n4457), .Z(
        n3362) );
  ND2I U2602 ( .A(\gpr[30][0] ), .B(n4489), .Z(n3360) );
  ND2I U2603 ( .A(\gpr[27][0] ), .B(n4501), .Z(n3359) );
  AN3 U2604 ( .A(n4453), .B(n3360), .C(n3359), .Z(n3361) );
  ND4 U2605 ( .A(n3364), .B(n3363), .C(n3362), .D(n3361), .Z(n3375) );
  IVI U2606 ( .A(n4054), .Z(n3660) );
  AO2 U2607 ( .A(\gpr[19][0] ), .B(n3660), .C(\gpr[16][0] ), .D(n4357), .Z(
        n3373) );
  IVI U2608 ( .A(n3365), .Z(n3366) );
  IVI U2609 ( .A(n3366), .Z(n4653) );
  AO2 U2610 ( .A(\gpr[18][0] ), .B(n4622), .C(\gpr[21][0] ), .D(n4653), .Z(
        n3372) );
  AO2 U2611 ( .A(\gpr[20][0] ), .B(n4624), .C(\gpr[22][0] ), .D(n4431), .Z(
        n3371) );
  IVI U2612 ( .A(n3897), .Z(n4374) );
  ND2I U2613 ( .A(\gpr[23][0] ), .B(n4374), .Z(n3369) );
  ND2I U2614 ( .A(\gpr[17][0] ), .B(n4001), .Z(n3368) );
  AN3 U2615 ( .A(n4628), .B(n3369), .C(n3368), .Z(n3370) );
  ND4 U2616 ( .A(n3373), .B(n3372), .C(n3371), .D(n3370), .Z(n3374) );
  AN2I U2617 ( .A(n3375), .B(n3374), .Z(n3395) );
  ND2I U2618 ( .A(\gpr[6][0] ), .B(n4674), .Z(n3378) );
  ND2I U2619 ( .A(n4777), .B(n3833), .Z(n3376) );
  AO3 U2620 ( .A(\gpr[15][0] ), .B(n4653), .C(n4652), .D(n3376), .Z(n3377) );
  AN3 U2621 ( .A(n3378), .B(n4561), .C(n3377), .Z(n3393) );
  B2IP U2622 ( .A(n4308), .Z2(n4666) );
  ND2I U2623 ( .A(\gpr[3][0] ), .B(n4657), .Z(n3380) );
  ND2I U2624 ( .A(\gpr[5][0] ), .B(n4658), .Z(n3379) );
  ND2I U2625 ( .A(n3380), .B(n3379), .Z(n3384) );
  ND2I U2626 ( .A(\gpr[1][0] ), .B(n4656), .Z(n3382) );
  ND2I U2627 ( .A(\gpr[2][0] ), .B(n4659), .Z(n3381) );
  ND2I U2628 ( .A(n3382), .B(n3381), .Z(n3383) );
  NR2I U2629 ( .A(n3384), .B(n3383), .Z(n3391) );
  IVI U2630 ( .A(n3485), .Z(n4432) );
  AO2 U2631 ( .A(\gpr[8][0] ), .B(n4432), .C(\gpr[14][0] ), .D(n4431), .Z(
        n3388) );
  AO2 U2632 ( .A(\gpr[11][0] ), .B(n3660), .C(\gpr[12][0] ), .D(n4498), .Z(
        n3387) );
  ND2I U2633 ( .A(\gpr[9][0] ), .B(n4490), .Z(n3386) );
  IVI U2634 ( .A(n3538), .Z(n4622) );
  ND2I U2635 ( .A(\gpr[10][0] ), .B(n4622), .Z(n3385) );
  ND4 U2636 ( .A(n3388), .B(n3387), .C(n3386), .D(n3385), .Z(n3389) );
  ND2I U2637 ( .A(n4442), .B(n3389), .Z(n3390) );
  ND4 U2638 ( .A(n3393), .B(n3392), .C(n3391), .D(n3390), .Z(n3394) );
  AN2I U2639 ( .A(n3395), .B(n3394), .Z(rd_data2[0]) );
  B4IP U2640 ( .A(wr_data[1]), .Z(n3399) );
  MUX21L U2641 ( .A(n4908), .B(n3399), .S(n3470), .Z(n2708) );
  MUX21L U2642 ( .A(n4909), .B(n3399), .S(n4537), .Z(n2740) );
  MUX21L U2643 ( .A(n4910), .B(n3399), .S(n4536), .Z(n2612) );
  B2IP U2644 ( .A(n3396), .Z1(n2349), .Z2(n4590) );
  MUX21L U2645 ( .A(n4841), .B(n3399), .S(n4590), .Z(n2676) );
  MUX21L U2646 ( .A(n5672), .B(n3399), .S(n3471), .Z(n2836) );
  B2IP U2647 ( .A(n3397), .Z1(n2350), .Z2(n4593) );
  MUX21L U2648 ( .A(n5673), .B(n3399), .S(n4593), .Z(n2804) );
  MUX21L U2649 ( .A(n5674), .B(n3399), .S(n4538), .Z(n2644) );
  MUX21L U2650 ( .A(n4836), .B(n3399), .S(n3978), .Z(n2772) );
  MUX21L U2651 ( .A(n4911), .B(n3399), .S(n3478), .Z(n2932) );
  MUX21L U2652 ( .A(n4912), .B(n3399), .S(n3477), .Z(n2868) );
  MUX21L U2653 ( .A(n4913), .B(n3399), .S(n3479), .Z(n3220) );
  MUX21L U2654 ( .A(n4914), .B(n3399), .S(n4540), .Z(n3284) );
  MUX21L U2655 ( .A(n4915), .B(n3399), .S(n4620), .Z(n3252) );
  MUX21L U2656 ( .A(n4916), .B(n3399), .S(n3472), .Z(n2964) );
  MUX21L U2657 ( .A(n5675), .B(n3399), .S(n3473), .Z(n3092) );
  MUX21L U2658 ( .A(n4917), .B(n3399), .S(n4539), .Z(n2996) );
  MUX21L U2659 ( .A(n4918), .B(n3399), .S(n3474), .Z(n3060) );
  MUX21L U2660 ( .A(n4760), .B(n3399), .S(n3475), .Z(n2900) );
  MUX21L U2661 ( .A(n4838), .B(n3399), .S(n3476), .Z(n3028) );
  MUX21L U2662 ( .A(n4837), .B(n3399), .S(n3480), .Z(n3124) );
  MUX21L U2663 ( .A(n4919), .B(n3399), .S(n3481), .Z(n3156) );
  MUX21L U2664 ( .A(n5676), .B(n3399), .S(n3482), .Z(n3188) );
  MUX21L U2665 ( .A(n4920), .B(n3399), .S(n3483), .Z(n3316) );
  MUX21L U2666 ( .A(n5677), .B(n3399), .S(n3975), .Z(n2356) );
  MUX21L U2667 ( .A(n4827), .B(n3399), .S(n3467), .Z(n2420) );
  MUX21L U2668 ( .A(n4921), .B(n3399), .S(n3468), .Z(n2452) );
  MUX21L U2669 ( .A(n4922), .B(n3399), .S(n3469), .Z(n2580) );
  MUX21L U2670 ( .A(n5678), .B(n3399), .S(n4535), .Z(n2484) );
  B2IP U2671 ( .A(n3398), .Z1(n2347), .Z2(n4601) );
  MUX21L U2672 ( .A(n5679), .B(n3399), .S(n4601), .Z(n2548) );
  MUX21L U2673 ( .A(n4923), .B(n3399), .S(n3976), .Z(n2388) );
  MUX21L U2674 ( .A(n4835), .B(n3399), .S(n3977), .Z(n2516) );
  IVI U2675 ( .A(n3400), .Z(n4636) );
  AO2 U2676 ( .A(\gpr[27][1] ), .B(n3660), .C(\gpr[25][1] ), .D(n4636), .Z(
        n3407) );
  IVI U2677 ( .A(n3485), .Z(n4542) );
  AO2 U2678 ( .A(\gpr[24][1] ), .B(n4542), .C(\gpr[28][1] ), .D(n220), .Z(
        n3406) );
  AO2 U2679 ( .A(\gpr[30][1] ), .B(n4431), .C(\gpr[29][1] ), .D(n4653), .Z(
        n3405) );
  B2IP U2680 ( .A(n3538), .Z1(n3703), .Z2(n4356) );
  ND2I U2681 ( .A(\gpr[31][1] ), .B(n4543), .Z(n3402) );
  AO3 U2682 ( .A(n4356), .B(n4835), .C(n4641), .D(n3402), .Z(n3403) );
  IVI U2683 ( .A(n3403), .Z(n3404) );
  IVI U2684 ( .A(n3485), .Z(n4626) );
  AO2 U2685 ( .A(\gpr[16][1] ), .B(n4626), .C(\gpr[17][1] ), .D(n4636), .Z(
        n3413) );
  AO2 U2686 ( .A(\gpr[19][1] ), .B(n3660), .C(\gpr[21][1] ), .D(n4653), .Z(
        n3412) );
  AO2 U2687 ( .A(\gpr[20][1] ), .B(n219), .C(\gpr[22][1] ), .D(n4431), .Z(
        n3411) );
  IVI U2688 ( .A(n4130), .Z(n4548) );
  ND2I U2689 ( .A(\gpr[23][1] ), .B(n4548), .Z(n3408) );
  AO3 U2690 ( .A(n4356), .B(n4836), .C(n4628), .D(n3408), .Z(n3409) );
  IVI U2691 ( .A(n3409), .Z(n3410) );
  AO2 U2692 ( .A(\gpr[6][1] ), .B(n4475), .C(\gpr[15][1] ), .D(n4572), .Z(
        n3420) );
  NR2I U2693 ( .A(n4837), .B(n3414), .Z(n3418) );
  ND2I U2694 ( .A(\gpr[5][1] ), .B(n4658), .Z(n3416) );
  ND2I U2695 ( .A(\gpr[1][1] ), .B(n4656), .Z(n3415) );
  ND2I U2696 ( .A(n3416), .B(n3415), .Z(n3417) );
  NR2I U2697 ( .A(n3418), .B(n3417), .Z(n3419) );
  AN2I U2698 ( .A(n3420), .B(n3419), .Z(n3432) );
  ND2I U2699 ( .A(\gpr[4][1] ), .B(n4666), .Z(n3422) );
  ND2I U2700 ( .A(n4578), .B(\gpr[13][1] ), .Z(n3421) );
  ND2I U2701 ( .A(\gpr[14][1] ), .B(n4489), .Z(n3423) );
  AO3 U2702 ( .A(n4838), .B(n4356), .C(n295), .D(n3423), .Z(n3430) );
  ND2I U2703 ( .A(\gpr[9][1] ), .B(n4490), .Z(n3427) );
  ND2I U2704 ( .A(\gpr[8][1] ), .B(n4357), .Z(n3426) );
  ND2I U2705 ( .A(\gpr[11][1] ), .B(n4501), .Z(n3425) );
  ND2I U2706 ( .A(\gpr[12][1] ), .B(n4624), .Z(n3424) );
  ND4 U2707 ( .A(n3427), .B(n3426), .C(n3425), .D(n3424), .Z(n3429) );
  ND2I U2708 ( .A(n3428), .B(n4561), .Z(n4362) );
  AO7 U2709 ( .A(n3430), .B(n3429), .C(n4362), .Z(n3431) );
  B4IP U2710 ( .A(wr_data[2]), .Z(n3433) );
  MUX21L U2711 ( .A(n4924), .B(n3433), .S(n3467), .Z(n2421) );
  MUX21L U2712 ( .A(n4925), .B(n3433), .S(n3468), .Z(n2453) );
  MUX21L U2713 ( .A(n4926), .B(n3433), .S(n3469), .Z(n2581) );
  MUX21L U2714 ( .A(n4927), .B(n3433), .S(n4535), .Z(n2485) );
  MUX21L U2715 ( .A(n4842), .B(n3433), .S(n3976), .Z(n2389) );
  MUX21L U2716 ( .A(n4928), .B(n3433), .S(n3977), .Z(n2517) );
  MUX21L U2717 ( .A(n4929), .B(n3433), .S(n3983), .Z(n2549) );
  MUX21L U2718 ( .A(n4930), .B(n3433), .S(n3975), .Z(n2357) );
  MUX21L U2719 ( .A(n4931), .B(n3433), .S(n4536), .Z(n2613) );
  MUX21L U2720 ( .A(n4932), .B(n3433), .S(n3996), .Z(n2677) );
  MUX21L U2721 ( .A(n4933), .B(n3433), .S(n4537), .Z(n2741) );
  MUX21L U2722 ( .A(n4934), .B(n3433), .S(n3999), .Z(n2805) );
  MUX21L U2723 ( .A(n4763), .B(n3433), .S(n4538), .Z(n2645) );
  MUX21L U2724 ( .A(n4935), .B(n3433), .S(n3978), .Z(n2773) );
  MUX21L U2725 ( .A(n4936), .B(n3433), .S(n3471), .Z(n2837) );
  MUX21L U2726 ( .A(n4937), .B(n3433), .S(n3470), .Z(n2709) );
  MUX21L U2727 ( .A(n5680), .B(n3433), .S(n3472), .Z(n2965) );
  MUX21L U2728 ( .A(n4938), .B(n3433), .S(n3473), .Z(n3093) );
  MUX21L U2729 ( .A(n4939), .B(n3433), .S(n4539), .Z(n2997) );
  MUX21L U2730 ( .A(n4940), .B(n3433), .S(n3474), .Z(n3061) );
  MUX21L U2731 ( .A(n4812), .B(n3433), .S(n3475), .Z(n2901) );
  MUX21L U2732 ( .A(n4941), .B(n3433), .S(n3476), .Z(n3029) );
  MUX21L U2733 ( .A(n4942), .B(n3433), .S(n3477), .Z(n2869) );
  MUX21L U2734 ( .A(n4778), .B(n3433), .S(n3478), .Z(n2933) );
  MUX21L U2735 ( .A(n5681), .B(n3433), .S(n3479), .Z(n3221) );
  MUX21L U2736 ( .A(n4943), .B(n3433), .S(n4540), .Z(n3285) );
  MUX21L U2737 ( .A(n4944), .B(n3433), .S(n3480), .Z(n3125) );
  MUX21L U2738 ( .A(n4945), .B(n3433), .S(n3481), .Z(n3157) );
  MUX21L U2739 ( .A(n4946), .B(n3433), .S(n3482), .Z(n3189) );
  MUX21L U2740 ( .A(n4947), .B(n3433), .S(n3483), .Z(n3317) );
  MUX21L U2741 ( .A(n4948), .B(n3433), .S(n4620), .Z(n3253) );
  AO2 U2742 ( .A(\gpr[26][2] ), .B(n4487), .C(\gpr[24][2] ), .D(n4637), .Z(
        n3439) );
  AO2 U2743 ( .A(\gpr[27][2] ), .B(n3660), .C(\gpr[28][2] ), .D(n4624), .Z(
        n3438) );
  AO2 U2744 ( .A(\gpr[29][2] ), .B(n4653), .C(\gpr[31][2] ), .D(n4374), .Z(
        n3437) );
  ND2I U2745 ( .A(\gpr[30][2] ), .B(n4625), .Z(n3435) );
  ND2I U2746 ( .A(\gpr[25][2] ), .B(n4490), .Z(n3434) );
  AN3 U2747 ( .A(n4641), .B(n3435), .C(n3434), .Z(n3436) );
  ND4 U2748 ( .A(n3439), .B(n3438), .C(n3437), .D(n3436), .Z(n3445) );
  AO2 U2749 ( .A(\gpr[20][2] ), .B(n4624), .C(\gpr[18][2] ), .D(n4622), .Z(
        n3443) );
  AO2 U2750 ( .A(\gpr[19][2] ), .B(n3660), .C(\gpr[17][2] ), .D(n4636), .Z(
        n3442) );
  AO2 U2751 ( .A(\gpr[21][2] ), .B(n4653), .C(\gpr[22][2] ), .D(n4431), .Z(
        n3441) );
  IVI U2752 ( .A(n3897), .Z(n4209) );
  IVI U2753 ( .A(n3485), .Z(n4497) );
  ND4 U2754 ( .A(n3443), .B(n3442), .C(n3441), .D(n3440), .Z(n3444) );
  AN2I U2755 ( .A(n3445), .B(n3444), .Z(n3466) );
  ND2I U2756 ( .A(n4625), .B(n4442), .Z(n3446) );
  IVI U2757 ( .A(n3446), .Z(n3589) );
  ND2I U2758 ( .A(n4778), .B(n3833), .Z(n3447) );
  AO3 U2759 ( .A(\gpr[15][2] ), .B(n4653), .C(n4652), .D(n3447), .Z(n3448) );
  AO3 U2760 ( .A(n4812), .B(n4108), .C(n295), .D(n3448), .Z(n3454) );
  ND2I U2761 ( .A(\gpr[3][2] ), .B(n4657), .Z(n3452) );
  ND2I U2762 ( .A(\gpr[5][2] ), .B(n4658), .Z(n3451) );
  ND2I U2763 ( .A(\gpr[1][2] ), .B(n4656), .Z(n3450) );
  ND2I U2764 ( .A(\gpr[4][2] ), .B(n4666), .Z(n3449) );
  ND4 U2765 ( .A(n3452), .B(n3451), .C(n3450), .D(n3449), .Z(n3453) );
  NR2I U2766 ( .A(n3454), .B(n3453), .Z(n3464) );
  ND2I U2767 ( .A(\gpr[2][2] ), .B(n4659), .Z(n3458) );
  AN2I U2768 ( .A(n3703), .B(n4442), .Z(n4473) );
  ND2I U2769 ( .A(n4473), .B(\gpr[10][2] ), .Z(n3457) );
  B2I U2770 ( .A(n3558), .Z2(n4668) );
  ND2I U2771 ( .A(\gpr[9][2] ), .B(n4668), .Z(n3456) );
  IVI U2772 ( .A(n3561), .Z(n4519) );
  ND2I U2773 ( .A(\gpr[8][2] ), .B(n4519), .Z(n3455) );
  ND2I U2774 ( .A(\gpr[11][2] ), .B(n4667), .Z(n3462) );
  ND2I U2775 ( .A(\gpr[12][2] ), .B(n4673), .Z(n3461) );
  ND2I U2776 ( .A(\gpr[7][2] ), .B(n4675), .Z(n3460) );
  IVI U2777 ( .A(n3562), .Z(n4197) );
  ND2I U2778 ( .A(\gpr[6][2] ), .B(n4197), .Z(n3459) );
  ND2I U2779 ( .A(n3464), .B(n3463), .Z(n3465) );
  AN2I U2780 ( .A(n3466), .B(n3465), .Z(rd_data2[2]) );
  B4IP U2781 ( .A(wr_data[3]), .Z(n3484) );
  MUX21L U2782 ( .A(n4949), .B(n3484), .S(n3467), .Z(n2422) );
  MUX21L U2783 ( .A(n4950), .B(n3484), .S(n3468), .Z(n2454) );
  MUX21L U2784 ( .A(n4951), .B(n3484), .S(n3469), .Z(n2582) );
  MUX21L U2785 ( .A(n4952), .B(n3484), .S(n4535), .Z(n2486) );
  MUX21L U2786 ( .A(n4953), .B(n3484), .S(n4601), .Z(n2550) );
  MUX21L U2787 ( .A(n4843), .B(n3484), .S(n3976), .Z(n2390) );
  MUX21L U2788 ( .A(n4779), .B(n3484), .S(n3977), .Z(n2518) );
  MUX21L U2789 ( .A(n4954), .B(n3484), .S(n3975), .Z(n2358) );
  MUX21L U2790 ( .A(n4955), .B(n3484), .S(n4590), .Z(n2678) );
  MUX21L U2791 ( .A(n4956), .B(n3484), .S(n3470), .Z(n2710) );
  MUX21L U2792 ( .A(n4957), .B(n3484), .S(n3471), .Z(n2838) );
  MUX21L U2793 ( .A(n4958), .B(n3484), .S(n4537), .Z(n2742) );
  MUX21L U2794 ( .A(n4764), .B(n3484), .S(n4538), .Z(n2646) );
  MUX21L U2795 ( .A(n299), .B(n3484), .S(n3978), .Z(n2774) );
  MUX21L U2796 ( .A(n4959), .B(n3484), .S(n4593), .Z(n2806) );
  MUX21L U2797 ( .A(n4960), .B(n3484), .S(n4536), .Z(n2614) );
  MUX21L U2798 ( .A(n4961), .B(n3484), .S(n3472), .Z(n2966) );
  MUX21L U2799 ( .A(n4962), .B(n3484), .S(n3473), .Z(n3094) );
  MUX21L U2800 ( .A(n4963), .B(n3484), .S(n4539), .Z(n2998) );
  MUX21L U2801 ( .A(n4964), .B(n3484), .S(n3474), .Z(n3062) );
  MUX21L U2802 ( .A(n4813), .B(n3484), .S(n3475), .Z(n2902) );
  MUX21L U2803 ( .A(n4965), .B(n3484), .S(n3476), .Z(n3030) );
  MUX21L U2804 ( .A(n4966), .B(n3484), .S(n3477), .Z(n2870) );
  MUX21L U2805 ( .A(n4780), .B(n3484), .S(n3478), .Z(n2934) );
  MUX21L U2806 ( .A(n4967), .B(n3484), .S(n3479), .Z(n3222) );
  MUX21L U2807 ( .A(n4968), .B(n3484), .S(n4540), .Z(n3286) );
  MUX21L U2808 ( .A(n4969), .B(n3484), .S(n3480), .Z(n3126) );
  MUX21L U2809 ( .A(n4970), .B(n3484), .S(n3481), .Z(n3158) );
  MUX21L U2810 ( .A(n4971), .B(n3484), .S(n3482), .Z(n3190) );
  MUX21L U2811 ( .A(n4972), .B(n3484), .S(n3483), .Z(n3318) );
  MUX21L U2812 ( .A(n4973), .B(n3484), .S(n4620), .Z(n3254) );
  IVI U2813 ( .A(n3485), .Z(n4549) );
  AO2 U2814 ( .A(\gpr[25][3] ), .B(n4296), .C(\gpr[24][3] ), .D(n4549), .Z(
        n3491) );
  AO2 U2815 ( .A(\gpr[27][3] ), .B(n3660), .C(\gpr[28][3] ), .D(n4498), .Z(
        n3490) );
  AO2 U2816 ( .A(\gpr[29][3] ), .B(n4653), .C(\gpr[31][3] ), .D(n4374), .Z(
        n3489) );
  ND2I U2817 ( .A(\gpr[30][3] ), .B(n4625), .Z(n3486) );
  AO3 U2818 ( .A(n4356), .B(n4779), .C(n4641), .D(n3486), .Z(n3487) );
  IVI U2819 ( .A(n3487), .Z(n3488) );
  ND4 U2820 ( .A(n3491), .B(n3490), .C(n3489), .D(n3488), .Z(n3499) );
  AO2 U2821 ( .A(\gpr[16][3] ), .B(n4450), .C(\gpr[18][3] ), .D(n4622), .Z(
        n3497) );
  AO2 U2822 ( .A(\gpr[19][3] ), .B(n3660), .C(\gpr[20][3] ), .D(n220), .Z(
        n3496) );
  AO2 U2823 ( .A(\gpr[21][3] ), .B(n4653), .C(\gpr[23][3] ), .D(n4209), .Z(
        n3495) );
  ND2I U2824 ( .A(\gpr[22][3] ), .B(n4625), .Z(n3493) );
  ND2I U2825 ( .A(\gpr[17][3] ), .B(n4490), .Z(n3492) );
  AN3 U2826 ( .A(n4628), .B(n3493), .C(n3492), .Z(n3494) );
  ND4 U2827 ( .A(n3497), .B(n3496), .C(n3495), .D(n3494), .Z(n3498) );
  AN2I U2828 ( .A(n3499), .B(n3498), .Z(n3524) );
  IVI U2829 ( .A(n3589), .Z(n4466) );
  ND2I U2830 ( .A(n4780), .B(n3833), .Z(n3500) );
  AO3 U2831 ( .A(\gpr[15][3] ), .B(n4653), .C(n4652), .D(n3500), .Z(n3501) );
  AO3 U2832 ( .A(n4813), .B(n4466), .C(n295), .D(n3501), .Z(n3507) );
  ND2I U2833 ( .A(\gpr[3][3] ), .B(n4657), .Z(n3505) );
  ND2I U2834 ( .A(\gpr[5][3] ), .B(n4658), .Z(n3504) );
  ND2I U2835 ( .A(\gpr[1][3] ), .B(n4656), .Z(n3503) );
  ND2I U2836 ( .A(\gpr[4][3] ), .B(n4666), .Z(n3502) );
  ND4 U2837 ( .A(n3505), .B(n3504), .C(n3503), .D(n3502), .Z(n3506) );
  NR2I U2838 ( .A(n3507), .B(n3506), .Z(n3522) );
  ND2I U2839 ( .A(\gpr[2][3] ), .B(n4659), .Z(n3512) );
  ND2I U2840 ( .A(n3679), .B(\gpr[10][3] ), .Z(n3511) );
  IVI U2841 ( .A(n3598), .Z(n4314) );
  B2I U2842 ( .A(n4314), .Z2(n4563) );
  ND2I U2843 ( .A(\gpr[9][3] ), .B(n4563), .Z(n3510) );
  IVI U2844 ( .A(n3508), .Z(n4315) );
  ND2I U2845 ( .A(\gpr[8][3] ), .B(n4315), .Z(n3509) );
  ND4 U2846 ( .A(n3512), .B(n3511), .C(n3510), .D(n3509), .Z(n3520) );
  IVI U2847 ( .A(n3513), .Z(n4571) );
  ND2I U2848 ( .A(\gpr[11][3] ), .B(n4571), .Z(n3518) );
  IVI U2849 ( .A(n3514), .Z(n4573) );
  ND2I U2850 ( .A(\gpr[12][3] ), .B(n4573), .Z(n3517) );
  ND2I U2851 ( .A(\gpr[7][3] ), .B(n4675), .Z(n3516) );
  IVI U2852 ( .A(n3562), .Z(n4354) );
  ND2I U2853 ( .A(\gpr[6][3] ), .B(n4354), .Z(n3515) );
  ND4 U2854 ( .A(n3518), .B(n3517), .C(n3516), .D(n3515), .Z(n3519) );
  NR2I U2855 ( .A(n3520), .B(n3519), .Z(n3521) );
  ND2I U2856 ( .A(n3522), .B(n3521), .Z(n3523) );
  AN2I U2857 ( .A(n3524), .B(n3523), .Z(rd_data2[3]) );
  MUX21L U2858 ( .A(n4974), .B(n3537), .S(n3975), .Z(n2359) );
  B4I U2859 ( .A(n3525), .Z(n3981) );
  MUX21L U2860 ( .A(n4975), .B(n3537), .S(n3981), .Z(n2423) );
  B4I U2861 ( .A(n4038), .Z(n3980) );
  MUX21L U2862 ( .A(n4976), .B(n3537), .S(n3980), .Z(n2455) );
  B5IP U2863 ( .A(n3526), .Z(n4600) );
  MUX21L U2864 ( .A(n4977), .B(n3537), .S(n4600), .Z(n2487) );
  MUX21L U2865 ( .A(n4806), .B(n3537), .S(n3976), .Z(n2391) );
  MUX21L U2866 ( .A(n4978), .B(n3537), .S(n3977), .Z(n2519) );
  B4I U2867 ( .A(n4037), .Z(n3982) );
  MUX21L U2868 ( .A(n4979), .B(n3537), .S(n3982), .Z(n2583) );
  MUX21L U2869 ( .A(n4980), .B(n3537), .S(n3983), .Z(n2551) );
  B5IP U2870 ( .A(n3527), .Z(n4597) );
  MUX21L U2871 ( .A(n4981), .B(n3537), .S(n4597), .Z(n2615) );
  MUX21L U2872 ( .A(n4982), .B(n3537), .S(n3996), .Z(n2679) );
  B4I U2873 ( .A(n4039), .Z(n3997) );
  MUX21L U2874 ( .A(n4983), .B(n3537), .S(n3997), .Z(n2711) );
  B4I U2875 ( .A(n4040), .Z(n3998) );
  MUX21L U2876 ( .A(n4984), .B(n3537), .S(n3998), .Z(n2839) );
  B2IP U2877 ( .A(n3528), .Z1(n3529), .Z2(n4538) );
  B4I U2878 ( .A(n3529), .Z(n4594) );
  MUX21L U2879 ( .A(n4805), .B(n3537), .S(n4594), .Z(n2647) );
  MUX21L U2880 ( .A(n4985), .B(n3537), .S(n3978), .Z(n2775) );
  MUX21L U2881 ( .A(n4986), .B(n3537), .S(n3999), .Z(n2807) );
  B5IP U2882 ( .A(n3530), .Z(n4592) );
  MUX21L U2883 ( .A(n4987), .B(n3537), .S(n4592), .Z(n2743) );
  B4I U2884 ( .A(n3531), .Z(n3985) );
  MUX21L U2885 ( .A(n5682), .B(n3537), .S(n3985), .Z(n2935) );
  B4I U2886 ( .A(n4046), .Z(n3984) );
  MUX21L U2887 ( .A(n5683), .B(n3537), .S(n3984), .Z(n2871) );
  B4I U2888 ( .A(n4041), .Z(n3988) );
  MUX21L U2889 ( .A(n4988), .B(n3537), .S(n3988), .Z(n2967) );
  B4I U2890 ( .A(n4042), .Z(n3989) );
  MUX21L U2891 ( .A(n4989), .B(n3537), .S(n3989), .Z(n3095) );
  B5IP U2892 ( .A(n3532), .Z(n4608) );
  MUX21L U2893 ( .A(n5684), .B(n3537), .S(n4608), .Z(n2999) );
  B4I U2894 ( .A(n3533), .Z(n3990) );
  MUX21L U2895 ( .A(n5685), .B(n3537), .S(n3990), .Z(n3063) );
  B4I U2896 ( .A(n4044), .Z(n3991) );
  MUX21L U2897 ( .A(n5686), .B(n3537), .S(n3991), .Z(n2903) );
  B4I U2898 ( .A(n4045), .Z(n3992) );
  MUX21L U2899 ( .A(n4990), .B(n3537), .S(n3992), .Z(n3031) );
  B4I U2900 ( .A(n4048), .Z(n3986) );
  MUX21L U2901 ( .A(n4991), .B(n3537), .S(n3986), .Z(n3223) );
  B5IP U2902 ( .A(n3534), .Z(n4615) );
  MUX21L U2903 ( .A(n4992), .B(n3537), .S(n4615), .Z(n3287) );
  B4I U2904 ( .A(n4049), .Z(n3993) );
  MUX21L U2905 ( .A(n5687), .B(n3537), .S(n3993), .Z(n3127) );
  B4I U2906 ( .A(n4050), .Z(n3994) );
  MUX21L U2907 ( .A(n5688), .B(n3537), .S(n3994), .Z(n3159) );
  B4I U2908 ( .A(n3535), .Z(n3995) );
  MUX21L U2909 ( .A(n5689), .B(n3537), .S(n3995), .Z(n3191) );
  B4I U2910 ( .A(n3536), .Z(n3987) );
  MUX21L U2911 ( .A(n5690), .B(n3537), .S(n3987), .Z(n3319) );
  MUX21L U2912 ( .A(n5691), .B(n3537), .S(n4620), .Z(n3255) );
  IVI U2913 ( .A(n3538), .Z(n4458) );
  AO2 U2914 ( .A(\gpr[26][4] ), .B(n4458), .C(\gpr[25][4] ), .D(n4296), .Z(
        n3546) );
  AO2 U2915 ( .A(\gpr[28][4] ), .B(n4624), .C(\gpr[27][4] ), .D(n3660), .Z(
        n3545) );
  AO2 U2916 ( .A(\gpr[29][4] ), .B(n4653), .C(\gpr[30][4] ), .D(n4431), .Z(
        n3544) );
  IVI U2917 ( .A(n3539), .Z(n3785) );
  IVI U2918 ( .A(n3785), .Z(n4060) );
  AN2I U2919 ( .A(\gpr[31][4] ), .B(n4060), .Z(n3542) );
  ND2I U2920 ( .A(\gpr[24][4] ), .B(n4542), .Z(n3540) );
  ND2I U2921 ( .A(n4641), .B(n3540), .Z(n3541) );
  NR2I U2922 ( .A(n3542), .B(n3541), .Z(n3543) );
  ND4 U2923 ( .A(n3546), .B(n3545), .C(n3544), .D(n3543), .Z(n3554) );
  AO2 U2924 ( .A(\gpr[19][4] ), .B(n3660), .C(\gpr[18][4] ), .D(n4622), .Z(
        n3552) );
  AO2 U2925 ( .A(\gpr[16][4] ), .B(n4450), .C(\gpr[20][4] ), .D(n4498), .Z(
        n3551) );
  AO2 U2926 ( .A(\gpr[21][4] ), .B(n4653), .C(\gpr[22][4] ), .D(n4431), .Z(
        n3550) );
  ND2I U2927 ( .A(\gpr[23][4] ), .B(n4060), .Z(n3548) );
  ND2I U2928 ( .A(\gpr[17][4] ), .B(n4490), .Z(n3547) );
  AN3 U2929 ( .A(n4628), .B(n3548), .C(n3547), .Z(n3549) );
  ND4 U2930 ( .A(n3552), .B(n3551), .C(n3550), .D(n3549), .Z(n3553) );
  AN2I U2931 ( .A(n3554), .B(n3553), .Z(n3572) );
  ND2I U2932 ( .A(\gpr[1][4] ), .B(n4656), .Z(n3557) );
  ND2I U2933 ( .A(\gpr[3][4] ), .B(n4657), .Z(n3556) );
  ND2I U2934 ( .A(\gpr[5][4] ), .B(n4658), .Z(n3555) );
  ND4 U2935 ( .A(n295), .B(n3557), .C(n3556), .D(n3555), .Z(n3560) );
  NR2I U2936 ( .A(n3560), .B(n3559), .Z(n3570) );
  IVI U2937 ( .A(n3562), .Z(n4475) );
  ND2I U2938 ( .A(\gpr[6][4] ), .B(n4475), .Z(n3566) );
  ND2I U2939 ( .A(\gpr[13][4] ), .B(n4578), .Z(n3565) );
  ND2I U2940 ( .A(\gpr[7][4] ), .B(n4675), .Z(n3564) );
  ND2I U2941 ( .A(\gpr[14][4] ), .B(n4579), .Z(n3563) );
  ND4 U2942 ( .A(n3566), .B(n3565), .C(n3564), .D(n3563), .Z(n3567) );
  NR2I U2943 ( .A(n3568), .B(n3567), .Z(n3569) );
  ND2I U2944 ( .A(n3570), .B(n3569), .Z(n3571) );
  AN2I U2945 ( .A(n3572), .B(n3571), .Z(rd_data2[4]) );
  B4IP U2946 ( .A(wr_data[5]), .Z(n3573) );
  MUX21L U2947 ( .A(n4993), .B(n3573), .S(n3996), .Z(n2680) );
  MUX21L U2948 ( .A(n300), .B(n3573), .S(n3997), .Z(n2712) );
  MUX21L U2949 ( .A(n4994), .B(n3573), .S(n3998), .Z(n2840) );
  MUX21L U2950 ( .A(n4995), .B(n3573), .S(n4592), .Z(n2744) );
  MUX21L U2951 ( .A(n4844), .B(n3573), .S(n4594), .Z(n2648) );
  MUX21L U2952 ( .A(n4996), .B(n3573), .S(n3978), .Z(n2776) );
  MUX21L U2953 ( .A(n4997), .B(n3573), .S(n3999), .Z(n2808) );
  MUX21L U2954 ( .A(n4998), .B(n3573), .S(n4597), .Z(n2616) );
  MUX21L U2955 ( .A(n4999), .B(n3573), .S(n3981), .Z(n2424) );
  MUX21L U2956 ( .A(n4845), .B(n3573), .S(n3980), .Z(n2456) );
  MUX21L U2957 ( .A(n5000), .B(n3573), .S(n3982), .Z(n2584) );
  MUX21L U2958 ( .A(n5001), .B(n3573), .S(n3983), .Z(n2552) );
  MUX21L U2959 ( .A(n5002), .B(n3573), .S(n3976), .Z(n2392) );
  MUX21L U2960 ( .A(n5003), .B(n3573), .S(n3977), .Z(n2520) );
  MUX21L U2961 ( .A(n5004), .B(n3573), .S(n4600), .Z(n2488) );
  MUX21L U2962 ( .A(n5005), .B(n3573), .S(n3975), .Z(n2360) );
  MUX21L U2963 ( .A(n5006), .B(n3573), .S(n3988), .Z(n2968) );
  MUX21L U2964 ( .A(n5007), .B(n3573), .S(n3989), .Z(n3096) );
  MUX21L U2965 ( .A(n5008), .B(n3573), .S(n4608), .Z(n3000) );
  MUX21L U2966 ( .A(n5009), .B(n3573), .S(n3990), .Z(n3064) );
  MUX21L U2967 ( .A(n4814), .B(n3573), .S(n3991), .Z(n2904) );
  MUX21L U2968 ( .A(n5010), .B(n3573), .S(n3992), .Z(n3032) );
  MUX21L U2969 ( .A(n5011), .B(n3573), .S(n3984), .Z(n2872) );
  MUX21L U2970 ( .A(n4781), .B(n3573), .S(n3985), .Z(n2936) );
  MUX21L U2971 ( .A(n5012), .B(n3573), .S(n3986), .Z(n3224) );
  MUX21L U2972 ( .A(n5013), .B(n3573), .S(n4615), .Z(n3288) );
  MUX21L U2973 ( .A(n5014), .B(n3573), .S(n3993), .Z(n3128) );
  MUX21L U2974 ( .A(n5015), .B(n3573), .S(n3994), .Z(n3160) );
  MUX21L U2975 ( .A(n5016), .B(n3573), .S(n3995), .Z(n3192) );
  MUX21L U2976 ( .A(n5017), .B(n3573), .S(n3987), .Z(n3320) );
  MUX21L U2977 ( .A(n5018), .B(n3573), .S(n4620), .Z(n3256) );
  AO2 U2978 ( .A(\gpr[18][5] ), .B(n4214), .C(\gpr[16][5] ), .D(n4637), .Z(
        n3579) );
  AO2 U2979 ( .A(\gpr[19][5] ), .B(n3660), .C(\gpr[20][5] ), .D(n4498), .Z(
        n3578) );
  IVI U2980 ( .A(n3785), .Z(n4002) );
  AO2 U2981 ( .A(\gpr[21][5] ), .B(n4653), .C(\gpr[23][5] ), .D(n4002), .Z(
        n3577) );
  ND2I U2982 ( .A(\gpr[22][5] ), .B(n4625), .Z(n3575) );
  ND2I U2983 ( .A(\gpr[17][5] ), .B(n4490), .Z(n3574) );
  AN3 U2984 ( .A(n4628), .B(n3575), .C(n3574), .Z(n3576) );
  ND4 U2985 ( .A(n3579), .B(n3578), .C(n3577), .D(n3576), .Z(n3588) );
  AO2 U2986 ( .A(\gpr[26][5] ), .B(n4487), .C(\gpr[24][5] ), .D(n4497), .Z(
        n3586) );
  AO2 U2987 ( .A(\gpr[25][5] ), .B(n4001), .C(\gpr[28][5] ), .D(n4498), .Z(
        n3585) );
  AO2 U2988 ( .A(\gpr[29][5] ), .B(n4097), .C(\gpr[31][5] ), .D(n4060), .Z(
        n3584) );
  AN2I U2989 ( .A(\gpr[30][5] ), .B(n4625), .Z(n3582) );
  ND2I U2990 ( .A(\gpr[27][5] ), .B(n4501), .Z(n3580) );
  ND2I U2991 ( .A(n4641), .B(n3580), .Z(n3581) );
  NR2I U2992 ( .A(n3582), .B(n3581), .Z(n3583) );
  ND4 U2993 ( .A(n3586), .B(n3585), .C(n3584), .D(n3583), .Z(n3587) );
  AN2I U2994 ( .A(n3588), .B(n3587), .Z(n3613) );
  IVI U2995 ( .A(n3589), .Z(n4655) );
  ND2I U2996 ( .A(n4781), .B(n3833), .Z(n3590) );
  AO3 U2997 ( .A(\gpr[15][5] ), .B(n4097), .C(n4652), .D(n3590), .Z(n3591) );
  AO3 U2998 ( .A(n4814), .B(n4655), .C(n295), .D(n3591), .Z(n3597) );
  ND2I U2999 ( .A(\gpr[3][5] ), .B(n4657), .Z(n3595) );
  ND2I U3000 ( .A(\gpr[5][5] ), .B(n4658), .Z(n3594) );
  ND2I U3001 ( .A(\gpr[1][5] ), .B(n4656), .Z(n3593) );
  ND2I U3002 ( .A(\gpr[4][5] ), .B(n4666), .Z(n3592) );
  ND4 U3003 ( .A(n3595), .B(n3594), .C(n3593), .D(n3592), .Z(n3596) );
  NR2I U3004 ( .A(n3597), .B(n3596), .Z(n3611) );
  ND2I U3005 ( .A(\gpr[2][5] ), .B(n4659), .Z(n3603) );
  ND2I U3006 ( .A(n3679), .B(\gpr[10][5] ), .Z(n3602) );
  IVI U3007 ( .A(n3598), .Z(n4474) );
  B2I U3008 ( .A(n4474), .Z2(n4518) );
  ND2I U3009 ( .A(\gpr[9][5] ), .B(n4518), .Z(n3601) );
  ND2I U3010 ( .A(\gpr[8][5] ), .B(n3599), .Z(n3600) );
  ND4 U3011 ( .A(n3603), .B(n3602), .C(n3601), .D(n3600), .Z(n3609) );
  ND2I U3012 ( .A(\gpr[11][5] ), .B(n4667), .Z(n3607) );
  ND2I U3013 ( .A(\gpr[12][5] ), .B(n4673), .Z(n3606) );
  ND2I U3014 ( .A(\gpr[7][5] ), .B(n4675), .Z(n3605) );
  ND2I U3015 ( .A(\gpr[6][5] ), .B(n4475), .Z(n3604) );
  ND4 U3016 ( .A(n3607), .B(n3606), .C(n3605), .D(n3604), .Z(n3608) );
  NR2I U3017 ( .A(n3609), .B(n3608), .Z(n3610) );
  ND2I U3018 ( .A(n3611), .B(n3610), .Z(n3612) );
  AN2I U3019 ( .A(n3613), .B(n3612), .Z(rd_data2[5]) );
  B5IP U3020 ( .A(wr_data[6]), .Z(n3614) );
  MUX21L U3021 ( .A(n5019), .B(n3614), .S(n4597), .Z(n2617) );
  MUX21L U3022 ( .A(n5020), .B(n3614), .S(n3996), .Z(n2681) );
  MUX21L U3023 ( .A(n5021), .B(n3614), .S(n3997), .Z(n2713) );
  MUX21L U3024 ( .A(n301), .B(n3614), .S(n3998), .Z(n2841) );
  MUX21L U3025 ( .A(n4846), .B(n3614), .S(n4594), .Z(n2649) );
  MUX21L U3026 ( .A(n5022), .B(n3614), .S(n3978), .Z(n2777) );
  MUX21L U3027 ( .A(n5023), .B(n3614), .S(n3999), .Z(n2809) );
  MUX21L U3028 ( .A(n5024), .B(n3614), .S(n4592), .Z(n2745) );
  MUX21L U3029 ( .A(n5025), .B(n3614), .S(n3975), .Z(n2361) );
  MUX21L U3030 ( .A(n5026), .B(n3614), .S(n3981), .Z(n2425) );
  MUX21L U3031 ( .A(n5027), .B(n3614), .S(n3982), .Z(n2585) );
  MUX21L U3032 ( .A(n5028), .B(n3614), .S(n3983), .Z(n2553) );
  MUX21L U3033 ( .A(n4847), .B(n3614), .S(n3976), .Z(n2393) );
  MUX21L U3034 ( .A(n5029), .B(n3614), .S(n3977), .Z(n2521) );
  MUX21L U3035 ( .A(n5030), .B(n3614), .S(n4600), .Z(n2489) );
  MUX21L U3036 ( .A(n5031), .B(n3614), .S(n3980), .Z(n2457) );
  MUX21L U3037 ( .A(n5032), .B(n3614), .S(n3985), .Z(n2937) );
  MUX21L U3038 ( .A(n5033), .B(n3614), .S(n3984), .Z(n2873) );
  MUX21L U3039 ( .A(n5034), .B(n3614), .S(n3988), .Z(n2969) );
  MUX21L U3040 ( .A(n5035), .B(n3614), .S(n3989), .Z(n3097) );
  MUX21L U3041 ( .A(n5036), .B(n3614), .S(n4608), .Z(n3001) );
  MUX21L U3042 ( .A(n5037), .B(n3614), .S(n3990), .Z(n3065) );
  MUX21L U3043 ( .A(n5038), .B(n3614), .S(n3991), .Z(n2905) );
  MUX21L U3044 ( .A(n5039), .B(n3614), .S(n3992), .Z(n3033) );
  MUX21L U3045 ( .A(n5040), .B(n3614), .S(n3986), .Z(n3225) );
  MUX21L U3046 ( .A(n5041), .B(n3614), .S(n4615), .Z(n3289) );
  MUX21L U3047 ( .A(n5042), .B(n3614), .S(n3993), .Z(n3129) );
  MUX21L U3048 ( .A(n5043), .B(n3614), .S(n3994), .Z(n3161) );
  MUX21L U3049 ( .A(n5044), .B(n3614), .S(n3995), .Z(n3193) );
  MUX21L U3050 ( .A(n5045), .B(n3614), .S(n3987), .Z(n3321) );
  MUX21L U3051 ( .A(n5046), .B(n3614), .S(n4620), .Z(n3257) );
  AO2 U3052 ( .A(\gpr[18][6] ), .B(n4458), .C(\gpr[19][6] ), .D(n3660), .Z(
        n3620) );
  AO2 U3053 ( .A(\gpr[20][6] ), .B(n4624), .C(\gpr[16][6] ), .D(n4626), .Z(
        n3619) );
  AO2 U3054 ( .A(\gpr[21][6] ), .B(n4097), .C(\gpr[22][6] ), .D(n4431), .Z(
        n3618) );
  ND2I U3055 ( .A(\gpr[23][6] ), .B(n4548), .Z(n3616) );
  ND2I U3056 ( .A(\gpr[17][6] ), .B(n4490), .Z(n3615) );
  AN3 U3057 ( .A(n4628), .B(n3616), .C(n3615), .Z(n3617) );
  ND4 U3058 ( .A(n3620), .B(n3619), .C(n3618), .D(n3617), .Z(n3629) );
  AO2 U3059 ( .A(\gpr[26][6] ), .B(n4622), .C(\gpr[28][6] ), .D(n4624), .Z(
        n3627) );
  AO2 U3060 ( .A(\gpr[24][6] ), .B(n4497), .C(\gpr[25][6] ), .D(n4001), .Z(
        n3626) );
  AO2 U3061 ( .A(\gpr[29][6] ), .B(n4097), .C(\gpr[30][6] ), .D(n4431), .Z(
        n3625) );
  IVI U3062 ( .A(n3897), .Z(n4543) );
  AN2I U3063 ( .A(\gpr[31][6] ), .B(n4543), .Z(n3623) );
  ND2I U3064 ( .A(\gpr[27][6] ), .B(n4501), .Z(n3621) );
  ND2I U3065 ( .A(n4641), .B(n3621), .Z(n3622) );
  NR2I U3066 ( .A(n3623), .B(n3622), .Z(n3624) );
  ND4 U3067 ( .A(n3627), .B(n3626), .C(n3625), .D(n3624), .Z(n3628) );
  AN2I U3068 ( .A(n3629), .B(n3628), .Z(n3652) );
  ND2I U3069 ( .A(\gpr[1][6] ), .B(n4656), .Z(n3632) );
  ND2I U3070 ( .A(\gpr[3][6] ), .B(n4657), .Z(n3631) );
  ND2I U3071 ( .A(\gpr[5][6] ), .B(n4658), .Z(n3630) );
  ND4 U3072 ( .A(n295), .B(n3632), .C(n3631), .D(n3630), .Z(n3638) );
  ND2I U3073 ( .A(\gpr[2][6] ), .B(n4659), .Z(n3636) );
  ND2I U3074 ( .A(\gpr[10][6] ), .B(n4268), .Z(n3635) );
  ND2I U3075 ( .A(\gpr[4][6] ), .B(n4666), .Z(n3634) );
  ND2I U3076 ( .A(\gpr[9][6] ), .B(n4518), .Z(n3633) );
  ND4 U3077 ( .A(n3636), .B(n3635), .C(n3634), .D(n3633), .Z(n3637) );
  NR2I U3078 ( .A(n3638), .B(n3637), .Z(n3650) );
  IVI U3079 ( .A(n3508), .Z(n4570) );
  ND2I U3080 ( .A(\gpr[8][6] ), .B(n4570), .Z(n3642) );
  ND2I U3081 ( .A(\gpr[11][6] ), .B(n4667), .Z(n3641) );
  ND2I U3082 ( .A(\gpr[15][6] ), .B(n4572), .Z(n3640) );
  ND2I U3083 ( .A(\gpr[12][6] ), .B(n4673), .Z(n3639) );
  ND4 U3084 ( .A(n3642), .B(n3641), .C(n3640), .D(n3639), .Z(n3648) );
  ND2I U3085 ( .A(\gpr[6][6] ), .B(n4475), .Z(n3646) );
  ND2I U3086 ( .A(\gpr[13][6] ), .B(n4578), .Z(n3645) );
  ND2I U3087 ( .A(\gpr[7][6] ), .B(n4675), .Z(n3644) );
  ND2I U3088 ( .A(\gpr[14][6] ), .B(n4579), .Z(n3643) );
  ND4 U3089 ( .A(n3646), .B(n3645), .C(n3644), .D(n3643), .Z(n3647) );
  NR2I U3090 ( .A(n3648), .B(n3647), .Z(n3649) );
  ND2I U3091 ( .A(n3650), .B(n3649), .Z(n3651) );
  AN2I U3092 ( .A(n3652), .B(n3651), .Z(rd_data2[6]) );
  B4IP U3093 ( .A(wr_data[7]), .Z(n3653) );
  MUX21L U3094 ( .A(n5047), .B(n3653), .S(n3975), .Z(n2362) );
  MUX21L U3095 ( .A(n5048), .B(n3653), .S(n3981), .Z(n2426) );
  MUX21L U3096 ( .A(n5049), .B(n3653), .S(n3982), .Z(n2586) );
  MUX21L U3097 ( .A(n5050), .B(n3653), .S(n4600), .Z(n2490) );
  MUX21L U3098 ( .A(n4849), .B(n3653), .S(n3976), .Z(n2394) );
  MUX21L U3099 ( .A(n5051), .B(n3653), .S(n3977), .Z(n2522) );
  MUX21L U3100 ( .A(n5052), .B(n3653), .S(n3983), .Z(n2554) );
  MUX21L U3101 ( .A(n302), .B(n3653), .S(n3980), .Z(n2458) );
  MUX21L U3102 ( .A(n5053), .B(n3653), .S(n3996), .Z(n2682) );
  MUX21L U3103 ( .A(n303), .B(n3653), .S(n3997), .Z(n2714) );
  MUX21L U3104 ( .A(n5054), .B(n3653), .S(n4592), .Z(n2746) );
  MUX21L U3105 ( .A(n5055), .B(n3653), .S(n3999), .Z(n2810) );
  MUX21L U3106 ( .A(n4848), .B(n3653), .S(n4594), .Z(n2650) );
  MUX21L U3107 ( .A(n5056), .B(n3653), .S(n3978), .Z(n2778) );
  MUX21L U3108 ( .A(n5057), .B(n3653), .S(n3998), .Z(n2842) );
  MUX21L U3109 ( .A(n5058), .B(n3653), .S(n4597), .Z(n2618) );
  MUX21L U3110 ( .A(n5059), .B(n3653), .S(n3988), .Z(n2970) );
  MUX21L U3111 ( .A(n5060), .B(n3653), .S(n3989), .Z(n3098) );
  MUX21L U3112 ( .A(n5061), .B(n3653), .S(n4608), .Z(n3002) );
  MUX21L U3113 ( .A(n5062), .B(n3653), .S(n3990), .Z(n3066) );
  MUX21L U3114 ( .A(n4815), .B(n3653), .S(n3991), .Z(n2906) );
  MUX21L U3115 ( .A(n5063), .B(n3653), .S(n3992), .Z(n3034) );
  MUX21L U3116 ( .A(n5064), .B(n3653), .S(n3984), .Z(n2874) );
  MUX21L U3117 ( .A(n4782), .B(n3653), .S(n3985), .Z(n2938) );
  MUX21L U3118 ( .A(n5065), .B(n3653), .S(n3986), .Z(n3226) );
  MUX21L U3119 ( .A(n5066), .B(n3653), .S(n4615), .Z(n3290) );
  MUX21L U3120 ( .A(n5067), .B(n3653), .S(n3993), .Z(n3130) );
  MUX21L U3121 ( .A(n5068), .B(n3653), .S(n3994), .Z(n3162) );
  MUX21L U3122 ( .A(n5069), .B(n3653), .S(n3995), .Z(n3194) );
  MUX21L U3123 ( .A(n5070), .B(n3653), .S(n3987), .Z(n3322) );
  MUX21L U3124 ( .A(n5071), .B(n3653), .S(n4620), .Z(n3258) );
  AO2 U3125 ( .A(\gpr[26][7] ), .B(n4458), .C(\gpr[28][7] ), .D(n4624), .Z(
        n3659) );
  AO2 U3126 ( .A(\gpr[27][7] ), .B(n3660), .C(\gpr[24][7] ), .D(n4549), .Z(
        n3658) );
  AO2 U3127 ( .A(\gpr[29][7] ), .B(n4097), .C(\gpr[30][7] ), .D(n4431), .Z(
        n3657) );
  ND2I U3128 ( .A(\gpr[31][7] ), .B(n4251), .Z(n3655) );
  ND2I U3129 ( .A(\gpr[25][7] ), .B(n4490), .Z(n3654) );
  AN3 U3130 ( .A(n4641), .B(n3655), .C(n3654), .Z(n3656) );
  ND4 U3131 ( .A(n3659), .B(n3658), .C(n3657), .D(n3656), .Z(n3670) );
  AO2 U3132 ( .A(\gpr[19][7] ), .B(n3660), .C(\gpr[18][7] ), .D(n4458), .Z(
        n3668) );
  AO2 U3133 ( .A(\gpr[20][7] ), .B(n4624), .C(\gpr[17][7] ), .D(n4001), .Z(
        n3667) );
  IVI U3134 ( .A(n3785), .Z(n4413) );
  AO2 U3135 ( .A(\gpr[21][7] ), .B(n4097), .C(\gpr[23][7] ), .D(n4413), .Z(
        n3666) );
  ND2I U3136 ( .A(\gpr[22][7] ), .B(n4431), .Z(n3661) );
  IVI U3137 ( .A(n3661), .Z(n3664) );
  ND2I U3138 ( .A(\gpr[16][7] ), .B(n4432), .Z(n3662) );
  ND2I U3139 ( .A(n4628), .B(n3662), .Z(n3663) );
  NR2I U3140 ( .A(n3664), .B(n3663), .Z(n3665) );
  ND4 U3141 ( .A(n3668), .B(n3667), .C(n3666), .D(n3665), .Z(n3669) );
  AN2I U3142 ( .A(n3670), .B(n3669), .Z(n3694) );
  ND2I U3143 ( .A(n4782), .B(n3833), .Z(n3671) );
  AO3 U3144 ( .A(\gpr[15][7] ), .B(n4097), .C(n4652), .D(n3671), .Z(n3672) );
  AO3 U3145 ( .A(n4815), .B(n4655), .C(n4561), .D(n3672), .Z(n3678) );
  ND2I U3146 ( .A(\gpr[3][7] ), .B(n4657), .Z(n3676) );
  ND2I U3147 ( .A(\gpr[5][7] ), .B(n4658), .Z(n3675) );
  ND2I U3148 ( .A(\gpr[1][7] ), .B(n4656), .Z(n3674) );
  ND2I U3149 ( .A(\gpr[4][7] ), .B(n4666), .Z(n3673) );
  ND4 U3150 ( .A(n3676), .B(n3675), .C(n3674), .D(n3673), .Z(n3677) );
  NR2I U3151 ( .A(n3678), .B(n3677), .Z(n3692) );
  ND2I U3152 ( .A(\gpr[2][7] ), .B(n4659), .Z(n3684) );
  ND2I U3153 ( .A(n3679), .B(\gpr[10][7] ), .Z(n3683) );
  ND2I U3154 ( .A(\gpr[9][7] ), .B(n4668), .Z(n3682) );
  IVI U3155 ( .A(n3680), .Z(n4158) );
  IVI U3156 ( .A(n4158), .Z(n3720) );
  ND2I U3157 ( .A(\gpr[8][7] ), .B(n3720), .Z(n3681) );
  ND4 U3158 ( .A(n3684), .B(n3683), .C(n3682), .D(n3681), .Z(n3690) );
  ND2I U3159 ( .A(\gpr[11][7] ), .B(n4571), .Z(n3688) );
  ND2I U3160 ( .A(\gpr[12][7] ), .B(n4573), .Z(n3687) );
  ND2I U3161 ( .A(\gpr[7][7] ), .B(n4675), .Z(n3686) );
  ND2I U3162 ( .A(\gpr[6][7] ), .B(n4475), .Z(n3685) );
  ND4 U3163 ( .A(n3688), .B(n3687), .C(n3686), .D(n3685), .Z(n3689) );
  NR2I U3164 ( .A(n3690), .B(n3689), .Z(n3691) );
  ND2I U3165 ( .A(n3692), .B(n3691), .Z(n3693) );
  AN2I U3166 ( .A(n3694), .B(n3693), .Z(rd_data2[7]) );
  B4IP U3167 ( .A(wr_data[8]), .Z(n3695) );
  MUX21L U3168 ( .A(n5072), .B(n3695), .S(n3996), .Z(n2683) );
  MUX21L U3169 ( .A(n5073), .B(n3695), .S(n3997), .Z(n2715) );
  MUX21L U3170 ( .A(n5074), .B(n3695), .S(n4592), .Z(n2747) );
  MUX21L U3171 ( .A(n5075), .B(n3695), .S(n3999), .Z(n2811) );
  MUX21L U3172 ( .A(n4850), .B(n3695), .S(n4594), .Z(n2651) );
  MUX21L U3173 ( .A(n5076), .B(n3695), .S(n3978), .Z(n2779) );
  MUX21L U3174 ( .A(n5077), .B(n3695), .S(n3998), .Z(n2843) );
  MUX21L U3175 ( .A(n5078), .B(n3695), .S(n4597), .Z(n2619) );
  MUX21L U3176 ( .A(n4828), .B(n3695), .S(n3981), .Z(n2427) );
  MUX21L U3177 ( .A(n5079), .B(n3695), .S(n3980), .Z(n2459) );
  MUX21L U3178 ( .A(n5080), .B(n3695), .S(n3982), .Z(n2587) );
  MUX21L U3179 ( .A(n5081), .B(n3695), .S(n4600), .Z(n2491) );
  MUX21L U3180 ( .A(n5082), .B(n3695), .S(n3976), .Z(n2395) );
  MUX21L U3181 ( .A(n5083), .B(n3695), .S(n3977), .Z(n2523) );
  MUX21L U3182 ( .A(n5084), .B(n3695), .S(n3983), .Z(n2555) );
  MUX21L U3183 ( .A(n5085), .B(n3695), .S(n3975), .Z(n2363) );
  MUX21L U3184 ( .A(n5086), .B(n3695), .S(n3988), .Z(n2971) );
  MUX21L U3185 ( .A(n5087), .B(n3695), .S(n3989), .Z(n3099) );
  MUX21L U3186 ( .A(n5088), .B(n3695), .S(n4608), .Z(n3003) );
  MUX21L U3187 ( .A(n5089), .B(n3695), .S(n3990), .Z(n3067) );
  MUX21L U3188 ( .A(n4771), .B(n3695), .S(n3991), .Z(n2907) );
  MUX21L U3189 ( .A(n5090), .B(n3695), .S(n3992), .Z(n3035) );
  MUX21L U3190 ( .A(n5091), .B(n3695), .S(n3984), .Z(n2875) );
  MUX21L U3191 ( .A(n4765), .B(n3695), .S(n3985), .Z(n2939) );
  MUX21L U3192 ( .A(n5092), .B(n3695), .S(n3986), .Z(n3227) );
  MUX21L U3193 ( .A(n5093), .B(n3695), .S(n4615), .Z(n3291) );
  MUX21L U3194 ( .A(n5094), .B(n3695), .S(n3993), .Z(n3131) );
  MUX21L U3195 ( .A(n5095), .B(n3695), .S(n3994), .Z(n3163) );
  MUX21L U3196 ( .A(n5096), .B(n3695), .S(n3995), .Z(n3195) );
  MUX21L U3197 ( .A(n5097), .B(n3695), .S(n3987), .Z(n3323) );
  MUX21L U3198 ( .A(n5098), .B(n3695), .S(n4620), .Z(n3259) );
  AO2 U3199 ( .A(\gpr[19][8] ), .B(n4009), .C(\gpr[18][8] ), .D(n4293), .Z(
        n3702) );
  AO2 U3200 ( .A(\gpr[17][8] ), .B(n4001), .C(\gpr[20][8] ), .D(n4498), .Z(
        n3701) );
  IVI U3201 ( .A(n3778), .Z(n4342) );
  AO2 U3202 ( .A(\gpr[21][8] ), .B(n4097), .C(\gpr[23][8] ), .D(n4342), .Z(
        n3700) );
  AN2I U3203 ( .A(\gpr[22][8] ), .B(n4431), .Z(n3698) );
  ND2I U3204 ( .A(\gpr[16][8] ), .B(n4549), .Z(n3696) );
  ND2I U3205 ( .A(n4628), .B(n3696), .Z(n3697) );
  NR2I U3206 ( .A(n3698), .B(n3697), .Z(n3699) );
  ND4 U3207 ( .A(n3702), .B(n3701), .C(n3700), .D(n3699), .Z(n3711) );
  AO2 U3208 ( .A(\gpr[26][8] ), .B(n3703), .C(\gpr[24][8] ), .D(n4497), .Z(
        n3709) );
  AO2 U3209 ( .A(\gpr[27][8] ), .B(n4009), .C(\gpr[28][8] ), .D(n4624), .Z(
        n3708) );
  AO2 U3210 ( .A(\gpr[31][8] ), .B(n3864), .C(\gpr[29][8] ), .D(n4097), .Z(
        n3707) );
  ND2I U3211 ( .A(\gpr[30][8] ), .B(n4625), .Z(n3705) );
  ND2I U3212 ( .A(\gpr[25][8] ), .B(n4490), .Z(n3704) );
  AN3 U3213 ( .A(n4641), .B(n3705), .C(n3704), .Z(n3706) );
  ND4 U3214 ( .A(n3709), .B(n3708), .C(n3707), .D(n3706), .Z(n3710) );
  AN2I U3215 ( .A(n3711), .B(n3710), .Z(n3734) );
  ND2I U3216 ( .A(n4765), .B(n3833), .Z(n3712) );
  AO3 U3217 ( .A(\gpr[15][8] ), .B(n4097), .C(n4652), .D(n3712), .Z(n3713) );
  AO3 U3218 ( .A(n4771), .B(n4466), .C(n295), .D(n3713), .Z(n3719) );
  ND2I U3219 ( .A(\gpr[3][8] ), .B(n4657), .Z(n3717) );
  ND2I U3220 ( .A(\gpr[5][8] ), .B(n4658), .Z(n3716) );
  ND2I U3221 ( .A(\gpr[1][8] ), .B(n4656), .Z(n3715) );
  ND2I U3222 ( .A(\gpr[4][8] ), .B(n4153), .Z(n3714) );
  ND4 U3223 ( .A(n3717), .B(n3716), .C(n3715), .D(n3714), .Z(n3718) );
  NR2I U3224 ( .A(n3719), .B(n3718), .Z(n3732) );
  ND2I U3225 ( .A(\gpr[2][8] ), .B(n4659), .Z(n3724) );
  ND2I U3226 ( .A(\gpr[10][8] ), .B(n4268), .Z(n3723) );
  ND2I U3227 ( .A(\gpr[9][8] ), .B(n4314), .Z(n3722) );
  ND2I U3228 ( .A(\gpr[8][8] ), .B(n3720), .Z(n3721) );
  ND4 U3229 ( .A(n3724), .B(n3723), .C(n3722), .D(n3721), .Z(n3730) );
  ND2I U3230 ( .A(\gpr[11][8] ), .B(n4571), .Z(n3728) );
  ND2I U3231 ( .A(\gpr[12][8] ), .B(n4573), .Z(n3727) );
  ND2I U3232 ( .A(\gpr[7][8] ), .B(n4675), .Z(n3726) );
  ND2I U3233 ( .A(\gpr[6][8] ), .B(n4354), .Z(n3725) );
  ND4 U3234 ( .A(n3728), .B(n3727), .C(n3726), .D(n3725), .Z(n3729) );
  NR2I U3235 ( .A(n3730), .B(n3729), .Z(n3731) );
  ND2I U3236 ( .A(n3732), .B(n3731), .Z(n3733) );
  AN2I U3237 ( .A(n3734), .B(n3733), .Z(rd_data2[8]) );
  B4IP U3238 ( .A(wr_data[9]), .Z(n3735) );
  MUX21L U3239 ( .A(n5099), .B(n3735), .S(n3975), .Z(n2364) );
  MUX21L U3240 ( .A(n5100), .B(n3735), .S(n3981), .Z(n2428) );
  MUX21L U3241 ( .A(n5101), .B(n3735), .S(n3982), .Z(n2588) );
  MUX21L U3242 ( .A(n5102), .B(n3735), .S(n3983), .Z(n2556) );
  MUX21L U3243 ( .A(n4851), .B(n3735), .S(n3976), .Z(n2396) );
  MUX21L U3244 ( .A(n5103), .B(n3735), .S(n3977), .Z(n2524) );
  MUX21L U3245 ( .A(n5104), .B(n3735), .S(n4600), .Z(n2492) );
  MUX21L U3246 ( .A(n5105), .B(n3735), .S(n3980), .Z(n2460) );
  MUX21L U3247 ( .A(n5106), .B(n3735), .S(n4597), .Z(n2620) );
  MUX21L U3248 ( .A(n5107), .B(n3735), .S(n3996), .Z(n2684) );
  MUX21L U3249 ( .A(n5108), .B(n3735), .S(n3998), .Z(n2844) );
  MUX21L U3250 ( .A(n5109), .B(n3735), .S(n3999), .Z(n2812) );
  MUX21L U3251 ( .A(n4852), .B(n3735), .S(n4594), .Z(n2652) );
  MUX21L U3252 ( .A(n5110), .B(n3735), .S(n3978), .Z(n2780) );
  MUX21L U3253 ( .A(n5111), .B(n3735), .S(n4592), .Z(n2748) );
  MUX21L U3254 ( .A(n5112), .B(n3735), .S(n3997), .Z(n2716) );
  MUX21L U3255 ( .A(n5113), .B(n3735), .S(n3988), .Z(n2972) );
  MUX21L U3256 ( .A(n5114), .B(n3735), .S(n3989), .Z(n3100) );
  MUX21L U3257 ( .A(n5115), .B(n3735), .S(n4608), .Z(n3004) );
  MUX21L U3258 ( .A(n5116), .B(n3735), .S(n3990), .Z(n3068) );
  MUX21L U3259 ( .A(n4816), .B(n3735), .S(n3991), .Z(n2908) );
  MUX21L U3260 ( .A(n5117), .B(n3735), .S(n3992), .Z(n3036) );
  MUX21L U3261 ( .A(n5118), .B(n3735), .S(n3984), .Z(n2876) );
  MUX21L U3262 ( .A(n4783), .B(n3735), .S(n3985), .Z(n2940) );
  MUX21L U3263 ( .A(n5119), .B(n3735), .S(n3986), .Z(n3228) );
  MUX21L U3264 ( .A(n5120), .B(n3735), .S(n4615), .Z(n3292) );
  MUX21L U3265 ( .A(n5121), .B(n3735), .S(n3993), .Z(n3132) );
  MUX21L U3266 ( .A(n5122), .B(n3735), .S(n3994), .Z(n3164) );
  MUX21L U3267 ( .A(n5123), .B(n3735), .S(n3995), .Z(n3196) );
  MUX21L U3268 ( .A(n5124), .B(n3735), .S(n3987), .Z(n3324) );
  MUX21L U3269 ( .A(n5125), .B(n3735), .S(n4620), .Z(n3260) );
  AO2 U3270 ( .A(\gpr[26][9] ), .B(n4458), .C(\gpr[28][9] ), .D(n4624), .Z(
        n3742) );
  AO2 U3271 ( .A(\gpr[25][9] ), .B(n4636), .C(\gpr[24][9] ), .D(n4357), .Z(
        n3741) );
  AO2 U3272 ( .A(\gpr[29][9] ), .B(n4097), .C(\gpr[30][9] ), .D(n4431), .Z(
        n3740) );
  AN2I U3273 ( .A(\gpr[31][9] ), .B(n4209), .Z(n3738) );
  ND2I U3274 ( .A(\gpr[27][9] ), .B(n4501), .Z(n3736) );
  ND2I U3275 ( .A(n4641), .B(n3736), .Z(n3737) );
  NR2I U3276 ( .A(n3738), .B(n3737), .Z(n3739) );
  ND4 U3277 ( .A(n3742), .B(n3741), .C(n3740), .D(n3739), .Z(n3748) );
  AO2 U3278 ( .A(\gpr[18][9] ), .B(n4622), .C(\gpr[20][9] ), .D(n4624), .Z(
        n3746) );
  AO2 U3279 ( .A(\gpr[17][9] ), .B(n4001), .C(\gpr[16][9] ), .D(n4549), .Z(
        n3745) );
  AO2 U3280 ( .A(\gpr[21][9] ), .B(n4097), .C(\gpr[22][9] ), .D(n4431), .Z(
        n3744) );
  IVI U3281 ( .A(n4054), .Z(n4623) );
  ND4 U3282 ( .A(n3746), .B(n3745), .C(n3744), .D(n3743), .Z(n3747) );
  AN2I U3283 ( .A(n3748), .B(n3747), .Z(n3770) );
  ND2I U3284 ( .A(n4783), .B(n3833), .Z(n3749) );
  AO3 U3285 ( .A(\gpr[15][9] ), .B(n4097), .C(n4652), .D(n3749), .Z(n3750) );
  AO3 U3286 ( .A(n4816), .B(n4655), .C(n295), .D(n3750), .Z(n3756) );
  ND2I U3287 ( .A(\gpr[3][9] ), .B(n4657), .Z(n3754) );
  ND2I U3288 ( .A(\gpr[5][9] ), .B(n4658), .Z(n3753) );
  ND2I U3289 ( .A(\gpr[1][9] ), .B(n4656), .Z(n3752) );
  ND2I U3290 ( .A(\gpr[4][9] ), .B(n4666), .Z(n3751) );
  ND4 U3291 ( .A(n3754), .B(n3753), .C(n3752), .D(n3751), .Z(n3755) );
  NR2I U3292 ( .A(n3756), .B(n3755), .Z(n3768) );
  ND2I U3293 ( .A(\gpr[2][9] ), .B(n4659), .Z(n3760) );
  ND2I U3294 ( .A(n3679), .B(\gpr[10][9] ), .Z(n3759) );
  ND2I U3295 ( .A(\gpr[9][9] ), .B(n4563), .Z(n3758) );
  IVI U3296 ( .A(n3561), .Z(n3960) );
  ND2I U3297 ( .A(\gpr[8][9] ), .B(n3960), .Z(n3757) );
  ND4 U3298 ( .A(n3760), .B(n3759), .C(n3758), .D(n3757), .Z(n3766) );
  ND2I U3299 ( .A(\gpr[11][9] ), .B(n4667), .Z(n3764) );
  ND2I U3300 ( .A(\gpr[12][9] ), .B(n4673), .Z(n3763) );
  ND2I U3301 ( .A(\gpr[7][9] ), .B(n4675), .Z(n3762) );
  ND2I U3302 ( .A(\gpr[6][9] ), .B(n4197), .Z(n3761) );
  ND4 U3303 ( .A(n3764), .B(n3763), .C(n3762), .D(n3761), .Z(n3765) );
  NR2I U3304 ( .A(n3766), .B(n3765), .Z(n3767) );
  ND2I U3305 ( .A(n3768), .B(n3767), .Z(n3769) );
  AN2I U3306 ( .A(n3770), .B(n3769), .Z(rd_data2[9]) );
  B4IP U3307 ( .A(wr_data[10]), .Z(n3775) );
  B5IP U3308 ( .A(n3771), .Z(n4605) );
  MUX21L U3309 ( .A(n5126), .B(n3775), .S(n4605), .Z(n2365) );
  MUX21L U3310 ( .A(n5127), .B(n3775), .S(n3980), .Z(n2461) );
  MUX21L U3311 ( .A(n5128), .B(n3775), .S(n3982), .Z(n2589) );
  MUX21L U3312 ( .A(n5129), .B(n3775), .S(n3983), .Z(n2557) );
  B5IP U3313 ( .A(n3772), .Z(n4602) );
  MUX21L U3314 ( .A(n5130), .B(n3775), .S(n4602), .Z(n2397) );
  B5IP U3315 ( .A(n3773), .Z(n4603) );
  MUX21L U3316 ( .A(n5131), .B(n3775), .S(n4603), .Z(n2525) );
  MUX21L U3317 ( .A(n5132), .B(n3775), .S(n4600), .Z(n2493) );
  MUX21L U3318 ( .A(n4829), .B(n3775), .S(n3981), .Z(n2429) );
  MUX21L U3319 ( .A(n4853), .B(n3775), .S(n4597), .Z(n2621) );
  MUX21L U3320 ( .A(n5133), .B(n3775), .S(n3996), .Z(n2685) );
  MUX21L U3321 ( .A(n5134), .B(n3775), .S(n3997), .Z(n2717) );
  MUX21L U3322 ( .A(n5135), .B(n3775), .S(n3999), .Z(n2813) );
  MUX21L U3323 ( .A(n5136), .B(n3775), .S(n4594), .Z(n2653) );
  B5IP U3324 ( .A(n3774), .Z(n4595) );
  MUX21L U3325 ( .A(n5137), .B(n3775), .S(n4595), .Z(n2781) );
  MUX21L U3326 ( .A(n5138), .B(n3775), .S(n3998), .Z(n2845) );
  MUX21L U3327 ( .A(n5139), .B(n3775), .S(n4592), .Z(n2749) );
  MUX21L U3328 ( .A(n5140), .B(n3775), .S(n3985), .Z(n2941) );
  MUX21L U3329 ( .A(n5141), .B(n3775), .S(n3984), .Z(n2877) );
  MUX21L U3330 ( .A(n5142), .B(n3775), .S(n3988), .Z(n2973) );
  MUX21L U3331 ( .A(n5143), .B(n3775), .S(n3989), .Z(n3101) );
  MUX21L U3332 ( .A(n5144), .B(n3775), .S(n4608), .Z(n3005) );
  MUX21L U3333 ( .A(n5145), .B(n3775), .S(n3990), .Z(n3069) );
  MUX21L U3334 ( .A(n5146), .B(n3775), .S(n3991), .Z(n2909) );
  MUX21L U3335 ( .A(n5147), .B(n3775), .S(n3992), .Z(n3037) );
  MUX21L U3336 ( .A(n5148), .B(n3775), .S(n3986), .Z(n3229) );
  MUX21L U3337 ( .A(n5149), .B(n3775), .S(n4615), .Z(n3293) );
  MUX21L U3338 ( .A(n5150), .B(n3775), .S(n3993), .Z(n3133) );
  MUX21L U3339 ( .A(n5151), .B(n3775), .S(n3994), .Z(n3165) );
  MUX21L U3340 ( .A(n5152), .B(n3775), .S(n3995), .Z(n3197) );
  MUX21L U3341 ( .A(n5153), .B(n3775), .S(n3987), .Z(n3325) );
  MUX21L U3342 ( .A(n5154), .B(n3775), .S(n4620), .Z(n3261) );
  B5IP U3343 ( .A(wr_data[11]), .Z(n3777) );
  MUX21L U3344 ( .A(n5155), .B(n3777), .S(n4597), .Z(n2622) );
  MUX21L U3345 ( .A(n5156), .B(n3777), .S(n3996), .Z(n2686) );
  MUX21L U3346 ( .A(n5157), .B(n3777), .S(n3998), .Z(n2846) );
  MUX21L U3347 ( .A(n5158), .B(n3777), .S(n4592), .Z(n2750) );
  MUX21L U3348 ( .A(n4854), .B(n3777), .S(n4594), .Z(n2654) );
  MUX21L U3349 ( .A(n5159), .B(n3777), .S(n3978), .Z(n2782) );
  MUX21L U3350 ( .A(n5160), .B(n3777), .S(n3999), .Z(n2814) );
  MUX21L U3351 ( .A(n5161), .B(n3777), .S(n3997), .Z(n2718) );
  MUX21L U3352 ( .A(n5162), .B(n3777), .S(n3981), .Z(n2430) );
  IVI U3353 ( .A(\gpr[28][11] ), .Z(n3776) );
  MUX21L U3354 ( .A(n3776), .B(n3777), .S(n3980), .Z(n2462) );
  MUX21L U3355 ( .A(n5163), .B(n3777), .S(n3982), .Z(n2590) );
  MUX21L U3356 ( .A(n5164), .B(n3777), .S(n4600), .Z(n2494) );
  MUX21L U3357 ( .A(n4855), .B(n3777), .S(n3976), .Z(n2398) );
  MUX21L U3358 ( .A(n5165), .B(n3777), .S(n3977), .Z(n2526) );
  MUX21L U3359 ( .A(n5166), .B(n3777), .S(n3983), .Z(n2558) );
  MUX21L U3360 ( .A(n5167), .B(n3777), .S(n3975), .Z(n2366) );
  MUX21L U3361 ( .A(n5168), .B(n3777), .S(n3988), .Z(n2974) );
  MUX21L U3362 ( .A(n5169), .B(n3777), .S(n3989), .Z(n3102) );
  MUX21L U3363 ( .A(n5170), .B(n3777), .S(n4608), .Z(n3006) );
  MUX21L U3364 ( .A(n5171), .B(n3777), .S(n3990), .Z(n3070) );
  MUX21L U3365 ( .A(n5172), .B(n3777), .S(n3991), .Z(n2910) );
  MUX21L U3366 ( .A(n5173), .B(n3777), .S(n3992), .Z(n3038) );
  MUX21L U3367 ( .A(n5174), .B(n3777), .S(n3984), .Z(n2878) );
  MUX21L U3368 ( .A(n4784), .B(n3777), .S(n3985), .Z(n2942) );
  MUX21L U3369 ( .A(n5175), .B(n3777), .S(n3986), .Z(n3230) );
  MUX21L U3370 ( .A(n5176), .B(n3777), .S(n4615), .Z(n3294) );
  MUX21L U3371 ( .A(n5177), .B(n3777), .S(n3993), .Z(n3134) );
  MUX21L U3372 ( .A(n5692), .B(n3777), .S(n3994), .Z(n3166) );
  MUX21L U3373 ( .A(n4761), .B(n3777), .S(n3995), .Z(n3198) );
  MUX21L U3374 ( .A(n5693), .B(n3777), .S(n3987), .Z(n3326) );
  MUX21L U3375 ( .A(n5694), .B(n3777), .S(n4620), .Z(n3262) );
  AO2 U3376 ( .A(\gpr[18][11] ), .B(n4487), .C(\gpr[20][11] ), .D(n4498), .Z(
        n3784) );
  AO2 U3377 ( .A(\gpr[19][11] ), .B(n4009), .C(\gpr[16][11] ), .D(n4450), .Z(
        n3783) );
  AO2 U3378 ( .A(\gpr[21][11] ), .B(n4090), .C(\gpr[22][11] ), .D(n4431), .Z(
        n3782) );
  IVI U3379 ( .A(n3778), .Z(n4333) );
  ND2I U3380 ( .A(\gpr[23][11] ), .B(n4333), .Z(n3780) );
  ND2I U3381 ( .A(\gpr[17][11] ), .B(n4490), .Z(n3779) );
  AN3 U3382 ( .A(n4628), .B(n3780), .C(n3779), .Z(n3781) );
  ND4 U3383 ( .A(n3784), .B(n3783), .C(n3782), .D(n3781), .Z(n3793) );
  AO2 U3384 ( .A(\gpr[26][11] ), .B(n4622), .C(\gpr[24][11] ), .D(n4637), .Z(
        n3791) );
  AO2 U3385 ( .A(\gpr[27][11] ), .B(n4009), .C(\gpr[28][11] ), .D(n4624), .Z(
        n3790) );
  IVI U3386 ( .A(n3785), .Z(n4488) );
  AO2 U3387 ( .A(\gpr[29][11] ), .B(n4090), .C(\gpr[31][11] ), .D(n4488), .Z(
        n3789) );
  ND2I U3388 ( .A(\gpr[30][11] ), .B(n4625), .Z(n3787) );
  ND2I U3389 ( .A(\gpr[25][11] ), .B(n4490), .Z(n3786) );
  AN3 U3390 ( .A(n4641), .B(n3787), .C(n3786), .Z(n3788) );
  ND4 U3391 ( .A(n3791), .B(n3790), .C(n3789), .D(n3788), .Z(n3792) );
  AN2I U3392 ( .A(n3793), .B(n3792), .Z(n3815) );
  ND2I U3393 ( .A(\gpr[6][11] ), .B(n4197), .Z(n3796) );
  ND2I U3394 ( .A(n4784), .B(n3833), .Z(n3794) );
  AO3 U3395 ( .A(\gpr[15][11] ), .B(n4090), .C(n4652), .D(n3794), .Z(n3795) );
  AN3 U3396 ( .A(n4561), .B(n3796), .C(n3795), .Z(n3813) );
  AO2 U3397 ( .A(\gpr[2][11] ), .B(n4659), .C(\gpr[7][11] ), .D(n4675), .Z(
        n3812) );
  AO2 U3398 ( .A(\gpr[1][11] ), .B(n4656), .C(\gpr[3][11] ), .D(n4657), .Z(
        n3800) );
  ND2I U3399 ( .A(\gpr[4][11] ), .B(n4153), .Z(n3798) );
  ND2I U3400 ( .A(n4658), .B(\gpr[5][11] ), .Z(n3797) );
  AN2I U3401 ( .A(n3798), .B(n3797), .Z(n3799) );
  AN2I U3402 ( .A(n3800), .B(n3799), .Z(n3811) );
  AO2 U3403 ( .A(\gpr[8][11] ), .B(n4637), .C(\gpr[14][11] ), .D(n4431), .Z(
        n3808) );
  ND2I U3404 ( .A(\gpr[10][11] ), .B(n4487), .Z(n3802) );
  ND2I U3405 ( .A(\gpr[9][11] ), .B(n4490), .Z(n3801) );
  ND2I U3406 ( .A(n3802), .B(n3801), .Z(n3806) );
  ND2I U3407 ( .A(\gpr[11][11] ), .B(n4623), .Z(n3804) );
  ND2I U3408 ( .A(\gpr[12][11] ), .B(n219), .Z(n3803) );
  ND2I U3409 ( .A(n3804), .B(n3803), .Z(n3805) );
  NR2I U3410 ( .A(n3806), .B(n3805), .Z(n3807) );
  ND2I U3411 ( .A(n3808), .B(n3807), .Z(n3809) );
  ND2I U3412 ( .A(n4442), .B(n3809), .Z(n3810) );
  ND4 U3413 ( .A(n3813), .B(n3812), .C(n3811), .D(n3810), .Z(n3814) );
  AN2I U3414 ( .A(n3815), .B(n3814), .Z(rd_data2[11]) );
  B4IP U3415 ( .A(wr_data[12]), .Z(n3816) );
  MUX21L U3416 ( .A(n5178), .B(n3816), .S(n3981), .Z(n2431) );
  MUX21L U3417 ( .A(n5179), .B(n3816), .S(n3980), .Z(n2463) );
  MUX21L U3418 ( .A(n5180), .B(n3816), .S(n4600), .Z(n2495) );
  MUX21L U3419 ( .A(n5181), .B(n3816), .S(n3983), .Z(n2559) );
  MUX21L U3420 ( .A(n4857), .B(n3816), .S(n4602), .Z(n2399) );
  MUX21L U3421 ( .A(n5182), .B(n3816), .S(n4603), .Z(n2527) );
  MUX21L U3422 ( .A(n5183), .B(n3816), .S(n3982), .Z(n2591) );
  MUX21L U3423 ( .A(n5184), .B(n3816), .S(n4605), .Z(n2367) );
  MUX21L U3424 ( .A(n5185), .B(n3816), .S(n3996), .Z(n2687) );
  MUX21L U3425 ( .A(n5186), .B(n3816), .S(n3997), .Z(n2719) );
  MUX21L U3426 ( .A(n5187), .B(n3816), .S(n3998), .Z(n2847) );
  MUX21L U3427 ( .A(n5188), .B(n3816), .S(n4592), .Z(n2751) );
  MUX21L U3428 ( .A(n4856), .B(n3816), .S(n4594), .Z(n2655) );
  MUX21L U3429 ( .A(n5189), .B(n3816), .S(n4595), .Z(n2783) );
  MUX21L U3430 ( .A(n5190), .B(n3816), .S(n3999), .Z(n2815) );
  MUX21L U3431 ( .A(n5191), .B(n3816), .S(n4597), .Z(n2623) );
  MUX21L U3432 ( .A(n5192), .B(n3816), .S(n3988), .Z(n2975) );
  MUX21L U3433 ( .A(n5193), .B(n3816), .S(n3989), .Z(n3103) );
  MUX21L U3434 ( .A(n5695), .B(n3816), .S(n4608), .Z(n3007) );
  MUX21L U3435 ( .A(n5696), .B(n3816), .S(n3990), .Z(n3071) );
  MUX21L U3436 ( .A(n4817), .B(n3816), .S(n3991), .Z(n2911) );
  MUX21L U3437 ( .A(n5194), .B(n3816), .S(n3992), .Z(n3039) );
  MUX21L U3438 ( .A(n5195), .B(n3816), .S(n3984), .Z(n2879) );
  MUX21L U3439 ( .A(n4785), .B(n3816), .S(n3985), .Z(n2943) );
  MUX21L U3440 ( .A(n5196), .B(n3816), .S(n3986), .Z(n3231) );
  MUX21L U3441 ( .A(n5197), .B(n3816), .S(n4615), .Z(n3295) );
  MUX21L U3442 ( .A(n5697), .B(n3816), .S(n3993), .Z(n3135) );
  MUX21L U3443 ( .A(n5698), .B(n3816), .S(n3994), .Z(n3167) );
  MUX21L U3444 ( .A(n5699), .B(n3816), .S(n3995), .Z(n3199) );
  MUX21L U3445 ( .A(n5700), .B(n3816), .S(n3987), .Z(n3327) );
  MUX21L U3446 ( .A(n5701), .B(n3816), .S(n4620), .Z(n3263) );
  AO2 U3447 ( .A(\gpr[26][12] ), .B(n4214), .C(\gpr[27][12] ), .D(n4009), .Z(
        n3824) );
  AO2 U3448 ( .A(\gpr[25][12] ), .B(n4001), .C(\gpr[28][12] ), .D(n4498), .Z(
        n3823) );
  AO2 U3449 ( .A(\gpr[29][12] ), .B(n4090), .C(\gpr[31][12] ), .D(n4413), .Z(
        n3822) );
  ND2I U3450 ( .A(\gpr[30][12] ), .B(n4431), .Z(n3817) );
  IVI U3451 ( .A(n3817), .Z(n3820) );
  ND2I U3452 ( .A(\gpr[24][12] ), .B(n4637), .Z(n3818) );
  ND2I U3453 ( .A(n4641), .B(n3818), .Z(n3819) );
  NR2I U3454 ( .A(n3820), .B(n3819), .Z(n3821) );
  ND4 U3455 ( .A(n3824), .B(n3823), .C(n3822), .D(n3821), .Z(n3832) );
  AO2 U3456 ( .A(\gpr[18][12] ), .B(n4214), .C(\gpr[16][12] ), .D(n4432), .Z(
        n3830) );
  AO2 U3457 ( .A(\gpr[19][12] ), .B(n4009), .C(\gpr[20][12] ), .D(n4624), .Z(
        n3829) );
  AO2 U3458 ( .A(\gpr[21][12] ), .B(n4090), .C(\gpr[23][12] ), .D(n4002), .Z(
        n3828) );
  ND2I U3459 ( .A(\gpr[22][12] ), .B(n4431), .Z(n3826) );
  ND2I U3460 ( .A(\gpr[17][12] ), .B(n4490), .Z(n3825) );
  AN3 U3461 ( .A(n4628), .B(n3826), .C(n3825), .Z(n3827) );
  ND4 U3462 ( .A(n3830), .B(n3829), .C(n3828), .D(n3827), .Z(n3831) );
  AN2I U3463 ( .A(n3832), .B(n3831), .Z(n3855) );
  ND2I U3464 ( .A(n4785), .B(n3833), .Z(n3834) );
  AO3 U3465 ( .A(\gpr[15][12] ), .B(n4090), .C(n4652), .D(n3834), .Z(n3835) );
  AO3 U3466 ( .A(n4817), .B(n3953), .C(n295), .D(n3835), .Z(n3841) );
  ND2I U3467 ( .A(\gpr[3][12] ), .B(n4657), .Z(n3839) );
  ND2I U3468 ( .A(\gpr[5][12] ), .B(n4658), .Z(n3838) );
  ND2I U3469 ( .A(\gpr[1][12] ), .B(n4656), .Z(n3837) );
  ND2I U3470 ( .A(\gpr[4][12] ), .B(n4153), .Z(n3836) );
  ND4 U3471 ( .A(n3839), .B(n3838), .C(n3837), .D(n3836), .Z(n3840) );
  NR2I U3472 ( .A(n3841), .B(n3840), .Z(n3853) );
  ND2I U3473 ( .A(\gpr[2][12] ), .B(n4659), .Z(n3845) );
  ND2I U3474 ( .A(n4473), .B(\gpr[10][12] ), .Z(n3844) );
  ND2I U3475 ( .A(\gpr[9][12] ), .B(n4314), .Z(n3843) );
  ND2I U3476 ( .A(\gpr[8][12] ), .B(n4570), .Z(n3842) );
  ND4 U3477 ( .A(n3845), .B(n3844), .C(n3843), .D(n3842), .Z(n3851) );
  ND2I U3478 ( .A(\gpr[11][12] ), .B(n4667), .Z(n3849) );
  ND2I U3479 ( .A(\gpr[12][12] ), .B(n4673), .Z(n3848) );
  ND2I U3480 ( .A(\gpr[7][12] ), .B(n4675), .Z(n3847) );
  ND2I U3481 ( .A(\gpr[6][12] ), .B(n4475), .Z(n3846) );
  ND4 U3482 ( .A(n3849), .B(n3848), .C(n3847), .D(n3846), .Z(n3850) );
  NR2I U3483 ( .A(n3851), .B(n3850), .Z(n3852) );
  ND2I U3484 ( .A(n3853), .B(n3852), .Z(n3854) );
  AN2I U3485 ( .A(n3855), .B(n3854), .Z(rd_data2[12]) );
  B4IP U3486 ( .A(wr_data[13]), .Z(n3856) );
  MUX21L U3487 ( .A(n5198), .B(n3856), .S(n4605), .Z(n2368) );
  MUX21L U3488 ( .A(n5199), .B(n3856), .S(n3981), .Z(n2432) );
  MUX21L U3489 ( .A(n5200), .B(n3856), .S(n3982), .Z(n2592) );
  MUX21L U3490 ( .A(n5201), .B(n3856), .S(n3983), .Z(n2560) );
  MUX21L U3491 ( .A(n4859), .B(n3856), .S(n4602), .Z(n2400) );
  MUX21L U3492 ( .A(n5202), .B(n3856), .S(n4603), .Z(n2528) );
  MUX21L U3493 ( .A(n5203), .B(n3856), .S(n4600), .Z(n2496) );
  MUX21L U3494 ( .A(n5204), .B(n3856), .S(n3980), .Z(n2464) );
  MUX21L U3495 ( .A(n4858), .B(n3856), .S(n4597), .Z(n2624) );
  MUX21L U3496 ( .A(n5205), .B(n3856), .S(n3996), .Z(n2688) );
  MUX21L U3497 ( .A(n5206), .B(n3856), .S(n3997), .Z(n2720) );
  MUX21L U3498 ( .A(n5207), .B(n3856), .S(n3998), .Z(n2848) );
  MUX21L U3499 ( .A(n5208), .B(n3856), .S(n4594), .Z(n2656) );
  MUX21L U3500 ( .A(n5209), .B(n3856), .S(n4595), .Z(n2784) );
  MUX21L U3501 ( .A(n5210), .B(n3856), .S(n3999), .Z(n2816) );
  MUX21L U3502 ( .A(n5211), .B(n3856), .S(n4592), .Z(n2752) );
  MUX21L U3503 ( .A(n5212), .B(n3856), .S(n3988), .Z(n2976) );
  MUX21L U3504 ( .A(n5213), .B(n3856), .S(n3989), .Z(n3104) );
  MUX21L U3505 ( .A(n5214), .B(n3856), .S(n4608), .Z(n3008) );
  MUX21L U3506 ( .A(n5215), .B(n3856), .S(n3990), .Z(n3072) );
  MUX21L U3507 ( .A(n4818), .B(n3856), .S(n3991), .Z(n2912) );
  MUX21L U3508 ( .A(n5216), .B(n3856), .S(n3992), .Z(n3040) );
  MUX21L U3509 ( .A(n5217), .B(n3856), .S(n3984), .Z(n2880) );
  MUX21L U3510 ( .A(n4786), .B(n3856), .S(n3985), .Z(n2944) );
  MUX21L U3511 ( .A(n5218), .B(n3856), .S(n3986), .Z(n3232) );
  MUX21L U3512 ( .A(n5219), .B(n3856), .S(n4615), .Z(n3296) );
  MUX21L U3513 ( .A(n5220), .B(n3856), .S(n3993), .Z(n3136) );
  MUX21L U3514 ( .A(n5221), .B(n3856), .S(n3994), .Z(n3168) );
  MUX21L U3515 ( .A(n5222), .B(n3856), .S(n3995), .Z(n3200) );
  MUX21L U3516 ( .A(n5223), .B(n3856), .S(n3987), .Z(n3328) );
  MUX21L U3517 ( .A(n5224), .B(n3856), .S(n4620), .Z(n3264) );
  AO2 U3518 ( .A(\gpr[28][13] ), .B(n4624), .C(\gpr[26][13] ), .D(n4487), .Z(
        n3863) );
  AO2 U3519 ( .A(\gpr[24][13] ), .B(n4497), .C(\gpr[25][13] ), .D(n4001), .Z(
        n3862) );
  AO2 U3520 ( .A(\gpr[29][13] ), .B(n4090), .C(\gpr[30][13] ), .D(n4431), .Z(
        n3861) );
  AN2I U3521 ( .A(\gpr[31][13] ), .B(n4374), .Z(n3859) );
  ND2I U3522 ( .A(\gpr[27][13] ), .B(n4623), .Z(n3857) );
  ND2I U3523 ( .A(n4453), .B(n3857), .Z(n3858) );
  NR2I U3524 ( .A(n3859), .B(n3858), .Z(n3860) );
  ND4 U3525 ( .A(n3863), .B(n3862), .C(n3861), .D(n3860), .Z(n3872) );
  AO2 U3526 ( .A(\gpr[19][13] ), .B(n4009), .C(\gpr[18][13] ), .D(n4458), .Z(
        n3870) );
  AO2 U3527 ( .A(\gpr[16][13] ), .B(n4542), .C(\gpr[20][13] ), .D(n219), .Z(
        n3869) );
  AO2 U3528 ( .A(\gpr[21][13] ), .B(n4090), .C(\gpr[22][13] ), .D(n4431), .Z(
        n3868) );
  ND2I U3529 ( .A(\gpr[23][13] ), .B(n3864), .Z(n3866) );
  ND2I U3530 ( .A(\gpr[17][13] ), .B(n4490), .Z(n3865) );
  AN3 U3531 ( .A(n4628), .B(n3866), .C(n3865), .Z(n3867) );
  ND4 U3532 ( .A(n3870), .B(n3869), .C(n3868), .D(n3867), .Z(n3871) );
  AN2I U3533 ( .A(n3872), .B(n3871), .Z(n3895) );
  IVI U3534 ( .A(n3873), .Z(n4108) );
  ND2I U3535 ( .A(n4786), .B(n4184), .Z(n3874) );
  AO3 U3536 ( .A(\gpr[15][13] ), .B(n4090), .C(n4652), .D(n3874), .Z(n3875) );
  AO3 U3537 ( .A(n4818), .B(n4108), .C(n295), .D(n3875), .Z(n3881) );
  ND2I U3538 ( .A(\gpr[3][13] ), .B(n4657), .Z(n3879) );
  ND2I U3539 ( .A(\gpr[5][13] ), .B(n4658), .Z(n3878) );
  ND2I U3540 ( .A(\gpr[1][13] ), .B(n4656), .Z(n3877) );
  ND2I U3541 ( .A(\gpr[4][13] ), .B(n4666), .Z(n3876) );
  ND4 U3542 ( .A(n3879), .B(n3878), .C(n3877), .D(n3876), .Z(n3880) );
  NR2I U3543 ( .A(n3881), .B(n3880), .Z(n3893) );
  ND2I U3544 ( .A(\gpr[2][13] ), .B(n4659), .Z(n3885) );
  ND2I U3545 ( .A(\gpr[10][13] ), .B(n4268), .Z(n3884) );
  ND2I U3546 ( .A(\gpr[9][13] ), .B(n4518), .Z(n3883) );
  ND2I U3547 ( .A(\gpr[8][13] ), .B(n4519), .Z(n3882) );
  ND4 U3548 ( .A(n3885), .B(n3884), .C(n3883), .D(n3882), .Z(n3891) );
  ND2I U3549 ( .A(\gpr[11][13] ), .B(n4571), .Z(n3889) );
  ND2I U3550 ( .A(\gpr[12][13] ), .B(n4573), .Z(n3888) );
  ND2I U3551 ( .A(\gpr[7][13] ), .B(n4675), .Z(n3887) );
  ND2I U3552 ( .A(\gpr[6][13] ), .B(n4524), .Z(n3886) );
  ND4 U3553 ( .A(n3889), .B(n3888), .C(n3887), .D(n3886), .Z(n3890) );
  NR2I U3554 ( .A(n3891), .B(n3890), .Z(n3892) );
  ND2I U3555 ( .A(n3893), .B(n3892), .Z(n3894) );
  AN2I U3556 ( .A(n3895), .B(n3894), .Z(rd_data2[13]) );
  B4IP U3557 ( .A(wr_data[14]), .Z(n3896) );
  MUX21L U3558 ( .A(n4830), .B(n3896), .S(n3981), .Z(n2433) );
  MUX21L U3559 ( .A(n5225), .B(n3896), .S(n3980), .Z(n2465) );
  MUX21L U3560 ( .A(n5226), .B(n3896), .S(n3982), .Z(n2593) );
  MUX21L U3561 ( .A(n5227), .B(n3896), .S(n3983), .Z(n2561) );
  MUX21L U3562 ( .A(n5228), .B(n3896), .S(n3976), .Z(n2401) );
  MUX21L U3563 ( .A(n5229), .B(n3896), .S(n3977), .Z(n2529) );
  MUX21L U3564 ( .A(n5230), .B(n3896), .S(n4600), .Z(n2497) );
  MUX21L U3565 ( .A(n5231), .B(n3896), .S(n3975), .Z(n2369) );
  MUX21L U3566 ( .A(n5232), .B(n3896), .S(n3996), .Z(n2689) );
  MUX21L U3567 ( .A(n5233), .B(n3896), .S(n3997), .Z(n2721) );
  MUX21L U3568 ( .A(n5234), .B(n3896), .S(n3998), .Z(n2849) );
  MUX21L U3569 ( .A(n5235), .B(n3896), .S(n3999), .Z(n2817) );
  MUX21L U3570 ( .A(n5236), .B(n3896), .S(n4594), .Z(n2657) );
  MUX21L U3571 ( .A(n5237), .B(n3896), .S(n3978), .Z(n2785) );
  MUX21L U3572 ( .A(n5238), .B(n3896), .S(n4592), .Z(n2753) );
  MUX21L U3573 ( .A(n4860), .B(n3896), .S(n4597), .Z(n2625) );
  MUX21L U3574 ( .A(n5239), .B(n3896), .S(n3988), .Z(n2977) );
  MUX21L U3575 ( .A(n5240), .B(n3896), .S(n3989), .Z(n3105) );
  MUX21L U3576 ( .A(n5241), .B(n3896), .S(n4608), .Z(n3009) );
  MUX21L U3577 ( .A(n5242), .B(n3896), .S(n3990), .Z(n3073) );
  MUX21L U3578 ( .A(n4772), .B(n3896), .S(n3991), .Z(n2913) );
  MUX21L U3579 ( .A(n5243), .B(n3896), .S(n3992), .Z(n3041) );
  MUX21L U3580 ( .A(n5244), .B(n3896), .S(n3984), .Z(n2881) );
  MUX21L U3581 ( .A(n4766), .B(n3896), .S(n3985), .Z(n2945) );
  MUX21L U3582 ( .A(n5245), .B(n3896), .S(n3986), .Z(n3233) );
  MUX21L U3583 ( .A(n5246), .B(n3896), .S(n4615), .Z(n3297) );
  MUX21L U3584 ( .A(n5247), .B(n3896), .S(n3993), .Z(n3137) );
  MUX21L U3585 ( .A(n5248), .B(n3896), .S(n3994), .Z(n3169) );
  MUX21L U3586 ( .A(n5249), .B(n3896), .S(n3995), .Z(n3201) );
  MUX21L U3587 ( .A(n5250), .B(n3896), .S(n3987), .Z(n3329) );
  MUX21L U3588 ( .A(n5251), .B(n3896), .S(n4620), .Z(n3265) );
  AO2 U3589 ( .A(\gpr[26][14] ), .B(n4293), .C(\gpr[24][14] ), .D(n4626), .Z(
        n3905) );
  AO2 U3590 ( .A(\gpr[25][14] ), .B(n4001), .C(\gpr[28][14] ), .D(n219), .Z(
        n3904) );
  AO2 U3591 ( .A(\gpr[31][14] ), .B(n4457), .C(\gpr[29][14] ), .D(n4090), .Z(
        n3903) );
  ND2I U3592 ( .A(\gpr[30][14] ), .B(n4431), .Z(n3898) );
  IVI U3593 ( .A(n3898), .Z(n3901) );
  ND2I U3594 ( .A(\gpr[27][14] ), .B(n3660), .Z(n3899) );
  ND2I U3595 ( .A(n4453), .B(n3899), .Z(n3900) );
  NR2I U3596 ( .A(n3901), .B(n3900), .Z(n3902) );
  ND4 U3597 ( .A(n3905), .B(n3904), .C(n3903), .D(n3902), .Z(n3915) );
  AO2 U3598 ( .A(\gpr[16][14] ), .B(n4357), .C(\gpr[18][14] ), .D(n4293), .Z(
        n3913) );
  AO2 U3599 ( .A(\gpr[17][14] ), .B(n4296), .C(\gpr[20][14] ), .D(n220), .Z(
        n3912) );
  AO2 U3600 ( .A(\gpr[21][14] ), .B(n4090), .C(\gpr[23][14] ), .D(n4251), .Z(
        n3911) );
  ND2I U3601 ( .A(\gpr[22][14] ), .B(n4431), .Z(n3906) );
  IVI U3602 ( .A(n3906), .Z(n3909) );
  ND2I U3603 ( .A(\gpr[19][14] ), .B(n4623), .Z(n3907) );
  ND2I U3604 ( .A(n4628), .B(n3907), .Z(n3908) );
  NR2I U3605 ( .A(n3909), .B(n3908), .Z(n3910) );
  ND4 U3606 ( .A(n3913), .B(n3912), .C(n3911), .D(n3910), .Z(n3914) );
  AN2I U3607 ( .A(n3915), .B(n3914), .Z(n3937) );
  ND2I U3608 ( .A(n4766), .B(n4184), .Z(n3916) );
  AO3 U3609 ( .A(\gpr[15][14] ), .B(n4090), .C(n4652), .D(n3916), .Z(n3917) );
  AO3 U3610 ( .A(n4772), .B(n4150), .C(n295), .D(n3917), .Z(n3923) );
  ND2I U3611 ( .A(\gpr[3][14] ), .B(n4657), .Z(n3921) );
  ND2I U3612 ( .A(\gpr[5][14] ), .B(n4658), .Z(n3920) );
  ND2I U3613 ( .A(\gpr[1][14] ), .B(n4656), .Z(n3919) );
  ND2I U3614 ( .A(\gpr[4][14] ), .B(n4308), .Z(n3918) );
  ND4 U3615 ( .A(n3921), .B(n3920), .C(n3919), .D(n3918), .Z(n3922) );
  NR2I U3616 ( .A(n3923), .B(n3922), .Z(n3935) );
  ND2I U3617 ( .A(\gpr[2][14] ), .B(n4659), .Z(n3927) );
  ND2I U3618 ( .A(n4473), .B(\gpr[10][14] ), .Z(n3926) );
  ND2I U3619 ( .A(\gpr[9][14] ), .B(n4474), .Z(n3925) );
  ND2I U3620 ( .A(\gpr[8][14] ), .B(n3720), .Z(n3924) );
  ND4 U3621 ( .A(n3927), .B(n3926), .C(n3925), .D(n3924), .Z(n3933) );
  ND2I U3622 ( .A(\gpr[11][14] ), .B(n4320), .Z(n3931) );
  ND2I U3623 ( .A(\gpr[12][14] ), .B(n4321), .Z(n3930) );
  ND2I U3624 ( .A(\gpr[7][14] ), .B(n4675), .Z(n3929) );
  ND2I U3625 ( .A(\gpr[6][14] ), .B(n4674), .Z(n3928) );
  ND4 U3626 ( .A(n3931), .B(n3930), .C(n3929), .D(n3928), .Z(n3932) );
  NR2I U3627 ( .A(n3933), .B(n3932), .Z(n3934) );
  ND2I U3628 ( .A(n3935), .B(n3934), .Z(n3936) );
  AN2I U3629 ( .A(n3937), .B(n3936), .Z(rd_data2[14]) );
  B4IP U3630 ( .A(wr_data[15]), .Z(n3938) );
  MUX21L U3631 ( .A(n5252), .B(n3938), .S(n4597), .Z(n2626) );
  MUX21L U3632 ( .A(n5253), .B(n3938), .S(n3996), .Z(n2690) );
  MUX21L U3633 ( .A(n5254), .B(n3938), .S(n4592), .Z(n2754) );
  MUX21L U3634 ( .A(n5255), .B(n3938), .S(n3999), .Z(n2818) );
  MUX21L U3635 ( .A(n4862), .B(n3938), .S(n4594), .Z(n2658) );
  MUX21L U3636 ( .A(n5256), .B(n3938), .S(n4595), .Z(n2786) );
  MUX21L U3637 ( .A(n5702), .B(n3938), .S(n3998), .Z(n2850) );
  MUX21L U3638 ( .A(n5257), .B(n3938), .S(n3997), .Z(n2722) );
  MUX21L U3639 ( .A(n5258), .B(n3938), .S(n4605), .Z(n2370) );
  MUX21L U3640 ( .A(n5259), .B(n3938), .S(n3981), .Z(n2434) );
  MUX21L U3641 ( .A(n5260), .B(n3938), .S(n3982), .Z(n2594) );
  MUX21L U3642 ( .A(n5261), .B(n3938), .S(n4600), .Z(n2498) );
  MUX21L U3643 ( .A(n4861), .B(n3938), .S(n4602), .Z(n2402) );
  MUX21L U3644 ( .A(n5262), .B(n3938), .S(n4603), .Z(n2530) );
  MUX21L U3645 ( .A(n5263), .B(n3938), .S(n3983), .Z(n2562) );
  MUX21L U3646 ( .A(n5264), .B(n3938), .S(n3980), .Z(n2466) );
  MUX21L U3647 ( .A(n5265), .B(n3938), .S(n3988), .Z(n2978) );
  MUX21L U3648 ( .A(n5266), .B(n3938), .S(n3989), .Z(n3106) );
  MUX21L U3649 ( .A(n5267), .B(n3938), .S(n4608), .Z(n3010) );
  MUX21L U3650 ( .A(n5268), .B(n3938), .S(n3990), .Z(n3074) );
  MUX21L U3651 ( .A(n4819), .B(n3938), .S(n3991), .Z(n2914) );
  MUX21L U3652 ( .A(n5269), .B(n3938), .S(n3992), .Z(n3042) );
  MUX21L U3653 ( .A(n5270), .B(n3938), .S(n3984), .Z(n2882) );
  MUX21L U3654 ( .A(n4787), .B(n3938), .S(n3985), .Z(n2946) );
  MUX21L U3655 ( .A(n5271), .B(n3938), .S(n3986), .Z(n3234) );
  MUX21L U3656 ( .A(n5272), .B(n3938), .S(n4615), .Z(n3298) );
  MUX21L U3657 ( .A(n5273), .B(n3938), .S(n3993), .Z(n3138) );
  MUX21L U3658 ( .A(n5274), .B(n3938), .S(n3994), .Z(n3170) );
  MUX21L U3659 ( .A(n5275), .B(n3938), .S(n3995), .Z(n3202) );
  MUX21L U3660 ( .A(n5276), .B(n3938), .S(n3987), .Z(n3330) );
  MUX21L U3661 ( .A(n5277), .B(n3938), .S(n4620), .Z(n3266) );
  AO2 U3662 ( .A(\gpr[20][15] ), .B(n4498), .C(\gpr[18][15] ), .D(n4622), .Z(
        n3942) );
  AO2 U3663 ( .A(\gpr[17][15] ), .B(n4001), .C(\gpr[19][15] ), .D(n4009), .Z(
        n3941) );
  AO2 U3664 ( .A(\gpr[21][15] ), .B(n4090), .C(\gpr[22][15] ), .D(n4431), .Z(
        n3940) );
  ND4 U3665 ( .A(n3942), .B(n3941), .C(n3940), .D(n3939), .Z(n3950) );
  AO2 U3666 ( .A(\gpr[28][15] ), .B(n4498), .C(\gpr[26][15] ), .D(n4458), .Z(
        n3948) );
  AO2 U3667 ( .A(\gpr[27][15] ), .B(n4009), .C(\gpr[24][15] ), .D(n4450), .Z(
        n3947) );
  AO2 U3668 ( .A(\gpr[29][15] ), .B(n4097), .C(\gpr[30][15] ), .D(n4431), .Z(
        n3946) );
  ND2I U3669 ( .A(\gpr[31][15] ), .B(n4543), .Z(n3944) );
  ND2I U3670 ( .A(\gpr[25][15] ), .B(n4490), .Z(n3943) );
  AN3 U3671 ( .A(n4453), .B(n3944), .C(n3943), .Z(n3945) );
  ND4 U3672 ( .A(n3948), .B(n3947), .C(n3946), .D(n3945), .Z(n3949) );
  AN2I U3673 ( .A(n3950), .B(n3949), .Z(n3974) );
  ND2I U3674 ( .A(n4787), .B(n4184), .Z(n3951) );
  AO3 U3675 ( .A(\gpr[15][15] ), .B(n4090), .C(n4652), .D(n3951), .Z(n3952) );
  AO3 U3676 ( .A(n4819), .B(n3953), .C(n295), .D(n3952), .Z(n3959) );
  ND2I U3677 ( .A(\gpr[3][15] ), .B(n4557), .Z(n3957) );
  ND2I U3678 ( .A(\gpr[5][15] ), .B(n4658), .Z(n3956) );
  ND2I U3679 ( .A(\gpr[1][15] ), .B(n4656), .Z(n3955) );
  ND2I U3680 ( .A(\gpr[4][15] ), .B(n4666), .Z(n3954) );
  ND4 U3681 ( .A(n3957), .B(n3956), .C(n3955), .D(n3954), .Z(n3958) );
  NR2I U3682 ( .A(n3959), .B(n3958), .Z(n3972) );
  ND2I U3683 ( .A(\gpr[2][15] ), .B(n4659), .Z(n3964) );
  ND2I U3684 ( .A(n4473), .B(\gpr[10][15] ), .Z(n3963) );
  ND2I U3685 ( .A(\gpr[9][15] ), .B(n4668), .Z(n3962) );
  ND2I U3686 ( .A(\gpr[8][15] ), .B(n3960), .Z(n3961) );
  ND4 U3687 ( .A(n3964), .B(n3963), .C(n3962), .D(n3961), .Z(n3970) );
  ND2I U3688 ( .A(\gpr[11][15] ), .B(n4667), .Z(n3968) );
  ND2I U3689 ( .A(\gpr[12][15] ), .B(n4673), .Z(n3967) );
  ND2I U3690 ( .A(\gpr[7][15] ), .B(n4675), .Z(n3966) );
  ND2I U3691 ( .A(\gpr[6][15] ), .B(n4674), .Z(n3965) );
  ND4 U3692 ( .A(n3968), .B(n3967), .C(n3966), .D(n3965), .Z(n3969) );
  NR2I U3693 ( .A(n3970), .B(n3969), .Z(n3971) );
  ND2I U3694 ( .A(n3972), .B(n3971), .Z(n3973) );
  AN2I U3695 ( .A(n3974), .B(n3973), .Z(rd_data2[15]) );
  B4IP U3696 ( .A(wr_data[16]), .Z(n3979) );
  MUX21L U3697 ( .A(n5278), .B(n3979), .S(n3975), .Z(n2371) );
  MUX21L U3698 ( .A(n4831), .B(n3979), .S(n3981), .Z(n2435) );
  MUX21L U3699 ( .A(n5279), .B(n3979), .S(n3982), .Z(n2595) );
  MUX21L U3700 ( .A(n5280), .B(n3979), .S(n4600), .Z(n2499) );
  MUX21L U3701 ( .A(n5281), .B(n3979), .S(n3976), .Z(n2403) );
  MUX21L U3702 ( .A(n5282), .B(n3979), .S(n3977), .Z(n2531) );
  MUX21L U3703 ( .A(n5283), .B(n3979), .S(n3983), .Z(n2563) );
  MUX21L U3704 ( .A(n5284), .B(n3979), .S(n3980), .Z(n2467) );
  MUX21L U3705 ( .A(n4807), .B(n3979), .S(n3996), .Z(n2691) );
  MUX21L U3706 ( .A(n5285), .B(n3979), .S(n3997), .Z(n2723) );
  MUX21L U3707 ( .A(n5286), .B(n3979), .S(n4592), .Z(n2755) );
  MUX21L U3708 ( .A(n5287), .B(n3979), .S(n3999), .Z(n2819) );
  MUX21L U3709 ( .A(n5288), .B(n3979), .S(n4594), .Z(n2659) );
  MUX21L U3710 ( .A(n5289), .B(n3979), .S(n3978), .Z(n2787) );
  MUX21L U3711 ( .A(n5290), .B(n3979), .S(n3998), .Z(n2851) );
  MUX21L U3712 ( .A(n5291), .B(n3979), .S(n4597), .Z(n2627) );
  MUX21L U3713 ( .A(n5292), .B(n3979), .S(n3988), .Z(n2979) );
  MUX21L U3714 ( .A(n5293), .B(n3979), .S(n3989), .Z(n3107) );
  MUX21L U3715 ( .A(n5294), .B(n3979), .S(n4608), .Z(n3011) );
  MUX21L U3716 ( .A(n5295), .B(n3979), .S(n3990), .Z(n3075) );
  MUX21L U3717 ( .A(n4773), .B(n3979), .S(n3991), .Z(n2915) );
  MUX21L U3718 ( .A(n5296), .B(n3979), .S(n3992), .Z(n3043) );
  MUX21L U3719 ( .A(n5297), .B(n3979), .S(n3984), .Z(n2883) );
  MUX21L U3720 ( .A(n4767), .B(n3979), .S(n3985), .Z(n2947) );
  MUX21L U3721 ( .A(n5298), .B(n3979), .S(n3986), .Z(n3235) );
  MUX21L U3722 ( .A(n5299), .B(n3979), .S(n4615), .Z(n3299) );
  MUX21L U3723 ( .A(n5300), .B(n3979), .S(n3993), .Z(n3139) );
  MUX21L U3724 ( .A(n5301), .B(n3979), .S(n3994), .Z(n3171) );
  MUX21L U3725 ( .A(n5302), .B(n3979), .S(n3995), .Z(n3203) );
  MUX21L U3726 ( .A(n5303), .B(n3979), .S(n3987), .Z(n3331) );
  MUX21L U3727 ( .A(n5304), .B(n3979), .S(n4620), .Z(n3267) );
  MUX21L U3728 ( .A(n304), .B(n4000), .S(n3980), .Z(n2468) );
  MUX21L U3729 ( .A(n5305), .B(n4000), .S(n4600), .Z(n2500) );
  MUX21L U3730 ( .A(n5306), .B(n4000), .S(n4605), .Z(n2372) );
  MUX21L U3731 ( .A(n5307), .B(n4000), .S(n3981), .Z(n2436) );
  MUX21L U3732 ( .A(n5308), .B(n4000), .S(n3982), .Z(n2596) );
  MUX21L U3733 ( .A(n5309), .B(n4000), .S(n3983), .Z(n2564) );
  MUX21L U3734 ( .A(n4864), .B(n4000), .S(n4602), .Z(n2404) );
  MUX21L U3735 ( .A(n4789), .B(n4000), .S(n4603), .Z(n2532) );
  MUX21L U3736 ( .A(n5310), .B(n4000), .S(n3984), .Z(n2884) );
  MUX21L U3737 ( .A(n4790), .B(n4000), .S(n3985), .Z(n2948) );
  MUX21L U3738 ( .A(n5311), .B(n4000), .S(n3986), .Z(n3236) );
  MUX21L U3739 ( .A(n5312), .B(n4000), .S(n3987), .Z(n3332) );
  MUX21L U3740 ( .A(n5313), .B(n4000), .S(n4620), .Z(n3268) );
  MUX21L U3741 ( .A(n5314), .B(n4000), .S(n3988), .Z(n2980) );
  MUX21L U3742 ( .A(n5315), .B(n4000), .S(n3989), .Z(n3108) );
  MUX21L U3743 ( .A(n5316), .B(n4000), .S(n4608), .Z(n3012) );
  MUX21L U3744 ( .A(n5317), .B(n4000), .S(n3990), .Z(n3076) );
  MUX21L U3745 ( .A(n5703), .B(n4000), .S(n3991), .Z(n2916) );
  MUX21L U3746 ( .A(n4839), .B(n4000), .S(n3992), .Z(n3044) );
  MUX21L U3747 ( .A(n5318), .B(n4000), .S(n4615), .Z(n3300) );
  MUX21L U3748 ( .A(n5319), .B(n4000), .S(n3993), .Z(n3140) );
  MUX21L U3749 ( .A(n5320), .B(n4000), .S(n3994), .Z(n3172) );
  MUX21L U3750 ( .A(n5321), .B(n4000), .S(n3995), .Z(n3204) );
  MUX21L U3751 ( .A(n5322), .B(n4000), .S(n4597), .Z(n2628) );
  MUX21L U3752 ( .A(n5323), .B(n4000), .S(n3996), .Z(n2692) );
  MUX21L U3753 ( .A(n305), .B(n4000), .S(n3997), .Z(n2724) );
  MUX21L U3754 ( .A(n5324), .B(n4000), .S(n3998), .Z(n2852) );
  MUX21L U3755 ( .A(n5325), .B(n4000), .S(n4592), .Z(n2756) );
  MUX21L U3756 ( .A(n5326), .B(n4000), .S(n3999), .Z(n2820) );
  MUX21L U3757 ( .A(n4863), .B(n4000), .S(n4594), .Z(n2660) );
  MUX21L U3758 ( .A(n4788), .B(n4000), .S(n4595), .Z(n2788) );
  AO2 U3759 ( .A(\gpr[17][17] ), .B(n4001), .C(\gpr[19][17] ), .D(n4009), .Z(
        n4008) );
  AO2 U3760 ( .A(\gpr[20][17] ), .B(n4498), .C(\gpr[16][17] ), .D(n4432), .Z(
        n4007) );
  AO2 U3761 ( .A(\gpr[21][17] ), .B(n4090), .C(\gpr[22][17] ), .D(n4431), .Z(
        n4006) );
  ND2I U3762 ( .A(\gpr[23][17] ), .B(n4002), .Z(n4003) );
  AO3 U3763 ( .A(n4356), .B(n4788), .C(n4628), .D(n4003), .Z(n4004) );
  IVI U3764 ( .A(n4004), .Z(n4005) );
  ND4 U3765 ( .A(n4008), .B(n4007), .C(n4006), .D(n4005), .Z(n4017) );
  AO2 U3766 ( .A(\gpr[25][17] ), .B(n4296), .C(\gpr[24][17] ), .D(n4626), .Z(
        n4015) );
  AO2 U3767 ( .A(\gpr[29][17] ), .B(n4097), .C(\gpr[27][17] ), .D(n4009), .Z(
        n4014) );
  AO2 U3768 ( .A(\gpr[28][17] ), .B(n4624), .C(\gpr[30][17] ), .D(n4431), .Z(
        n4013) );
  ND2I U3769 ( .A(\gpr[31][17] ), .B(n4342), .Z(n4010) );
  AO3 U3770 ( .A(n4356), .B(n4789), .C(n4641), .D(n4010), .Z(n4011) );
  IVI U3771 ( .A(n4011), .Z(n4012) );
  ND4 U3772 ( .A(n4015), .B(n4014), .C(n4013), .D(n4012), .Z(n4016) );
  AN2I U3773 ( .A(n4017), .B(n4016), .Z(n4035) );
  ND2I U3774 ( .A(\gpr[5][17] ), .B(n4658), .Z(n4022) );
  ND2I U3775 ( .A(n4790), .B(n4184), .Z(n4018) );
  AO3 U3776 ( .A(\gpr[15][17] ), .B(n4097), .C(n4652), .D(n4018), .Z(n4021) );
  ND2I U3777 ( .A(\gpr[2][17] ), .B(n4659), .Z(n4020) );
  ND2I U3778 ( .A(\gpr[3][17] ), .B(n4557), .Z(n4019) );
  ND4 U3779 ( .A(n4022), .B(n4021), .C(n4020), .D(n4019), .Z(n4024) );
  NR2I U3780 ( .A(n4024), .B(n4023), .Z(n4033) );
  ND2I U3781 ( .A(\gpr[14][17] ), .B(n4625), .Z(n4025) );
  AO3 U3782 ( .A(n4839), .B(n4356), .C(n4561), .D(n4025), .Z(n4031) );
  ND2I U3783 ( .A(\gpr[9][17] ), .B(n4490), .Z(n4029) );
  ND2I U3784 ( .A(\gpr[8][17] ), .B(n4542), .Z(n4028) );
  ND2I U3785 ( .A(\gpr[11][17] ), .B(n4623), .Z(n4027) );
  ND2I U3786 ( .A(\gpr[12][17] ), .B(n4498), .Z(n4026) );
  ND4 U3787 ( .A(n4029), .B(n4028), .C(n4027), .D(n4026), .Z(n4030) );
  AO7 U3788 ( .A(n4031), .B(n4030), .C(n4362), .Z(n4032) );
  ND2I U3789 ( .A(n4033), .B(n4032), .Z(n4034) );
  AN2I U3790 ( .A(n4035), .B(n4034), .Z(rd_data2[17]) );
  B4IP U3791 ( .A(wr_data[18]), .Z(n4053) );
  B2IP U3792 ( .A(n4036), .Z1(n3525), .Z2(n4598) );
  MUX21L U3793 ( .A(n5327), .B(n4053), .S(n4598), .Z(n2437) );
  B4I U3794 ( .A(n4037), .Z(n4599) );
  MUX21L U3795 ( .A(n5328), .B(n4053), .S(n4599), .Z(n2597) );
  MUX21L U3796 ( .A(n5329), .B(n4053), .S(n4600), .Z(n2501) );
  MUX21L U3797 ( .A(n5330), .B(n4053), .S(n4601), .Z(n2565) );
  MUX21L U3798 ( .A(n5331), .B(n4053), .S(n4602), .Z(n2405) );
  MUX21L U3799 ( .A(n5332), .B(n4053), .S(n4603), .Z(n2533) );
  B4I U3800 ( .A(n4038), .Z(n4604) );
  MUX21L U3801 ( .A(n4770), .B(n4053), .S(n4604), .Z(n2469) );
  MUX21L U3802 ( .A(n5333), .B(n4053), .S(n4605), .Z(n2373) );
  MUX21L U3803 ( .A(n5334), .B(n4053), .S(n4536), .Z(n2629) );
  MUX21L U3804 ( .A(n5335), .B(n4053), .S(n4590), .Z(n2693) );
  B4I U3805 ( .A(n4039), .Z(n4591) );
  MUX21L U3806 ( .A(n5336), .B(n4053), .S(n4591), .Z(n2725) );
  MUX21L U3807 ( .A(n5337), .B(n4053), .S(n4592), .Z(n2757) );
  MUX21L U3808 ( .A(n4865), .B(n4053), .S(n4538), .Z(n2661) );
  MUX21L U3809 ( .A(n5338), .B(n4053), .S(n4595), .Z(n2789) );
  B4I U3810 ( .A(n4040), .Z(n4596) );
  MUX21L U3811 ( .A(n5339), .B(n4053), .S(n4596), .Z(n2853) );
  MUX21L U3812 ( .A(n5340), .B(n4053), .S(n4593), .Z(n2821) );
  B4I U3813 ( .A(n4041), .Z(n4606) );
  MUX21L U3814 ( .A(n306), .B(n4053), .S(n4606), .Z(n2981) );
  B4I U3815 ( .A(n4042), .Z(n4607) );
  MUX21L U3816 ( .A(n5341), .B(n4053), .S(n4607), .Z(n3109) );
  MUX21L U3817 ( .A(n307), .B(n4053), .S(n4608), .Z(n3013) );
  B2IP U3818 ( .A(n4043), .Z1(n3533), .Z2(n4609) );
  MUX21L U3819 ( .A(n308), .B(n4053), .S(n4609), .Z(n3077) );
  B4I U3820 ( .A(n4044), .Z(n4610) );
  MUX21L U3821 ( .A(n5342), .B(n4053), .S(n4610), .Z(n2917) );
  B4I U3822 ( .A(n4045), .Z(n4611) );
  MUX21L U3823 ( .A(n309), .B(n4053), .S(n4611), .Z(n3045) );
  B4I U3824 ( .A(n4046), .Z(n4612) );
  MUX21L U3825 ( .A(n5343), .B(n4053), .S(n4612), .Z(n2885) );
  B2IP U3826 ( .A(n4047), .Z1(n3531), .Z2(n4613) );
  MUX21L U3827 ( .A(n4791), .B(n4053), .S(n4613), .Z(n2949) );
  B4I U3828 ( .A(n4048), .Z(n4614) );
  MUX21L U3829 ( .A(n5704), .B(n4053), .S(n4614), .Z(n3237) );
  MUX21L U3830 ( .A(n5344), .B(n4053), .S(n4540), .Z(n3301) );
  B4I U3831 ( .A(n4049), .Z(n4616) );
  MUX21L U3832 ( .A(n5345), .B(n4053), .S(n4616), .Z(n3141) );
  B4I U3833 ( .A(n4050), .Z(n4617) );
  MUX21L U3834 ( .A(n310), .B(n4053), .S(n4617), .Z(n3173) );
  B2IP U3835 ( .A(n4051), .Z1(n3535), .Z2(n4618) );
  MUX21L U3836 ( .A(n4759), .B(n4053), .S(n4618), .Z(n3205) );
  B2IP U3837 ( .A(n4052), .Z1(n3536), .Z2(n4619) );
  MUX21L U3838 ( .A(n311), .B(n4053), .S(n4619), .Z(n3333) );
  MUX21L U3839 ( .A(n5346), .B(n4053), .S(n4620), .Z(n3269) );
  IVI U3840 ( .A(n4054), .Z(n4635) );
  AO2 U3841 ( .A(\gpr[25][18] ), .B(n4296), .C(\gpr[24][18] ), .D(n4357), .Z(
        n4059) );
  IVI U3842 ( .A(n4498), .Z(n4056) );
  ND2I U3843 ( .A(\gpr[30][18] ), .B(n4625), .Z(n4055) );
  AO3P U3844 ( .A(n4056), .B(n4770), .C(n4641), .D(n4055), .Z(n4057) );
  IVI U3845 ( .A(n4057), .Z(n4058) );
  AO2 U3846 ( .A(\gpr[18][18] ), .B(n4214), .C(\gpr[17][18] ), .D(n4296), .Z(
        n4067) );
  AO2 U3847 ( .A(\gpr[20][18] ), .B(n4498), .C(\gpr[19][18] ), .D(n4635), .Z(
        n4066) );
  AO2 U3848 ( .A(\gpr[21][18] ), .B(n4097), .C(\gpr[22][18] ), .D(n4431), .Z(
        n4065) );
  AN2I U3849 ( .A(\gpr[23][18] ), .B(n4060), .Z(n4063) );
  ND2I U3850 ( .A(\gpr[16][18] ), .B(n4549), .Z(n4061) );
  ND2I U3851 ( .A(n4628), .B(n4061), .Z(n4062) );
  NR2I U3852 ( .A(n4063), .B(n4062), .Z(n4064) );
  ND4 U3853 ( .A(n4067), .B(n4066), .C(n4065), .D(n4064), .Z(n4068) );
  AN2I U3854 ( .A(n4069), .B(n4068), .Z(n4088) );
  AO2 U3855 ( .A(\gpr[2][18] ), .B(n4659), .C(\gpr[7][18] ), .D(n4675), .Z(
        n4085) );
  AO2 U3856 ( .A(\gpr[1][18] ), .B(n4656), .C(\gpr[3][18] ), .D(n4657), .Z(
        n4073) );
  ND2I U3857 ( .A(\gpr[4][18] ), .B(n4308), .Z(n4071) );
  ND2I U3858 ( .A(n4658), .B(\gpr[5][18] ), .Z(n4070) );
  AN2I U3859 ( .A(n4071), .B(n4070), .Z(n4072) );
  AN2I U3860 ( .A(n4073), .B(n4072), .Z(n4084) );
  AO2 U3861 ( .A(\gpr[8][18] ), .B(n4542), .C(\gpr[14][18] ), .D(n4431), .Z(
        n4081) );
  ND2I U3862 ( .A(\gpr[10][18] ), .B(n4487), .Z(n4075) );
  ND2I U3863 ( .A(\gpr[9][18] ), .B(n4490), .Z(n4074) );
  ND2I U3864 ( .A(n4075), .B(n4074), .Z(n4079) );
  ND2I U3865 ( .A(\gpr[11][18] ), .B(n4501), .Z(n4077) );
  ND2I U3866 ( .A(\gpr[12][18] ), .B(n4498), .Z(n4076) );
  ND2I U3867 ( .A(n4077), .B(n4076), .Z(n4078) );
  NR2I U3868 ( .A(n4079), .B(n4078), .Z(n4080) );
  ND2I U3869 ( .A(n4081), .B(n4080), .Z(n4082) );
  ND2I U3870 ( .A(n4442), .B(n4082), .Z(n4083) );
  ND4 U3871 ( .A(n4086), .B(n4085), .C(n4084), .D(n4083), .Z(n4087) );
  AN2I U3872 ( .A(n4088), .B(n4087), .Z(rd_data2[18]) );
  B4IP U3873 ( .A(wr_data[19]), .Z(n4089) );
  MUX21L U3874 ( .A(n5347), .B(n4089), .S(n4590), .Z(n2694) );
  MUX21L U3875 ( .A(n312), .B(n4089), .S(n4591), .Z(n2726) );
  MUX21L U3876 ( .A(n5348), .B(n4089), .S(n4596), .Z(n2854) );
  MUX21L U3877 ( .A(n5349), .B(n4089), .S(n4592), .Z(n2758) );
  MUX21L U3878 ( .A(n4867), .B(n4089), .S(n4538), .Z(n2662) );
  MUX21L U3879 ( .A(n5350), .B(n4089), .S(n4595), .Z(n2790) );
  MUX21L U3880 ( .A(n5351), .B(n4089), .S(n4593), .Z(n2822) );
  MUX21L U3881 ( .A(n5352), .B(n4089), .S(n4536), .Z(n2630) );
  MUX21L U3882 ( .A(n5353), .B(n4089), .S(n4598), .Z(n2438) );
  MUX21L U3883 ( .A(n313), .B(n4089), .S(n4604), .Z(n2470) );
  MUX21L U3884 ( .A(n5354), .B(n4089), .S(n4600), .Z(n2502) );
  MUX21L U3885 ( .A(n5355), .B(n4089), .S(n4601), .Z(n2566) );
  MUX21L U3886 ( .A(n4866), .B(n4089), .S(n4602), .Z(n2406) );
  MUX21L U3887 ( .A(n5356), .B(n4089), .S(n4603), .Z(n2534) );
  MUX21L U3888 ( .A(n5705), .B(n4089), .S(n4599), .Z(n2598) );
  MUX21L U3889 ( .A(n5357), .B(n4089), .S(n4605), .Z(n2374) );
  MUX21L U3890 ( .A(n5358), .B(n4089), .S(n4606), .Z(n2982) );
  MUX21L U3891 ( .A(n5359), .B(n4089), .S(n4607), .Z(n3110) );
  MUX21L U3892 ( .A(n5360), .B(n4089), .S(n4608), .Z(n3014) );
  MUX21L U3893 ( .A(n5361), .B(n4089), .S(n4609), .Z(n3078) );
  MUX21L U3894 ( .A(n4820), .B(n4089), .S(n4610), .Z(n2918) );
  MUX21L U3895 ( .A(n5362), .B(n4089), .S(n4611), .Z(n3046) );
  MUX21L U3896 ( .A(n5363), .B(n4089), .S(n4612), .Z(n2886) );
  MUX21L U3897 ( .A(n4792), .B(n4089), .S(n4613), .Z(n2950) );
  MUX21L U3898 ( .A(n5364), .B(n4089), .S(n4614), .Z(n3238) );
  MUX21L U3899 ( .A(n5365), .B(n4089), .S(n4540), .Z(n3302) );
  MUX21L U3900 ( .A(n5366), .B(n4089), .S(n4616), .Z(n3142) );
  MUX21L U3901 ( .A(n5367), .B(n4089), .S(n4617), .Z(n3174) );
  MUX21L U3902 ( .A(n5368), .B(n4089), .S(n4618), .Z(n3206) );
  MUX21L U3903 ( .A(n5369), .B(n4089), .S(n4619), .Z(n3334) );
  MUX21L U3904 ( .A(n5370), .B(n4089), .S(n4620), .Z(n3270) );
  AO2 U3905 ( .A(\gpr[18][19] ), .B(n4487), .C(\gpr[16][19] ), .D(n4357), .Z(
        n4096) );
  AO2 U3906 ( .A(\gpr[20][19] ), .B(n4498), .C(\gpr[19][19] ), .D(n4635), .Z(
        n4095) );
  AO2 U3907 ( .A(\gpr[21][19] ), .B(n4090), .C(\gpr[23][19] ), .D(n4543), .Z(
        n4094) );
  ND2I U3908 ( .A(\gpr[22][19] ), .B(n4625), .Z(n4092) );
  ND2I U3909 ( .A(\gpr[17][19] ), .B(n4490), .Z(n4091) );
  AN3 U3910 ( .A(n4628), .B(n4092), .C(n4091), .Z(n4093) );
  ND4 U3911 ( .A(n4096), .B(n4095), .C(n4094), .D(n4093), .Z(n4103) );
  AO2 U3912 ( .A(\gpr[26][19] ), .B(n4622), .C(\gpr[27][19] ), .D(n4635), .Z(
        n4101) );
  AO2 U3913 ( .A(\gpr[28][19] ), .B(n4624), .C(\gpr[25][19] ), .D(n4296), .Z(
        n4100) );
  AO2 U3914 ( .A(\gpr[29][19] ), .B(n4097), .C(\gpr[31][19] ), .D(n4548), .Z(
        n4099) );
  ND4 U3915 ( .A(n4101), .B(n4100), .C(n4099), .D(n4098), .Z(n4102) );
  AN2I U3916 ( .A(n4103), .B(n4102), .Z(n4128) );
  IVI U3917 ( .A(n4104), .Z(n4105) );
  B4IP U3918 ( .A(n4105), .Z(n4639) );
  ND2I U3919 ( .A(n4792), .B(n4184), .Z(n4106) );
  AO3 U3920 ( .A(\gpr[15][19] ), .B(n4639), .C(n4652), .D(n4106), .Z(n4107) );
  AO3 U3921 ( .A(n4820), .B(n4108), .C(n4561), .D(n4107), .Z(n4114) );
  ND2I U3922 ( .A(\gpr[3][19] ), .B(n4557), .Z(n4112) );
  ND2I U3923 ( .A(\gpr[5][19] ), .B(n4658), .Z(n4111) );
  ND2I U3924 ( .A(\gpr[1][19] ), .B(n4556), .Z(n4110) );
  ND2I U3925 ( .A(\gpr[4][19] ), .B(n4666), .Z(n4109) );
  ND4 U3926 ( .A(n4112), .B(n4111), .C(n4110), .D(n4109), .Z(n4113) );
  NR2I U3927 ( .A(n4114), .B(n4113), .Z(n4126) );
  ND2I U3928 ( .A(\gpr[2][19] ), .B(n4659), .Z(n4118) );
  B2I U3929 ( .A(n4473), .Z2(n4562) );
  ND2I U3930 ( .A(n4562), .B(\gpr[10][19] ), .Z(n4117) );
  ND2I U3931 ( .A(\gpr[9][19] ), .B(n4563), .Z(n4116) );
  ND2I U3932 ( .A(\gpr[8][19] ), .B(n3960), .Z(n4115) );
  ND4 U3933 ( .A(n4118), .B(n4117), .C(n4116), .D(n4115), .Z(n4124) );
  ND2I U3934 ( .A(\gpr[11][19] ), .B(n4571), .Z(n4122) );
  ND2I U3935 ( .A(\gpr[12][19] ), .B(n4573), .Z(n4121) );
  ND2I U3936 ( .A(\gpr[7][19] ), .B(n4675), .Z(n4120) );
  ND2I U3937 ( .A(\gpr[6][19] ), .B(n4197), .Z(n4119) );
  ND4 U3938 ( .A(n4122), .B(n4121), .C(n4120), .D(n4119), .Z(n4123) );
  NR2I U3939 ( .A(n4124), .B(n4123), .Z(n4125) );
  ND2I U3940 ( .A(n4126), .B(n4125), .Z(n4127) );
  AN2I U3941 ( .A(n4128), .B(n4127), .Z(rd_data2[19]) );
  B4IP U3942 ( .A(wr_data[20]), .Z(n4129) );
  MUX21L U3943 ( .A(n4833), .B(n4129), .S(n4598), .Z(n2439) );
  MUX21L U3944 ( .A(n5371), .B(n4129), .S(n4599), .Z(n2599) );
  MUX21L U3945 ( .A(n5372), .B(n4129), .S(n4600), .Z(n2503) );
  MUX21L U3946 ( .A(n5373), .B(n4129), .S(n4601), .Z(n2567) );
  MUX21L U3947 ( .A(n5374), .B(n4129), .S(n4602), .Z(n2407) );
  MUX21L U3948 ( .A(n5375), .B(n4129), .S(n4603), .Z(n2535) );
  MUX21L U3949 ( .A(n5376), .B(n4129), .S(n4604), .Z(n2471) );
  MUX21L U3950 ( .A(n5377), .B(n4129), .S(n4605), .Z(n2375) );
  MUX21L U3951 ( .A(n4832), .B(n4129), .S(n4590), .Z(n2695) );
  MUX21L U3952 ( .A(n5378), .B(n4129), .S(n4591), .Z(n2727) );
  MUX21L U3953 ( .A(n5379), .B(n4129), .S(n4596), .Z(n2855) );
  MUX21L U3954 ( .A(n5380), .B(n4129), .S(n4593), .Z(n2823) );
  MUX21L U3955 ( .A(n5381), .B(n4129), .S(n4538), .Z(n2663) );
  MUX21L U3956 ( .A(n5382), .B(n4129), .S(n4595), .Z(n2791) );
  MUX21L U3957 ( .A(n5383), .B(n4129), .S(n4592), .Z(n2759) );
  MUX21L U3958 ( .A(n5384), .B(n4129), .S(n4536), .Z(n2631) );
  MUX21L U3959 ( .A(n5385), .B(n4129), .S(n4606), .Z(n2983) );
  MUX21L U3960 ( .A(n5386), .B(n4129), .S(n4608), .Z(n3015) );
  MUX21L U3961 ( .A(n5387), .B(n4129), .S(n4609), .Z(n3079) );
  MUX21L U3962 ( .A(n4774), .B(n4129), .S(n4610), .Z(n2919) );
  MUX21L U3963 ( .A(n5388), .B(n4129), .S(n4611), .Z(n3047) );
  MUX21L U3964 ( .A(n5389), .B(n4129), .S(n4612), .Z(n2887) );
  MUX21L U3965 ( .A(n4768), .B(n4129), .S(n4613), .Z(n2951) );
  MUX21L U3966 ( .A(n5390), .B(n4129), .S(n4614), .Z(n3239) );
  MUX21L U3967 ( .A(n5391), .B(n4129), .S(n4540), .Z(n3303) );
  MUX21L U3968 ( .A(n5392), .B(n4129), .S(n4616), .Z(n3143) );
  MUX21L U3969 ( .A(n5393), .B(n4129), .S(n4617), .Z(n3175) );
  MUX21L U3970 ( .A(n5394), .B(n4129), .S(n4618), .Z(n3207) );
  MUX21L U3971 ( .A(n5395), .B(n4129), .S(n4619), .Z(n3335) );
  MUX21L U3972 ( .A(n5396), .B(n4129), .S(n4620), .Z(n3271) );
  AO2 U3973 ( .A(\gpr[27][20] ), .B(n4635), .C(\gpr[26][20] ), .D(n4293), .Z(
        n4137) );
  AO2 U3974 ( .A(\gpr[25][20] ), .B(n4296), .C(\gpr[24][20] ), .D(n4549), .Z(
        n4136) );
  IVI U3975 ( .A(n4130), .Z(n4638) );
  AO2 U3976 ( .A(\gpr[31][20] ), .B(n4638), .C(\gpr[29][20] ), .D(n4639), .Z(
        n4135) );
  AN2I U3977 ( .A(\gpr[30][20] ), .B(n4625), .Z(n4133) );
  ND2I U3978 ( .A(\gpr[28][20] ), .B(n219), .Z(n4131) );
  ND2I U3979 ( .A(n4453), .B(n4131), .Z(n4132) );
  NR2I U3980 ( .A(n4133), .B(n4132), .Z(n4134) );
  ND4 U3981 ( .A(n4137), .B(n4136), .C(n4135), .D(n4134), .Z(n4149) );
  AO2 U3982 ( .A(\gpr[18][20] ), .B(n4293), .C(\gpr[16][20] ), .D(n4497), .Z(
        n4147) );
  ND2I U3983 ( .A(n4138), .B(\gpr[20][20] ), .Z(n4140) );
  ND2I U3984 ( .A(n4296), .B(\gpr[17][20] ), .Z(n4139) );
  AN2I U3985 ( .A(n4140), .B(n4139), .Z(n4146) );
  AO2 U3986 ( .A(\gpr[23][20] ), .B(n4499), .C(\gpr[21][20] ), .D(n4639), .Z(
        n4145) );
  AN2I U3987 ( .A(\gpr[22][20] ), .B(n4625), .Z(n4143) );
  ND2I U3988 ( .A(\gpr[19][20] ), .B(n4623), .Z(n4141) );
  ND2I U3989 ( .A(n4628), .B(n4141), .Z(n4142) );
  NR2I U3990 ( .A(n4143), .B(n4142), .Z(n4144) );
  ND4 U3991 ( .A(n4147), .B(n4146), .C(n4145), .D(n4144), .Z(n4148) );
  AN2I U3992 ( .A(n4149), .B(n4148), .Z(n4170) );
  ND2I U3993 ( .A(n4768), .B(n4184), .Z(n4151) );
  AO3 U3994 ( .A(\gpr[15][20] ), .B(n4639), .C(n4652), .D(n4151), .Z(n4152) );
  ND2I U3995 ( .A(\gpr[3][20] ), .B(n4557), .Z(n4157) );
  ND2I U3996 ( .A(\gpr[5][20] ), .B(n4658), .Z(n4156) );
  ND2I U3997 ( .A(\gpr[1][20] ), .B(n4556), .Z(n4155) );
  ND2I U3998 ( .A(\gpr[4][20] ), .B(n4153), .Z(n4154) );
  ND2I U3999 ( .A(\gpr[2][20] ), .B(n4659), .Z(n4162) );
  ND2I U4000 ( .A(\gpr[10][20] ), .B(n4313), .Z(n4161) );
  ND2I U4001 ( .A(\gpr[9][20] ), .B(n4474), .Z(n4160) );
  ND2I U4002 ( .A(\gpr[8][20] ), .B(n4315), .Z(n4159) );
  ND2I U4003 ( .A(\gpr[11][20] ), .B(n4320), .Z(n4166) );
  ND2I U4004 ( .A(\gpr[12][20] ), .B(n4321), .Z(n4165) );
  ND2I U4005 ( .A(\gpr[7][20] ), .B(n4675), .Z(n4164) );
  ND2I U4006 ( .A(\gpr[6][20] ), .B(n4197), .Z(n4163) );
  ND2I U4007 ( .A(n4168), .B(n4167), .Z(n4169) );
  AN2I U4008 ( .A(n4170), .B(n4169), .Z(rd_data2[20]) );
  B5IP U4009 ( .A(wr_data[21]), .Z(n4171) );
  MUX21L U4010 ( .A(n5397), .B(n4171), .S(n4598), .Z(n2440) );
  MUX21L U4011 ( .A(n5706), .B(n4171), .S(n4604), .Z(n2472) );
  MUX21L U4012 ( .A(n5398), .B(n4171), .S(n4599), .Z(n2600) );
  MUX21L U4013 ( .A(n5399), .B(n4171), .S(n4535), .Z(n2504) );
  MUX21L U4014 ( .A(n4869), .B(n4171), .S(n4602), .Z(n2408) );
  MUX21L U4015 ( .A(n5400), .B(n4171), .S(n4603), .Z(n2536) );
  MUX21L U4016 ( .A(n5401), .B(n4171), .S(n4601), .Z(n2568) );
  MUX21L U4017 ( .A(n5402), .B(n4171), .S(n4605), .Z(n2376) );
  MUX21L U4018 ( .A(n5403), .B(n4171), .S(n4590), .Z(n2696) );
  MUX21L U4019 ( .A(n4868), .B(n4171), .S(n4591), .Z(n2728) );
  MUX21L U4020 ( .A(n5404), .B(n4171), .S(n4537), .Z(n2760) );
  MUX21L U4021 ( .A(n5405), .B(n4171), .S(n4593), .Z(n2824) );
  MUX21L U4022 ( .A(n5406), .B(n4171), .S(n4538), .Z(n2664) );
  MUX21L U4023 ( .A(n5407), .B(n4171), .S(n4595), .Z(n2792) );
  MUX21L U4024 ( .A(n5408), .B(n4171), .S(n4596), .Z(n2856) );
  MUX21L U4025 ( .A(n5409), .B(n4171), .S(n4536), .Z(n2632) );
  MUX21L U4026 ( .A(n5410), .B(n4171), .S(n4606), .Z(n2984) );
  MUX21L U4027 ( .A(n5411), .B(n4171), .S(n4607), .Z(n3112) );
  MUX21L U4028 ( .A(n5412), .B(n4171), .S(n4539), .Z(n3016) );
  MUX21L U4029 ( .A(n5413), .B(n4171), .S(n4609), .Z(n3080) );
  MUX21L U4030 ( .A(n4821), .B(n4171), .S(n4610), .Z(n2920) );
  MUX21L U4031 ( .A(n5414), .B(n4171), .S(n4611), .Z(n3048) );
  MUX21L U4032 ( .A(n5415), .B(n4171), .S(n4612), .Z(n2888) );
  MUX21L U4033 ( .A(n4793), .B(n4171), .S(n4613), .Z(n2952) );
  MUX21L U4034 ( .A(n5416), .B(n4171), .S(n4614), .Z(n3240) );
  MUX21L U4035 ( .A(n5417), .B(n4171), .S(n4540), .Z(n3304) );
  MUX21L U4036 ( .A(n5418), .B(n4171), .S(n4616), .Z(n3144) );
  MUX21L U4037 ( .A(n5419), .B(n4171), .S(n4617), .Z(n3176) );
  MUX21L U4038 ( .A(n5420), .B(n4171), .S(n4618), .Z(n3208) );
  MUX21L U4039 ( .A(n5421), .B(n4171), .S(n4619), .Z(n3336) );
  MUX21L U4040 ( .A(n5422), .B(n4171), .S(n4620), .Z(n3272) );
  AO2 U4041 ( .A(\gpr[26][21] ), .B(n4622), .C(\gpr[24][21] ), .D(n4432), .Z(
        n4177) );
  AO2 U4042 ( .A(\gpr[28][21] ), .B(n4498), .C(\gpr[27][21] ), .D(n4635), .Z(
        n4176) );
  AO2 U4043 ( .A(\gpr[29][21] ), .B(n4639), .C(\gpr[31][21] ), .D(n4548), .Z(
        n4175) );
  ND2I U4044 ( .A(\gpr[30][21] ), .B(n4625), .Z(n4173) );
  ND2I U4045 ( .A(\gpr[25][21] ), .B(n4636), .Z(n4172) );
  AN3 U4046 ( .A(n4453), .B(n4173), .C(n4172), .Z(n4174) );
  ND4 U4047 ( .A(n4177), .B(n4176), .C(n4175), .D(n4174), .Z(n4183) );
  AO2 U4048 ( .A(\gpr[18][21] ), .B(n4487), .C(\gpr[19][21] ), .D(n4635), .Z(
        n4181) );
  AO2 U4049 ( .A(\gpr[17][21] ), .B(n4296), .C(\gpr[20][21] ), .D(n4624), .Z(
        n4180) );
  AO2 U4050 ( .A(\gpr[21][21] ), .B(n4639), .C(\gpr[23][21] ), .D(n4638), .Z(
        n4179) );
  ND4 U4051 ( .A(n4181), .B(n4180), .C(n4179), .D(n4178), .Z(n4182) );
  AN2I U4052 ( .A(n4183), .B(n4182), .Z(n4207) );
  ND2I U4053 ( .A(n4793), .B(n4184), .Z(n4185) );
  AO3 U4054 ( .A(\gpr[15][21] ), .B(n4639), .C(n4652), .D(n4185), .Z(n4186) );
  AO3 U4055 ( .A(n4821), .B(n4108), .C(n4561), .D(n4186), .Z(n4192) );
  ND2I U4056 ( .A(\gpr[3][21] ), .B(n4557), .Z(n4190) );
  ND2I U4057 ( .A(\gpr[5][21] ), .B(n4658), .Z(n4189) );
  ND2I U4058 ( .A(\gpr[1][21] ), .B(n4556), .Z(n4188) );
  ND2I U4059 ( .A(\gpr[4][21] ), .B(n4666), .Z(n4187) );
  ND4 U4060 ( .A(n4190), .B(n4189), .C(n4188), .D(n4187), .Z(n4191) );
  NR2I U4061 ( .A(n4192), .B(n4191), .Z(n4205) );
  ND2I U4062 ( .A(\gpr[2][21] ), .B(n4659), .Z(n4196) );
  ND2I U4063 ( .A(\gpr[10][21] ), .B(n4268), .Z(n4195) );
  ND2I U4064 ( .A(\gpr[9][21] ), .B(n4668), .Z(n4194) );
  ND2I U4065 ( .A(\gpr[8][21] ), .B(n4519), .Z(n4193) );
  ND4 U4066 ( .A(n4196), .B(n4195), .C(n4194), .D(n4193), .Z(n4203) );
  ND2I U4067 ( .A(\gpr[11][21] ), .B(n4571), .Z(n4201) );
  ND2I U4068 ( .A(\gpr[12][21] ), .B(n4573), .Z(n4200) );
  ND2I U4069 ( .A(\gpr[7][21] ), .B(n4675), .Z(n4199) );
  ND2I U4070 ( .A(\gpr[6][21] ), .B(n4197), .Z(n4198) );
  ND4 U4071 ( .A(n4201), .B(n4200), .C(n4199), .D(n4198), .Z(n4202) );
  NR2I U4072 ( .A(n4203), .B(n4202), .Z(n4204) );
  ND2I U4073 ( .A(n4205), .B(n4204), .Z(n4206) );
  AN2I U4074 ( .A(n4207), .B(n4206), .Z(rd_data2[21]) );
  B4IP U4075 ( .A(wr_data[22]), .Z(n4208) );
  MUX21L U4076 ( .A(n5423), .B(n4208), .S(n4536), .Z(n2633) );
  MUX21L U4077 ( .A(n5424), .B(n4208), .S(n4590), .Z(n2697) );
  MUX21L U4078 ( .A(n5425), .B(n4208), .S(n4591), .Z(n2729) );
  MUX21L U4079 ( .A(n5426), .B(n4208), .S(n4592), .Z(n2761) );
  MUX21L U4080 ( .A(n4870), .B(n4208), .S(n4538), .Z(n2665) );
  MUX21L U4081 ( .A(n5427), .B(n4208), .S(n4595), .Z(n2793) );
  MUX21L U4082 ( .A(n5428), .B(n4208), .S(n4596), .Z(n2857) );
  MUX21L U4083 ( .A(n5429), .B(n4208), .S(n4593), .Z(n2825) );
  MUX21L U4084 ( .A(n5430), .B(n4208), .S(n4598), .Z(n2441) );
  MUX21L U4085 ( .A(n5431), .B(n4208), .S(n4604), .Z(n2473) );
  MUX21L U4086 ( .A(n5432), .B(n4208), .S(n4599), .Z(n2601) );
  MUX21L U4087 ( .A(n5433), .B(n4208), .S(n4600), .Z(n2505) );
  MUX21L U4088 ( .A(n4871), .B(n4208), .S(n4602), .Z(n2409) );
  MUX21L U4089 ( .A(n5434), .B(n4208), .S(n4603), .Z(n2537) );
  MUX21L U4090 ( .A(n5435), .B(n4208), .S(n4601), .Z(n2569) );
  MUX21L U4091 ( .A(n5436), .B(n4208), .S(n4605), .Z(n2377) );
  MUX21L U4092 ( .A(n5437), .B(n4208), .S(n4606), .Z(n2985) );
  MUX21L U4093 ( .A(n5438), .B(n4208), .S(n4607), .Z(n3113) );
  MUX21L U4094 ( .A(n5707), .B(n4208), .S(n4608), .Z(n3017) );
  MUX21L U4095 ( .A(n5708), .B(n4208), .S(n4609), .Z(n3081) );
  MUX21L U4096 ( .A(n4822), .B(n4208), .S(n4610), .Z(n2921) );
  MUX21L U4097 ( .A(n5439), .B(n4208), .S(n4611), .Z(n3049) );
  MUX21L U4098 ( .A(n5440), .B(n4208), .S(n4612), .Z(n2889) );
  MUX21L U4099 ( .A(n4794), .B(n4208), .S(n4613), .Z(n2953) );
  MUX21L U4100 ( .A(n5441), .B(n4208), .S(n4614), .Z(n3241) );
  MUX21L U4101 ( .A(n5442), .B(n4208), .S(n4540), .Z(n3305) );
  MUX21L U4102 ( .A(n5709), .B(n4208), .S(n4616), .Z(n3145) );
  MUX21L U4103 ( .A(n5710), .B(n4208), .S(n4617), .Z(n3177) );
  MUX21L U4104 ( .A(n5711), .B(n4208), .S(n4618), .Z(n3209) );
  MUX21L U4105 ( .A(n5712), .B(n4208), .S(n4619), .Z(n3337) );
  MUX21L U4106 ( .A(n5713), .B(n4208), .S(n4620), .Z(n3273) );
  AO2 U4107 ( .A(\gpr[17][22] ), .B(n4296), .C(\gpr[18][22] ), .D(n4214), .Z(
        n4213) );
  AO2 U4108 ( .A(\gpr[19][22] ), .B(n4635), .C(\gpr[20][22] ), .D(n4624), .Z(
        n4212) );
  AO2 U4109 ( .A(\gpr[21][22] ), .B(n4639), .C(\gpr[22][22] ), .D(n4431), .Z(
        n4211) );
  ND4 U4110 ( .A(n4213), .B(n4212), .C(n4211), .D(n4210), .Z(n4222) );
  AO2 U4111 ( .A(\gpr[26][22] ), .B(n4214), .C(\gpr[24][22] ), .D(n4626), .Z(
        n4220) );
  AO2 U4112 ( .A(\gpr[27][22] ), .B(n4635), .C(\gpr[28][22] ), .D(n4498), .Z(
        n4219) );
  AO2 U4113 ( .A(\gpr[29][22] ), .B(n4639), .C(\gpr[31][22] ), .D(n4333), .Z(
        n4218) );
  ND2I U4114 ( .A(\gpr[30][22] ), .B(n4625), .Z(n4216) );
  ND2I U4115 ( .A(\gpr[25][22] ), .B(n4636), .Z(n4215) );
  AN3 U4116 ( .A(n4453), .B(n4216), .C(n4215), .Z(n4217) );
  ND4 U4117 ( .A(n4220), .B(n4219), .C(n4218), .D(n4217), .Z(n4221) );
  AN2I U4118 ( .A(n4222), .B(n4221), .Z(n4245) );
  IVI U4119 ( .A(n4223), .Z(n4650) );
  ND2I U4120 ( .A(n4794), .B(n4650), .Z(n4224) );
  AO3 U4121 ( .A(\gpr[15][22] ), .B(n4639), .C(n4652), .D(n4224), .Z(n4225) );
  AO3 U4122 ( .A(n4822), .B(n4108), .C(n4561), .D(n4225), .Z(n4231) );
  ND2I U4123 ( .A(\gpr[3][22] ), .B(n4557), .Z(n4229) );
  ND2I U4124 ( .A(\gpr[5][22] ), .B(n4658), .Z(n4228) );
  ND2I U4125 ( .A(\gpr[1][22] ), .B(n4556), .Z(n4227) );
  ND2I U4126 ( .A(\gpr[4][22] ), .B(n4666), .Z(n4226) );
  ND4 U4127 ( .A(n4229), .B(n4228), .C(n4227), .D(n4226), .Z(n4230) );
  NR2I U4128 ( .A(n4231), .B(n4230), .Z(n4243) );
  ND2I U4129 ( .A(\gpr[2][22] ), .B(n4659), .Z(n4235) );
  ND2I U4130 ( .A(n4562), .B(\gpr[10][22] ), .Z(n4234) );
  ND2I U4131 ( .A(\gpr[9][22] ), .B(n4518), .Z(n4233) );
  ND2I U4132 ( .A(\gpr[8][22] ), .B(n3960), .Z(n4232) );
  ND4 U4133 ( .A(n4235), .B(n4234), .C(n4233), .D(n4232), .Z(n4241) );
  ND2I U4134 ( .A(\gpr[11][22] ), .B(n4667), .Z(n4239) );
  ND2I U4135 ( .A(\gpr[12][22] ), .B(n4673), .Z(n4238) );
  ND2I U4136 ( .A(\gpr[7][22] ), .B(n4675), .Z(n4237) );
  ND2I U4137 ( .A(\gpr[6][22] ), .B(n4354), .Z(n4236) );
  ND4 U4138 ( .A(n4239), .B(n4238), .C(n4237), .D(n4236), .Z(n4240) );
  NR2I U4139 ( .A(n4241), .B(n4240), .Z(n4242) );
  ND2I U4140 ( .A(n4243), .B(n4242), .Z(n4244) );
  AN2I U4141 ( .A(n4245), .B(n4244), .Z(rd_data2[22]) );
  B4IP U4142 ( .A(wr_data[23]), .Z(n4246) );
  MUX21L U4143 ( .A(n5443), .B(n4246), .S(n4605), .Z(n2378) );
  MUX21L U4144 ( .A(n5444), .B(n4246), .S(n4598), .Z(n2442) );
  MUX21L U4145 ( .A(n5445), .B(n4246), .S(n4600), .Z(n2506) );
  MUX21L U4146 ( .A(n4873), .B(n4246), .S(n4602), .Z(n2410) );
  MUX21L U4147 ( .A(n5446), .B(n4246), .S(n4603), .Z(n2538) );
  MUX21L U4148 ( .A(n5714), .B(n4246), .S(n4599), .Z(n2602) );
  MUX21L U4149 ( .A(n5447), .B(n4246), .S(n4601), .Z(n2570) );
  MUX21L U4150 ( .A(n5448), .B(n4246), .S(n4536), .Z(n2634) );
  MUX21L U4151 ( .A(n5449), .B(n4246), .S(n4590), .Z(n2698) );
  MUX21L U4152 ( .A(n5450), .B(n4246), .S(n4596), .Z(n2858) );
  MUX21L U4153 ( .A(n4872), .B(n4246), .S(n4538), .Z(n2666) );
  MUX21L U4154 ( .A(n5451), .B(n4246), .S(n4595), .Z(n2794) );
  MUX21L U4155 ( .A(n5452), .B(n4246), .S(n4593), .Z(n2826) );
  MUX21L U4156 ( .A(n5453), .B(n4246), .S(n4592), .Z(n2762) );
  MUX21L U4157 ( .A(n5454), .B(n4246), .S(n4606), .Z(n2986) );
  MUX21L U4158 ( .A(n5455), .B(n4246), .S(n4607), .Z(n3114) );
  MUX21L U4159 ( .A(n5456), .B(n4246), .S(n4608), .Z(n3018) );
  MUX21L U4160 ( .A(n5457), .B(n4246), .S(n4609), .Z(n3082) );
  MUX21L U4161 ( .A(n4823), .B(n4246), .S(n4610), .Z(n2922) );
  MUX21L U4162 ( .A(n5458), .B(n4246), .S(n4611), .Z(n3050) );
  MUX21L U4163 ( .A(n5459), .B(n4246), .S(n4612), .Z(n2890) );
  MUX21L U4164 ( .A(n4795), .B(n4246), .S(n4613), .Z(n2954) );
  MUX21L U4165 ( .A(n5460), .B(n4246), .S(n4614), .Z(n3242) );
  MUX21L U4166 ( .A(n5461), .B(n4246), .S(n4540), .Z(n3306) );
  MUX21L U4167 ( .A(n5462), .B(n4246), .S(n4616), .Z(n3146) );
  MUX21L U4168 ( .A(n5463), .B(n4246), .S(n4617), .Z(n3178) );
  MUX21L U4169 ( .A(n5464), .B(n4246), .S(n4618), .Z(n3210) );
  MUX21L U4170 ( .A(n5465), .B(n4246), .S(n4619), .Z(n3338) );
  MUX21L U4171 ( .A(n5466), .B(n4246), .S(n4620), .Z(n3274) );
  AO2 U4172 ( .A(\gpr[25][23] ), .B(n4296), .C(\gpr[26][23] ), .D(n4622), .Z(
        n4250) );
  AO2 U4173 ( .A(\gpr[27][23] ), .B(n4635), .C(\gpr[28][23] ), .D(n4498), .Z(
        n4249) );
  AO2 U4174 ( .A(\gpr[29][23] ), .B(n4639), .C(\gpr[30][23] ), .D(n4431), .Z(
        n4248) );
  ND4 U4175 ( .A(n4250), .B(n4249), .C(n4248), .D(n4247), .Z(n4259) );
  AO2 U4176 ( .A(\gpr[18][23] ), .B(n4458), .C(\gpr[19][23] ), .D(n4635), .Z(
        n4257) );
  AO2 U4177 ( .A(\gpr[20][23] ), .B(n4624), .C(\gpr[16][23] ), .D(n4542), .Z(
        n4256) );
  AO2 U4178 ( .A(\gpr[21][23] ), .B(n4639), .C(\gpr[22][23] ), .D(n4431), .Z(
        n4255) );
  ND2I U4179 ( .A(\gpr[23][23] ), .B(n4251), .Z(n4253) );
  ND2I U4180 ( .A(\gpr[17][23] ), .B(n4636), .Z(n4252) );
  AN3 U4181 ( .A(n4628), .B(n4253), .C(n4252), .Z(n4254) );
  ND4 U4182 ( .A(n4257), .B(n4256), .C(n4255), .D(n4254), .Z(n4258) );
  AN2I U4183 ( .A(n4259), .B(n4258), .Z(n4282) );
  ND2I U4184 ( .A(n4795), .B(n4650), .Z(n4260) );
  AO3 U4185 ( .A(\gpr[15][23] ), .B(n4639), .C(n4652), .D(n4260), .Z(n4261) );
  AO3 U4186 ( .A(n4823), .B(n4466), .C(n4561), .D(n4261), .Z(n4267) );
  ND2I U4187 ( .A(\gpr[3][23] ), .B(n4557), .Z(n4265) );
  ND2I U4188 ( .A(\gpr[5][23] ), .B(n4658), .Z(n4264) );
  ND2I U4189 ( .A(\gpr[1][23] ), .B(n4556), .Z(n4263) );
  ND2I U4190 ( .A(\gpr[4][23] ), .B(n4666), .Z(n4262) );
  ND4 U4191 ( .A(n4265), .B(n4264), .C(n4263), .D(n4262), .Z(n4266) );
  NR2I U4192 ( .A(n4267), .B(n4266), .Z(n4280) );
  ND2I U4193 ( .A(\gpr[2][23] ), .B(n4659), .Z(n4272) );
  ND2I U4194 ( .A(\gpr[10][23] ), .B(n4268), .Z(n4271) );
  ND2I U4195 ( .A(\gpr[9][23] ), .B(n4563), .Z(n4270) );
  ND2I U4196 ( .A(\gpr[8][23] ), .B(n4519), .Z(n4269) );
  ND4 U4197 ( .A(n4272), .B(n4271), .C(n4270), .D(n4269), .Z(n4278) );
  ND2I U4198 ( .A(\gpr[11][23] ), .B(n4667), .Z(n4276) );
  ND2I U4199 ( .A(\gpr[12][23] ), .B(n4673), .Z(n4275) );
  ND2I U4200 ( .A(\gpr[7][23] ), .B(n4675), .Z(n4274) );
  ND2I U4201 ( .A(\gpr[6][23] ), .B(n4354), .Z(n4273) );
  ND4 U4202 ( .A(n4276), .B(n4275), .C(n4274), .D(n4273), .Z(n4277) );
  NR2I U4203 ( .A(n4278), .B(n4277), .Z(n4279) );
  ND2I U4204 ( .A(n4280), .B(n4279), .Z(n4281) );
  AN2I U4205 ( .A(n4282), .B(n4281), .Z(rd_data2[23]) );
  B4IP U4206 ( .A(wr_data[24]), .Z(n4283) );
  MUX21L U4207 ( .A(n5467), .B(n4283), .S(n4598), .Z(n2443) );
  MUX21L U4208 ( .A(n5468), .B(n4283), .S(n4604), .Z(n2475) );
  MUX21L U4209 ( .A(n5469), .B(n4283), .S(n4599), .Z(n2603) );
  MUX21L U4210 ( .A(n5470), .B(n4283), .S(n4600), .Z(n2507) );
  MUX21L U4211 ( .A(n5471), .B(n4283), .S(n4602), .Z(n2411) );
  MUX21L U4212 ( .A(n5472), .B(n4283), .S(n4603), .Z(n2539) );
  MUX21L U4213 ( .A(n5473), .B(n4283), .S(n4601), .Z(n2571) );
  MUX21L U4214 ( .A(n4808), .B(n4283), .S(n4605), .Z(n2379) );
  MUX21L U4215 ( .A(n4776), .B(n4283), .S(n4590), .Z(n2699) );
  MUX21L U4216 ( .A(n5474), .B(n4283), .S(n4591), .Z(n2731) );
  MUX21L U4217 ( .A(n5475), .B(n4283), .S(n4592), .Z(n2763) );
  MUX21L U4218 ( .A(n5476), .B(n4283), .S(n4593), .Z(n2827) );
  MUX21L U4219 ( .A(n5477), .B(n4283), .S(n4538), .Z(n2667) );
  MUX21L U4220 ( .A(n5478), .B(n4283), .S(n4595), .Z(n2795) );
  MUX21L U4221 ( .A(n5479), .B(n4283), .S(n4596), .Z(n2859) );
  MUX21L U4222 ( .A(n5480), .B(n4283), .S(n4597), .Z(n2635) );
  MUX21L U4223 ( .A(n5481), .B(n4283), .S(n4606), .Z(n2987) );
  MUX21L U4224 ( .A(n5482), .B(n4283), .S(n4607), .Z(n3115) );
  MUX21L U4225 ( .A(n5483), .B(n4283), .S(n4608), .Z(n3019) );
  MUX21L U4226 ( .A(n5484), .B(n4283), .S(n4609), .Z(n3083) );
  MUX21L U4227 ( .A(n4775), .B(n4283), .S(n4610), .Z(n2923) );
  MUX21L U4228 ( .A(n5485), .B(n4283), .S(n4611), .Z(n3051) );
  MUX21L U4229 ( .A(n5486), .B(n4283), .S(n4612), .Z(n2891) );
  MUX21L U4230 ( .A(n4769), .B(n4283), .S(n4613), .Z(n2955) );
  MUX21L U4231 ( .A(n5487), .B(n4283), .S(n4614), .Z(n3243) );
  MUX21L U4232 ( .A(n5488), .B(n4283), .S(n4615), .Z(n3307) );
  MUX21L U4233 ( .A(n5489), .B(n4283), .S(n4616), .Z(n3147) );
  MUX21L U4234 ( .A(n5490), .B(n4283), .S(n4617), .Z(n3179) );
  MUX21L U4235 ( .A(n5491), .B(n4283), .S(n4618), .Z(n3211) );
  MUX21L U4236 ( .A(n5492), .B(n4283), .S(n4619), .Z(n3339) );
  MUX21L U4237 ( .A(n5493), .B(n4283), .S(n4620), .Z(n3275) );
  AO2 U4238 ( .A(\gpr[24][24] ), .B(n4432), .C(\gpr[26][24] ), .D(n4293), .Z(
        n4292) );
  ND2I U4239 ( .A(\gpr[27][24] ), .B(n4623), .Z(n4285) );
  ND2I U4240 ( .A(n219), .B(\gpr[28][24] ), .Z(n4284) );
  AN2I U4241 ( .A(n4285), .B(n4284), .Z(n4291) );
  AO2 U4242 ( .A(\gpr[29][24] ), .B(n4639), .C(\gpr[31][24] ), .D(n4488), .Z(
        n4290) );
  ND2I U4243 ( .A(\gpr[30][24] ), .B(n4625), .Z(n4288) );
  ND2I U4244 ( .A(\gpr[25][24] ), .B(n4286), .Z(n4287) );
  AN3 U4245 ( .A(n4453), .B(n4288), .C(n4287), .Z(n4289) );
  ND4 U4246 ( .A(n4292), .B(n4291), .C(n4290), .D(n4289), .Z(n4305) );
  ND2I U4247 ( .A(\gpr[19][24] ), .B(n4623), .Z(n4295) );
  ND2I U4248 ( .A(n4293), .B(\gpr[18][24] ), .Z(n4294) );
  AN2I U4249 ( .A(n4295), .B(n4294), .Z(n4303) );
  AO2 U4250 ( .A(\gpr[17][24] ), .B(n4296), .C(\gpr[20][24] ), .D(n219), .Z(
        n4302) );
  AO2 U4251 ( .A(\gpr[23][24] ), .B(n4499), .C(\gpr[21][24] ), .D(n4639), .Z(
        n4301) );
  AN2I U4252 ( .A(\gpr[22][24] ), .B(n4625), .Z(n4299) );
  ND2I U4253 ( .A(\gpr[16][24] ), .B(n4542), .Z(n4297) );
  ND2I U4254 ( .A(n4628), .B(n4297), .Z(n4298) );
  NR2I U4255 ( .A(n4299), .B(n4298), .Z(n4300) );
  ND4 U4256 ( .A(n4303), .B(n4302), .C(n4301), .D(n4300), .Z(n4304) );
  AN2I U4257 ( .A(n4305), .B(n4304), .Z(n4331) );
  ND2I U4258 ( .A(n4769), .B(n4650), .Z(n4306) );
  AO3 U4259 ( .A(\gpr[15][24] ), .B(n4639), .C(n4652), .D(n4306), .Z(n4307) );
  ND2I U4260 ( .A(\gpr[3][24] ), .B(n4557), .Z(n4312) );
  ND2I U4261 ( .A(\gpr[5][24] ), .B(n4658), .Z(n4311) );
  ND2I U4262 ( .A(\gpr[1][24] ), .B(n4556), .Z(n4310) );
  ND2I U4263 ( .A(\gpr[4][24] ), .B(n4308), .Z(n4309) );
  ND2I U4264 ( .A(\gpr[2][24] ), .B(n4659), .Z(n4319) );
  ND2I U4265 ( .A(\gpr[10][24] ), .B(n4313), .Z(n4318) );
  ND2I U4266 ( .A(\gpr[9][24] ), .B(n4314), .Z(n4317) );
  ND2I U4267 ( .A(\gpr[8][24] ), .B(n4315), .Z(n4316) );
  ND4 U4268 ( .A(n4319), .B(n4318), .C(n4317), .D(n4316), .Z(n4327) );
  ND2I U4269 ( .A(\gpr[11][24] ), .B(n4320), .Z(n4325) );
  ND2I U4270 ( .A(\gpr[12][24] ), .B(n4321), .Z(n4324) );
  ND2I U4271 ( .A(\gpr[7][24] ), .B(n4675), .Z(n4323) );
  ND2I U4272 ( .A(\gpr[6][24] ), .B(n4354), .Z(n4322) );
  ND4 U4273 ( .A(n4325), .B(n4324), .C(n4323), .D(n4322), .Z(n4326) );
  NR2I U4274 ( .A(n4327), .B(n4326), .Z(n4328) );
  ND2I U4275 ( .A(n4329), .B(n4328), .Z(n4330) );
  AN2I U4276 ( .A(n4331), .B(n4330), .Z(rd_data2[24]) );
  B4IP U4277 ( .A(wr_data[25]), .Z(n4332) );
  MUX21L U4278 ( .A(n314), .B(n4332), .S(n4604), .Z(n2476) );
  MUX21L U4279 ( .A(n5494), .B(n4332), .S(n4600), .Z(n2508) );
  MUX21L U4280 ( .A(n5495), .B(n4332), .S(n4605), .Z(n2380) );
  MUX21L U4281 ( .A(n5496), .B(n4332), .S(n4598), .Z(n2444) );
  MUX21L U4282 ( .A(n5497), .B(n4332), .S(n4599), .Z(n2604) );
  MUX21L U4283 ( .A(n5498), .B(n4332), .S(n4601), .Z(n2572) );
  MUX21L U4284 ( .A(n4874), .B(n4332), .S(n4602), .Z(n2412) );
  MUX21L U4285 ( .A(n4797), .B(n4332), .S(n4603), .Z(n2540) );
  MUX21L U4286 ( .A(n5499), .B(n4332), .S(n4612), .Z(n2892) );
  MUX21L U4287 ( .A(n4798), .B(n4332), .S(n4613), .Z(n2956) );
  MUX21L U4288 ( .A(n5500), .B(n4332), .S(n4616), .Z(n3148) );
  MUX21L U4289 ( .A(n5501), .B(n4332), .S(n4617), .Z(n3180) );
  MUX21L U4290 ( .A(n5502), .B(n4332), .S(n4618), .Z(n3212) );
  MUX21L U4291 ( .A(n5503), .B(n4332), .S(n4606), .Z(n2988) );
  MUX21L U4292 ( .A(n315), .B(n4332), .S(n4607), .Z(n3116) );
  MUX21L U4293 ( .A(n5504), .B(n4332), .S(n4608), .Z(n3020) );
  MUX21L U4294 ( .A(n5505), .B(n4332), .S(n4609), .Z(n3084) );
  MUX21L U4295 ( .A(n5506), .B(n4332), .S(n4610), .Z(n2924) );
  MUX21L U4296 ( .A(n4799), .B(n4332), .S(n4611), .Z(n3052) );
  MUX21L U4297 ( .A(n5507), .B(n4332), .S(n4614), .Z(n3244) );
  MUX21L U4298 ( .A(n5508), .B(n4332), .S(n4540), .Z(n3308) );
  MUX21L U4299 ( .A(n5509), .B(n4332), .S(n4619), .Z(n3340) );
  MUX21L U4300 ( .A(n5510), .B(n4332), .S(n4620), .Z(n3276) );
  MUX21L U4301 ( .A(n5511), .B(n4332), .S(n4536), .Z(n2636) );
  MUX21L U4302 ( .A(n5512), .B(n4332), .S(n4590), .Z(n2700) );
  MUX21L U4303 ( .A(n316), .B(n4332), .S(n4591), .Z(n2732) );
  MUX21L U4304 ( .A(n5513), .B(n4332), .S(n4596), .Z(n2860) );
  MUX21L U4305 ( .A(n5514), .B(n4332), .S(n4592), .Z(n2764) );
  MUX21L U4306 ( .A(n5515), .B(n4332), .S(n4593), .Z(n2828) );
  MUX21L U4307 ( .A(n4875), .B(n4332), .S(n4538), .Z(n2668) );
  MUX21L U4308 ( .A(n4796), .B(n4332), .S(n4595), .Z(n2796) );
  AO2 U4309 ( .A(\gpr[19][25] ), .B(n4635), .C(\gpr[17][25] ), .D(n4636), .Z(
        n4339) );
  AO2 U4310 ( .A(\gpr[16][25] ), .B(n4626), .C(\gpr[20][25] ), .D(n4498), .Z(
        n4338) );
  AO2 U4311 ( .A(\gpr[21][25] ), .B(n4639), .C(\gpr[22][25] ), .D(n4431), .Z(
        n4337) );
  ND2I U4312 ( .A(\gpr[23][25] ), .B(n4333), .Z(n4334) );
  AO3 U4313 ( .A(n4356), .B(n4796), .C(n4628), .D(n4334), .Z(n4335) );
  IVI U4314 ( .A(n4335), .Z(n4336) );
  ND4 U4315 ( .A(n4339), .B(n4338), .C(n4337), .D(n4336), .Z(n4346) );
  ND2I U4316 ( .A(\gpr[27][25] ), .B(n4623), .Z(n4341) );
  ND2I U4317 ( .A(n4639), .B(\gpr[29][25] ), .Z(n4340) );
  ND2I U4318 ( .A(\gpr[31][25] ), .B(n4342), .Z(n4343) );
  AO3 U4319 ( .A(n4356), .B(n4797), .C(n4641), .D(n4343), .Z(n4344) );
  AN2I U4320 ( .A(n4346), .B(n4345), .Z(n4370) );
  ND2I U4321 ( .A(\gpr[1][25] ), .B(n4556), .Z(n4349) );
  ND2I U4322 ( .A(n4798), .B(n4650), .Z(n4347) );
  AO3 U4323 ( .A(\gpr[15][25] ), .B(n4639), .C(n4652), .D(n4347), .Z(n4348) );
  ND2I U4324 ( .A(n4349), .B(n4348), .Z(n4353) );
  ND2I U4325 ( .A(\gpr[3][25] ), .B(n4557), .Z(n4351) );
  ND2I U4326 ( .A(\gpr[4][25] ), .B(n4666), .Z(n4350) );
  ND2I U4327 ( .A(n4351), .B(n4350), .Z(n4352) );
  NR2I U4328 ( .A(n4353), .B(n4352), .Z(n4368) );
  AO2 U4329 ( .A(\gpr[2][25] ), .B(n4659), .C(\gpr[5][25] ), .D(n4658), .Z(
        n4367) );
  AO2 U4330 ( .A(\gpr[6][25] ), .B(n4354), .C(\gpr[7][25] ), .D(n4675), .Z(
        n4366) );
  ND2I U4331 ( .A(\gpr[14][25] ), .B(n4489), .Z(n4355) );
  AO3 U4332 ( .A(n4799), .B(n4356), .C(n4561), .D(n4355), .Z(n4364) );
  ND2I U4333 ( .A(\gpr[9][25] ), .B(n4636), .Z(n4361) );
  ND2I U4334 ( .A(\gpr[8][25] ), .B(n4357), .Z(n4360) );
  ND2I U4335 ( .A(\gpr[11][25] ), .B(n4501), .Z(n4359) );
  ND2I U4336 ( .A(\gpr[12][25] ), .B(n4624), .Z(n4358) );
  ND4 U4337 ( .A(n4361), .B(n4360), .C(n4359), .D(n4358), .Z(n4363) );
  AO7 U4338 ( .A(n4364), .B(n4363), .C(n4362), .Z(n4365) );
  ND4 U4339 ( .A(n4368), .B(n4367), .C(n4366), .D(n4365), .Z(n4369) );
  AN2I U4340 ( .A(n4370), .B(n4369), .Z(rd_data2[25]) );
  B4IP U4341 ( .A(wr_data[26]), .Z(n4371) );
  MUX21L U4342 ( .A(n5516), .B(n4371), .S(n4605), .Z(n2381) );
  MUX21L U4343 ( .A(n5517), .B(n4371), .S(n4598), .Z(n2445) );
  MUX21L U4344 ( .A(n5518), .B(n4371), .S(n4604), .Z(n2477) );
  MUX21L U4345 ( .A(n5519), .B(n4371), .S(n4599), .Z(n2605) );
  MUX21L U4346 ( .A(n4809), .B(n4371), .S(n4602), .Z(n2413) );
  MUX21L U4347 ( .A(n5520), .B(n4371), .S(n4603), .Z(n2541) );
  MUX21L U4348 ( .A(n5521), .B(n4371), .S(n4601), .Z(n2573) );
  MUX21L U4349 ( .A(n5522), .B(n4371), .S(n4535), .Z(n2509) );
  MUX21L U4350 ( .A(n4876), .B(n4371), .S(n4590), .Z(n2701) );
  MUX21L U4351 ( .A(n5523), .B(n4371), .S(n4591), .Z(n2733) );
  MUX21L U4352 ( .A(n5524), .B(n4371), .S(n4596), .Z(n2861) );
  MUX21L U4353 ( .A(n5525), .B(n4371), .S(n4593), .Z(n2829) );
  MUX21L U4354 ( .A(n5526), .B(n4371), .S(n4538), .Z(n2669) );
  MUX21L U4355 ( .A(n5527), .B(n4371), .S(n4595), .Z(n2797) );
  MUX21L U4356 ( .A(n5528), .B(n4371), .S(n4537), .Z(n2765) );
  MUX21L U4357 ( .A(n5529), .B(n4371), .S(n4597), .Z(n2637) );
  MUX21L U4358 ( .A(n5715), .B(n4371), .S(n4606), .Z(n2989) );
  MUX21L U4359 ( .A(n5530), .B(n4371), .S(n4607), .Z(n3117) );
  MUX21L U4360 ( .A(n5531), .B(n4371), .S(n4539), .Z(n3021) );
  MUX21L U4361 ( .A(n5532), .B(n4371), .S(n4609), .Z(n3085) );
  MUX21L U4362 ( .A(n5533), .B(n4371), .S(n4610), .Z(n2925) );
  MUX21L U4363 ( .A(n5534), .B(n4371), .S(n4611), .Z(n3053) );
  MUX21L U4364 ( .A(n5535), .B(n4371), .S(n4612), .Z(n2893) );
  MUX21L U4365 ( .A(n4800), .B(n4371), .S(n4613), .Z(n2957) );
  MUX21L U4366 ( .A(n5536), .B(n4371), .S(n4615), .Z(n3309) );
  MUX21L U4367 ( .A(n5537), .B(n4371), .S(n4616), .Z(n3149) );
  MUX21L U4368 ( .A(n5538), .B(n4371), .S(n4617), .Z(n3181) );
  MUX21L U4369 ( .A(n5539), .B(n4371), .S(n4618), .Z(n3213) );
  MUX21L U4370 ( .A(n5540), .B(n4371), .S(n4619), .Z(n3341) );
  MUX21L U4371 ( .A(n5541), .B(n4371), .S(n4620), .Z(n3277) );
  ND2I U4372 ( .A(\gpr[27][26] ), .B(n4623), .Z(n4373) );
  ND2I U4373 ( .A(n4487), .B(\gpr[26][26] ), .Z(n4372) );
  AN2I U4374 ( .A(n4373), .B(n4372), .Z(n4380) );
  AO2 U4375 ( .A(\gpr[28][26] ), .B(n4624), .C(\gpr[24][26] ), .D(n4432), .Z(
        n4379) );
  AO2 U4376 ( .A(\gpr[29][26] ), .B(n4639), .C(\gpr[30][26] ), .D(n4431), .Z(
        n4378) );
  ND2I U4377 ( .A(\gpr[31][26] ), .B(n4374), .Z(n4376) );
  ND2I U4378 ( .A(\gpr[25][26] ), .B(n4636), .Z(n4375) );
  AN3 U4379 ( .A(n4453), .B(n4376), .C(n4375), .Z(n4377) );
  ND4 U4380 ( .A(n4380), .B(n4379), .C(n4378), .D(n4377), .Z(n4389) );
  AO2 U4381 ( .A(\gpr[18][26] ), .B(n4458), .C(\gpr[16][26] ), .D(n4626), .Z(
        n4387) );
  AO2 U4382 ( .A(\gpr[17][26] ), .B(n4636), .C(\gpr[20][26] ), .D(n4624), .Z(
        n4386) );
  AO2 U4383 ( .A(\gpr[23][26] ), .B(n4543), .C(\gpr[21][26] ), .D(n4639), .Z(
        n4385) );
  AN2I U4384 ( .A(\gpr[22][26] ), .B(n4625), .Z(n4383) );
  ND2I U4385 ( .A(\gpr[19][26] ), .B(n4501), .Z(n4381) );
  ND2I U4386 ( .A(n4628), .B(n4381), .Z(n4382) );
  NR2I U4387 ( .A(n4383), .B(n4382), .Z(n4384) );
  ND4 U4388 ( .A(n4387), .B(n4386), .C(n4385), .D(n4384), .Z(n4388) );
  AN2I U4389 ( .A(n4389), .B(n4388), .Z(n4411) );
  ND2I U4390 ( .A(\gpr[6][26] ), .B(n4524), .Z(n4392) );
  ND2I U4391 ( .A(n4800), .B(n4650), .Z(n4390) );
  AO3 U4392 ( .A(\gpr[15][26] ), .B(n4639), .C(n4652), .D(n4390), .Z(n4391) );
  AN3 U4393 ( .A(n4561), .B(n4392), .C(n4391), .Z(n4409) );
  AO2 U4394 ( .A(\gpr[2][26] ), .B(n4659), .C(\gpr[7][26] ), .D(n4675), .Z(
        n4408) );
  AO2 U4395 ( .A(\gpr[1][26] ), .B(n4656), .C(\gpr[3][26] ), .D(n4657), .Z(
        n4396) );
  ND2I U4396 ( .A(\gpr[4][26] ), .B(n4153), .Z(n4394) );
  ND2I U4397 ( .A(n4658), .B(\gpr[5][26] ), .Z(n4393) );
  AN2I U4398 ( .A(n4394), .B(n4393), .Z(n4395) );
  AN2I U4399 ( .A(n4396), .B(n4395), .Z(n4407) );
  AO2 U4400 ( .A(\gpr[8][26] ), .B(n4450), .C(\gpr[14][26] ), .D(n4431), .Z(
        n4404) );
  ND2I U4401 ( .A(\gpr[10][26] ), .B(n4487), .Z(n4398) );
  ND2I U4402 ( .A(\gpr[9][26] ), .B(n4636), .Z(n4397) );
  ND2I U4403 ( .A(n4398), .B(n4397), .Z(n4402) );
  ND2I U4404 ( .A(\gpr[11][26] ), .B(n4501), .Z(n4400) );
  ND2I U4405 ( .A(\gpr[12][26] ), .B(n4498), .Z(n4399) );
  ND2I U4406 ( .A(n4400), .B(n4399), .Z(n4401) );
  NR2I U4407 ( .A(n4402), .B(n4401), .Z(n4403) );
  ND2I U4408 ( .A(n4404), .B(n4403), .Z(n4405) );
  ND2I U4409 ( .A(n4442), .B(n4405), .Z(n4406) );
  ND4 U4410 ( .A(n4409), .B(n4408), .C(n4407), .D(n4406), .Z(n4410) );
  AN2I U4411 ( .A(n4411), .B(n4410), .Z(rd_data2[26]) );
  B4IP U4412 ( .A(wr_data[27]), .Z(n4412) );
  MUX21L U4413 ( .A(n5542), .B(n4412), .S(n4590), .Z(n2702) );
  MUX21L U4414 ( .A(n4877), .B(n4412), .S(n4591), .Z(n2734) );
  MUX21L U4415 ( .A(n5543), .B(n4412), .S(n4596), .Z(n2862) );
  MUX21L U4416 ( .A(n5544), .B(n4412), .S(n4593), .Z(n2830) );
  MUX21L U4417 ( .A(n5545), .B(n4412), .S(n4538), .Z(n2670) );
  MUX21L U4418 ( .A(n5546), .B(n4412), .S(n4595), .Z(n2798) );
  MUX21L U4419 ( .A(n5547), .B(n4412), .S(n4592), .Z(n2766) );
  MUX21L U4420 ( .A(n5548), .B(n4412), .S(n4597), .Z(n2638) );
  MUX21L U4421 ( .A(n5549), .B(n4412), .S(n4605), .Z(n2382) );
  MUX21L U4422 ( .A(n5550), .B(n4412), .S(n4599), .Z(n2606) );
  MUX21L U4423 ( .A(n5551), .B(n4412), .S(n4600), .Z(n2510) );
  MUX21L U4424 ( .A(n5552), .B(n4412), .S(n4601), .Z(n2574) );
  MUX21L U4425 ( .A(n5553), .B(n4412), .S(n4602), .Z(n2414) );
  MUX21L U4426 ( .A(n5554), .B(n4412), .S(n4603), .Z(n2542) );
  MUX21L U4427 ( .A(n5555), .B(n4412), .S(n4604), .Z(n2478) );
  MUX21L U4428 ( .A(n4834), .B(n4412), .S(n4598), .Z(n2446) );
  MUX21L U4429 ( .A(n5556), .B(n4412), .S(n4606), .Z(n2990) );
  MUX21L U4430 ( .A(n5557), .B(n4412), .S(n4607), .Z(n3118) );
  MUX21L U4431 ( .A(n5558), .B(n4412), .S(n4608), .Z(n3022) );
  MUX21L U4432 ( .A(n5559), .B(n4412), .S(n4609), .Z(n3086) );
  MUX21L U4433 ( .A(n5560), .B(n4412), .S(n4610), .Z(n2926) );
  MUX21L U4434 ( .A(n5561), .B(n4412), .S(n4611), .Z(n3054) );
  MUX21L U4435 ( .A(n5562), .B(n4412), .S(n4612), .Z(n2894) );
  MUX21L U4436 ( .A(n4801), .B(n4412), .S(n4613), .Z(n2958) );
  MUX21L U4437 ( .A(n5563), .B(n4412), .S(n4614), .Z(n3246) );
  MUX21L U4438 ( .A(n5564), .B(n4412), .S(n4615), .Z(n3310) );
  MUX21L U4439 ( .A(n5565), .B(n4412), .S(n4616), .Z(n3150) );
  MUX21L U4440 ( .A(n5716), .B(n4412), .S(n4617), .Z(n3182) );
  MUX21L U4441 ( .A(n5717), .B(n4412), .S(n4619), .Z(n3342) );
  MUX21L U4442 ( .A(n5718), .B(n4412), .S(n4620), .Z(n3278) );
  AO2 U4443 ( .A(\gpr[18][27] ), .B(n4458), .C(\gpr[16][27] ), .D(n4626), .Z(
        n4420) );
  AO2 U4444 ( .A(\gpr[17][27] ), .B(n4636), .C(\gpr[20][27] ), .D(n4498), .Z(
        n4419) );
  AO2 U4445 ( .A(\gpr[21][27] ), .B(n4639), .C(\gpr[23][27] ), .D(n4413), .Z(
        n4418) );
  AN2I U4446 ( .A(\gpr[22][27] ), .B(n4489), .Z(n4416) );
  ND2I U4447 ( .A(\gpr[19][27] ), .B(n4501), .Z(n4414) );
  ND2I U4448 ( .A(n4628), .B(n4414), .Z(n4415) );
  NR2I U4449 ( .A(n4416), .B(n4415), .Z(n4417) );
  ND4 U4450 ( .A(n4420), .B(n4419), .C(n4418), .D(n4417), .Z(n4426) );
  AO2 U4451 ( .A(\gpr[26][27] ), .B(n4458), .C(\gpr[29][27] ), .D(n4639), .Z(
        n4424) );
  AO2 U4452 ( .A(\gpr[24][27] ), .B(n4450), .C(\gpr[30][27] ), .D(n4431), .Z(
        n4422) );
  ND4 U4453 ( .A(n4424), .B(n4423), .C(n4422), .D(n4421), .Z(n4425) );
  AN2I U4454 ( .A(n4426), .B(n4425), .Z(n4448) );
  AO2 U4455 ( .A(\gpr[2][27] ), .B(n4659), .C(\gpr[7][27] ), .D(n4675), .Z(
        n4445) );
  AO2 U4456 ( .A(\gpr[1][27] ), .B(n4656), .C(\gpr[3][27] ), .D(n4657), .Z(
        n4430) );
  ND2I U4457 ( .A(\gpr[4][27] ), .B(n4666), .Z(n4428) );
  ND2I U4458 ( .A(n4658), .B(\gpr[5][27] ), .Z(n4427) );
  AN2I U4459 ( .A(n4428), .B(n4427), .Z(n4429) );
  AN2I U4460 ( .A(n4430), .B(n4429), .Z(n4444) );
  AO2 U4461 ( .A(\gpr[8][27] ), .B(n4432), .C(\gpr[14][27] ), .D(n4431), .Z(
        n4440) );
  ND2I U4462 ( .A(\gpr[10][27] ), .B(n4458), .Z(n4434) );
  ND2I U4463 ( .A(\gpr[9][27] ), .B(n4636), .Z(n4433) );
  ND2I U4464 ( .A(n4434), .B(n4433), .Z(n4438) );
  ND2I U4465 ( .A(\gpr[11][27] ), .B(n4501), .Z(n4436) );
  ND2I U4466 ( .A(\gpr[12][27] ), .B(n4498), .Z(n4435) );
  ND2I U4467 ( .A(n4436), .B(n4435), .Z(n4437) );
  NR2I U4468 ( .A(n4438), .B(n4437), .Z(n4439) );
  ND2I U4469 ( .A(n4440), .B(n4439), .Z(n4441) );
  ND2I U4470 ( .A(n4442), .B(n4441), .Z(n4443) );
  ND4 U4471 ( .A(n4446), .B(n4445), .C(n4444), .D(n4443), .Z(n4447) );
  AN2I U4472 ( .A(n4448), .B(n4447), .Z(rd_data2[27]) );
  B4IP U4473 ( .A(wr_data[28]), .Z(n4449) );
  MUX21L U4474 ( .A(n5566), .B(n4449), .S(n4605), .Z(n2383) );
  MUX21L U4475 ( .A(n5567), .B(n4449), .S(n4598), .Z(n2447) );
  MUX21L U4476 ( .A(n5568), .B(n4449), .S(n4604), .Z(n2479) );
  MUX21L U4477 ( .A(n5569), .B(n4449), .S(n4599), .Z(n2607) );
  MUX21L U4478 ( .A(n4878), .B(n4449), .S(n4602), .Z(n2415) );
  MUX21L U4479 ( .A(n5570), .B(n4449), .S(n4603), .Z(n2543) );
  MUX21L U4480 ( .A(n5571), .B(n4449), .S(n4601), .Z(n2575) );
  MUX21L U4481 ( .A(n5572), .B(n4449), .S(n4600), .Z(n2511) );
  MUX21L U4482 ( .A(n4879), .B(n4449), .S(n4536), .Z(n2639) );
  MUX21L U4483 ( .A(n5573), .B(n4449), .S(n4590), .Z(n2703) );
  MUX21L U4484 ( .A(n5574), .B(n4449), .S(n4591), .Z(n2735) );
  MUX21L U4485 ( .A(n5575), .B(n4449), .S(n4596), .Z(n2863) );
  MUX21L U4486 ( .A(n5576), .B(n4449), .S(n4538), .Z(n2671) );
  MUX21L U4487 ( .A(n5577), .B(n4449), .S(n4595), .Z(n2799) );
  MUX21L U4488 ( .A(n5578), .B(n4449), .S(n4593), .Z(n2831) );
  MUX21L U4489 ( .A(n5579), .B(n4449), .S(n4592), .Z(n2767) );
  MUX21L U4490 ( .A(n5580), .B(n4449), .S(n4606), .Z(n2991) );
  MUX21L U4491 ( .A(n5581), .B(n4449), .S(n4607), .Z(n3119) );
  MUX21L U4492 ( .A(n5582), .B(n4449), .S(n4608), .Z(n3023) );
  MUX21L U4493 ( .A(n5583), .B(n4449), .S(n4609), .Z(n3087) );
  MUX21L U4494 ( .A(n4824), .B(n4449), .S(n4610), .Z(n2927) );
  MUX21L U4495 ( .A(n5584), .B(n4449), .S(n4611), .Z(n3055) );
  MUX21L U4496 ( .A(n5585), .B(n4449), .S(n4612), .Z(n2895) );
  MUX21L U4497 ( .A(n4802), .B(n4449), .S(n4613), .Z(n2959) );
  MUX21L U4498 ( .A(n5586), .B(n4449), .S(n4614), .Z(n3247) );
  MUX21L U4499 ( .A(n5587), .B(n4449), .S(n4540), .Z(n3311) );
  MUX21L U4500 ( .A(n5588), .B(n4449), .S(n4616), .Z(n3151) );
  MUX21L U4501 ( .A(n5589), .B(n4449), .S(n4617), .Z(n3183) );
  MUX21L U4502 ( .A(n5590), .B(n4449), .S(n4618), .Z(n3215) );
  MUX21L U4503 ( .A(n5591), .B(n4449), .S(n4619), .Z(n3343) );
  MUX21L U4504 ( .A(n5592), .B(n4449), .S(n4620), .Z(n3279) );
  ND2I U4505 ( .A(\gpr[31][28] ), .B(n4457), .Z(n4452) );
  ND2I U4506 ( .A(\gpr[25][28] ), .B(n4636), .Z(n4451) );
  AN3 U4507 ( .A(n4453), .B(n4452), .C(n4451), .Z(n4456) );
  AO2 U4508 ( .A(\gpr[29][28] ), .B(n4639), .C(\gpr[30][28] ), .D(n4431), .Z(
        n4455) );
  AO2 U4509 ( .A(\gpr[16][28] ), .B(n4549), .C(\gpr[20][28] ), .D(n4498), .Z(
        n4461) );
  AO2 U4510 ( .A(\gpr[21][28] ), .B(n4639), .C(\gpr[22][28] ), .D(n4431), .Z(
        n4460) );
  AO2 U4511 ( .A(\gpr[19][28] ), .B(n4635), .C(\gpr[18][28] ), .D(n4458), .Z(
        n4459) );
  AN2I U4512 ( .A(n4463), .B(n4462), .Z(n4485) );
  ND2I U4513 ( .A(n4802), .B(n4650), .Z(n4464) );
  AO3 U4514 ( .A(\gpr[15][28] ), .B(n4639), .C(n4652), .D(n4464), .Z(n4465) );
  AO3 U4515 ( .A(n4824), .B(n4466), .C(n4561), .D(n4465), .Z(n4472) );
  ND2I U4516 ( .A(\gpr[3][28] ), .B(n4557), .Z(n4470) );
  ND2I U4517 ( .A(\gpr[5][28] ), .B(n4658), .Z(n4469) );
  ND2I U4518 ( .A(\gpr[1][28] ), .B(n4556), .Z(n4468) );
  ND2I U4519 ( .A(\gpr[4][28] ), .B(n4666), .Z(n4467) );
  ND4 U4520 ( .A(n4470), .B(n4469), .C(n4468), .D(n4467), .Z(n4471) );
  NR2I U4521 ( .A(n4472), .B(n4471), .Z(n4483) );
  ND2I U4522 ( .A(\gpr[11][28] ), .B(n4571), .Z(n4479) );
  ND2I U4523 ( .A(\gpr[12][28] ), .B(n4573), .Z(n4478) );
  ND2I U4524 ( .A(\gpr[7][28] ), .B(n4675), .Z(n4477) );
  ND2I U4525 ( .A(\gpr[6][28] ), .B(n4475), .Z(n4476) );
  ND4 U4526 ( .A(n4479), .B(n4478), .C(n4477), .D(n4476), .Z(n4480) );
  NR2I U4527 ( .A(n4481), .B(n4480), .Z(n4482) );
  ND2I U4528 ( .A(n4483), .B(n4482), .Z(n4484) );
  AN2I U4529 ( .A(n4485), .B(n4484), .Z(rd_data2[28]) );
  MUX21L U4530 ( .A(n5593), .B(n4486), .S(n4590), .Z(n2704) );
  MUX21L U4531 ( .A(n5719), .B(n4486), .S(n4591), .Z(n2736) );
  MUX21L U4532 ( .A(n5594), .B(n4486), .S(n4596), .Z(n2864) );
  MUX21L U4533 ( .A(n5595), .B(n4486), .S(n4592), .Z(n2768) );
  MUX21L U4534 ( .A(n4880), .B(n4486), .S(n4538), .Z(n2672) );
  MUX21L U4535 ( .A(n5596), .B(n4486), .S(n4595), .Z(n2800) );
  MUX21L U4536 ( .A(n5597), .B(n4486), .S(n4593), .Z(n2832) );
  MUX21L U4537 ( .A(n5598), .B(n4486), .S(n4597), .Z(n2640) );
  MUX21L U4538 ( .A(n5599), .B(n4486), .S(n4598), .Z(n2448) );
  MUX21L U4539 ( .A(n5720), .B(n4486), .S(n4604), .Z(n2480) );
  MUX21L U4540 ( .A(n5600), .B(n4486), .S(n4599), .Z(n2608) );
  MUX21L U4541 ( .A(n5721), .B(n4486), .S(n4601), .Z(n2576) );
  MUX21L U4542 ( .A(n4810), .B(n4486), .S(n4602), .Z(n2416) );
  MUX21L U4543 ( .A(n5601), .B(n4486), .S(n4603), .Z(n2544) );
  MUX21L U4544 ( .A(n5722), .B(n4486), .S(n4600), .Z(n2512) );
  MUX21L U4545 ( .A(n5602), .B(n4486), .S(n4605), .Z(n2384) );
  MUX21L U4546 ( .A(n5603), .B(n4486), .S(n4606), .Z(n2992) );
  MUX21L U4547 ( .A(n5604), .B(n4486), .S(n4607), .Z(n3120) );
  MUX21L U4548 ( .A(n5605), .B(n4486), .S(n4608), .Z(n3024) );
  MUX21L U4549 ( .A(n5606), .B(n4486), .S(n4609), .Z(n3088) );
  MUX21L U4550 ( .A(n4825), .B(n4486), .S(n4610), .Z(n2928) );
  MUX21L U4551 ( .A(n5607), .B(n4486), .S(n4611), .Z(n3056) );
  MUX21L U4552 ( .A(n5608), .B(n4486), .S(n4612), .Z(n2896) );
  MUX21L U4553 ( .A(n4803), .B(n4486), .S(n4613), .Z(n2960) );
  MUX21L U4554 ( .A(n5609), .B(n4486), .S(n4614), .Z(n3248) );
  MUX21L U4555 ( .A(n5610), .B(n4486), .S(n4615), .Z(n3312) );
  MUX21L U4556 ( .A(n5611), .B(n4486), .S(n4616), .Z(n3152) );
  MUX21L U4557 ( .A(n5612), .B(n4486), .S(n4617), .Z(n3184) );
  MUX21L U4558 ( .A(n5613), .B(n4486), .S(n4618), .Z(n3216) );
  MUX21L U4559 ( .A(n5614), .B(n4486), .S(n4619), .Z(n3344) );
  MUX21L U4560 ( .A(n5615), .B(n4486), .S(n4620), .Z(n3280) );
  AO2 U4561 ( .A(\gpr[18][29] ), .B(n4487), .C(\gpr[16][29] ), .D(n4542), .Z(
        n4496) );
  AO2 U4562 ( .A(\gpr[21][29] ), .B(n4639), .C(\gpr[23][29] ), .D(n4488), .Z(
        n4494) );
  ND2I U4563 ( .A(\gpr[22][29] ), .B(n4489), .Z(n4492) );
  ND2I U4564 ( .A(\gpr[17][29] ), .B(n4490), .Z(n4491) );
  AN3 U4565 ( .A(n4628), .B(n4492), .C(n4491), .Z(n4493) );
  ND4 U4566 ( .A(n4496), .B(n4495), .C(n4494), .D(n4493), .Z(n4509) );
  AO2 U4567 ( .A(\gpr[26][29] ), .B(n4622), .C(\gpr[24][29] ), .D(n4497), .Z(
        n4507) );
  AO2 U4568 ( .A(\gpr[28][29] ), .B(n4498), .C(\gpr[25][29] ), .D(n4636), .Z(
        n4506) );
  AO2 U4569 ( .A(\gpr[29][29] ), .B(n4639), .C(\gpr[31][29] ), .D(n4499), .Z(
        n4505) );
  IVI U4570 ( .A(n4500), .Z(n4642) );
  ND2I U4571 ( .A(\gpr[27][29] ), .B(n4501), .Z(n4502) );
  AO3 U4572 ( .A(n4642), .B(n4810), .C(n4641), .D(n4502), .Z(n4503) );
  IVI U4573 ( .A(n4503), .Z(n4504) );
  ND4 U4574 ( .A(n4507), .B(n4506), .C(n4505), .D(n4504), .Z(n4508) );
  AN2I U4575 ( .A(n4509), .B(n4508), .Z(n4534) );
  ND2I U4576 ( .A(n4803), .B(n4650), .Z(n4510) );
  AO3 U4577 ( .A(\gpr[15][29] ), .B(n4639), .C(n4652), .D(n4510), .Z(n4511) );
  AO3 U4578 ( .A(n4825), .B(n4655), .C(n4561), .D(n4511), .Z(n4517) );
  ND2I U4579 ( .A(\gpr[3][29] ), .B(n4557), .Z(n4515) );
  ND2I U4580 ( .A(\gpr[5][29] ), .B(n4658), .Z(n4514) );
  ND2I U4581 ( .A(\gpr[1][29] ), .B(n4556), .Z(n4513) );
  ND2I U4582 ( .A(\gpr[4][29] ), .B(n4666), .Z(n4512) );
  ND4 U4583 ( .A(n4515), .B(n4514), .C(n4513), .D(n4512), .Z(n4516) );
  NR2I U4584 ( .A(n4517), .B(n4516), .Z(n4532) );
  ND2I U4585 ( .A(\gpr[2][29] ), .B(n4659), .Z(n4523) );
  ND2I U4586 ( .A(n4562), .B(\gpr[10][29] ), .Z(n4522) );
  ND2I U4587 ( .A(\gpr[9][29] ), .B(n4518), .Z(n4521) );
  ND2I U4588 ( .A(\gpr[8][29] ), .B(n4519), .Z(n4520) );
  ND4 U4589 ( .A(n4523), .B(n4522), .C(n4521), .D(n4520), .Z(n4530) );
  ND2I U4590 ( .A(\gpr[11][29] ), .B(n4571), .Z(n4528) );
  ND2I U4591 ( .A(\gpr[12][29] ), .B(n4573), .Z(n4527) );
  ND2I U4592 ( .A(\gpr[7][29] ), .B(n4675), .Z(n4526) );
  ND2I U4593 ( .A(\gpr[6][29] ), .B(n4524), .Z(n4525) );
  ND4 U4594 ( .A(n4528), .B(n4527), .C(n4526), .D(n4525), .Z(n4529) );
  NR2I U4595 ( .A(n4530), .B(n4529), .Z(n4531) );
  ND2I U4596 ( .A(n4532), .B(n4531), .Z(n4533) );
  AN2I U4597 ( .A(n4534), .B(n4533), .Z(rd_data2[29]) );
  B4IP U4598 ( .A(wr_data[30]), .Z(n4541) );
  MUX21L U4599 ( .A(n5616), .B(n4541), .S(n4605), .Z(n2385) );
  MUX21L U4600 ( .A(n5617), .B(n4541), .S(n4599), .Z(n2609) );
  MUX21L U4601 ( .A(n5618), .B(n4541), .S(n4535), .Z(n2513) );
  MUX21L U4602 ( .A(n5619), .B(n4541), .S(n4601), .Z(n2577) );
  MUX21L U4603 ( .A(n4881), .B(n4541), .S(n4602), .Z(n2417) );
  MUX21L U4604 ( .A(n5620), .B(n4541), .S(n4603), .Z(n2545) );
  MUX21L U4605 ( .A(n5621), .B(n4541), .S(n4604), .Z(n2481) );
  MUX21L U4606 ( .A(n5622), .B(n4541), .S(n4598), .Z(n2449) );
  MUX21L U4607 ( .A(n5623), .B(n4541), .S(n4536), .Z(n2641) );
  MUX21L U4608 ( .A(n5624), .B(n4541), .S(n4590), .Z(n2705) );
  MUX21L U4609 ( .A(n5625), .B(n4541), .S(n4537), .Z(n2769) );
  MUX21L U4610 ( .A(n5626), .B(n4541), .S(n4593), .Z(n2833) );
  MUX21L U4611 ( .A(n4882), .B(n4541), .S(n4538), .Z(n2673) );
  MUX21L U4612 ( .A(n5627), .B(n4541), .S(n4595), .Z(n2801) );
  MUX21L U4613 ( .A(n5723), .B(n4541), .S(n4596), .Z(n2865) );
  MUX21L U4614 ( .A(n5628), .B(n4541), .S(n4591), .Z(n2737) );
  MUX21L U4615 ( .A(n5629), .B(n4541), .S(n4613), .Z(n2961) );
  MUX21L U4616 ( .A(n5630), .B(n4541), .S(n4612), .Z(n2897) );
  MUX21L U4617 ( .A(n5631), .B(n4541), .S(n4606), .Z(n2993) );
  MUX21L U4618 ( .A(n5632), .B(n4541), .S(n4607), .Z(n3121) );
  MUX21L U4619 ( .A(n5633), .B(n4541), .S(n4539), .Z(n3025) );
  MUX21L U4620 ( .A(n5634), .B(n4541), .S(n4609), .Z(n3089) );
  MUX21L U4621 ( .A(n5635), .B(n4541), .S(n4610), .Z(n2929) );
  MUX21L U4622 ( .A(n5636), .B(n4541), .S(n4611), .Z(n3057) );
  MUX21L U4623 ( .A(n5637), .B(n4541), .S(n4614), .Z(n3249) );
  MUX21L U4624 ( .A(n5638), .B(n4541), .S(n4540), .Z(n3313) );
  MUX21L U4625 ( .A(n5639), .B(n4541), .S(n4616), .Z(n3153) );
  MUX21L U4626 ( .A(n5640), .B(n4541), .S(n4617), .Z(n3185) );
  MUX21L U4627 ( .A(n5641), .B(n4541), .S(n4618), .Z(n3217) );
  MUX21L U4628 ( .A(n5642), .B(n4541), .S(n4619), .Z(n3345) );
  MUX21L U4629 ( .A(n5643), .B(n4541), .S(n4620), .Z(n3281) );
  AO2 U4630 ( .A(\gpr[29][30] ), .B(n4639), .C(\gpr[26][30] ), .D(n4458), .Z(
        n4547) );
  AO2 U4631 ( .A(\gpr[24][30] ), .B(n4542), .C(\gpr[30][30] ), .D(n4431), .Z(
        n4545) );
  ND4 U4632 ( .A(n4547), .B(n4546), .C(n4545), .D(n4544), .Z(n4555) );
  AO2 U4633 ( .A(\gpr[20][30] ), .B(n4624), .C(\gpr[18][30] ), .D(n4622), .Z(
        n4553) );
  AO2 U4634 ( .A(\gpr[21][30] ), .B(n4639), .C(\gpr[22][30] ), .D(n4431), .Z(
        n4551) );
  ND4 U4635 ( .A(n4553), .B(n4552), .C(n4551), .D(n4550), .Z(n4554) );
  AN2I U4636 ( .A(n4555), .B(n4554), .Z(n4589) );
  ND2I U4637 ( .A(\gpr[1][30] ), .B(n4556), .Z(n4560) );
  ND2I U4638 ( .A(\gpr[3][30] ), .B(n4557), .Z(n4559) );
  ND2I U4639 ( .A(\gpr[5][30] ), .B(n4658), .Z(n4558) );
  ND4 U4640 ( .A(n4561), .B(n4560), .C(n4559), .D(n4558), .Z(n4569) );
  ND2I U4641 ( .A(\gpr[2][30] ), .B(n4659), .Z(n4567) );
  ND2I U4642 ( .A(n4562), .B(\gpr[10][30] ), .Z(n4566) );
  ND2I U4643 ( .A(\gpr[4][30] ), .B(n4666), .Z(n4565) );
  ND2I U4644 ( .A(\gpr[9][30] ), .B(n4563), .Z(n4564) );
  ND4 U4645 ( .A(n4567), .B(n4566), .C(n4565), .D(n4564), .Z(n4568) );
  NR2I U4646 ( .A(n4569), .B(n4568), .Z(n4587) );
  ND2I U4647 ( .A(\gpr[8][30] ), .B(n4570), .Z(n4577) );
  ND2I U4648 ( .A(\gpr[11][30] ), .B(n4571), .Z(n4576) );
  ND2I U4649 ( .A(\gpr[15][30] ), .B(n4572), .Z(n4575) );
  ND2I U4650 ( .A(\gpr[12][30] ), .B(n4573), .Z(n4574) );
  ND4 U4651 ( .A(n4577), .B(n4576), .C(n4575), .D(n4574), .Z(n4585) );
  ND2I U4652 ( .A(\gpr[6][30] ), .B(n4674), .Z(n4583) );
  ND2I U4653 ( .A(\gpr[13][30] ), .B(n4578), .Z(n4582) );
  ND2I U4654 ( .A(\gpr[7][30] ), .B(n4675), .Z(n4581) );
  ND2I U4655 ( .A(\gpr[14][30] ), .B(n4579), .Z(n4580) );
  ND4 U4656 ( .A(n4583), .B(n4582), .C(n4581), .D(n4580), .Z(n4584) );
  NR2I U4657 ( .A(n4585), .B(n4584), .Z(n4586) );
  ND2I U4658 ( .A(n4587), .B(n4586), .Z(n4588) );
  AN2I U4659 ( .A(n4589), .B(n4588), .Z(rd_data2[30]) );
  B4IP U4660 ( .A(wr_data[31]), .Z(n4621) );
  MUX21L U4661 ( .A(n5644), .B(n4621), .S(n4590), .Z(n2706) );
  MUX21L U4662 ( .A(n317), .B(n4621), .S(n4591), .Z(n2738) );
  MUX21L U4663 ( .A(n5645), .B(n4621), .S(n4592), .Z(n2770) );
  MUX21L U4664 ( .A(n5646), .B(n4621), .S(n4593), .Z(n2834) );
  MUX21L U4665 ( .A(n4883), .B(n4621), .S(n4594), .Z(n2674) );
  MUX21L U4666 ( .A(n5647), .B(n4621), .S(n4595), .Z(n2802) );
  MUX21L U4667 ( .A(n5648), .B(n4621), .S(n4596), .Z(n2866) );
  MUX21L U4668 ( .A(n5649), .B(n4621), .S(n4597), .Z(n2642) );
  MUX21L U4669 ( .A(n5650), .B(n4621), .S(n4598), .Z(n2450) );
  MUX21L U4670 ( .A(n5651), .B(n4621), .S(n4599), .Z(n2610) );
  MUX21L U4671 ( .A(n5652), .B(n4621), .S(n4600), .Z(n2514) );
  MUX21L U4672 ( .A(n5653), .B(n4621), .S(n4601), .Z(n2578) );
  MUX21L U4673 ( .A(n4811), .B(n4621), .S(n4602), .Z(n2418) );
  MUX21L U4674 ( .A(n5654), .B(n4621), .S(n4603), .Z(n2546) );
  MUX21L U4675 ( .A(n318), .B(n4621), .S(n4604), .Z(n2482) );
  MUX21L U4676 ( .A(n5655), .B(n4621), .S(n4605), .Z(n2386) );
  MUX21L U4677 ( .A(n5656), .B(n4621), .S(n4606), .Z(n2994) );
  MUX21L U4678 ( .A(n5657), .B(n4621), .S(n4607), .Z(n3122) );
  MUX21L U4679 ( .A(n5658), .B(n4621), .S(n4608), .Z(n3026) );
  MUX21L U4680 ( .A(n5659), .B(n4621), .S(n4609), .Z(n3090) );
  MUX21L U4681 ( .A(n4826), .B(n4621), .S(n4610), .Z(n2930) );
  MUX21L U4682 ( .A(n5660), .B(n4621), .S(n4611), .Z(n3058) );
  MUX21L U4683 ( .A(n5661), .B(n4621), .S(n4612), .Z(n2898) );
  MUX21L U4684 ( .A(n4804), .B(n4621), .S(n4613), .Z(n2962) );
  MUX21L U4685 ( .A(n5662), .B(n4621), .S(n4614), .Z(n3250) );
  MUX21L U4686 ( .A(n5663), .B(n4621), .S(n4615), .Z(n3314) );
  MUX21L U4687 ( .A(n5664), .B(n4621), .S(n4616), .Z(n3154) );
  MUX21L U4688 ( .A(n5665), .B(n4621), .S(n4617), .Z(n3186) );
  MUX21L U4689 ( .A(n5666), .B(n4621), .S(n4618), .Z(n3218) );
  MUX21L U4690 ( .A(n5667), .B(n4621), .S(n4619), .Z(n3346) );
  MUX21L U4691 ( .A(n5668), .B(n4621), .S(n4620), .Z(n3282) );
  AO2 U4692 ( .A(\gpr[17][31] ), .B(n4636), .C(\gpr[20][31] ), .D(n4624), .Z(
        n4633) );
  AO2 U4693 ( .A(\gpr[21][31] ), .B(n4639), .C(\gpr[23][31] ), .D(n4638), .Z(
        n4632) );
  AN2I U4694 ( .A(\gpr[22][31] ), .B(n4625), .Z(n4630) );
  ND2I U4695 ( .A(\gpr[16][31] ), .B(n4626), .Z(n4627) );
  ND2I U4696 ( .A(n4628), .B(n4627), .Z(n4629) );
  NR2I U4697 ( .A(n4630), .B(n4629), .Z(n4631) );
  ND4 U4698 ( .A(n4634), .B(n4633), .C(n4632), .D(n4631), .Z(n4649) );
  AO2 U4699 ( .A(\gpr[26][31] ), .B(n4622), .C(\gpr[27][31] ), .D(n4635), .Z(
        n4647) );
  AO2 U4700 ( .A(\gpr[24][31] ), .B(n4637), .C(\gpr[25][31] ), .D(n4636), .Z(
        n4646) );
  AO2 U4701 ( .A(\gpr[29][31] ), .B(n4639), .C(\gpr[31][31] ), .D(n4638), .Z(
        n4645) );
  ND2I U4702 ( .A(\gpr[28][31] ), .B(n219), .Z(n4640) );
  AO3 U4703 ( .A(n4642), .B(n4811), .C(n4641), .D(n4640), .Z(n4643) );
  IVI U4704 ( .A(n4643), .Z(n4644) );
  ND4 U4705 ( .A(n4647), .B(n4646), .C(n4645), .D(n4644), .Z(n4648) );
  AN2I U4706 ( .A(n4649), .B(n4648), .Z(n4685) );
  ND2I U4707 ( .A(n4804), .B(n4650), .Z(n4651) );
  AO3 U4708 ( .A(\gpr[15][31] ), .B(n4653), .C(n4652), .D(n4651), .Z(n4654) );
  AO3 U4709 ( .A(n4826), .B(n4655), .C(n295), .D(n4654), .Z(n4665) );
  ND2I U4710 ( .A(\gpr[1][31] ), .B(n4656), .Z(n4663) );
  ND2I U4711 ( .A(\gpr[3][31] ), .B(n4657), .Z(n4662) );
  ND2I U4712 ( .A(\gpr[5][31] ), .B(n4658), .Z(n4661) );
  ND2I U4713 ( .A(\gpr[2][31] ), .B(n4659), .Z(n4660) );
  ND4 U4714 ( .A(n4663), .B(n4662), .C(n4661), .D(n4660), .Z(n4664) );
  NR2I U4715 ( .A(n4665), .B(n4664), .Z(n4683) );
  ND2I U4716 ( .A(\gpr[4][31] ), .B(n4666), .Z(n4672) );
  ND2I U4717 ( .A(n3679), .B(\gpr[10][31] ), .Z(n4671) );
  ND2I U4718 ( .A(\gpr[11][31] ), .B(n4667), .Z(n4670) );
  ND2I U4719 ( .A(\gpr[9][31] ), .B(n4668), .Z(n4669) );
  ND4 U4720 ( .A(n4672), .B(n4671), .C(n4670), .D(n4669), .Z(n4681) );
  ND2I U4721 ( .A(\gpr[12][31] ), .B(n4673), .Z(n4679) );
  ND2I U4722 ( .A(\gpr[8][31] ), .B(n3960), .Z(n4678) );
  ND2I U4723 ( .A(\gpr[6][31] ), .B(n4674), .Z(n4677) );
  ND2I U4724 ( .A(\gpr[7][31] ), .B(n4675), .Z(n4676) );
  ND4 U4725 ( .A(n4679), .B(n4678), .C(n4677), .D(n4676), .Z(n4680) );
  NR2I U4726 ( .A(n4681), .B(n4680), .Z(n4682) );
  ND2I U4727 ( .A(n4683), .B(n4682), .Z(n4684) );
  AN2I U4728 ( .A(n4685), .B(n4684), .Z(rd_data2[31]) );
  AO2 U4729 ( .A(n4726), .B(\gpr[26][25] ), .C(n2231), .D(\gpr[25][25] ), .Z(
        n4700) );
  NR2I U4730 ( .A(n4687), .B(n4874), .Z(n4692) );
  ND2I U4731 ( .A(n4688), .B(\gpr[27][25] ), .Z(n4689) );
  ND2I U4732 ( .A(n2079), .B(n4689), .Z(n4691) );
  NR2I U4733 ( .A(n4692), .B(n4691), .Z(n4699) );
  ND2I U4734 ( .A(n2268), .B(\gpr[29][25] ), .Z(n4696) );
  ND2I U4735 ( .A(\gpr[28][25] ), .B(n4694), .Z(n4695) );
  ND2I U4736 ( .A(n4696), .B(n4695), .Z(n4697) );
  IVI U4737 ( .A(n4697), .Z(n4698) );
  AO2 U4738 ( .A(n4702), .B(\gpr[18][25] ), .C(n4701), .D(\gpr[21][25] ), .Z(
        n4715) );
  AO2P U4739 ( .A(n878), .B(\gpr[16][25] ), .C(n4703), .D(\gpr[19][25] ), .Z(
        n4714) );
  ND2I U4740 ( .A(\gpr[20][25] ), .B(n2158), .Z(n4706) );
  ND2I U4741 ( .A(\gpr[23][25] ), .B(n4704), .Z(n4705) );
  AN2I U4742 ( .A(n4706), .B(n4705), .Z(n4713) );
  NR2I U4743 ( .A(n4707), .B(n4875), .Z(n4711) );
  ND2I U4744 ( .A(n1466), .B(\gpr[17][25] ), .Z(n4708) );
  ND2I U4745 ( .A(n4709), .B(n4708), .Z(n4710) );
  NR2I U4746 ( .A(n4711), .B(n4710), .Z(n4712) );
  ND4 U4747 ( .A(n4715), .B(n4714), .C(n4713), .D(n4712), .Z(n4716) );
  AN2I U4748 ( .A(n4717), .B(n4716), .Z(n4758) );
  ND2I U4749 ( .A(\gpr[13][25] ), .B(n4718), .Z(n4722) );
  ND2I U4750 ( .A(\gpr[1][25] ), .B(n4719), .Z(n4721) );
  ND2I U4751 ( .A(n2115), .B(\gpr[2][25] ), .Z(n4720) );
  ND4 U4752 ( .A(n498), .B(n4722), .C(n4721), .D(n4720), .Z(n4736) );
  ND2I U4753 ( .A(n4723), .B(\gpr[5][25] ), .Z(n4730) );
  ND2I U4754 ( .A(n4724), .B(\gpr[3][25] ), .Z(n4728) );
  ND2I U4755 ( .A(n4726), .B(n297), .Z(n4727) );
  AN2I U4756 ( .A(n4728), .B(n4727), .Z(n4729) );
  ND2I U4757 ( .A(n4730), .B(n4729), .Z(n4731) );
  IVI U4758 ( .A(n4731), .Z(n4734) );
  ND2I U4759 ( .A(\gpr[4][25] ), .B(n4732), .Z(n4733) );
  ND2I U4760 ( .A(n4734), .B(n4733), .Z(n4735) );
  NR2I U4761 ( .A(n4736), .B(n4735), .Z(n4756) );
  ND2I U4762 ( .A(n4737), .B(\gpr[9][25] ), .Z(n4744) );
  ND2I U4763 ( .A(n4738), .B(\gpr[8][25] ), .Z(n4743) );
  ND2I U4764 ( .A(n4739), .B(\gpr[11][25] ), .Z(n4742) );
  ND2I U4765 ( .A(n106), .B(\gpr[12][25] ), .Z(n4741) );
  ND4 U4766 ( .A(n4744), .B(n4743), .C(n4742), .D(n4741), .Z(n4754) );
  ND2I U4767 ( .A(\gpr[15][25] ), .B(n4745), .Z(n4752) );
  ND2I U4768 ( .A(n4746), .B(\gpr[6][25] ), .Z(n4751) );
  ND2I U4769 ( .A(n4747), .B(\gpr[7][25] ), .Z(n4750) );
  ND2I U4770 ( .A(n4748), .B(\gpr[14][25] ), .Z(n4749) );
  ND4 U4771 ( .A(n4752), .B(n4751), .C(n4750), .D(n4749), .Z(n4753) );
  NR2I U4772 ( .A(n4754), .B(n4753), .Z(n4755) );
  ND2I U4773 ( .A(n4756), .B(n4755), .Z(n4757) );
  AN2I U4774 ( .A(n4758), .B(n4757), .Z(rd_data1[25]) );
endmodule


module processor ( clock, reset, PC, Inst, MemRead, MemWrite, Addr, Din, Dout
 );
  output [31:0] PC;
  input [31:0] Inst;
  output [31:0] Addr;
  output [31:0] Din;
  input [31:0] Dout;
  input clock, reset;
  output MemRead, MemWrite;
  wire   mw_Inst_5, mw_Inst_4, mw_Inst_2, mw_Inst_1, mw_Inst_0, xm_Inst_5,
         xm_Inst_4, xm_Inst_2, xm_Inst_1, xm_Inst_0, w_RegWrite, \pc_u0/N31 ,
         \pc_u0/N30 , \pc_u0/N29 , \pc_u0/N28 , \pc_u0/N27 , \pc_u0/N26 ,
         \pc_u0/N25 , \pc_u0/N24 , \pc_u0/N23 , \pc_u0/N22 , \pc_u0/N21 ,
         \pc_u0/N20 , \pc_u0/N19 , \pc_u0/N18 , \pc_u0/N17 , \pc_u0/N16 ,
         \pc_u0/N15 , \pc_u0/N14 , \pc_u0/N13 , \pc_u0/N12 , \pc_u0/N11 ,
         \pc_u0/N10 , \pc_u0/N9 , \pc_u0/N8 , \pc_u0/N7 , \pc_u0/N6 ,
         \pc_u0/N5 , \pc_u0/N4 , n1137, n1139, n1140, n1141, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874;
  wire   [31:0] fd_Inst;
  wire   [31:0] Inst_stall_b_j;
  wire   [31:0] gpr_rd_data2;
  wire   [31:11] dx_Inst;
  wire   [31:0] dx_pc_plus_8;
  wire   [31:0] x_ALU_Result;
  wire   [31:0] dx_Inst_15_0_signext;
  wire   [31:0] dx_gpr_rd_data1;
  wire   [4:0] dx_gpr_rd_addr1;
  wire   [31:11] mw_Inst;
  wire   [31:0] mw_pc_plus_8;
  wire   [31:0] xm_pc_plus_8;
  wire   [31:11] xm_Inst;
  wire   [31:0] dx_gpr_rd_data2;
  wire   [31:0] gpr_rd_data1;
  wire   [4:0] gpr_rd_addr1;
  wire   [4:0] gpr_wr_addr;
  wire   [31:0] gpr_wr_data;
  wire   [31:0] \pc_u0/pc_plus_4 ;
  assign PC[1] = \pc_u0/pc_plus_4  [1];
  assign PC[0] = \pc_u0/pc_plus_4  [0];

  gpr gpr_u0 ( .clk(clock), .RegWrite(w_RegWrite), .rd_addr1(gpr_rd_addr1), 
        .rd_addr2({fd_Inst[20:19], n4714, fd_Inst[17], n4713}), .wr_addr({
        n4874, gpr_wr_addr[3:2], n4712, n4797}), .wr_data(gpr_wr_data), 
        .rd_data2(gpr_rd_data2), .\rd_data1[31]_BAR (gpr_rd_data1[31]), 
        .\rd_data1[30] (gpr_rd_data1[30]), .\rd_data1[29] (gpr_rd_data1[29]), 
        .\rd_data1[28] (gpr_rd_data1[28]), .\rd_data1[27] (gpr_rd_data1[27]), 
        .\rd_data1[26] (gpr_rd_data1[26]), .\rd_data1[25] (gpr_rd_data1[25]), 
        .\rd_data1[24] (gpr_rd_data1[24]), .\rd_data1[23] (gpr_rd_data1[23]), 
        .\rd_data1[22] (gpr_rd_data1[22]), .\rd_data1[21] (gpr_rd_data1[21]), 
        .\rd_data1[20] (gpr_rd_data1[20]), .\rd_data1[19] (gpr_rd_data1[19]), 
        .\rd_data1[17] (gpr_rd_data1[17]), .\rd_data1[16] (gpr_rd_data1[16]), 
        .\rd_data1[15] (gpr_rd_data1[15]), .\rd_data1[14] (gpr_rd_data1[14]), 
        .\rd_data1[13] (gpr_rd_data1[13]), .\rd_data1[12] (gpr_rd_data1[12]), 
        .\rd_data1[11] (gpr_rd_data1[11]), .\rd_data1[10] (gpr_rd_data1[10]), 
        .\rd_data1[9] (gpr_rd_data1[9]), .\rd_data1[8] (gpr_rd_data1[8]), 
        .\rd_data1[7] (gpr_rd_data1[7]), .\rd_data1[6] (gpr_rd_data1[6]), 
        .\rd_data1[5] (gpr_rd_data1[5]), .\rd_data1[4] (gpr_rd_data1[4]), 
        .\rd_data1[3] (gpr_rd_data1[3]), .\rd_data1[2] (gpr_rd_data1[2]), 
        .\rd_data1[1] (gpr_rd_data1[1]), .\rd_data1[0] (gpr_rd_data1[0]), 
        .\rd_data1[18]_BAR (gpr_rd_data1[18]) );
  FD2 \mw_Dout_reg[31]  ( .D(Dout[31]), .CP(clock), .CD(n4873), .QN(n4801) );
  FD2 \mw_Dout_reg[30]  ( .D(Dout[30]), .CP(clock), .CD(n4873), .QN(n4807) );
  FD2 \mw_Dout_reg[29]  ( .D(Dout[29]), .CP(clock), .CD(n4873), .QN(n4783) );
  FD2 \mw_Dout_reg[28]  ( .D(Dout[28]), .CP(clock), .CD(n4873), .QN(n4787) );
  FD2 \mw_Dout_reg[27]  ( .D(Dout[27]), .CP(clock), .CD(n4873), .QN(n4808) );
  FD2 \mw_Dout_reg[26]  ( .D(Dout[26]), .CP(clock), .CD(n4873), .QN(n4802) );
  FD2 \mw_Dout_reg[25]  ( .D(Dout[25]), .CP(clock), .CD(n4873), .QN(n4800) );
  FD2 \mw_Dout_reg[24]  ( .D(Dout[24]), .CP(clock), .CD(n4873), .QN(n4810) );
  FD2 \mw_Dout_reg[23]  ( .D(Dout[23]), .CP(clock), .CD(n4873), .QN(n4809) );
  FD2 \mw_Dout_reg[22]  ( .D(Dout[22]), .CP(clock), .CD(n4873), .QN(n4799) );
  FD2 \mw_Dout_reg[21]  ( .D(Dout[21]), .CP(clock), .CD(n4873), .QN(n4811) );
  FD2 \mw_Dout_reg[20]  ( .D(Dout[20]), .CP(clock), .CD(n4873), .QN(n4812) );
  FD2 \mw_Dout_reg[19]  ( .D(Dout[19]), .CP(clock), .CD(n4873), .QN(n4798) );
  FD2 \mw_Dout_reg[18]  ( .D(Dout[18]), .CP(clock), .CD(n4873), .QN(n4786) );
  FD2 \mw_Dout_reg[17]  ( .D(Dout[17]), .CP(clock), .CD(n4873), .QN(n4813) );
  FD2 \mw_Dout_reg[16]  ( .D(Dout[16]), .CP(clock), .CD(n4873), .QN(n4785) );
  FD2 \mw_Dout_reg[15]  ( .D(Dout[15]), .CP(clock), .CD(n4873), .QN(n4790) );
  FD2 \mw_Dout_reg[14]  ( .D(Dout[14]), .CP(clock), .CD(n4873), .QN(n4814) );
  FD2 \mw_Dout_reg[13]  ( .D(Dout[13]), .CP(clock), .CD(n4873), .QN(n4815) );
  FD2 \mw_Dout_reg[12]  ( .D(Dout[12]), .CP(clock), .CD(n4873), .QN(n4816) );
  FD2 \mw_Dout_reg[11]  ( .D(Dout[11]), .CP(clock), .CD(n4873), .QN(n4817) );
  FD2 \mw_Dout_reg[10]  ( .D(Dout[10]), .CP(clock), .CD(n4873), .QN(n4804) );
  FD2 \mw_Dout_reg[9]  ( .D(Dout[9]), .CP(clock), .CD(n4873), .QN(n4803) );
  FD2 \mw_Dout_reg[8]  ( .D(Dout[8]), .CP(clock), .CD(n4873), .QN(n4805) );
  FD2 \mw_Dout_reg[7]  ( .D(Dout[7]), .CP(clock), .CD(n4873), .QN(n4789) );
  FD2 \mw_Dout_reg[6]  ( .D(Dout[6]), .CP(clock), .CD(n4873), .QN(n4806) );
  FD2 \mw_Dout_reg[5]  ( .D(Dout[5]), .CP(clock), .CD(n4873), .QN(n4788) );
  FD2 \mw_Dout_reg[4]  ( .D(Dout[4]), .CP(clock), .CD(n4873), .QN(n4791) );
  FD2 \mw_Dout_reg[3]  ( .D(Dout[3]), .CP(clock), .CD(n4873), .QN(n4793) );
  FD2 \mw_Dout_reg[2]  ( .D(Dout[2]), .CP(clock), .CD(n4873), .QN(n4818) );
  FD2 \mw_Dout_reg[1]  ( .D(Dout[1]), .CP(clock), .CD(n4873), .QN(n4792) );
  FD2 \mw_Dout_reg[0]  ( .D(Dout[0]), .CP(clock), .CD(n4873), .QN(n4784) );
  FD2 \dx_pc_plus_8_reg[31]  ( .D(\pc_u0/pc_plus_4 [31]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[31]) );
  FD2 \xm_pc_plus_8_reg[31]  ( .D(dx_pc_plus_8[31]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[31]) );
  FD2 \dx_pc_plus_8_reg[30]  ( .D(\pc_u0/pc_plus_4 [30]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[30]) );
  FD2 \xm_pc_plus_8_reg[30]  ( .D(dx_pc_plus_8[30]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[30]) );
  FD2 \dx_pc_plus_8_reg[29]  ( .D(\pc_u0/pc_plus_4 [29]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[29]) );
  FD2 \xm_pc_plus_8_reg[29]  ( .D(dx_pc_plus_8[29]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[29]) );
  FD2 \dx_pc_plus_8_reg[28]  ( .D(\pc_u0/pc_plus_4 [28]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[28]) );
  FD2 \xm_pc_plus_8_reg[28]  ( .D(dx_pc_plus_8[28]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[28]) );
  FD2 \dx_pc_plus_8_reg[27]  ( .D(\pc_u0/pc_plus_4 [27]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[27]) );
  FD2 \xm_pc_plus_8_reg[27]  ( .D(dx_pc_plus_8[27]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[27]) );
  FD2 \dx_pc_plus_8_reg[26]  ( .D(\pc_u0/pc_plus_4 [26]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[26]) );
  FD2 \xm_pc_plus_8_reg[26]  ( .D(dx_pc_plus_8[26]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[26]) );
  FD2 \dx_pc_plus_8_reg[25]  ( .D(\pc_u0/pc_plus_4 [25]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[25]) );
  FD2 \xm_pc_plus_8_reg[25]  ( .D(dx_pc_plus_8[25]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[25]) );
  FD2 \dx_pc_plus_8_reg[24]  ( .D(\pc_u0/pc_plus_4 [24]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[24]) );
  FD2 \xm_pc_plus_8_reg[24]  ( .D(dx_pc_plus_8[24]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[24]) );
  FD2 \dx_pc_plus_8_reg[23]  ( .D(\pc_u0/pc_plus_4 [23]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[23]) );
  FD2 \xm_pc_plus_8_reg[23]  ( .D(dx_pc_plus_8[23]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[23]) );
  FD2 \dx_pc_plus_8_reg[22]  ( .D(\pc_u0/pc_plus_4 [22]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[22]) );
  FD2 \xm_pc_plus_8_reg[22]  ( .D(dx_pc_plus_8[22]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[22]) );
  FD2 \dx_pc_plus_8_reg[21]  ( .D(\pc_u0/pc_plus_4 [21]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[21]) );
  FD2 \xm_pc_plus_8_reg[21]  ( .D(dx_pc_plus_8[21]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[21]) );
  FD2 \dx_pc_plus_8_reg[20]  ( .D(\pc_u0/pc_plus_4 [20]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[20]) );
  FD2 \xm_pc_plus_8_reg[20]  ( .D(dx_pc_plus_8[20]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[20]) );
  FD2 \dx_pc_plus_8_reg[19]  ( .D(\pc_u0/pc_plus_4 [19]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[19]) );
  FD2 \xm_pc_plus_8_reg[19]  ( .D(dx_pc_plus_8[19]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[19]) );
  FD2 \dx_pc_plus_8_reg[18]  ( .D(\pc_u0/pc_plus_4 [18]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[18]) );
  FD2 \xm_pc_plus_8_reg[18]  ( .D(dx_pc_plus_8[18]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[18]) );
  FD2 \dx_pc_plus_8_reg[17]  ( .D(\pc_u0/pc_plus_4 [17]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[17]) );
  FD2 \xm_pc_plus_8_reg[17]  ( .D(dx_pc_plus_8[17]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[17]) );
  FD2 \dx_pc_plus_8_reg[16]  ( .D(\pc_u0/pc_plus_4 [16]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[16]) );
  FD2 \xm_pc_plus_8_reg[16]  ( .D(dx_pc_plus_8[16]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[16]) );
  FD2 \dx_pc_plus_8_reg[15]  ( .D(\pc_u0/pc_plus_4 [15]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[15]) );
  FD2 \xm_pc_plus_8_reg[15]  ( .D(dx_pc_plus_8[15]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[15]) );
  FD2 \dx_pc_plus_8_reg[14]  ( .D(\pc_u0/pc_plus_4 [14]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[14]) );
  FD2 \xm_pc_plus_8_reg[14]  ( .D(dx_pc_plus_8[14]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[14]) );
  FD2 \dx_pc_plus_8_reg[13]  ( .D(\pc_u0/pc_plus_4 [13]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[13]) );
  FD2 \xm_pc_plus_8_reg[13]  ( .D(dx_pc_plus_8[13]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[13]) );
  FD2 \dx_pc_plus_8_reg[12]  ( .D(\pc_u0/pc_plus_4 [12]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[12]) );
  FD2 \xm_pc_plus_8_reg[12]  ( .D(dx_pc_plus_8[12]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[12]) );
  FD2 \dx_pc_plus_8_reg[11]  ( .D(\pc_u0/pc_plus_4 [11]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[11]) );
  FD2 \xm_pc_plus_8_reg[11]  ( .D(dx_pc_plus_8[11]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[11]) );
  FD2 \dx_pc_plus_8_reg[10]  ( .D(\pc_u0/pc_plus_4 [10]), .CP(clock), .CD(
        n4873), .Q(dx_pc_plus_8[10]) );
  FD2 \xm_pc_plus_8_reg[10]  ( .D(dx_pc_plus_8[10]), .CP(clock), .CD(n4873), 
        .Q(xm_pc_plus_8[10]) );
  FD2 \dx_pc_plus_8_reg[9]  ( .D(\pc_u0/pc_plus_4 [9]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[9]) );
  FD2 \xm_pc_plus_8_reg[9]  ( .D(dx_pc_plus_8[9]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[9]) );
  FD2 \dx_pc_plus_8_reg[8]  ( .D(\pc_u0/pc_plus_4 [8]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[8]) );
  FD2 \xm_pc_plus_8_reg[8]  ( .D(dx_pc_plus_8[8]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[8]) );
  FD2 \dx_pc_plus_8_reg[7]  ( .D(\pc_u0/pc_plus_4 [7]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[7]) );
  FD2 \xm_pc_plus_8_reg[7]  ( .D(dx_pc_plus_8[7]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[7]) );
  FD2 \dx_pc_plus_8_reg[6]  ( .D(\pc_u0/pc_plus_4 [6]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[6]) );
  FD2 \xm_pc_plus_8_reg[6]  ( .D(dx_pc_plus_8[6]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[6]) );
  FD2 \dx_pc_plus_8_reg[5]  ( .D(\pc_u0/pc_plus_4 [5]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[5]) );
  FD2 \xm_pc_plus_8_reg[5]  ( .D(dx_pc_plus_8[5]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[5]) );
  FD2 \dx_pc_plus_8_reg[4]  ( .D(\pc_u0/pc_plus_4 [4]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[4]) );
  FD2 \xm_pc_plus_8_reg[4]  ( .D(dx_pc_plus_8[4]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[4]) );
  FD2 \dx_pc_plus_8_reg[3]  ( .D(\pc_u0/pc_plus_4 [3]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[3]) );
  FD2 \xm_pc_plus_8_reg[3]  ( .D(dx_pc_plus_8[3]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[3]) );
  FD2 \dx_pc_plus_8_reg[2]  ( .D(n1462), .CP(clock), .CD(n4873), .Q(
        dx_pc_plus_8[2]) );
  FD2 \xm_pc_plus_8_reg[2]  ( .D(dx_pc_plus_8[2]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[2]) );
  FD2 \dx_pc_plus_8_reg[1]  ( .D(\pc_u0/pc_plus_4 [1]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[1]) );
  FD2 \xm_pc_plus_8_reg[1]  ( .D(dx_pc_plus_8[1]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[1]) );
  FD2 \dx_pc_plus_8_reg[0]  ( .D(\pc_u0/pc_plus_4 [0]), .CP(clock), .CD(n4873), 
        .Q(dx_pc_plus_8[0]) );
  FD2 \xm_pc_plus_8_reg[0]  ( .D(dx_pc_plus_8[0]), .CP(clock), .CD(n4873), .Q(
        xm_pc_plus_8[0]) );
  FD2 \mw_pc_plus_8_reg[31]  ( .D(xm_pc_plus_8[31]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[31]) );
  FD2 \mw_pc_plus_8_reg[30]  ( .D(xm_pc_plus_8[30]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[30]) );
  FD2 \mw_pc_plus_8_reg[29]  ( .D(xm_pc_plus_8[29]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[29]) );
  FD2 \mw_pc_plus_8_reg[28]  ( .D(xm_pc_plus_8[28]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[28]) );
  FD2 \mw_pc_plus_8_reg[27]  ( .D(xm_pc_plus_8[27]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[27]) );
  FD2 \mw_pc_plus_8_reg[26]  ( .D(xm_pc_plus_8[26]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[26]) );
  FD2 \mw_pc_plus_8_reg[25]  ( .D(xm_pc_plus_8[25]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[25]) );
  FD2 \mw_pc_plus_8_reg[24]  ( .D(xm_pc_plus_8[24]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[24]) );
  FD2 \mw_pc_plus_8_reg[23]  ( .D(xm_pc_plus_8[23]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[23]) );
  FD2 \mw_pc_plus_8_reg[22]  ( .D(xm_pc_plus_8[22]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[22]) );
  FD2 \mw_pc_plus_8_reg[21]  ( .D(xm_pc_plus_8[21]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[21]) );
  FD2 \mw_pc_plus_8_reg[20]  ( .D(xm_pc_plus_8[20]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[20]) );
  FD2 \mw_pc_plus_8_reg[19]  ( .D(xm_pc_plus_8[19]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[19]) );
  FD2 \mw_pc_plus_8_reg[18]  ( .D(xm_pc_plus_8[18]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[18]) );
  FD2 \mw_pc_plus_8_reg[17]  ( .D(xm_pc_plus_8[17]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[17]) );
  FD2 \mw_pc_plus_8_reg[16]  ( .D(xm_pc_plus_8[16]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[16]) );
  FD2 \mw_pc_plus_8_reg[15]  ( .D(xm_pc_plus_8[15]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[15]) );
  FD2 \mw_pc_plus_8_reg[14]  ( .D(xm_pc_plus_8[14]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[14]) );
  FD2 \mw_pc_plus_8_reg[13]  ( .D(xm_pc_plus_8[13]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[13]) );
  FD2 \mw_pc_plus_8_reg[12]  ( .D(xm_pc_plus_8[12]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[12]) );
  FD2 \mw_pc_plus_8_reg[11]  ( .D(xm_pc_plus_8[11]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[11]) );
  FD2 \mw_pc_plus_8_reg[10]  ( .D(xm_pc_plus_8[10]), .CP(clock), .CD(n4873), 
        .Q(mw_pc_plus_8[10]) );
  FD2 \mw_pc_plus_8_reg[9]  ( .D(xm_pc_plus_8[9]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[9]) );
  FD2 \mw_pc_plus_8_reg[8]  ( .D(xm_pc_plus_8[8]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[8]) );
  FD2 \mw_pc_plus_8_reg[7]  ( .D(xm_pc_plus_8[7]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[7]) );
  FD2 \mw_pc_plus_8_reg[6]  ( .D(xm_pc_plus_8[6]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[6]) );
  FD2 \mw_pc_plus_8_reg[5]  ( .D(xm_pc_plus_8[5]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[5]) );
  FD2 \mw_pc_plus_8_reg[4]  ( .D(xm_pc_plus_8[4]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[4]) );
  FD2 \mw_pc_plus_8_reg[3]  ( .D(xm_pc_plus_8[3]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[3]) );
  FD2 \mw_pc_plus_8_reg[2]  ( .D(xm_pc_plus_8[2]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[2]) );
  FD2 \mw_pc_plus_8_reg[1]  ( .D(xm_pc_plus_8[1]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[1]) );
  FD2 \mw_pc_plus_8_reg[0]  ( .D(xm_pc_plus_8[0]), .CP(clock), .CD(n4873), .Q(
        mw_pc_plus_8[0]) );
  FD2 \dx_gpr_rd_data2_reg[0]  ( .D(gpr_rd_data2[0]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[0]), .QN(n1459) );
  FD2 \xm_gpr_rd_data2_reg[0]  ( .D(dx_gpr_rd_data2[0]), .CP(clock), .CD(n4873), .Q(Din[0]) );
  FD2 \dx_gpr_rd_data2_reg[1]  ( .D(gpr_rd_data2[1]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[1]) );
  FD2 \xm_gpr_rd_data2_reg[1]  ( .D(dx_gpr_rd_data2[1]), .CP(clock), .CD(n4873), .Q(Din[1]) );
  FD2 \xm_gpr_rd_data2_reg[2]  ( .D(dx_gpr_rd_data2[2]), .CP(clock), .CD(n4873), .Q(Din[2]) );
  FD2 \dx_gpr_rd_data2_reg[3]  ( .D(gpr_rd_data2[3]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[3]) );
  FD2 \xm_gpr_rd_data2_reg[3]  ( .D(dx_gpr_rd_data2[3]), .CP(clock), .CD(n4873), .Q(Din[3]) );
  FD2 \xm_gpr_rd_data2_reg[4]  ( .D(dx_gpr_rd_data2[4]), .CP(clock), .CD(n4873), .Q(Din[4]) );
  FD2 \dx_gpr_rd_data2_reg[5]  ( .D(gpr_rd_data2[5]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[5]) );
  FD2 \xm_gpr_rd_data2_reg[5]  ( .D(dx_gpr_rd_data2[5]), .CP(clock), .CD(n4873), .Q(Din[5]) );
  FD2 \dx_gpr_rd_data2_reg[6]  ( .D(gpr_rd_data2[6]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[6]) );
  FD2 \xm_gpr_rd_data2_reg[6]  ( .D(dx_gpr_rd_data2[6]), .CP(clock), .CD(n4873), .Q(Din[6]) );
  FD2 \xm_gpr_rd_data2_reg[7]  ( .D(dx_gpr_rd_data2[7]), .CP(clock), .CD(n4873), .Q(Din[7]) );
  FD2 \dx_gpr_rd_data2_reg[8]  ( .D(gpr_rd_data2[8]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[8]) );
  FD2 \xm_gpr_rd_data2_reg[8]  ( .D(dx_gpr_rd_data2[8]), .CP(clock), .CD(n4873), .Q(Din[8]) );
  FD2 \dx_gpr_rd_data2_reg[9]  ( .D(gpr_rd_data2[9]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[9]) );
  FD2 \xm_gpr_rd_data2_reg[9]  ( .D(dx_gpr_rd_data2[9]), .CP(clock), .CD(n4873), .Q(Din[9]) );
  FD2 \dx_gpr_rd_data2_reg[10]  ( .D(gpr_rd_data2[10]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[10]) );
  FD2 \xm_gpr_rd_data2_reg[10]  ( .D(dx_gpr_rd_data2[10]), .CP(clock), .CD(
        n4873), .Q(Din[10]) );
  FD2 \dx_gpr_rd_data2_reg[11]  ( .D(gpr_rd_data2[11]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[11]) );
  FD2 \xm_gpr_rd_data2_reg[11]  ( .D(dx_gpr_rd_data2[11]), .CP(clock), .CD(
        n4873), .Q(Din[11]) );
  FD2 \dx_gpr_rd_data2_reg[12]  ( .D(gpr_rd_data2[12]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[12]) );
  FD2 \xm_gpr_rd_data2_reg[12]  ( .D(dx_gpr_rd_data2[12]), .CP(clock), .CD(
        n4873), .Q(Din[12]) );
  FD2 \dx_gpr_rd_data2_reg[13]  ( .D(gpr_rd_data2[13]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[13]) );
  FD2 \xm_gpr_rd_data2_reg[13]  ( .D(dx_gpr_rd_data2[13]), .CP(clock), .CD(
        n4873), .Q(Din[13]) );
  FD2 \dx_gpr_rd_data2_reg[14]  ( .D(gpr_rd_data2[14]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[14]) );
  FD2 \xm_gpr_rd_data2_reg[14]  ( .D(dx_gpr_rd_data2[14]), .CP(clock), .CD(
        n4873), .Q(Din[14]) );
  FD2 \xm_gpr_rd_data2_reg[15]  ( .D(dx_gpr_rd_data2[15]), .CP(clock), .CD(
        n4873), .Q(Din[15]) );
  FD2 \dx_gpr_rd_data2_reg[16]  ( .D(gpr_rd_data2[16]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[16]) );
  FD2 \xm_gpr_rd_data2_reg[16]  ( .D(dx_gpr_rd_data2[16]), .CP(clock), .CD(
        n4873), .Q(Din[16]) );
  FD2 \dx_gpr_rd_data2_reg[17]  ( .D(gpr_rd_data2[17]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[17]) );
  FD2 \xm_gpr_rd_data2_reg[17]  ( .D(dx_gpr_rd_data2[17]), .CP(clock), .CD(
        n4873), .Q(Din[17]) );
  FD2 \dx_gpr_rd_data2_reg[18]  ( .D(gpr_rd_data2[18]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[18]) );
  FD2 \xm_gpr_rd_data2_reg[18]  ( .D(dx_gpr_rd_data2[18]), .CP(clock), .CD(
        n4873), .Q(Din[18]) );
  FD2 \dx_gpr_rd_data2_reg[19]  ( .D(gpr_rd_data2[19]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[19]) );
  FD2 \xm_gpr_rd_data2_reg[19]  ( .D(dx_gpr_rd_data2[19]), .CP(clock), .CD(
        n4873), .Q(Din[19]) );
  FD2 \dx_gpr_rd_data2_reg[20]  ( .D(gpr_rd_data2[20]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[20]) );
  FD2 \xm_gpr_rd_data2_reg[20]  ( .D(dx_gpr_rd_data2[20]), .CP(clock), .CD(
        n4873), .Q(Din[20]) );
  FD2 \dx_gpr_rd_data2_reg[21]  ( .D(gpr_rd_data2[21]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[21]) );
  FD2 \xm_gpr_rd_data2_reg[21]  ( .D(dx_gpr_rd_data2[21]), .CP(clock), .CD(
        n4873), .Q(Din[21]) );
  FD2 \dx_gpr_rd_data2_reg[22]  ( .D(gpr_rd_data2[22]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[22]) );
  FD2 \xm_gpr_rd_data2_reg[22]  ( .D(dx_gpr_rd_data2[22]), .CP(clock), .CD(
        n4873), .Q(Din[22]) );
  FD2 \dx_gpr_rd_data2_reg[23]  ( .D(gpr_rd_data2[23]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[23]) );
  FD2 \xm_gpr_rd_data2_reg[23]  ( .D(dx_gpr_rd_data2[23]), .CP(clock), .CD(
        n4873), .Q(Din[23]) );
  FD2 \dx_gpr_rd_data2_reg[24]  ( .D(gpr_rd_data2[24]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[24]) );
  FD2 \xm_gpr_rd_data2_reg[24]  ( .D(dx_gpr_rd_data2[24]), .CP(clock), .CD(
        n4873), .Q(Din[24]) );
  FD2 \dx_gpr_rd_data2_reg[25]  ( .D(gpr_rd_data2[25]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[25]) );
  FD2 \xm_gpr_rd_data2_reg[25]  ( .D(dx_gpr_rd_data2[25]), .CP(clock), .CD(
        n4873), .Q(Din[25]) );
  FD2 \dx_gpr_rd_data2_reg[26]  ( .D(gpr_rd_data2[26]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[26]) );
  FD2 \xm_gpr_rd_data2_reg[26]  ( .D(dx_gpr_rd_data2[26]), .CP(clock), .CD(
        n4873), .Q(Din[26]) );
  FD2 \dx_gpr_rd_data2_reg[27]  ( .D(gpr_rd_data2[27]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[27]) );
  FD2 \xm_gpr_rd_data2_reg[27]  ( .D(dx_gpr_rd_data2[27]), .CP(clock), .CD(
        n4873), .Q(Din[27]) );
  FD2 \dx_gpr_rd_data2_reg[28]  ( .D(gpr_rd_data2[28]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[28]) );
  FD2 \xm_gpr_rd_data2_reg[28]  ( .D(dx_gpr_rd_data2[28]), .CP(clock), .CD(
        n4873), .Q(Din[28]) );
  FD2 \dx_gpr_rd_data2_reg[29]  ( .D(gpr_rd_data2[29]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[29]) );
  FD2 \xm_gpr_rd_data2_reg[29]  ( .D(dx_gpr_rd_data2[29]), .CP(clock), .CD(
        n4873), .Q(Din[29]) );
  FD2 \dx_gpr_rd_data2_reg[30]  ( .D(gpr_rd_data2[30]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[30]) );
  FD2 \xm_gpr_rd_data2_reg[30]  ( .D(dx_gpr_rd_data2[30]), .CP(clock), .CD(
        n4873), .Q(Din[30]) );
  FD2 \dx_gpr_rd_data2_reg[31]  ( .D(gpr_rd_data2[31]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[31]) );
  FD2 \xm_gpr_rd_data2_reg[31]  ( .D(dx_gpr_rd_data2[31]), .CP(clock), .CD(
        n4873), .Q(Din[31]) );
  FD2 \fd_Inst_reg[0]  ( .D(Inst_stall_b_j[0]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[0]), .QN(n4870) );
  FD2 \dx_Inst_15_0_signext_reg[0]  ( .D(fd_Inst[0]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[0]) );
  FD2 \xm_Inst_reg[0]  ( .D(dx_Inst_15_0_signext[0]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst_0) );
  FD2 \mw_Inst_reg[0]  ( .D(xm_Inst_0), .CP(clock), .CD(n4873), .Q(mw_Inst_0)
         );
  FD2 \fd_Inst_reg[1]  ( .D(Inst_stall_b_j[1]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[1]), .QN(n4828) );
  FD2 \dx_Inst_15_0_signext_reg[1]  ( .D(fd_Inst[1]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[1]), .QN(n4773) );
  FD2 \xm_Inst_reg[1]  ( .D(dx_Inst_15_0_signext[1]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst_1) );
  FD2 \mw_Inst_reg[1]  ( .D(xm_Inst_1), .CP(clock), .CD(n4873), .Q(mw_Inst_1)
         );
  FD2 \fd_Inst_reg[2]  ( .D(Inst_stall_b_j[2]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[2]), .QN(n4868) );
  FD2 \dx_Inst_15_0_signext_reg[2]  ( .D(fd_Inst[2]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[2]), .QN(n4770) );
  FD2 \xm_Inst_reg[2]  ( .D(dx_Inst_15_0_signext[2]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst_2) );
  FD2 \mw_Inst_reg[2]  ( .D(xm_Inst_2), .CP(clock), .CD(n4873), .Q(mw_Inst_2)
         );
  FD2 \fd_Inst_reg[3]  ( .D(Inst_stall_b_j[3]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[3]), .QN(n4871) );
  FD2 \dx_Inst_15_0_signext_reg[3]  ( .D(fd_Inst[3]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[3]) );
  FD2 \xm_Inst_reg[3]  ( .D(dx_Inst_15_0_signext[3]), .CP(clock), .CD(n4873), 
        .QN(n1463) );
  FD2 \fd_Inst_reg[4]  ( .D(Inst_stall_b_j[4]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[4]), .QN(n4872) );
  FD2 \dx_Inst_15_0_signext_reg[4]  ( .D(fd_Inst[4]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[4]), .QN(n4769) );
  FD2 \xm_Inst_reg[4]  ( .D(dx_Inst_15_0_signext[4]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst_4) );
  FD2 \mw_Inst_reg[4]  ( .D(xm_Inst_4), .CP(clock), .CD(n4873), .Q(mw_Inst_4)
         );
  FD2 \fd_Inst_reg[5]  ( .D(Inst_stall_b_j[5]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[5]), .QN(n4867) );
  FD2 \dx_Inst_15_0_signext_reg[5]  ( .D(fd_Inst[5]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[5]), .QN(n4771) );
  FD2 \xm_Inst_reg[5]  ( .D(dx_Inst_15_0_signext[5]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst_5) );
  FD2 \mw_Inst_reg[5]  ( .D(xm_Inst_5), .CP(clock), .CD(n4873), .Q(mw_Inst_5)
         );
  FD2 \dx_Inst_15_0_signext_reg[6]  ( .D(fd_Inst[6]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[6]), .QN(n4796) );
  FD2 \dx_Inst_15_0_signext_reg[7]  ( .D(fd_Inst[7]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[7]), .QN(n4795) );
  FD2 \dx_Inst_15_0_signext_reg[8]  ( .D(fd_Inst[8]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[8]) );
  FD2 \dx_Inst_15_0_signext_reg[9]  ( .D(fd_Inst[9]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[9]), .QN(n4822) );
  FD2 \dx_Inst_15_0_signext_reg[10]  ( .D(fd_Inst[10]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[10]), .QN(n4820) );
  FD2 \dx_Inst_15_0_signext_reg[11]  ( .D(fd_Inst[11]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[11]) );
  FD2 \xm_Inst_reg[11]  ( .D(dx_Inst_15_0_signext[11]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst[11]), .QN(n4781) );
  FD2 \dx_Inst_15_0_signext_reg[12]  ( .D(fd_Inst[12]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[12]) );
  FD2 \xm_Inst_reg[12]  ( .D(dx_Inst_15_0_signext[12]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst[12]), .QN(n4766) );
  FD2 \mw_Inst_reg[12]  ( .D(xm_Inst[12]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[12]) );
  FD2 \dx_Inst_15_0_signext_reg[13]  ( .D(fd_Inst[13]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[13]) );
  FD2 \xm_Inst_reg[13]  ( .D(dx_Inst_15_0_signext[13]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst[13]), .QN(n4778) );
  FD2 \mw_Inst_reg[13]  ( .D(xm_Inst[13]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[13]), .QN(n1458) );
  FD2 \dx_Inst_15_0_signext_reg[14]  ( .D(fd_Inst[14]), .CP(clock), .CD(n4873), 
        .Q(dx_Inst_15_0_signext[14]) );
  FD2 \xm_Inst_reg[14]  ( .D(dx_Inst_15_0_signext[14]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst[14]), .QN(n4779) );
  FD2 \mw_Inst_reg[14]  ( .D(xm_Inst[14]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[14]) );
  FD2 \fd_Inst_reg[15]  ( .D(Inst_stall_b_j[15]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[15]), .QN(n4715) );
  FD2 \xm_Inst_reg[15]  ( .D(dx_Inst_15_0_signext[31]), .CP(clock), .CD(n4873), 
        .Q(xm_Inst[15]), .QN(n4780) );
  FD2 \mw_Inst_reg[15]  ( .D(xm_Inst[15]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[15]) );
  FD2 \fd_Inst_reg[16]  ( .D(Inst_stall_b_j[16]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[16]), .QN(n1446) );
  FD2 \dx_Inst_reg[16]  ( .D(n4713), .CP(clock), .CD(n4873), .Q(dx_Inst[16]), 
        .QN(n4762) );
  FD2 \xm_Inst_reg[16]  ( .D(dx_Inst[16]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[16]), .QN(n4768) );
  FD2 \mw_Inst_reg[16]  ( .D(xm_Inst[16]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[16]) );
  FD2 \fd_Inst_reg[17]  ( .D(Inst_stall_b_j[17]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[17]), .QN(n4861) );
  FD2 \dx_Inst_reg[17]  ( .D(n4862), .CP(clock), .CD(n4873), .Q(dx_Inst[17]), 
        .QN(n4716) );
  FD2 \xm_Inst_reg[17]  ( .D(dx_Inst[17]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[17]), .QN(n4763) );
  FD2 \mw_Inst_reg[17]  ( .D(xm_Inst[17]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[17]) );
  FD2 \fd_Inst_reg[18]  ( .D(Inst_stall_b_j[18]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[18]), .QN(n1448) );
  FD2 \dx_Inst_reg[18]  ( .D(n4714), .CP(clock), .CD(n4873), .Q(dx_Inst[18]), 
        .QN(n4777) );
  FD2 \xm_Inst_reg[18]  ( .D(dx_Inst[18]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[18]), .QN(n4764) );
  FD2 \mw_Inst_reg[18]  ( .D(xm_Inst[18]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[18]), .QN(n1457) );
  FD2 \fd_Inst_reg[19]  ( .D(Inst_stall_b_j[19]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[19]), .QN(n4858) );
  FD2 \dx_Inst_reg[19]  ( .D(n4859), .CP(clock), .CD(n4873), .Q(dx_Inst[19]), 
        .QN(n4782) );
  FD2 \xm_Inst_reg[19]  ( .D(dx_Inst[19]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[19]), .QN(n4767) );
  FD2 \mw_Inst_reg[19]  ( .D(xm_Inst[19]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[19]) );
  FD2 \fd_Inst_reg[20]  ( .D(Inst_stall_b_j[20]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[20]), .QN(n4772) );
  FD2 \dx_Inst_reg[20]  ( .D(fd_Inst[20]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[20]), .QN(n4756) );
  FD2 \xm_Inst_reg[20]  ( .D(dx_Inst[20]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[20]), .QN(n4765) );
  FD2 \mw_Inst_reg[20]  ( .D(xm_Inst[20]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[20]) );
  FD2 \fd_Inst_reg[21]  ( .D(Inst_stall_b_j[21]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[21]), .QN(n4759) );
  FD2 \dx_Inst_reg[21]  ( .D(fd_Inst[21]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[21]) );
  FD2 \xm_Inst_reg[21]  ( .D(dx_Inst[21]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[21]) );
  FD2 \mw_Inst_reg[21]  ( .D(xm_Inst[21]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[21]) );
  FD2 \fd_Inst_reg[22]  ( .D(Inst_stall_b_j[22]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[22]), .QN(n4752) );
  FD2 \dx_Inst_reg[22]  ( .D(fd_Inst[22]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[22]) );
  FD2 \xm_Inst_reg[22]  ( .D(dx_Inst[22]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[22]) );
  FD2 \mw_Inst_reg[22]  ( .D(xm_Inst[22]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[22]) );
  FD2 \fd_Inst_reg[23]  ( .D(Inst_stall_b_j[23]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[23]), .QN(n4757) );
  FD2 \dx_Inst_reg[23]  ( .D(fd_Inst[23]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[23]) );
  FD2 \xm_Inst_reg[23]  ( .D(dx_Inst[23]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[23]) );
  FD2 \mw_Inst_reg[23]  ( .D(xm_Inst[23]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[23]) );
  FD2 \fd_Inst_reg[24]  ( .D(Inst_stall_b_j[24]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[24]), .QN(n4758) );
  FD2 \dx_Inst_reg[24]  ( .D(fd_Inst[24]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[24]) );
  FD2 \xm_Inst_reg[24]  ( .D(dx_Inst[24]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[24]) );
  FD2 \mw_Inst_reg[24]  ( .D(xm_Inst[24]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[24]) );
  FD2 \fd_Inst_reg[25]  ( .D(Inst_stall_b_j[25]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[25]), .QN(n4717) );
  FD2 \dx_Inst_reg[25]  ( .D(fd_Inst[25]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[25]) );
  FD2 \xm_Inst_reg[25]  ( .D(dx_Inst[25]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[25]) );
  FD2 \mw_Inst_reg[25]  ( .D(xm_Inst[25]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[25]) );
  FD2 \fd_Inst_reg[26]  ( .D(Inst_stall_b_j[26]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[26]), .QN(n4865) );
  FD2 \dx_Inst_reg[26]  ( .D(fd_Inst[26]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[26]), .QN(n4761) );
  FD2 \xm_Inst_reg[26]  ( .D(dx_Inst[26]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[26]), .QN(n4708) );
  FD2 \mw_Inst_reg[26]  ( .D(n4709), .CP(clock), .CD(n4873), .Q(mw_Inst[26]), 
        .QN(n4824) );
  FD2 \fd_Inst_reg[27]  ( .D(Inst_stall_b_j[27]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[27]), .QN(n4866) );
  FD2 \dx_Inst_reg[27]  ( .D(fd_Inst[27]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[27]) );
  FD2 \xm_Inst_reg[27]  ( .D(dx_Inst[27]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[27]), .QN(n4710) );
  FD2 \mw_Inst_reg[27]  ( .D(n4711), .CP(clock), .CD(n4873), .Q(mw_Inst[27]), 
        .QN(n4825) );
  FD2 \fd_Inst_reg[28]  ( .D(Inst_stall_b_j[28]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[28]), .QN(n4869) );
  FD2 \dx_Inst_reg[28]  ( .D(fd_Inst[28]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[28]), .QN(n4760) );
  FD2 \xm_Inst_reg[28]  ( .D(dx_Inst[28]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[28]), .QN(n4860) );
  FD2 \mw_Inst_reg[28]  ( .D(xm_Inst[28]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[28]), .QN(n4701) );
  FD2 \fd_Inst_reg[29]  ( .D(Inst_stall_b_j[29]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[29]), .QN(n4753) );
  FD2 \dx_Inst_reg[29]  ( .D(fd_Inst[29]), .CP(clock), .CD(n4873), .Q(
        dx_Inst[29]), .QN(n4754) );
  FD2 \xm_Inst_reg[29]  ( .D(dx_Inst[29]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[29]), .QN(n4855) );
  FD2 \mw_Inst_reg[29]  ( .D(n1994), .CP(clock), .CD(n4873), .Q(mw_Inst[29]), 
        .QN(n4864) );
  FD2 \fd_Inst_reg[30]  ( .D(Inst_stall_b_j[30]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[30]), .QN(n4704) );
  FD2 \dx_Inst_reg[30]  ( .D(n4705), .CP(clock), .CD(n4873), .Q(dx_Inst[30])
         );
  FD2 \xm_Inst_reg[30]  ( .D(dx_Inst[30]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[30]), .QN(n4854) );
  FD2 \mw_Inst_reg[30]  ( .D(n4702), .CP(clock), .CD(n4873), .Q(mw_Inst[30]), 
        .QN(n4826) );
  FD2 \fd_Inst_reg[31]  ( .D(Inst_stall_b_j[31]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[31]), .QN(n4706) );
  FD2 \dx_Inst_reg[31]  ( .D(n4707), .CP(clock), .CD(n4873), .Q(dx_Inst[31])
         );
  FD2 \xm_Inst_reg[31]  ( .D(dx_Inst[31]), .CP(clock), .CD(n4873), .Q(
        xm_Inst[31]), .QN(n4755) );
  FD2 \mw_Inst_reg[31]  ( .D(xm_Inst[31]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[31]), .QN(n4863) );
  FD2 \dx_gpr_rd_addr1_reg[0]  ( .D(gpr_rd_addr1[0]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_addr1[0]), .QN(n4774) );
  FD2 \dx_gpr_rd_addr1_reg[1]  ( .D(gpr_rd_addr1[1]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_addr1[1]), .QN(n4776) );
  FD2 \dx_gpr_rd_addr1_reg[3]  ( .D(gpr_rd_addr1[3]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_addr1[3]) );
  FD2 \dx_gpr_rd_addr1_reg[4]  ( .D(gpr_rd_addr1[4]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_addr1[4]), .QN(n4775) );
  FD2 \mw_ALU_Result_reg[31]  ( .D(Addr[31]), .CP(clock), .CD(n4873), .QN(
        n4733) );
  FD2 \mw_ALU_Result_reg[0]  ( .D(Addr[0]), .CP(clock), .CD(n4873), .QN(n4719)
         );
  FD2 \mw_ALU_Result_reg[16]  ( .D(Addr[16]), .CP(clock), .CD(n4873), .QN(
        n4720) );
  FD2 \mw_ALU_Result_reg[24]  ( .D(Addr[24]), .CP(clock), .CD(n4873), .QN(
        n4741) );
  FD2 \xm_ALU_Result_reg[28]  ( .D(x_ALU_Result[28]), .CP(clock), .CD(n4873), 
        .Q(Addr[28]) );
  FD2 \mw_ALU_Result_reg[28]  ( .D(Addr[28]), .CP(clock), .CD(n4873), .QN(
        n4722) );
  FD2 \mw_ALU_Result_reg[30]  ( .D(Addr[30]), .CP(clock), .CD(n4873), .QN(
        n4738) );
  FD2 \mw_ALU_Result_reg[8]  ( .D(Addr[8]), .CP(clock), .CD(n4873), .QN(n4737)
         );
  FD2 \mw_ALU_Result_reg[10]  ( .D(Addr[10]), .CP(clock), .CD(n4873), .QN(
        n4736) );
  FD2 \mw_ALU_Result_reg[12]  ( .D(Addr[12]), .CP(clock), .CD(n4873), .QN(
        n4747) );
  FD2 \mw_ALU_Result_reg[14]  ( .D(Addr[14]), .CP(clock), .CD(n4873), .QN(
        n4745) );
  FD2 \mw_ALU_Result_reg[15]  ( .D(Addr[15]), .CP(clock), .CD(n4873), .QN(
        n4726) );
  FD2 \mw_ALU_Result_reg[4]  ( .D(Addr[4]), .CP(clock), .CD(n4873), .QN(n4727)
         );
  FD2 \mw_ALU_Result_reg[22]  ( .D(Addr[22]), .CP(clock), .CD(n4873), .QN(
        n4731) );
  FD2 \mw_ALU_Result_reg[26]  ( .D(Addr[26]), .CP(clock), .CD(n4873), .QN(
        n4734) );
  FD2 \mw_ALU_Result_reg[27]  ( .D(Addr[27]), .CP(clock), .CD(n4873), .QN(
        n4739) );
  FD2 \mw_ALU_Result_reg[20]  ( .D(Addr[20]), .CP(clock), .CD(n4873), .QN(
        n4743) );
  FD2 \mw_ALU_Result_reg[21]  ( .D(Addr[21]), .CP(clock), .CD(n4873), .QN(
        n4742) );
  FD2 \mw_ALU_Result_reg[18]  ( .D(Addr[18]), .CP(clock), .CD(n4873), .QN(
        n4721) );
  FD2 \mw_ALU_Result_reg[19]  ( .D(Addr[19]), .CP(clock), .CD(n4873), .QN(
        n4730) );
  FD2 \mw_ALU_Result_reg[11]  ( .D(Addr[11]), .CP(clock), .CD(n4873), .QN(
        n4748) );
  FD2 \mw_ALU_Result_reg[13]  ( .D(Addr[13]), .CP(clock), .CD(n4873), .QN(
        n4746) );
  FD2 \mw_ALU_Result_reg[2]  ( .D(Addr[2]), .CP(clock), .CD(n4873), .QN(n4749)
         );
  FD2 \mw_ALU_Result_reg[3]  ( .D(Addr[3]), .CP(clock), .CD(n4873), .QN(n4729)
         );
  FD2 \xm_ALU_Result_reg[1]  ( .D(x_ALU_Result[1]), .CP(clock), .CD(n4873), 
        .Q(Addr[1]) );
  FD2 \mw_ALU_Result_reg[1]  ( .D(Addr[1]), .CP(clock), .CD(n4873), .QN(n4728)
         );
  FD2 \mw_ALU_Result_reg[5]  ( .D(Addr[5]), .CP(clock), .CD(n4873), .QN(n4724)
         );
  FD2 \mw_ALU_Result_reg[25]  ( .D(Addr[25]), .CP(clock), .CD(n4873), .QN(
        n4732) );
  FD2 \mw_ALU_Result_reg[6]  ( .D(Addr[6]), .CP(clock), .CD(n4873), .QN(n4723)
         );
  FD2 \mw_ALU_Result_reg[17]  ( .D(Addr[17]), .CP(clock), .CD(n4873), .QN(
        n4744) );
  FD2 \mw_ALU_Result_reg[7]  ( .D(Addr[7]), .CP(clock), .CD(n4873), .QN(n4725)
         );
  FD2 \mw_ALU_Result_reg[29]  ( .D(Addr[29]), .CP(clock), .CD(n4873), .QN(
        n4718) );
  FD2 \mw_ALU_Result_reg[9]  ( .D(Addr[9]), .CP(clock), .CD(n4873), .QN(n4735)
         );
  FD2 \pc_u0/pc_val_reg[4]  ( .D(\pc_u0/N8 ), .CP(clock), .CD(n4873), .Q(PC[4]), .QN(n4853) );
  FD2 \pc_u0/pc_val_reg[5]  ( .D(\pc_u0/N9 ), .CP(clock), .CD(n4873), .Q(PC[5]), .QN(n4844) );
  FD2 \pc_u0/pc_val_reg[6]  ( .D(\pc_u0/N10 ), .CP(clock), .CD(n4873), .Q(
        PC[6]), .QN(n4852) );
  FD2 \pc_u0/pc_val_reg[7]  ( .D(\pc_u0/N11 ), .CP(clock), .CD(n4873), .Q(
        PC[7]), .QN(n4851) );
  FD2 \pc_u0/pc_val_reg[8]  ( .D(\pc_u0/N12 ), .CP(clock), .CD(n4873), .Q(
        PC[8]), .QN(n4850) );
  FD2 \pc_u0/pc_val_reg[9]  ( .D(\pc_u0/N13 ), .CP(clock), .CD(n4873), .Q(
        PC[9]), .QN(n4845) );
  FD2 \pc_u0/pc_val_reg[10]  ( .D(\pc_u0/N14 ), .CP(clock), .CD(n4873), .Q(
        PC[10]), .QN(n4849) );
  FD2 \pc_u0/pc_val_reg[11]  ( .D(\pc_u0/N15 ), .CP(clock), .CD(n4873), .Q(
        PC[11]), .QN(n4751) );
  FD2 \pc_u0/pc_val_reg[12]  ( .D(\pc_u0/N16 ), .CP(clock), .CD(n4873), .Q(
        PC[12]), .QN(n4848) );
  FD2 \pc_u0/pc_val_reg[13]  ( .D(\pc_u0/N17 ), .CP(clock), .CD(n4873), .Q(
        PC[13]), .QN(n4840) );
  FD2 \pc_u0/pc_val_reg[14]  ( .D(\pc_u0/N18 ), .CP(clock), .CD(n4873), .Q(
        PC[14]), .QN(n4847) );
  FD2 \pc_u0/pc_val_reg[15]  ( .D(\pc_u0/N19 ), .CP(clock), .CD(n4873), .Q(
        PC[15]), .QN(n4839) );
  FD2 \pc_u0/pc_val_reg[16]  ( .D(\pc_u0/N20 ), .CP(clock), .CD(n4873), .Q(
        PC[16]), .QN(n4838) );
  FD2 \pc_u0/pc_val_reg[17]  ( .D(\pc_u0/N21 ), .CP(clock), .CD(n4873), .Q(
        PC[17]), .QN(n4832) );
  FD2 \pc_u0/pc_val_reg[18]  ( .D(\pc_u0/N22 ), .CP(clock), .CD(n4873), .Q(
        PC[18]), .QN(n4846) );
  FD2 \pc_u0/pc_val_reg[19]  ( .D(\pc_u0/N23 ), .CP(clock), .CD(n4873), .Q(
        PC[19]), .QN(n4750) );
  FD2 \pc_u0/pc_val_reg[20]  ( .D(\pc_u0/N24 ), .CP(clock), .CD(n4873), .Q(
        PC[20]), .QN(n4843) );
  FD2 \pc_u0/pc_val_reg[21]  ( .D(\pc_u0/N25 ), .CP(clock), .CD(n4873), .Q(
        PC[21]), .QN(n4837) );
  FD2 \pc_u0/pc_val_reg[22]  ( .D(\pc_u0/N26 ), .CP(clock), .CD(n4873), .Q(
        PC[22]), .QN(n4842) );
  FD2 \pc_u0/pc_val_reg[23]  ( .D(\pc_u0/N27 ), .CP(clock), .CD(n4873), .Q(
        PC[23]), .QN(n4836) );
  FD2 \pc_u0/pc_val_reg[24]  ( .D(\pc_u0/N28 ), .CP(clock), .CD(n4873), .Q(
        PC[24]), .QN(n4831) );
  FD2 \pc_u0/pc_val_reg[25]  ( .D(\pc_u0/N29 ), .CP(clock), .CD(n4873), .Q(
        PC[25]), .QN(n4829) );
  FD2 \pc_u0/pc_val_reg[26]  ( .D(\pc_u0/N30 ), .CP(clock), .CD(n4873), .Q(
        PC[26]), .QN(n4841) );
  FD2 \pc_u0/pc_val_reg[27]  ( .D(\pc_u0/N31 ), .CP(clock), .CD(n4873), .Q(
        PC[27]), .QN(n4835) );
  FD2 \pc_u0/pc_val_reg[28]  ( .D(n1137), .CP(clock), .CD(n4873), .Q(PC[28]), 
        .QN(n4834) );
  FD2 \pc_u0/pc_val_reg[29]  ( .D(n1139), .CP(clock), .CD(n4873), .Q(PC[29]), 
        .QN(n4830) );
  FD2 \pc_u0/pc_val_reg[30]  ( .D(n1140), .CP(clock), .CD(n4873), .Q(PC[30]), 
        .QN(n4827) );
  FD2 \pc_u0/pc_val_reg[31]  ( .D(n1141), .CP(clock), .CD(n4873), .Q(PC[31]), 
        .QN(n4833) );
  FD4 \mw_Inst_reg[3]  ( .D(n1463), .CP(clock), .SD(n4873), .Q(n4823) );
  FD2 \dx_gpr_rd_data2_reg[15]  ( .D(gpr_rd_data2[15]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[15]) );
  FD2 \dx_gpr_rd_data2_reg[7]  ( .D(gpr_rd_data2[7]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data2[7]) );
  FD2 \dx_gpr_rd_data1_reg[28]  ( .D(gpr_rd_data1[28]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[28]) );
  FD2 \dx_gpr_rd_data1_reg[10]  ( .D(gpr_rd_data1[10]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[10]) );
  FD2 \dx_gpr_rd_data1_reg[2]  ( .D(gpr_rd_data1[2]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[2]) );
  FD2 \dx_gpr_rd_data1_reg[18]  ( .D(n1432), .CP(clock), .CD(n4873), .Q(
        dx_gpr_rd_data1[18]) );
  FD2 \dx_gpr_rd_data1_reg[12]  ( .D(gpr_rd_data1[12]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[12]) );
  FD2 \dx_gpr_rd_data1_reg[8]  ( .D(gpr_rd_data1[8]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[8]) );
  FD2 \dx_gpr_rd_data1_reg[31]  ( .D(n1434), .CP(clock), .CD(n4873), .Q(
        dx_gpr_rd_data1[31]) );
  FD2 \dx_gpr_rd_data1_reg[11]  ( .D(gpr_rd_data1[11]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[11]) );
  FD2 \dx_gpr_rd_data1_reg[4]  ( .D(gpr_rd_data1[4]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[4]) );
  FD2 \dx_gpr_rd_data1_reg[7]  ( .D(gpr_rd_data1[7]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[7]) );
  FD2 \dx_gpr_rd_data1_reg[15]  ( .D(gpr_rd_data1[15]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[15]) );
  FD2 \dx_gpr_rd_data1_reg[1]  ( .D(gpr_rd_data1[1]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[1]) );
  FD2 \dx_gpr_rd_data1_reg[29]  ( .D(gpr_rd_data1[29]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[29]) );
  FD2 \dx_gpr_rd_data1_reg[30]  ( .D(gpr_rd_data1[30]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[30]) );
  FD2 \dx_gpr_rd_data1_reg[27]  ( .D(gpr_rd_data1[27]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[27]) );
  FD2 \dx_gpr_rd_data1_reg[9]  ( .D(gpr_rd_data1[9]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[9]) );
  FD2 \dx_gpr_rd_data1_reg[0]  ( .D(gpr_rd_data1[0]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[0]) );
  FD2 \dx_gpr_rd_data1_reg[24]  ( .D(gpr_rd_data1[24]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[24]) );
  FD2 \dx_gpr_rd_data1_reg[21]  ( .D(gpr_rd_data1[21]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[21]) );
  FD2 \dx_gpr_rd_data1_reg[16]  ( .D(gpr_rd_data1[16]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[16]) );
  FD2 \dx_gpr_rd_data1_reg[23]  ( .D(gpr_rd_data1[23]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[23]) );
  FD2 \dx_gpr_rd_data1_reg[13]  ( .D(gpr_rd_data1[13]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[13]) );
  FD2 \dx_gpr_rd_data1_reg[22]  ( .D(gpr_rd_data1[22]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[22]) );
  FD2 \dx_gpr_rd_data1_reg[3]  ( .D(gpr_rd_data1[3]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[3]) );
  FD2 \dx_gpr_rd_data1_reg[19]  ( .D(gpr_rd_data1[19]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[19]) );
  FD2 \dx_gpr_rd_data1_reg[5]  ( .D(gpr_rd_data1[5]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[5]) );
  FD2 \dx_gpr_rd_data1_reg[25]  ( .D(gpr_rd_data1[25]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[25]) );
  FD2 \dx_gpr_rd_data1_reg[26]  ( .D(gpr_rd_data1[26]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[26]) );
  FD2 \dx_gpr_rd_data1_reg[6]  ( .D(gpr_rd_data1[6]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[6]) );
  FD2 \dx_gpr_rd_data1_reg[20]  ( .D(n1195), .CP(clock), .CD(n4873), .Q(
        dx_gpr_rd_data1[20]) );
  FD2 \dx_gpr_rd_data1_reg[17]  ( .D(gpr_rd_data1[17]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[17]) );
  FD2 \dx_gpr_rd_data1_reg[14]  ( .D(gpr_rd_data1[14]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_data1[14]) );
  FD2 \pc_u0/pc_val_reg[0]  ( .D(\pc_u0/N4 ), .CP(clock), .CD(n4873), .Q(
        \pc_u0/pc_plus_4 [0]) );
  FD4 \dx_gpr_rd_data2_reg[2]  ( .D(n4856), .CP(clock), .SD(n4873), .Q(n4821), 
        .QN(dx_gpr_rd_data2[2]) );
  FD4 \dx_gpr_rd_data2_reg[4]  ( .D(n4857), .CP(clock), .SD(n4873), .Q(n4819), 
        .QN(dx_gpr_rd_data2[4]) );
  FD4 \dx_Inst_15_0_signext_reg[31]  ( .D(n4715), .CP(clock), .SD(n4873), .Q(
        n4794), .QN(dx_Inst_15_0_signext[31]) );
  FD4 \mw_ALU_Result_reg[23]  ( .D(n4700), .CP(clock), .SD(n4873), .Q(n4740)
         );
  FD2 \mw_Inst_reg[11]  ( .D(xm_Inst[11]), .CP(clock), .CD(n4873), .Q(
        mw_Inst[11]) );
  FD2 \dx_gpr_rd_addr1_reg[2]  ( .D(gpr_rd_addr1[2]), .CP(clock), .CD(n4873), 
        .Q(dx_gpr_rd_addr1[2]) );
  FD2 \xm_ALU_Result_reg[2]  ( .D(x_ALU_Result[2]), .CP(clock), .CD(n4873), 
        .Q(Addr[2]) );
  FD2 \xm_ALU_Result_reg[7]  ( .D(x_ALU_Result[7]), .CP(clock), .CD(n4873), 
        .Q(Addr[7]) );
  FD2 \xm_ALU_Result_reg[3]  ( .D(x_ALU_Result[3]), .CP(clock), .CD(n4873), 
        .Q(Addr[3]) );
  FD2 \xm_ALU_Result_reg[11]  ( .D(x_ALU_Result[11]), .CP(clock), .CD(n4873), 
        .Q(Addr[11]) );
  FD2 \xm_ALU_Result_reg[4]  ( .D(x_ALU_Result[4]), .CP(clock), .CD(n4873), 
        .Q(Addr[4]) );
  FD2 \xm_ALU_Result_reg[0]  ( .D(x_ALU_Result[0]), .CP(clock), .CD(n4873), 
        .Q(Addr[0]) );
  FD2 \fd_Inst_reg[12]  ( .D(Inst_stall_b_j[12]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[12]) );
  FD2 \fd_Inst_reg[9]  ( .D(Inst_stall_b_j[9]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[9]) );
  FD2 \xm_ALU_Result_reg[17]  ( .D(x_ALU_Result[17]), .CP(clock), .CD(n4873), 
        .Q(Addr[17]) );
  FD2 \xm_ALU_Result_reg[10]  ( .D(x_ALU_Result[10]), .CP(clock), .CD(n4873), 
        .Q(Addr[10]) );
  FD2 \xm_ALU_Result_reg[16]  ( .D(x_ALU_Result[16]), .CP(clock), .CD(n4873), 
        .Q(Addr[16]) );
  FD2 \fd_Inst_reg[14]  ( .D(Inst_stall_b_j[14]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[14]) );
  FD2 \fd_Inst_reg[13]  ( .D(Inst_stall_b_j[13]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[13]) );
  FD2 \fd_Inst_reg[11]  ( .D(Inst_stall_b_j[11]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[11]) );
  FD2 \fd_Inst_reg[10]  ( .D(Inst_stall_b_j[10]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[10]) );
  FD2 \fd_Inst_reg[8]  ( .D(Inst_stall_b_j[8]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[8]) );
  FD2 \fd_Inst_reg[7]  ( .D(Inst_stall_b_j[7]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[7]) );
  FD2 \fd_Inst_reg[6]  ( .D(Inst_stall_b_j[6]), .CP(clock), .CD(n4873), .Q(
        fd_Inst[6]) );
  FD2 \xm_ALU_Result_reg[5]  ( .D(x_ALU_Result[5]), .CP(clock), .CD(n4873), 
        .Q(Addr[5]), .QN(n4703) );
  FD2 \xm_ALU_Result_reg[15]  ( .D(x_ALU_Result[15]), .CP(clock), .CD(n4873), 
        .Q(Addr[15]) );
  FD2 \xm_ALU_Result_reg[14]  ( .D(x_ALU_Result[14]), .CP(clock), .CD(n4873), 
        .Q(Addr[14]) );
  FD2 \xm_ALU_Result_reg[9]  ( .D(x_ALU_Result[9]), .CP(clock), .CD(n4873), 
        .Q(Addr[9]) );
  FD2 \xm_ALU_Result_reg[6]  ( .D(x_ALU_Result[6]), .CP(clock), .CD(n4873), 
        .Q(Addr[6]) );
  FD2 \xm_ALU_Result_reg[8]  ( .D(x_ALU_Result[8]), .CP(clock), .CD(n4873), 
        .Q(Addr[8]) );
  FD2 \pc_u0/pc_val_reg[2]  ( .D(\pc_u0/N6 ), .CP(clock), .CD(n4873), .Q(PC[2]), .QN(n1462) );
  FD2 \xm_ALU_Result_reg[23]  ( .D(x_ALU_Result[23]), .CP(clock), .CD(n4873), 
        .Q(Addr[23]), .QN(n4700) );
  FD2 \pc_u0/pc_val_reg[3]  ( .D(\pc_u0/N7 ), .CP(clock), .CD(n4873), .Q(PC[3]) );
  FD2 \pc_u0/pc_val_reg[1]  ( .D(\pc_u0/N5 ), .CP(clock), .CD(n4873), .Q(
        \pc_u0/pc_plus_4 [1]) );
  FD2 \xm_ALU_Result_reg[13]  ( .D(x_ALU_Result[13]), .CP(clock), .CD(n4873), 
        .Q(Addr[13]) );
  FD2 \xm_ALU_Result_reg[12]  ( .D(x_ALU_Result[12]), .CP(clock), .CD(n4873), 
        .Q(Addr[12]) );
  FD2 \xm_ALU_Result_reg[31]  ( .D(x_ALU_Result[31]), .CP(clock), .CD(n4873), 
        .Q(Addr[31]) );
  FD2 \xm_ALU_Result_reg[30]  ( .D(x_ALU_Result[30]), .CP(clock), .CD(n4873), 
        .Q(Addr[30]) );
  FD2 \xm_ALU_Result_reg[29]  ( .D(x_ALU_Result[29]), .CP(clock), .CD(n4873), 
        .Q(Addr[29]) );
  FD2 \xm_ALU_Result_reg[27]  ( .D(x_ALU_Result[27]), .CP(clock), .CD(n4873), 
        .Q(Addr[27]) );
  FD2 \xm_ALU_Result_reg[26]  ( .D(x_ALU_Result[26]), .CP(clock), .CD(n4873), 
        .Q(Addr[26]) );
  FD2 \xm_ALU_Result_reg[25]  ( .D(x_ALU_Result[25]), .CP(clock), .CD(n4873), 
        .Q(Addr[25]) );
  FD2 \xm_ALU_Result_reg[24]  ( .D(x_ALU_Result[24]), .CP(clock), .CD(n4873), 
        .Q(Addr[24]) );
  FD2 \xm_ALU_Result_reg[22]  ( .D(x_ALU_Result[22]), .CP(clock), .CD(n4873), 
        .Q(Addr[22]) );
  FD2 \xm_ALU_Result_reg[21]  ( .D(x_ALU_Result[21]), .CP(clock), .CD(n4873), 
        .Q(Addr[21]) );
  FD2 \xm_ALU_Result_reg[20]  ( .D(x_ALU_Result[20]), .CP(clock), .CD(n4873), 
        .Q(Addr[20]) );
  FD2 \xm_ALU_Result_reg[18]  ( .D(x_ALU_Result[18]), .CP(clock), .CD(n4873), 
        .Q(Addr[18]) );
  FD2 \xm_ALU_Result_reg[19]  ( .D(x_ALU_Result[19]), .CP(clock), .CD(n4873), 
        .Q(Addr[19]) );
  MUX21LP U1348 ( .A(n2901), .B(n2900), .S(n4626), .Z(n2915) );
  B4I U1349 ( .A(n2302), .Z(n2307) );
  B2IP U1350 ( .A(n2664), .Z2(n3918) );
  B2IP U1351 ( .A(n3118), .Z2(n1144) );
  IVI U1352 ( .A(n2300), .Z(n1145) );
  AO3P U1353 ( .A(n3908), .B(n4621), .C(n3131), .D(n3130), .Z(n3132) );
  AO3P U1354 ( .A(n4621), .B(n3837), .C(n2953), .D(n2952), .Z(n2954) );
  B4I U1355 ( .A(n4412), .Z(n4621) );
  ND2I U1356 ( .A(n2283), .B(n2098), .Z(n1146) );
  B4IP U1357 ( .A(n1146), .Z(n2296) );
  ND4P U1358 ( .A(n2875), .B(n2876), .C(n2873), .D(n2874), .Z(n3905) );
  ND4P U1359 ( .A(n4490), .B(n4299), .C(n4072), .D(n4015), .Z(n4257) );
  ND2I U1360 ( .A(n4490), .B(n4412), .Z(n1219) );
  IVDA U1361 ( .A(n3836), .Y(n1148), .Z(n1147) );
  ND2I U1362 ( .A(n1145), .B(n2668), .Z(n1149) );
  IVI U1363 ( .A(n2994), .Z(n1150) );
  IVI U1364 ( .A(n2994), .Z(n1151) );
  ND2I U1365 ( .A(n3876), .B(n3875), .Z(n1152) );
  B2I U1366 ( .A(n3900), .Z2(n1153) );
  ND2I U1367 ( .A(n2133), .B(n2132), .Z(n1154) );
  AO6 U1368 ( .A(n4353), .B(n4513), .C(n4371), .Z(n4384) );
  ND4P U1369 ( .A(n3177), .B(n3176), .C(n3175), .D(n3174), .Z(x_ALU_Result[8])
         );
  B2I U1370 ( .A(n4079), .Z2(n1155) );
  IVI U1371 ( .A(n2223), .Z(n1156) );
  IVI U1372 ( .A(n3925), .Z(n1157) );
  ND4P U1373 ( .A(n3794), .B(n3793), .C(n3792), .D(n3791), .Z(x_ALU_Result[13]) );
  B2I U1374 ( .A(n3796), .Z2(n1158) );
  AN2I U1375 ( .A(n2623), .B(n2624), .Z(n1159) );
  NR2I U1376 ( .A(n2212), .B(n1160), .Z(n2448) );
  ND2I U1377 ( .A(n1161), .B(n2214), .Z(n1160) );
  AN2I U1378 ( .A(n3221), .B(n3215), .Z(n1161) );
  ND2I U1379 ( .A(n1499), .B(n1498), .Z(n1162) );
  ND2I U1380 ( .A(n1484), .B(n2006), .Z(n1163) );
  ND2I U1381 ( .A(n4303), .B(n3013), .Z(n1217) );
  B2I U1382 ( .A(n4460), .Z2(n1164) );
  ND4P U1383 ( .A(n3055), .B(n3054), .C(n3053), .D(n3052), .Z(n1165) );
  ND4P U1384 ( .A(n2803), .B(n2804), .C(n1383), .D(n1384), .Z(n3185) );
  IVDA U1385 ( .A(n4220), .Z(n1166) );
  ND4 U1386 ( .A(n3111), .B(n3110), .C(n3109), .D(n3108), .Z(x_ALU_Result[9])
         );
  AN2I U1387 ( .A(n4637), .B(n4022), .Z(n1167) );
  IVI U1388 ( .A(n2109), .Z(n1168) );
  NR2I U1389 ( .A(n2842), .B(n2259), .Z(n1169) );
  AN2I U1390 ( .A(n4626), .B(n2409), .Z(n1170) );
  IVI U1391 ( .A(n3831), .Z(n1171) );
  ND4P U1392 ( .A(n4117), .B(n4555), .C(n4446), .D(n1217), .Z(n3874) );
  MUX21LP U1393 ( .A(n3133), .B(n3132), .S(n4626), .Z(n3134) );
  NR2I U1394 ( .A(n2045), .B(n2041), .Z(n2066) );
  IVI U1395 ( .A(n2116), .Z(n1172) );
  B2I U1396 ( .A(n4552), .Z2(n1173) );
  B2I U1397 ( .A(n3188), .Z1(n1175), .Z2(n1174) );
  IVI U1398 ( .A(n3807), .Z(n1176) );
  ND2I U1399 ( .A(n2903), .B(n2846), .Z(n1177) );
  IVI U1400 ( .A(n2861), .Z(n1178) );
  ND4 U1401 ( .A(n3082), .B(n3081), .C(n3080), .D(n3079), .Z(x_ALU_Result[15])
         );
  IVI U1402 ( .A(n3499), .Z(n1179) );
  ND2I U1403 ( .A(n2393), .B(n2392), .Z(n1180) );
  ND2I U1404 ( .A(n2393), .B(n2392), .Z(n1181) );
  MUX21LP U1405 ( .A(n2594), .B(n2595), .S(n2828), .Z(n2606) );
  ND2I U1406 ( .A(n2387), .B(n2386), .Z(n1182) );
  ND2I U1407 ( .A(n2387), .B(n2386), .Z(n1183) );
  ND2I U1408 ( .A(n2596), .B(n2607), .Z(n1184) );
  AN2I U1409 ( .A(n1309), .B(n1310), .Z(n1185) );
  B4IP U1410 ( .A(n1185), .Z(n4086) );
  B2I U1411 ( .A(n4191), .Z2(n4480) );
  B4I U1412 ( .A(n2365), .Z(n3118) );
  AO6P U1413 ( .A(n4357), .B(n4281), .C(n4250), .Z(n4253) );
  ND2I U1414 ( .A(n2525), .B(n2524), .Z(n1186) );
  ND2I U1415 ( .A(n2525), .B(n2524), .Z(n1187) );
  ND2I U1416 ( .A(n2614), .B(n2617), .Z(n1188) );
  IVI U1417 ( .A(n3831), .Z(n1189) );
  NR2I U1418 ( .A(n4344), .B(n4343), .Z(n1190) );
  MUX21LP U1419 ( .A(n2610), .B(n2609), .S(n3041), .Z(n2686) );
  MUX21LP U1420 ( .A(n2610), .B(n2609), .S(n3040), .Z(n2687) );
  IVI U1421 ( .A(n3697), .Z(n1191) );
  IVI U1422 ( .A(n3722), .Z(n1192) );
  IVDA U1423 ( .A(n4146), .Z(n1193) );
  MUX21LP U1424 ( .A(n4165), .B(n4164), .S(n4571), .Z(n1194) );
  AN2I U1425 ( .A(n4824), .B(n4825), .Z(n1516) );
  IVDA U1426 ( .A(gpr_rd_data1[20]), .Z(n1195) );
  AO6P U1427 ( .A(n4635), .B(n1387), .C(n1175), .Z(n2957) );
  IVI U1428 ( .A(n4471), .Z(n4169) );
  ENI U1429 ( .A(n4436), .B(n1196), .Z(n4471) );
  IVI U1430 ( .A(n1436), .Z(n1196) );
  ND2I U1431 ( .A(n1197), .B(n3259), .Z(n4436) );
  IVI U1432 ( .A(n3253), .Z(n3259) );
  AN2I U1433 ( .A(n3258), .B(n4146), .Z(n1197) );
  ND2I U1434 ( .A(n2683), .B(n3895), .Z(n1198) );
  ND2I U1435 ( .A(n1212), .B(n2362), .Z(n1199) );
  IVI U1436 ( .A(n2389), .Z(n1200) );
  IVI U1437 ( .A(n2389), .Z(n1201) );
  IVI U1438 ( .A(n2389), .Z(n1202) );
  IVI U1439 ( .A(n2389), .Z(n1203) );
  IVI U1440 ( .A(n2389), .Z(n1204) );
  IVI U1441 ( .A(n2389), .Z(n1205) );
  IVI U1442 ( .A(n1199), .Z(n1206) );
  IVI U1443 ( .A(n1199), .Z(n1207) );
  IVI U1444 ( .A(n1199), .Z(n1208) );
  IVI U1445 ( .A(n1199), .Z(n1209) );
  IVI U1446 ( .A(n1199), .Z(n1210) );
  IVI U1447 ( .A(n1199), .Z(n1211) );
  ND2I U1448 ( .A(n2340), .B(n2341), .Z(n1212) );
  ND2I U1449 ( .A(n2340), .B(n2341), .Z(n1213) );
  MUX21LP U1450 ( .A(n2641), .B(n2640), .S(n3891), .Z(n2683) );
  IVDA U1451 ( .A(n3762), .Z(n4797) );
  AO7 U1452 ( .A(n4398), .B(n4208), .C(n4642), .Z(n4209) );
  AO7 U1453 ( .A(n4644), .B(n4497), .C(n4643), .Z(n4498) );
  AO7 U1454 ( .A(n2197), .B(n2196), .C(n2262), .Z(n2198) );
  IVI U1455 ( .A(n1537), .Z(n3829) );
  IVI U1456 ( .A(n2781), .Z(n4672) );
  ND4 U1457 ( .A(n3050), .B(n3049), .C(n3048), .D(n3047), .Z(x_ALU_Result[14])
         );
  AO3 U1458 ( .A(n4669), .B(n2776), .C(n4041), .D(n2775), .Z(n2777) );
  IVI U1459 ( .A(n4854), .Z(n4702) );
  NR2 U1460 ( .A(dx_Inst_15_0_signext[3]), .B(dx_Inst_15_0_signext[4]), .Z(
        n1214) );
  ND4P U1461 ( .A(n2182), .B(n1214), .C(dx_Inst_15_0_signext[5]), .D(n2174), 
        .Z(n2197) );
  AO2P U1462 ( .A(Addr[29]), .B(n2544), .C(n4691), .D(n2539), .Z(n1215) );
  ND2 U1463 ( .A(n1211), .B(dx_gpr_rd_data1[29]), .Z(n1216) );
  ND2P U1464 ( .A(n1215), .B(n1216), .Z(n4601) );
  IVI U1465 ( .A(n4491), .Z(n1218) );
  AO3P U1466 ( .A(n1218), .B(n1219), .C(n4416), .D(n4415), .Z(n4417) );
  AO7 U1467 ( .A(n4021), .B(n4020), .C(n4642), .Z(n1220) );
  IVI U1468 ( .A(n4037), .Z(n1221) );
  AO2 U1469 ( .A(n4037), .B(n4313), .C(n4314), .D(n1221), .Z(n1222) );
  ND2I U1470 ( .A(n1222), .B(n4642), .Z(n1223) );
  AO2 U1471 ( .A(n4037), .B(n1220), .C(n4019), .D(n1223), .Z(n4025) );
  AO2 U1472 ( .A(n2526), .B(n2500), .C(n2514), .D(Addr[30]), .Z(n1224) );
  ND2I U1473 ( .A(n1200), .B(dx_gpr_rd_data1[30]), .Z(n1225) );
  ND2I U1474 ( .A(n1224), .B(n1225), .Z(n4653) );
  IVI U1475 ( .A(n3008), .Z(n1226) );
  AO2 U1476 ( .A(n3008), .B(n4640), .C(n4641), .D(n1226), .Z(n1227) );
  ND2I U1477 ( .A(n4642), .B(n1227), .Z(n1228) );
  ND2I U1478 ( .A(n2110), .B(n1228), .Z(n2974) );
  AN3 U1479 ( .A(n2707), .B(n3386), .C(n2491), .Z(n2908) );
  AO2 U1480 ( .A(n4632), .B(n4631), .C(n4630), .D(n4629), .Z(n1229) );
  AO2 U1481 ( .A(n4403), .B(n4633), .C(n4634), .D(n1144), .Z(n1230) );
  ND2I U1482 ( .A(n1229), .B(n1230), .Z(n1231) );
  ND2I U1483 ( .A(n4635), .B(n1231), .Z(n4636) );
  ND3 U1484 ( .A(n1540), .B(fd_Inst[27]), .C(n1538), .Z(n3418) );
  IVI U1485 ( .A(n2491), .Z(n1232) );
  NR2I U1486 ( .A(n3386), .B(n1232), .Z(n2706) );
  AO2 U1487 ( .A(n4634), .B(n3117), .C(n4631), .D(n4591), .Z(n1233) );
  AO2 U1488 ( .A(n4629), .B(n4592), .C(n4593), .D(n1144), .Z(n1234) );
  ND2I U1489 ( .A(n1233), .B(n1234), .Z(n4594) );
  AO2 U1490 ( .A(n2526), .B(n2504), .C(n2514), .D(Addr[31]), .Z(n1235) );
  ND2 U1491 ( .A(n1210), .B(dx_gpr_rd_data1[31]), .Z(n1236) );
  ND2I U1492 ( .A(n1235), .B(n1236), .Z(n4650) );
  ND2I U1493 ( .A(n3739), .B(PC[18]), .Z(n1237) );
  EOI U1494 ( .A(n4750), .B(n1237), .Z(\pc_u0/pc_plus_4 [19]) );
  IVI U1495 ( .A(n4565), .Z(n1238) );
  AO2 U1496 ( .A(n4565), .B(n4640), .C(n4641), .D(n1238), .Z(n1239) );
  ND2I U1497 ( .A(n1239), .B(n4642), .Z(n1240) );
  ND2I U1498 ( .A(n4534), .B(n1240), .Z(n4537) );
  ND4 U1499 ( .A(n4014), .B(n3166), .C(n3163), .D(n3164), .Z(n3937) );
  IV U1500 ( .A(n3554), .Z(n1241) );
  IVI U1501 ( .A(n3739), .Z(n1242) );
  MUX31L U1502 ( .D0(n3554), .D1(n1241), .D2(n4843), .A(PC[20]), .B(n1242), 
        .Z(\pc_u0/pc_plus_4 [20]) );
  ND4 U1503 ( .A(n3016), .B(n3015), .C(n2949), .D(n2950), .Z(n3849) );
  AO7 U1504 ( .A(n3271), .B(n4020), .C(n4642), .Z(n1243) );
  IVI U1505 ( .A(n2945), .Z(n1244) );
  AO2 U1506 ( .A(n2945), .B(n4313), .C(n4314), .D(n1244), .Z(n1245) );
  ND2I U1507 ( .A(n1245), .B(n4642), .Z(n1246) );
  AO2 U1508 ( .A(n2945), .B(n1243), .C(n3271), .D(n1246), .Z(n2745) );
  AO2 U1509 ( .A(n3350), .B(n3117), .C(n4591), .D(n3371), .Z(n1247) );
  AO2 U1510 ( .A(n4592), .B(n3365), .C(n3351), .D(n1144), .Z(n1248) );
  ND2I U1511 ( .A(n1247), .B(n1248), .Z(n3119) );
  AO2 U1512 ( .A(n2515), .B(n4677), .C(n2514), .D(Addr[1]), .Z(n1249) );
  ND2 U1513 ( .A(dx_gpr_rd_data1[1]), .B(n1202), .Z(n1250) );
  ND2I U1514 ( .A(n1249), .B(n1250), .Z(n2966) );
  ND2I U1515 ( .A(n4295), .B(n4646), .Z(n1251) );
  ND2I U1516 ( .A(n4331), .B(n4511), .Z(n1252) );
  ND3P U1517 ( .A(n4296), .B(n1251), .C(n1252), .Z(n4301) );
  IV U1518 ( .A(n4837), .Z(n1253) );
  MUX31L U1519 ( .D0(n1253), .D1(n4837), .D2(PC[21]), .A(PC[20]), .B(n3554), 
        .Z(n1254) );
  EO1 U1520 ( .A(n3739), .B(n1254), .C(n1253), .D(n3739), .Z(
        \pc_u0/pc_plus_4 [21]) );
  ND2I U1521 ( .A(dx_gpr_rd_data1[13]), .B(n1205), .Z(n1255) );
  ND3P U1522 ( .A(n2417), .B(n2416), .C(n1255), .Z(n3781) );
  AO7P U1523 ( .A(n3210), .B(n3205), .C(n3204), .Z(n1256) );
  ND2I U1524 ( .A(n3212), .B(n1256), .Z(n1257) );
  ND2I U1525 ( .A(n1257), .B(n3207), .Z(n1258) );
  NR2 U1526 ( .A(n3208), .B(n3209), .Z(n1259) );
  NR2I U1527 ( .A(n1258), .B(n1259), .Z(n3237) );
  IVI U1528 ( .A(n3929), .Z(n1260) );
  AO2 U1529 ( .A(n3929), .B(n4640), .C(n4641), .D(n1260), .Z(n1261) );
  ND2I U1530 ( .A(n1261), .B(n4642), .Z(n1262) );
  AO7 U1531 ( .A(n3928), .B(n4020), .C(n4643), .Z(n1263) );
  AO2 U1532 ( .A(n3928), .B(n1262), .C(n3929), .D(n1263), .Z(n3934) );
  IVI U1533 ( .A(n2708), .Z(n1264) );
  AO6 U1534 ( .A(n2707), .B(n2706), .C(n1264), .Z(n2781) );
  IVI U1535 ( .A(n2781), .Z(n4041) );
  AO2 U1536 ( .A(n2951), .B(n3364), .C(n4591), .D(n3358), .Z(n1265) );
  AO2 U1537 ( .A(n3186), .B(n3356), .C(n3365), .D(n3013), .Z(n1266) );
  ND2I U1538 ( .A(n1265), .B(n1266), .Z(n1267) );
  ND2I U1539 ( .A(n4635), .B(n1267), .Z(n3187) );
  IV U1540 ( .A(n4836), .Z(n1268) );
  MUX31L U1541 ( .D0(n1268), .D1(n4836), .D2(PC[23]), .A(PC[22]), .B(n3580), 
        .Z(n1269) );
  EO1 U1542 ( .A(n3739), .B(n1269), .C(n1268), .D(n3739), .Z(
        \pc_u0/pc_plus_4 [23]) );
  IVI U1543 ( .A(n2319), .Z(n1270) );
  ND2I U1544 ( .A(n4686), .B(n1270), .Z(n2136) );
  IV U1545 ( .A(n4653), .Z(n1271) );
  AO2 U1546 ( .A(n4653), .B(n4640), .C(n4641), .D(n1271), .Z(n1272) );
  ND2 U1547 ( .A(n1272), .B(n4643), .Z(n1273) );
  AO7 U1548 ( .A(n4604), .B(n4644), .C(n4643), .Z(n1274) );
  AO2 U1549 ( .A(n4604), .B(n1273), .C(n4653), .D(n1274), .Z(n1275) );
  ND2I U1550 ( .A(n4598), .B(n4646), .Z(n1276) );
  ND2I U1551 ( .A(n1275), .B(n1276), .Z(n4599) );
  ND4 U1552 ( .A(n3169), .B(n3170), .C(n3167), .D(n3168), .Z(n3942) );
  IV U1553 ( .A(n2959), .Z(n1277) );
  AO2 U1554 ( .A(n2959), .B(n1440), .C(n3138), .D(n1277), .Z(n1278) );
  ENI U1555 ( .A(n3137), .B(n1278), .Z(n1279) );
  ENI U1556 ( .A(n1279), .B(n3136), .Z(n3139) );
  IV U1557 ( .A(n4831), .Z(n1280) );
  MUX31L U1558 ( .D0(n4831), .D1(n1280), .D2(PC[24]), .A(n3596), .B(n3580), 
        .Z(n1281) );
  EO1 U1559 ( .A(n3739), .B(n1281), .C(n1280), .D(n3739), .Z(
        \pc_u0/pc_plus_4 [24]) );
  AN4P U1560 ( .A(n4297), .B(n4299), .C(n4300), .D(n4298), .Z(n4584) );
  AO2 U1561 ( .A(n2526), .B(n2499), .C(n2514), .D(Addr[27]), .Z(n1282) );
  ND2 U1562 ( .A(n1202), .B(dx_gpr_rd_data1[27]), .Z(n1283) );
  ND2I U1563 ( .A(n1282), .B(n1283), .Z(n4565) );
  AO7 U1564 ( .A(n3361), .B(n3360), .C(n3359), .Z(n1284) );
  AN2I U1565 ( .A(n3370), .B(n1284), .Z(n1285) );
  NR2 U1566 ( .A(n3928), .B(n3371), .Z(n1286) );
  NR2 U1567 ( .A(n3372), .B(n1286), .Z(n1287) );
  AO3 U1568 ( .A(n1285), .B(n3369), .C(n3373), .D(n1287), .Z(n3374) );
  ND4 U1569 ( .A(n2888), .B(n2889), .C(n2886), .D(n2887), .Z(n3763) );
  AO7 U1570 ( .A(n4649), .B(n4644), .C(n4643), .Z(n1288) );
  IVI U1571 ( .A(n4650), .Z(n1289) );
  AO2 U1572 ( .A(n4650), .B(n4640), .C(n4641), .D(n1289), .Z(n1290) );
  ND2I U1573 ( .A(n1290), .B(n4642), .Z(n1291) );
  AO2 U1574 ( .A(n4650), .B(n1288), .C(n4649), .D(n1291), .Z(n1292) );
  ND2I U1575 ( .A(n4646), .B(n4645), .Z(n1293) );
  ND2I U1576 ( .A(n1292), .B(n1293), .Z(n4647) );
  ND2I U1577 ( .A(n4630), .B(n2966), .Z(n1294) );
  ND3P U1578 ( .A(n2965), .B(n2964), .C(n1294), .Z(n4336) );
  IV U1579 ( .A(n3482), .Z(n1295) );
  IV U1580 ( .A(n3754), .Z(n1296) );
  MUX31L U1581 ( .D0(n1295), .D1(n3482), .D2(n3483), .A(n3751), .B(n1296), .Z(
        n1297) );
  ND2I U1582 ( .A(n3637), .B(n1297), .Z(n3484) );
  ND2 U1583 ( .A(n3514), .B(PC[10]), .Z(n1298) );
  EO U1584 ( .A(n4751), .B(n1298), .Z(\pc_u0/pc_plus_4 [11]) );
  IV U1585 ( .A(n4829), .Z(n1299) );
  MUX31L U1586 ( .D0(n1299), .D1(n4829), .D2(PC[25]), .A(PC[24]), .B(n3596), 
        .Z(n1300) );
  ND2I U1587 ( .A(n3597), .B(n3739), .Z(n1301) );
  MUX21L U1588 ( .A(n1300), .B(n4829), .S(n1301), .Z(\pc_u0/pc_plus_4 [25]) );
  IVI U1589 ( .A(n2827), .Z(n1302) );
  ND2I U1590 ( .A(n2595), .B(n1302), .Z(n1303) );
  ND2I U1591 ( .A(n2827), .B(n2594), .Z(n1304) );
  ND2I U1592 ( .A(n1303), .B(n1304), .Z(n2607) );
  ND2 U1593 ( .A(n2110), .B(n3350), .Z(n1305) );
  ND2 U1594 ( .A(n3371), .B(n3928), .Z(n1306) );
  AO7 U1595 ( .A(n3372), .B(n1306), .C(n1305), .Z(n1307) );
  AO7 U1596 ( .A(n3355), .B(n3354), .C(n3353), .Z(n1308) );
  AO6 U1597 ( .A(n3373), .B(n1307), .C(n1308), .Z(n3375) );
  AN2I U1598 ( .A(n4297), .B(n4277), .Z(n3921) );
  AO2 U1599 ( .A(n2545), .B(n2450), .C(n2544), .D(Addr[19]), .Z(n1309) );
  ND2 U1600 ( .A(dx_gpr_rd_data1[19]), .B(n1208), .Z(n1310) );
  AO2 U1601 ( .A(n2292), .B(n4690), .C(n2310), .D(Addr[28]), .Z(n1311) );
  AN2I U1602 ( .A(n1311), .B(n4146), .Z(n4139) );
  ND4 U1603 ( .A(n4013), .B(n3014), .C(n4071), .D(n2946), .Z(n3836) );
  EN U1604 ( .A(n3747), .B(n3631), .Z(n3632) );
  EN U1605 ( .A(n3519), .B(n3521), .Z(n3525) );
  AO2 U1606 ( .A(n4402), .B(n4401), .C(n4400), .D(n4593), .Z(n1312) );
  AO2 U1607 ( .A(n4403), .B(n4634), .C(n4404), .D(n3013), .Z(n1313) );
  ND2I U1608 ( .A(n1312), .B(n1313), .Z(n1314) );
  ND2I U1609 ( .A(n4635), .B(n1314), .Z(n4405) );
  AO2P U1610 ( .A(n4517), .B(n3795), .C(n4512), .D(n3161), .Z(n1315) );
  AN2I U1611 ( .A(n3162), .B(n1315), .Z(n3177) );
  IVI U1612 ( .A(n2963), .Z(n1316) );
  AO2 U1613 ( .A(n2963), .B(n4640), .C(n4641), .D(n1316), .Z(n1317) );
  ND2I U1614 ( .A(n4643), .B(n1317), .Z(n1318) );
  ND2I U1615 ( .A(n3918), .B(n1318), .Z(n2917) );
  IV U1616 ( .A(n3463), .Z(n1319) );
  IV U1617 ( .A(n3526), .Z(n1320) );
  MUX31L U1618 ( .D0(n1319), .D1(n3463), .D2(n3464), .A(n3523), .B(n1320), .Z(
        n1321) );
  ND2I U1619 ( .A(n3576), .B(n1321), .Z(n3465) );
  IVI U1620 ( .A(n2903), .Z(n1322) );
  NR2I U1621 ( .A(n2902), .B(n1322), .Z(n3188) );
  IV U1622 ( .A(PC[9]), .Z(n1323) );
  MUX31L U1623 ( .D0(n1323), .D1(PC[9]), .D2(n4845), .A(PC[8]), .B(n3723), .Z(
        n1324) );
  EO1 U1624 ( .A(n3724), .B(n1324), .C(n1323), .D(n3724), .Z(n3958) );
  IV U1625 ( .A(n4840), .Z(n1325) );
  MUX31L U1626 ( .D0(n1325), .D1(n4840), .D2(PC[13]), .A(PC[12]), .B(n3487), 
        .Z(n1326) );
  EO1 U1627 ( .A(n3514), .B(n1326), .C(n1325), .D(n3514), .Z(
        \pc_u0/pc_plus_4 [13]) );
  IV U1628 ( .A(n3738), .Z(n1327) );
  IVI U1629 ( .A(n3739), .Z(n1328) );
  MUX31L U1630 ( .D0(n3738), .D1(n1327), .D2(n4841), .A(PC[26]), .B(n1328), 
        .Z(\pc_u0/pc_plus_4 [26]) );
  IVI U1631 ( .A(n4504), .Z(n1329) );
  ND2 U1632 ( .A(n4502), .B(n4334), .Z(n1330) );
  AO3P U1633 ( .A(n1329), .B(n1330), .C(n4024), .D(n4025), .Z(n4026) );
  ENI U1634 ( .A(n4571), .B(n4305), .Z(n4306) );
  EN U1635 ( .A(n3746), .B(n3631), .Z(n3633) );
  EN U1636 ( .A(n3520), .B(n3521), .Z(n3524) );
  AO2 U1637 ( .A(n2526), .B(n4690), .C(n2521), .D(Addr[28]), .Z(n1331) );
  ND2 U1638 ( .A(n1206), .B(dx_gpr_rd_data1[28]), .Z(n1332) );
  ND2I U1639 ( .A(n1331), .B(n1332), .Z(n4424) );
  IV U1640 ( .A(n1461), .Z(n1333) );
  ND2 U1641 ( .A(mw_pc_plus_8[17]), .B(n1333), .Z(n1334) );
  ND2I U1642 ( .A(n1461), .B(n4685), .Z(n1335) );
  ND2I U1643 ( .A(n1334), .B(n1335), .Z(gpr_wr_data[17]) );
  AO7 U1644 ( .A(n4142), .B(n4398), .C(n4642), .Z(n1336) );
  AO2 U1645 ( .A(n4142), .B(n4136), .C(n4601), .D(n1336), .Z(n1337) );
  ND2I U1646 ( .A(n1151), .B(n4353), .Z(n1338) );
  ND2I U1647 ( .A(n1337), .B(n1338), .Z(n4137) );
  EO U1648 ( .A(fd_Inst[1]), .B(PC[3]), .Z(n1339) );
  EN U1649 ( .A(n3668), .B(n1339), .Z(n3669) );
  ND4 U1650 ( .A(n2892), .B(n2893), .C(n2890), .D(n2891), .Z(n3097) );
  IVI U1651 ( .A(n4541), .Z(n4254) );
  AO2 U1652 ( .A(n3007), .B(n3365), .C(n4124), .D(n3364), .Z(n1340) );
  AO2 U1653 ( .A(n2904), .B(n3358), .C(n3013), .D(n3371), .Z(n1341) );
  ND2I U1654 ( .A(n1340), .B(n1341), .Z(n1342) );
  ND2I U1655 ( .A(n4635), .B(n1342), .Z(n2905) );
  IV U1656 ( .A(PC[6]), .Z(n1343) );
  MUX31L U1657 ( .D0(n1343), .D1(PC[6]), .D2(n4851), .A(PC[7]), .B(n3709), .Z(
        \pc_u0/pc_plus_4 [7]) );
  IV U1658 ( .A(n4839), .Z(n1344) );
  MUX31L U1659 ( .D0(n1344), .D1(n4839), .D2(PC[15]), .A(PC[14]), .B(n3513), 
        .Z(n1345) );
  EO1 U1660 ( .A(n3514), .B(n1345), .C(n1344), .D(n3514), .Z(
        \pc_u0/pc_plus_4 [15]) );
  IV U1661 ( .A(n4835), .Z(n1346) );
  MUX31L U1662 ( .D0(n1346), .D1(n4835), .D2(PC[27]), .A(PC[26]), .B(n3738), 
        .Z(n1347) );
  EO1 U1663 ( .A(n3739), .B(n1347), .C(n1346), .D(n3739), .Z(
        \pc_u0/pc_plus_4 [27]) );
  NR2I U1664 ( .A(mw_Inst[29]), .B(mw_Inst[28]), .Z(n1348) );
  AN2I U1665 ( .A(n1466), .B(n1348), .Z(n1515) );
  ND2I U1666 ( .A(dx_gpr_rd_data2[24]), .B(n3254), .Z(n1349) );
  AN2I U1667 ( .A(n4146), .B(n1349), .Z(n3220) );
  IV U1668 ( .A(n2147), .Z(n1350) );
  NR2I U1669 ( .A(n3303), .B(n1350), .Z(n3318) );
  ND2I U1670 ( .A(n3330), .B(n4246), .Z(n1351) );
  EON1 U1671 ( .A(n3333), .B(n1351), .C(n3332), .D(n3331), .Z(n3334) );
  ND2I U1672 ( .A(n2668), .B(n1145), .Z(n1352) );
  ENI U1673 ( .A(n1436), .B(n1352), .Z(n3189) );
  ND4P U1674 ( .A(n2878), .B(n2879), .C(n4110), .D(n2877), .Z(n3907) );
  IV U1675 ( .A(n3600), .Z(n1353) );
  AO1 U1676 ( .A(PC[25]), .B(n3599), .C(n3604), .D(n1353), .Z(n1354) );
  ND2I U1677 ( .A(n1354), .B(n3608), .Z(n3751) );
  EOI U1678 ( .A(n4662), .B(n4426), .Z(n4427) );
  IV U1679 ( .A(n1461), .Z(n1355) );
  ND2 U1680 ( .A(mw_pc_plus_8[29]), .B(n1355), .Z(n1356) );
  ND2I U1681 ( .A(n1461), .B(n4691), .Z(n1357) );
  ND2I U1682 ( .A(n1356), .B(n1357), .Z(gpr_wr_data[29]) );
  AO6 U1683 ( .A(n4492), .B(n4493), .C(n4509), .Z(n4523) );
  EO U1684 ( .A(n2998), .B(n3008), .Z(n1358) );
  IV U1685 ( .A(n2999), .Z(n1359) );
  MUX21L U1686 ( .A(n1359), .B(n3000), .S(n1451), .Z(n1360) );
  ENI U1687 ( .A(n1358), .B(n1360), .Z(n3002) );
  IVI U1688 ( .A(n4548), .Z(n4261) );
  AN3 U1689 ( .A(n4048), .B(n4046), .C(n4047), .Z(n1361) );
  IV U1690 ( .A(n1177), .Z(n1362) );
  AO2 U1691 ( .A(n3927), .B(n4251), .C(n1361), .D(n1362), .Z(n3941) );
  EN U1692 ( .A(fd_Inst[3]), .B(PC[5]), .Z(n1363) );
  MUX21L U1693 ( .A(n3681), .B(n3682), .S(n3683), .Z(n1364) );
  EN U1694 ( .A(n1363), .B(n1364), .Z(n3684) );
  IVI U1695 ( .A(n2966), .Z(n1365) );
  AO2 U1696 ( .A(n2966), .B(n4640), .C(n4641), .D(n1365), .Z(n1366) );
  AO7 U1697 ( .A(n3357), .B(n4317), .C(n4643), .Z(n1367) );
  ND2 U1698 ( .A(n2966), .B(n1367), .Z(n1368) );
  ND2I U1699 ( .A(n1366), .B(n4642), .Z(n1369) );
  ND2I U1700 ( .A(n3357), .B(n1369), .Z(n1370) );
  ND2I U1701 ( .A(n1370), .B(n1368), .Z(n2910) );
  IV U1702 ( .A(PC[8]), .Z(n1371) );
  MUX31L U1703 ( .D0(PC[8]), .D1(n1371), .D2(n4850), .A(n3723), .B(n3709), .Z(
        \pc_u0/pc_plus_4 [8]) );
  IV U1704 ( .A(n4838), .Z(n1372) );
  MUX31L U1705 ( .D0(n4838), .D1(n1372), .D2(PC[16]), .A(n3512), .B(n3513), 
        .Z(n1373) );
  EO1 U1706 ( .A(n3514), .B(n1373), .C(n1372), .D(n3514), .Z(
        \pc_u0/pc_plus_4 [16]) );
  IV U1707 ( .A(n4834), .Z(n1374) );
  MUX31L U1708 ( .D0(n4834), .D1(n1374), .D2(PC[28]), .A(n3737), .B(n3738), 
        .Z(n1375) );
  EO1 U1709 ( .A(n3739), .B(n1375), .C(n1374), .D(n3739), .Z(
        \pc_u0/pc_plus_4 [28]) );
  NR4 U1710 ( .A(fd_Inst[23]), .B(fd_Inst[25]), .C(fd_Inst[24]), .D(
        fd_Inst[22]), .Z(n1376) );
  ND2I U1711 ( .A(n1376), .B(n4759), .Z(n1532) );
  ND2 U1712 ( .A(PC[30]), .B(n3742), .Z(n1377) );
  EO U1713 ( .A(n3648), .B(n1377), .Z(n3651) );
  ENI U1714 ( .A(n4090), .B(n2691), .Z(n2713) );
  ENI U1715 ( .A(n4476), .B(n4345), .Z(n4346) );
  ND2I U1716 ( .A(n3248), .B(dx_gpr_rd_data2[29]), .Z(n1378) );
  ND4P U1717 ( .A(n4146), .B(n2069), .C(n2070), .D(n1378), .Z(n4142) );
  ENI U1718 ( .A(n3784), .B(n3785), .Z(n3786) );
  EOI U1719 ( .A(n1436), .B(n3194), .Z(n1379) );
  ENI U1720 ( .A(n3189), .B(n1379), .Z(n3190) );
  ENI U1721 ( .A(n2828), .B(n2829), .Z(n2853) );
  EN U1722 ( .A(n3603), .B(n3585), .Z(n3588) );
  EN U1723 ( .A(n3730), .B(n3714), .Z(n3716) );
  IV U1724 ( .A(n1461), .Z(n1380) );
  ND2 U1725 ( .A(mw_pc_plus_8[4]), .B(n1380), .Z(n1381) );
  ND2I U1726 ( .A(n1461), .B(n4678), .Z(n1382) );
  ND2I U1727 ( .A(n1381), .B(n1382), .Z(gpr_wr_data[4]) );
  ND4P U1728 ( .A(n3850), .B(n3851), .C(n3838), .D(n3839), .Z(n3866) );
  ND2 U1729 ( .A(n1445), .B(n4517), .Z(n1383) );
  ND2I U1730 ( .A(n4583), .B(n4512), .Z(n1384) );
  AO2 U1731 ( .A(n4591), .B(n3365), .C(n3371), .D(n3117), .Z(n1385) );
  AO2 U1732 ( .A(n1144), .B(n3350), .C(n2922), .D(n3364), .Z(n1386) );
  ND2I U1733 ( .A(n1386), .B(n1385), .Z(n1387) );
  EOI U1734 ( .A(n2906), .B(n2907), .Z(n1388) );
  ENI U1735 ( .A(n2966), .B(n1388), .Z(n2911) );
  IV U1736 ( .A(n4424), .Z(n1389) );
  AO2 U1737 ( .A(n4424), .B(n4640), .C(n4641), .D(n1389), .Z(n1390) );
  ND2I U1738 ( .A(n4642), .B(n1390), .Z(n1391) );
  AO7 U1739 ( .A(n4399), .B(n4398), .C(n4643), .Z(n1392) );
  AO2 U1740 ( .A(n4397), .B(n1391), .C(n4424), .D(n1392), .Z(n4423) );
  IV U1741 ( .A(PC[4]), .Z(n1393) );
  MUX31L U1742 ( .D0(n1393), .D1(PC[4]), .D2(PC[5]), .A(n4844), .B(n3679), .Z(
        n3957) );
  IVI U1743 ( .A(PC[17]), .Z(n1394) );
  MUX31L U1744 ( .D0(n1394), .D1(PC[17]), .D2(n4832), .A(PC[16]), .B(n3512), 
        .Z(n1395) );
  EO1 U1745 ( .A(n3456), .B(n1395), .C(n1394), .D(n3456), .Z(n1396) );
  IV U1746 ( .A(n3414), .Z(n1397) );
  AO2 U1747 ( .A(n3414), .B(n4832), .C(n1396), .D(n1397), .Z(
        \pc_u0/pc_plus_4 [17]) );
  NR2I U1748 ( .A(n3737), .B(n3738), .Z(n1398) );
  ND2 U1749 ( .A(n4830), .B(PC[28]), .Z(n1399) );
  AO3 U1750 ( .A(n4830), .B(PC[28]), .C(n1398), .D(n1399), .Z(n1400) );
  AO7 U1751 ( .A(PC[29]), .B(n1398), .C(n1400), .Z(n1401) );
  IVI U1752 ( .A(n3739), .Z(n1402) );
  AO2 U1753 ( .A(n3739), .B(n1401), .C(n4830), .D(n1402), .Z(
        \pc_u0/pc_plus_4 [29]) );
  IVI U1754 ( .A(gpr_rd_data1[14]), .Z(n1596) );
  IV U1755 ( .A(n4695), .Z(n1403) );
  ND2 U1756 ( .A(n4696), .B(n4825), .Z(n1404) );
  ND2 U1757 ( .A(n4701), .B(n4694), .Z(n1405) );
  AO4 U1758 ( .A(n4701), .B(n1404), .C(n1403), .D(n1405), .Z(n1406) );
  NR4 U1759 ( .A(mw_Inst[16]), .B(mw_Inst[17]), .C(mw_Inst[11]), .D(
        mw_Inst[13]), .Z(n1407) );
  NR4 U1760 ( .A(mw_Inst[15]), .B(mw_Inst[20]), .C(mw_Inst[14]), .D(
        mw_Inst[18]), .Z(n1408) );
  NR4 U1761 ( .A(mw_Inst[19]), .B(mw_Inst[23]), .C(mw_Inst[24]), .D(
        mw_Inst[25]), .Z(n1409) );
  ND3 U1762 ( .A(n1407), .B(n1408), .C(n1409), .Z(n1410) );
  NR4 U1763 ( .A(mw_Inst[12]), .B(mw_Inst[22]), .C(mw_Inst[21]), .D(n1410), 
        .Z(n1411) );
  OR3 U1764 ( .A(n4823), .B(mw_Inst_2), .C(mw_Inst_4), .Z(n1412) );
  NR4 U1765 ( .A(mw_Inst_5), .B(mw_Inst_0), .C(mw_Inst_1), .D(n1412), .Z(n1413) );
  ND2 U1766 ( .A(n4693), .B(n4824), .Z(n1414) );
  NR2 U1767 ( .A(n1413), .B(n4692), .Z(n1415) );
  NR2 U1768 ( .A(n1414), .B(n1415), .Z(n1416) );
  AO1 U1769 ( .A(n1406), .B(n4826), .C(n1411), .D(n1416), .Z(w_RegWrite) );
  IV U1770 ( .A(n3342), .Z(n1417) );
  IV U1771 ( .A(n3343), .Z(n1418) );
  AO3 U1772 ( .A(n3341), .B(n1417), .C(n3344), .D(n1418), .Z(n3346) );
  NR2 U1773 ( .A(n3742), .B(PC[30]), .Z(n1419) );
  EO U1774 ( .A(n1419), .B(n3648), .Z(n3652) );
  EN U1775 ( .A(n4036), .B(n4037), .Z(n4038) );
  EN U1776 ( .A(n4475), .B(n4345), .Z(n4347) );
  EN U1777 ( .A(n4570), .B(n4305), .Z(n4307) );
  EN U1778 ( .A(n3604), .B(n3585), .Z(n3589) );
  NR4 U1779 ( .A(fd_Inst[0]), .B(fd_Inst[2]), .C(fd_Inst[5]), .D(fd_Inst[27]), 
        .Z(n1420) );
  IV U1780 ( .A(fd_Inst[3]), .Z(n1421) );
  NR4 U1781 ( .A(fd_Inst[4]), .B(fd_Inst[28]), .C(n1465), .D(n1421), .Z(n1422)
         );
  IV U1782 ( .A(fd_Inst[26]), .Z(n1423) );
  ND4 U1783 ( .A(n4828), .B(n1420), .C(n1422), .D(n1423), .Z(n1537) );
  EN U1784 ( .A(n2770), .B(n2773), .Z(n2776) );
  AO2 U1785 ( .A(n4511), .B(n3943), .C(n4513), .D(n3942), .Z(n3946) );
  EO U1786 ( .A(PC[9]), .B(fd_Inst[7]), .Z(n1424) );
  EN U1787 ( .A(n3729), .B(n1424), .Z(n1425) );
  EN U1788 ( .A(n3728), .B(n1424), .Z(n1426) );
  IV U1789 ( .A(n3731), .Z(n1427) );
  AO2 U1790 ( .A(n3731), .B(n1425), .C(n1426), .D(n1427), .Z(n1428) );
  IV U1791 ( .A(n3730), .Z(n1429) );
  AO2 U1792 ( .A(n3730), .B(n1425), .C(n1426), .D(n1429), .Z(n1430) );
  IV U1793 ( .A(n3732), .Z(n1431) );
  AO2 U1794 ( .A(n3732), .B(n1428), .C(n1430), .D(n1431), .Z(n3733) );
  EO U1795 ( .A(n3679), .B(n4853), .Z(\pc_u0/pc_plus_4 [4]) );
  IVI U1796 ( .A(gpr_rd_data1[18]), .Z(n1432) );
  IVI U1797 ( .A(gpr_rd_data1[18]), .Z(n1433) );
  IVI U1798 ( .A(gpr_rd_data1[31]), .Z(n1434) );
  IVI U1799 ( .A(gpr_rd_data1[31]), .Z(n1435) );
  B4IP U1800 ( .A(n2669), .Z(n1436) );
  AN2I U1801 ( .A(n2682), .B(n2681), .Z(n1437) );
  OR2P U1802 ( .A(n2907), .B(n2966), .Z(n1438) );
  B4IP U1803 ( .A(n2908), .Z(n4642) );
  B4IP U1804 ( .A(n2908), .Z(n4643) );
  AN2I U1805 ( .A(n2844), .B(n2449), .Z(n1439) );
  AN2I U1806 ( .A(n2677), .B(n3364), .Z(n1440) );
  IVDA U1807 ( .A(mw_Inst[31]), .Y(n1441), .Z(n1526) );
  AN2I U1808 ( .A(n2111), .B(n3348), .Z(n1442) );
  ND2I U1809 ( .A(n2485), .B(n2213), .Z(n1443) );
  AN2I U1810 ( .A(n4506), .B(n4505), .Z(n1444) );
  AN2I U1811 ( .A(n3871), .B(n3031), .Z(n1445) );
  IVDA U1812 ( .A(n3843), .Y(n1451) );
  AN2I U1813 ( .A(n2695), .B(n2692), .Z(n1452) );
  AN2I U1814 ( .A(n2292), .B(n2401), .Z(n1453) );
  MUX21L U1815 ( .A(n1188), .B(n2641), .S(n3840), .Z(n2832) );
  AN2I U1816 ( .A(n4075), .B(n4074), .Z(n1455) );
  IVI U1817 ( .A(n2110), .Z(n3348) );
  B2IP U1818 ( .A(n2060), .Z1(n1460), .Z2(n1461) );
  IVI U1819 ( .A(n4855), .Z(n1994) );
  IVI U1820 ( .A(n4101), .Z(n4102) );
  IVI U1821 ( .A(n2680), .Z(n2681) );
  IVI U1822 ( .A(n2671), .Z(n2672) );
  IVI U1823 ( .A(n2650), .Z(n2642) );
  IVI U1824 ( .A(n2832), .Z(n2684) );
  IVI U1825 ( .A(n2589), .Z(n2590) );
  IVI U1826 ( .A(n3324), .Z(n2597) );
  IVI U1827 ( .A(n3100), .Z(n2598) );
  NR2I U1828 ( .A(fd_Inst[31]), .B(fd_Inst[30]), .Z(n1464) );
  AN2I U1829 ( .A(n1464), .B(n4753), .Z(n2019) );
  AN2I U1830 ( .A(n4863), .B(n4864), .Z(n4696) );
  NR2I U1831 ( .A(mw_Inst[30]), .B(mw_Inst[28]), .Z(n1529) );
  AN2I U1832 ( .A(n4696), .B(n1529), .Z(n4693) );
  AN2I U1833 ( .A(mw_Inst[26]), .B(mw_Inst[27]), .Z(n1514) );
  ND2I U1834 ( .A(n4693), .B(n1514), .Z(n1992) );
  NR2I U1835 ( .A(mw_Inst[31]), .B(mw_Inst[30]), .Z(n1466) );
  ND2I U1836 ( .A(n1515), .B(n1516), .Z(n1468) );
  MUX21LP U1837 ( .A(mw_Inst[15]), .B(mw_Inst[20]), .S(n1468), .Z(n2059) );
  ND2I U1838 ( .A(n1992), .B(n2059), .Z(n4874) );
  ENI U1839 ( .A(n4874), .B(fd_Inst[25]), .Z(n1473) );
  ND2I U1840 ( .A(n4693), .B(n1514), .Z(n2060) );
  ND2I U1841 ( .A(n1468), .B(mw_Inst[16]), .Z(n1467) );
  AN2I U1842 ( .A(n1992), .B(n1467), .Z(n1471) );
  IVI U1843 ( .A(n1468), .Z(n1469) );
  ND2I U1844 ( .A(n1469), .B(mw_Inst[11]), .Z(n1470) );
  ND2I U1845 ( .A(n1471), .B(n1470), .Z(n3762) );
  ENI U1846 ( .A(n3762), .B(fd_Inst[21]), .Z(n1472) );
  AN2I U1847 ( .A(n1473), .B(n1472), .Z(n1507) );
  NR2I U1848 ( .A(xm_Inst[30]), .B(xm_Inst[29]), .Z(n1474) );
  IVI U1849 ( .A(xm_Inst[28]), .Z(n4698) );
  AN2I U1850 ( .A(n1474), .B(n4698), .Z(n1485) );
  NR2I U1851 ( .A(xm_Inst[27]), .B(xm_Inst[26]), .Z(n1486) );
  ND2I U1852 ( .A(n1485), .B(n1486), .Z(n1498) );
  IVI U1853 ( .A(n1498), .Z(n1475) );
  ND2I U1854 ( .A(n4766), .B(n1475), .Z(n1481) );
  NR2I U1855 ( .A(xm_Inst[30]), .B(xm_Inst[29]), .Z(n1483) );
  ND2I U1856 ( .A(xm_Inst[27]), .B(xm_Inst[26]), .Z(n1476) );
  IVI U1857 ( .A(n1476), .Z(n1477) );
  ND2I U1858 ( .A(n4860), .B(n1477), .Z(n1478) );
  IVI U1859 ( .A(n1478), .Z(n1482) );
  ND2I U1860 ( .A(n1483), .B(n1482), .Z(n1493) );
  ND2I U1861 ( .A(n4763), .B(n1493), .Z(n1479) );
  IVI U1862 ( .A(n1479), .Z(n2004) );
  ND2I U1863 ( .A(n2004), .B(n1498), .Z(n1480) );
  ND2I U1864 ( .A(n1481), .B(n1480), .Z(n2326) );
  ENI U1865 ( .A(n2326), .B(fd_Inst[22]), .Z(n1488) );
  ND2I U1866 ( .A(n1483), .B(n1482), .Z(n1497) );
  AN2I U1867 ( .A(n1497), .B(n4768), .Z(n1484) );
  ND2I U1868 ( .A(n1485), .B(n1486), .Z(n2006) );
  ND2I U1869 ( .A(n1484), .B(n2006), .Z(n2023) );
  ND2I U1870 ( .A(n1486), .B(n1485), .Z(n1496) );
  IVI U1871 ( .A(n1496), .Z(n1491) );
  ND2I U1872 ( .A(n1491), .B(n4781), .Z(n2022) );
  ND2I U1873 ( .A(n1163), .B(n2022), .Z(n2325) );
  ENI U1874 ( .A(n2325), .B(fd_Inst[21]), .Z(n1487) );
  NR2I U1875 ( .A(n1488), .B(n1487), .Z(n1506) );
  ND2I U1876 ( .A(n4765), .B(n1493), .Z(n1489) );
  IVI U1877 ( .A(n1489), .Z(n1490) );
  ND2I U1878 ( .A(n1490), .B(n2006), .Z(n2034) );
  ND2I U1879 ( .A(n1491), .B(n4780), .Z(n2033) );
  ND2I U1880 ( .A(n2034), .B(n2033), .Z(n2323) );
  ENI U1881 ( .A(n2323), .B(n4717), .Z(n1492) );
  ND2I U1882 ( .A(n4755), .B(n1492), .Z(n1504) );
  ND2I U1883 ( .A(n4764), .B(n1493), .Z(n1494) );
  IVI U1884 ( .A(n1494), .Z(n1495) );
  ND2I U1885 ( .A(n1495), .B(n1498), .Z(n2031) );
  IVI U1886 ( .A(n1496), .Z(n1500) );
  ND2I U1887 ( .A(n1500), .B(n4778), .Z(n2030) );
  ND2I U1888 ( .A(n2031), .B(n2030), .Z(n2331) );
  ENI U1889 ( .A(n2331), .B(n4757), .Z(n1502) );
  AN2I U1890 ( .A(n1497), .B(n4767), .Z(n1499) );
  ND2I U1891 ( .A(n1499), .B(n1498), .Z(n2026) );
  ND2I U1892 ( .A(n1500), .B(n4779), .Z(n2025) );
  ND2I U1893 ( .A(n1162), .B(n2025), .Z(n2332) );
  ENI U1894 ( .A(n2332), .B(n4758), .Z(n1501) );
  ND2I U1895 ( .A(n1502), .B(n1501), .Z(n1503) );
  NR2I U1896 ( .A(n1504), .B(n1503), .Z(n1505) );
  ND2I U1897 ( .A(n1506), .B(n1505), .Z(n1531) );
  AN2I U1898 ( .A(n1507), .B(n1531), .Z(n1525) );
  ND2I U1899 ( .A(n1516), .B(n1515), .Z(n1508) );
  ND2I U1900 ( .A(n1457), .B(n1508), .Z(n1510) );
  IVI U1901 ( .A(n1508), .Z(n1519) );
  ND2I U1902 ( .A(n1519), .B(n1458), .Z(n1509) );
  ND2I U1903 ( .A(n1510), .B(n1509), .Z(n1511) );
  ND2I U1904 ( .A(n2060), .B(n1511), .Z(gpr_wr_addr[2]) );
  ENI U1905 ( .A(gpr_wr_addr[2]), .B(fd_Inst[23]), .Z(n1513) );
  B2I U1906 ( .A(mw_Inst[29]), .Z2(n1527) );
  ND2I U1907 ( .A(n1527), .B(n1526), .Z(n2342) );
  AN2I U1908 ( .A(n2342), .B(n1532), .Z(n1512) );
  ND2I U1909 ( .A(n1513), .B(n1512), .Z(n1523) );
  ND2I U1910 ( .A(n4693), .B(n1514), .Z(n2038) );
  ND2I U1911 ( .A(n1516), .B(n1515), .Z(n1517) );
  MUX21LP U1912 ( .A(mw_Inst[12]), .B(mw_Inst[17]), .S(n1517), .Z(n2037) );
  ND2I U1913 ( .A(n1992), .B(n2037), .Z(n4712) );
  ENI U1914 ( .A(n4712), .B(fd_Inst[22]), .Z(n1521) );
  ND2I U1915 ( .A(n1517), .B(mw_Inst[19]), .Z(n1518) );
  AN2I U1916 ( .A(n2038), .B(n1518), .Z(n2056) );
  ND2I U1917 ( .A(mw_Inst[14]), .B(n1519), .Z(n2053) );
  ND2I U1918 ( .A(n2056), .B(n2053), .Z(gpr_wr_addr[3]) );
  ENI U1919 ( .A(gpr_wr_addr[3]), .B(fd_Inst[24]), .Z(n1520) );
  ND2I U1920 ( .A(n1521), .B(n1520), .Z(n1522) );
  NR2I U1921 ( .A(n1523), .B(n1522), .Z(n1524) );
  ND2I U1922 ( .A(n1525), .B(n1524), .Z(n1534) );
  B4IP U1923 ( .A(n1534), .Z(n1866) );
  NR2I U1924 ( .A(n1527), .B(n1441), .Z(n1528) );
  AN2I U1925 ( .A(n1529), .B(n1528), .Z(n1530) );
  B2I U1926 ( .A(mw_Inst[27]), .Z2(n4692) );
  ENI U1927 ( .A(mw_Inst[26]), .B(n4692), .Z(n4694) );
  AN2I U1928 ( .A(n1530), .B(n4694), .Z(n1757) );
  B4IP U1929 ( .A(n1757), .Z(n1806) );
  MUX21L U1930 ( .A(n4807), .B(n4738), .S(n1806), .Z(n2500) );
  IVI U1931 ( .A(n1531), .Z(n1533) );
  AN2I U1932 ( .A(n1533), .B(n1532), .Z(n1617) );
  B2IP U1933 ( .A(n1617), .Z1(n1450), .Z2(n1865) );
  AO2 U1934 ( .A(n1866), .B(n2500), .C(n1865), .D(Addr[30]), .Z(n1536) );
  ND2I U1935 ( .A(n1450), .B(n1534), .Z(n1665) );
  IVI U1936 ( .A(n1665), .Z(n1573) );
  IVI U1937 ( .A(n1573), .Z(n1773) );
  IVI U1938 ( .A(n1773), .Z(n1810) );
  ND2I U1939 ( .A(n1810), .B(gpr_rd_data1[30]), .Z(n1535) );
  ND2I U1940 ( .A(n1536), .B(n1535), .Z(n1673) );
  IVDA U1941 ( .A(n2019), .Y(n1465), .Z(n1540) );
  IVI U1942 ( .A(fd_Inst[28]), .Z(n1538) );
  AO2 U1943 ( .A(n3829), .B(n1673), .C(n3740), .D(PC[30]), .Z(n1929) );
  AN2I U1944 ( .A(n1537), .B(n3418), .Z(n3824) );
  NR2I U1945 ( .A(fd_Inst[27]), .B(n1538), .Z(n1539) );
  AN2I U1946 ( .A(n1540), .B(n1539), .Z(n3544) );
  AN2I U1947 ( .A(fd_Inst[26]), .B(n3544), .Z(n1909) );
  IVI U1948 ( .A(gpr_rd_data2[4]), .Z(n4857) );
  IVI U1949 ( .A(n4861), .Z(n4862) );
  IVI U1950 ( .A(n4862), .Z(n3955) );
  ENI U1951 ( .A(n2326), .B(n3955), .Z(n1541) );
  ND2I U1952 ( .A(n4755), .B(n1541), .Z(n1545) );
  B2IP U1953 ( .A(fd_Inst[18]), .Z1(n1449), .Z2(n4714) );
  ENI U1954 ( .A(n2331), .B(n1449), .Z(n1543) );
  B2IP U1955 ( .A(fd_Inst[16]), .Z1(n1447), .Z2(n4713) );
  ENI U1956 ( .A(n2325), .B(n1447), .Z(n1542) );
  ND2I U1957 ( .A(n1543), .B(n1542), .Z(n1544) );
  NR2I U1958 ( .A(n1545), .B(n1544), .Z(n1549) );
  IVI U1959 ( .A(n4858), .Z(n4859) );
  ENI U1960 ( .A(n2332), .B(n4859), .Z(n1547) );
  ENI U1961 ( .A(n2323), .B(fd_Inst[20]), .Z(n1546) );
  NR2I U1962 ( .A(n1547), .B(n1546), .Z(n1548) );
  ND2I U1963 ( .A(n1549), .B(n1548), .Z(n1558) );
  IVI U1964 ( .A(n1558), .Z(n1553) );
  NR2I U1965 ( .A(n4714), .B(fd_Inst[20]), .Z(n1552) );
  NR2I U1966 ( .A(n4862), .B(n4713), .Z(n1550) );
  IVI U1967 ( .A(n4859), .Z(n3951) );
  AN2I U1968 ( .A(n1550), .B(n3951), .Z(n1551) );
  ND2I U1969 ( .A(n1552), .B(n1551), .Z(n1554) );
  ND2I U1970 ( .A(n1553), .B(n1554), .Z(n1574) );
  ENI U1971 ( .A(gpr_wr_addr[2]), .B(n4714), .Z(n1556) );
  AN2I U1972 ( .A(n2342), .B(n1554), .Z(n1555) );
  AN2I U1973 ( .A(n1556), .B(n1555), .Z(n1557) );
  AN2I U1974 ( .A(n1558), .B(n1557), .Z(n1566) );
  ENI U1975 ( .A(gpr_wr_addr[3]), .B(n4859), .Z(n1560) );
  ENI U1976 ( .A(n4712), .B(n4862), .Z(n1559) );
  ND2I U1977 ( .A(n1560), .B(n1559), .Z(n1564) );
  ENI U1978 ( .A(n3762), .B(n4713), .Z(n1562) );
  ENI U1979 ( .A(n4874), .B(fd_Inst[20]), .Z(n1561) );
  ND2I U1980 ( .A(n1562), .B(n1561), .Z(n1563) );
  NR2I U1981 ( .A(n1564), .B(n1563), .Z(n1565) );
  ND2I U1982 ( .A(n1566), .B(n1565), .Z(n1567) );
  ND2I U1983 ( .A(n1574), .B(n1567), .Z(n1760) );
  B4I U1984 ( .A(n1767), .Z(n1797) );
  B5IP U1985 ( .A(n1567), .Z(n1867) );
  MUX21LP U1986 ( .A(n4791), .B(n4727), .S(n1806), .Z(n4678) );
  ND2I U1987 ( .A(n1867), .B(n4678), .Z(n1569) );
  IVI U1988 ( .A(n1574), .Z(n1868) );
  ND2I U1989 ( .A(n1868), .B(Addr[4]), .Z(n1568) );
  AO3 U1990 ( .A(n4857), .B(n1797), .C(n1569), .D(n1568), .Z(n1572) );
  AO2 U1991 ( .A(n1866), .B(n4678), .C(n1865), .D(Addr[4]), .Z(n1571) );
  ND2I U1992 ( .A(n1810), .B(gpr_rd_data1[4]), .Z(n1570) );
  ND2I U1993 ( .A(n1571), .B(n1570), .Z(n3672) );
  ENI U1994 ( .A(n1572), .B(n3672), .Z(n1589) );
  IVI U1995 ( .A(n1573), .Z(n1735) );
  MUX21LP U1996 ( .A(n4785), .B(n4720), .S(n1806), .Z(n2534) );
  ND2I U1997 ( .A(n1867), .B(n2534), .Z(n1576) );
  IVI U1998 ( .A(n1574), .Z(n1740) );
  ND2I U1999 ( .A(n1740), .B(Addr[16]), .Z(n1575) );
  AN2I U2000 ( .A(n1576), .B(n1575), .Z(n1578) );
  IVI U2001 ( .A(n1760), .Z(n1767) );
  ND2I U2002 ( .A(n1767), .B(gpr_rd_data2[16]), .Z(n1577) );
  ND2I U2003 ( .A(n1578), .B(n1577), .Z(n1713) );
  NR2I U2004 ( .A(n1735), .B(n1713), .Z(n1579) );
  ND2I U2005 ( .A(gpr_rd_data1[16]), .B(n1579), .Z(n1587) );
  IVI U2006 ( .A(n1665), .Z(n1722) );
  ND2I U2007 ( .A(n1722), .B(gpr_rd_data1[10]), .Z(n3393) );
  ND2I U2008 ( .A(n1617), .B(Addr[10]), .Z(n1581) );
  MUX21LP U2009 ( .A(n4804), .B(n4736), .S(n1806), .Z(n4682) );
  ND2I U2010 ( .A(n1866), .B(n4682), .Z(n1580) );
  ND2I U2011 ( .A(n1581), .B(n1580), .Z(n1685) );
  IVI U2012 ( .A(n1685), .Z(n3394) );
  AO2 U2013 ( .A(n1867), .B(n4682), .C(n1868), .D(Addr[10]), .Z(n1583) );
  ND2I U2014 ( .A(n1767), .B(gpr_rd_data2[10]), .Z(n1582) );
  AN2I U2015 ( .A(n1583), .B(n1582), .Z(n1686) );
  IVI U2016 ( .A(n1686), .Z(n1584) );
  AN2I U2017 ( .A(n3394), .B(n1584), .Z(n1585) );
  ND2I U2018 ( .A(n3393), .B(n1585), .Z(n1586) );
  AN2I U2019 ( .A(n1587), .B(n1586), .Z(n1588) );
  ND2I U2020 ( .A(n1589), .B(n1588), .Z(n1590) );
  IVI U2021 ( .A(n1590), .Z(n1608) );
  ND2I U2022 ( .A(n1865), .B(Addr[14]), .Z(n1592) );
  MUX21LP U2023 ( .A(n4814), .B(n4745), .S(n1806), .Z(n4684) );
  ND2I U2024 ( .A(n1866), .B(n4684), .Z(n1591) );
  ND2I U2025 ( .A(n1592), .B(n1591), .Z(n1712) );
  IVI U2026 ( .A(n1712), .Z(n3459) );
  ND2I U2027 ( .A(n1867), .B(n4684), .Z(n1594) );
  ND2I U2028 ( .A(n1740), .B(Addr[14]), .Z(n1593) );
  AN2I U2029 ( .A(n1594), .B(n1593), .Z(n1709) );
  ND2I U2030 ( .A(n1767), .B(gpr_rd_data2[14]), .Z(n1708) );
  ND2I U2031 ( .A(n1709), .B(n1708), .Z(n1652) );
  AN2I U2032 ( .A(n3459), .B(n1652), .Z(n1595) );
  ND2I U2033 ( .A(n1596), .B(n1595), .Z(n1606) );
  ND2I U2034 ( .A(n1722), .B(gpr_rd_data1[8]), .Z(n3710) );
  ND2I U2035 ( .A(n1865), .B(Addr[8]), .Z(n1598) );
  IVI U2036 ( .A(n1757), .Z(n1632) );
  MUX21LP U2037 ( .A(n4805), .B(n4737), .S(n1632), .Z(n2396) );
  ND2I U2038 ( .A(n1866), .B(n2396), .Z(n1597) );
  ND2I U2039 ( .A(n1598), .B(n1597), .Z(n1687) );
  IVI U2040 ( .A(n1687), .Z(n3711) );
  ND2I U2041 ( .A(n3710), .B(n3711), .Z(n1602) );
  AO2 U2042 ( .A(n1867), .B(n2396), .C(n1868), .D(Addr[8]), .Z(n1600) );
  ND2I U2043 ( .A(n1767), .B(gpr_rd_data2[8]), .Z(n1599) );
  AN2I U2044 ( .A(n1600), .B(n1599), .Z(n1688) );
  IVI U2045 ( .A(n1688), .Z(n1601) );
  ND2I U2046 ( .A(n1602), .B(n1601), .Z(n1604) );
  ND2I U2047 ( .A(n1688), .B(n3710), .Z(n1603) );
  ND2I U2048 ( .A(n1604), .B(n1603), .Z(n1605) );
  AN2I U2049 ( .A(n1606), .B(n1605), .Z(n1607) );
  ND2I U2050 ( .A(n1608), .B(n1607), .Z(n1645) );
  ND2I U2051 ( .A(n1810), .B(gpr_rd_data1[12]), .Z(n1610) );
  MUX21LP U2052 ( .A(n4816), .B(n4747), .S(n1806), .Z(n2418) );
  AO2 U2053 ( .A(n1866), .B(n2418), .C(n1865), .D(Addr[12]), .Z(n1609) );
  ND2I U2054 ( .A(n1610), .B(n1609), .Z(n3489) );
  IVI U2055 ( .A(gpr_rd_data2[12]), .Z(n1613) );
  ND2I U2056 ( .A(n1867), .B(n2418), .Z(n1612) );
  ND2I U2057 ( .A(n1868), .B(Addr[12]), .Z(n1611) );
  AO3 U2058 ( .A(n1613), .B(n1797), .C(n1612), .D(n1611), .Z(n1614) );
  IVI U2059 ( .A(n1614), .Z(n1615) );
  ENI U2060 ( .A(n3489), .B(n1615), .Z(n1626) );
  IVI U2061 ( .A(n3393), .Z(n1616) );
  ND2I U2062 ( .A(n1616), .B(n1686), .Z(n1624) );
  MUX21LP U2063 ( .A(n4818), .B(n4749), .S(n1632), .Z(n2372) );
  B2I U2064 ( .A(n1617), .Z2(n1856) );
  AO2 U2065 ( .A(n1866), .B(n2372), .C(n1856), .D(Addr[2]), .Z(n1619) );
  ND2I U2066 ( .A(gpr_rd_data1[2]), .B(n1722), .Z(n1618) );
  ND2I U2067 ( .A(n1619), .B(n1618), .Z(n3661) );
  IVI U2068 ( .A(gpr_rd_data2[2]), .Z(n4856) );
  ND2I U2069 ( .A(n1867), .B(n2372), .Z(n1621) );
  ND2I U2070 ( .A(n1868), .B(Addr[2]), .Z(n1620) );
  AO3P U2071 ( .A(n4856), .B(n1797), .C(n1621), .D(n1620), .Z(n1622) );
  ENI U2072 ( .A(n3661), .B(n1622), .Z(n1623) );
  ND2I U2073 ( .A(n1624), .B(n1623), .Z(n1625) );
  NR2I U2074 ( .A(n1626), .B(n1625), .Z(n1643) );
  MUX21LP U2075 ( .A(n4806), .B(n4723), .S(n1632), .Z(n4680) );
  AO2 U2076 ( .A(n1866), .B(n4680), .C(n1865), .D(Addr[6]), .Z(n3689) );
  ND2I U2077 ( .A(gpr_rd_data1[6]), .B(n1722), .Z(n3688) );
  ND2I U2078 ( .A(n3689), .B(n3688), .Z(n1631) );
  IVI U2079 ( .A(gpr_rd_data2[6]), .Z(n1629) );
  ND2I U2080 ( .A(n1867), .B(n4680), .Z(n1628) );
  ND2I U2081 ( .A(n1740), .B(Addr[6]), .Z(n1627) );
  AO3 U2082 ( .A(n1629), .B(n1797), .C(n1628), .D(n1627), .Z(n1630) );
  ENI U2083 ( .A(n1631), .B(n1630), .Z(n1640) );
  MUX21LP U2084 ( .A(n4784), .B(n4719), .S(n1632), .Z(n4676) );
  AO2 U2085 ( .A(n1866), .B(n4676), .C(n1865), .D(Addr[0]), .Z(n1634) );
  ND2I U2086 ( .A(n1722), .B(gpr_rd_data1[0]), .Z(n1633) );
  ND2I U2087 ( .A(n1634), .B(n1633), .Z(n3825) );
  IVI U2088 ( .A(gpr_rd_data2[0]), .Z(n1637) );
  ND2I U2089 ( .A(n1867), .B(n4676), .Z(n1636) );
  ND2I U2090 ( .A(n1740), .B(Addr[0]), .Z(n1635) );
  AO3 U2091 ( .A(n1637), .B(n1797), .C(n1636), .D(n1635), .Z(n1638) );
  ENI U2092 ( .A(n3825), .B(n1638), .Z(n1639) );
  ND2I U2093 ( .A(n1640), .B(n1639), .Z(n1641) );
  IVI U2094 ( .A(n1641), .Z(n1642) );
  ND2I U2095 ( .A(n1643), .B(n1642), .Z(n1644) );
  NR2I U2096 ( .A(n1645), .B(n1644), .Z(n1755) );
  MUX21L U2097 ( .A(n4802), .B(n4734), .S(n1806), .Z(n2478) );
  AO2 U2098 ( .A(n1866), .B(n2478), .C(n1865), .D(Addr[26]), .Z(n1647) );
  ND2I U2099 ( .A(n1810), .B(gpr_rd_data1[26]), .Z(n1646) );
  ND2I U2100 ( .A(n1647), .B(n1646), .Z(n3481) );
  IVI U2101 ( .A(gpr_rd_data2[26]), .Z(n1650) );
  ND2I U2102 ( .A(n1867), .B(n2478), .Z(n1649) );
  ND2I U2103 ( .A(n1740), .B(Addr[26]), .Z(n1648) );
  AO3 U2104 ( .A(n1650), .B(n1797), .C(n1649), .D(n1648), .Z(n1651) );
  ENI U2105 ( .A(n3481), .B(n1651), .Z(n1655) );
  NR2I U2106 ( .A(n1665), .B(n1652), .Z(n1653) );
  ND2I U2107 ( .A(n1653), .B(gpr_rd_data1[14]), .Z(n1654) );
  ND2I U2108 ( .A(n1655), .B(n1654), .Z(n1656) );
  IVI U2109 ( .A(n1656), .Z(n1678) );
  IVI U2110 ( .A(gpr_rd_data1[16]), .Z(n1660) );
  ND2I U2111 ( .A(n1865), .B(Addr[16]), .Z(n1658) );
  ND2I U2112 ( .A(n1866), .B(n2534), .Z(n1657) );
  ND2I U2113 ( .A(n1658), .B(n1657), .Z(n1715) );
  IVI U2114 ( .A(n1715), .Z(n3516) );
  AN2I U2115 ( .A(n3516), .B(n1713), .Z(n1659) );
  ND2I U2116 ( .A(n1660), .B(n1659), .Z(n1668) );
  MUX21LP U2117 ( .A(n4812), .B(n4743), .S(n1806), .Z(n2459) );
  ND2I U2118 ( .A(n1867), .B(n2459), .Z(n1662) );
  ND2I U2119 ( .A(n1740), .B(Addr[20]), .Z(n1661) );
  AN2I U2120 ( .A(n1662), .B(n1661), .Z(n1664) );
  ND2I U2121 ( .A(n1767), .B(gpr_rd_data2[20]), .Z(n1663) );
  ND2I U2122 ( .A(n1664), .B(n1663), .Z(n1731) );
  NR2I U2123 ( .A(n1665), .B(n1731), .Z(n1666) );
  ND2I U2124 ( .A(n1666), .B(gpr_rd_data1[20]), .Z(n1667) );
  AN2I U2125 ( .A(n1668), .B(n1667), .Z(n1675) );
  IVI U2126 ( .A(gpr_rd_data2[30]), .Z(n1671) );
  ND2I U2127 ( .A(n1867), .B(n2500), .Z(n1670) );
  ND2I U2128 ( .A(n1740), .B(Addr[30]), .Z(n1669) );
  AO3P U2129 ( .A(n1671), .B(n1797), .C(n1670), .D(n1669), .Z(n1672) );
  ENI U2130 ( .A(n1673), .B(n1672), .Z(n1674) );
  ND2I U2131 ( .A(n1675), .B(n1674), .Z(n1676) );
  IVI U2132 ( .A(n1676), .Z(n1677) );
  ND2I U2133 ( .A(n1678), .B(n1677), .Z(n1753) );
  MUX21LP U2134 ( .A(n4799), .B(n4731), .S(n1806), .Z(n4688) );
  AO2 U2135 ( .A(n1866), .B(n4688), .C(n1865), .D(Addr[22]), .Z(n1680) );
  ND2I U2136 ( .A(n1810), .B(gpr_rd_data1[22]), .Z(n1679) );
  ND2I U2137 ( .A(n1680), .B(n1679), .Z(n3570) );
  IVI U2138 ( .A(gpr_rd_data2[22]), .Z(n1683) );
  ND2I U2139 ( .A(n1867), .B(n4688), .Z(n1682) );
  ND2I U2140 ( .A(n1740), .B(Addr[22]), .Z(n1681) );
  AO3 U2141 ( .A(n1683), .B(n1797), .C(n1682), .D(n1681), .Z(n1684) );
  ENI U2142 ( .A(n3570), .B(n1684), .Z(n1700) );
  AO2P U2143 ( .A(n1688), .B(n1687), .C(n1686), .D(n1685), .Z(n1698) );
  ND2I U2144 ( .A(n1865), .B(Addr[24]), .Z(n1690) );
  MUX21LP U2145 ( .A(n4810), .B(n4741), .S(n1806), .Z(n2473) );
  ND2I U2146 ( .A(n1866), .B(n2473), .Z(n1689) );
  ND2I U2147 ( .A(n1690), .B(n1689), .Z(n1719) );
  IVI U2148 ( .A(n1719), .Z(n3583) );
  ND2I U2149 ( .A(n1867), .B(n2473), .Z(n1692) );
  ND2I U2150 ( .A(n1740), .B(Addr[24]), .Z(n1691) );
  AN2I U2151 ( .A(n1692), .B(n1691), .Z(n1694) );
  ND2I U2152 ( .A(n1767), .B(gpr_rd_data2[24]), .Z(n1693) );
  ND2I U2153 ( .A(n1694), .B(n1693), .Z(n1734) );
  AN2I U2154 ( .A(n3583), .B(n1734), .Z(n1696) );
  IVI U2155 ( .A(gpr_rd_data1[24]), .Z(n1695) );
  ND2I U2156 ( .A(n1696), .B(n1695), .Z(n1697) );
  AN2I U2157 ( .A(n1698), .B(n1697), .Z(n1699) );
  ND2I U2158 ( .A(n1700), .B(n1699), .Z(n1701) );
  IVI U2159 ( .A(n1701), .Z(n1751) );
  MUX21LP U2160 ( .A(n4787), .B(n4722), .S(n1806), .Z(n4690) );
  AO2 U2161 ( .A(n1866), .B(n4690), .C(n1865), .D(Addr[28]), .Z(n1703) );
  ND2I U2162 ( .A(n1810), .B(gpr_rd_data1[28]), .Z(n1702) );
  ND2I U2163 ( .A(n1703), .B(n1702), .Z(n3629) );
  IVI U2164 ( .A(gpr_rd_data2[28]), .Z(n1706) );
  ND2I U2165 ( .A(n1867), .B(n4690), .Z(n1705) );
  ND2I U2166 ( .A(n1740), .B(Addr[28]), .Z(n1704) );
  AO3P U2167 ( .A(n1706), .B(n1797), .C(n1705), .D(n1704), .Z(n1707) );
  ENI U2168 ( .A(n3629), .B(n1707), .Z(n1729) );
  NR2I U2169 ( .A(n1722), .B(n1712), .Z(n1711) );
  ND2I U2170 ( .A(n1709), .B(n1708), .Z(n1710) );
  MUX21L U2171 ( .A(n1712), .B(n1711), .S(n1710), .Z(n1717) );
  NR2I U2172 ( .A(n1722), .B(n1715), .Z(n1714) );
  MUX21L U2173 ( .A(n1715), .B(n1714), .S(n1713), .Z(n1716) );
  AN2I U2174 ( .A(n1717), .B(n1716), .Z(n1727) );
  NR2I U2175 ( .A(n1722), .B(n1719), .Z(n1718) );
  MUX21L U2176 ( .A(n1719), .B(n1718), .S(n1734), .Z(n1725) );
  ND2I U2177 ( .A(n1865), .B(Addr[20]), .Z(n1721) );
  ND2I U2178 ( .A(n1866), .B(n2459), .Z(n1720) );
  ND2I U2179 ( .A(n1721), .B(n1720), .Z(n1730) );
  NR2I U2180 ( .A(n1722), .B(n1730), .Z(n1723) );
  MUX21L U2181 ( .A(n1730), .B(n1723), .S(n1731), .Z(n1724) );
  AN2I U2182 ( .A(n1725), .B(n1724), .Z(n1726) );
  AN2I U2183 ( .A(n1727), .B(n1726), .Z(n1728) );
  ND2I U2184 ( .A(n1729), .B(n1728), .Z(n1749) );
  IVI U2185 ( .A(gpr_rd_data1[20]), .Z(n1733) );
  IVI U2186 ( .A(n1730), .Z(n3435) );
  AN2I U2187 ( .A(n3435), .B(n1731), .Z(n1732) );
  ND2I U2188 ( .A(n1733), .B(n1732), .Z(n1738) );
  NR2I U2189 ( .A(n1735), .B(n1734), .Z(n1736) );
  ND2I U2190 ( .A(n1736), .B(gpr_rd_data1[24]), .Z(n1737) );
  ND2I U2191 ( .A(n1738), .B(n1737), .Z(n1739) );
  IVI U2192 ( .A(n1739), .Z(n1747) );
  MUX21LP U2193 ( .A(n4786), .B(n4721), .S(n1806), .Z(n4686) );
  AO2 U2194 ( .A(n1866), .B(n4686), .C(n1865), .D(Addr[18]), .Z(n3534) );
  ND2I U2195 ( .A(n1810), .B(n1433), .Z(n3533) );
  ND2I U2196 ( .A(n3534), .B(n3533), .Z(n1745) );
  IVI U2197 ( .A(gpr_rd_data2[18]), .Z(n1743) );
  ND2I U2198 ( .A(n1867), .B(n4686), .Z(n1742) );
  ND2I U2199 ( .A(n1740), .B(Addr[18]), .Z(n1741) );
  AO3 U2200 ( .A(n1743), .B(n1797), .C(n1742), .D(n1741), .Z(n1744) );
  ENI U2201 ( .A(n1745), .B(n1744), .Z(n1746) );
  ND2I U2202 ( .A(n1747), .B(n1746), .Z(n1748) );
  NR2I U2203 ( .A(n1749), .B(n1748), .Z(n1750) );
  ND2I U2204 ( .A(n1751), .B(n1750), .Z(n1752) );
  NR2I U2205 ( .A(n1753), .B(n1752), .Z(n1754) );
  ND2I U2206 ( .A(n1755), .B(n1754), .Z(n1883) );
  ND2I U2207 ( .A(n1909), .B(n1883), .Z(n1756) );
  AN2I U2208 ( .A(n3824), .B(n1756), .Z(n3403) );
  B4IP U2209 ( .A(n1757), .Z(n1864) );
  MUX21LP U2210 ( .A(n4789), .B(n4725), .S(n1864), .Z(n4681) );
  AO2 U2211 ( .A(n1866), .B(n4681), .C(n1856), .D(Addr[7]), .Z(n1759) );
  IVI U2212 ( .A(n1773), .Z(n3581) );
  ND2I U2213 ( .A(n3581), .B(gpr_rd_data1[7]), .Z(n1758) );
  ND2I U2214 ( .A(n1759), .B(n1758), .Z(n3698) );
  IVI U2215 ( .A(gpr_rd_data2[7]), .Z(n1763) );
  B2IP U2216 ( .A(n1760), .Z2(n1871) );
  ND2I U2217 ( .A(n1867), .B(n4681), .Z(n1762) );
  ND2I U2218 ( .A(n1868), .B(Addr[7]), .Z(n1761) );
  AO3 U2219 ( .A(n1763), .B(n1871), .C(n1762), .D(n1761), .Z(n1764) );
  ENI U2220 ( .A(n3698), .B(n1764), .Z(n1772) );
  MUX21LP U2221 ( .A(n4792), .B(n4728), .S(n1864), .Z(n4677) );
  AO2 U2222 ( .A(n1866), .B(n4677), .C(n1856), .D(Addr[1]), .Z(n1766) );
  ND2I U2223 ( .A(n3581), .B(gpr_rd_data1[1]), .Z(n1765) );
  ND2I U2224 ( .A(n1766), .B(n1765), .Z(n3828) );
  AO2 U2225 ( .A(n4677), .B(n1867), .C(Addr[1]), .D(n1868), .Z(n1769) );
  ND2I U2226 ( .A(n1767), .B(gpr_rd_data2[1]), .Z(n1768) );
  ND2I U2227 ( .A(n1769), .B(n1768), .Z(n1770) );
  ENI U2228 ( .A(n3828), .B(n1770), .Z(n1771) );
  ND2I U2229 ( .A(n1772), .B(n1771), .Z(n1886) );
  MUX21LP U2230 ( .A(n4817), .B(n4748), .S(n1864), .Z(n4683) );
  AO2 U2231 ( .A(n1866), .B(n4683), .C(n1856), .D(Addr[11]), .Z(n1775) );
  IVI U2232 ( .A(n1773), .Z(n3415) );
  ND2I U2233 ( .A(n3415), .B(gpr_rd_data1[11]), .Z(n1774) );
  ND2I U2234 ( .A(n1775), .B(n1774), .Z(n3404) );
  IVI U2235 ( .A(gpr_rd_data2[11]), .Z(n1778) );
  ND2I U2236 ( .A(n1867), .B(n4683), .Z(n1777) );
  ND2I U2237 ( .A(n1868), .B(Addr[11]), .Z(n1776) );
  AO3 U2238 ( .A(n1778), .B(n1871), .C(n1777), .D(n1776), .Z(n1779) );
  ENI U2239 ( .A(n3404), .B(n1779), .Z(n1786) );
  MUX21LP U2240 ( .A(n4803), .B(n4735), .S(n1864), .Z(n2401) );
  AO2 U2241 ( .A(n1866), .B(n2401), .C(n1856), .D(Addr[9]), .Z(n3726) );
  ND2I U2242 ( .A(n3415), .B(gpr_rd_data1[9]), .Z(n3725) );
  ND2I U2243 ( .A(n3726), .B(n3725), .Z(n1784) );
  IVI U2244 ( .A(gpr_rd_data2[9]), .Z(n1782) );
  ND2I U2245 ( .A(n1867), .B(n2401), .Z(n1781) );
  ND2I U2246 ( .A(n1868), .B(Addr[9]), .Z(n1780) );
  AO3 U2247 ( .A(n1782), .B(n1871), .C(n1781), .D(n1780), .Z(n1783) );
  ENI U2248 ( .A(n1784), .B(n1783), .Z(n1785) );
  ND2I U2249 ( .A(n1786), .B(n1785), .Z(n1885) );
  NR2I U2250 ( .A(n1886), .B(n1885), .Z(n1817) );
  IVI U2251 ( .A(gpr_rd_data2[23]), .Z(n1789) );
  MUX21L U2252 ( .A(n4809), .B(n4740), .S(n1864), .Z(n2464) );
  ND2I U2253 ( .A(n1867), .B(n2464), .Z(n1788) );
  ND2I U2254 ( .A(n1868), .B(Addr[23]), .Z(n1787) );
  AO3 U2255 ( .A(n1789), .B(n1871), .C(n1788), .D(n1787), .Z(n1792) );
  AO2 U2256 ( .A(n1866), .B(n2464), .C(n1856), .D(Addr[23]), .Z(n1791) );
  ND2I U2257 ( .A(n3415), .B(gpr_rd_data1[23]), .Z(n1790) );
  ND2I U2258 ( .A(n1791), .B(n1790), .Z(n3468) );
  ENI U2259 ( .A(n1792), .B(n3468), .Z(n1896) );
  MUX21LP U2260 ( .A(n4800), .B(n4732), .S(n1806), .Z(n4689) );
  AO2 U2261 ( .A(n1866), .B(n4689), .C(n1865), .D(Addr[25]), .Z(n1794) );
  ND2I U2262 ( .A(n1810), .B(gpr_rd_data1[25]), .Z(n1793) );
  ND2I U2263 ( .A(n1794), .B(n1793), .Z(n3598) );
  IVI U2264 ( .A(gpr_rd_data2[25]), .Z(n1798) );
  ND2I U2265 ( .A(n4689), .B(n1867), .Z(n1796) );
  ND2I U2266 ( .A(Addr[25]), .B(n1868), .Z(n1795) );
  AO3 U2267 ( .A(n1798), .B(n1797), .C(n1796), .D(n1795), .Z(n1799) );
  ENI U2268 ( .A(n3598), .B(n1799), .Z(n1902) );
  ND2I U2269 ( .A(n1896), .B(n1902), .Z(n1815) );
  ND2I U2270 ( .A(n3415), .B(gpr_rd_data1[13]), .Z(n1801) );
  MUX21LP U2271 ( .A(n4815), .B(n4746), .S(n1864), .Z(n2415) );
  AO2 U2272 ( .A(n1866), .B(n2415), .C(n1856), .D(Addr[13]), .Z(n1800) );
  ND2I U2273 ( .A(n1801), .B(n1800), .Z(n3444) );
  IVI U2274 ( .A(gpr_rd_data2[13]), .Z(n1804) );
  ND2I U2275 ( .A(n1867), .B(n2415), .Z(n1803) );
  ND2I U2276 ( .A(n1868), .B(Addr[13]), .Z(n1802) );
  AO3 U2277 ( .A(n1804), .B(n1871), .C(n1803), .D(n1802), .Z(n1805) );
  ENI U2278 ( .A(n3444), .B(n1805), .Z(n1901) );
  IVI U2279 ( .A(gpr_rd_data2[27]), .Z(n1809) );
  MUX21L U2280 ( .A(n4808), .B(n4739), .S(n1806), .Z(n2499) );
  ND2I U2281 ( .A(n1867), .B(n2499), .Z(n1808) );
  ND2I U2282 ( .A(n1868), .B(Addr[27]), .Z(n1807) );
  AO3 U2283 ( .A(n1809), .B(n1871), .C(n1808), .D(n1807), .Z(n1813) );
  AO2 U2284 ( .A(n1866), .B(n2499), .C(n1865), .D(Addr[27]), .Z(n1812) );
  ND2I U2285 ( .A(n1810), .B(gpr_rd_data1[27]), .Z(n1811) );
  ND2I U2286 ( .A(n1812), .B(n1811), .Z(n3617) );
  ENI U2287 ( .A(n1813), .B(n3617), .Z(n1904) );
  ND2I U2288 ( .A(n1901), .B(n1904), .Z(n1814) );
  NR2I U2289 ( .A(n1815), .B(n1814), .Z(n1816) );
  ND2I U2290 ( .A(n1817), .B(n1816), .Z(n1882) );
  MUX21LP U2291 ( .A(n4793), .B(n4729), .S(n1864), .Z(n2355) );
  AO2 U2292 ( .A(n1866), .B(n2355), .C(n1856), .D(Addr[3]), .Z(n1819) );
  ND2I U2293 ( .A(n3581), .B(gpr_rd_data1[3]), .Z(n1818) );
  ND2I U2294 ( .A(n1819), .B(n1818), .Z(n3667) );
  IVI U2295 ( .A(gpr_rd_data2[3]), .Z(n1822) );
  ND2I U2296 ( .A(n1867), .B(n2355), .Z(n1821) );
  ND2I U2297 ( .A(n1868), .B(Addr[3]), .Z(n1820) );
  AO3 U2298 ( .A(n1822), .B(n1871), .C(n1821), .D(n1820), .Z(n1823) );
  ENI U2299 ( .A(n3667), .B(n1823), .Z(n1895) );
  IVI U2300 ( .A(gpr_rd_data2[21]), .Z(n1826) );
  MUX21L U2301 ( .A(n4811), .B(n4742), .S(n1864), .Z(n4687) );
  ND2I U2302 ( .A(n1867), .B(n4687), .Z(n1825) );
  ND2I U2303 ( .A(n1868), .B(Addr[21]), .Z(n1824) );
  AO3 U2304 ( .A(n1826), .B(n1871), .C(n1825), .D(n1824), .Z(n1829) );
  AO2 U2305 ( .A(n1866), .B(n4687), .C(n1856), .D(Addr[21]), .Z(n1828) );
  ND2I U2306 ( .A(n3415), .B(gpr_rd_data1[21]), .Z(n1827) );
  ND2I U2307 ( .A(n1828), .B(n1827), .Z(n3555) );
  ENI U2308 ( .A(n1829), .B(n3555), .Z(n1898) );
  ND2I U2309 ( .A(n1895), .B(n1898), .Z(n1843) );
  MUX21LP U2310 ( .A(n4788), .B(n4724), .S(n1864), .Z(n4679) );
  AO2 U2311 ( .A(n1866), .B(n4679), .C(n1856), .D(Addr[5]), .Z(n1831) );
  ND2I U2312 ( .A(n3415), .B(gpr_rd_data1[5]), .Z(n1830) );
  ND2I U2313 ( .A(n1831), .B(n1830), .Z(n3680) );
  IVI U2314 ( .A(gpr_rd_data2[5]), .Z(n1834) );
  ND2I U2315 ( .A(n1867), .B(n4679), .Z(n1833) );
  ND2I U2316 ( .A(n1868), .B(Addr[5]), .Z(n1832) );
  AO3 U2317 ( .A(n1834), .B(n1871), .C(n1833), .D(n1832), .Z(n1835) );
  ENI U2318 ( .A(n3680), .B(n1835), .Z(n1897) );
  IVI U2319 ( .A(gpr_rd_data2[15]), .Z(n1838) );
  MUX21LP U2320 ( .A(n4790), .B(n4726), .S(n1864), .Z(n2424) );
  ND2I U2321 ( .A(n1867), .B(n2424), .Z(n1837) );
  ND2I U2322 ( .A(n1868), .B(Addr[15]), .Z(n1836) );
  AO3 U2323 ( .A(n1838), .B(n1871), .C(n1837), .D(n1836), .Z(n1841) );
  AO2 U2324 ( .A(n1866), .B(n2424), .C(n1856), .D(Addr[15]), .Z(n1840) );
  ND2I U2325 ( .A(n3415), .B(gpr_rd_data1[15]), .Z(n1839) );
  ND2I U2326 ( .A(n1840), .B(n1839), .Z(n3500) );
  ENI U2327 ( .A(n1841), .B(n3500), .Z(n1903) );
  ND2I U2328 ( .A(n1897), .B(n1903), .Z(n1842) );
  NR2I U2329 ( .A(n1843), .B(n1842), .Z(n1880) );
  MUX21L U2330 ( .A(n4813), .B(n4744), .S(n1864), .Z(n4685) );
  AO2 U2331 ( .A(n1866), .B(n4685), .C(n1856), .D(Addr[17]), .Z(n3417) );
  ND2I U2332 ( .A(n3415), .B(gpr_rd_data1[17]), .Z(n1844) );
  ND2I U2333 ( .A(n3417), .B(n1844), .Z(n1849) );
  IVI U2334 ( .A(gpr_rd_data2[17]), .Z(n1847) );
  ND2I U2335 ( .A(n1867), .B(n4685), .Z(n1846) );
  ND2I U2336 ( .A(n1868), .B(Addr[17]), .Z(n1845) );
  AO3 U2337 ( .A(n1847), .B(n1871), .C(n1846), .D(n1845), .Z(n1848) );
  ENI U2338 ( .A(n1849), .B(n1848), .Z(n1888) );
  IVI U2339 ( .A(gpr_rd_data2[29]), .Z(n1852) );
  MUX21LP U2340 ( .A(n4783), .B(n4718), .S(n1864), .Z(n4691) );
  ND2I U2341 ( .A(n1867), .B(n4691), .Z(n1851) );
  ND2I U2342 ( .A(n1868), .B(Addr[29]), .Z(n1850) );
  AO3 U2343 ( .A(n1852), .B(n1871), .C(n1851), .D(n1850), .Z(n1855) );
  AO2 U2344 ( .A(n1866), .B(n4691), .C(n1856), .D(Addr[29]), .Z(n1854) );
  ND2I U2345 ( .A(n3581), .B(gpr_rd_data1[29]), .Z(n1853) );
  ND2I U2346 ( .A(n1854), .B(n1853), .Z(n3741) );
  ENI U2347 ( .A(n1855), .B(n3741), .Z(n1890) );
  ND2I U2348 ( .A(n1888), .B(n1890), .Z(n1878) );
  MUX21L U2349 ( .A(n4798), .B(n4730), .S(n1864), .Z(n2450) );
  AO2 U2350 ( .A(n1866), .B(n2450), .C(n1856), .D(Addr[19]), .Z(n1858) );
  ND2I U2351 ( .A(gpr_rd_data1[19]), .B(n3415), .Z(n1857) );
  ND2I U2352 ( .A(n1858), .B(n1857), .Z(n3542) );
  IVI U2353 ( .A(gpr_rd_data2[19]), .Z(n1861) );
  ND2I U2354 ( .A(n1867), .B(n2450), .Z(n1860) );
  ND2I U2355 ( .A(n1868), .B(Addr[19]), .Z(n1859) );
  AO3 U2356 ( .A(n1861), .B(n1871), .C(n1860), .D(n1859), .Z(n1862) );
  ENI U2357 ( .A(n3542), .B(n1862), .Z(n1889) );
  IVI U2358 ( .A(n3544), .Z(n1863) );
  NR2I U2359 ( .A(fd_Inst[26]), .B(n1863), .Z(n1875) );
  MUX21L U2360 ( .A(n4801), .B(n4733), .S(n1864), .Z(n2504) );
  AO2 U2361 ( .A(n1866), .B(n2504), .C(n1865), .D(Addr[31]), .Z(n3646) );
  ND2I U2362 ( .A(n3581), .B(n1435), .Z(n3645) );
  ND2I U2363 ( .A(n3646), .B(n3645), .Z(n1874) );
  IVI U2364 ( .A(gpr_rd_data2[31]), .Z(n1872) );
  ND2I U2365 ( .A(n1867), .B(n2504), .Z(n1870) );
  ND2I U2366 ( .A(n1868), .B(Addr[31]), .Z(n1869) );
  AO3P U2367 ( .A(n1872), .B(n1871), .C(n1870), .D(n1869), .Z(n1873) );
  ENI U2368 ( .A(n1874), .B(n1873), .Z(n1887) );
  AN2I U2369 ( .A(n1875), .B(n1887), .Z(n1876) );
  ND2I U2370 ( .A(n1889), .B(n1876), .Z(n1877) );
  NR2I U2371 ( .A(n1878), .B(n1877), .Z(n1879) );
  ND2I U2372 ( .A(n1880), .B(n1879), .Z(n1881) );
  NR2I U2373 ( .A(n1882), .B(n1881), .Z(n1884) );
  IVI U2374 ( .A(n1883), .Z(n1987) );
  ND2I U2375 ( .A(n1884), .B(n1987), .Z(n1912) );
  NR2I U2376 ( .A(n1886), .B(n1885), .Z(n1894) );
  ND2I U2377 ( .A(n1888), .B(n1887), .Z(n1892) );
  ND2I U2378 ( .A(n1890), .B(n1889), .Z(n1891) );
  NR2I U2379 ( .A(n1892), .B(n1891), .Z(n1893) );
  AN2I U2380 ( .A(n1894), .B(n1893), .Z(n1985) );
  ND2I U2381 ( .A(n1896), .B(n1895), .Z(n1900) );
  ND2I U2382 ( .A(n1898), .B(n1897), .Z(n1899) );
  NR2I U2383 ( .A(n1900), .B(n1899), .Z(n1908) );
  ND2I U2384 ( .A(n1902), .B(n1901), .Z(n1906) );
  ND2I U2385 ( .A(n1904), .B(n1903), .Z(n1905) );
  NR2I U2386 ( .A(n1906), .B(n1905), .Z(n1907) );
  AN2I U2387 ( .A(n1908), .B(n1907), .Z(n1984) );
  ND2I U2388 ( .A(n1985), .B(n1984), .Z(n1910) );
  ND2I U2389 ( .A(n1910), .B(n1909), .Z(n1911) );
  ND2I U2390 ( .A(n1912), .B(n1911), .Z(n1913) );
  IVI U2391 ( .A(n1913), .Z(n3402) );
  ND2I U2392 ( .A(n3403), .B(n3402), .Z(n3974) );
  IVI U2393 ( .A(n3974), .Z(n3831) );
  ND2I U2394 ( .A(PC[28]), .B(PC[29]), .Z(n1914) );
  ND2I U2395 ( .A(PC[26]), .B(PC[27]), .Z(n3737) );
  NR2I U2396 ( .A(n1914), .B(n3737), .Z(n3641) );
  ENI U2397 ( .A(n3641), .B(n4827), .Z(n1918) );
  ND2I U2398 ( .A(PC[18]), .B(PC[19]), .Z(n3554) );
  ND2I U2399 ( .A(PC[20]), .B(PC[21]), .Z(n1915) );
  NR2I U2400 ( .A(n3554), .B(n1915), .Z(n3597) );
  ND2I U2401 ( .A(PC[22]), .B(PC[23]), .Z(n3596) );
  ND2I U2402 ( .A(PC[24]), .B(PC[25]), .Z(n1916) );
  NR2I U2403 ( .A(n3596), .B(n1916), .Z(n1917) );
  ND2I U2404 ( .A(n3597), .B(n1917), .Z(n3738) );
  MUX21L U2405 ( .A(n1918), .B(PC[30]), .S(n3738), .Z(n1927) );
  ND2I U2406 ( .A(PC[10]), .B(PC[11]), .Z(n3487) );
  ND2I U2407 ( .A(PC[12]), .B(PC[13]), .Z(n1919) );
  NR2I U2408 ( .A(n3487), .B(n1919), .Z(n3456) );
  ND2I U2409 ( .A(PC[14]), .B(PC[15]), .Z(n3512) );
  ND2I U2410 ( .A(PC[16]), .B(PC[17]), .Z(n1920) );
  NR2I U2411 ( .A(n3512), .B(n1920), .Z(n1921) );
  ND2I U2412 ( .A(n3456), .B(n1921), .Z(n1925) );
  ND2I U2413 ( .A(PC[6]), .B(PC[7]), .Z(n3723) );
  ND2I U2414 ( .A(PC[8]), .B(PC[9]), .Z(n1922) );
  NR2I U2415 ( .A(n3723), .B(n1922), .Z(n1924) );
  ND2I U2416 ( .A(PC[4]), .B(PC[5]), .Z(n1923) );
  ND2I U2417 ( .A(PC[3]), .B(PC[2]), .Z(n3679) );
  NR2I U2418 ( .A(n1923), .B(n3679), .Z(n3724) );
  ND2I U2419 ( .A(n1924), .B(n3724), .Z(n3414) );
  NR2I U2420 ( .A(n1925), .B(n3414), .Z(n1926) );
  B2IP U2421 ( .A(n1926), .Z2(n3739) );
  MUX21L U2422 ( .A(n4827), .B(n1927), .S(n3739), .Z(\pc_u0/pc_plus_4 [30]) );
  ND2I U2423 ( .A(n3666), .B(\pc_u0/pc_plus_4 [30]), .Z(n1928) );
  ND2I U2424 ( .A(n1929), .B(n1928), .Z(n1930) );
  IVI U2425 ( .A(n1930), .Z(n1991) );
  IVI U2426 ( .A(fd_Inst[15]), .Z(n1938) );
  IVI U2427 ( .A(n1938), .Z(n3630) );
  ND2I U2428 ( .A(n3630), .B(PC[28]), .Z(n3743) );
  IVI U2429 ( .A(n1938), .Z(n3742) );
  ND2I U2430 ( .A(n3742), .B(PC[29]), .Z(n1931) );
  ND2I U2431 ( .A(n3743), .B(n1931), .Z(n1933) );
  ND2I U2432 ( .A(n3630), .B(PC[26]), .Z(n3618) );
  ND2I U2433 ( .A(n3630), .B(PC[27]), .Z(n1932) );
  ND2I U2434 ( .A(n3618), .B(n1932), .Z(n3746) );
  NR2I U2435 ( .A(n1933), .B(n3746), .Z(n3649) );
  ENI U2436 ( .A(n3742), .B(PC[30]), .Z(n1937) );
  EOI U2437 ( .A(n3649), .B(n1937), .Z(n1951) );
  NR2I U2438 ( .A(n3630), .B(PC[27]), .Z(n1934) );
  NR2I U2439 ( .A(n3630), .B(PC[26]), .Z(n3620) );
  NR2I U2440 ( .A(n1934), .B(n3620), .Z(n3747) );
  NR2I U2441 ( .A(n3742), .B(PC[29]), .Z(n1935) );
  NR2I U2442 ( .A(n3630), .B(PC[28]), .Z(n3745) );
  NR2I U2443 ( .A(n1935), .B(n3745), .Z(n1936) );
  ND2I U2444 ( .A(n3747), .B(n1936), .Z(n3650) );
  EOI U2445 ( .A(n3650), .B(n1937), .Z(n1950) );
  IVI U2446 ( .A(n1938), .Z(n3599) );
  NR2I U2447 ( .A(n3599), .B(PC[23]), .Z(n1939) );
  IVI U2448 ( .A(n4715), .Z(n3571) );
  NR2I U2449 ( .A(n3571), .B(PC[22]), .Z(n3471) );
  NR2I U2450 ( .A(n1939), .B(n3471), .Z(n3603) );
  NR2I U2451 ( .A(n3599), .B(PC[25]), .Z(n1940) );
  NR2I U2452 ( .A(n3599), .B(PC[24]), .Z(n3602) );
  NR2I U2453 ( .A(n1940), .B(n3602), .Z(n1941) );
  ND2I U2454 ( .A(n3603), .B(n1941), .Z(n1945) );
  NR2I U2455 ( .A(n3571), .B(PC[19]), .Z(n1942) );
  NR2I U2456 ( .A(n3571), .B(PC[18]), .Z(n3545) );
  NR2I U2457 ( .A(n1942), .B(n3545), .Z(n3559) );
  NR2I U2458 ( .A(n3571), .B(PC[21]), .Z(n1943) );
  NR2I U2459 ( .A(n3571), .B(PC[20]), .Z(n3558) );
  NR2I U2460 ( .A(n1943), .B(n3558), .Z(n1944) );
  ND2I U2461 ( .A(n3559), .B(n1944), .Z(n3607) );
  NR2I U2462 ( .A(n1945), .B(n3607), .Z(n3750) );
  MUX21L U2463 ( .A(n1951), .B(n1950), .S(n3750), .Z(n1983) );
  ND2I U2464 ( .A(n3571), .B(PC[20]), .Z(n3556) );
  ND2I U2465 ( .A(n3571), .B(PC[21]), .Z(n1946) );
  ND2I U2466 ( .A(n3556), .B(n1946), .Z(n1948) );
  ND2I U2467 ( .A(n3742), .B(PC[18]), .Z(n3546) );
  ND2I U2468 ( .A(n3630), .B(PC[19]), .Z(n1947) );
  ND2I U2469 ( .A(n3546), .B(n1947), .Z(n3560) );
  NR2I U2470 ( .A(n1948), .B(n3560), .Z(n3608) );
  ND2I U2471 ( .A(n3599), .B(PC[24]), .Z(n3600) );
  ND2I U2472 ( .A(n3571), .B(PC[22]), .Z(n3469) );
  ND2I U2473 ( .A(n3599), .B(PC[23]), .Z(n1949) );
  ND2I U2474 ( .A(n3469), .B(n1949), .Z(n3604) );
  MUX21L U2475 ( .A(n1951), .B(n1950), .S(n3751), .Z(n1982) );
  NR2I U2476 ( .A(n3630), .B(PC[17]), .Z(n1953) );
  ND2I U2477 ( .A(n3742), .B(PC[17]), .Z(n1952) );
  ND2I U2478 ( .A(PC[16]), .B(fd_Inst[14]), .Z(n3420) );
  MUX21L U2479 ( .A(n1953), .B(n1952), .S(n3420), .Z(n1957) );
  NR2I U2480 ( .A(PC[16]), .B(fd_Inst[14]), .Z(n3421) );
  MUX21L U2481 ( .A(n1953), .B(n1952), .S(n3421), .Z(n1956) );
  NR2I U2482 ( .A(PC[15]), .B(fd_Inst[13]), .Z(n1955) );
  ND2I U2483 ( .A(PC[15]), .B(fd_Inst[13]), .Z(n1954) );
  NR2I U2484 ( .A(PC[14]), .B(fd_Inst[12]), .Z(n3503) );
  MUX21L U2485 ( .A(n1955), .B(n1954), .S(n3503), .Z(n3520) );
  MUX21L U2486 ( .A(n1957), .B(n1956), .S(n3520), .Z(n1965) );
  ND2I U2487 ( .A(PC[14]), .B(fd_Inst[12]), .Z(n3501) );
  MUX21L U2488 ( .A(n1955), .B(n1954), .S(n3501), .Z(n3519) );
  MUX21L U2489 ( .A(n1957), .B(n1956), .S(n3519), .Z(n1964) );
  NR2I U2490 ( .A(PC[13]), .B(fd_Inst[11]), .Z(n1959) );
  ND2I U2491 ( .A(PC[13]), .B(fd_Inst[11]), .Z(n1958) );
  ND2I U2492 ( .A(PC[12]), .B(fd_Inst[10]), .Z(n3445) );
  MUX21L U2493 ( .A(n1959), .B(n1958), .S(n3445), .Z(n1963) );
  NR2I U2494 ( .A(PC[12]), .B(fd_Inst[10]), .Z(n3447) );
  MUX21L U2495 ( .A(n1959), .B(n1958), .S(n3447), .Z(n1962) );
  NR2I U2496 ( .A(PC[11]), .B(fd_Inst[9]), .Z(n1961) );
  ND2I U2497 ( .A(PC[11]), .B(fd_Inst[9]), .Z(n1960) );
  ND2I U2498 ( .A(PC[10]), .B(fd_Inst[8]), .Z(n3406) );
  MUX21L U2499 ( .A(n1961), .B(n1960), .S(n3406), .Z(n3492) );
  MUX21L U2500 ( .A(n1963), .B(n1962), .S(n3492), .Z(n3462) );
  MUX21L U2501 ( .A(n1965), .B(n1964), .S(n3462), .Z(n1981) );
  NR2I U2502 ( .A(PC[10]), .B(fd_Inst[8]), .Z(n3405) );
  MUX21L U2503 ( .A(n1961), .B(n1960), .S(n3405), .Z(n3490) );
  MUX21L U2504 ( .A(n1963), .B(n1962), .S(n3490), .Z(n3461) );
  MUX21L U2505 ( .A(n1965), .B(n1964), .S(n3461), .Z(n1980) );
  NR2I U2506 ( .A(PC[9]), .B(fd_Inst[7]), .Z(n1967) );
  ND2I U2507 ( .A(PC[9]), .B(fd_Inst[7]), .Z(n1966) );
  ND2I U2508 ( .A(PC[8]), .B(fd_Inst[6]), .Z(n3728) );
  MUX21L U2509 ( .A(n1967), .B(n1966), .S(n3728), .Z(n1971) );
  NR2I U2510 ( .A(PC[8]), .B(fd_Inst[6]), .Z(n3729) );
  MUX21L U2511 ( .A(n1967), .B(n1966), .S(n3729), .Z(n1970) );
  NR2I U2512 ( .A(fd_Inst[5]), .B(PC[7]), .Z(n1969) );
  ND2I U2513 ( .A(fd_Inst[5]), .B(PC[7]), .Z(n1968) );
  NR2I U2514 ( .A(PC[6]), .B(fd_Inst[4]), .Z(n3700) );
  MUX21L U2515 ( .A(n1969), .B(n1968), .S(n3700), .Z(n3730) );
  MUX21L U2516 ( .A(n1971), .B(n1970), .S(n3730), .Z(n1979) );
  ND2I U2517 ( .A(PC[6]), .B(fd_Inst[4]), .Z(n3699) );
  MUX21L U2518 ( .A(n1969), .B(n1968), .S(n3699), .Z(n3731) );
  MUX21L U2519 ( .A(n1971), .B(n1970), .S(n3731), .Z(n1978) );
  NR2I U2520 ( .A(fd_Inst[3]), .B(PC[5]), .Z(n1973) );
  ND2I U2521 ( .A(fd_Inst[3]), .B(PC[5]), .Z(n1972) );
  ND2I U2522 ( .A(PC[4]), .B(fd_Inst[2]), .Z(n3681) );
  MUX21L U2523 ( .A(n1973), .B(n1972), .S(n3681), .Z(n1977) );
  NR2I U2524 ( .A(PC[4]), .B(fd_Inst[2]), .Z(n3682) );
  MUX21L U2525 ( .A(n1973), .B(n1972), .S(n3682), .Z(n1976) );
  NR2I U2526 ( .A(PC[3]), .B(fd_Inst[1]), .Z(n1975) );
  ND2I U2527 ( .A(PC[3]), .B(fd_Inst[1]), .Z(n1974) );
  ND2I U2528 ( .A(PC[2]), .B(fd_Inst[0]), .Z(n3668) );
  MUX21L U2529 ( .A(n1975), .B(n1974), .S(n3668), .Z(n3683) );
  MUX21L U2530 ( .A(n1977), .B(n1976), .S(n3683), .Z(n3732) );
  MUX21L U2531 ( .A(n1979), .B(n1978), .S(n3732), .Z(n3427) );
  MUX21LP U2532 ( .A(n1981), .B(n1980), .S(n3427), .Z(n3754) );
  MUX21L U2533 ( .A(n1983), .B(n1982), .S(n3754), .Z(n1989) );
  ND2I U2534 ( .A(n1985), .B(n1984), .Z(n1986) );
  IVI U2535 ( .A(n1986), .Z(n1988) );
  ND2I U2536 ( .A(n1988), .B(n1987), .Z(n3396) );
  ENI U2537 ( .A(n3396), .B(fd_Inst[26]), .Z(n3543) );
  AN2I U2538 ( .A(n3544), .B(n3543), .Z(n3637) );
  ND2I U2539 ( .A(n1989), .B(n3637), .Z(n1990) );
  ND2I U2540 ( .A(n1991), .B(n1990), .Z(n1140) );
  IVI U2541 ( .A(n1460), .Z(n1993) );
  MUX21H U2542 ( .A(mw_pc_plus_8[26]), .B(n2478), .S(n1993), .Z(
        gpr_wr_data[26]) );
  MUX21H U2543 ( .A(mw_pc_plus_8[24]), .B(n2473), .S(n1461), .Z(
        gpr_wr_data[24]) );
  MUX21H U2544 ( .A(mw_pc_plus_8[27]), .B(n2499), .S(n1993), .Z(
        gpr_wr_data[27]) );
  MUX21H U2545 ( .A(mw_pc_plus_8[30]), .B(n2500), .S(n1993), .Z(
        gpr_wr_data[30]) );
  MUX21H U2546 ( .A(mw_pc_plus_8[31]), .B(n2504), .S(n1461), .Z(
        gpr_wr_data[31]) );
  MUX21H U2547 ( .A(mw_pc_plus_8[2]), .B(n2372), .S(n1993), .Z(gpr_wr_data[2])
         );
  MUX21H U2548 ( .A(mw_pc_plus_8[15]), .B(n2424), .S(n1993), .Z(
        gpr_wr_data[15]) );
  MUX21H U2549 ( .A(mw_pc_plus_8[3]), .B(n2355), .S(n1461), .Z(gpr_wr_data[3])
         );
  MUX21H U2550 ( .A(mw_pc_plus_8[16]), .B(n2534), .S(n1461), .Z(
        gpr_wr_data[16]) );
  MUX21H U2551 ( .A(mw_pc_plus_8[19]), .B(n2450), .S(n1993), .Z(
        gpr_wr_data[19]) );
  MUX21H U2552 ( .A(mw_pc_plus_8[9]), .B(n2401), .S(n1993), .Z(gpr_wr_data[9])
         );
  MUX21H U2553 ( .A(mw_pc_plus_8[23]), .B(n2464), .S(n1993), .Z(
        gpr_wr_data[23]) );
  MUX21H U2554 ( .A(mw_pc_plus_8[20]), .B(n2459), .S(n1993), .Z(
        gpr_wr_data[20]) );
  MUX21H U2555 ( .A(mw_pc_plus_8[12]), .B(n2418), .S(n1993), .Z(
        gpr_wr_data[12]) );
  MUX21H U2556 ( .A(mw_pc_plus_8[13]), .B(n2415), .S(n1461), .Z(
        gpr_wr_data[13]) );
  MUX21H U2557 ( .A(mw_pc_plus_8[8]), .B(n2396), .S(n1993), .Z(gpr_wr_data[8])
         );
  IVI U2558 ( .A(n4706), .Z(n4707) );
  IVI U2559 ( .A(n4704), .Z(n4705) );
  IVI U2560 ( .A(n4708), .Z(n4709) );
  IVI U2561 ( .A(n4710), .Z(n4711) );
  NR2I U2562 ( .A(dx_Inst[29]), .B(dx_Inst[30]), .Z(n2010) );
  NR2I U2563 ( .A(dx_Inst[31]), .B(dx_Inst[27]), .Z(n1995) );
  AN2I U2564 ( .A(n2010), .B(n1995), .Z(n2182) );
  ND2I U2565 ( .A(dx_Inst[26]), .B(n4760), .Z(n1996) );
  ND2I U2566 ( .A(n2182), .B(n1996), .Z(n2098) );
  IVI U2567 ( .A(n2098), .Z(n2001) );
  NR2I U2568 ( .A(dx_Inst_15_0_signext[0]), .B(dx_Inst_15_0_signext[2]), .Z(
        n1997) );
  ND2I U2569 ( .A(n1997), .B(n4769), .Z(n2183) );
  NR2I U2570 ( .A(dx_Inst[28]), .B(dx_Inst[26]), .Z(n2174) );
  NR2I U2571 ( .A(dx_Inst_15_0_signext[3]), .B(dx_Inst_15_0_signext[5]), .Z(
        n1998) );
  ND2I U2572 ( .A(n2174), .B(n1998), .Z(n1999) );
  NR2I U2573 ( .A(n2183), .B(n1999), .Z(n2000) );
  ND2I U2574 ( .A(n2182), .B(n2000), .Z(n2262) );
  AN2I U2575 ( .A(n2001), .B(n2262), .Z(n2260) );
  ENI U2576 ( .A(dx_Inst[17]), .B(xm_Inst[12]), .Z(n2002) );
  AO7P U2577 ( .A(n2002), .B(n2006), .C(n4755), .Z(n2003) );
  IVI U2578 ( .A(n2003), .Z(n2008) );
  ENI U2579 ( .A(n2004), .B(dx_Inst[17]), .Z(n2005) );
  ND2I U2580 ( .A(n2006), .B(n2005), .Z(n2007) );
  ND2I U2581 ( .A(n2008), .B(n2007), .Z(n2045) );
  NR2I U2582 ( .A(dx_Inst[16]), .B(dx_Inst[18]), .Z(n2009) );
  ND4 U2583 ( .A(n2009), .B(n4716), .C(n4756), .D(n4782), .Z(n2012) );
  ND2I U2584 ( .A(n2010), .B(dx_Inst[31]), .Z(n2011) );
  AN2I U2585 ( .A(n2012), .B(n2011), .Z(n2021) );
  AN2I U2586 ( .A(n4867), .B(n4868), .Z(n2014) );
  AN2I U2587 ( .A(n4865), .B(n4866), .Z(n2013) );
  ND2I U2588 ( .A(n2014), .B(n2013), .Z(n2015) );
  IVI U2589 ( .A(n2015), .Z(n3950) );
  ND2I U2590 ( .A(n4870), .B(n4869), .Z(n2017) );
  ND2I U2591 ( .A(n4872), .B(n4871), .Z(n2016) );
  NR2I U2592 ( .A(n2017), .B(n2016), .Z(n2018) );
  ND2I U2593 ( .A(n2019), .B(n2018), .Z(n2020) );
  IVI U2594 ( .A(n2020), .Z(n3949) );
  ND2I U2595 ( .A(n3950), .B(n3949), .Z(n3952) );
  ND2I U2596 ( .A(n2021), .B(n3952), .Z(n2041) );
  ND2I U2597 ( .A(n2023), .B(n2022), .Z(n2024) );
  ENI U2598 ( .A(n2024), .B(n4762), .Z(n2029) );
  ND2I U2599 ( .A(n2026), .B(n2025), .Z(n2027) );
  ENI U2600 ( .A(n2027), .B(n4782), .Z(n2028) );
  ND2I U2601 ( .A(n2029), .B(n2028), .Z(n2046) );
  ND2I U2602 ( .A(n2031), .B(n2030), .Z(n2032) );
  ENI U2603 ( .A(n2032), .B(n4777), .Z(n2042) );
  ND2I U2604 ( .A(n2034), .B(n2033), .Z(n2035) );
  ENI U2605 ( .A(n2035), .B(n4756), .Z(n2043) );
  ND2I U2606 ( .A(n2042), .B(n2043), .Z(n2036) );
  NR2I U2607 ( .A(n2046), .B(n2036), .Z(n2065) );
  ND2I U2608 ( .A(n2066), .B(n2065), .Z(n2068) );
  ND2I U2609 ( .A(n2260), .B(n2068), .Z(n2302) );
  ENI U2610 ( .A(n3762), .B(dx_Inst[16]), .Z(n2073) );
  IVI U2611 ( .A(n2073), .Z(n2040) );
  ENI U2612 ( .A(gpr_wr_addr[2]), .B(dx_Inst[18]), .Z(n2074) );
  ND2I U2613 ( .A(n2060), .B(n2037), .Z(n2349) );
  ENI U2614 ( .A(n2349), .B(dx_Inst[17]), .Z(n2075) );
  ND2I U2615 ( .A(n2074), .B(n2075), .Z(n2039) );
  NR2I U2616 ( .A(n2040), .B(n2039), .Z(n2064) );
  IVI U2617 ( .A(n2342), .Z(n4695) );
  NR2I U2618 ( .A(n4695), .B(n2041), .Z(n2050) );
  ND2I U2619 ( .A(n2043), .B(n2042), .Z(n2044) );
  NR2I U2620 ( .A(n2045), .B(n2044), .Z(n2048) );
  IVI U2621 ( .A(n2046), .Z(n2047) );
  ND2I U2622 ( .A(n2048), .B(n2047), .Z(n2049) );
  ND2I U2623 ( .A(n2050), .B(n2049), .Z(n2072) );
  IVI U2624 ( .A(n2053), .Z(n2052) );
  IVI U2625 ( .A(n2056), .Z(n2051) );
  AO7P U2626 ( .A(n2052), .B(n2051), .C(dx_Inst[19]), .Z(n2058) );
  ND2I U2627 ( .A(n2053), .B(n4782), .Z(n2054) );
  IVI U2628 ( .A(n2054), .Z(n2055) );
  ND2I U2629 ( .A(n2056), .B(n2055), .Z(n2057) );
  ND2I U2630 ( .A(n2058), .B(n2057), .Z(n2078) );
  ND2I U2631 ( .A(n1992), .B(n2059), .Z(n2061) );
  ENI U2632 ( .A(n2061), .B(dx_Inst[20]), .Z(n2076) );
  ND2I U2633 ( .A(n2078), .B(n2076), .Z(n2062) );
  NR2I U2634 ( .A(n2072), .B(n2062), .Z(n2063) );
  AN2I U2635 ( .A(n2064), .B(n2063), .Z(n2309) );
  IVI U2636 ( .A(n2309), .Z(n2254) );
  ND2I U2637 ( .A(n2307), .B(n2254), .Z(n2204) );
  IVI U2638 ( .A(n2204), .Z(n3248) );
  ND2I U2639 ( .A(n2066), .B(n2065), .Z(n2283) );
  ND2I U2640 ( .A(n2283), .B(n2098), .Z(n2318) );
  NR2I U2641 ( .A(n2318), .B(n4794), .Z(n2067) );
  IVI U2642 ( .A(n2309), .Z(n2106) );
  ND2I U2643 ( .A(n2067), .B(n2106), .Z(n3246) );
  IVI U2644 ( .A(n2309), .Z(n2289) );
  IVI U2645 ( .A(n2254), .Z(n2155) );
  ND2I U2646 ( .A(n4691), .B(n2155), .Z(n2070) );
  IVI U2647 ( .A(n2068), .Z(n2293) );
  B4I U2648 ( .A(n2293), .Z(n2102) );
  IVI U2649 ( .A(n2102), .Z(n2278) );
  ND2I U2650 ( .A(n2278), .B(Addr[29]), .Z(n2069) );
  ND2I U2651 ( .A(n3248), .B(dx_gpr_rd_data2[30]), .Z(n2071) );
  AN2I U2652 ( .A(n2071), .B(n4146), .Z(n2087) );
  IVI U2653 ( .A(n2072), .Z(n2083) );
  ND2I U2654 ( .A(n2074), .B(n2073), .Z(n2081) );
  ND2I U2655 ( .A(n2076), .B(n2075), .Z(n2077) );
  IVI U2656 ( .A(n2077), .Z(n2079) );
  ND2I U2657 ( .A(n2079), .B(n2078), .Z(n2080) );
  NR2I U2658 ( .A(n2081), .B(n2080), .Z(n2082) );
  ND2I U2659 ( .A(n2083), .B(n2082), .Z(n2161) );
  IVI U2660 ( .A(n2319), .Z(n2249) );
  ND2I U2661 ( .A(n2500), .B(n2249), .Z(n2085) );
  ND2I U2662 ( .A(n2278), .B(Addr[30]), .Z(n2084) );
  AN2I U2663 ( .A(n2085), .B(n2084), .Z(n2086) );
  ND2I U2664 ( .A(n2087), .B(n2086), .Z(n4604) );
  NR2I U2665 ( .A(n4142), .B(n4604), .Z(n2115) );
  IVI U2666 ( .A(n2102), .Z(n2310) );
  B2IP U2667 ( .A(n2161), .Z1(n2292), .Z2(n2319) );
  IVI U2668 ( .A(n2204), .Z(n2700) );
  ND2I U2669 ( .A(dx_gpr_rd_data2[28]), .B(n3254), .Z(n4140) );
  ND2I U2670 ( .A(n4139), .B(n4140), .Z(n4397) );
  ND2I U2671 ( .A(n2278), .B(Addr[26]), .Z(n2089) );
  IVI U2672 ( .A(n2319), .Z(n2215) );
  ND2I U2673 ( .A(n2478), .B(n2215), .Z(n2088) );
  ND2I U2674 ( .A(n2089), .B(n2088), .Z(n3216) );
  NR2I U2675 ( .A(n4397), .B(n3216), .Z(n2112) );
  ND2I U2676 ( .A(n2504), .B(n2215), .Z(n2091) );
  ND2I U2677 ( .A(n2278), .B(Addr[31]), .Z(n2090) );
  ND2I U2678 ( .A(n2091), .B(n2090), .Z(n2092) );
  IVI U2679 ( .A(n2092), .Z(n2093) );
  ND2I U2680 ( .A(n4146), .B(n2093), .Z(n3200) );
  B5IP U2681 ( .A(n2102), .Z(n2291) );
  ND2I U2682 ( .A(Addr[7]), .B(n2291), .Z(n2095) );
  ND2I U2683 ( .A(n4681), .B(n2155), .Z(n2094) );
  ND2I U2684 ( .A(n2095), .B(n2094), .Z(n2096) );
  IVI U2685 ( .A(n2096), .Z(n2612) );
  AN2I U2686 ( .A(n2307), .B(dx_gpr_rd_data2[7]), .Z(n2097) );
  ND2I U2687 ( .A(n2319), .B(n2097), .Z(n2101) );
  AN2I U2688 ( .A(n2296), .B(dx_Inst_15_0_signext[7]), .Z(n2099) );
  ND2I U2689 ( .A(n2319), .B(n2099), .Z(n2100) );
  AN2I U2690 ( .A(n2101), .B(n2100), .Z(n2611) );
  ND2I U2691 ( .A(n2612), .B(n2611), .Z(n3880) );
  NR2I U2692 ( .A(n3200), .B(n3880), .Z(n2111) );
  OR2I U2693 ( .A(n4703), .B(n2102), .Z(n2104) );
  ND2I U2694 ( .A(n2292), .B(n4679), .Z(n2103) );
  ND2I U2695 ( .A(n2104), .B(n2103), .Z(n2105) );
  IVI U2696 ( .A(n2105), .Z(n2108) );
  AN2I U2697 ( .A(n2296), .B(n2106), .Z(n2252) );
  ND2I U2698 ( .A(n2252), .B(dx_Inst_15_0_signext[5]), .Z(n2107) );
  ND2I U2699 ( .A(n2108), .B(n2107), .Z(n2109) );
  IVI U2700 ( .A(n2109), .Z(n2631) );
  ND2I U2701 ( .A(n2700), .B(dx_gpr_rd_data2[5]), .Z(n2632) );
  ND2I U2702 ( .A(n2631), .B(n2632), .Z(n2110) );
  ND2I U2703 ( .A(n2112), .B(n1442), .Z(n2113) );
  IVI U2704 ( .A(n2113), .Z(n2114) );
  ND2I U2705 ( .A(n2115), .B(n2114), .Z(n2116) );
  IVI U2706 ( .A(n2116), .Z(n2442) );
  ND2I U2707 ( .A(n2252), .B(dx_Inst_15_0_signext[14]), .Z(n2118) );
  IVI U2708 ( .A(n2204), .Z(n3254) );
  ND2I U2709 ( .A(n2700), .B(dx_gpr_rd_data2[14]), .Z(n2117) );
  AN2I U2710 ( .A(n2118), .B(n2117), .Z(n2123) );
  ND2I U2711 ( .A(n2278), .B(Addr[14]), .Z(n2120) );
  ND2I U2712 ( .A(n4684), .B(n1270), .Z(n2119) );
  ND2I U2713 ( .A(n2120), .B(n2119), .Z(n2121) );
  IVI U2714 ( .A(n2121), .Z(n2122) );
  ND2I U2715 ( .A(n2123), .B(n2122), .Z(n3024) );
  IVI U2716 ( .A(n3024), .Z(n2124) );
  ND2I U2717 ( .A(Addr[17]), .B(n2291), .Z(n2695) );
  ND2I U2718 ( .A(n4685), .B(n2249), .Z(n2692) );
  ND2I U2719 ( .A(n2124), .B(n1452), .Z(n2134) );
  IVI U2720 ( .A(n2418), .Z(n2125) );
  OR2I U2721 ( .A(n2125), .B(n2319), .Z(n2127) );
  ND2I U2722 ( .A(Addr[12]), .B(n2291), .Z(n2126) );
  ND2I U2723 ( .A(n2127), .B(n2126), .Z(n2128) );
  IVI U2724 ( .A(n2128), .Z(n2133) );
  ND2I U2725 ( .A(dx_gpr_rd_data2[12]), .B(n3218), .Z(n2130) );
  ND2I U2726 ( .A(n2252), .B(dx_Inst_15_0_signext[12]), .Z(n2129) );
  ND2I U2727 ( .A(n2130), .B(n2129), .Z(n2131) );
  IVI U2728 ( .A(n2131), .Z(n2132) );
  ND2I U2729 ( .A(n2133), .B(n2132), .Z(n2569) );
  NR2I U2730 ( .A(n2134), .B(n1154), .Z(n2171) );
  ND2I U2731 ( .A(n2278), .B(Addr[18]), .Z(n2135) );
  ND2I U2732 ( .A(n2136), .B(n2135), .Z(n2137) );
  IVI U2733 ( .A(n2137), .Z(n2138) );
  ND2I U2734 ( .A(n4146), .B(n2138), .Z(n2688) );
  ND2I U2735 ( .A(n2252), .B(dx_Inst_15_0_signext[13]), .Z(n2140) );
  ND2I U2736 ( .A(Addr[13]), .B(n2291), .Z(n2139) );
  AN2I U2737 ( .A(n2140), .B(n2139), .Z(n2146) );
  ND2I U2738 ( .A(n3218), .B(dx_gpr_rd_data2[13]), .Z(n2143) );
  IVI U2739 ( .A(n2415), .Z(n2141) );
  OR2I U2740 ( .A(n2141), .B(n2319), .Z(n2142) );
  ND2I U2741 ( .A(n2143), .B(n2142), .Z(n2144) );
  IVI U2742 ( .A(n2144), .Z(n2145) );
  ND2I U2743 ( .A(n2146), .B(n2145), .Z(n3302) );
  IVI U2744 ( .A(n3302), .Z(n2147) );
  ND2I U2745 ( .A(n2689), .B(n2147), .Z(n2169) );
  ND2I U2746 ( .A(Addr[11]), .B(n2291), .Z(n2149) );
  ND2I U2747 ( .A(dx_gpr_rd_data2[11]), .B(n3218), .Z(n2148) );
  AN2I U2748 ( .A(n2149), .B(n2148), .Z(n2153) );
  IVI U2749 ( .A(n2319), .Z(n2270) );
  ND2I U2750 ( .A(n4683), .B(n2270), .Z(n2151) );
  ND2I U2751 ( .A(n2252), .B(dx_Inst_15_0_signext[11]), .Z(n2150) );
  AN2I U2752 ( .A(n2151), .B(n2150), .Z(n2152) );
  ND2I U2753 ( .A(n2153), .B(n2152), .Z(n2855) );
  IVI U2754 ( .A(n2855), .Z(n2167) );
  AN2I U2755 ( .A(n2307), .B(dx_gpr_rd_data2[15]), .Z(n2154) );
  ND2I U2756 ( .A(n2289), .B(n2154), .Z(n2160) );
  ND2I U2757 ( .A(n2424), .B(n2155), .Z(n2157) );
  ND2I U2758 ( .A(Addr[15]), .B(n2291), .Z(n2156) );
  ND2I U2759 ( .A(n2157), .B(n2156), .Z(n2158) );
  IVI U2760 ( .A(n2158), .Z(n2159) );
  AN2I U2761 ( .A(n2160), .B(n2159), .Z(n3056) );
  ND2I U2762 ( .A(n3056), .B(n4146), .Z(n2560) );
  ND2I U2763 ( .A(Addr[16]), .B(n2291), .Z(n2164) );
  IVI U2764 ( .A(n2534), .Z(n2162) );
  OR2I U2765 ( .A(n2162), .B(n2319), .Z(n2163) );
  AN2I U2766 ( .A(n2164), .B(n2163), .Z(n2165) );
  ND2I U2767 ( .A(n2165), .B(n4146), .Z(n2701) );
  NR2I U2768 ( .A(n2560), .B(n2701), .Z(n2166) );
  ND2I U2769 ( .A(n2167), .B(n2166), .Z(n2168) );
  NR2I U2770 ( .A(n2169), .B(n2168), .Z(n2170) );
  ND2I U2771 ( .A(n2171), .B(n2170), .Z(n2443) );
  NR2I U2772 ( .A(dx_Inst[30]), .B(dx_Inst[31]), .Z(n2192) );
  NR2I U2773 ( .A(dx_Inst[26]), .B(n4754), .Z(n2172) );
  AN2I U2774 ( .A(n2192), .B(n2172), .Z(n2178) );
  ND2I U2775 ( .A(dx_Inst[28]), .B(n2178), .Z(n2173) );
  AN2I U2776 ( .A(n2262), .B(n2173), .Z(n2177) );
  IVI U2777 ( .A(n2197), .Z(n2190) );
  NR2I U2778 ( .A(dx_Inst_15_0_signext[0]), .B(n4770), .Z(n2175) );
  ND2I U2779 ( .A(n2190), .B(n2175), .Z(n2176) );
  AN2I U2780 ( .A(n2177), .B(n2176), .Z(n2707) );
  ND2I U2781 ( .A(dx_Inst[27]), .B(n2178), .Z(n2188) );
  ND2I U2782 ( .A(dx_Inst_15_0_signext[1]), .B(n4760), .Z(n2181) );
  ND2I U2783 ( .A(dx_Inst_15_0_signext[3]), .B(n4771), .Z(n2179) );
  ND2I U2784 ( .A(n4761), .B(n2179), .Z(n2180) );
  NR2I U2785 ( .A(n2181), .B(n2180), .Z(n2186) );
  IVI U2786 ( .A(n2182), .Z(n2184) );
  NR2I U2787 ( .A(n2184), .B(n2183), .Z(n2185) );
  ND2I U2788 ( .A(n2186), .B(n2185), .Z(n2187) );
  AN2I U2789 ( .A(n2188), .B(n2187), .Z(n2191) );
  NR2I U2790 ( .A(dx_Inst_15_0_signext[0]), .B(n4773), .Z(n2189) );
  ND2I U2791 ( .A(n2190), .B(n2189), .Z(n2195) );
  ND2I U2792 ( .A(n2191), .B(n2195), .Z(n2558) );
  NR2I U2793 ( .A(n2707), .B(n2558), .Z(n2201) );
  ENI U2794 ( .A(n4761), .B(dx_Inst[27]), .Z(n2193) );
  ND4 U2795 ( .A(n2193), .B(n2192), .C(dx_Inst[29]), .D(dx_Inst[28]), .Z(n2194) );
  AN2I U2796 ( .A(n2195), .B(n2194), .Z(n2200) );
  ND2I U2797 ( .A(dx_Inst_15_0_signext[0]), .B(dx_Inst_15_0_signext[2]), .Z(
        n2196) );
  ND2I U2798 ( .A(n4773), .B(n2198), .Z(n2199) );
  ND2I U2799 ( .A(n2200), .B(n2199), .Z(n3386) );
  ND2I U2800 ( .A(n2201), .B(n3386), .Z(n2202) );
  NR2I U2801 ( .A(n2443), .B(n2202), .Z(n2203) );
  AN2I U2802 ( .A(n2442), .B(n2203), .Z(n2807) );
  IVI U2803 ( .A(n2204), .Z(n3218) );
  ND2I U2804 ( .A(dx_gpr_rd_data2[27]), .B(n2700), .Z(n2205) );
  ND2I U2805 ( .A(n4146), .B(n2205), .Z(n2206) );
  IVI U2806 ( .A(n2206), .Z(n3214) );
  ND2I U2807 ( .A(n3220), .B(n3214), .Z(n2212) );
  ND2I U2808 ( .A(n2278), .B(Addr[24]), .Z(n2208) );
  ND2I U2809 ( .A(n2473), .B(n2270), .Z(n2207) );
  ND2I U2810 ( .A(n2208), .B(n2207), .Z(n2209) );
  IVI U2811 ( .A(n2209), .Z(n3221) );
  ND2I U2812 ( .A(n2499), .B(n1270), .Z(n2211) );
  ND2I U2813 ( .A(n2278), .B(Addr[27]), .Z(n2210) );
  AN2I U2814 ( .A(n2211), .B(n2210), .Z(n3215) );
  ND2I U2815 ( .A(n2450), .B(n2249), .Z(n2485) );
  AN2I U2816 ( .A(n2291), .B(Addr[19]), .Z(n2483) );
  IVI U2817 ( .A(n2483), .Z(n2213) );
  ND2I U2818 ( .A(Addr[20]), .B(n2291), .Z(n4054) );
  ND2I U2819 ( .A(n2459), .B(n2215), .Z(n4058) );
  ND2I U2820 ( .A(n4054), .B(n4058), .Z(n3247) );
  NR2I U2821 ( .A(n1443), .B(n3247), .Z(n2214) );
  ND2I U2822 ( .A(Addr[21]), .B(n2291), .Z(n2217) );
  ND2I U2823 ( .A(n4687), .B(n2215), .Z(n2216) );
  ND2I U2824 ( .A(n2217), .B(n2216), .Z(n2218) );
  NR2I U2825 ( .A(n2218), .B(n4056), .Z(n3244) );
  ND2I U2826 ( .A(Addr[23]), .B(n2291), .Z(n2220) );
  ND2I U2827 ( .A(n2464), .B(n2249), .Z(n2219) );
  ND2I U2828 ( .A(n2220), .B(n2219), .Z(n3253) );
  AN2I U2829 ( .A(n3244), .B(n3259), .Z(n2444) );
  ND2I U2830 ( .A(n4688), .B(n1270), .Z(n2222) );
  ND2I U2831 ( .A(n2278), .B(Addr[22]), .Z(n2221) );
  ND2I U2832 ( .A(n2222), .B(n2221), .Z(n2223) );
  IVI U2833 ( .A(n2223), .Z(n4171) );
  AN2I U2834 ( .A(n4171), .B(n4146), .Z(n3252) );
  ND2I U2835 ( .A(n2278), .B(Addr[25]), .Z(n2225) );
  ND2I U2836 ( .A(n4689), .B(n1270), .Z(n2224) );
  ND2I U2837 ( .A(n2225), .B(n2224), .Z(n2226) );
  IVI U2838 ( .A(n2226), .Z(n2227) );
  AN2I U2839 ( .A(n4146), .B(n2227), .Z(n3222) );
  ND2I U2840 ( .A(n3252), .B(n3222), .Z(n2446) );
  IVI U2841 ( .A(n2446), .Z(n2228) );
  ND2I U2842 ( .A(n2444), .B(n2228), .Z(n2229) );
  IVI U2843 ( .A(n2229), .Z(n2230) );
  ND2I U2844 ( .A(n2448), .B(n2230), .Z(n2842) );
  ND2I U2845 ( .A(dx_Inst_15_0_signext[9]), .B(n2252), .Z(n2237) );
  ND2I U2846 ( .A(n2307), .B(dx_gpr_rd_data2[9]), .Z(n2231) );
  IVI U2847 ( .A(n2231), .Z(n2232) );
  ND2I U2848 ( .A(n2289), .B(n2232), .Z(n2234) );
  ND2I U2849 ( .A(n2291), .B(Addr[9]), .Z(n2233) );
  ND2I U2850 ( .A(n2234), .B(n2233), .Z(n2235) );
  NR2I U2851 ( .A(n1453), .B(n2235), .Z(n2236) );
  ND2I U2852 ( .A(n2237), .B(n2236), .Z(n3088) );
  ND2I U2853 ( .A(dx_gpr_rd_data2[10]), .B(n3218), .Z(n2239) );
  ND2I U2854 ( .A(n2252), .B(dx_Inst_15_0_signext[10]), .Z(n2238) );
  ND2I U2855 ( .A(n2239), .B(n2238), .Z(n2240) );
  IVI U2856 ( .A(n2240), .Z(n2245) );
  ND2I U2857 ( .A(Addr[10]), .B(n2291), .Z(n2242) );
  ND2I U2858 ( .A(n2270), .B(n4682), .Z(n2241) );
  ND2I U2859 ( .A(n2242), .B(n2241), .Z(n2243) );
  IVI U2860 ( .A(n2243), .Z(n2244) );
  ND2I U2861 ( .A(n2245), .B(n2244), .Z(n3322) );
  NR2I U2862 ( .A(n3088), .B(n3322), .Z(n2440) );
  ND2I U2863 ( .A(Addr[8]), .B(n2291), .Z(n2582) );
  ND2I U2864 ( .A(n2396), .B(n2249), .Z(n2583) );
  ND2I U2865 ( .A(n2582), .B(n2583), .Z(n2247) );
  ND2I U2866 ( .A(n2252), .B(dx_Inst_15_0_signext[8]), .Z(n2581) );
  IVI U2867 ( .A(n2581), .Z(n2246) );
  NR2I U2868 ( .A(n2247), .B(n2246), .Z(n2248) );
  ND2I U2869 ( .A(dx_gpr_rd_data2[8]), .B(n3248), .Z(n2584) );
  ND2I U2870 ( .A(n2248), .B(n2584), .Z(n2437) );
  ND2I U2871 ( .A(Addr[6]), .B(n2291), .Z(n2251) );
  ND2I U2872 ( .A(n2249), .B(n4680), .Z(n2250) );
  AN2I U2873 ( .A(n2251), .B(n2250), .Z(n2435) );
  ND2I U2874 ( .A(dx_Inst_15_0_signext[6]), .B(n2252), .Z(n2257) );
  ND2I U2875 ( .A(n2307), .B(dx_gpr_rd_data2[6]), .Z(n2253) );
  IVI U2876 ( .A(n2253), .Z(n2255) );
  ND2I U2877 ( .A(n2255), .B(n2289), .Z(n2256) );
  AN2I U2878 ( .A(n2257), .B(n2256), .Z(n2434) );
  ND2I U2879 ( .A(n2435), .B(n2434), .Z(n3861) );
  NR2I U2880 ( .A(n2437), .B(n3861), .Z(n2258) );
  ND2I U2881 ( .A(n2440), .B(n2258), .Z(n2259) );
  NR2I U2882 ( .A(n2842), .B(n2259), .Z(n2409) );
  ND2I U2883 ( .A(n2807), .B(n1169), .Z(n2382) );
  IVI U2884 ( .A(n2382), .Z(n4029) );
  ND2I U2885 ( .A(dx_Inst_15_0_signext[4]), .B(n2296), .Z(n2268) );
  ND2I U2886 ( .A(n2260), .B(n2283), .Z(n2271) );
  NR2I U2887 ( .A(n2271), .B(n4819), .Z(n2261) );
  IVI U2888 ( .A(n2261), .Z(n2265) );
  IVI U2889 ( .A(n2262), .Z(n2284) );
  ND2I U2890 ( .A(n2284), .B(n2283), .Z(n2316) );
  NR2I U2891 ( .A(n2316), .B(n4820), .Z(n2263) );
  IVI U2892 ( .A(n2263), .Z(n2264) );
  ND2I U2893 ( .A(n2265), .B(n2264), .Z(n2266) );
  IVI U2894 ( .A(n2266), .Z(n2267) );
  ND2I U2895 ( .A(n2268), .B(n2267), .Z(n2269) );
  ND2I U2896 ( .A(n2319), .B(n2269), .Z(n2623) );
  ND2I U2897 ( .A(n4678), .B(n2270), .Z(n2627) );
  ND2I U2898 ( .A(Addr[4]), .B(n2278), .Z(n2624) );
  ND2I U2899 ( .A(n2627), .B(n1159), .Z(n3928) );
  IVDA U2900 ( .A(n3928), .Y(n1456), .Z(n2752) );
  NR2I U2901 ( .A(n2271), .B(n4821), .Z(n2276) );
  IVI U2902 ( .A(n2316), .Z(n2272) );
  ND2I U2903 ( .A(n2272), .B(dx_Inst_15_0_signext[8]), .Z(n2274) );
  ND2I U2904 ( .A(dx_Inst_15_0_signext[2]), .B(n2296), .Z(n2273) );
  ND2I U2905 ( .A(n2274), .B(n2273), .Z(n2275) );
  AO7 U2906 ( .A(n2276), .B(n2275), .C(n2319), .Z(n2282) );
  IVI U2907 ( .A(n2319), .Z(n2277) );
  ND2I U2908 ( .A(n2372), .B(n2277), .Z(n2280) );
  ND2I U2909 ( .A(n2278), .B(Addr[2]), .Z(n2279) );
  AN2I U2910 ( .A(n2280), .B(n2279), .Z(n2281) );
  ND2I U2911 ( .A(n2282), .B(n2281), .Z(n2664) );
  IVI U2912 ( .A(n2664), .Z(n3871) );
  AN2I U2913 ( .A(n2307), .B(dx_gpr_rd_data2[3]), .Z(n2286) );
  ND2I U2914 ( .A(n2284), .B(n2283), .Z(n2301) );
  NR2I U2915 ( .A(n2301), .B(n4822), .Z(n2285) );
  NR2I U2916 ( .A(n2286), .B(n2285), .Z(n2287) );
  IVI U2917 ( .A(n2287), .Z(n2288) );
  ND2I U2918 ( .A(n2289), .B(n2288), .Z(n2646) );
  AN2I U2919 ( .A(dx_Inst_15_0_signext[3]), .B(n2296), .Z(n2290) );
  ND2I U2920 ( .A(n2290), .B(n2289), .Z(n2653) );
  AN2I U2921 ( .A(n2646), .B(n2653), .Z(n2502) );
  ND2I U2922 ( .A(Addr[3]), .B(n2291), .Z(n2649) );
  ND2I U2923 ( .A(n2355), .B(n2292), .Z(n2650) );
  AN2I U2924 ( .A(n2649), .B(n2650), .Z(n2501) );
  ND2I U2925 ( .A(n2502), .B(n2501), .Z(n3920) );
  IVI U2926 ( .A(n3920), .Z(n2533) );
  AN2I U2927 ( .A(n3871), .B(n2533), .Z(n3856) );
  AN2I U2928 ( .A(n2752), .B(n3856), .Z(n4027) );
  AN2I U2929 ( .A(n4029), .B(n4027), .Z(n4461) );
  ND2I U2930 ( .A(n4676), .B(n2309), .Z(n2295) );
  ND2I U2931 ( .A(Addr[0]), .B(n2293), .Z(n2294) );
  AN2I U2932 ( .A(n2295), .B(n2294), .Z(n2299) );
  AN2I U2933 ( .A(dx_Inst_15_0_signext[0]), .B(n2296), .Z(n2297) );
  ND2I U2934 ( .A(n2319), .B(n2297), .Z(n2298) );
  ND2I U2935 ( .A(n2299), .B(n2298), .Z(n2300) );
  IVI U2936 ( .A(n2300), .Z(n2667) );
  NR2I U2937 ( .A(n2301), .B(n4796), .Z(n2304) );
  NR2I U2938 ( .A(n1459), .B(n2302), .Z(n2303) );
  NR2I U2939 ( .A(n2304), .B(n2303), .Z(n2305) );
  IVI U2940 ( .A(n2305), .Z(n2306) );
  ND2I U2941 ( .A(n2319), .B(n2306), .Z(n2668) );
  ND2I U2942 ( .A(n2667), .B(n2668), .Z(n2919) );
  IVI U2943 ( .A(n2919), .Z(n2379) );
  AN2I U2944 ( .A(n2307), .B(dx_gpr_rd_data2[1]), .Z(n2308) );
  ND2I U2945 ( .A(n2319), .B(n2308), .Z(n2315) );
  ND2I U2946 ( .A(n4677), .B(n2309), .Z(n2312) );
  ND2I U2947 ( .A(n2310), .B(Addr[1]), .Z(n2311) );
  ND2I U2948 ( .A(n2312), .B(n2311), .Z(n2313) );
  IVI U2949 ( .A(n2313), .Z(n2314) );
  AN2I U2950 ( .A(n2315), .B(n2314), .Z(n2378) );
  NR2I U2951 ( .A(n2316), .B(n4795), .Z(n2317) );
  ND2I U2952 ( .A(n2317), .B(n2319), .Z(n2322) );
  NR2I U2953 ( .A(n4773), .B(n2318), .Z(n2320) );
  ND2I U2954 ( .A(n2320), .B(n2319), .Z(n2321) );
  AN2I U2955 ( .A(n2322), .B(n2321), .Z(n2377) );
  ND2I U2956 ( .A(n2378), .B(n2377), .Z(n2666) );
  IVI U2957 ( .A(n2666), .Z(n2921) );
  AN2I U2958 ( .A(n2379), .B(n2921), .Z(n2503) );
  IVI U2959 ( .A(n2720), .Z(n2922) );
  ENI U2960 ( .A(n2323), .B(n4775), .Z(n2324) );
  ND2I U2961 ( .A(n4755), .B(n2324), .Z(n2330) );
  ENI U2962 ( .A(n2325), .B(n4774), .Z(n2328) );
  ENI U2963 ( .A(n2326), .B(n4776), .Z(n2327) );
  ND2I U2964 ( .A(n2328), .B(n2327), .Z(n2329) );
  NR2I U2965 ( .A(n2330), .B(n2329), .Z(n2336) );
  ENI U2966 ( .A(n2331), .B(dx_gpr_rd_addr1[2]), .Z(n2334) );
  ENI U2967 ( .A(n2332), .B(dx_gpr_rd_addr1[3]), .Z(n2333) );
  NR2I U2968 ( .A(n2334), .B(n2333), .Z(n2335) );
  ND2I U2969 ( .A(n2336), .B(n2335), .Z(n2347) );
  IVI U2970 ( .A(n2347), .Z(n2340) );
  NR2I U2971 ( .A(dx_gpr_rd_addr1[2]), .B(dx_gpr_rd_addr1[1]), .Z(n2339) );
  NR2I U2972 ( .A(dx_gpr_rd_addr1[4]), .B(dx_gpr_rd_addr1[3]), .Z(n2337) );
  AN2I U2973 ( .A(n2337), .B(n4774), .Z(n2338) );
  ND2I U2974 ( .A(n2339), .B(n2338), .Z(n2341) );
  ND2I U2975 ( .A(n2340), .B(n2341), .Z(n2394) );
  IVI U2976 ( .A(n2394), .Z(n2514) );
  ND2I U2977 ( .A(Addr[3]), .B(n2514), .Z(n2357) );
  ENI U2978 ( .A(gpr_wr_addr[3]), .B(dx_gpr_rd_addr1[3]), .Z(n2344) );
  AN2I U2979 ( .A(n2342), .B(n2341), .Z(n2343) );
  ND2I U2980 ( .A(n2344), .B(n2343), .Z(n2345) );
  IVI U2981 ( .A(n2345), .Z(n2346) );
  ND2I U2982 ( .A(n2347), .B(n2346), .Z(n2348) );
  IVI U2983 ( .A(n2348), .Z(n2361) );
  ENI U2984 ( .A(n2349), .B(dx_gpr_rd_addr1[1]), .Z(n2351) );
  ENI U2985 ( .A(gpr_wr_addr[2]), .B(dx_gpr_rd_addr1[2]), .Z(n2350) );
  ND2I U2986 ( .A(n2351), .B(n2350), .Z(n2359) );
  ENI U2987 ( .A(n3762), .B(dx_gpr_rd_addr1[0]), .Z(n2353) );
  ENI U2988 ( .A(n4874), .B(dx_gpr_rd_addr1[4]), .Z(n2352) );
  ND2I U2989 ( .A(n2353), .B(n2352), .Z(n2358) );
  NR2I U2990 ( .A(n2359), .B(n2358), .Z(n2354) );
  ND2I U2991 ( .A(n2361), .B(n2354), .Z(n2383) );
  IVI U2992 ( .A(n2383), .Z(n2515) );
  ND2I U2993 ( .A(n2355), .B(n2515), .Z(n2356) );
  AN2I U2994 ( .A(n2357), .B(n2356), .Z(n2364) );
  NR2I U2995 ( .A(n2359), .B(n2358), .Z(n2360) );
  ND2I U2996 ( .A(n2361), .B(n2360), .Z(n2362) );
  ND2I U2997 ( .A(n1213), .B(n2362), .Z(n2389) );
  ND2I U2998 ( .A(n1208), .B(dx_gpr_rd_data1[3]), .Z(n2363) );
  ND2I U2999 ( .A(n2364), .B(n2363), .Z(n3136) );
  ND2I U3000 ( .A(n2922), .B(n3136), .Z(n2371) );
  ND2I U3001 ( .A(n2666), .B(n2919), .Z(n2365) );
  B5IP U3002 ( .A(n2365), .Z(n3013) );
  IVI U3003 ( .A(n2383), .Z(n2526) );
  ND2I U3004 ( .A(n4676), .B(n2526), .Z(n2367) );
  IVI U3005 ( .A(n2394), .Z(n2521) );
  ND2I U3006 ( .A(Addr[0]), .B(n2521), .Z(n2366) );
  AN2I U3007 ( .A(n2367), .B(n2366), .Z(n2369) );
  ND2I U3008 ( .A(n1206), .B(dx_gpr_rd_data1[0]), .Z(n2368) );
  ND2I U3009 ( .A(n2369), .B(n2368), .Z(n3194) );
  ND2I U3010 ( .A(n3118), .B(n3194), .Z(n2370) );
  AN2I U3011 ( .A(n2371), .B(n2370), .Z(n3141) );
  AN2I U3012 ( .A(n2921), .B(n2919), .Z(n2520) );
  IVI U3013 ( .A(n2520), .Z(n2783) );
  ND2I U3014 ( .A(Addr[2]), .B(n2514), .Z(n2374) );
  ND2I U3015 ( .A(n2372), .B(n2515), .Z(n2373) );
  AN2I U3016 ( .A(n2374), .B(n2373), .Z(n2376) );
  ND2I U3017 ( .A(n1201), .B(dx_gpr_rd_data1[2]), .Z(n2375) );
  ND2I U3018 ( .A(n2376), .B(n2375), .Z(n2963) );
  ND2I U3019 ( .A(n2793), .B(n2963), .Z(n2381) );
  ND2I U3020 ( .A(n2378), .B(n2377), .Z(n3357) );
  AN2I U3021 ( .A(n2379), .B(n3357), .Z(n2740) );
  IVI U3022 ( .A(n2740), .Z(n2809) );
  IVI U3023 ( .A(n2809), .Z(n4632) );
  ND2I U3024 ( .A(n4632), .B(n2966), .Z(n2380) );
  AN2I U3025 ( .A(n2381), .B(n2380), .Z(n3140) );
  ND2I U3026 ( .A(n3141), .B(n3140), .Z(n2836) );
  ND2I U3027 ( .A(n4461), .B(n2836), .Z(n2433) );
  IVI U3028 ( .A(n2382), .Z(n4637) );
  IVI U3029 ( .A(n3928), .Z(n4626) );
  ND2I U3030 ( .A(n2502), .B(n2501), .Z(n3031) );
  AN2I U3031 ( .A(n4626), .B(n1445), .Z(n4022) );
  AN2I U3032 ( .A(n4637), .B(n4022), .Z(n4549) );
  IVI U3033 ( .A(n1212), .Z(n2544) );
  ND2I U3034 ( .A(Addr[11]), .B(n2544), .Z(n2385) );
  IVI U3035 ( .A(n2383), .Z(n2395) );
  IVI U3036 ( .A(n2395), .Z(n2388) );
  IVI U3037 ( .A(n2388), .Z(n2545) );
  ND2I U3038 ( .A(n4683), .B(n2545), .Z(n2384) );
  AN2I U3039 ( .A(n2385), .B(n2384), .Z(n2387) );
  ND2I U3040 ( .A(n1200), .B(dx_gpr_rd_data1[11]), .Z(n2386) );
  ND2I U3041 ( .A(n2387), .B(n2386), .Z(n3012) );
  ND2I U3042 ( .A(n4403), .B(n1183), .Z(n2876) );
  IVI U3043 ( .A(n2783), .Z(n4630) );
  IVI U3044 ( .A(n2388), .Z(n2539) );
  ND2I U3045 ( .A(n2539), .B(n4682), .Z(n2393) );
  ND2I U3046 ( .A(n1203), .B(dx_gpr_rd_data1[10]), .Z(n2391) );
  ND2I U3047 ( .A(Addr[10]), .B(n2521), .Z(n2390) );
  AN2I U3048 ( .A(n2391), .B(n2390), .Z(n2392) );
  ND2I U3049 ( .A(n2393), .B(n2392), .Z(n4265) );
  ND2I U3050 ( .A(n4630), .B(n4265), .Z(n2893) );
  AN2I U3051 ( .A(n2876), .B(n2893), .Z(n2408) );
  ND2I U3052 ( .A(n1209), .B(dx_gpr_rd_data1[8]), .Z(n2400) );
  IVI U3053 ( .A(n1213), .Z(n2419) );
  ND2I U3054 ( .A(Addr[8]), .B(n2419), .Z(n2398) );
  ND2I U3055 ( .A(n2396), .B(n2395), .Z(n2397) );
  AN2I U3056 ( .A(n2398), .B(n2397), .Z(n2399) );
  ND2I U3057 ( .A(n2400), .B(n2399), .Z(n3156) );
  ND2I U3058 ( .A(n3013), .B(n3156), .Z(n2896) );
  ND2I U3059 ( .A(n2401), .B(n2545), .Z(n2405) );
  ND2I U3060 ( .A(n1200), .B(dx_gpr_rd_data1[9]), .Z(n2403) );
  ND2I U3061 ( .A(Addr[9]), .B(n2419), .Z(n2402) );
  AN2I U3062 ( .A(n2403), .B(n2402), .Z(n2404) );
  ND2I U3063 ( .A(n2405), .B(n2404), .Z(n3324) );
  ND2I U3064 ( .A(n4632), .B(n3324), .Z(n3126) );
  ND2I U3065 ( .A(n2896), .B(n3126), .Z(n2406) );
  IVI U3066 ( .A(n2406), .Z(n2407) );
  ND2I U3067 ( .A(n2408), .B(n2407), .Z(n4453) );
  ND2I U3068 ( .A(n1167), .B(n4453), .Z(n2430) );
  AN2I U3069 ( .A(n1170), .B(n2807), .Z(n4357) );
  ND2I U3070 ( .A(n3918), .B(n2533), .Z(n2410) );
  B4IP U3071 ( .A(n2410), .Z(n4412) );
  AN2I U3072 ( .A(n4357), .B(n4412), .Z(n4511) );
  IVI U3073 ( .A(n2520), .Z(n2728) );
  ND2I U3074 ( .A(Addr[14]), .B(n2419), .Z(n2412) );
  ND2I U3075 ( .A(n4684), .B(n2545), .Z(n2411) );
  AN2I U3076 ( .A(n2412), .B(n2411), .Z(n2414) );
  ND2I U3077 ( .A(n1201), .B(dx_gpr_rd_data1[14]), .Z(n2413) );
  ND2I U3078 ( .A(n2414), .B(n2413), .Z(n3035) );
  ND2I U3079 ( .A(n4591), .B(n3035), .Z(n2889) );
  IVI U3080 ( .A(n2725), .Z(n2761) );
  ND2I U3081 ( .A(Addr[13]), .B(n2419), .Z(n2417) );
  ND2I U3082 ( .A(n2415), .B(n2545), .Z(n2416) );
  ND2I U3083 ( .A(n2761), .B(n3781), .Z(n2875) );
  ND2I U3084 ( .A(n2545), .B(n2418), .Z(n2423) );
  ND2I U3085 ( .A(Addr[12]), .B(n2419), .Z(n2421) );
  ND2I U3086 ( .A(n1211), .B(dx_gpr_rd_data1[12]), .Z(n2420) );
  AN2I U3087 ( .A(n2421), .B(n2420), .Z(n2422) );
  ND2I U3088 ( .A(n2423), .B(n2422), .Z(n3813) );
  ND2I U3089 ( .A(n3118), .B(n3813), .Z(n2892) );
  IVI U3090 ( .A(n2503), .Z(n2762) );
  IVI U3091 ( .A(n2762), .Z(n2904) );
  ND2I U3092 ( .A(Addr[15]), .B(n2544), .Z(n2426) );
  ND2I U3093 ( .A(n2424), .B(n2545), .Z(n2425) );
  AN2I U3094 ( .A(n2426), .B(n2425), .Z(n2428) );
  ND2I U3095 ( .A(n1204), .B(dx_gpr_rd_data1[15]), .Z(n2427) );
  ND2I U3096 ( .A(n2428), .B(n2427), .Z(n3165) );
  ND2I U3097 ( .A(n2904), .B(n3165), .Z(n2879) );
  ND4P U3098 ( .A(n2889), .B(n2875), .C(n2892), .D(n2879), .Z(n4552) );
  ND2I U3099 ( .A(n4511), .B(n1173), .Z(n2429) );
  ND2I U3100 ( .A(n2430), .B(n2429), .Z(n2431) );
  IVI U3101 ( .A(n2431), .Z(n2432) );
  ND2I U3102 ( .A(n2433), .B(n2432), .Z(n2557) );
  IVI U3103 ( .A(n2707), .Z(n2492) );
  ND2I U3104 ( .A(n2492), .B(n2558), .Z(n2489) );
  OR2I U3105 ( .A(n3386), .B(n2489), .Z(n2436) );
  ND2I U3106 ( .A(n2435), .B(n2434), .Z(n2615) );
  NR2I U3107 ( .A(n2436), .B(n2615), .Z(n2438) );
  IVI U3108 ( .A(n2437), .Z(n3153) );
  AN2I U3109 ( .A(n2438), .B(n3153), .Z(n2439) );
  AN2I U3110 ( .A(n2440), .B(n2439), .Z(n2441) );
  ND2I U3111 ( .A(n1172), .B(n2441), .Z(n2841) );
  IVI U3112 ( .A(n2841), .Z(n2498) );
  IVI U3113 ( .A(n2443), .Z(n2844) );
  ND2I U3114 ( .A(n2444), .B(n1456), .Z(n2445) );
  NR2I U3115 ( .A(n2446), .B(n2445), .Z(n2447) );
  AN2I U3116 ( .A(n2448), .B(n2447), .Z(n2449) );
  ND2I U3117 ( .A(n2498), .B(n1439), .Z(n4445) );
  AN2I U3118 ( .A(n3871), .B(n2533), .Z(n4239) );
  IVI U3119 ( .A(n2503), .Z(n2729) );
  IVI U3120 ( .A(n2729), .Z(n2816) );
  ND2I U3121 ( .A(n2816), .B(n4086), .Z(n2550) );
  ND2I U3122 ( .A(Addr[21]), .B(n2544), .Z(n2452) );
  ND2I U3123 ( .A(n4687), .B(n2539), .Z(n2451) );
  AN2I U3124 ( .A(n2452), .B(n2451), .Z(n2454) );
  ND2I U3125 ( .A(n1206), .B(dx_gpr_rd_data1[21]), .Z(n2453) );
  ND2I U3126 ( .A(n2454), .B(n2453), .Z(n4227) );
  ND2I U3127 ( .A(n2761), .B(n4227), .Z(n4448) );
  ND2I U3128 ( .A(Addr[22]), .B(n2521), .Z(n2456) );
  ND2I U3129 ( .A(n4688), .B(n2539), .Z(n2455) );
  AN2I U3130 ( .A(n2456), .B(n2455), .Z(n2458) );
  ND2I U3131 ( .A(n1207), .B(dx_gpr_rd_data1[22]), .Z(n2457) );
  ND2I U3132 ( .A(n2458), .B(n2457), .Z(n4343) );
  ND2I U3133 ( .A(n3013), .B(n4343), .Z(n4116) );
  IVI U3134 ( .A(n2728), .Z(n2793) );
  ND2I U3135 ( .A(n2459), .B(n2539), .Z(n2463) );
  ND2I U3136 ( .A(Addr[20]), .B(n2544), .Z(n2461) );
  ND2I U3137 ( .A(n1210), .B(dx_gpr_rd_data1[20]), .Z(n2460) );
  AN2I U3138 ( .A(n2461), .B(n2460), .Z(n2462) );
  ND2I U3139 ( .A(n2463), .B(n2462), .Z(n4181) );
  ND2I U3140 ( .A(n2793), .B(n4181), .Z(n4112) );
  ND4P U3141 ( .A(n2550), .B(n4448), .C(n4116), .D(n4112), .Z(n3900) );
  ND2I U3142 ( .A(Addr[23]), .B(n2419), .Z(n2466) );
  ND2I U3143 ( .A(n2464), .B(n2526), .Z(n2465) );
  AN2I U3144 ( .A(n2466), .B(n2465), .Z(n2468) );
  ND2I U3145 ( .A(dx_gpr_rd_data1[23]), .B(n1208), .Z(n2467) );
  ND2I U3146 ( .A(n2468), .B(n2467), .Z(n4470) );
  ND2I U3147 ( .A(n2904), .B(n4470), .Z(n4446) );
  ND2I U3148 ( .A(Addr[25]), .B(n2419), .Z(n2470) );
  ND2I U3149 ( .A(n4689), .B(n2526), .Z(n2469) );
  AN2I U3150 ( .A(n2470), .B(n2469), .Z(n2472) );
  ND2I U3151 ( .A(dx_gpr_rd_data1[25]), .B(n1211), .Z(n2471) );
  ND2I U3152 ( .A(n2472), .B(n2471), .Z(n4385) );
  ND2I U3153 ( .A(n4402), .B(n4385), .Z(n4555) );
  ND2I U3154 ( .A(Addr[24]), .B(n2514), .Z(n2475) );
  ND2I U3155 ( .A(n2473), .B(n2526), .Z(n2474) );
  AN2I U3156 ( .A(n2475), .B(n2474), .Z(n2477) );
  ND2I U3157 ( .A(dx_gpr_rd_data1[24]), .B(n1203), .Z(n2476) );
  ND2I U3158 ( .A(n2477), .B(n2476), .Z(n4524) );
  ND2I U3159 ( .A(n2793), .B(n4524), .Z(n4117) );
  ND2I U3160 ( .A(Addr[26]), .B(n2521), .Z(n2480) );
  ND2I U3161 ( .A(n2478), .B(n2539), .Z(n2479) );
  AN2I U3162 ( .A(n2480), .B(n2479), .Z(n2482) );
  ND2I U3163 ( .A(n1210), .B(dx_gpr_rd_data1[26]), .Z(n2481) );
  ND2I U3164 ( .A(n2482), .B(n2481), .Z(n4303) );
  AO2 U3165 ( .A(n4239), .B(n3900), .C(n4412), .D(n3874), .Z(n3123) );
  NR2I U3166 ( .A(n4056), .B(n2483), .Z(n2488) );
  ND2I U3167 ( .A(dx_gpr_rd_data2[19]), .B(n2700), .Z(n2484) );
  ND2I U3168 ( .A(n2485), .B(n2484), .Z(n2486) );
  IVI U3169 ( .A(n2486), .Z(n2487) );
  ND2I U3170 ( .A(n2488), .B(n2487), .Z(n3277) );
  IVI U3171 ( .A(n2558), .Z(n2491) );
  IVI U3172 ( .A(n2489), .Z(n2490) );
  ND2I U3173 ( .A(n2490), .B(n3386), .Z(n3022) );
  IVI U3174 ( .A(n3022), .Z(n4314) );
  ND2I U3175 ( .A(n2706), .B(n2492), .Z(n2909) );
  IVI U3176 ( .A(n2909), .Z(n4313) );
  MUX21L U3177 ( .A(n4314), .B(n4313), .S(n4086), .Z(n2493) );
  ND2I U3178 ( .A(n4642), .B(n2493), .Z(n2494) );
  ND2I U3179 ( .A(n3277), .B(n2494), .Z(n2497) );
  IVI U3180 ( .A(n3022), .Z(n4496) );
  IVI U3181 ( .A(n4496), .Z(n4020) );
  AO7 U3182 ( .A(n3277), .B(n4020), .C(n4643), .Z(n2495) );
  ND2I U3183 ( .A(n4086), .B(n2495), .Z(n2496) );
  AN2I U3184 ( .A(n2497), .B(n2496), .Z(n2508) );
  ND2I U3185 ( .A(n2498), .B(n1439), .Z(n2871) );
  IVI U3186 ( .A(n2871), .Z(n3098) );
  IVI U3187 ( .A(n2729), .Z(n2942) );
  ND2I U3188 ( .A(n2942), .B(n4565), .Z(n4556) );
  IVI U3189 ( .A(n2520), .Z(n2736) );
  ND2I U3190 ( .A(n2923), .B(n4424), .Z(n2864) );
  ND2I U3191 ( .A(n4632), .B(n4601), .Z(n2863) );
  ND2I U3192 ( .A(n3013), .B(n4653), .Z(n2862) );
  ND4P U3193 ( .A(n4556), .B(n2864), .C(n2863), .D(n2862), .Z(n3870) );
  ND2I U3194 ( .A(n1445), .B(n3870), .Z(n2506) );
  ND2I U3195 ( .A(n2502), .B(n2501), .Z(n3362) );
  ND2I U3196 ( .A(n3918), .B(n3362), .Z(n4619) );
  IVI U3197 ( .A(n2503), .Z(n2720) );
  IVI U3198 ( .A(n2720), .Z(n4403) );
  AN2I U3199 ( .A(n4403), .B(n4650), .Z(n4540) );
  ND2I U3200 ( .A(n4502), .B(n4540), .Z(n2505) );
  ND2I U3201 ( .A(n2506), .B(n2505), .Z(n3121) );
  ND2I U3202 ( .A(n3098), .B(n3121), .Z(n2507) );
  AO3 U3203 ( .A(n4445), .B(n3123), .C(n2508), .D(n2507), .Z(n2509) );
  IVI U3204 ( .A(n2509), .Z(n2555) );
  AN2I U3205 ( .A(n1170), .B(n2807), .Z(n4504) );
  IVI U3206 ( .A(n4619), .Z(n4502) );
  AN2I U3207 ( .A(n4504), .B(n4502), .Z(n4553) );
  IVI U3208 ( .A(n2740), .Z(n2730) );
  IVI U3209 ( .A(n2730), .Z(n3007) );
  ND2I U3210 ( .A(Addr[5]), .B(n2514), .Z(n2511) );
  ND2I U3211 ( .A(n4679), .B(n2515), .Z(n2510) );
  AN2I U3212 ( .A(n2511), .B(n2510), .Z(n2513) );
  ND2I U3213 ( .A(n1207), .B(dx_gpr_rd_data1[5]), .Z(n2512) );
  ND2I U3214 ( .A(n2513), .B(n2512), .Z(n3008) );
  ND2I U3215 ( .A(n3007), .B(n3008), .Z(n2532) );
  ND2I U3216 ( .A(Addr[4]), .B(n2514), .Z(n2517) );
  ND2I U3217 ( .A(n4678), .B(n2515), .Z(n2516) );
  AN2I U3218 ( .A(n2517), .B(n2516), .Z(n2519) );
  ND2I U3219 ( .A(n1204), .B(dx_gpr_rd_data1[4]), .Z(n2518) );
  ND2I U3220 ( .A(n2519), .B(n2518), .Z(n3929) );
  ND2I U3221 ( .A(n3118), .B(n3929), .Z(n2531) );
  IVI U3222 ( .A(n2520), .Z(n2756) );
  ND2I U3223 ( .A(Addr[6]), .B(n2521), .Z(n2523) );
  ND2I U3224 ( .A(n4680), .B(n2539), .Z(n2522) );
  AN2I U3225 ( .A(n2523), .B(n2522), .Z(n2525) );
  ND2I U3226 ( .A(n1205), .B(dx_gpr_rd_data1[6]), .Z(n2524) );
  ND2I U3227 ( .A(n2525), .B(n2524), .Z(n3886) );
  ND2I U3228 ( .A(n2796), .B(n1187), .Z(n2897) );
  IVI U3229 ( .A(n2762), .Z(n3186) );
  ND2I U3230 ( .A(dx_gpr_rd_data1[7]), .B(n1209), .Z(n2528) );
  ND2I U3231 ( .A(n4681), .B(n2526), .Z(n2527) );
  AN2I U3232 ( .A(n2528), .B(n2527), .Z(n2530) );
  ND2I U3233 ( .A(n2521), .B(Addr[7]), .Z(n2529) );
  ND2I U3234 ( .A(n2530), .B(n2529), .Z(n3883) );
  ND2I U3235 ( .A(n3186), .B(n3883), .Z(n3127) );
  ND4P U3236 ( .A(n2532), .B(n2531), .C(n2897), .D(n3127), .Z(n4460) );
  ND2I U3237 ( .A(n4553), .B(n1164), .Z(n2552) );
  AN2I U3238 ( .A(n3871), .B(n2533), .Z(n4356) );
  AN2I U3239 ( .A(n4356), .B(n4357), .Z(n4452) );
  ND2I U3240 ( .A(n1209), .B(dx_gpr_rd_data1[16]), .Z(n2538) );
  ND2I U3241 ( .A(Addr[16]), .B(n2544), .Z(n2536) );
  ND2I U3242 ( .A(n2534), .B(n2539), .Z(n2535) );
  AN2I U3243 ( .A(n2536), .B(n2535), .Z(n2537) );
  ND2I U3244 ( .A(n2538), .B(n2537), .Z(n2947) );
  ND2I U3245 ( .A(n3013), .B(n2947), .Z(n2888) );
  IVI U3246 ( .A(n2740), .Z(n2725) );
  IVI U3247 ( .A(n2725), .Z(n2802) );
  ND2I U3248 ( .A(Addr[17]), .B(n2544), .Z(n2541) );
  ND2I U3249 ( .A(n4685), .B(n2539), .Z(n2540) );
  AN2I U3250 ( .A(n2541), .B(n2540), .Z(n2543) );
  ND2I U3251 ( .A(n1207), .B(dx_gpr_rd_data1[17]), .Z(n2542) );
  ND2I U3252 ( .A(n2543), .B(n2542), .Z(n2945) );
  ND2I U3253 ( .A(n2802), .B(n2945), .Z(n2878) );
  IVI U3254 ( .A(n2736), .Z(n4400) );
  ND2I U3255 ( .A(Addr[18]), .B(n2544), .Z(n2547) );
  ND2I U3256 ( .A(n4686), .B(n2545), .Z(n2546) );
  AN2I U3257 ( .A(n2547), .B(n2546), .Z(n2549) );
  ND2I U3258 ( .A(n1201), .B(dx_gpr_rd_data1[18]), .Z(n2548) );
  ND2I U3259 ( .A(n2549), .B(n2548), .Z(n4037) );
  ND2I U3260 ( .A(n4400), .B(n4037), .Z(n2741) );
  ND4 U3261 ( .A(n2888), .B(n2878), .C(n2741), .D(n2550), .Z(n4618) );
  ND2I U3262 ( .A(n4452), .B(n4618), .Z(n2551) );
  ND2I U3263 ( .A(n2552), .B(n2551), .Z(n2553) );
  IVI U3264 ( .A(n2553), .Z(n2554) );
  ND2I U3265 ( .A(n2555), .B(n2554), .Z(n2556) );
  NR2I U3266 ( .A(n2557), .B(n2556), .Z(n2719) );
  AN2I U3267 ( .A(n2707), .B(n2558), .Z(n3384) );
  ND2I U3268 ( .A(n3384), .B(n3386), .Z(n2708) );
  IVI U3269 ( .A(n2708), .Z(n2633) );
  IVI U3270 ( .A(n2633), .Z(n2669) );
  IVI U3271 ( .A(n1436), .Z(n2559) );
  ENI U3272 ( .A(n2560), .B(n2559), .Z(n3065) );
  IVI U3273 ( .A(n3065), .Z(n2561) );
  IVI U3274 ( .A(n3165), .Z(n3310) );
  AN2I U3275 ( .A(n2561), .B(n3310), .Z(n2564) );
  ND2I U3276 ( .A(n3065), .B(n3165), .Z(n2562) );
  IVI U3277 ( .A(n1436), .Z(n4183) );
  ENI U3278 ( .A(n3024), .B(n4183), .Z(n3036) );
  ND2I U3279 ( .A(n3036), .B(n3035), .Z(n3066) );
  MUX21L U3280 ( .A(n2564), .B(n2562), .S(n3066), .Z(n2578) );
  IVI U3281 ( .A(n3036), .Z(n2563) );
  IVI U3282 ( .A(n3035), .Z(n3308) );
  ND2I U3283 ( .A(n2563), .B(n3308), .Z(n3067) );
  IVI U3284 ( .A(n2564), .Z(n2565) );
  ND2I U3285 ( .A(n3067), .B(n2565), .Z(n2566) );
  ND2I U3286 ( .A(n2562), .B(n2566), .Z(n2577) );
  IVI U3287 ( .A(n1436), .Z(n2568) );
  ENI U3288 ( .A(n3302), .B(n2568), .Z(n3782) );
  ND2I U3289 ( .A(n3782), .B(n3781), .Z(n2567) );
  ENI U3290 ( .A(n2569), .B(n2568), .Z(n3814) );
  ND2I U3291 ( .A(n3813), .B(n3814), .Z(n3783) );
  IVI U3292 ( .A(n3783), .Z(n2572) );
  IVI U3293 ( .A(n3782), .Z(n2571) );
  IVI U3294 ( .A(n3781), .Z(n2570) );
  ND2I U3295 ( .A(n2571), .B(n2570), .Z(n2575) );
  ND2I U3296 ( .A(n2572), .B(n2575), .Z(n2573) );
  ND2I U3297 ( .A(n2567), .B(n2573), .Z(n3069) );
  MUX21LP U3298 ( .A(n2578), .B(n2577), .S(n3069), .Z(n2610) );
  IVI U3299 ( .A(n3813), .Z(n3317) );
  IVI U3300 ( .A(n3814), .Z(n2574) );
  ND2I U3301 ( .A(n3317), .B(n2574), .Z(n3784) );
  ND2I U3302 ( .A(n2575), .B(n3784), .Z(n2576) );
  ND2I U3303 ( .A(n2567), .B(n2576), .Z(n3070) );
  MUX21LP U3304 ( .A(n2578), .B(n2577), .S(n3070), .Z(n2609) );
  IVI U3305 ( .A(n1436), .Z(n2663) );
  ENI U3306 ( .A(n2855), .B(n1436), .Z(n2579) );
  IVI U3307 ( .A(n2579), .Z(n2826) );
  ND2I U3308 ( .A(n2826), .B(n1183), .Z(n2594) );
  IVI U3309 ( .A(n3012), .Z(n3332) );
  AN2I U3310 ( .A(n3332), .B(n2579), .Z(n2595) );
  ENI U3311 ( .A(n3322), .B(n1436), .Z(n2593) );
  IVI U3312 ( .A(n4265), .Z(n2580) );
  ND2I U3313 ( .A(n2593), .B(n2580), .Z(n2828) );
  IVI U3314 ( .A(n2633), .Z(n2628) );
  ENI U3315 ( .A(n3088), .B(n2628), .Z(n3100) );
  ND2I U3316 ( .A(n3100), .B(n3324), .Z(n2602) );
  IVI U3317 ( .A(n3156), .Z(n3341) );
  AN2I U3318 ( .A(n2582), .B(n2581), .Z(n2587) );
  ND2I U3319 ( .A(n2584), .B(n2583), .Z(n2585) );
  IVI U3320 ( .A(n2585), .Z(n2586) );
  ND2I U3321 ( .A(n2587), .B(n2586), .Z(n2599) );
  ENI U3322 ( .A(n2599), .B(n1436), .Z(n3171) );
  ND2I U3323 ( .A(n3341), .B(n3171), .Z(n3099) );
  IVI U3324 ( .A(n3099), .Z(n2588) );
  ND2I U3325 ( .A(n2602), .B(n2588), .Z(n2591) );
  NR2I U3326 ( .A(n3100), .B(n3324), .Z(n2589) );
  ND2I U3327 ( .A(n2591), .B(n2590), .Z(n2592) );
  IVI U3328 ( .A(n2592), .Z(n2830) );
  ND2I U3329 ( .A(n2606), .B(n2830), .Z(n2596) );
  IVI U3330 ( .A(n2593), .Z(n4266) );
  ND2I U3331 ( .A(n4266), .B(n1180), .Z(n2827) );
  ND2I U3332 ( .A(n2596), .B(n2607), .Z(n3040) );
  ND2I U3333 ( .A(n2598), .B(n2597), .Z(n2604) );
  ENI U3334 ( .A(n2599), .B(n1436), .Z(n2600) );
  IVI U3335 ( .A(n2600), .Z(n2601) );
  ND2I U3336 ( .A(n2601), .B(n3156), .Z(n3104) );
  ND2I U3337 ( .A(n2602), .B(n3104), .Z(n2603) );
  ND2I U3338 ( .A(n2604), .B(n2603), .Z(n2851) );
  IVI U3339 ( .A(n2851), .Z(n2605) );
  ND2I U3340 ( .A(n2606), .B(n2605), .Z(n2608) );
  ND2I U3341 ( .A(n2608), .B(n2607), .Z(n3041) );
  ND2I U3342 ( .A(n2612), .B(n2611), .Z(n2613) );
  ENI U3343 ( .A(n2613), .B(n2628), .Z(n3884) );
  ND2I U3344 ( .A(n3884), .B(n3883), .Z(n2614) );
  ENI U3345 ( .A(n2615), .B(n2628), .Z(n3887) );
  ND2I U3346 ( .A(n3887), .B(n3886), .Z(n3885) );
  IVI U3347 ( .A(n3885), .Z(n2616) );
  OR2P U3348 ( .A(n3884), .B(n3883), .Z(n2620) );
  ND2I U3349 ( .A(n2616), .B(n2620), .Z(n2617) );
  ND2I U3350 ( .A(n2614), .B(n2617), .Z(n2640) );
  IVI U3351 ( .A(n3886), .Z(n2619) );
  IVI U3352 ( .A(n3887), .Z(n2618) );
  ND2I U3353 ( .A(n2619), .B(n2618), .Z(n2621) );
  ND2I U3354 ( .A(n2621), .B(n2620), .Z(n2622) );
  ND2I U3355 ( .A(n2614), .B(n2622), .Z(n2641) );
  IVI U3356 ( .A(n3929), .Z(n3371) );
  ND2I U3357 ( .A(n2624), .B(n2623), .Z(n2625) );
  IVI U3358 ( .A(n2625), .Z(n2626) );
  ND2I U3359 ( .A(n2627), .B(n2626), .Z(n2629) );
  ENI U3360 ( .A(n2629), .B(n2628), .Z(n3930) );
  IVI U3361 ( .A(n3930), .Z(n2630) );
  ND2I U3362 ( .A(n3371), .B(n2630), .Z(n3000) );
  IVI U3363 ( .A(n3008), .Z(n3350) );
  ND2I U3364 ( .A(n2632), .B(n1168), .Z(n2635) );
  IVI U3365 ( .A(n2633), .Z(n2654) );
  IVI U3366 ( .A(n2654), .Z(n2647) );
  ENI U3367 ( .A(n2635), .B(n2647), .Z(n2634) );
  ND2I U3368 ( .A(n3350), .B(n2634), .Z(n2638) );
  ND2I U3369 ( .A(n3000), .B(n2638), .Z(n2636) );
  ENI U3370 ( .A(n2635), .B(n2654), .Z(n2998) );
  ND2I U3371 ( .A(n3008), .B(n2998), .Z(n2637) );
  ND2I U3372 ( .A(n2636), .B(n2637), .Z(n3840) );
  ND2I U3373 ( .A(n3930), .B(n3929), .Z(n2999) );
  ND2I U3374 ( .A(n2999), .B(n2637), .Z(n2639) );
  ND2I U3375 ( .A(n2639), .B(n2638), .Z(n3891) );
  ND2I U3376 ( .A(n2647), .B(n2649), .Z(n2643) );
  NR2I U3377 ( .A(n2643), .B(n2642), .Z(n2644) );
  ND2I U3378 ( .A(n2646), .B(n2644), .Z(n2659) );
  IVI U3379 ( .A(n3136), .Z(n2645) );
  ND2I U3380 ( .A(n2659), .B(n2645), .Z(n2657) );
  IVI U3381 ( .A(n2646), .Z(n2648) );
  ND2I U3382 ( .A(n2648), .B(n2628), .Z(n2662) );
  ND2I U3383 ( .A(n2650), .B(n2649), .Z(n2651) );
  IVI U3384 ( .A(n2651), .Z(n2652) );
  ND2I U3385 ( .A(n2653), .B(n2652), .Z(n2655) );
  ND2I U3386 ( .A(n2655), .B(n2654), .Z(n2658) );
  ND2I U3387 ( .A(n2662), .B(n2658), .Z(n2656) );
  NR2I U3388 ( .A(n2657), .B(n2656), .Z(n2680) );
  IVI U3389 ( .A(n2680), .Z(n2665) );
  ND2I U3390 ( .A(n2659), .B(n2658), .Z(n2660) );
  IVI U3391 ( .A(n2660), .Z(n2661) );
  ND2I U3392 ( .A(n2662), .B(n2661), .Z(n3137) );
  AN2I U3393 ( .A(n3137), .B(n3136), .Z(n2678) );
  ENI U3394 ( .A(n2664), .B(n2663), .Z(n2960) );
  ND2I U3395 ( .A(n2963), .B(n2960), .Z(n3138) );
  MUX21L U3396 ( .A(n2665), .B(n2678), .S(n3138), .Z(n2676) );
  ENI U3397 ( .A(n3357), .B(n2628), .Z(n2907) );
  ND2I U3398 ( .A(n2907), .B(n2966), .Z(n2674) );
  ND2I U3399 ( .A(n3194), .B(n1436), .Z(n2670) );
  ND2I U3400 ( .A(n3189), .B(n2670), .Z(n2673) );
  NR2I U3401 ( .A(n3194), .B(n1436), .Z(n2671) );
  ND2I U3402 ( .A(n2673), .B(n2672), .Z(n2906) );
  ND2I U3403 ( .A(n2674), .B(n2906), .Z(n2675) );
  ND2I U3404 ( .A(n2675), .B(n1438), .Z(n2958) );
  ND2I U3405 ( .A(n2676), .B(n2958), .Z(n3001) );
  IVI U3406 ( .A(n2960), .Z(n2677) );
  IVI U3407 ( .A(n2963), .Z(n3364) );
  IVI U3408 ( .A(n2678), .Z(n2679) );
  ND2I U3409 ( .A(n1440), .B(n2679), .Z(n2682) );
  ND2I U3410 ( .A(n3001), .B(n1437), .Z(n3895) );
  ND2I U3411 ( .A(n2683), .B(n3895), .Z(n2833) );
  ND2I U3412 ( .A(n2684), .B(n2833), .Z(n2685) );
  MUX21LP U3413 ( .A(n2687), .B(n2686), .S(n2685), .Z(n4483) );
  IVI U3414 ( .A(n1436), .Z(n4177) );
  ENI U3415 ( .A(n3277), .B(n4177), .Z(n4087) );
  ENI U3416 ( .A(n4087), .B(n4086), .Z(n2691) );
  IVI U3417 ( .A(n2688), .Z(n2689) );
  ND2I U3418 ( .A(dx_gpr_rd_data2[18]), .B(n3248), .Z(n3269) );
  ND2I U3419 ( .A(n2689), .B(n3269), .Z(n4021) );
  IVI U3420 ( .A(n1436), .Z(n2698) );
  ENI U3421 ( .A(n4021), .B(n2698), .Z(n2690) );
  ND2I U3422 ( .A(n2690), .B(n4037), .Z(n4094) );
  EOI U3423 ( .A(n2691), .B(n4094), .Z(n2714) );
  ENI U3424 ( .A(n4021), .B(n4153), .Z(n4036) );
  IVI U3425 ( .A(n4037), .Z(n3276) );
  ND2I U3426 ( .A(n4036), .B(n3276), .Z(n4090) );
  IVI U3427 ( .A(n2692), .Z(n2693) );
  NR2I U3428 ( .A(n4056), .B(n2693), .Z(n2697) );
  ND2I U3429 ( .A(n3254), .B(dx_gpr_rd_data2[17]), .Z(n2694) );
  AN2I U3430 ( .A(n2695), .B(n2694), .Z(n2696) );
  ND2I U3431 ( .A(n2697), .B(n2696), .Z(n2724) );
  ENI U3432 ( .A(n2724), .B(n2698), .Z(n2771) );
  ND2I U3433 ( .A(n2771), .B(n2945), .Z(n2709) );
  IVI U3434 ( .A(n2771), .Z(n2699) );
  IVI U3435 ( .A(n2945), .Z(n3272) );
  ND2I U3436 ( .A(n2699), .B(n3272), .Z(n2711) );
  ND2I U3437 ( .A(dx_gpr_rd_data2[16]), .B(n3254), .Z(n2703) );
  IVI U3438 ( .A(n2701), .Z(n2702) );
  ND2I U3439 ( .A(n2703), .B(n2702), .Z(n2786) );
  ENI U3440 ( .A(n2786), .B(n4141), .Z(n2779) );
  IVI U3441 ( .A(n2779), .Z(n2704) );
  IVI U3442 ( .A(n2947), .Z(n3292) );
  ND2I U3443 ( .A(n2704), .B(n3292), .Z(n2770) );
  ND2I U3444 ( .A(n2711), .B(n2770), .Z(n2705) );
  ND2I U3445 ( .A(n2709), .B(n2705), .Z(n4092) );
  MUX21H U3446 ( .A(n2714), .B(n2713), .S(n4092), .Z(n2717) );
  ND2I U3447 ( .A(n2779), .B(n2947), .Z(n2772) );
  IVI U3448 ( .A(n2772), .Z(n2710) );
  ND2I U3449 ( .A(n2711), .B(n2710), .Z(n2712) );
  ND2I U3450 ( .A(n2709), .B(n2712), .Z(n4099) );
  MUX21L U3451 ( .A(n2714), .B(n2713), .S(n4099), .Z(n2715) );
  ND2I U3452 ( .A(n4669), .B(n2715), .Z(n2716) );
  AO3 U3453 ( .A(n4669), .B(n2717), .C(n4041), .D(n2716), .Z(n2718) );
  ND2I U3454 ( .A(n2719), .B(n2718), .Z(x_ALU_Result[19]) );
  ND2I U3455 ( .A(n4400), .B(n3929), .Z(n2723) );
  IVI U3456 ( .A(n2725), .Z(n4402) );
  ND2I U3457 ( .A(n4402), .B(n3136), .Z(n2722) );
  IVI U3458 ( .A(n2720), .Z(n2936) );
  ND2I U3459 ( .A(n2936), .B(n3008), .Z(n2894) );
  ND2I U3460 ( .A(n3013), .B(n2963), .Z(n2721) );
  ND4P U3461 ( .A(n2723), .B(n2722), .C(n2894), .D(n2721), .Z(n4220) );
  ND2I U3462 ( .A(n4553), .B(n1166), .Z(n2751) );
  B2I U3463 ( .A(n2724), .Z2(n3271) );
  ND2I U3464 ( .A(n2745), .B(n4445), .Z(n2749) );
  IVI U3465 ( .A(n2725), .Z(n3117) );
  ND2I U3466 ( .A(n3117), .B(n4565), .Z(n2727) );
  ND2I U3467 ( .A(n3013), .B(n4424), .Z(n2726) );
  AN2I U3468 ( .A(n2727), .B(n2726), .Z(n2983) );
  IVI U3469 ( .A(n2728), .Z(n2796) );
  ND2I U3470 ( .A(n2796), .B(n4303), .Z(n4557) );
  ND2I U3471 ( .A(n2922), .B(n4385), .Z(n4119) );
  AN2I U3472 ( .A(n4557), .B(n4119), .Z(n2982) );
  ND2I U3473 ( .A(n2983), .B(n2982), .Z(n4372) );
  ND2I U3474 ( .A(n4372), .B(n1445), .Z(n2734) );
  IVI U3475 ( .A(n2730), .Z(n2948) );
  ND2I U3476 ( .A(n2948), .B(n4650), .Z(n2732) );
  ND2I U3477 ( .A(n4403), .B(n4601), .Z(n2731) );
  AN2I U3478 ( .A(n2732), .B(n2731), .Z(n2979) );
  ND2I U3479 ( .A(n4400), .B(n4653), .Z(n2978) );
  ND2I U3480 ( .A(n2979), .B(n2978), .Z(n4353) );
  IVI U3481 ( .A(n4619), .Z(n4583) );
  ND2I U3482 ( .A(n4353), .B(n4583), .Z(n2733) );
  AN2I U3483 ( .A(n2734), .B(n2733), .Z(n2885) );
  IVI U3484 ( .A(n2809), .Z(n2951) );
  ND2I U3485 ( .A(n2951), .B(n4470), .Z(n4118) );
  ND2I U3486 ( .A(n2904), .B(n4227), .Z(n4111) );
  ND2I U3487 ( .A(n4118), .B(n4111), .Z(n2735) );
  IVI U3488 ( .A(n2735), .Z(n2739) );
  IVI U3489 ( .A(n2736), .Z(n2923) );
  ND2I U3490 ( .A(n2923), .B(n4343), .Z(n4447) );
  ND2I U3491 ( .A(n3013), .B(n4524), .Z(n4554) );
  ND2I U3492 ( .A(n4447), .B(n4554), .Z(n2737) );
  IVI U3493 ( .A(n2737), .Z(n2738) );
  AN2I U3494 ( .A(n2739), .B(n2738), .Z(n2976) );
  IVI U3495 ( .A(n2976), .Z(n3777) );
  ND2I U3496 ( .A(n3777), .B(n4412), .Z(n2743) );
  ND2I U3497 ( .A(n3013), .B(n4181), .Z(n4449) );
  ND2I U3498 ( .A(n2936), .B(n2945), .Z(n2757) );
  ND2I U3499 ( .A(n3007), .B(n4086), .Z(n4113) );
  ND4P U3500 ( .A(n2741), .B(n4449), .C(n2757), .D(n4113), .Z(n3780) );
  ND2I U3501 ( .A(n3780), .B(n4356), .Z(n2742) );
  ND2I U3502 ( .A(n2743), .B(n2742), .Z(n2744) );
  IVI U3503 ( .A(n2744), .Z(n2884) );
  ND2I U3504 ( .A(n2745), .B(n2884), .Z(n2746) );
  IVI U3505 ( .A(n2746), .Z(n2747) );
  ND2I U3506 ( .A(n2885), .B(n2747), .Z(n2748) );
  ND2I U3507 ( .A(n2749), .B(n2748), .Z(n2750) );
  ND2I U3508 ( .A(n2751), .B(n2750), .Z(n2769) );
  AN2I U3509 ( .A(n2752), .B(n4029), .Z(n4532) );
  ND2I U3510 ( .A(n2816), .B(n2966), .Z(n2754) );
  IVI U3511 ( .A(n2756), .Z(n4124) );
  ND2I U3512 ( .A(n4124), .B(n3194), .Z(n2753) );
  AN2I U3513 ( .A(n2754), .B(n2753), .Z(n4202) );
  IVI U3514 ( .A(n4202), .Z(n3765) );
  AN2I U3515 ( .A(n3856), .B(n3765), .Z(n2755) );
  ND2I U3516 ( .A(n4532), .B(n2755), .Z(n2759) );
  AN2I U3517 ( .A(n4504), .B(n4356), .Z(n4558) );
  ND2I U3518 ( .A(n4402), .B(n3165), .Z(n2886) );
  ND2I U3519 ( .A(n3013), .B(n3035), .Z(n2873) );
  IVI U3520 ( .A(n2756), .Z(n2929) );
  ND2I U3521 ( .A(n2929), .B(n2947), .Z(n2877) );
  ND4 U3522 ( .A(n2757), .B(n2886), .C(n2873), .D(n2877), .Z(n4377) );
  ND2I U3523 ( .A(n4558), .B(n4377), .Z(n2758) );
  AN2I U3524 ( .A(n2759), .B(n2758), .Z(n2767) );
  ND2I U3525 ( .A(n2802), .B(n3883), .Z(n2895) );
  ND2I U3526 ( .A(n3013), .B(n1186), .Z(n2760) );
  ND2I U3527 ( .A(n2796), .B(n3156), .Z(n3125) );
  ND2I U3528 ( .A(n2942), .B(n3324), .Z(n2891) );
  ND4P U3529 ( .A(n2895), .B(n2760), .C(n3125), .D(n2891), .Z(n3764) );
  ND2I U3530 ( .A(n4549), .B(n3764), .Z(n2764) );
  ND2I U3531 ( .A(n2761), .B(n1182), .Z(n2890) );
  ND2I U3532 ( .A(n2923), .B(n3813), .Z(n2874) );
  IVI U3533 ( .A(n2762), .Z(n4126) );
  ND2I U3534 ( .A(n4126), .B(n3781), .Z(n2887) );
  ND2I U3535 ( .A(n3118), .B(n1181), .Z(n3124) );
  ND4P U3536 ( .A(n2890), .B(n2874), .C(n2887), .D(n3124), .Z(n4374) );
  ND2I U3537 ( .A(n4374), .B(n4511), .Z(n2763) );
  ND2I U3538 ( .A(n2764), .B(n2763), .Z(n2765) );
  IVI U3539 ( .A(n2765), .Z(n2766) );
  ND2I U3540 ( .A(n2767), .B(n2766), .Z(n2768) );
  NR2I U3541 ( .A(n2769), .B(n2768), .Z(n2778) );
  ENI U3542 ( .A(n2771), .B(n2945), .Z(n2773) );
  ENI U3543 ( .A(n2773), .B(n2772), .Z(n2774) );
  ND2I U3544 ( .A(n2774), .B(n4576), .Z(n2775) );
  ND2I U3545 ( .A(n2778), .B(n2777), .Z(x_ALU_Result[17]) );
  ENI U3546 ( .A(n2779), .B(n2947), .Z(n2780) );
  ENI U3547 ( .A(n4484), .B(n2780), .Z(n2782) );
  ND2I U3548 ( .A(n2782), .B(n4672), .Z(n2825) );
  ND2I U3549 ( .A(n3007), .B(n1186), .Z(n3179) );
  ND2I U3550 ( .A(n3118), .B(n3008), .Z(n2784) );
  IVI U3551 ( .A(n2783), .Z(n4591) );
  ND2I U3552 ( .A(n4591), .B(n3883), .Z(n2944) );
  ND2I U3553 ( .A(n2922), .B(n3156), .Z(n3168) );
  ND4P U3554 ( .A(n3179), .B(n2784), .C(n2944), .D(n3168), .Z(n3796) );
  ND2I U3555 ( .A(n4549), .B(n1158), .Z(n2792) );
  MUX21L U3556 ( .A(n4314), .B(n4313), .S(n2947), .Z(n2785) );
  ND2I U3557 ( .A(n4642), .B(n2785), .Z(n2787) );
  IVDA U3558 ( .A(n2786), .Z(n3291) );
  ND2I U3559 ( .A(n2787), .B(n3291), .Z(n2790) );
  AO7 U3560 ( .A(n4317), .B(n3291), .C(n4642), .Z(n2788) );
  ND2I U3561 ( .A(n2947), .B(n2788), .Z(n2789) );
  AN2I U3562 ( .A(n2790), .B(n2789), .Z(n2791) );
  AN2I U3563 ( .A(n2792), .B(n2791), .Z(n2806) );
  IVI U3564 ( .A(n2871), .Z(n4293) );
  AO2 U3565 ( .A(n3013), .B(n4650), .C(n2816), .D(n4424), .Z(n2795) );
  AO2 U3566 ( .A(n2951), .B(n4653), .C(n2793), .D(n4601), .Z(n2794) );
  AN2I U3567 ( .A(n2795), .B(n2794), .Z(n3919) );
  IVI U3568 ( .A(n3919), .Z(n4512) );
  ND2I U3569 ( .A(n2796), .B(n4385), .Z(n4280) );
  ND2I U3570 ( .A(n4126), .B(n4524), .Z(n4408) );
  AN2I U3571 ( .A(n4280), .B(n4408), .Z(n2800) );
  ND2I U3572 ( .A(n2948), .B(n4303), .Z(n2798) );
  ND2I U3573 ( .A(n3013), .B(n4565), .Z(n2797) );
  AN2I U3574 ( .A(n2798), .B(n2797), .Z(n2799) );
  ND2I U3575 ( .A(n2800), .B(n2799), .Z(n4517) );
  ND2I U3576 ( .A(n4126), .B(n4181), .Z(n4074) );
  ND2I U3577 ( .A(n4632), .B(n4343), .Z(n4407) );
  ND2I U3578 ( .A(n4074), .B(n4407), .Z(n2801) );
  IVI U3579 ( .A(n2801), .Z(n3923) );
  ND2I U3580 ( .A(n3013), .B(n4470), .Z(n4277) );
  ND2I U3581 ( .A(n2923), .B(n4227), .Z(n4297) );
  ND2I U3582 ( .A(n3923), .B(n3921), .Z(n3810) );
  ND2I U3583 ( .A(n4412), .B(n3810), .Z(n2804) );
  ND2I U3584 ( .A(n2929), .B(n2945), .Z(n4016) );
  ND2I U3585 ( .A(n3013), .B(n4086), .Z(n4300) );
  ND2I U3586 ( .A(n2936), .B(n2947), .Z(n2815) );
  ND2I U3587 ( .A(n2802), .B(n4037), .Z(n4075) );
  ND4 U3588 ( .A(n4016), .B(n4300), .C(n2815), .D(n4075), .Z(n3927) );
  ND2I U3589 ( .A(n4356), .B(n3927), .Z(n2803) );
  ND2I U3590 ( .A(n4293), .B(n3185), .Z(n2805) );
  ND2I U3591 ( .A(n2806), .B(n2805), .Z(n2823) );
  AN2I U3592 ( .A(n2807), .B(n4412), .Z(n2808) );
  AN2I U3593 ( .A(n1170), .B(n2808), .Z(n4542) );
  ND2I U3594 ( .A(n2951), .B(n1181), .Z(n3167) );
  ND2I U3595 ( .A(n2923), .B(n1182), .Z(n2950) );
  ND2I U3596 ( .A(n2936), .B(n3813), .Z(n3164) );
  ND2I U3597 ( .A(n3013), .B(n3324), .Z(n2943) );
  ND4P U3598 ( .A(n3167), .B(n2950), .C(n3164), .D(n2943), .Z(n4501) );
  ND2I U3599 ( .A(n4542), .B(n4501), .Z(n2814) );
  ND2I U3600 ( .A(n2793), .B(n3136), .Z(n2812) );
  IVI U3601 ( .A(n2809), .Z(n4125) );
  ND2I U3602 ( .A(n4125), .B(n2963), .Z(n2811) );
  ND2I U3603 ( .A(n3186), .B(n3929), .Z(n3178) );
  ND2I U3604 ( .A(n3118), .B(n2966), .Z(n2810) );
  ND4P U3605 ( .A(n2812), .B(n2811), .C(n3178), .D(n2810), .Z(n4079) );
  ND2I U3606 ( .A(n4553), .B(n1155), .Z(n2813) );
  AN2I U3607 ( .A(n2814), .B(n2813), .Z(n2821) );
  ND2I U3608 ( .A(n2948), .B(n3035), .Z(n3163) );
  ND2I U3609 ( .A(n2929), .B(n3165), .Z(n2946) );
  ND2I U3610 ( .A(n3013), .B(n3781), .Z(n2949) );
  ND4P U3611 ( .A(n3163), .B(n2946), .C(n2815), .D(n2949), .Z(n4516) );
  ND2I U3612 ( .A(n4452), .B(n4516), .Z(n2818) );
  ND2I U3613 ( .A(n2816), .B(n3194), .Z(n4045) );
  IVI U3614 ( .A(n4045), .Z(n3943) );
  ND2I U3615 ( .A(n3943), .B(n4461), .Z(n2817) );
  ND2I U3616 ( .A(n2818), .B(n2817), .Z(n2819) );
  IVI U3617 ( .A(n2819), .Z(n2820) );
  ND2I U3618 ( .A(n2821), .B(n2820), .Z(n2822) );
  NR2I U3619 ( .A(n2823), .B(n2822), .Z(n2824) );
  ND2I U3620 ( .A(n2825), .B(n2824), .Z(x_ALU_Result[16]) );
  ENI U3621 ( .A(n2826), .B(n1182), .Z(n2829) );
  EOI U3622 ( .A(n2827), .B(n2829), .Z(n2852) );
  B2I U3623 ( .A(n2830), .Z2(n4268) );
  MUX21L U3624 ( .A(n2852), .B(n2853), .S(n4268), .Z(n2831) );
  NR2I U3625 ( .A(n2831), .B(n2781), .Z(n2835) );
  ND2I U3626 ( .A(n1198), .B(n2684), .Z(n4271) );
  IVI U3627 ( .A(n4271), .Z(n2834) );
  ND2I U3628 ( .A(n2835), .B(n2834), .Z(n2850) );
  ND2I U3629 ( .A(n1445), .B(n2836), .Z(n2838) );
  ND2I U3630 ( .A(n4239), .B(n4453), .Z(n2837) );
  AN2I U3631 ( .A(n2838), .B(n2837), .Z(n2840) );
  ND2I U3632 ( .A(n4412), .B(n4460), .Z(n2839) );
  ND2I U3633 ( .A(n2840), .B(n2839), .Z(n4533) );
  ND2I U3634 ( .A(n4504), .B(n4533), .Z(n2848) );
  IVI U3635 ( .A(n2841), .Z(n2903) );
  IVI U3636 ( .A(n2842), .Z(n2843) );
  ND2I U3637 ( .A(n2844), .B(n2843), .Z(n2902) );
  IVI U3638 ( .A(n2902), .Z(n2845) );
  AN2I U3639 ( .A(n3928), .B(n2845), .Z(n2846) );
  ND2I U3640 ( .A(n2903), .B(n2846), .Z(n3925) );
  IVI U3641 ( .A(n3925), .Z(n2860) );
  AN2I U3642 ( .A(n4412), .B(n2860), .Z(n3161) );
  ND2I U3643 ( .A(n4540), .B(n3161), .Z(n2847) );
  AN2I U3644 ( .A(n2848), .B(n2847), .Z(n2849) );
  ND2I U3645 ( .A(n2850), .B(n2849), .Z(n2870) );
  ND2I U3646 ( .A(n4271), .B(n4041), .Z(n2868) );
  IVDA U3647 ( .A(n2851), .Z(n4269) );
  MUX21L U3648 ( .A(n2853), .B(n2852), .S(n4269), .Z(n2867) );
  MUX21L U3649 ( .A(n4314), .B(n4313), .S(n1183), .Z(n2854) );
  ND2I U3650 ( .A(n4642), .B(n2854), .Z(n2856) );
  B2I U3651 ( .A(n2855), .Z2(n3331) );
  ND2I U3652 ( .A(n2856), .B(n3331), .Z(n2859) );
  IVI U3653 ( .A(n4496), .Z(n4317) );
  AO7 U3654 ( .A(n4317), .B(n3331), .C(n4642), .Z(n2857) );
  ND2I U3655 ( .A(n1182), .B(n2857), .Z(n2858) );
  AN2I U3656 ( .A(n2859), .B(n2858), .Z(n2866) );
  ND2I U3657 ( .A(n1157), .B(n3856), .Z(n2861) );
  IVI U3658 ( .A(n2861), .Z(n3795) );
  ND4P U3659 ( .A(n4556), .B(n2864), .C(n2863), .D(n2862), .Z(n4547) );
  ND2I U3660 ( .A(n1178), .B(n4547), .Z(n2865) );
  AO3P U3661 ( .A(n2868), .B(n2867), .C(n2866), .D(n2865), .Z(n2869) );
  NR2I U3662 ( .A(n2870), .B(n2869), .Z(n2883) );
  IVI U3663 ( .A(n2871), .Z(n2872) );
  ND2I U3664 ( .A(n2872), .B(n4583), .Z(n3807) );
  IVI U3665 ( .A(n3807), .Z(n4251) );
  IVDA U3666 ( .A(n3874), .Y(n1454), .Z(n3051) );
  AN2I U3667 ( .A(n4293), .B(n1445), .Z(n3906) );
  AO2 U3668 ( .A(n4251), .B(n3051), .C(n3906), .D(n1153), .Z(n2881) );
  ND2I U3669 ( .A(n2872), .B(n4239), .Z(n2994) );
  IVI U3670 ( .A(n2994), .Z(n4373) );
  AN2I U3671 ( .A(n4293), .B(n4412), .Z(n4541) );
  ND2I U3672 ( .A(n3118), .B(n4037), .Z(n4110) );
  AO2 U3673 ( .A(n4373), .B(n3905), .C(n4541), .D(n3907), .Z(n2880) );
  AN2I U3674 ( .A(n2881), .B(n2880), .Z(n2882) );
  ND2I U3675 ( .A(n2883), .B(n2882), .Z(x_ALU_Result[11]) );
  ND2I U3676 ( .A(n2885), .B(n2884), .Z(n2901) );
  NR2I U3677 ( .A(n4619), .B(n3763), .Z(n2899) );
  IVI U3678 ( .A(n1445), .Z(n4623) );
  ND4 U3679 ( .A(n2897), .B(n2896), .C(n2895), .D(n2894), .Z(n2995) );
  AO4 U3680 ( .A(n4623), .B(n3097), .C(n4621), .D(n2995), .Z(n2898) );
  NR2I U3681 ( .A(n2899), .B(n2898), .Z(n2900) );
  AN2I U3682 ( .A(n3856), .B(n4626), .Z(n4635) );
  IVI U3683 ( .A(n3136), .Z(n3365) );
  IVI U3684 ( .A(n2966), .Z(n3358) );
  ND2I U3685 ( .A(n1174), .B(n2905), .Z(n2914) );
  IVI U3686 ( .A(n3022), .Z(n4641) );
  IVI U3687 ( .A(n2909), .Z(n4640) );
  AO6 U3688 ( .A(n2911), .B(n4672), .C(n2910), .Z(n2913) );
  ND2I U3689 ( .A(n4452), .B(n3765), .Z(n2912) );
  AO3P U3690 ( .A(n2915), .B(n2914), .C(n2913), .D(n2912), .Z(x_ALU_Result[1])
         );
  AO7 U3691 ( .A(n4020), .B(n3918), .C(n4643), .Z(n2916) );
  ND2I U3692 ( .A(n2963), .B(n2916), .Z(n2918) );
  AN2I U3693 ( .A(n2918), .B(n2917), .Z(n2970) );
  IVI U3694 ( .A(n4653), .Z(n4629) );
  IVI U3695 ( .A(n4650), .Z(n4633) );
  MUX21L U3696 ( .A(n4629), .B(n4633), .S(n1149), .Z(n2920) );
  AN2I U3697 ( .A(n2921), .B(n2920), .Z(n3030) );
  IVI U3698 ( .A(n3030), .Z(n2928) );
  ND2I U3699 ( .A(n2922), .B(n4303), .Z(n4279) );
  ND2I U3700 ( .A(n2923), .B(n4565), .Z(n2926) );
  ND2I U3701 ( .A(n3117), .B(n4424), .Z(n2925) );
  ND2I U3702 ( .A(n3013), .B(n4601), .Z(n2924) );
  ND4P U3703 ( .A(n4279), .B(n2926), .C(n2925), .D(n2924), .Z(n3852) );
  IVI U3704 ( .A(n3852), .Z(n2927) );
  MUX21L U3705 ( .A(n2928), .B(n2927), .S(n3871), .Z(n4295) );
  ND2I U3706 ( .A(n4295), .B(n3031), .Z(n2941) );
  ND2I U3707 ( .A(n2929), .B(n4470), .Z(n4410) );
  ND2I U3708 ( .A(n3013), .B(n4385), .Z(n2930) );
  ND2I U3709 ( .A(n4410), .B(n2930), .Z(n2931) );
  IVI U3710 ( .A(n2931), .Z(n2934) );
  ND2I U3711 ( .A(n3117), .B(n4524), .Z(n4278) );
  ND2I U3712 ( .A(n4403), .B(n4343), .Z(n4298) );
  ND2I U3713 ( .A(n4278), .B(n4298), .Z(n2932) );
  IVI U3714 ( .A(n2932), .Z(n2933) );
  AN2I U3715 ( .A(n2934), .B(n2933), .Z(n3855) );
  IVI U3716 ( .A(n3855), .Z(n2935) );
  ND2I U3717 ( .A(n4412), .B(n2935), .Z(n2938) );
  ND2I U3718 ( .A(n2936), .B(n4037), .Z(n4015) );
  ND2I U3719 ( .A(n4591), .B(n4086), .Z(n4072) );
  ND2I U3720 ( .A(n4632), .B(n4181), .Z(n4299) );
  ND2I U3721 ( .A(n3013), .B(n4227), .Z(n4490) );
  ND2I U3722 ( .A(n4257), .B(n3856), .Z(n2937) );
  ND2I U3723 ( .A(n2938), .B(n2937), .Z(n2939) );
  IVI U3724 ( .A(n2939), .Z(n2940) );
  ND2I U3725 ( .A(n2941), .B(n2940), .Z(n4012) );
  IVI U3726 ( .A(n4012), .Z(n2955) );
  ND2I U3727 ( .A(n2942), .B(n1187), .Z(n3009) );
  ND2I U3728 ( .A(n4125), .B(n3156), .Z(n3017) );
  ND4 U3729 ( .A(n3009), .B(n3017), .C(n2944), .D(n2943), .Z(n3837) );
  ND2I U3730 ( .A(n3013), .B(n2945), .Z(n4071) );
  ND2I U3731 ( .A(n3186), .B(n3035), .Z(n3014) );
  ND2I U3732 ( .A(n2948), .B(n2947), .Z(n4013) );
  IVI U3733 ( .A(n3836), .Z(n4255) );
  ND2I U3734 ( .A(n4583), .B(n4255), .Z(n2953) );
  ND2I U3735 ( .A(n2951), .B(n3813), .Z(n3015) );
  ND2I U3736 ( .A(n2942), .B(n4265), .Z(n3016) );
  IVI U3737 ( .A(n3849), .Z(n4262) );
  ND2I U3738 ( .A(n1445), .B(n4262), .Z(n2952) );
  MUX21L U3739 ( .A(n2955), .B(n2954), .S(n4626), .Z(n2956) );
  ND2I U3740 ( .A(n2957), .B(n2956), .Z(n2969) );
  IVI U3741 ( .A(n2958), .Z(n2959) );
  ENI U3742 ( .A(n2960), .B(n2963), .Z(n2961) );
  ENI U3743 ( .A(n2959), .B(n2961), .Z(n2962) );
  ND2I U3744 ( .A(n2962), .B(n4672), .Z(n2968) );
  ND2I U3745 ( .A(n4125), .B(n3194), .Z(n2965) );
  IVI U3746 ( .A(n2762), .Z(n4592) );
  ND2I U3747 ( .A(n4592), .B(n2963), .Z(n2964) );
  ND2I U3748 ( .A(n4558), .B(n4336), .Z(n2967) );
  ND4P U3749 ( .A(n2970), .B(n2969), .C(n2968), .D(n2967), .Z(x_ALU_Result[2])
         );
  ND2I U3750 ( .A(n4542), .B(n3765), .Z(n2993) );
  IVI U3751 ( .A(n3807), .Z(n3926) );
  AN2I U3752 ( .A(n3926), .B(n3780), .Z(n2991) );
  IVI U3753 ( .A(n4644), .Z(n2971) );
  ND2I U3754 ( .A(n3348), .B(n2971), .Z(n2972) );
  ND2I U3755 ( .A(n4643), .B(n2972), .Z(n2973) );
  ND2I U3756 ( .A(n3008), .B(n2973), .Z(n2975) );
  AN2I U3757 ( .A(n2975), .B(n2974), .Z(n2989) );
  ND2I U3758 ( .A(n4356), .B(n2976), .Z(n2977) );
  AN2I U3759 ( .A(n4619), .B(n2977), .Z(n4204) );
  ND2I U3760 ( .A(n2979), .B(n2978), .Z(n2980) );
  IVI U3761 ( .A(n2980), .Z(n2981) );
  ND2I U3762 ( .A(n2981), .B(n3031), .Z(n2986) );
  AN2I U3763 ( .A(n3918), .B(n2982), .Z(n2984) );
  ND2I U3764 ( .A(n2984), .B(n2983), .Z(n2985) );
  AN2I U3765 ( .A(n2986), .B(n2985), .Z(n4203) );
  IVI U3766 ( .A(n1177), .Z(n3032) );
  AN2I U3767 ( .A(n4203), .B(n3032), .Z(n2987) );
  ND2I U3768 ( .A(n4204), .B(n2987), .Z(n2988) );
  ND2I U3769 ( .A(n2989), .B(n2988), .Z(n2990) );
  NR2I U3770 ( .A(n2991), .B(n2990), .Z(n2992) );
  AN2I U3771 ( .A(n2993), .B(n2992), .Z(n3006) );
  AN2I U3772 ( .A(n3098), .B(n4412), .Z(n4513) );
  AN2I U3773 ( .A(n3856), .B(n4504), .Z(n4493) );
  AO2 U3774 ( .A(n4513), .B(n3097), .C(n4493), .D(n1166), .Z(n3005) );
  ND2I U3775 ( .A(n3763), .B(n3906), .Z(n2997) );
  IVI U3776 ( .A(n2994), .Z(n4548) );
  ND2I U3777 ( .A(n2995), .B(n4373), .Z(n2996) );
  AN2I U3778 ( .A(n2997), .B(n2996), .Z(n3004) );
  ND2I U3779 ( .A(n1437), .B(n3001), .Z(n3843) );
  ND2I U3780 ( .A(n3002), .B(n4672), .Z(n3003) );
  ND4P U3781 ( .A(n3006), .B(n3005), .C(n3004), .D(n3003), .Z(x_ALU_Result[5])
         );
  AO2 U3782 ( .A(n3906), .B(n2935), .C(n4541), .D(n4257), .Z(n3050) );
  ND2I U3783 ( .A(n3007), .B(n3929), .Z(n3011) );
  ND2I U3784 ( .A(n3118), .B(n3136), .Z(n3010) );
  ND2I U3785 ( .A(n4124), .B(n3008), .Z(n3181) );
  ND4P U3786 ( .A(n3011), .B(n3010), .C(n3181), .D(n3009), .Z(n4334) );
  ND2I U3787 ( .A(n1445), .B(n4334), .Z(n3021) );
  ND2I U3788 ( .A(n4583), .B(n4336), .Z(n3020) );
  ND2I U3789 ( .A(n4400), .B(n3781), .Z(n3166) );
  ND2I U3790 ( .A(n3013), .B(n1183), .Z(n3170) );
  ND4P U3791 ( .A(n3166), .B(n3015), .C(n3170), .D(n3014), .Z(n4330) );
  ND2I U3792 ( .A(n4239), .B(n4330), .Z(n3019) );
  ND2I U3793 ( .A(n4630), .B(n3324), .Z(n3169) );
  ND2I U3794 ( .A(n3118), .B(n3883), .Z(n3180) );
  ND4P U3795 ( .A(n3169), .B(n3017), .C(n3180), .D(n3016), .Z(n4324) );
  ND2I U3796 ( .A(n4412), .B(n4324), .Z(n3018) );
  ND4P U3797 ( .A(n3021), .B(n3020), .C(n3019), .D(n3018), .Z(n4590) );
  MUX21L U3798 ( .A(n4496), .B(n4313), .S(n3035), .Z(n3023) );
  ND2I U3799 ( .A(n4642), .B(n3023), .Z(n3025) );
  IVDA U3800 ( .A(n3024), .Z(n3307) );
  ND2I U3801 ( .A(n3025), .B(n3307), .Z(n3028) );
  AO7 U3802 ( .A(n4644), .B(n3307), .C(n4643), .Z(n3026) );
  ND2I U3803 ( .A(n3035), .B(n3026), .Z(n3027) );
  ND2I U3804 ( .A(n3028), .B(n3027), .Z(n3029) );
  AO6 U3805 ( .A(n4357), .B(n4590), .C(n3029), .Z(n3034) );
  AN2I U3806 ( .A(n3871), .B(n3030), .Z(n4598) );
  IVI U3807 ( .A(n3031), .Z(n4294) );
  AN2I U3808 ( .A(n4294), .B(n3032), .Z(n4256) );
  ND2I U3809 ( .A(n4598), .B(n4256), .Z(n3033) );
  AN2I U3810 ( .A(n3034), .B(n3033), .Z(n3049) );
  AO2 U3811 ( .A(n1151), .B(n1147), .C(n1176), .D(n3852), .Z(n3048) );
  IVI U3812 ( .A(n3069), .Z(n3037) );
  ENI U3813 ( .A(n3036), .B(n3035), .Z(n3038) );
  EOI U3814 ( .A(n3037), .B(n3038), .Z(n3043) );
  EOI U3815 ( .A(n3039), .B(n3038), .Z(n3042) );
  MUX21L U3816 ( .A(n3043), .B(n3042), .S(n1184), .Z(n3045) );
  B2I U3817 ( .A(n3041), .Z2(n3816) );
  MUX21L U3818 ( .A(n3043), .B(n3042), .S(n3816), .Z(n3044) );
  MUX21L U3819 ( .A(n3045), .B(n3044), .S(n4271), .Z(n3046) );
  ND2I U3820 ( .A(n3046), .B(n4041), .Z(n3047) );
  AO2 U3821 ( .A(n3906), .B(n3051), .C(n4513), .D(n1153), .Z(n3082) );
  ND2I U3822 ( .A(n1445), .B(n4460), .Z(n3055) );
  ND2I U3823 ( .A(n3141), .B(n3140), .Z(n3869) );
  ND2I U3824 ( .A(n4583), .B(n3869), .Z(n3054) );
  ND2I U3825 ( .A(n4412), .B(n4453), .Z(n3053) );
  ND2I U3826 ( .A(n3856), .B(n4552), .Z(n3052) );
  ND4P U3827 ( .A(n3055), .B(n3054), .C(n3053), .D(n3052), .Z(n4628) );
  ND2I U3828 ( .A(n3056), .B(n1193), .Z(n3309) );
  MUX21L U3829 ( .A(n4314), .B(n4313), .S(n3165), .Z(n3057) );
  ND2I U3830 ( .A(n4642), .B(n3057), .Z(n3058) );
  ND2I U3831 ( .A(n3309), .B(n3058), .Z(n3061) );
  AO7 U3832 ( .A(n4317), .B(n3309), .C(n4643), .Z(n3059) );
  ND2I U3833 ( .A(n3165), .B(n3059), .Z(n3060) );
  ND2I U3834 ( .A(n3061), .B(n3060), .Z(n3062) );
  AO6 U3835 ( .A(n4357), .B(n4628), .C(n3062), .Z(n3064) );
  ND2I U3836 ( .A(n3871), .B(n4540), .Z(n3873) );
  IVI U3837 ( .A(n3873), .Z(n4645) );
  ND2I U3838 ( .A(n4645), .B(n4256), .Z(n3063) );
  AN2I U3839 ( .A(n3064), .B(n3063), .Z(n3081) );
  AO2 U3840 ( .A(n4548), .B(n3907), .C(n4251), .D(n4547), .Z(n3080) );
  EOI U3841 ( .A(n3065), .B(n3165), .Z(n3068) );
  EOI U3842 ( .A(n3066), .B(n3068), .Z(n3073) );
  ENI U3843 ( .A(n3068), .B(n3067), .Z(n3072) );
  MUX21LP U3844 ( .A(n3073), .B(n3072), .S(n3069), .Z(n3075) );
  IVDA U3845 ( .A(n3070), .Y(n3039), .Z(n3071) );
  MUX21L U3846 ( .A(n3073), .B(n3072), .S(n3071), .Z(n3074) );
  MUX21L U3847 ( .A(n3075), .B(n3074), .S(n1184), .Z(n3077) );
  MUX21L U3848 ( .A(n3075), .B(n3074), .S(n3816), .Z(n3076) );
  MUX21L U3849 ( .A(n3077), .B(n3076), .S(n4271), .Z(n3078) );
  ND2I U3850 ( .A(n3078), .B(n4041), .Z(n3079) );
  ND2I U3851 ( .A(n4412), .B(n4220), .Z(n3086) );
  ND2I U3852 ( .A(n3856), .B(n3764), .Z(n3084) );
  ND2I U3853 ( .A(n1445), .B(n3765), .Z(n3083) );
  AN2I U3854 ( .A(n3084), .B(n3083), .Z(n3085) );
  ND2I U3855 ( .A(n3086), .B(n3085), .Z(n4354) );
  MUX21L U3856 ( .A(n2971), .B(n4313), .S(n3324), .Z(n3087) );
  ND2I U3857 ( .A(n4642), .B(n3087), .Z(n3089) );
  IVDA U3858 ( .A(n3088), .Z(n3326) );
  ND2I U3859 ( .A(n3089), .B(n3326), .Z(n3092) );
  AO7 U3860 ( .A(n4438), .B(n3326), .C(n4643), .Z(n3090) );
  ND2I U3861 ( .A(n3324), .B(n3090), .Z(n3091) );
  ND2I U3862 ( .A(n3092), .B(n3091), .Z(n3093) );
  AO6P U3863 ( .A(n4357), .B(n4354), .C(n3093), .Z(n3096) );
  ND2I U3864 ( .A(n3795), .B(n4372), .Z(n3095) );
  ND2I U3865 ( .A(n3161), .B(n4353), .Z(n3094) );
  AN3 U3866 ( .A(n3096), .B(n3095), .C(n3094), .Z(n3111) );
  AO2 U3867 ( .A(n1150), .B(n3097), .C(n4251), .D(n3777), .Z(n3110) );
  AN2I U3868 ( .A(n3098), .B(n1445), .Z(n4258) );
  AO2 U3869 ( .A(n4541), .B(n3763), .C(n4258), .D(n3780), .Z(n3109) );
  IVI U3870 ( .A(n3099), .Z(n3101) );
  ENI U3871 ( .A(n3100), .B(n3324), .Z(n3102) );
  ENI U3872 ( .A(n3101), .B(n3102), .Z(n3106) );
  IVI U3873 ( .A(n3102), .Z(n3103) );
  EOI U3874 ( .A(n3104), .B(n3103), .Z(n3105) );
  MUX21L U3875 ( .A(n3106), .B(n3105), .S(n4271), .Z(n3107) );
  ND2I U3876 ( .A(n3107), .B(n4041), .Z(n3108) );
  AO7 U3877 ( .A(n3362), .B(n4644), .C(n4643), .Z(n3112) );
  ND2I U3878 ( .A(n3136), .B(n3112), .Z(n3116) );
  MUX21L U3879 ( .A(n4641), .B(n4640), .S(n3136), .Z(n3113) );
  ND2I U3880 ( .A(n4643), .B(n3113), .Z(n3114) );
  ND2I U3881 ( .A(n3920), .B(n3114), .Z(n3115) );
  AN2I U3882 ( .A(n3116), .B(n3115), .Z(n3145) );
  IVI U3883 ( .A(n1187), .Z(n3351) );
  ND2I U3884 ( .A(n4635), .B(n3119), .Z(n3120) );
  AN2I U3885 ( .A(n1174), .B(n3120), .Z(n3135) );
  IVI U3886 ( .A(n3121), .Z(n3122) );
  AN2I U3887 ( .A(n3123), .B(n3122), .Z(n3133) );
  ND4 U3888 ( .A(n3127), .B(n3126), .C(n3125), .D(n3124), .Z(n3908) );
  IVI U3889 ( .A(n3907), .Z(n3128) );
  ND2I U3890 ( .A(n4583), .B(n3128), .Z(n3131) );
  IVI U3891 ( .A(n3905), .Z(n3129) );
  ND2I U3892 ( .A(n1445), .B(n3129), .Z(n3130) );
  ND2I U3893 ( .A(n3135), .B(n3134), .Z(n3144) );
  ND2I U3894 ( .A(n3139), .B(n4672), .Z(n3143) );
  ND2I U3895 ( .A(n3141), .B(n3140), .Z(n4462) );
  ND2I U3896 ( .A(n4493), .B(n4462), .Z(n3142) );
  ND4P U3897 ( .A(n3145), .B(n3144), .C(n3143), .D(n3142), .Z(x_ALU_Result[3])
         );
  ND2I U3898 ( .A(n4412), .B(n4079), .Z(n3150) );
  ND2I U3899 ( .A(n4356), .B(n3796), .Z(n3147) );
  ND2I U3900 ( .A(n3943), .B(n1445), .Z(n3146) );
  ND2I U3901 ( .A(n3147), .B(n3146), .Z(n3148) );
  IVI U3902 ( .A(n3148), .Z(n3149) );
  ND2I U3903 ( .A(n3150), .B(n3149), .Z(n4507) );
  ND2I U3904 ( .A(n4357), .B(n4507), .Z(n3160) );
  MUX21L U3905 ( .A(n4496), .B(n4313), .S(n3156), .Z(n3151) );
  ND2I U3906 ( .A(n4642), .B(n3151), .Z(n3152) );
  ND2I U3907 ( .A(n3152), .B(n3325), .Z(n3158) );
  IVDA U3908 ( .A(n3153), .Y(n3325), .Z(n3342) );
  ND2I U3909 ( .A(n3342), .B(n2971), .Z(n3154) );
  ND2I U3910 ( .A(n4643), .B(n3154), .Z(n3155) );
  ND2I U3911 ( .A(n3156), .B(n3155), .Z(n3157) );
  AN2I U3912 ( .A(n3158), .B(n3157), .Z(n3159) );
  AN2I U3913 ( .A(n3160), .B(n3159), .Z(n3162) );
  ND2I U3914 ( .A(n3118), .B(n3165), .Z(n4014) );
  AO2 U3915 ( .A(n4513), .B(n3937), .C(n1176), .D(n3810), .Z(n3176) );
  AO2 U3916 ( .A(n4548), .B(n3942), .C(n4258), .D(n3927), .Z(n3175) );
  EOI U3917 ( .A(n3171), .B(n3341), .Z(n3172) );
  ENI U3918 ( .A(n4271), .B(n3172), .Z(n3173) );
  ND2I U3919 ( .A(n3173), .B(n4041), .Z(n3174) );
  NR2I U3920 ( .A(n4619), .B(n3937), .Z(n3183) );
  ND4 U3921 ( .A(n3181), .B(n3180), .C(n3179), .D(n3178), .Z(n3944) );
  AO4 U3922 ( .A(n4623), .B(n3942), .C(n4621), .D(n3944), .Z(n3182) );
  NR2I U3923 ( .A(n3183), .B(n3182), .Z(n3184) );
  MUX21L U3924 ( .A(n3185), .B(n3184), .S(n4626), .Z(n3392) );
  IVI U3925 ( .A(n3194), .Z(n3356) );
  ND2I U3926 ( .A(n1174), .B(n3187), .Z(n3391) );
  ND2I U3927 ( .A(n3190), .B(n4672), .Z(n3197) );
  MUX21L U3928 ( .A(n4641), .B(n4640), .S(n3194), .Z(n3191) );
  ND2I U3929 ( .A(n4642), .B(n3191), .Z(n3192) );
  ND2I U3930 ( .A(n1149), .B(n3192), .Z(n3196) );
  AO7 U3931 ( .A(n1149), .B(n4438), .C(n4643), .Z(n3193) );
  ND2I U3932 ( .A(n3194), .B(n3193), .Z(n3195) );
  AN3 U3933 ( .A(n3197), .B(n3196), .C(n3195), .Z(n3199) );
  ND2I U3934 ( .A(n3943), .B(n4452), .Z(n3198) );
  AN2I U3935 ( .A(n3199), .B(n3198), .Z(n3390) );
  NR2I U3936 ( .A(n4629), .B(n4604), .Z(n3203) );
  IVI U3937 ( .A(n3200), .Z(n3202) );
  ND2I U3938 ( .A(dx_gpr_rd_data2[31]), .B(n3248), .Z(n3201) );
  ND2I U3939 ( .A(n3202), .B(n3201), .Z(n4649) );
  IVI U3940 ( .A(n4649), .Z(n3206) );
  NR2I U3941 ( .A(n3206), .B(n4650), .Z(n3209) );
  NR2I U3942 ( .A(n3203), .B(n3209), .Z(n3212) );
  IVI U3943 ( .A(n4601), .Z(n4631) );
  NR2I U3944 ( .A(n4631), .B(n4142), .Z(n3210) );
  IVI U3945 ( .A(n4424), .Z(n4634) );
  ND2I U3946 ( .A(n4634), .B(n4397), .Z(n3205) );
  ND2I U3947 ( .A(n4631), .B(n4142), .Z(n3204) );
  ND2I U3948 ( .A(n4629), .B(n4604), .Z(n3208) );
  ND2I U3949 ( .A(n3206), .B(n4650), .Z(n3207) );
  NR2I U3950 ( .A(n4634), .B(n4397), .Z(n3211) );
  NR2I U3951 ( .A(n3211), .B(n3210), .Z(n3213) );
  ND2I U3952 ( .A(n3213), .B(n3212), .Z(n3242) );
  IVI U3953 ( .A(n3242), .Z(n3235) );
  IVI U3954 ( .A(n4565), .Z(n4593) );
  ND2I U3955 ( .A(n3215), .B(n3214), .Z(n4534) );
  NR2I U3956 ( .A(n4593), .B(n4534), .Z(n3230) );
  IVI U3957 ( .A(n4303), .Z(n4401) );
  IVI U3958 ( .A(n3216), .Z(n4148) );
  ND2I U3959 ( .A(n4148), .B(n1193), .Z(n3217) );
  IVI U3960 ( .A(n3217), .Z(n3227) );
  ND2I U3961 ( .A(dx_gpr_rd_data2[26]), .B(n3218), .Z(n4145) );
  ND2I U3962 ( .A(n3227), .B(n4145), .Z(n4285) );
  NR2I U3963 ( .A(n4401), .B(n4285), .Z(n3219) );
  NR2I U3964 ( .A(n3230), .B(n3219), .Z(n3241) );
  IVI U3965 ( .A(n4385), .Z(n4404) );
  ND2I U3966 ( .A(dx_gpr_rd_data2[25]), .B(n2700), .Z(n3223) );
  ND2I U3967 ( .A(n3222), .B(n3223), .Z(n4362) );
  NR2I U3968 ( .A(n4404), .B(n4362), .Z(n3238) );
  IVI U3969 ( .A(n4524), .Z(n4160) );
  ND2I U3970 ( .A(n3221), .B(n3220), .Z(n4152) );
  B2I U3971 ( .A(n4152), .Z2(n4497) );
  ND2I U3972 ( .A(n4160), .B(n4497), .Z(n3225) );
  ND2I U3973 ( .A(n3223), .B(n3222), .Z(n4361) );
  ND2I U3974 ( .A(n4404), .B(n4361), .Z(n3224) );
  AO7 U3975 ( .A(n3238), .B(n3225), .C(n3224), .Z(n3226) );
  ND2I U3976 ( .A(n3241), .B(n3226), .Z(n3233) );
  ND2I U3977 ( .A(n3227), .B(n4145), .Z(n4284) );
  ND2I U3978 ( .A(n4401), .B(n4284), .Z(n3229) );
  ND2I U3979 ( .A(n4593), .B(n4534), .Z(n3228) );
  AO7 U3980 ( .A(n3230), .B(n3229), .C(n3228), .Z(n3231) );
  IVI U3981 ( .A(n3231), .Z(n3232) );
  ND2I U3982 ( .A(n3233), .B(n3232), .Z(n3234) );
  ND2I U3983 ( .A(n3235), .B(n3234), .Z(n3236) );
  AN2I U3984 ( .A(n3237), .B(n3236), .Z(n3290) );
  NR2I U3985 ( .A(n4160), .B(n4497), .Z(n3239) );
  NR2I U3986 ( .A(n3239), .B(n3238), .Z(n3240) );
  ND2I U3987 ( .A(n3241), .B(n3240), .Z(n3243) );
  NR2I U3988 ( .A(n3243), .B(n3242), .Z(n3300) );
  IVI U3989 ( .A(n4227), .Z(n4180) );
  ND2I U3990 ( .A(n2700), .B(dx_gpr_rd_data2[21]), .Z(n3245) );
  ND2I U3991 ( .A(n3245), .B(n3244), .Z(n4178) );
  NR2I U3992 ( .A(n4180), .B(n4208), .Z(n3266) );
  IVI U3993 ( .A(n4181), .Z(n4186) );
  B2IP U3994 ( .A(n3246), .Z1(n4056), .Z2(n4146) );
  NR2I U3995 ( .A(n3247), .B(n4056), .Z(n3249) );
  ND2I U3996 ( .A(n3254), .B(dx_gpr_rd_data2[20]), .Z(n4057) );
  ND2I U3997 ( .A(n3249), .B(n4057), .Z(n4053) );
  ND2I U3998 ( .A(n4186), .B(n4053), .Z(n3251) );
  B2I U3999 ( .A(n4178), .Z2(n4208) );
  ND2I U4000 ( .A(n4180), .B(n4208), .Z(n3250) );
  AO7 U4001 ( .A(n3266), .B(n3251), .C(n3250), .Z(n3264) );
  IVI U4002 ( .A(n4343), .Z(n3257) );
  ND2I U4003 ( .A(n3254), .B(dx_gpr_rd_data2[22]), .Z(n4170) );
  ND2I U4004 ( .A(n3252), .B(n4170), .Z(n4318) );
  NR2I U4005 ( .A(n3257), .B(n4318), .Z(n3256) );
  IVI U4006 ( .A(n4470), .Z(n4168) );
  NR2I U4007 ( .A(n3253), .B(n4056), .Z(n3255) );
  ND2I U4008 ( .A(n3248), .B(dx_gpr_rd_data2[23]), .Z(n3258) );
  ND2I U4009 ( .A(n3255), .B(n3258), .Z(n4439) );
  NR2I U4010 ( .A(n4168), .B(n4439), .Z(n3262) );
  NR2I U4011 ( .A(n3256), .B(n3262), .Z(n3267) );
  ND2I U4012 ( .A(n3257), .B(n4318), .Z(n3261) );
  ND2I U4013 ( .A(n4168), .B(n4436), .Z(n3260) );
  AO7 U4014 ( .A(n3262), .B(n3261), .C(n3260), .Z(n3263) );
  AO6 U4015 ( .A(n3264), .B(n3267), .C(n3263), .Z(n3287) );
  NR2I U4016 ( .A(n4186), .B(n4053), .Z(n3265) );
  NR2I U4017 ( .A(n3266), .B(n3265), .Z(n3268) );
  ND2I U4018 ( .A(n3268), .B(n3267), .Z(n3297) );
  IVI U4019 ( .A(n3297), .Z(n3285) );
  ND2I U4020 ( .A(n2689), .B(n3269), .Z(n4019) );
  NR2I U4021 ( .A(n3276), .B(n4019), .Z(n3270) );
  IVI U4022 ( .A(n4086), .Z(n4089) );
  NR2I U4023 ( .A(n4089), .B(n3277), .Z(n3280) );
  NR2I U4024 ( .A(n3270), .B(n3280), .Z(n3295) );
  NR2I U4025 ( .A(n3272), .B(n3271), .Z(n3293) );
  ND2I U4026 ( .A(n3292), .B(n3291), .Z(n3274) );
  ND2I U4027 ( .A(n3272), .B(n3271), .Z(n3273) );
  AO7 U4028 ( .A(n3293), .B(n3274), .C(n3273), .Z(n3275) );
  ND2I U4029 ( .A(n3295), .B(n3275), .Z(n3283) );
  ND2I U4030 ( .A(n3276), .B(n4019), .Z(n3279) );
  ND2I U4031 ( .A(n4089), .B(n3277), .Z(n3278) );
  AO7 U4032 ( .A(n3280), .B(n3279), .C(n3278), .Z(n3281) );
  IVI U4033 ( .A(n3281), .Z(n3282) );
  ND2I U4034 ( .A(n3283), .B(n3282), .Z(n3284) );
  ND2I U4035 ( .A(n3285), .B(n3284), .Z(n3286) );
  ND2I U4036 ( .A(n3287), .B(n3286), .Z(n3288) );
  ND2I U4037 ( .A(n3300), .B(n3288), .Z(n3289) );
  AN2I U4038 ( .A(n3290), .B(n3289), .Z(n3383) );
  NR2I U4039 ( .A(n3292), .B(n3291), .Z(n3294) );
  NR2I U4040 ( .A(n3294), .B(n3293), .Z(n3296) );
  ND2I U4041 ( .A(n3296), .B(n3295), .Z(n3298) );
  NR2I U4042 ( .A(n3298), .B(n3297), .Z(n3299) );
  AN2I U4043 ( .A(n3300), .B(n3299), .Z(n3381) );
  NR2I U4044 ( .A(n3308), .B(n3307), .Z(n3301) );
  NR2I U4045 ( .A(n3310), .B(n3309), .Z(n3313) );
  NR2I U4046 ( .A(n3301), .B(n3313), .Z(n3320) );
  IVI U4047 ( .A(n3781), .Z(n3303) );
  ND2I U4048 ( .A(n3317), .B(n1154), .Z(n3305) );
  B2I U4049 ( .A(n3302), .Z2(n3772) );
  ND2I U4050 ( .A(n3303), .B(n3772), .Z(n3304) );
  AO7P U4051 ( .A(n3318), .B(n3305), .C(n3304), .Z(n3306) );
  ND2I U4052 ( .A(n3320), .B(n3306), .Z(n3316) );
  ND2I U4053 ( .A(n3308), .B(n3307), .Z(n3312) );
  ND2I U4054 ( .A(n3310), .B(n3309), .Z(n3311) );
  AO7 U4055 ( .A(n3313), .B(n3312), .C(n3311), .Z(n3314) );
  IVI U4056 ( .A(n3314), .Z(n3315) );
  AN2I U4057 ( .A(n3316), .B(n3315), .Z(n3340) );
  NR2I U4058 ( .A(n3317), .B(n1154), .Z(n3319) );
  NR2I U4059 ( .A(n3319), .B(n3318), .Z(n3321) );
  ND2I U4060 ( .A(n3321), .B(n3320), .Z(n3345) );
  IVI U4061 ( .A(n3345), .Z(n3338) );
  IVI U4062 ( .A(n1180), .Z(n3330) );
  B2I U4063 ( .A(n3322), .Z2(n4246) );
  NR2I U4064 ( .A(n3330), .B(n4246), .Z(n3323) );
  NR2I U4065 ( .A(n3332), .B(n3331), .Z(n3333) );
  NR2I U4066 ( .A(n3323), .B(n3333), .Z(n3344) );
  NR2I U4067 ( .A(n2597), .B(n3326), .Z(n3343) );
  ND2I U4068 ( .A(n3341), .B(n3325), .Z(n3328) );
  ND2I U4069 ( .A(n2597), .B(n3326), .Z(n3327) );
  AO7 U4070 ( .A(n3343), .B(n3328), .C(n3327), .Z(n3329) );
  ND2I U4071 ( .A(n3344), .B(n3329), .Z(n3336) );
  IVI U4072 ( .A(n3334), .Z(n3335) );
  ND2I U4073 ( .A(n3336), .B(n3335), .Z(n3337) );
  ND2I U4074 ( .A(n3338), .B(n3337), .Z(n3339) );
  AN2I U4075 ( .A(n3340), .B(n3339), .Z(n3379) );
  NR2I U4076 ( .A(n3346), .B(n3345), .Z(n3377) );
  NR2I U4077 ( .A(n3351), .B(n3861), .Z(n3347) );
  IVI U4078 ( .A(n3883), .Z(n3352) );
  NR2I U4079 ( .A(n3352), .B(n3880), .Z(n3355) );
  NR2I U4080 ( .A(n3347), .B(n3355), .Z(n3373) );
  ND2I U4081 ( .A(n3348), .B(n3008), .Z(n3349) );
  IVI U4082 ( .A(n3349), .Z(n3372) );
  ND2I U4083 ( .A(n3351), .B(n3861), .Z(n3354) );
  ND2I U4084 ( .A(n3352), .B(n3880), .Z(n3353) );
  NR2I U4085 ( .A(n3358), .B(n3357), .Z(n3361) );
  ND2I U4086 ( .A(n3356), .B(n1149), .Z(n3360) );
  ND2I U4087 ( .A(n3358), .B(n3357), .Z(n3359) );
  NR2I U4088 ( .A(n3365), .B(n3362), .Z(n3368) );
  NR2I U4089 ( .A(n3364), .B(n3918), .Z(n3363) );
  NR2I U4090 ( .A(n3368), .B(n3363), .Z(n3370) );
  ND2I U4091 ( .A(n3364), .B(n3918), .Z(n3367) );
  ND2I U4092 ( .A(n3365), .B(n3920), .Z(n3366) );
  AO7 U4093 ( .A(n3368), .B(n3367), .C(n3366), .Z(n3369) );
  ND2I U4094 ( .A(n3375), .B(n3374), .Z(n3376) );
  ND2I U4095 ( .A(n3377), .B(n3376), .Z(n3378) );
  ND2I U4096 ( .A(n3379), .B(n3378), .Z(n3380) );
  ND2I U4097 ( .A(n3381), .B(n3380), .Z(n3382) );
  ND2I U4098 ( .A(n3383), .B(n3382), .Z(n3388) );
  IVI U4099 ( .A(n3384), .Z(n3385) );
  NR2I U4100 ( .A(n3386), .B(n3385), .Z(n3387) );
  ND2I U4101 ( .A(n3388), .B(n3387), .Z(n3389) );
  AO3P U4102 ( .A(n3392), .B(n3391), .C(n3390), .D(n3389), .Z(x_ALU_Result[0])
         );
  ND2I U4103 ( .A(n3403), .B(n3402), .Z(n3541) );
  IVI U4104 ( .A(n3541), .Z(n3708) );
  IVI U4105 ( .A(n3708), .Z(n3979) );
  IVI U4106 ( .A(n3414), .Z(n3514) );
  ENI U4107 ( .A(n3514), .B(n4849), .Z(\pc_u0/pc_plus_4 [10]) );
  IVI U4108 ( .A(\pc_u0/pc_plus_4 [10]), .Z(n3401) );
  ND2I U4109 ( .A(n3394), .B(n3393), .Z(n3395) );
  AO2 U4110 ( .A(n3829), .B(n3395), .C(n3740), .D(fd_Inst[8]), .Z(n3400) );
  ENI U4111 ( .A(n3396), .B(fd_Inst[26]), .Z(n3518) );
  AN2I U4112 ( .A(n3544), .B(n3518), .Z(n3830) );
  IVI U4113 ( .A(n3427), .Z(n3526) );
  ENI U4114 ( .A(PC[10]), .B(fd_Inst[8]), .Z(n3397) );
  EOI U4115 ( .A(n3526), .B(n3397), .Z(n3398) );
  ND2I U4116 ( .A(n3830), .B(n3398), .Z(n3399) );
  AO3P U4117 ( .A(n3979), .B(n3401), .C(n3400), .D(n3399), .Z(\pc_u0/N14 ) );
  ND2I U4118 ( .A(n3403), .B(n3402), .Z(n3480) );
  IVI U4119 ( .A(n3480), .Z(n3687) );
  IVI U4120 ( .A(n3687), .Z(n3998) );
  IVI U4121 ( .A(\pc_u0/pc_plus_4 [11]), .Z(n3413) );
  AO2 U4122 ( .A(n3829), .B(n3404), .C(n3740), .D(fd_Inst[9]), .Z(n3412) );
  AN2I U4123 ( .A(n3544), .B(n3543), .Z(n3576) );
  ENI U4124 ( .A(PC[11]), .B(fd_Inst[9]), .Z(n3407) );
  ENI U4125 ( .A(n3405), .B(n3407), .Z(n3409) );
  ENI U4126 ( .A(n3407), .B(n3406), .Z(n3408) );
  MUX21L U4127 ( .A(n3409), .B(n3408), .S(n3526), .Z(n3410) );
  ND2I U4128 ( .A(n3576), .B(n3410), .Z(n3411) );
  AO3P U4129 ( .A(n3998), .B(n3413), .C(n3412), .D(n3411), .Z(\pc_u0/N15 ) );
  IVI U4130 ( .A(n3480), .Z(n3499) );
  IVI U4131 ( .A(n3499), .Z(n4009) );
  IVI U4132 ( .A(\pc_u0/pc_plus_4 [17]), .Z(n3433) );
  ND2I U4133 ( .A(n3415), .B(gpr_rd_data1[17]), .Z(n3416) );
  ND2I U4134 ( .A(n3417), .B(n3416), .Z(n3419) );
  IVI U4135 ( .A(n3418), .Z(n3740) );
  AO2 U4136 ( .A(n3829), .B(n3419), .C(n3740), .D(n3571), .Z(n3432) );
  AN2I U4137 ( .A(n3544), .B(n3518), .Z(n3663) );
  EOI U4138 ( .A(n3630), .B(PC[17]), .Z(n3422) );
  EOI U4139 ( .A(n3422), .B(n3420), .Z(n3424) );
  EOI U4140 ( .A(n3422), .B(n3421), .Z(n3423) );
  MUX21L U4141 ( .A(n3424), .B(n3423), .S(n3520), .Z(n3426) );
  MUX21L U4142 ( .A(n3424), .B(n3423), .S(n3519), .Z(n3425) );
  MUX21L U4143 ( .A(n3426), .B(n3425), .S(n3462), .Z(n3429) );
  MUX21L U4144 ( .A(n3426), .B(n3425), .S(n3461), .Z(n3428) );
  MUX21L U4145 ( .A(n3429), .B(n3428), .S(n3427), .Z(n3430) );
  ND2I U4146 ( .A(n3663), .B(n3430), .Z(n3431) );
  AO3P U4147 ( .A(n3981), .B(n3433), .C(n3432), .D(n3431), .Z(\pc_u0/N21 ) );
  IVI U4148 ( .A(n3541), .Z(n3666) );
  IVI U4149 ( .A(n3831), .Z(n3965) );
  IVI U4150 ( .A(\pc_u0/pc_plus_4 [20]), .Z(n3443) );
  ND2I U4151 ( .A(n3581), .B(n1195), .Z(n3434) );
  ND2I U4152 ( .A(n3435), .B(n3434), .Z(n3436) );
  AO2 U4153 ( .A(n3829), .B(n3436), .C(n4714), .D(n3740), .Z(n3442) );
  EOI U4154 ( .A(n3571), .B(PC[20]), .Z(n3437) );
  ENI U4155 ( .A(n3559), .B(n3437), .Z(n3439) );
  ENI U4156 ( .A(n3560), .B(n3437), .Z(n3438) );
  MUX21L U4157 ( .A(n3439), .B(n3438), .S(n3754), .Z(n3440) );
  ND2I U4158 ( .A(n3637), .B(n3440), .Z(n3441) );
  AO3P U4159 ( .A(n1189), .B(n3443), .C(n3442), .D(n3441), .Z(\pc_u0/N24 ) );
  IVI U4160 ( .A(n3708), .Z(n3960) );
  IVI U4161 ( .A(\pc_u0/pc_plus_4 [13]), .Z(n3455) );
  AO2 U4162 ( .A(n3829), .B(n3444), .C(n3740), .D(fd_Inst[11]), .Z(n3454) );
  ENI U4163 ( .A(PC[13]), .B(fd_Inst[11]), .Z(n3446) );
  EOI U4164 ( .A(n3446), .B(n3445), .Z(n3449) );
  EOI U4165 ( .A(n3447), .B(n3446), .Z(n3448) );
  MUX21L U4166 ( .A(n3449), .B(n3448), .S(n3490), .Z(n3451) );
  MUX21L U4167 ( .A(n3449), .B(n3448), .S(n3492), .Z(n3450) );
  MUX21L U4168 ( .A(n3451), .B(n3450), .S(n3526), .Z(n3452) );
  ND2I U4169 ( .A(n3576), .B(n3452), .Z(n3453) );
  AO3P U4170 ( .A(n3960), .B(n3455), .C(n3454), .D(n3453), .Z(\pc_u0/N17 ) );
  IVI U4171 ( .A(n3499), .Z(n3981) );
  IVI U4172 ( .A(n3456), .Z(n3513) );
  EOI U4173 ( .A(n3513), .B(PC[14]), .Z(n3457) );
  MUX21L U4174 ( .A(n4847), .B(n3457), .S(n3514), .Z(\pc_u0/pc_plus_4 [14]) );
  IVI U4175 ( .A(\pc_u0/pc_plus_4 [14]), .Z(n3467) );
  ND2I U4176 ( .A(n3581), .B(gpr_rd_data1[14]), .Z(n3458) );
  ND2I U4177 ( .A(n3459), .B(n3458), .Z(n3460) );
  AO2 U4178 ( .A(n3829), .B(n3460), .C(n3740), .D(fd_Inst[12]), .Z(n3466) );
  IVI U4179 ( .A(n3461), .Z(n3522) );
  EOI U4180 ( .A(PC[14]), .B(fd_Inst[12]), .Z(n3463) );
  ENI U4181 ( .A(n3522), .B(n3463), .Z(n3464) );
  IVI U4182 ( .A(n3462), .Z(n3523) );
  AO3P U4183 ( .A(n1179), .B(n3467), .C(n3466), .D(n3465), .Z(\pc_u0/N18 ) );
  IVI U4184 ( .A(n3974), .Z(n3722) );
  IVI U4185 ( .A(n3722), .Z(n3970) );
  IVI U4186 ( .A(n3597), .Z(n3580) );
  IVI U4187 ( .A(\pc_u0/pc_plus_4 [23]), .Z(n3479) );
  AO2 U4188 ( .A(fd_Inst[21]), .B(n3740), .C(n3829), .D(n3468), .Z(n3478) );
  ENI U4189 ( .A(n3599), .B(PC[23]), .Z(n3470) );
  EOI U4190 ( .A(n3470), .B(n3469), .Z(n3473) );
  EOI U4191 ( .A(n3471), .B(n3470), .Z(n3472) );
  IVI U4192 ( .A(n3607), .Z(n3586) );
  MUX21L U4193 ( .A(n3473), .B(n3472), .S(n3586), .Z(n3475) );
  IVI U4194 ( .A(n3608), .Z(n3587) );
  MUX21L U4195 ( .A(n3473), .B(n3472), .S(n3587), .Z(n3474) );
  MUX21L U4196 ( .A(n3475), .B(n3474), .S(n3754), .Z(n3476) );
  ND2I U4197 ( .A(n3576), .B(n3476), .Z(n3477) );
  AO3P U4198 ( .A(n1192), .B(n3479), .C(n3478), .D(n3477), .Z(\pc_u0/N27 ) );
  IVI U4199 ( .A(n3480), .Z(n3697) );
  IVI U4200 ( .A(n3697), .Z(n3962) );
  IVI U4201 ( .A(\pc_u0/pc_plus_4 [26]), .Z(n3486) );
  AO2 U4202 ( .A(fd_Inst[24]), .B(n3740), .C(n3829), .D(n3481), .Z(n3485) );
  EOI U4203 ( .A(n3630), .B(PC[26]), .Z(n3482) );
  ENI U4204 ( .A(n3750), .B(n3482), .Z(n3483) );
  AO3P U4205 ( .A(n1191), .B(n3486), .C(n3485), .D(n3484), .Z(\pc_u0/N30 ) );
  EOI U4206 ( .A(n3487), .B(PC[12]), .Z(n3488) );
  MUX21L U4207 ( .A(n4848), .B(n3488), .S(n3514), .Z(\pc_u0/pc_plus_4 [12]) );
  IVI U4208 ( .A(\pc_u0/pc_plus_4 [12]), .Z(n3498) );
  AO2 U4209 ( .A(n3829), .B(n3489), .C(n3740), .D(fd_Inst[10]), .Z(n3497) );
  EOI U4210 ( .A(PC[12]), .B(fd_Inst[10]), .Z(n3491) );
  ENI U4211 ( .A(n3490), .B(n3491), .Z(n3494) );
  ENI U4212 ( .A(n3492), .B(n3491), .Z(n3493) );
  MUX21L U4213 ( .A(n3494), .B(n3493), .S(n3526), .Z(n3495) );
  ND2I U4214 ( .A(n3637), .B(n3495), .Z(n3496) );
  AO3P U4215 ( .A(n3987), .B(n3498), .C(n3497), .D(n3496), .Z(\pc_u0/N16 ) );
  IVI U4216 ( .A(n3499), .Z(n4011) );
  IVI U4217 ( .A(\pc_u0/pc_plus_4 [15]), .Z(n3511) );
  AO2 U4218 ( .A(n3829), .B(n3500), .C(n3740), .D(fd_Inst[13]), .Z(n3510) );
  ENI U4219 ( .A(PC[15]), .B(fd_Inst[13]), .Z(n3502) );
  EOI U4220 ( .A(n3502), .B(n3501), .Z(n3505) );
  EOI U4221 ( .A(n3503), .B(n3502), .Z(n3504) );
  MUX21L U4222 ( .A(n3505), .B(n3504), .S(n3522), .Z(n3507) );
  MUX21L U4223 ( .A(n3505), .B(n3504), .S(n3523), .Z(n3506) );
  MUX21L U4224 ( .A(n3507), .B(n3506), .S(n3526), .Z(n3508) );
  ND2I U4225 ( .A(n3576), .B(n3508), .Z(n3509) );
  AO3P U4226 ( .A(n4011), .B(n3511), .C(n3510), .D(n3509), .Z(\pc_u0/N19 ) );
  IVI U4227 ( .A(n3697), .Z(n4005) );
  IVI U4228 ( .A(\pc_u0/pc_plus_4 [16]), .Z(n3532) );
  ND2I U4229 ( .A(n3581), .B(gpr_rd_data1[16]), .Z(n3515) );
  ND2I U4230 ( .A(n3516), .B(n3515), .Z(n3517) );
  AO2 U4231 ( .A(n3829), .B(n3517), .C(n3740), .D(fd_Inst[14]), .Z(n3531) );
  AN2I U4232 ( .A(n3544), .B(n3518), .Z(n3758) );
  ENI U4233 ( .A(PC[16]), .B(fd_Inst[14]), .Z(n3521) );
  MUX21L U4234 ( .A(n3525), .B(n3524), .S(n3522), .Z(n3528) );
  MUX21L U4235 ( .A(n3525), .B(n3524), .S(n3523), .Z(n3527) );
  MUX21L U4236 ( .A(n3528), .B(n3527), .S(n3526), .Z(n3529) );
  ND2I U4237 ( .A(n3758), .B(n3529), .Z(n3530) );
  AO3P U4238 ( .A(n4009), .B(n3532), .C(n3531), .D(n3530), .Z(\pc_u0/N20 ) );
  IVI U4239 ( .A(n3687), .Z(n4007) );
  ENI U4240 ( .A(n3739), .B(n4846), .Z(\pc_u0/pc_plus_4 [18]) );
  IVI U4241 ( .A(\pc_u0/pc_plus_4 [18]), .Z(n3540) );
  ND2I U4242 ( .A(n3534), .B(n3533), .Z(n3535) );
  AO2 U4243 ( .A(n3829), .B(n3535), .C(n4713), .D(n3740), .Z(n3539) );
  ENI U4244 ( .A(n3630), .B(PC[18]), .Z(n3536) );
  EOI U4245 ( .A(n3754), .B(n3536), .Z(n3537) );
  ND2I U4246 ( .A(n3637), .B(n3537), .Z(n3538) );
  AO3P U4247 ( .A(n3996), .B(n3540), .C(n3539), .D(n3538), .Z(\pc_u0/N22 ) );
  IVI U4248 ( .A(n3541), .Z(n3736) );
  IVI U4249 ( .A(n3736), .Z(n4000) );
  IVI U4250 ( .A(\pc_u0/pc_plus_4 [19]), .Z(n3553) );
  AO2 U4251 ( .A(n3829), .B(n3542), .C(n4862), .D(n3740), .Z(n3552) );
  AN2I U4252 ( .A(n3544), .B(n3543), .Z(n3693) );
  ENI U4253 ( .A(n3742), .B(PC[19]), .Z(n3547) );
  ENI U4254 ( .A(n3545), .B(n3547), .Z(n3549) );
  ENI U4255 ( .A(n3547), .B(n3546), .Z(n3548) );
  MUX21L U4256 ( .A(n3549), .B(n3548), .S(n3754), .Z(n3550) );
  ND2I U4257 ( .A(n3693), .B(n3550), .Z(n3551) );
  AO3P U4258 ( .A(n4000), .B(n3553), .C(n3552), .D(n3551), .Z(\pc_u0/N23 ) );
  IVI U4259 ( .A(\pc_u0/pc_plus_4 [21]), .Z(n3568) );
  AO2 U4260 ( .A(n3829), .B(n3555), .C(n4859), .D(n3740), .Z(n3567) );
  ENI U4261 ( .A(n3571), .B(PC[21]), .Z(n3557) );
  EOI U4262 ( .A(n3557), .B(n3556), .Z(n3562) );
  EOI U4263 ( .A(n3558), .B(n3557), .Z(n3561) );
  MUX21L U4264 ( .A(n3562), .B(n3561), .S(n3559), .Z(n3564) );
  MUX21L U4265 ( .A(n3562), .B(n3561), .S(n3560), .Z(n3563) );
  MUX21L U4266 ( .A(n3564), .B(n3563), .S(n3754), .Z(n3565) );
  ND2I U4267 ( .A(n3663), .B(n3565), .Z(n3566) );
  AO3P U4268 ( .A(n3979), .B(n3568), .C(n3567), .D(n3566), .Z(\pc_u0/N25 ) );
  EOI U4269 ( .A(n3580), .B(PC[22]), .Z(n3569) );
  MUX21L U4270 ( .A(n4842), .B(n3569), .S(n3739), .Z(\pc_u0/pc_plus_4 [22]) );
  IVI U4271 ( .A(\pc_u0/pc_plus_4 [22]), .Z(n3579) );
  AO2 U4272 ( .A(n3829), .B(n3570), .C(fd_Inst[20]), .D(n3740), .Z(n3578) );
  EOI U4273 ( .A(n3571), .B(PC[22]), .Z(n3572) );
  ENI U4274 ( .A(n3586), .B(n3572), .Z(n3574) );
  ENI U4275 ( .A(n3587), .B(n3572), .Z(n3573) );
  MUX21L U4276 ( .A(n3574), .B(n3573), .S(n3754), .Z(n3575) );
  ND2I U4277 ( .A(n3576), .B(n3575), .Z(n3577) );
  AO3P U4278 ( .A(n4005), .B(n3579), .C(n3578), .D(n3577), .Z(\pc_u0/N26 ) );
  IVI U4279 ( .A(n3736), .Z(n3984) );
  IVI U4280 ( .A(\pc_u0/pc_plus_4 [24]), .Z(n3595) );
  ND2I U4281 ( .A(n3581), .B(gpr_rd_data1[24]), .Z(n3582) );
  ND2I U4282 ( .A(n3583), .B(n3582), .Z(n3584) );
  AO2 U4283 ( .A(fd_Inst[22]), .B(n3740), .C(n3829), .D(n3584), .Z(n3594) );
  ENI U4284 ( .A(n3599), .B(PC[24]), .Z(n3585) );
  MUX21L U4285 ( .A(n3589), .B(n3588), .S(n3586), .Z(n3591) );
  MUX21L U4286 ( .A(n3589), .B(n3588), .S(n3587), .Z(n3590) );
  MUX21L U4287 ( .A(n3591), .B(n3590), .S(n3754), .Z(n3592) );
  ND2I U4288 ( .A(n3693), .B(n3592), .Z(n3593) );
  AO3P U4289 ( .A(n3984), .B(n3595), .C(n3594), .D(n3593), .Z(\pc_u0/N28 ) );
  IVI U4290 ( .A(n3666), .Z(n3993) );
  IVI U4291 ( .A(\pc_u0/pc_plus_4 [25]), .Z(n3616) );
  AO2 U4292 ( .A(fd_Inst[23]), .B(n3740), .C(n3829), .D(n3598), .Z(n3615) );
  ENI U4293 ( .A(n3599), .B(PC[25]), .Z(n3601) );
  EOI U4294 ( .A(n3601), .B(n3600), .Z(n3606) );
  EOI U4295 ( .A(n3602), .B(n3601), .Z(n3605) );
  MUX21L U4296 ( .A(n3606), .B(n3605), .S(n3603), .Z(n3610) );
  MUX21L U4297 ( .A(n3606), .B(n3605), .S(n3604), .Z(n3609) );
  MUX21H U4298 ( .A(n3610), .B(n3609), .S(n3607), .Z(n3612) );
  MUX21H U4299 ( .A(n3610), .B(n3609), .S(n3608), .Z(n3611) );
  MUX21L U4300 ( .A(n3612), .B(n3611), .S(n3754), .Z(n3613) );
  ND2I U4301 ( .A(n3693), .B(n3613), .Z(n3614) );
  AO3P U4302 ( .A(n3993), .B(n3616), .C(n3615), .D(n3614), .Z(\pc_u0/N29 ) );
  IVI U4303 ( .A(n3687), .Z(n3972) );
  IVI U4304 ( .A(\pc_u0/pc_plus_4 [27]), .Z(n3628) );
  AO2 U4305 ( .A(fd_Inst[25]), .B(n3740), .C(n3829), .D(n3617), .Z(n3627) );
  ENI U4306 ( .A(n3630), .B(PC[27]), .Z(n3619) );
  EOI U4307 ( .A(n3619), .B(n3618), .Z(n3622) );
  EOI U4308 ( .A(n3620), .B(n3619), .Z(n3621) );
  MUX21L U4309 ( .A(n3622), .B(n3621), .S(n3750), .Z(n3624) );
  MUX21L U4310 ( .A(n3622), .B(n3621), .S(n3751), .Z(n3623) );
  MUX21L U4311 ( .A(n3624), .B(n3623), .S(n3754), .Z(n3625) );
  ND2I U4312 ( .A(n3663), .B(n3625), .Z(n3626) );
  AO3P U4313 ( .A(n3967), .B(n3628), .C(n3627), .D(n3626), .Z(\pc_u0/N31 ) );
  IVI U4314 ( .A(n3736), .Z(n4002) );
  IVI U4315 ( .A(\pc_u0/pc_plus_4 [28]), .Z(n3640) );
  AO2 U4316 ( .A(n3829), .B(n3629), .C(n3740), .D(PC[28]), .Z(n3639) );
  ENI U4317 ( .A(n3630), .B(PC[28]), .Z(n3631) );
  MUX21L U4318 ( .A(n3633), .B(n3632), .S(n3750), .Z(n3635) );
  MUX21L U4319 ( .A(n3633), .B(n3632), .S(n3751), .Z(n3634) );
  MUX21L U4320 ( .A(n3635), .B(n3634), .S(n3754), .Z(n3636) );
  ND2I U4321 ( .A(n3637), .B(n3636), .Z(n3638) );
  AO3P U4322 ( .A(n4002), .B(n3640), .C(n3639), .D(n3638), .Z(n1137) );
  EOI U4323 ( .A(n4827), .B(PC[31]), .Z(n3642) );
  MUX21L U4324 ( .A(n4833), .B(n3642), .S(n3641), .Z(n3643) );
  MUX21L U4325 ( .A(n3643), .B(PC[31]), .S(n3738), .Z(n3644) );
  MUX21L U4326 ( .A(n4833), .B(n3644), .S(n3739), .Z(\pc_u0/pc_plus_4 [31]) );
  IVI U4327 ( .A(\pc_u0/pc_plus_4 [31]), .Z(n3660) );
  ND2I U4328 ( .A(n3646), .B(n3645), .Z(n3647) );
  AO2 U4329 ( .A(n3829), .B(n3647), .C(n3740), .D(PC[31]), .Z(n3659) );
  EOI U4330 ( .A(n3742), .B(PC[31]), .Z(n3648) );
  MUX21L U4331 ( .A(n3652), .B(n3651), .S(n3649), .Z(n3654) );
  MUX21L U4332 ( .A(n3652), .B(n3651), .S(n3650), .Z(n3653) );
  MUX21L U4333 ( .A(n3654), .B(n3653), .S(n3750), .Z(n3656) );
  MUX21L U4334 ( .A(n3654), .B(n3653), .S(n3751), .Z(n3655) );
  MUX21L U4335 ( .A(n3656), .B(n3655), .S(n3754), .Z(n3657) );
  ND2I U4336 ( .A(n3693), .B(n3657), .Z(n3658) );
  AO3P U4337 ( .A(n3967), .B(n3660), .C(n3659), .D(n3658), .Z(n1141) );
  IVI U4338 ( .A(n3666), .Z(n3991) );
  AO2 U4339 ( .A(fd_Inst[0]), .B(n3740), .C(n3829), .D(n3661), .Z(n3665) );
  EOI U4340 ( .A(PC[2]), .B(fd_Inst[0]), .Z(n3662) );
  ND2I U4341 ( .A(n3663), .B(n3662), .Z(n3664) );
  AO3P U4342 ( .A(n1192), .B(PC[2]), .C(n3665), .D(n3664), .Z(\pc_u0/N6 ) );
  ENI U4343 ( .A(PC[3]), .B(PC[2]), .Z(n3956) );
  AO2 U4344 ( .A(fd_Inst[1]), .B(n3740), .C(n3829), .D(n3667), .Z(n3671) );
  ND2I U4345 ( .A(n3758), .B(n3669), .Z(n3670) );
  AO3P U4346 ( .A(n3993), .B(n3956), .C(n3671), .D(n3670), .Z(\pc_u0/N7 ) );
  IVI U4347 ( .A(\pc_u0/pc_plus_4 [4]), .Z(n3678) );
  AO2 U4348 ( .A(fd_Inst[2]), .B(n3740), .C(n3829), .D(n3672), .Z(n3677) );
  IVI U4349 ( .A(n3683), .Z(n3674) );
  ENI U4350 ( .A(PC[4]), .B(fd_Inst[2]), .Z(n3673) );
  EOI U4351 ( .A(n3674), .B(n3673), .Z(n3675) );
  ND2I U4352 ( .A(n3830), .B(n3675), .Z(n3676) );
  AO3P U4353 ( .A(n3996), .B(n3678), .C(n3677), .D(n3676), .Z(\pc_u0/N8 ) );
  IVI U4354 ( .A(n3708), .Z(n3987) );
  AO2 U4355 ( .A(fd_Inst[3]), .B(n3740), .C(n3829), .D(n3680), .Z(n3686) );
  ND2I U4356 ( .A(n3693), .B(n3684), .Z(n3685) );
  AO3P U4357 ( .A(n3987), .B(n3957), .C(n3686), .D(n3685), .Z(\pc_u0/N9 ) );
  IVI U4358 ( .A(n3724), .Z(n3709) );
  EOI U4359 ( .A(n3709), .B(n4852), .Z(\pc_u0/pc_plus_4 [6]) );
  IVI U4360 ( .A(\pc_u0/pc_plus_4 [6]), .Z(n3696) );
  ND2I U4361 ( .A(n3689), .B(n3688), .Z(n3690) );
  AO2 U4362 ( .A(fd_Inst[4]), .B(n3740), .C(n3829), .D(n3690), .Z(n3695) );
  IVI U4363 ( .A(n3732), .Z(n3715) );
  ENI U4364 ( .A(PC[6]), .B(fd_Inst[4]), .Z(n3691) );
  ENI U4365 ( .A(n3715), .B(n3691), .Z(n3692) );
  ND2I U4366 ( .A(n3693), .B(n3692), .Z(n3694) );
  AO3P U4367 ( .A(n3960), .B(n3696), .C(n3695), .D(n3694), .Z(\pc_u0/N10 ) );
  IVI U4368 ( .A(\pc_u0/pc_plus_4 [7]), .Z(n3707) );
  AO2 U4369 ( .A(fd_Inst[5]), .B(n3740), .C(n3829), .D(n3698), .Z(n3706) );
  EOI U4370 ( .A(fd_Inst[5]), .B(PC[7]), .Z(n3701) );
  EOI U4371 ( .A(n3701), .B(n3699), .Z(n3703) );
  EOI U4372 ( .A(n3701), .B(n3700), .Z(n3702) );
  MUX21L U4373 ( .A(n3703), .B(n3702), .S(n3715), .Z(n3704) );
  ND2I U4374 ( .A(n3758), .B(n3704), .Z(n3705) );
  AO3P U4375 ( .A(n4005), .B(n3707), .C(n3706), .D(n3705), .Z(\pc_u0/N11 ) );
  IVI U4376 ( .A(\pc_u0/pc_plus_4 [8]), .Z(n3721) );
  ND2I U4377 ( .A(n3711), .B(n3710), .Z(n3712) );
  AO2 U4378 ( .A(n3829), .B(n3712), .C(n3740), .D(fd_Inst[6]), .Z(n3720) );
  IVI U4379 ( .A(n3731), .Z(n3713) );
  EOI U4380 ( .A(PC[8]), .B(fd_Inst[6]), .Z(n3714) );
  EOI U4381 ( .A(n3713), .B(n3714), .Z(n3717) );
  MUX21L U4382 ( .A(n3717), .B(n3716), .S(n3715), .Z(n3718) );
  ND2I U4383 ( .A(n3830), .B(n3718), .Z(n3719) );
  AO3P U4384 ( .A(n3970), .B(n3721), .C(n3720), .D(n3719), .Z(\pc_u0/N12 ) );
  IVI U4385 ( .A(n3722), .Z(n3996) );
  ND2I U4386 ( .A(n3726), .B(n3725), .Z(n3727) );
  AO2 U4387 ( .A(n3829), .B(n3727), .C(n3740), .D(fd_Inst[7]), .Z(n3735) );
  ND2I U4388 ( .A(n3758), .B(n3733), .Z(n3734) );
  AO3P U4389 ( .A(n1192), .B(n3958), .C(n3735), .D(n3734), .Z(\pc_u0/N13 ) );
  IVI U4390 ( .A(\pc_u0/pc_plus_4 [29]), .Z(n3761) );
  AO2 U4391 ( .A(n3829), .B(n3741), .C(n3740), .D(PC[29]), .Z(n3760) );
  ENI U4392 ( .A(n3742), .B(PC[29]), .Z(n3744) );
  EOI U4393 ( .A(n3744), .B(n3743), .Z(n3749) );
  EOI U4394 ( .A(n3745), .B(n3744), .Z(n3748) );
  MUX21H U4395 ( .A(n3749), .B(n3748), .S(n3746), .Z(n3753) );
  MUX21H U4396 ( .A(n3749), .B(n3748), .S(n3747), .Z(n3752) );
  MUX21L U4397 ( .A(n3753), .B(n3752), .S(n3750), .Z(n3756) );
  MUX21L U4398 ( .A(n3753), .B(n3752), .S(n3751), .Z(n3755) );
  MUX21L U4399 ( .A(n3756), .B(n3755), .S(n3754), .Z(n3757) );
  ND2I U4400 ( .A(n3758), .B(n3757), .Z(n3759) );
  AO3P U4401 ( .A(n3996), .B(n3761), .C(n3760), .D(n3759), .Z(n1139) );
  AO2 U4402 ( .A(n4373), .B(n3763), .C(n1178), .D(n4353), .Z(n3794) );
  ND2I U4403 ( .A(n4412), .B(n3764), .Z(n3769) );
  ND2I U4404 ( .A(n4583), .B(n3765), .Z(n3768) );
  ND2I U4405 ( .A(n1445), .B(n4220), .Z(n3767) );
  ND2I U4406 ( .A(n4356), .B(n4374), .Z(n3766) );
  ND4P U4407 ( .A(n3769), .B(n3768), .C(n3767), .D(n3766), .Z(n4123) );
  MUX21L U4408 ( .A(n2971), .B(n4313), .S(n3781), .Z(n3770) );
  ND2I U4409 ( .A(n4642), .B(n3770), .Z(n3771) );
  ND2I U4410 ( .A(n3771), .B(n3772), .Z(n3775) );
  AO7 U4411 ( .A(n4317), .B(n3772), .C(n4643), .Z(n3773) );
  ND2I U4412 ( .A(n3781), .B(n3773), .Z(n3774) );
  ND2I U4413 ( .A(n3775), .B(n3774), .Z(n3776) );
  AO6 U4414 ( .A(n4357), .B(n4123), .C(n3776), .Z(n3779) );
  ND2I U4415 ( .A(n3906), .B(n3777), .Z(n3778) );
  AN2I U4416 ( .A(n3779), .B(n3778), .Z(n3793) );
  AO2 U4417 ( .A(n1176), .B(n4372), .C(n4513), .D(n3780), .Z(n3792) );
  ENI U4418 ( .A(n3782), .B(n3781), .Z(n3785) );
  ENI U4419 ( .A(n3785), .B(n2572), .Z(n3787) );
  MUX21L U4420 ( .A(n3787), .B(n3786), .S(n1184), .Z(n3789) );
  MUX21L U4421 ( .A(n3787), .B(n3786), .S(n3816), .Z(n3788) );
  MUX21L U4422 ( .A(n3789), .B(n3788), .S(n4271), .Z(n3790) );
  ND2I U4423 ( .A(n3790), .B(n4041), .Z(n3791) );
  AO2 U4424 ( .A(n4541), .B(n3927), .C(n1178), .D(n4512), .Z(n3823) );
  ND2I U4425 ( .A(n4239), .B(n4501), .Z(n3800) );
  ND2I U4426 ( .A(n4412), .B(n3796), .Z(n3799) );
  ND2I U4427 ( .A(n1445), .B(n4079), .Z(n3798) );
  ND2I U4428 ( .A(n4502), .B(n3943), .Z(n3797) );
  ND4P U4429 ( .A(n3800), .B(n3799), .C(n3798), .D(n3797), .Z(n4406) );
  MUX21L U4430 ( .A(n4314), .B(n4313), .S(n3813), .Z(n3801) );
  ND2I U4431 ( .A(n4642), .B(n3801), .Z(n3802) );
  ND2I U4432 ( .A(n3802), .B(n1154), .Z(n3805) );
  AO7 U4433 ( .A(n4020), .B(n1154), .C(n4643), .Z(n3803) );
  ND2I U4434 ( .A(n3813), .B(n3803), .Z(n3804) );
  ND2I U4435 ( .A(n3805), .B(n3804), .Z(n3806) );
  AO6 U4436 ( .A(n4357), .B(n4406), .C(n3806), .Z(n3809) );
  IVI U4437 ( .A(n4517), .Z(n3917) );
  OR2I U4438 ( .A(n3807), .B(n3917), .Z(n3808) );
  AN2I U4439 ( .A(n3809), .B(n3808), .Z(n3822) );
  ND2I U4440 ( .A(n3810), .B(n4258), .Z(n3812) );
  ND2I U4441 ( .A(n3937), .B(n1150), .Z(n3811) );
  AN2I U4442 ( .A(n3812), .B(n3811), .Z(n3821) );
  EOI U4443 ( .A(n3814), .B(n3813), .Z(n3815) );
  ENI U4444 ( .A(n1184), .B(n3815), .Z(n3818) );
  ENI U4445 ( .A(n3816), .B(n3815), .Z(n3817) );
  MUX21L U4446 ( .A(n3818), .B(n3817), .S(n4271), .Z(n3819) );
  ND2I U4447 ( .A(n3819), .B(n4041), .Z(n3820) );
  ND4 U4448 ( .A(n3823), .B(n3822), .C(n3821), .D(n3820), .Z(x_ALU_Result[12])
         );
  ND2I U4449 ( .A(n3824), .B(\pc_u0/pc_plus_4 [0]), .Z(n3827) );
  ND2I U4450 ( .A(n3829), .B(n3825), .Z(n3826) );
  ND2I U4451 ( .A(n3827), .B(n3826), .Z(\pc_u0/N4 ) );
  ND2I U4452 ( .A(n3829), .B(n3828), .Z(n3835) );
  IVI U4453 ( .A(n3830), .Z(n3832) );
  IVI U4454 ( .A(n3831), .Z(n3967) );
  ND2I U4455 ( .A(n3832), .B(n3972), .Z(n3833) );
  ND2I U4456 ( .A(\pc_u0/pc_plus_4 [1]), .B(n3833), .Z(n3834) );
  ND2I U4457 ( .A(n3835), .B(n3834), .Z(\pc_u0/N5 ) );
  AO2 U4458 ( .A(n4511), .B(n4336), .C(n4493), .D(n4334), .Z(n3868) );
  ND2I U4459 ( .A(n1147), .B(n4258), .Z(n3839) );
  ND2I U4460 ( .A(n3837), .B(n1151), .Z(n3838) );
  B2I U4461 ( .A(n3840), .Z2(n3890) );
  EOI U4462 ( .A(n3887), .B(n1186), .Z(n3841) );
  ENI U4463 ( .A(n3890), .B(n3841), .Z(n3845) );
  ENI U4464 ( .A(n3842), .B(n3841), .Z(n3844) );
  MUX21L U4465 ( .A(n3845), .B(n3844), .S(n3843), .Z(n3846) );
  ND2I U4466 ( .A(n3846), .B(n4672), .Z(n3848) );
  ND2I U4467 ( .A(n4257), .B(n3926), .Z(n3847) );
  AN2I U4468 ( .A(n3848), .B(n3847), .Z(n3851) );
  ND2I U4469 ( .A(n3849), .B(n4513), .Z(n3850) );
  IVI U4470 ( .A(n4598), .Z(n3854) );
  AO7 U4471 ( .A(n3871), .B(n3852), .C(n4294), .Z(n3853) );
  ND2I U4472 ( .A(n3854), .B(n3853), .Z(n3858) );
  ND2I U4473 ( .A(n3856), .B(n3855), .Z(n3857) );
  ND2I U4474 ( .A(n3858), .B(n3857), .Z(n4323) );
  AO7 U4475 ( .A(n4317), .B(n3861), .C(n4643), .Z(n3859) );
  ND2I U4476 ( .A(n1186), .B(n3859), .Z(n3864) );
  MUX21L U4477 ( .A(n4314), .B(n4313), .S(n1187), .Z(n3860) );
  ND2I U4478 ( .A(n4642), .B(n3860), .Z(n3862) );
  ND2I U4479 ( .A(n3862), .B(n3861), .Z(n3863) );
  AO3 U4480 ( .A(n1177), .B(n4323), .C(n3864), .D(n3863), .Z(n3865) );
  NR2I U4481 ( .A(n3866), .B(n3865), .Z(n3867) );
  ND2I U4482 ( .A(n3868), .B(n3867), .Z(x_ALU_Result[6]) );
  AO2 U4483 ( .A(n4542), .B(n3869), .C(n4558), .D(n1164), .Z(n3916) );
  AO7 U4484 ( .A(n3871), .B(n3870), .C(n4294), .Z(n3872) );
  ND2I U4485 ( .A(n3873), .B(n3872), .Z(n3876) );
  ND2I U4486 ( .A(n4356), .B(n1454), .Z(n3875) );
  ND2I U4487 ( .A(n3876), .B(n3875), .Z(n4444) );
  IVI U4488 ( .A(n4496), .Z(n4438) );
  AO7 U4489 ( .A(n3880), .B(n4438), .C(n4643), .Z(n3877) );
  ND2I U4490 ( .A(n3883), .B(n3877), .Z(n3882) );
  MUX21L U4491 ( .A(n4641), .B(n4640), .S(n3883), .Z(n3878) );
  ND2I U4492 ( .A(n4642), .B(n3878), .Z(n3879) );
  ND2I U4493 ( .A(n3880), .B(n3879), .Z(n3881) );
  AO3 U4494 ( .A(n1177), .B(n4444), .C(n3882), .D(n3881), .Z(n3904) );
  EOI U4495 ( .A(n3884), .B(n3883), .Z(n3888) );
  EOI U4496 ( .A(n3885), .B(n3888), .Z(n3893) );
  NR2I U4497 ( .A(n3887), .B(n1186), .Z(n3889) );
  EOI U4498 ( .A(n3889), .B(n3888), .Z(n3894) );
  MUX21L U4499 ( .A(n3893), .B(n3894), .S(n3890), .Z(n3897) );
  IVDA U4500 ( .A(n3891), .Y(n3842), .Z(n3892) );
  MUX21L U4501 ( .A(n3894), .B(n3893), .S(n3892), .Z(n3896) );
  MUX21L U4502 ( .A(n3897), .B(n3896), .S(n3895), .Z(n3898) );
  IVI U4503 ( .A(n3898), .Z(n3899) );
  ND2I U4504 ( .A(n3899), .B(n4672), .Z(n3902) );
  ND2I U4505 ( .A(n4251), .B(n1153), .Z(n3901) );
  ND2I U4506 ( .A(n3902), .B(n3901), .Z(n3903) );
  NR2I U4507 ( .A(n3904), .B(n3903), .Z(n3914) );
  AN2I U4508 ( .A(n3905), .B(n4541), .Z(n3912) );
  ND2I U4509 ( .A(n3907), .B(n3906), .Z(n3910) );
  ND2I U4510 ( .A(n3908), .B(n1151), .Z(n3909) );
  ND2I U4511 ( .A(n3910), .B(n3909), .Z(n3911) );
  NR2I U4512 ( .A(n3912), .B(n3911), .Z(n3913) );
  AN2I U4513 ( .A(n3914), .B(n3913), .Z(n3915) );
  ND2I U4514 ( .A(n3916), .B(n3915), .Z(x_ALU_Result[7]) );
  ND2I U4515 ( .A(n3918), .B(n3917), .Z(n4047) );
  ND2I U4516 ( .A(n3920), .B(n3919), .Z(n4046) );
  AN2I U4517 ( .A(n3921), .B(n4239), .Z(n3922) );
  ND2I U4518 ( .A(n3923), .B(n3922), .Z(n3924) );
  AN2I U4519 ( .A(n4619), .B(n3924), .Z(n4048) );
  ENI U4520 ( .A(n3930), .B(n3929), .Z(n3931) );
  ENI U4521 ( .A(n1451), .B(n3931), .Z(n3932) );
  ND2I U4522 ( .A(n3932), .B(n4672), .Z(n3933) );
  AN2I U4523 ( .A(n3934), .B(n3933), .Z(n3936) );
  ND2I U4524 ( .A(n4452), .B(n1155), .Z(n3935) );
  ND2I U4525 ( .A(n3936), .B(n3935), .Z(n3939) );
  AN2I U4526 ( .A(n3937), .B(n4258), .Z(n3938) );
  NR2I U4527 ( .A(n3939), .B(n3938), .Z(n3940) );
  AN2I U4528 ( .A(n3941), .B(n3940), .Z(n3948) );
  ND2I U4529 ( .A(n3944), .B(n4548), .Z(n3945) );
  AN2I U4530 ( .A(n3946), .B(n3945), .Z(n3947) );
  ND2I U4531 ( .A(n3948), .B(n3947), .Z(x_ALU_Result[4]) );
  ND2I U4532 ( .A(n3950), .B(n3949), .Z(n3953) );
  MUX21LP U4533 ( .A(n4772), .B(n4717), .S(n3953), .Z(gpr_rd_addr1[4]) );
  ND2I U4534 ( .A(n3950), .B(n3949), .Z(n3954) );
  MUX21LP U4535 ( .A(n3951), .B(n4758), .S(n3954), .Z(gpr_rd_addr1[3]) );
  MUX21LP U4536 ( .A(n1446), .B(n4759), .S(n3952), .Z(gpr_rd_addr1[0]) );
  MUX21LP U4537 ( .A(n1448), .B(n4757), .S(n3953), .Z(gpr_rd_addr1[2]) );
  MUX21LP U4538 ( .A(n3955), .B(n4752), .S(n3954), .Z(gpr_rd_addr1[1]) );
  IVI U4539 ( .A(n3956), .Z(\pc_u0/pc_plus_4 [3]) );
  IVI U4540 ( .A(n3957), .Z(\pc_u0/pc_plus_4 [5]) );
  IVI U4541 ( .A(n3958), .Z(\pc_u0/pc_plus_4 [9]) );
  IVI U4542 ( .A(reset), .Z(n4873) );
  IVI U4543 ( .A(Inst[21]), .Z(n3959) );
  NR2I U4544 ( .A(n4007), .B(n3959), .Z(Inst_stall_b_j[21]) );
  IVI U4545 ( .A(Inst[11]), .Z(n3961) );
  NR2I U4546 ( .A(n3962), .B(n3961), .Z(Inst_stall_b_j[11]) );
  IVI U4547 ( .A(Inst[16]), .Z(n3963) );
  NR2I U4548 ( .A(n1171), .B(n3963), .Z(Inst_stall_b_j[16]) );
  IVI U4549 ( .A(Inst[28]), .Z(n3964) );
  NR2I U4550 ( .A(n3965), .B(n3964), .Z(Inst_stall_b_j[28]) );
  IVI U4551 ( .A(Inst[30]), .Z(n3966) );
  NR2I U4552 ( .A(n1171), .B(n3966), .Z(Inst_stall_b_j[30]) );
  IVI U4553 ( .A(Inst[26]), .Z(n3968) );
  NR2I U4554 ( .A(n3970), .B(n3968), .Z(Inst_stall_b_j[26]) );
  IVI U4555 ( .A(Inst[27]), .Z(n3969) );
  NR2I U4556 ( .A(n3970), .B(n3969), .Z(Inst_stall_b_j[27]) );
  IVI U4557 ( .A(Inst[31]), .Z(n3971) );
  NR2I U4558 ( .A(n3972), .B(n3971), .Z(Inst_stall_b_j[31]) );
  IVI U4559 ( .A(Inst[29]), .Z(n3973) );
  NR2I U4560 ( .A(n3965), .B(n3973), .Z(Inst_stall_b_j[29]) );
  IVI U4561 ( .A(Inst[24]), .Z(n3975) );
  NR2I U4562 ( .A(n4000), .B(n3975), .Z(Inst_stall_b_j[24]) );
  IVI U4563 ( .A(Inst[14]), .Z(n3976) );
  NR2I U4564 ( .A(n3965), .B(n3976), .Z(Inst_stall_b_j[14]) );
  IVI U4565 ( .A(Inst[19]), .Z(n3977) );
  NR2I U4566 ( .A(n1191), .B(n3977), .Z(Inst_stall_b_j[19]) );
  IVI U4567 ( .A(Inst[22]), .Z(n3978) );
  NR2I U4568 ( .A(n3972), .B(n3978), .Z(Inst_stall_b_j[22]) );
  IVI U4569 ( .A(Inst[12]), .Z(n3980) );
  NR2I U4570 ( .A(n1179), .B(n3980), .Z(Inst_stall_b_j[12]) );
  IVI U4571 ( .A(Inst[17]), .Z(n3982) );
  NR2I U4572 ( .A(n3962), .B(n3982), .Z(Inst_stall_b_j[17]) );
  IVI U4573 ( .A(Inst[23]), .Z(n3983) );
  NR2I U4574 ( .A(n3984), .B(n3983), .Z(Inst_stall_b_j[23]) );
  IVI U4575 ( .A(Inst[13]), .Z(n3985) );
  NR2I U4576 ( .A(n4011), .B(n3985), .Z(Inst_stall_b_j[13]) );
  IVI U4577 ( .A(Inst[18]), .Z(n3986) );
  NR2I U4578 ( .A(n1171), .B(n3986), .Z(Inst_stall_b_j[18]) );
  IVI U4579 ( .A(Inst[25]), .Z(n3988) );
  NR2I U4580 ( .A(n3991), .B(n3988), .Z(Inst_stall_b_j[25]) );
  IVI U4581 ( .A(Inst[15]), .Z(n3989) );
  NR2I U4582 ( .A(n3998), .B(n3989), .Z(Inst_stall_b_j[15]) );
  IVI U4583 ( .A(Inst[20]), .Z(n3990) );
  NR2I U4584 ( .A(n1189), .B(n3990), .Z(Inst_stall_b_j[20]) );
  IVI U4585 ( .A(Inst[2]), .Z(n3992) );
  NR2I U4586 ( .A(n3991), .B(n3992), .Z(Inst_stall_b_j[2]) );
  IVI U4587 ( .A(Inst[5]), .Z(n3994) );
  NR2I U4588 ( .A(n3991), .B(n3994), .Z(Inst_stall_b_j[5]) );
  IVI U4589 ( .A(Inst[0]), .Z(n3995) );
  NR2I U4590 ( .A(n4002), .B(n3995), .Z(Inst_stall_b_j[0]) );
  IVI U4591 ( .A(Inst[4]), .Z(n3997) );
  NR2I U4592 ( .A(n3998), .B(n3997), .Z(Inst_stall_b_j[4]) );
  IVI U4593 ( .A(Inst[3]), .Z(n3999) );
  NR2I U4594 ( .A(n4000), .B(n3999), .Z(Inst_stall_b_j[3]) );
  IVI U4595 ( .A(Inst[1]), .Z(n4001) );
  NR2I U4596 ( .A(n4002), .B(n4001), .Z(Inst_stall_b_j[1]) );
  IVI U4597 ( .A(Inst[7]), .Z(n4003) );
  NR2I U4598 ( .A(n4009), .B(n4003), .Z(Inst_stall_b_j[7]) );
  IVI U4599 ( .A(Inst[10]), .Z(n4004) );
  NR2I U4600 ( .A(n3984), .B(n4004), .Z(Inst_stall_b_j[10]) );
  IVI U4601 ( .A(Inst[8]), .Z(n4006) );
  NR2I U4602 ( .A(n4007), .B(n4006), .Z(Inst_stall_b_j[8]) );
  IVI U4603 ( .A(Inst[9]), .Z(n4008) );
  NR2I U4604 ( .A(n1189), .B(n4008), .Z(Inst_stall_b_j[9]) );
  IVI U4605 ( .A(Inst[6]), .Z(n4010) );
  NR2I U4606 ( .A(n3981), .B(n4010), .Z(Inst_stall_b_j[6]) );
  NR2I U4607 ( .A(n2955), .B(n4445), .Z(n4035) );
  AN2I U4608 ( .A(n4014), .B(n4013), .Z(n4018) );
  AN2I U4609 ( .A(n4016), .B(n4015), .Z(n4017) );
  AN2I U4610 ( .A(n4018), .B(n4017), .Z(n4582) );
  IVI U4611 ( .A(n4582), .Z(n4325) );
  ND2I U4612 ( .A(n4558), .B(n4325), .Z(n4033) );
  AN2I U4613 ( .A(n4324), .B(n4022), .Z(n4023) );
  ND2I U4614 ( .A(n4637), .B(n4023), .Z(n4024) );
  IVI U4615 ( .A(n4026), .Z(n4032) );
  ND2I U4616 ( .A(n4542), .B(n4330), .Z(n4031) );
  AN2I U4617 ( .A(n4027), .B(n4336), .Z(n4028) );
  ND2I U4618 ( .A(n4029), .B(n4028), .Z(n4030) );
  ND4P U4619 ( .A(n4033), .B(n4032), .C(n4031), .D(n4030), .Z(n4034) );
  NR2I U4620 ( .A(n4035), .B(n4034), .Z(n4044) );
  ENI U4621 ( .A(n4092), .B(n4038), .Z(n4040) );
  ENI U4622 ( .A(n4099), .B(n4038), .Z(n4039) );
  MUX21L U4623 ( .A(n4040), .B(n4039), .S(n4669), .Z(n4042) );
  ND2I U4624 ( .A(n4042), .B(n4041), .Z(n4043) );
  ND2I U4625 ( .A(n4044), .B(n4043), .Z(x_ALU_Result[18]) );
  ND2I U4626 ( .A(n4412), .B(n4532), .Z(n4335) );
  NR2I U4627 ( .A(n4045), .B(n4335), .Z(n4070) );
  ND2I U4628 ( .A(n4046), .B(n4293), .Z(n4050) );
  ND2I U4629 ( .A(n4048), .B(n4047), .Z(n4049) );
  NR2I U4630 ( .A(n4050), .B(n4049), .Z(n4066) );
  MUX21L U4631 ( .A(n4314), .B(n4313), .S(n4181), .Z(n4051) );
  ND2I U4632 ( .A(n4642), .B(n4051), .Z(n4052) );
  ND2I U4633 ( .A(n4053), .B(n4052), .Z(n4064) );
  IVI U4634 ( .A(n4054), .Z(n4055) );
  NR2I U4635 ( .A(n4056), .B(n4055), .Z(n4061) );
  ND2I U4636 ( .A(n4058), .B(n4057), .Z(n4059) );
  IVI U4637 ( .A(n4059), .Z(n4060) );
  ND2I U4638 ( .A(n4061), .B(n4060), .Z(n4184) );
  AO7 U4639 ( .A(n4184), .B(n4644), .C(n4642), .Z(n4062) );
  ND2I U4640 ( .A(n4181), .B(n4062), .Z(n4063) );
  ND2I U4641 ( .A(n4064), .B(n4063), .Z(n4065) );
  NR2I U4642 ( .A(n4066), .B(n4065), .Z(n4068) );
  ND2I U4643 ( .A(n1167), .B(n4501), .Z(n4067) );
  ND2I U4644 ( .A(n4068), .B(n4067), .Z(n4069) );
  NR2I U4645 ( .A(n4070), .B(n4069), .Z(n4085) );
  ND2I U4646 ( .A(n4072), .B(n4071), .Z(n4073) );
  IVI U4647 ( .A(n4073), .Z(n4076) );
  AN2I U4648 ( .A(n4076), .B(n1455), .Z(n4414) );
  IVI U4649 ( .A(n4414), .Z(n4510) );
  ND2I U4650 ( .A(n4493), .B(n4510), .Z(n4078) );
  ND2I U4651 ( .A(n4542), .B(n4516), .Z(n4077) );
  ND2I U4652 ( .A(n4078), .B(n4077), .Z(n4083) );
  ND2I U4653 ( .A(n4553), .B(n1158), .Z(n4081) );
  ND2I U4654 ( .A(n4461), .B(n1155), .Z(n4080) );
  ND2I U4655 ( .A(n4081), .B(n4080), .Z(n4082) );
  NR2I U4656 ( .A(n4083), .B(n4082), .Z(n4084) );
  AN2I U4657 ( .A(n4085), .B(n4084), .Z(n4109) );
  ND2I U4658 ( .A(n4087), .B(n4086), .Z(n4093) );
  IVI U4659 ( .A(n4087), .Z(n4088) );
  ND2I U4660 ( .A(n4089), .B(n4088), .Z(n4095) );
  ND2I U4661 ( .A(n4090), .B(n4095), .Z(n4091) );
  ND2I U4662 ( .A(n4093), .B(n4091), .Z(n4100) );
  ND2I U4663 ( .A(n4092), .B(n4100), .Z(n4098) );
  IVI U4664 ( .A(n4094), .Z(n4096) );
  ND2I U4665 ( .A(n4096), .B(n4095), .Z(n4097) );
  ND2I U4666 ( .A(n4093), .B(n4097), .Z(n4101) );
  ND2I U4667 ( .A(n4098), .B(n4102), .Z(n4191) );
  ENI U4668 ( .A(n4184), .B(n4183), .Z(n4182) );
  EOI U4669 ( .A(n4182), .B(n4181), .Z(n4104) );
  ENI U4670 ( .A(n4480), .B(n4104), .Z(n4106) );
  ND2I U4671 ( .A(n4100), .B(n4099), .Z(n4103) );
  ND2I U4672 ( .A(n4103), .B(n4102), .Z(n4192) );
  B2IP U4673 ( .A(n4192), .Z2(n4479) );
  ENI U4674 ( .A(n4479), .B(n4104), .Z(n4105) );
  MUX21L U4675 ( .A(n4106), .B(n4105), .S(n4576), .Z(n4107) );
  ND2I U4676 ( .A(n4107), .B(n4672), .Z(n4108) );
  ND2I U4677 ( .A(n4109), .B(n4108), .Z(x_ALU_Result[20]) );
  NR2I U4678 ( .A(n4619), .B(n4377), .Z(n4121) );
  AN2I U4679 ( .A(n4111), .B(n4110), .Z(n4115) );
  AN2I U4680 ( .A(n4113), .B(n4112), .Z(n4114) );
  ND2I U4681 ( .A(n4115), .B(n4114), .Z(n4378) );
  ND4 U4682 ( .A(n4119), .B(n4118), .C(n4117), .D(n4116), .Z(n4355) );
  AO4 U4683 ( .A(n4623), .B(n4378), .C(n4621), .D(n4355), .Z(n4120) );
  NR2I U4684 ( .A(n4121), .B(n4120), .Z(n4122) );
  MUX21L U4685 ( .A(n4123), .B(n4122), .S(n4626), .Z(n4134) );
  ND2I U4686 ( .A(n4124), .B(n4634), .Z(n4130) );
  ND2I U4687 ( .A(n4125), .B(n4593), .Z(n4129) );
  ND2I U4688 ( .A(n4126), .B(n4631), .Z(n4128) );
  ND2I U4689 ( .A(n1144), .B(n4401), .Z(n4127) );
  ND4 U4690 ( .A(n4130), .B(n4129), .C(n4128), .D(n4127), .Z(n4131) );
  ND2I U4691 ( .A(n4635), .B(n4131), .Z(n4132) );
  ND2I U4692 ( .A(n4637), .B(n4132), .Z(n4133) );
  NR2I U4693 ( .A(n4134), .B(n4133), .Z(n4138) );
  MUX21L U4694 ( .A(n4314), .B(n4313), .S(n4601), .Z(n4135) );
  ND2I U4695 ( .A(n4642), .B(n4135), .Z(n4136) );
  NR2I U4696 ( .A(n4138), .B(n4137), .Z(n4201) );
  ND2I U4697 ( .A(n4140), .B(n4139), .Z(n4399) );
  IVI U4698 ( .A(n1436), .Z(n4141) );
  ENI U4699 ( .A(n4399), .B(n4141), .Z(n4425) );
  NR2I U4700 ( .A(n4425), .B(n4424), .Z(n4603) );
  IVI U4701 ( .A(n1436), .Z(n4144) );
  ENI U4702 ( .A(n4142), .B(n4144), .Z(n4602) );
  ENI U4703 ( .A(n4602), .B(n4601), .Z(n4143) );
  ENI U4704 ( .A(n4603), .B(n4143), .Z(n4167) );
  ND2I U4705 ( .A(n4425), .B(n4424), .Z(n4605) );
  ENI U4706 ( .A(n4143), .B(n4605), .Z(n4166) );
  ENI U4707 ( .A(n4534), .B(n4144), .Z(n4566) );
  NR2I U4708 ( .A(n4566), .B(n4565), .Z(n4151) );
  ND2I U4709 ( .A(n4566), .B(n4565), .Z(n4150) );
  AN2I U4710 ( .A(n4146), .B(n4145), .Z(n4147) );
  ND2I U4711 ( .A(n4148), .B(n4147), .Z(n4149) );
  IVI U4712 ( .A(n1436), .Z(n4173) );
  ENI U4713 ( .A(n4149), .B(n4173), .Z(n4304) );
  ND2I U4714 ( .A(n4304), .B(n4303), .Z(n4567) );
  MUX21LP U4715 ( .A(n4151), .B(n4150), .S(n4567), .Z(n4165) );
  NR2I U4716 ( .A(n4304), .B(n4303), .Z(n4569) );
  MUX21LP U4717 ( .A(n4151), .B(n4150), .S(n4569), .Z(n4164) );
  ENI U4718 ( .A(n4152), .B(n1436), .Z(n4161) );
  IVI U4719 ( .A(n4161), .Z(n4525) );
  ND2I U4720 ( .A(n4525), .B(n4524), .Z(n4387) );
  IVI U4721 ( .A(n4387), .Z(n4154) );
  IVI U4722 ( .A(n4173), .Z(n4153) );
  ENI U4723 ( .A(n4361), .B(n4153), .Z(n4155) );
  ND2I U4724 ( .A(n4155), .B(n4404), .Z(n4159) );
  ND2I U4725 ( .A(n4154), .B(n4159), .Z(n4158) );
  IVI U4726 ( .A(n4155), .Z(n4386) );
  IVI U4727 ( .A(n4404), .Z(n4156) );
  ND2I U4728 ( .A(n4386), .B(n4156), .Z(n4157) );
  ND2I U4729 ( .A(n4158), .B(n4157), .Z(n4570) );
  MUX21LP U4730 ( .A(n4165), .B(n4164), .S(n4570), .Z(n4661) );
  MUX21L U4731 ( .A(n4167), .B(n4166), .S(n4661), .Z(n4196) );
  IVI U4732 ( .A(n4159), .Z(n4163) );
  ND2I U4733 ( .A(n4386), .B(n4385), .Z(n4162) );
  AN2I U4734 ( .A(n4161), .B(n4160), .Z(n4389) );
  MUX21LP U4735 ( .A(n4163), .B(n4162), .S(n4389), .Z(n4571) );
  MUX21LP U4736 ( .A(n4165), .B(n4164), .S(n4571), .Z(n4662) );
  MUX21LP U4737 ( .A(n4167), .B(n4166), .S(n1194), .Z(n4195) );
  AN2I U4738 ( .A(n4169), .B(n4168), .Z(n4176) );
  ND2I U4739 ( .A(n4471), .B(n4470), .Z(n4175) );
  AN2I U4740 ( .A(n4170), .B(n4146), .Z(n4172) );
  ND2I U4741 ( .A(n4172), .B(n1156), .Z(n4174) );
  ENI U4742 ( .A(n4174), .B(n4173), .Z(n4344) );
  ND2I U4743 ( .A(n4344), .B(n4343), .Z(n4472) );
  MUX21LP U4744 ( .A(n4176), .B(n4175), .S(n4472), .Z(n4190) );
  NR2I U4745 ( .A(n4344), .B(n4343), .Z(n4474) );
  MUX21LP U4746 ( .A(n4176), .B(n4175), .S(n4474), .Z(n4189) );
  ENI U4747 ( .A(n4178), .B(n4177), .Z(n4228) );
  IVI U4748 ( .A(n4228), .Z(n4179) );
  AN2I U4749 ( .A(n4180), .B(n4179), .Z(n4188) );
  ND2I U4750 ( .A(n4227), .B(n4228), .Z(n4187) );
  ND2I U4751 ( .A(n4182), .B(n4181), .Z(n4229) );
  MUX21LP U4752 ( .A(n4188), .B(n4187), .S(n4229), .Z(n4475) );
  MUX21LP U4753 ( .A(n4190), .B(n4189), .S(n4475), .Z(n4194) );
  ENI U4754 ( .A(n4184), .B(n1436), .Z(n4185) );
  AN2I U4755 ( .A(n4186), .B(n4185), .Z(n4231) );
  MUX21LP U4756 ( .A(n4188), .B(n4187), .S(n4231), .Z(n4476) );
  MUX21LP U4757 ( .A(n4190), .B(n4189), .S(n4476), .Z(n4193) );
  MUX21LP U4758 ( .A(n4194), .B(n4193), .S(n4191), .Z(n4665) );
  MUX21L U4759 ( .A(n4196), .B(n4195), .S(n4665), .Z(n4198) );
  MUX21LP U4760 ( .A(n4194), .B(n4193), .S(n4192), .Z(n4666) );
  MUX21L U4761 ( .A(n4196), .B(n4195), .S(n4666), .Z(n4197) );
  MUX21L U4762 ( .A(n4198), .B(n4197), .S(n4669), .Z(n4199) );
  ND2I U4763 ( .A(n4199), .B(n4672), .Z(n4200) );
  ND2I U4764 ( .A(n4201), .B(n4200), .Z(x_ALU_Result[29]) );
  NR2I U4765 ( .A(n4202), .B(n4335), .Z(n4217) );
  ND2I U4766 ( .A(n4204), .B(n4203), .Z(n4205) );
  NR2I U4767 ( .A(n4445), .B(n4205), .Z(n4213) );
  MUX21L U4768 ( .A(n4314), .B(n4313), .S(n4227), .Z(n4206) );
  ND2I U4769 ( .A(n4642), .B(n4206), .Z(n4207) );
  ND2I U4770 ( .A(n4207), .B(n4208), .Z(n4211) );
  ND2I U4771 ( .A(n4227), .B(n4209), .Z(n4210) );
  ND2I U4772 ( .A(n4211), .B(n4210), .Z(n4212) );
  NR2I U4773 ( .A(n4213), .B(n4212), .Z(n4215) );
  ND2I U4774 ( .A(n4553), .B(n3764), .Z(n4214) );
  ND2I U4775 ( .A(n4215), .B(n4214), .Z(n4216) );
  NR2I U4776 ( .A(n4217), .B(n4216), .Z(n4226) );
  ND2I U4777 ( .A(n4558), .B(n4378), .Z(n4219) );
  ND2I U4778 ( .A(n4549), .B(n4374), .Z(n4218) );
  ND2I U4779 ( .A(n4219), .B(n4218), .Z(n4224) );
  ND2I U4780 ( .A(n4542), .B(n4377), .Z(n4222) );
  ND2I U4781 ( .A(n4461), .B(n1166), .Z(n4221) );
  ND2I U4782 ( .A(n4222), .B(n4221), .Z(n4223) );
  NR2I U4783 ( .A(n4224), .B(n4223), .Z(n4225) );
  AN2I U4784 ( .A(n4226), .B(n4225), .Z(n4238) );
  ENI U4785 ( .A(n4228), .B(n4227), .Z(n4230) );
  EOI U4786 ( .A(n4230), .B(n4229), .Z(n4233) );
  EOI U4787 ( .A(n4231), .B(n4230), .Z(n4232) );
  MUX21L U4788 ( .A(n4233), .B(n4232), .S(n4480), .Z(n4235) );
  MUX21L U4789 ( .A(n4233), .B(n4232), .S(n4479), .Z(n4234) );
  MUX21L U4790 ( .A(n4235), .B(n4234), .S(n4576), .Z(n4236) );
  ND2I U4791 ( .A(n4236), .B(n4672), .Z(n4237) );
  ND2I U4792 ( .A(n4238), .B(n4237), .Z(x_ALU_Result[21]) );
  ND2I U4793 ( .A(n1445), .B(n4336), .Z(n4241) );
  ND2I U4794 ( .A(n4239), .B(n4324), .Z(n4240) );
  AN2I U4795 ( .A(n4241), .B(n4240), .Z(n4243) );
  ND2I U4796 ( .A(n4412), .B(n4334), .Z(n4242) );
  ND2I U4797 ( .A(n4243), .B(n4242), .Z(n4281) );
  MUX21L U4798 ( .A(n4314), .B(n4313), .S(n1180), .Z(n4244) );
  ND2I U4799 ( .A(n4642), .B(n4244), .Z(n4245) );
  ND2I U4800 ( .A(n4245), .B(n4246), .Z(n4249) );
  AO7 U4801 ( .A(n4438), .B(n4246), .C(n4642), .Z(n4247) );
  ND2I U4802 ( .A(n1181), .B(n4247), .Z(n4248) );
  ND2I U4803 ( .A(n4249), .B(n4248), .Z(n4250) );
  ND2I U4804 ( .A(n1176), .B(n2935), .Z(n4252) );
  AO3 U4805 ( .A(n1148), .B(n4254), .C(n4253), .D(n4252), .Z(n4264) );
  ND2I U4806 ( .A(n4295), .B(n4256), .Z(n4260) );
  ND2I U4807 ( .A(n4258), .B(n4257), .Z(n4259) );
  AO3 U4808 ( .A(n4262), .B(n4261), .C(n4260), .D(n4259), .Z(n4263) );
  NR2I U4809 ( .A(n4264), .B(n4263), .Z(n4276) );
  ENI U4810 ( .A(n4266), .B(n4265), .Z(n4270) );
  IVI U4811 ( .A(n4270), .Z(n4267) );
  ENI U4812 ( .A(n4268), .B(n4267), .Z(n4273) );
  ENI U4813 ( .A(n4270), .B(n4269), .Z(n4272) );
  MUX21L U4814 ( .A(n4273), .B(n4272), .S(n4271), .Z(n4274) );
  ND2I U4815 ( .A(n4274), .B(n4672), .Z(n4275) );
  ND2I U4816 ( .A(n4276), .B(n4275), .Z(x_ALU_Result[10]) );
  ND2I U4817 ( .A(n4549), .B(n4325), .Z(n4292) );
  ND4 U4818 ( .A(n4280), .B(n4279), .C(n4278), .D(n4277), .Z(n4587) );
  ND2I U4819 ( .A(n4452), .B(n4587), .Z(n4291) );
  ND2I U4820 ( .A(n4532), .B(n4281), .Z(n4290) );
  MUX21L U4821 ( .A(n4314), .B(n4313), .S(n4303), .Z(n4282) );
  ND2I U4822 ( .A(n4642), .B(n4282), .Z(n4283) );
  ND2I U4823 ( .A(n4284), .B(n4283), .Z(n4288) );
  AO7 U4824 ( .A(n4285), .B(n4438), .C(n4643), .Z(n4286) );
  ND2I U4825 ( .A(n4303), .B(n4286), .Z(n4287) );
  AN2I U4826 ( .A(n4288), .B(n4287), .Z(n4289) );
  ND4P U4827 ( .A(n4292), .B(n4291), .C(n4290), .D(n4289), .Z(n4302) );
  AN2I U4828 ( .A(n4294), .B(n4293), .Z(n4646) );
  ND2I U4829 ( .A(n4553), .B(n4330), .Z(n4296) );
  IVI U4830 ( .A(n4584), .Z(n4331) );
  NR2I U4831 ( .A(n4302), .B(n4301), .Z(n4312) );
  ENI U4832 ( .A(n4304), .B(n4303), .Z(n4305) );
  MUX21L U4833 ( .A(n4307), .B(n4306), .S(n4665), .Z(n4309) );
  MUX21L U4834 ( .A(n4307), .B(n4306), .S(n4666), .Z(n4308) );
  MUX21L U4835 ( .A(n4309), .B(n4308), .S(n4576), .Z(n4310) );
  ND2I U4836 ( .A(n4310), .B(n4672), .Z(n4311) );
  ND2I U4837 ( .A(n4312), .B(n4311), .Z(x_ALU_Result[26]) );
  MUX21L U4838 ( .A(n4314), .B(n4313), .S(n4343), .Z(n4315) );
  ND2I U4839 ( .A(n4642), .B(n4315), .Z(n4316) );
  ND2I U4840 ( .A(n4318), .B(n4316), .Z(n4321) );
  AO7 U4841 ( .A(n4318), .B(n4317), .C(n4643), .Z(n4319) );
  ND2I U4842 ( .A(n4343), .B(n4319), .Z(n4320) );
  AN2I U4843 ( .A(n4321), .B(n4320), .Z(n4322) );
  AO7 U4844 ( .A(n4445), .B(n4323), .C(n4322), .Z(n4329) );
  ND2I U4845 ( .A(n4553), .B(n4324), .Z(n4327) );
  ND2I U4846 ( .A(n4542), .B(n4325), .Z(n4326) );
  ND2I U4847 ( .A(n4327), .B(n4326), .Z(n4328) );
  NR2I U4848 ( .A(n4329), .B(n4328), .Z(n4342) );
  ND2I U4849 ( .A(n1167), .B(n4330), .Z(n4333) );
  ND2I U4850 ( .A(n4493), .B(n4331), .Z(n4332) );
  ND2I U4851 ( .A(n4333), .B(n4332), .Z(n4340) );
  ND2I U4852 ( .A(n4461), .B(n4334), .Z(n4338) );
  IVI U4853 ( .A(n4335), .Z(n4463) );
  ND2I U4854 ( .A(n4463), .B(n4336), .Z(n4337) );
  ND2I U4855 ( .A(n4338), .B(n4337), .Z(n4339) );
  NR2I U4856 ( .A(n4340), .B(n4339), .Z(n4341) );
  AN2I U4857 ( .A(n4342), .B(n4341), .Z(n4352) );
  ENI U4858 ( .A(n4344), .B(n4343), .Z(n4345) );
  MUX21L U4859 ( .A(n4347), .B(n4346), .S(n4480), .Z(n4349) );
  MUX21L U4860 ( .A(n4347), .B(n4346), .S(n4479), .Z(n4348) );
  MUX21L U4861 ( .A(n4349), .B(n4348), .S(n4669), .Z(n4350) );
  ND2I U4862 ( .A(n4350), .B(n4672), .Z(n4351) );
  ND2I U4863 ( .A(n4352), .B(n4351), .Z(x_ALU_Result[22]) );
  ND2I U4864 ( .A(n4532), .B(n4354), .Z(n4370) );
  AN2I U4865 ( .A(n4356), .B(n4355), .Z(n4358) );
  ND2I U4866 ( .A(n4358), .B(n4357), .Z(n4367) );
  MUX21L U4867 ( .A(n4641), .B(n4640), .S(n4385), .Z(n4359) );
  ND2I U4868 ( .A(n4642), .B(n4359), .Z(n4360) );
  ND2I U4869 ( .A(n4361), .B(n4360), .Z(n4365) );
  IVI U4870 ( .A(n4496), .Z(n4398) );
  AO7 U4871 ( .A(n4362), .B(n4398), .C(n4643), .Z(n4363) );
  ND2I U4872 ( .A(n4385), .B(n4363), .Z(n4364) );
  AN2I U4873 ( .A(n4365), .B(n4364), .Z(n4366) );
  ND2I U4874 ( .A(n4367), .B(n4366), .Z(n4368) );
  IVI U4875 ( .A(n4368), .Z(n4369) );
  ND2I U4876 ( .A(n4370), .B(n4369), .Z(n4371) );
  ND2I U4877 ( .A(n4548), .B(n4372), .Z(n4376) );
  ND2I U4878 ( .A(n4553), .B(n4374), .Z(n4375) );
  ND2I U4879 ( .A(n4376), .B(n4375), .Z(n4382) );
  ND2I U4880 ( .A(n4549), .B(n4377), .Z(n4380) );
  ND2I U4881 ( .A(n4542), .B(n4378), .Z(n4379) );
  ND2I U4882 ( .A(n4380), .B(n4379), .Z(n4381) );
  NR2I U4883 ( .A(n4382), .B(n4381), .Z(n4383) );
  AN2I U4884 ( .A(n4384), .B(n4383), .Z(n4396) );
  ENI U4885 ( .A(n4386), .B(n4385), .Z(n4388) );
  EOI U4886 ( .A(n4388), .B(n4387), .Z(n4391) );
  EOI U4887 ( .A(n4389), .B(n4388), .Z(n4390) );
  MUX21L U4888 ( .A(n4391), .B(n4390), .S(n4665), .Z(n4393) );
  MUX21L U4889 ( .A(n4391), .B(n4390), .S(n4666), .Z(n4392) );
  MUX21L U4890 ( .A(n4393), .B(n4392), .S(n4576), .Z(n4394) );
  ND2I U4891 ( .A(n4394), .B(n4672), .Z(n4395) );
  ND2I U4892 ( .A(n4396), .B(n4395), .Z(x_ALU_Result[25]) );
  AN2I U4893 ( .A(n4637), .B(n4405), .Z(n4420) );
  IVI U4894 ( .A(n4406), .Z(n4418) );
  ND2I U4895 ( .A(n4408), .B(n4407), .Z(n4409) );
  IVI U4896 ( .A(n4409), .Z(n4411) );
  AN2I U4897 ( .A(n4411), .B(n4410), .Z(n4491) );
  IVI U4898 ( .A(n4516), .Z(n4413) );
  ND2I U4899 ( .A(n4583), .B(n4413), .Z(n4416) );
  ND2I U4900 ( .A(n1445), .B(n4414), .Z(n4415) );
  MUX21L U4901 ( .A(n4418), .B(n4417), .S(n4626), .Z(n4419) );
  ND2I U4902 ( .A(n4420), .B(n4419), .Z(n4422) );
  ND2I U4903 ( .A(n1150), .B(n4512), .Z(n4421) );
  AN3 U4904 ( .A(n4423), .B(n4422), .C(n4421), .Z(n4434) );
  ENI U4905 ( .A(n4425), .B(n4424), .Z(n4426) );
  EOI U4906 ( .A(n4661), .B(n4426), .Z(n4428) );
  MUX21L U4907 ( .A(n4428), .B(n4427), .S(n4666), .Z(n4431) );
  MUX21L U4908 ( .A(n4428), .B(n4427), .S(n4665), .Z(n4430) );
  B2IP U4909 ( .A(n4483), .Z1(n4429), .Z2(n4669) );
  MUX21LP U4910 ( .A(n4431), .B(n4430), .S(n4429), .Z(n4432) );
  ND2I U4911 ( .A(n4432), .B(n4672), .Z(n4433) );
  ND2I U4912 ( .A(n4434), .B(n4433), .Z(x_ALU_Result[28]) );
  MUX21L U4913 ( .A(n4641), .B(n4640), .S(n4470), .Z(n4435) );
  ND2I U4914 ( .A(n4642), .B(n4435), .Z(n4437) );
  ND2I U4915 ( .A(n4437), .B(n4436), .Z(n4442) );
  AO7 U4916 ( .A(n4439), .B(n4438), .C(n4643), .Z(n4440) );
  ND2I U4917 ( .A(n4470), .B(n4440), .Z(n4441) );
  AN2I U4918 ( .A(n4442), .B(n4441), .Z(n4443) );
  AO7 U4919 ( .A(n4445), .B(n1152), .C(n4443), .Z(n4457) );
  AN2I U4920 ( .A(n4447), .B(n4446), .Z(n4451) );
  AN2I U4921 ( .A(n4449), .B(n4448), .Z(n4450) );
  ND2I U4922 ( .A(n4451), .B(n4450), .Z(n4622) );
  ND2I U4923 ( .A(n4452), .B(n4622), .Z(n4455) );
  ND2I U4924 ( .A(n4553), .B(n4453), .Z(n4454) );
  ND2I U4925 ( .A(n4455), .B(n4454), .Z(n4456) );
  NR2I U4926 ( .A(n4457), .B(n4456), .Z(n4469) );
  ND2I U4927 ( .A(n1167), .B(n1173), .Z(n4459) );
  ND2I U4928 ( .A(n4542), .B(n4618), .Z(n4458) );
  ND2I U4929 ( .A(n4459), .B(n4458), .Z(n4467) );
  ND2I U4930 ( .A(n4461), .B(n1164), .Z(n4465) );
  ND2I U4931 ( .A(n4463), .B(n4462), .Z(n4464) );
  ND2I U4932 ( .A(n4465), .B(n4464), .Z(n4466) );
  NR2I U4933 ( .A(n4467), .B(n4466), .Z(n4468) );
  AN2I U4934 ( .A(n4469), .B(n4468), .Z(n4489) );
  ENI U4935 ( .A(n4471), .B(n4470), .Z(n4473) );
  EOI U4936 ( .A(n4473), .B(n4472), .Z(n4478) );
  EOI U4937 ( .A(n1190), .B(n4473), .Z(n4477) );
  MUX21L U4938 ( .A(n4478), .B(n4477), .S(n4475), .Z(n4482) );
  MUX21L U4939 ( .A(n4478), .B(n4477), .S(n4476), .Z(n4481) );
  MUX21H U4940 ( .A(n4482), .B(n4481), .S(n4479), .Z(n4486) );
  MUX21H U4941 ( .A(n4482), .B(n4481), .S(n4480), .Z(n4485) );
  B2IP U4942 ( .A(n4483), .Z1(n4484), .Z2(n4576) );
  MUX21L U4943 ( .A(n4486), .B(n4485), .S(n4484), .Z(n4487) );
  ND2I U4944 ( .A(n4487), .B(n4672), .Z(n4488) );
  ND2I U4945 ( .A(n4489), .B(n4488), .Z(x_ALU_Result[23]) );
  ND2I U4946 ( .A(n4491), .B(n4490), .Z(n4492) );
  MUX21L U4947 ( .A(n4641), .B(n4640), .S(n4524), .Z(n4494) );
  ND2I U4948 ( .A(n4642), .B(n4494), .Z(n4495) );
  ND2I U4949 ( .A(n4495), .B(n4497), .Z(n4500) );
  IVI U4950 ( .A(n4496), .Z(n4644) );
  ND2I U4951 ( .A(n4524), .B(n4498), .Z(n4499) );
  AN2I U4952 ( .A(n4500), .B(n4499), .Z(n4506) );
  AN2I U4953 ( .A(n4502), .B(n4501), .Z(n4503) );
  ND2I U4954 ( .A(n4504), .B(n4503), .Z(n4505) );
  ND2I U4955 ( .A(n4507), .B(n4532), .Z(n4508) );
  ND2I U4956 ( .A(n1444), .B(n4508), .Z(n4509) );
  ND2I U4957 ( .A(n4511), .B(n4510), .Z(n4515) );
  ND2I U4958 ( .A(n4513), .B(n4512), .Z(n4514) );
  ND2I U4959 ( .A(n4515), .B(n4514), .Z(n4521) );
  ND2I U4960 ( .A(n4549), .B(n4516), .Z(n4519) );
  ND2I U4961 ( .A(n1150), .B(n4517), .Z(n4518) );
  ND2I U4962 ( .A(n4519), .B(n4518), .Z(n4520) );
  NR2I U4963 ( .A(n4521), .B(n4520), .Z(n4522) );
  AN2I U4964 ( .A(n4523), .B(n4522), .Z(n4531) );
  EOI U4965 ( .A(n4525), .B(n4524), .Z(n4526) );
  ENI U4966 ( .A(n4665), .B(n4526), .Z(n4528) );
  ENI U4967 ( .A(n4666), .B(n4526), .Z(n4527) );
  MUX21L U4968 ( .A(n4528), .B(n4527), .S(n4576), .Z(n4529) );
  ND2I U4969 ( .A(n4529), .B(n4672), .Z(n4530) );
  ND2I U4970 ( .A(n4531), .B(n4530), .Z(x_ALU_Result[24]) );
  ND2I U4971 ( .A(n4533), .B(n4532), .Z(n4539) );
  AO7 U4972 ( .A(n4534), .B(n4438), .C(n4643), .Z(n4535) );
  ND2I U4973 ( .A(n4565), .B(n4535), .Z(n4536) );
  AN2I U4974 ( .A(n4537), .B(n4536), .Z(n4538) );
  ND2I U4975 ( .A(n4539), .B(n4538), .Z(n4546) );
  ND2I U4976 ( .A(n4541), .B(n4540), .Z(n4544) );
  ND2I U4977 ( .A(n4622), .B(n4542), .Z(n4543) );
  ND2I U4978 ( .A(n4544), .B(n4543), .Z(n4545) );
  NR2I U4979 ( .A(n4546), .B(n4545), .Z(n4564) );
  ND2I U4980 ( .A(n4373), .B(n4547), .Z(n4551) );
  ND2I U4981 ( .A(n1167), .B(n4618), .Z(n4550) );
  ND2I U4982 ( .A(n4551), .B(n4550), .Z(n4562) );
  ND2I U4983 ( .A(n4553), .B(n1173), .Z(n4560) );
  ND4 U4984 ( .A(n4557), .B(n4556), .C(n4555), .D(n4554), .Z(n4620) );
  ND2I U4985 ( .A(n4558), .B(n4620), .Z(n4559) );
  ND2I U4986 ( .A(n4560), .B(n4559), .Z(n4561) );
  NR2I U4987 ( .A(n4562), .B(n4561), .Z(n4563) );
  AN2I U4988 ( .A(n4564), .B(n4563), .Z(n4581) );
  ENI U4989 ( .A(n4566), .B(n4565), .Z(n4568) );
  EOI U4990 ( .A(n4568), .B(n4567), .Z(n4573) );
  EOI U4991 ( .A(n4569), .B(n4568), .Z(n4572) );
  MUX21H U4992 ( .A(n4573), .B(n4572), .S(n4570), .Z(n4575) );
  MUX21H U4993 ( .A(n4573), .B(n4572), .S(n4571), .Z(n4574) );
  MUX21L U4994 ( .A(n4575), .B(n4574), .S(n4665), .Z(n4578) );
  MUX21L U4995 ( .A(n4575), .B(n4574), .S(n4666), .Z(n4577) );
  MUX21L U4996 ( .A(n4578), .B(n4577), .S(n4576), .Z(n4579) );
  ND2I U4997 ( .A(n4579), .B(n4672), .Z(n4580) );
  ND2I U4998 ( .A(n4581), .B(n4580), .Z(x_ALU_Result[27]) );
  ND2I U4999 ( .A(n4583), .B(n4582), .Z(n4586) );
  ND2I U5000 ( .A(n1445), .B(n4584), .Z(n4585) );
  AO3 U5001 ( .A(n4621), .B(n4587), .C(n4586), .D(n4585), .Z(n4588) );
  IVI U5002 ( .A(n4588), .Z(n4589) );
  MUX21L U5003 ( .A(n4590), .B(n4589), .S(n4626), .Z(n4597) );
  ND2I U5004 ( .A(n4635), .B(n4594), .Z(n4595) );
  ND2I U5005 ( .A(n4637), .B(n4595), .Z(n4596) );
  NR2I U5006 ( .A(n4597), .B(n4596), .Z(n4600) );
  NR2I U5007 ( .A(n4600), .B(n4599), .Z(n4617) );
  NR2I U5008 ( .A(n4602), .B(n4601), .Z(n4607) );
  ND2I U5009 ( .A(n4602), .B(n4601), .Z(n4606) );
  MUX21LP U5010 ( .A(n4607), .B(n4606), .S(n4603), .Z(n4657) );
  EOI U5011 ( .A(n4604), .B(n1436), .Z(n4654) );
  EOI U5012 ( .A(n4654), .B(n4653), .Z(n4608) );
  ENI U5013 ( .A(n4657), .B(n4608), .Z(n4610) );
  MUX21LP U5014 ( .A(n4607), .B(n4606), .S(n4605), .Z(n4658) );
  ENI U5015 ( .A(n4658), .B(n4608), .Z(n4609) );
  MUX21L U5016 ( .A(n4610), .B(n4609), .S(n4661), .Z(n4612) );
  MUX21LP U5017 ( .A(n4610), .B(n4609), .S(n4662), .Z(n4611) );
  MUX21L U5018 ( .A(n4612), .B(n4611), .S(n4665), .Z(n4614) );
  MUX21L U5019 ( .A(n4612), .B(n4611), .S(n4666), .Z(n4613) );
  MUX21L U5020 ( .A(n4614), .B(n4613), .S(n4669), .Z(n4615) );
  ND2I U5021 ( .A(n4615), .B(n4672), .Z(n4616) );
  ND2I U5022 ( .A(n4617), .B(n4616), .Z(x_ALU_Result[30]) );
  NR2I U5023 ( .A(n4619), .B(n4618), .Z(n4625) );
  AO4 U5024 ( .A(n4623), .B(n4622), .C(n4621), .D(n4620), .Z(n4624) );
  NR2I U5025 ( .A(n4625), .B(n4624), .Z(n4627) );
  MUX21L U5026 ( .A(n1165), .B(n4627), .S(n4626), .Z(n4639) );
  ND2I U5027 ( .A(n4637), .B(n4636), .Z(n4638) );
  NR2I U5028 ( .A(n4639), .B(n4638), .Z(n4648) );
  NR2I U5029 ( .A(n4648), .B(n4647), .Z(n4675) );
  EOI U5030 ( .A(n4649), .B(n1436), .Z(n4651) );
  ENI U5031 ( .A(n4651), .B(n4650), .Z(n4655) );
  ND2I U5032 ( .A(n4654), .B(n4653), .Z(n4652) );
  EOI U5033 ( .A(n4655), .B(n4652), .Z(n4660) );
  NR2I U5034 ( .A(n4654), .B(n4653), .Z(n4656) );
  EOI U5035 ( .A(n4656), .B(n4655), .Z(n4659) );
  MUX21LP U5036 ( .A(n4660), .B(n4659), .S(n4657), .Z(n4664) );
  MUX21L U5037 ( .A(n4660), .B(n4659), .S(n4658), .Z(n4663) );
  MUX21LP U5038 ( .A(n4664), .B(n4663), .S(n4661), .Z(n4668) );
  MUX21LP U5039 ( .A(n4664), .B(n4663), .S(n1194), .Z(n4667) );
  MUX21L U5040 ( .A(n4668), .B(n4667), .S(n4665), .Z(n4671) );
  MUX21L U5041 ( .A(n4668), .B(n4667), .S(n4666), .Z(n4670) );
  MUX21L U5042 ( .A(n4671), .B(n4670), .S(n4669), .Z(n4673) );
  ND2I U5043 ( .A(n4673), .B(n4672), .Z(n4674) );
  ND2I U5044 ( .A(n4675), .B(n4674), .Z(x_ALU_Result[31]) );
  MUX21H U5045 ( .A(mw_pc_plus_8[0]), .B(n4676), .S(n1461), .Z(gpr_wr_data[0])
         );
  MUX21H U5046 ( .A(mw_pc_plus_8[1]), .B(n4677), .S(n1461), .Z(gpr_wr_data[1])
         );
  MUX21H U5047 ( .A(mw_pc_plus_8[5]), .B(n4679), .S(n1461), .Z(gpr_wr_data[5])
         );
  MUX21H U5048 ( .A(mw_pc_plus_8[6]), .B(n4680), .S(n1461), .Z(gpr_wr_data[6])
         );
  MUX21H U5049 ( .A(mw_pc_plus_8[7]), .B(n4681), .S(n1461), .Z(gpr_wr_data[7])
         );
  MUX21H U5050 ( .A(mw_pc_plus_8[10]), .B(n4682), .S(n1461), .Z(
        gpr_wr_data[10]) );
  MUX21H U5051 ( .A(mw_pc_plus_8[11]), .B(n4683), .S(n1461), .Z(
        gpr_wr_data[11]) );
  MUX21H U5052 ( .A(mw_pc_plus_8[14]), .B(n4684), .S(n1461), .Z(
        gpr_wr_data[14]) );
  MUX21H U5053 ( .A(mw_pc_plus_8[18]), .B(n4686), .S(n1461), .Z(
        gpr_wr_data[18]) );
  MUX21H U5054 ( .A(mw_pc_plus_8[21]), .B(n4687), .S(n1461), .Z(
        gpr_wr_data[21]) );
  MUX21H U5055 ( .A(mw_pc_plus_8[22]), .B(n4688), .S(n1461), .Z(
        gpr_wr_data[22]) );
  MUX21H U5056 ( .A(mw_pc_plus_8[25]), .B(n4689), .S(n1461), .Z(
        gpr_wr_data[25]) );
  MUX21H U5057 ( .A(mw_pc_plus_8[28]), .B(n4690), .S(n1461), .Z(
        gpr_wr_data[28]) );
  ENI U5058 ( .A(n4711), .B(n4709), .Z(n4697) );
  ND4 U5059 ( .A(xm_Inst[31]), .B(n4698), .C(n4854), .D(n4697), .Z(n4699) );
  NR2I U5060 ( .A(n4855), .B(n4699), .Z(MemWrite) );
  NR2I U5061 ( .A(n1994), .B(n4699), .Z(MemRead) );
endmodule

