
module signext ( ip, op );
  input [15:0] ip;
  output [31:0] op;
  wire   op_31, \op[15] , \op[28] , n3;
  assign op_31 = ip[15];
  assign op[14] = ip[14];
  assign op[13] = ip[13];
  assign op[12] = ip[12];
  assign op[11] = ip[11];
  assign op[10] = ip[10];
  assign op[9] = ip[9];
  assign op[8] = ip[8];
  assign op[7] = ip[7];
  assign op[6] = ip[6];
  assign op[5] = ip[5];
  assign op[4] = ip[4];
  assign op[3] = ip[3];
  assign op[2] = ip[2];
  assign op[1] = ip[1];
  assign op[0] = ip[0];
  assign op[27] = \op[15] ;
  assign op[26] = \op[15] ;
  assign op[25] = \op[15] ;
  assign op[24] = \op[15] ;
  assign op[23] = \op[15] ;
  assign op[22] = \op[15] ;
  assign op[21] = \op[15] ;
  assign op[20] = \op[15] ;
  assign op[19] = \op[15] ;
  assign op[18] = \op[15] ;
  assign op[17] = \op[15] ;
  assign op[16] = \op[15] ;
  assign op[15] = \op[15] ;
  assign op[31] = \op[28] ;
  assign op[30] = \op[28] ;
  assign op[29] = \op[28] ;
  assign op[28] = \op[28] ;

  B4IP U1 ( .A(n3), .Z(\op[15] ) );
  IVI U2 ( .A(n3), .Z(\op[28] ) );
  IVI U3 ( .A(op_31), .Z(n3) );
endmodule


module lshift ( ip, op );
  input [31:0] ip;
  output [31:0] op;
  wire   \ip[29] , \ip[28] , \ip[27] , \ip[26] , \ip[25] , \ip[24] , \ip[23] ,
         \ip[22] , \ip[21] , \ip[20] , \ip[19] , \ip[18] , \ip[17] , \ip[16] ,
         \ip[15] , \ip[14] , \ip[13] , \ip[12] , \ip[11] , \ip[10] , \ip[9] ,
         \ip[8] , \ip[7] , \ip[6] , \ip[5] , \ip[4] , \ip[3] , \ip[2] ,
         \ip[1] , \ip[0] ;
  assign op[0] = 1'b0;
  assign op[1] = 1'b0;
  assign op[31] = \ip[29] ;
  assign \ip[29]  = ip[29];
  assign op[30] = \ip[28] ;
  assign \ip[28]  = ip[28];
  assign op[29] = \ip[27] ;
  assign \ip[27]  = ip[27];
  assign op[28] = \ip[26] ;
  assign \ip[26]  = ip[26];
  assign op[27] = \ip[25] ;
  assign \ip[25]  = ip[25];
  assign op[26] = \ip[24] ;
  assign \ip[24]  = ip[24];
  assign op[25] = \ip[23] ;
  assign \ip[23]  = ip[23];
  assign op[24] = \ip[22] ;
  assign \ip[22]  = ip[22];
  assign op[23] = \ip[21] ;
  assign \ip[21]  = ip[21];
  assign op[22] = \ip[20] ;
  assign \ip[20]  = ip[20];
  assign op[21] = \ip[19] ;
  assign \ip[19]  = ip[19];
  assign op[20] = \ip[18] ;
  assign \ip[18]  = ip[18];
  assign op[19] = \ip[17] ;
  assign \ip[17]  = ip[17];
  assign op[18] = \ip[16] ;
  assign \ip[16]  = ip[16];
  assign op[17] = \ip[15] ;
  assign \ip[15]  = ip[15];
  assign op[16] = \ip[14] ;
  assign \ip[14]  = ip[14];
  assign op[15] = \ip[13] ;
  assign \ip[13]  = ip[13];
  assign op[14] = \ip[12] ;
  assign \ip[12]  = ip[12];
  assign op[13] = \ip[11] ;
  assign \ip[11]  = ip[11];
  assign op[12] = \ip[10] ;
  assign \ip[10]  = ip[10];
  assign op[11] = \ip[9] ;
  assign \ip[9]  = ip[9];
  assign op[10] = \ip[8] ;
  assign \ip[8]  = ip[8];
  assign op[9] = \ip[7] ;
  assign \ip[7]  = ip[7];
  assign op[8] = \ip[6] ;
  assign \ip[6]  = ip[6];
  assign op[7] = \ip[5] ;
  assign \ip[5]  = ip[5];
  assign op[6] = \ip[4] ;
  assign \ip[4]  = ip[4];
  assign op[5] = \ip[3] ;
  assign \ip[3]  = ip[3];
  assign op[4] = \ip[2] ;
  assign \ip[2]  = ip[2];
  assign op[3] = \ip[1] ;
  assign \ip[1]  = ip[1];
  assign op[2] = \ip[0] ;
  assign \ip[0]  = ip[0];

endmodule


module mux_2x1_DATA_WIDTH32_0 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;

  IVI U1 ( .A(ip1[24]), .Z(n12) );
  IVI U2 ( .A(ip1[27]), .Z(n2) );
  IVI U3 ( .A(ip1[23]), .Z(n6) );
  IVI U4 ( .A(ip1[13]), .Z(n22) );
  IVI U5 ( .A(ip1[11]), .Z(n4) );
  IVI U6 ( .A(ip1[9]), .Z(n29) );
  IVI U7 ( .A(ip1[4]), .Z(n10) );
  IVI U8 ( .A(ip0[21]), .Z(n7) );
  IVI U9 ( .A(ip0[17]), .Z(n19) );
  IVI U10 ( .A(ip0[24]), .Z(n11) );
  IVI U11 ( .A(ip1[21]), .Z(n8) );
  IVI U12 ( .A(ip1[17]), .Z(n20) );
  IVI U13 ( .A(ip0[27]), .Z(n1) );
  IVI U14 ( .A(ip0[23]), .Z(n5) );
  IVI U15 ( .A(ip0[13]), .Z(n21) );
  IVI U16 ( .A(ip0[11]), .Z(n3) );
  IVI U17 ( .A(ip0[9]), .Z(n28) );
  IVI U18 ( .A(ip0[4]), .Z(n9) );
  MUX21L U19 ( .A(n1), .B(n2), .S(n17), .Z(out[27]) );
  MUX21L U20 ( .A(n3), .B(n4), .S(n17), .Z(out[11]) );
  MUX21L U21 ( .A(n5), .B(n6), .S(n31), .Z(out[23]) );
  MUX21L U22 ( .A(n7), .B(n8), .S(n31), .Z(out[21]) );
  MUX21L U23 ( .A(n9), .B(n10), .S(n32), .Z(out[4]) );
  MUX21L U24 ( .A(n12), .B(n11), .S(n23), .Z(out[24]) );
  IVI U25 ( .A(n33), .Z(n13) );
  IVI U26 ( .A(sel), .Z(n14) );
  IVI U27 ( .A(n14), .Z(n15) );
  IVI U28 ( .A(n30), .Z(n16) );
  IVI U29 ( .A(n30), .Z(n17) );
  IVI U30 ( .A(n30), .Z(n18) );
  IVI U31 ( .A(n14), .Z(n32) );
  MUX21L U32 ( .A(n19), .B(n20), .S(n25), .Z(out[17]) );
  MUX21L U33 ( .A(n22), .B(n21), .S(n23), .Z(out[13]) );
  IVI U34 ( .A(n15), .Z(n23) );
  IVI U35 ( .A(n23), .Z(n24) );
  IVI U36 ( .A(sel), .Z(n30) );
  IVI U37 ( .A(n33), .Z(n25) );
  IVI U38 ( .A(n30), .Z(n26) );
  IVI U39 ( .A(n33), .Z(n27) );
  IVI U40 ( .A(n33), .Z(n31) );
  MUX21L U41 ( .A(n28), .B(n29), .S(n18), .Z(out[9]) );
  IVI U42 ( .A(sel), .Z(n33) );
  MUX21H U43 ( .A(ip0[0]), .B(ip1[0]), .S(n24), .Z(out[0]) );
  MUX21H U44 ( .A(ip0[1]), .B(ip1[1]), .S(n24), .Z(out[1]) );
  MUX21H U45 ( .A(ip0[2]), .B(ip1[2]), .S(n25), .Z(out[2]) );
  MUX21H U46 ( .A(ip0[3]), .B(ip1[3]), .S(n18), .Z(out[3]) );
  MUX21H U47 ( .A(ip0[5]), .B(ip1[5]), .S(n27), .Z(out[5]) );
  MUX21H U48 ( .A(ip0[6]), .B(ip1[6]), .S(n16), .Z(out[6]) );
  MUX21H U49 ( .A(ip0[7]), .B(ip1[7]), .S(n31), .Z(out[7]) );
  MUX21H U50 ( .A(ip0[8]), .B(ip1[8]), .S(n24), .Z(out[8]) );
  MUX21H U51 ( .A(ip0[10]), .B(ip1[10]), .S(n26), .Z(out[10]) );
  MUX21H U52 ( .A(ip0[12]), .B(ip1[12]), .S(n16), .Z(out[12]) );
  MUX21H U53 ( .A(ip0[14]), .B(ip1[14]), .S(n25), .Z(out[14]) );
  MUX21H U54 ( .A(ip0[15]), .B(ip1[15]), .S(n31), .Z(out[15]) );
  MUX21H U55 ( .A(ip0[16]), .B(ip1[16]), .S(n32), .Z(out[16]) );
  MUX21H U56 ( .A(ip0[18]), .B(ip1[18]), .S(n13), .Z(out[18]) );
  MUX21H U57 ( .A(ip0[19]), .B(ip1[19]), .S(n27), .Z(out[19]) );
  MUX21H U58 ( .A(ip0[20]), .B(ip1[20]), .S(n25), .Z(out[20]) );
  MUX21H U59 ( .A(ip0[22]), .B(ip1[22]), .S(n15), .Z(out[22]) );
  MUX21H U60 ( .A(ip0[25]), .B(ip1[25]), .S(n13), .Z(out[25]) );
  MUX21H U61 ( .A(ip0[26]), .B(ip1[26]), .S(n26), .Z(out[26]) );
  MUX21H U62 ( .A(ip0[28]), .B(ip1[28]), .S(n26), .Z(out[28]) );
  MUX21H U63 ( .A(ip0[29]), .B(ip1[29]), .S(n18), .Z(out[29]) );
  MUX21H U64 ( .A(ip0[30]), .B(ip1[30]), .S(n16), .Z(out[30]) );
  MUX21H U65 ( .A(ip0[31]), .B(ip1[31]), .S(n17), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_11 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4, n6, n7, n9, n10, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59;

  B2I U1 ( .A(n35), .Z1(n1), .Z2(n2) );
  B2I U2 ( .A(n35), .Z1(n3), .Z2(n4) );
  B5IP U3 ( .A(n14), .Z(n30) );
  B4IP U4 ( .A(n31), .Z(n33) );
  ND2I U5 ( .A(n6), .B(n7), .Z(out[7]) );
  ND2I U6 ( .A(ip0[7]), .B(n36), .Z(n6) );
  ND2I U7 ( .A(ip1[7]), .B(n33), .Z(n7) );
  ND2I U8 ( .A(n9), .B(n10), .Z(out[2]) );
  ND2I U9 ( .A(ip0[2]), .B(n31), .Z(n9) );
  ND2I U10 ( .A(ip1[2]), .B(n33), .Z(n10) );
  ND2I U11 ( .A(n17), .B(n18), .Z(out[15]) );
  ND2I U12 ( .A(n15), .B(n16), .Z(out[8]) );
  ND2I U13 ( .A(n19), .B(n20), .Z(out[10]) );
  IVI U14 ( .A(n35), .Z(n14) );
  ND2I U15 ( .A(ip0[8]), .B(n36), .Z(n15) );
  ND2I U16 ( .A(ip1[8]), .B(n33), .Z(n16) );
  ND2I U17 ( .A(ip0[15]), .B(n4), .Z(n17) );
  ND2I U18 ( .A(ip1[15]), .B(n14), .Z(n18) );
  AO2P U19 ( .A(ip0[19]), .B(n30), .C(ip1[19]), .D(n33), .Z(n47) );
  AO2P U20 ( .A(ip0[26]), .B(n2), .C(ip1[26]), .D(n33), .Z(n54) );
  ND2I U21 ( .A(ip0[10]), .B(n31), .Z(n19) );
  ND2I U22 ( .A(ip1[10]), .B(n33), .Z(n20) );
  AO2P U23 ( .A(ip0[16]), .B(n4), .C(ip1[16]), .D(n3), .Z(n44) );
  AO2P U24 ( .A(ip0[11]), .B(n2), .C(ip1[11]), .D(n34), .Z(n41) );
  AO2P U25 ( .A(ip0[6]), .B(n35), .C(ip1[6]), .D(n32), .Z(n39) );
  ND2I U26 ( .A(n23), .B(n24), .Z(out[14]) );
  MUX21LP U27 ( .A(ip0[17]), .B(ip1[17]), .S(n32), .Z(n45) );
  MUX21LP U28 ( .A(ip0[20]), .B(ip1[20]), .S(n14), .Z(n48) );
  ND2I U29 ( .A(n26), .B(n27), .Z(out[0]) );
  ND2I U30 ( .A(n21), .B(n22), .Z(out[1]) );
  AO2P U31 ( .A(ip0[13]), .B(n4), .C(ip1[13]), .D(n34), .Z(n43) );
  AO2P U32 ( .A(ip0[30]), .B(n30), .C(ip1[30]), .D(n33), .Z(n58) );
  AO2P U33 ( .A(ip0[28]), .B(n30), .C(ip1[28]), .D(n14), .Z(n56) );
  AO2P U34 ( .A(ip0[25]), .B(n2), .C(ip1[25]), .D(n34), .Z(n53) );
  AO2P U35 ( .A(ip0[18]), .B(n30), .C(ip1[18]), .D(n33), .Z(n46) );
  AO2P U36 ( .A(ip0[12]), .B(n4), .C(ip1[12]), .D(n34), .Z(n42) );
  AO2P U37 ( .A(ip0[5]), .B(n30), .C(ip1[5]), .D(n25), .Z(n38) );
  AO2P U38 ( .A(ip0[29]), .B(n30), .C(ip1[29]), .D(n33), .Z(n57) );
  ND2I U39 ( .A(ip0[1]), .B(n35), .Z(n21) );
  ND2I U40 ( .A(ip1[1]), .B(n3), .Z(n22) );
  AO2P U41 ( .A(ip0[31]), .B(n2), .C(ip1[31]), .D(n33), .Z(n59) );
  AO2P U42 ( .A(ip0[27]), .B(n2), .C(ip1[27]), .D(n33), .Z(n55) );
  ND2I U43 ( .A(ip0[14]), .B(n4), .Z(n23) );
  ND2I U44 ( .A(ip1[14]), .B(n1), .Z(n24) );
  IVI U45 ( .A(n36), .Z(n25) );
  AO2P U46 ( .A(ip0[22]), .B(n2), .C(ip1[22]), .D(n33), .Z(n50) );
  AO2P U47 ( .A(ip0[24]), .B(n2), .C(ip1[24]), .D(n25), .Z(n52) );
  AO2P U48 ( .A(ip0[23]), .B(n2), .C(ip1[23]), .D(n34), .Z(n51) );
  AO2P U49 ( .A(ip0[21]), .B(n30), .C(ip1[21]), .D(n33), .Z(n49) );
  ND2I U50 ( .A(ip0[0]), .B(n31), .Z(n26) );
  ND2I U51 ( .A(ip1[0]), .B(n1), .Z(n27) );
  IVI U52 ( .A(sel), .Z(n31) );
  AO2P U53 ( .A(ip0[3]), .B(n4), .C(ip1[3]), .D(n25), .Z(n37) );
  IVI U54 ( .A(ip0[4]), .Z(n29) );
  AO2P U55 ( .A(ip0[9]), .B(n30), .C(ip1[9]), .D(n32), .Z(n40) );
  EON1P U56 ( .A(n29), .B(n25), .C(ip1[4]), .D(n32), .Z(out[4]) );
  IVI U57 ( .A(n36), .Z(n32) );
  IVI U58 ( .A(n31), .Z(n34) );
  IVI U59 ( .A(sel), .Z(n35) );
  IVI U60 ( .A(sel), .Z(n36) );
  IVI U61 ( .A(n37), .Z(out[3]) );
  IVI U62 ( .A(n38), .Z(out[5]) );
  IVI U63 ( .A(n39), .Z(out[6]) );
  IVI U64 ( .A(n40), .Z(out[9]) );
  IVI U65 ( .A(n41), .Z(out[11]) );
  IVI U66 ( .A(n42), .Z(out[12]) );
  IVI U67 ( .A(n43), .Z(out[13]) );
  IVI U68 ( .A(n44), .Z(out[16]) );
  IVI U69 ( .A(n45), .Z(out[17]) );
  IVI U70 ( .A(n46), .Z(out[18]) );
  IVI U71 ( .A(n47), .Z(out[19]) );
  IVI U72 ( .A(n48), .Z(out[20]) );
  IVI U73 ( .A(n49), .Z(out[21]) );
  IVI U74 ( .A(n50), .Z(out[22]) );
  IVI U75 ( .A(n51), .Z(out[23]) );
  IVI U76 ( .A(n52), .Z(out[24]) );
  IVI U77 ( .A(n53), .Z(out[25]) );
  IVI U78 ( .A(n54), .Z(out[26]) );
  IVI U79 ( .A(n55), .Z(out[27]) );
  IVI U80 ( .A(n56), .Z(out[28]) );
  IVI U81 ( .A(n57), .Z(out[29]) );
  IVI U82 ( .A(n58), .Z(out[30]) );
  IVI U83 ( .A(n59), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_10 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34;

  IVI U1 ( .A(ip1[16]), .Z(n2) );
  IVI U2 ( .A(ip0[14]), .Z(n3) );
  IVI U3 ( .A(ip1[14]), .Z(n4) );
  IVI U4 ( .A(ip0[29]), .Z(n5) );
  IVI U5 ( .A(ip1[29]), .Z(n6) );
  IVI U6 ( .A(ip0[16]), .Z(n1) );
  MUX21L U7 ( .A(n1), .B(n2), .S(n32), .Z(out[16]) );
  MUX21L U8 ( .A(n3), .B(n4), .S(n29), .Z(out[14]) );
  MUX21L U9 ( .A(n5), .B(n6), .S(n32), .Z(out[29]) );
  IVI U10 ( .A(ip1[24]), .Z(n18) );
  IVI U11 ( .A(ip0[1]), .Z(n9) );
  IVI U12 ( .A(ip1[1]), .Z(n10) );
  IVI U13 ( .A(ip0[3]), .Z(n13) );
  IVI U14 ( .A(ip1[3]), .Z(n14) );
  IVI U15 ( .A(ip0[26]), .Z(n7) );
  IVI U16 ( .A(ip1[26]), .Z(n8) );
  IVI U17 ( .A(ip1[27]), .Z(n16) );
  IVI U18 ( .A(ip0[27]), .Z(n15) );
  IVI U19 ( .A(ip0[28]), .Z(n26) );
  IVI U20 ( .A(ip1[28]), .Z(n27) );
  IVI U21 ( .A(ip1[31]), .Z(n20) );
  IVI U22 ( .A(ip0[31]), .Z(n19) );
  IVI U23 ( .A(ip0[30]), .Z(n24) );
  IVI U24 ( .A(ip1[30]), .Z(n25) );
  IVI U25 ( .A(ip0[24]), .Z(n17) );
  MUX21L U26 ( .A(n7), .B(n8), .S(n32), .Z(out[26]) );
  MUX21L U27 ( .A(n9), .B(n10), .S(n32), .Z(out[1]) );
  IVI U28 ( .A(n34), .Z(n11) );
  IVI U29 ( .A(sel), .Z(n12) );
  MUX21L U30 ( .A(n13), .B(n14), .S(n30), .Z(out[3]) );
  MUX21L U31 ( .A(n15), .B(n16), .S(n33), .Z(out[27]) );
  MUX21L U32 ( .A(n17), .B(n18), .S(n33), .Z(out[24]) );
  MUX21L U33 ( .A(n19), .B(n20), .S(n11), .Z(out[31]) );
  IVI U34 ( .A(n12), .Z(n21) );
  IVI U35 ( .A(n31), .Z(n22) );
  IVI U36 ( .A(n12), .Z(n23) );
  MUX21L U37 ( .A(n24), .B(n25), .S(n32), .Z(out[30]) );
  MUX21L U38 ( .A(n26), .B(n27), .S(n32), .Z(out[28]) );
  IVI U39 ( .A(n12), .Z(n28) );
  IVI U40 ( .A(n34), .Z(n29) );
  IVI U41 ( .A(n34), .Z(n30) );
  IVI U42 ( .A(sel), .Z(n34) );
  B2IP U43 ( .A(sel), .Z1(n31), .Z2(n32) );
  IVI U44 ( .A(n34), .Z(n33) );
  MUX21H U45 ( .A(ip1[7]), .B(ip0[7]), .S(n31), .Z(out[7]) );
  MUX21H U46 ( .A(ip0[0]), .B(ip1[0]), .S(n23), .Z(out[0]) );
  MUX21H U47 ( .A(ip0[2]), .B(ip1[2]), .S(n21), .Z(out[2]) );
  MUX21H U48 ( .A(ip0[4]), .B(ip1[4]), .S(n21), .Z(out[4]) );
  MUX21H U49 ( .A(ip0[5]), .B(ip1[5]), .S(n22), .Z(out[5]) );
  MUX21H U50 ( .A(ip0[6]), .B(ip1[6]), .S(n33), .Z(out[6]) );
  MUX21H U51 ( .A(ip0[8]), .B(ip1[8]), .S(n32), .Z(out[8]) );
  MUX21H U52 ( .A(ip0[9]), .B(ip1[9]), .S(n29), .Z(out[9]) );
  MUX21H U53 ( .A(ip0[10]), .B(ip1[10]), .S(n11), .Z(out[10]) );
  MUX21H U54 ( .A(ip0[11]), .B(ip1[11]), .S(n32), .Z(out[11]) );
  MUX21H U55 ( .A(ip0[12]), .B(ip1[12]), .S(n28), .Z(out[12]) );
  MUX21H U56 ( .A(ip0[13]), .B(ip1[13]), .S(n32), .Z(out[13]) );
  MUX21H U57 ( .A(ip0[15]), .B(ip1[15]), .S(n28), .Z(out[15]) );
  MUX21H U58 ( .A(ip0[17]), .B(ip1[17]), .S(n28), .Z(out[17]) );
  MUX21H U59 ( .A(ip0[18]), .B(ip1[18]), .S(n11), .Z(out[18]) );
  MUX21H U60 ( .A(ip0[19]), .B(ip1[19]), .S(n32), .Z(out[19]) );
  MUX21H U61 ( .A(ip0[20]), .B(ip1[20]), .S(n30), .Z(out[20]) );
  MUX21H U62 ( .A(ip0[21]), .B(ip1[21]), .S(n32), .Z(out[21]) );
  MUX21H U63 ( .A(ip0[22]), .B(ip1[22]), .S(n28), .Z(out[22]) );
  MUX21H U64 ( .A(ip0[23]), .B(ip1[23]), .S(n32), .Z(out[23]) );
  MUX21H U65 ( .A(ip0[25]), .B(ip1[25]), .S(n32), .Z(out[25]) );
endmodule


module mux_2x1_DATA_WIDTH32_9 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  MUX21L U1 ( .A(n18), .B(n19), .S(n2), .Z(out[14]) );
  B2IP U2 ( .A(sel), .Z2(n1) );
  B2IP U3 ( .A(sel), .Z2(n2) );
  IVI U4 ( .A(ip0[9]), .Z(n20) );
  IVI U5 ( .A(n27), .Z(out[12]) );
  MUX21L U6 ( .A(ip0[12]), .B(ip1[12]), .S(n2), .Z(n27) );
  IVI U7 ( .A(ip0[14]), .Z(n18) );
  IVI U8 ( .A(ip0[10]), .Z(n3) );
  IVI U9 ( .A(n25), .Z(out[18]) );
  MUX21L U10 ( .A(ip0[18]), .B(ip1[18]), .S(n1), .Z(n25) );
  IVI U11 ( .A(n24), .Z(out[20]) );
  MUX21L U12 ( .A(ip0[20]), .B(ip1[20]), .S(n1), .Z(n24) );
  IVI U13 ( .A(n23), .Z(out[22]) );
  MUX21L U14 ( .A(ip0[22]), .B(ip1[22]), .S(n1), .Z(n23) );
  MUX21L U15 ( .A(ip0[23]), .B(ip1[23]), .S(n1), .Z(n9) );
  MUX21L U16 ( .A(ip0[19]), .B(ip1[19]), .S(n1), .Z(n11) );
  MUX21L U17 ( .A(ip0[16]), .B(ip1[16]), .S(n2), .Z(n12) );
  MUX21LP U18 ( .A(ip0[1]), .B(ip1[1]), .S(n1), .Z(n17) );
  MUX21L U19 ( .A(ip0[5]), .B(ip1[5]), .S(n2), .Z(n28) );
  IVI U20 ( .A(n9), .Z(out[23]) );
  IVI U21 ( .A(n10), .Z(out[21]) );
  MUX21L U22 ( .A(ip0[21]), .B(ip1[21]), .S(n1), .Z(n10) );
  IVI U23 ( .A(n11), .Z(out[19]) );
  IVI U24 ( .A(n12), .Z(out[16]) );
  IVI U25 ( .A(n28), .Z(out[5]) );
  IVI U26 ( .A(n7), .Z(out[15]) );
  MUX21L U27 ( .A(ip0[15]), .B(ip1[15]), .S(n2), .Z(n7) );
  MUX21L U28 ( .A(ip0[17]), .B(ip1[17]), .S(n2), .Z(n26) );
  MUX21L U29 ( .A(ip0[8]), .B(ip1[8]), .S(n2), .Z(n15) );
  MUX21L U30 ( .A(ip0[11]), .B(ip1[11]), .S(n2), .Z(n14) );
  MUX21L U31 ( .A(ip0[13]), .B(ip1[13]), .S(n2), .Z(n13) );
  IVI U32 ( .A(n26), .Z(out[17]) );
  IVI U33 ( .A(n5), .Z(out[30]) );
  MUX21L U34 ( .A(ip0[30]), .B(ip1[30]), .S(n1), .Z(n5) );
  IVI U35 ( .A(n6), .Z(out[28]) );
  MUX21L U36 ( .A(ip0[28]), .B(ip1[28]), .S(n1), .Z(n6) );
  IVI U37 ( .A(ip1[10]), .Z(n4) );
  IVI U38 ( .A(n8), .Z(out[26]) );
  MUX21L U39 ( .A(ip0[26]), .B(ip1[26]), .S(n1), .Z(n8) );
  IVI U40 ( .A(n14), .Z(out[11]) );
  IVI U41 ( .A(n15), .Z(out[8]) );
  IVI U42 ( .A(n13), .Z(out[13]) );
  MUX21LP U43 ( .A(n3), .B(n4), .S(n2), .Z(out[10]) );
  IVI U44 ( .A(n16), .Z(out[25]) );
  MUX21L U45 ( .A(ip0[25]), .B(ip1[25]), .S(n1), .Z(n16) );
  MUX21L U46 ( .A(ip0[29]), .B(ip1[29]), .S(n1), .Z(n22) );
  IVI U47 ( .A(n22), .Z(out[29]) );
  IVI U48 ( .A(n17), .Z(out[1]) );
  IVI U49 ( .A(ip1[14]), .Z(n19) );
  IVI U50 ( .A(ip1[9]), .Z(n21) );
  MUX21LP U51 ( .A(n20), .B(n21), .S(n2), .Z(out[9]) );
  MUX21H U52 ( .A(ip0[0]), .B(ip1[0]), .S(n1), .Z(out[0]) );
  MUX21H U53 ( .A(ip0[2]), .B(ip1[2]), .S(n1), .Z(out[2]) );
  MUX21H U54 ( .A(ip0[3]), .B(ip1[3]), .S(n1), .Z(out[3]) );
  MUX21H U55 ( .A(ip0[4]), .B(ip1[4]), .S(n2), .Z(out[4]) );
  MUX21H U56 ( .A(ip0[6]), .B(ip1[6]), .S(n2), .Z(out[6]) );
  MUX21H U57 ( .A(ip0[7]), .B(ip1[7]), .S(n2), .Z(out[7]) );
  MUX21H U58 ( .A(ip0[24]), .B(ip1[24]), .S(n1), .Z(out[24]) );
  MUX21H U59 ( .A(ip0[27]), .B(ip1[27]), .S(n1), .Z(out[27]) );
  MUX21H U60 ( .A(ip0[31]), .B(ip1[31]), .S(n1), .Z(out[31]) );
endmodule


module pc_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n4, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n26, n27, n28, n29, n30, n31, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n85, n86, n89, n90, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n106, n107,
         n108, n109, n110, n113, n115, n116, n117, n118, n119, n120, n121,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n149,
         n150, n151, n152, n153, n154, n155, n157, n158, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n216, n217, n220, n221, n222, n223, n224,
         n225, n226, n228, n229, n230, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n260, n261,
         n262, n264, n267, n268, n269, n270, n271, n272, n273, n274, n277,
         n279, n280, n281, n384, n385, n386, n387, n389, n390, n391, n392,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n404, n405,
         n406, n407, n408, n409, n410, n411, n412;

  MUX21LP U9 ( .A(n9), .B(n10), .S(n412), .Z(SUM[31]) );
  EOI U16 ( .A(n26), .B(n17), .Z(n15) );
  EOI U17 ( .A(n17), .B(n27), .Z(n16) );
  ENI U18 ( .A(B[31]), .B(A[31]), .Z(n17) );
  ENI U24 ( .A(n36), .B(n407), .Z(n22) );
  ENI U25 ( .A(n37), .B(n407), .Z(n23) );
  NR2I U28 ( .A(B[30]), .B(A[30]), .Z(n26) );
  ND2I U29 ( .A(B[30]), .B(A[30]), .Z(n27) );
  MUX21LP U30 ( .A(n28), .B(n29), .S(n410), .Z(SUM[29]) );
  ENI U41 ( .A(B[29]), .B(A[29]), .Z(n38) );
  NR2I U42 ( .A(B[29]), .B(A[29]), .Z(n39) );
  ND2I U43 ( .A(B[29]), .B(A[29]), .Z(n40) );
  EOI U47 ( .A(n54), .B(n45), .Z(n43) );
  EOI U48 ( .A(n55), .B(n45), .Z(n44) );
  ENI U49 ( .A(B[28]), .B(A[28]), .Z(n45) );
  NR2I U50 ( .A(B[28]), .B(A[28]), .Z(n46) );
  ND2I U51 ( .A(B[28]), .B(A[28]), .Z(n47) );
  EOI U61 ( .A(n68), .B(n60), .Z(n56) );
  EOI U62 ( .A(n60), .B(n69), .Z(n57) );
  ENI U65 ( .A(B[27]), .B(A[27]), .Z(n60) );
  NR2I U66 ( .A(B[27]), .B(A[27]), .Z(n61) );
  ND2I U67 ( .A(B[27]), .B(A[27]), .Z(n62) );
  EOI U71 ( .A(n72), .B(n67), .Z(n65) );
  ENI U73 ( .A(B[26]), .B(A[26]), .Z(n67) );
  NR2I U74 ( .A(B[26]), .B(A[26]), .Z(n68) );
  ND2I U75 ( .A(B[26]), .B(A[26]), .Z(n69) );
  EOI U81 ( .A(n85), .B(n78), .Z(n74) );
  EOI U82 ( .A(n78), .B(n86), .Z(n75) );
  MUX21LP U83 ( .A(n79), .B(n80), .S(n85), .Z(n76) );
  MUX21LP U84 ( .A(n79), .B(n80), .S(n86), .Z(n77) );
  ENI U85 ( .A(B[25]), .B(A[25]), .Z(n78) );
  NR2I U86 ( .A(B[25]), .B(A[25]), .Z(n79) );
  ND2I U87 ( .A(B[25]), .B(A[25]), .Z(n80) );
  ENI U89 ( .A(n8), .B(n390), .Z(n81) );
  ENI U90 ( .A(n6), .B(n390), .Z(n82) );
  NR2I U93 ( .A(B[24]), .B(A[24]), .Z(n85) );
  ND2I U94 ( .A(B[24]), .B(A[24]), .Z(n86) );
  MUX21LP U101 ( .A(n95), .B(n96), .S(n133), .Z(n6) );
  MUX21LP U104 ( .A(n100), .B(n99), .S(n117), .Z(n95) );
  MUX21LP U105 ( .A(n100), .B(n99), .S(n118), .Z(n96) );
  EOI U106 ( .A(n109), .B(n101), .Z(n97) );
  EOI U107 ( .A(n101), .B(n110), .Z(n98) );
  MUX21LP U108 ( .A(n102), .B(n103), .S(n109), .Z(n99) );
  MUX21LP U109 ( .A(n102), .B(n103), .S(n110), .Z(n100) );
  ENI U110 ( .A(B[23]), .B(A[23]), .Z(n101) );
  NR2I U111 ( .A(B[23]), .B(A[23]), .Z(n102) );
  ND2I U112 ( .A(B[23]), .B(A[23]), .Z(n103) );
  EOI U116 ( .A(n113), .B(n108), .Z(n106) );
  ENI U118 ( .A(B[22]), .B(A[22]), .Z(n108) );
  NR2I U119 ( .A(B[22]), .B(A[22]), .Z(n109) );
  ND2I U120 ( .A(B[22]), .B(A[22]), .Z(n110) );
  EOI U126 ( .A(n126), .B(n119), .Z(n115) );
  EOI U127 ( .A(n119), .B(n127), .Z(n116) );
  MUX21LP U128 ( .A(n120), .B(n121), .S(n126), .Z(n117) );
  MUX21LP U129 ( .A(n120), .B(n121), .S(n127), .Z(n118) );
  ENI U130 ( .A(B[21]), .B(A[21]), .Z(n119) );
  NR2I U131 ( .A(B[21]), .B(A[21]), .Z(n120) );
  ND2I U132 ( .A(B[21]), .B(A[21]), .Z(n121) );
  NR2I U138 ( .A(B[20]), .B(A[20]), .Z(n126) );
  ND2I U139 ( .A(B[20]), .B(A[20]), .Z(n127) );
  MUX21LP U145 ( .A(n137), .B(n136), .S(n151), .Z(n132) );
  MUX21LP U146 ( .A(n137), .B(n136), .S(n152), .Z(n133) );
  EOI U147 ( .A(n145), .B(n138), .Z(n134) );
  EOI U148 ( .A(n138), .B(n146), .Z(n135) );
  MUX21LP U149 ( .A(n139), .B(n140), .S(n145), .Z(n136) );
  MUX21LP U150 ( .A(n139), .B(n140), .S(n146), .Z(n137) );
  ENI U151 ( .A(B[19]), .B(A[19]), .Z(n138) );
  NR2I U152 ( .A(B[19]), .B(A[19]), .Z(n139) );
  ND2I U153 ( .A(B[19]), .B(A[19]), .Z(n140) );
  ENI U155 ( .A(n151), .B(n143), .Z(n141) );
  ENI U156 ( .A(n152), .B(n143), .Z(n142) );
  ENI U158 ( .A(B[18]), .B(A[18]), .Z(n144) );
  NR2I U159 ( .A(B[18]), .B(A[18]), .Z(n145) );
  ND2I U160 ( .A(B[18]), .B(A[18]), .Z(n146) );
  EOI U164 ( .A(n157), .B(n153), .Z(n149) );
  EOI U165 ( .A(n153), .B(n158), .Z(n150) );
  MUX21LP U166 ( .A(n154), .B(n155), .S(n157), .Z(n151) );
  MUX21LP U167 ( .A(n154), .B(n155), .S(n158), .Z(n152) );
  ENI U168 ( .A(B[17]), .B(A[17]), .Z(n153) );
  NR2I U169 ( .A(B[17]), .B(A[17]), .Z(n154) );
  ND2I U170 ( .A(B[17]), .B(A[17]), .Z(n155) );
  NR2I U173 ( .A(B[16]), .B(A[16]), .Z(n157) );
  ND2I U174 ( .A(B[16]), .B(A[16]), .Z(n158) );
  MUX21LP U176 ( .A(n163), .B(n162), .S(n232), .Z(n4) );
  MUX21LP U183 ( .A(n171), .B(n170), .S(n188), .Z(n166) );
  EOI U185 ( .A(n172), .B(n180), .Z(n168) );
  EOI U186 ( .A(n172), .B(n181), .Z(n169) );
  MUX21LP U187 ( .A(n173), .B(n174), .S(n180), .Z(n170) );
  MUX21LP U188 ( .A(n173), .B(n174), .S(n181), .Z(n171) );
  EOI U189 ( .A(B[15]), .B(A[15]), .Z(n172) );
  NR2I U190 ( .A(B[15]), .B(A[15]), .Z(n173) );
  ND2I U191 ( .A(B[15]), .B(A[15]), .Z(n174) );
  EOI U195 ( .A(n184), .B(n179), .Z(n177) );
  ENI U197 ( .A(B[14]), .B(A[14]), .Z(n179) );
  NR2I U198 ( .A(B[14]), .B(A[14]), .Z(n180) );
  ND2I U199 ( .A(B[14]), .B(A[14]), .Z(n181) );
  EOI U205 ( .A(n197), .B(n190), .Z(n186) );
  EOI U206 ( .A(n190), .B(n198), .Z(n187) );
  MUX21LP U207 ( .A(n191), .B(n192), .S(n197), .Z(n188) );
  MUX21LP U208 ( .A(n191), .B(n192), .S(n198), .Z(n189) );
  ENI U209 ( .A(B[13]), .B(A[13]), .Z(n190) );
  NR2I U210 ( .A(B[13]), .B(A[13]), .Z(n191) );
  ND2I U211 ( .A(B[13]), .B(A[13]), .Z(n192) );
  ENI U213 ( .A(n199), .B(n392), .Z(n193) );
  ENI U214 ( .A(n200), .B(n392), .Z(n194) );
  NR2I U217 ( .A(B[12]), .B(A[12]), .Z(n197) );
  ND2I U218 ( .A(B[12]), .B(A[12]), .Z(n198) );
  MUX21LP U225 ( .A(n208), .B(n207), .S(n223), .Z(n204) );
  EOI U226 ( .A(n216), .B(n209), .Z(n205) );
  EOI U227 ( .A(n209), .B(n217), .Z(n206) );
  MUX21LP U228 ( .A(n210), .B(n211), .S(n216), .Z(n207) );
  MUX21LP U229 ( .A(n210), .B(n211), .S(n217), .Z(n208) );
  ENI U230 ( .A(B[11]), .B(A[11]), .Z(n209) );
  NR2I U231 ( .A(B[11]), .B(A[11]), .Z(n210) );
  ND2I U232 ( .A(B[11]), .B(A[11]), .Z(n211) );
  ENI U234 ( .A(n222), .B(n391), .Z(n212) );
  ENI U235 ( .A(n223), .B(n391), .Z(n213) );
  NR2I U238 ( .A(B[10]), .B(A[10]), .Z(n216) );
  ND2I U239 ( .A(B[10]), .B(A[10]), .Z(n217) );
  EOI U243 ( .A(n228), .B(n224), .Z(n220) );
  EOI U244 ( .A(n224), .B(n229), .Z(n221) );
  MUX21LP U245 ( .A(n225), .B(n226), .S(n228), .Z(n222) );
  MUX21LP U246 ( .A(n225), .B(n226), .S(n229), .Z(n223) );
  ENI U247 ( .A(B[9]), .B(A[9]), .Z(n224) );
  NR2I U248 ( .A(B[9]), .B(A[9]), .Z(n225) );
  ND2I U249 ( .A(B[9]), .B(A[9]), .Z(n226) );
  NR2I U252 ( .A(B[8]), .B(A[8]), .Z(n228) );
  ND2I U253 ( .A(B[8]), .B(A[8]), .Z(n229) );
  MUX21LP U257 ( .A(n235), .B(n236), .S(n264), .Z(n232) );
  EOI U262 ( .A(n241), .B(n247), .Z(n237) );
  EOI U263 ( .A(n241), .B(n248), .Z(n238) );
  MUX21LP U264 ( .A(n242), .B(n243), .S(n247), .Z(n239) );
  MUX21LP U265 ( .A(n242), .B(n243), .S(n248), .Z(n240) );
  EOI U266 ( .A(B[7]), .B(A[7]), .Z(n241) );
  NR2I U267 ( .A(B[7]), .B(A[7]), .Z(n242) );
  ND2I U268 ( .A(B[7]), .B(A[7]), .Z(n243) );
  EOI U270 ( .A(n249), .B(n246), .Z(n244) );
  EOI U271 ( .A(n250), .B(n246), .Z(n245) );
  EOI U272 ( .A(B[6]), .B(A[6]), .Z(n246) );
  NR2I U273 ( .A(B[6]), .B(A[6]), .Z(n247) );
  ND2I U274 ( .A(B[6]), .B(A[6]), .Z(n248) );
  EOI U278 ( .A(n255), .B(n260), .Z(n251) );
  EOI U279 ( .A(n255), .B(n261), .Z(n252) );
  MUX21LP U280 ( .A(n256), .B(n257), .S(n260), .Z(n253) );
  MUX21LP U281 ( .A(n256), .B(n257), .S(n261), .Z(n254) );
  EOI U282 ( .A(B[5]), .B(A[5]), .Z(n255) );
  NR2I U283 ( .A(B[5]), .B(A[5]), .Z(n256) );
  ND2I U284 ( .A(B[5]), .B(A[5]), .Z(n257) );
  ENI U285 ( .A(n262), .B(n408), .Z(SUM[4]) );
  NR2I U288 ( .A(B[4]), .B(A[4]), .Z(n260) );
  ND2I U289 ( .A(B[4]), .B(A[4]), .Z(n261) );
  MUX21LP U293 ( .A(n268), .B(n267), .S(n277), .Z(n264) );
  ENI U298 ( .A(B[3]), .B(A[3]), .Z(n269) );
  NR2I U299 ( .A(B[3]), .B(A[3]), .Z(n270) );
  ND2I U300 ( .A(B[3]), .B(A[3]), .Z(n271) );
  ENI U302 ( .A(B[2]), .B(A[2]), .Z(n272) );
  NR2I U303 ( .A(B[2]), .B(A[2]), .Z(n273) );
  ND2I U304 ( .A(B[2]), .B(A[2]), .Z(n274) );
  NR2I U310 ( .A(A[1]), .B(B[1]), .Z(n279) );
  ND2I U311 ( .A(A[1]), .B(B[1]), .Z(n280) );
  EOI U312 ( .A(A[0]), .B(B[0]), .Z(SUM[0]) );
  ND2I U313 ( .A(A[0]), .B(B[0]), .Z(n281) );
  IVDAP U317 ( .A(n4), .Y(n400), .Z(n412) );
  EOI U318 ( .A(n128), .B(n389), .Z(n384) );
  EOI U319 ( .A(n129), .B(n389), .Z(n385) );
  MUX21H U320 ( .A(n57), .B(n56), .S(n76), .Z(n386) );
  MUX21H U321 ( .A(n57), .B(n56), .S(n77), .Z(n387) );
  MUX21H U322 ( .A(n233), .B(n234), .S(n264), .Z(SUM[7]) );
  EOI U323 ( .A(B[20]), .B(A[20]), .Z(n389) );
  EOI U324 ( .A(B[24]), .B(A[24]), .Z(n390) );
  EOI U325 ( .A(B[10]), .B(A[10]), .Z(n391) );
  EOI U326 ( .A(B[12]), .B(A[12]), .Z(n392) );
  EOI U327 ( .A(n409), .B(n281), .Z(SUM[1]) );
  B2IP U328 ( .A(n4), .Z1(n396), .Z2(n411) );
  MUX21LP U329 ( .A(n95), .B(n96), .S(n132), .Z(n8) );
  MUX21LP U330 ( .A(n59), .B(n58), .S(n77), .Z(n55) );
  MUX21LP U331 ( .A(n59), .B(n58), .S(n76), .Z(n54) );
  MUX21LP U332 ( .A(n208), .B(n207), .S(n222), .Z(n203) );
  MUX21LP U333 ( .A(n171), .B(n170), .S(n189), .Z(n167) );
  MUX21H U334 ( .A(n394), .B(n395), .S(n396), .Z(SUM[21]) );
  MUX21H U335 ( .A(n116), .B(n115), .S(n129), .Z(n394) );
  MUX21H U336 ( .A(n116), .B(n115), .S(n128), .Z(n395) );
  MUX21H U337 ( .A(n385), .B(n384), .S(n400), .Z(SUM[20]) );
  ENI U338 ( .A(n400), .B(n397), .Z(SUM[16]) );
  ENI U339 ( .A(B[16]), .B(A[16]), .Z(n397) );
  MUX21L U340 ( .A(n21), .B(n20), .S(n6), .Z(n19) );
  MUX21L U341 ( .A(n21), .B(n20), .S(n8), .Z(n18) );
  MUX21L U342 ( .A(n31), .B(n30), .S(n6), .Z(n29) );
  MUX21L U343 ( .A(n31), .B(n30), .S(n8), .Z(n28) );
  MUX21L U344 ( .A(n12), .B(n11), .S(n6), .Z(n10) );
  MUX21L U345 ( .A(n12), .B(n11), .S(n8), .Z(n9) );
  MUX21L U346 ( .A(n48), .B(n49), .S(n411), .Z(SUM[27]) );
  MUX21L U347 ( .A(n387), .B(n386), .S(n8), .Z(n48) );
  MUX21L U348 ( .A(n387), .B(n386), .S(n6), .Z(n49) );
  MUX21H U349 ( .A(n89), .B(n90), .S(n410), .Z(SUM[23]) );
  MUX21L U350 ( .A(n93), .B(n94), .S(n132), .Z(n89) );
  MUX21L U351 ( .A(n93), .B(n94), .S(n133), .Z(n90) );
  MUX21L U352 ( .A(n44), .B(n43), .S(n6), .Z(n42) );
  MUX21L U353 ( .A(n44), .B(n43), .S(n8), .Z(n41) );
  MUX21L U354 ( .A(n22), .B(n23), .S(n55), .Z(n21) );
  MUX21L U355 ( .A(n402), .B(n401), .S(n55), .Z(n31) );
  MUX21L U356 ( .A(n13), .B(n14), .S(n55), .Z(n12) );
  MUX21L U357 ( .A(n22), .B(n23), .S(n54), .Z(n20) );
  MUX21L U358 ( .A(n402), .B(n401), .S(n54), .Z(n30) );
  MUX21L U359 ( .A(n13), .B(n14), .S(n54), .Z(n11) );
  MUX21L U360 ( .A(n166), .B(n167), .S(n203), .Z(n162) );
  MUX21L U361 ( .A(n166), .B(n167), .S(n204), .Z(n163) );
  MUX21L U362 ( .A(n98), .B(n97), .S(n118), .Z(n94) );
  MUX21L U363 ( .A(n98), .B(n97), .S(n117), .Z(n93) );
  MUX21L U364 ( .A(n169), .B(n168), .S(n189), .Z(n165) );
  MUX21L U365 ( .A(n161), .B(n160), .S(n232), .Z(SUM[15]) );
  MUX21L U366 ( .A(n164), .B(n165), .S(n203), .Z(n160) );
  MUX21L U367 ( .A(n164), .B(n165), .S(n204), .Z(n161) );
  MUX21L U368 ( .A(n169), .B(n168), .S(n188), .Z(n164) );
  MUX21L U369 ( .A(n240), .B(n239), .S(n254), .Z(n236) );
  MUX21L U370 ( .A(n240), .B(n239), .S(n253), .Z(n235) );
  MUX21L U371 ( .A(n61), .B(n62), .S(n69), .Z(n59) );
  MUX21L U372 ( .A(n61), .B(n62), .S(n68), .Z(n58) );
  MUX21H U373 ( .A(n398), .B(n399), .S(n396), .Z(SUM[22]) );
  MUX21H U374 ( .A(n107), .B(n106), .S(n129), .Z(n398) );
  MUX21H U375 ( .A(n107), .B(n106), .S(n128), .Z(n399) );
  MUX21L U376 ( .A(n81), .B(n82), .S(n411), .Z(SUM[24]) );
  MUX21L U377 ( .A(n63), .B(n64), .S(n410), .Z(SUM[26]) );
  MUX21L U378 ( .A(n66), .B(n65), .S(n8), .Z(n63) );
  MUX21L U379 ( .A(n66), .B(n65), .S(n6), .Z(n64) );
  MUX21L U380 ( .A(n130), .B(n131), .S(n410), .Z(SUM[19]) );
  MUX21L U381 ( .A(n135), .B(n134), .S(n151), .Z(n130) );
  MUX21L U382 ( .A(n135), .B(n134), .S(n152), .Z(n131) );
  MUX21L U383 ( .A(n70), .B(n71), .S(n412), .Z(SUM[25]) );
  MUX21L U384 ( .A(n75), .B(n74), .S(n8), .Z(n70) );
  MUX21L U385 ( .A(n75), .B(n74), .S(n6), .Z(n71) );
  MUX21L U386 ( .A(n141), .B(n142), .S(n411), .Z(SUM[18]) );
  MUX21H U387 ( .A(n150), .B(n149), .S(n400), .Z(SUM[17]) );
  ENI U388 ( .A(n38), .B(n47), .Z(n401) );
  ENI U389 ( .A(n46), .B(n38), .Z(n402) );
  ENI U390 ( .A(n118), .B(n108), .Z(n107) );
  ENI U391 ( .A(n77), .B(n67), .Z(n66) );
  MUX21L U392 ( .A(n16), .B(n15), .S(n37), .Z(n14) );
  MUX21L U393 ( .A(n16), .B(n15), .S(n36), .Z(n13) );
  MUX21L U394 ( .A(n39), .B(n40), .S(n47), .Z(n37) );
  MUX21L U395 ( .A(n39), .B(n40), .S(n46), .Z(n36) );
  MUX21L U396 ( .A(n175), .B(n176), .S(n230), .Z(SUM[14]) );
  MUX21L U397 ( .A(n178), .B(n177), .S(n199), .Z(n175) );
  MUX21L U398 ( .A(n178), .B(n177), .S(n200), .Z(n176) );
  MUX21L U399 ( .A(n193), .B(n194), .S(n230), .Z(SUM[12]) );
  MUX21L U400 ( .A(n212), .B(n213), .S(n230), .Z(SUM[10]) );
  MUX21L U401 ( .A(n182), .B(n183), .S(n230), .Z(SUM[13]) );
  MUX21L U402 ( .A(n187), .B(n186), .S(n199), .Z(n182) );
  MUX21L U403 ( .A(n187), .B(n186), .S(n200), .Z(n183) );
  MUX21L U404 ( .A(n201), .B(n202), .S(n230), .Z(SUM[11]) );
  MUX21L U405 ( .A(n206), .B(n205), .S(n222), .Z(n201) );
  MUX21L U406 ( .A(n206), .B(n205), .S(n223), .Z(n202) );
  MUX21H U407 ( .A(n220), .B(n221), .S(n230), .Z(SUM[9]) );
  ENI U408 ( .A(n189), .B(n179), .Z(n178) );
  MUX21L U409 ( .A(n238), .B(n237), .S(n253), .Z(n233) );
  MUX21L U410 ( .A(n238), .B(n237), .S(n254), .Z(n234) );
  MUX21L U411 ( .A(n404), .B(n405), .S(n277), .Z(SUM[3]) );
  ENI U412 ( .A(n269), .B(n274), .Z(n404) );
  ENI U413 ( .A(n273), .B(n269), .Z(n405) );
  MUX21L U414 ( .A(n18), .B(n19), .S(n411), .Z(SUM[30]) );
  MUX21L U415 ( .A(n41), .B(n42), .S(n412), .Z(SUM[28]) );
  MUX21L U416 ( .A(n270), .B(n271), .S(n273), .Z(n267) );
  MUX21L U417 ( .A(n270), .B(n271), .S(n274), .Z(n268) );
  ENI U418 ( .A(n230), .B(n406), .Z(SUM[8]) );
  EOI U419 ( .A(B[8]), .B(A[8]), .Z(n406) );
  EOI U420 ( .A(B[30]), .B(A[30]), .Z(n407) );
  ENI U421 ( .A(B[4]), .B(A[4]), .Z(n408) );
  MUX21L U422 ( .A(n245), .B(n244), .S(n262), .Z(SUM[6]) );
  MUX21L U423 ( .A(n252), .B(n251), .S(n262), .Z(SUM[5]) );
  ENI U424 ( .A(A[1]), .B(B[1]), .Z(n409) );
  ENI U425 ( .A(n277), .B(n272), .Z(SUM[2]) );
  MUX21L U426 ( .A(n279), .B(n280), .S(n281), .Z(n277) );
  B2IP U427 ( .A(n4), .Z2(n410) );
  IVI U428 ( .A(n76), .Z(n72) );
  IVI U429 ( .A(n264), .Z(n262) );
  IVI U430 ( .A(n254), .Z(n250) );
  IVI U431 ( .A(n253), .Z(n249) );
  IVI U432 ( .A(n232), .Z(n230) );
  IVI U433 ( .A(n204), .Z(n200) );
  IVI U434 ( .A(n203), .Z(n199) );
  IVI U435 ( .A(n188), .Z(n184) );
  IVI U436 ( .A(n144), .Z(n143) );
  IVI U437 ( .A(n133), .Z(n129) );
  IVI U438 ( .A(n132), .Z(n128) );
  IVI U439 ( .A(n117), .Z(n113) );
endmodule


module pc_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n16, n18, n21, n23, n24, n25, n28, n30, n31,
         n32, n33, n34, n36, n37, n39, n45, n46, n47, n48, n49, n51, n53, n55,
         n57, n58, n59, n60, n64, n69, n70, n71, n72, n73, n74, n76, n77, n79,
         n81, n82, n83, n84, n85, n86, n90, n92, n93, n94, n95, n96, n97, n98,
         n102, n105, n106, n107, n110, n112, n113, n115, n116, n117, n118,
         n119, n121, n123, n125, n129, n130, n131, n132, n133, n134, n136,
         n139, n140, n141, n142, n143, n144, n145, n146, n148, n152, n153,
         n155, n157, n160, n161, n162, n163, n164, n166, n167, n170, n172,
         n174, n175, n176, n179, n181, n183, n185, n186, n187, n191, n192,
         \A[0] , \A[1] , n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n306, n308, n310;
  assign n31 = A[31];
  assign n37 = A[30];
  assign n47 = A[29];
  assign n53 = A[28];
  assign n57 = A[27];
  assign n64 = A[26];
  assign n73 = A[25];
  assign n79 = A[24];
  assign n83 = A[23];
  assign n90 = A[22];
  assign n97 = A[21];
  assign n102 = A[20];
  assign n107 = A[18];
  assign n119 = A[17];
  assign n125 = A[16];
  assign n129 = A[15];
  assign n136 = A[14];
  assign n143 = A[13];
  assign n148 = A[12];
  assign n153 = A[10];
  assign n164 = A[9];
  assign n170 = A[8];
  assign n176 = A[7];
  assign n179 = A[6];
  assign n185 = A[5];
  assign n187 = A[4];
  assign n192 = A[2];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];

  EOI U10 ( .A(n5), .B(n31), .Z(n32) );
  ENI U15 ( .A(n45), .B(n5), .Z(n36) );
  NR2I U26 ( .A(n60), .B(n48), .Z(n45) );
  ENI U27 ( .A(n53), .B(n6), .Z(n46) );
  ND2I U29 ( .A(n53), .B(n47), .Z(n48) );
  ENI U34 ( .A(n58), .B(n7), .Z(n51) );
  ENI U44 ( .A(n64), .B(n8), .Z(n59) );
  ND2I U45 ( .A(n57), .B(n64), .Z(n60) );
  ND2I U57 ( .A(n95), .B(n71), .Z(n4) );
  NR2I U60 ( .A(n86), .B(n74), .Z(n71) );
  ENI U61 ( .A(n79), .B(n70), .Z(n72) );
  ND2I U63 ( .A(n73), .B(n79), .Z(n74) );
  ENI U68 ( .A(n84), .B(n76), .Z(n77) );
  ENI U78 ( .A(n90), .B(n82), .Z(n85) );
  ND2I U79 ( .A(n83), .B(n90), .Z(n86) );
  NR2I U92 ( .A(n106), .B(n98), .Z(n95) );
  ENI U93 ( .A(n102), .B(n92), .Z(n96) );
  ND2I U95 ( .A(n97), .B(n102), .Z(n98) );
  ENI U106 ( .A(n107), .B(n16), .Z(n105) );
  ND2I U107 ( .A(A[19]), .B(n107), .Z(n106) );
  NR2I U114 ( .A(n112), .B(n157), .Z(n2) );
  ND2I U117 ( .A(n141), .B(n115), .Z(n112) );
  NR2I U120 ( .A(n132), .B(n118), .Z(n115) );
  ENI U121 ( .A(n125), .B(n119), .Z(n116) );
  ND2I U123 ( .A(n119), .B(n125), .Z(n118) );
  ENI U129 ( .A(n130), .B(n18), .Z(n123) );
  ENI U139 ( .A(n136), .B(n294), .Z(n131) );
  ND2I U140 ( .A(n129), .B(n136), .Z(n132) );
  EOI U143 ( .A(n139), .B(n136), .Z(n133) );
  NR2I U153 ( .A(n152), .B(n144), .Z(n141) );
  ENI U154 ( .A(n148), .B(n21), .Z(n142) );
  ND2I U156 ( .A(n143), .B(n148), .Z(n144) );
  EOI U159 ( .A(n152), .B(n148), .Z(n145) );
  ND2I U168 ( .A(A[11]), .B(n153), .Z(n152) );
  ENI U170 ( .A(n155), .B(n24), .Z(SUM[10]) );
  ND2I U177 ( .A(n160), .B(n183), .Z(n157) );
  NR2I U180 ( .A(n175), .B(n163), .Z(n160) );
  ENI U181 ( .A(n170), .B(n164), .Z(n161) );
  ND2I U183 ( .A(n164), .B(n170), .Z(n163) );
  ENI U196 ( .A(n179), .B(n176), .Z(n174) );
  ND2I U197 ( .A(n176), .B(n179), .Z(n175) );
  NR2I U207 ( .A(n186), .B(n191), .Z(n183) );
  ND2I U210 ( .A(n185), .B(n187), .Z(n186) );
  ND2I U219 ( .A(A[3]), .B(n192), .Z(n191) );
  MUX21L U227 ( .A(n82), .B(n81), .S(n310), .Z(SUM[23]) );
  MUX21L U228 ( .A(n21), .B(n140), .S(n155), .Z(SUM[13]) );
  MUX21L U229 ( .A(n166), .B(n167), .S(n181), .Z(SUM[8]) );
  IVDA U230 ( .A(n129), .Y(n294), .Z(n295) );
  MUX21LP U231 ( .A(n174), .B(n172), .S(n181), .Z(SUM[7]) );
  MUX21LP U232 ( .A(n162), .B(n306), .S(n183), .Z(SUM[9]) );
  MUX21LP U233 ( .A(n146), .B(n145), .S(n155), .Z(SUM[12]) );
  MUX21H U234 ( .A(n70), .B(n69), .S(n95), .Z(n296) );
  MUX21H U235 ( .A(n46), .B(n47), .S(n60), .Z(n297) );
  EOI U236 ( .A(n153), .B(n23), .Z(n298) );
  B2IP U237 ( .A(n2), .Z1(n304), .Z2(n310) );
  MUX21H U238 ( .A(n295), .B(n299), .S(n155), .Z(SUM[15]) );
  MUX21H U239 ( .A(n131), .B(n129), .S(n139), .Z(n299) );
  MUX21L U240 ( .A(n8), .B(n55), .S(n310), .Z(SUM[27]) );
  MUX21L U241 ( .A(n59), .B(n57), .S(n4), .Z(n55) );
  MUX21H U242 ( .A(n300), .B(n79), .S(n304), .Z(SUM[24]) );
  MUX21H U243 ( .A(n77), .B(n79), .S(n93), .Z(n300) );
  MUX21H U244 ( .A(n301), .B(n90), .S(n304), .Z(SUM[22]) );
  ENI U245 ( .A(n93), .B(n90), .Z(n301) );
  MUX21H U246 ( .A(n302), .B(n102), .S(n304), .Z(SUM[20]) );
  ENI U247 ( .A(n106), .B(n102), .Z(n302) );
  MUX21H U248 ( .A(n303), .B(n64), .S(n304), .Z(SUM[26]) );
  ENI U249 ( .A(n4), .B(n64), .Z(n303) );
  MUX21L U250 ( .A(n70), .B(n296), .S(n310), .Z(SUM[25]) );
  MUX21L U251 ( .A(n72), .B(n73), .S(n86), .Z(n69) );
  MUX21L U252 ( .A(n85), .B(n83), .S(n93), .Z(n81) );
  MUX21L U253 ( .A(n92), .B(n94), .S(n310), .Z(SUM[21]) );
  MUX21L U254 ( .A(n96), .B(n97), .S(n106), .Z(n94) );
  MUX21H U255 ( .A(n105), .B(A[19]), .S(n304), .Z(SUM[19]) );
  ENI U256 ( .A(n304), .B(n107), .Z(SUM[18]) );
  MUX21L U257 ( .A(n33), .B(n28), .S(n310), .Z(SUM[31]) );
  MUX21L U258 ( .A(n30), .B(n31), .S(n4), .Z(n28) );
  MUX21L U259 ( .A(n33), .B(n32), .S(n45), .Z(n30) );
  MUX21L U260 ( .A(n5), .B(n34), .S(n310), .Z(SUM[30]) );
  MUX21L U261 ( .A(n36), .B(n37), .S(n4), .Z(n34) );
  MUX21L U262 ( .A(n6), .B(n39), .S(n310), .Z(SUM[29]) );
  MUX21L U263 ( .A(n297), .B(n47), .S(n4), .Z(n39) );
  MUX21L U264 ( .A(n7), .B(n49), .S(n310), .Z(SUM[28]) );
  MUX21L U265 ( .A(n51), .B(n53), .S(n4), .Z(n49) );
  ENI U266 ( .A(n181), .B(n179), .Z(SUM[6]) );
  MUX21L U267 ( .A(n134), .B(n133), .S(n155), .Z(SUM[14]) );
  MUX21L U268 ( .A(n18), .B(n121), .S(n155), .Z(SUM[16]) );
  MUX21L U269 ( .A(n123), .B(n125), .S(n139), .Z(n121) );
  MUX21L U270 ( .A(n142), .B(n143), .S(n152), .Z(n140) );
  MUX21L U271 ( .A(n23), .B(n298), .S(n155), .Z(SUM[11]) );
  MUX21L U272 ( .A(n110), .B(n117), .S(n157), .Z(SUM[17]) );
  MUX21L U273 ( .A(n119), .B(n113), .S(n141), .Z(n110) );
  MUX21L U274 ( .A(n116), .B(n117), .S(n132), .Z(n113) );
  MUX21H U275 ( .A(n161), .B(n162), .S(n175), .Z(n306) );
  ENI U276 ( .A(n175), .B(n167), .Z(n166) );
  MUX21L U277 ( .A(n308), .B(n25), .S(n191), .Z(SUM[5]) );
  EOI U278 ( .A(n187), .B(n25), .Z(n308) );
  ENI U279 ( .A(n191), .B(n187), .Z(SUM[4]) );
  EOI U280 ( .A(n192), .B(A[3]), .Z(SUM[3]) );
  IVI U281 ( .A(n95), .Z(n93) );
  IVI U282 ( .A(n86), .Z(n84) );
  IVI U283 ( .A(n60), .Z(n58) );
  IVI U284 ( .A(n57), .Z(n8) );
  IVI U285 ( .A(n53), .Z(n7) );
  IVI U286 ( .A(n47), .Z(n6) );
  IVI U287 ( .A(n37), .Z(n5) );
  IVI U288 ( .A(n31), .Z(n33) );
  IVI U289 ( .A(n185), .Z(n25) );
  IVI U290 ( .A(n153), .Z(n24) );
  IVI U291 ( .A(A[11]), .Z(n23) );
  IVI U292 ( .A(n183), .Z(n181) );
  IVI U293 ( .A(n176), .Z(n172) );
  IVI U294 ( .A(n170), .Z(n167) );
  IVI U295 ( .A(n164), .Z(n162) );
  IVI U296 ( .A(A[19]), .Z(n16) );
  IVI U297 ( .A(n157), .Z(n155) );
  IVI U298 ( .A(n148), .Z(n146) );
  IVI U299 ( .A(n97), .Z(n92) );
  IVI U300 ( .A(n141), .Z(n139) );
  IVI U301 ( .A(n143), .Z(n21) );
  IVI U302 ( .A(n136), .Z(n134) );
  IVI U303 ( .A(n132), .Z(n130) );
  IVI U304 ( .A(n125), .Z(n18) );
  IVI U305 ( .A(n83), .Z(n82) );
  IVI U306 ( .A(n119), .Z(n117) );
  IVI U307 ( .A(n79), .Z(n76) );
  IVI U308 ( .A(n73), .Z(n70) );
  IVI U309 ( .A(n192), .Z(SUM[2]) );
endmodule


module pc ( clk, rst, fd_br_signext_sl2, fd_Inst_25_0, fwd_gpr_rd_data1, 
        d_stall, jump, branch, jump_reg, pc, d_pc_plus_8 );
  input [31:0] fd_br_signext_sl2;
  input [25:0] fd_Inst_25_0;
  input [31:0] fwd_gpr_rd_data1;
  output [31:0] pc;
  output [31:0] d_pc_plus_8;
  input clk, rst, d_stall, jump, branch, jump_reg;
  wire   n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n140, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n139, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235;
  wire   [31:0] pc_plus_4;
  wire   [31:0] br_loc;
  assign d_pc_plus_8[31] = pc_plus_4[31];
  assign d_pc_plus_8[30] = pc_plus_4[30];
  assign d_pc_plus_8[29] = pc_plus_4[29];
  assign d_pc_plus_8[28] = pc_plus_4[28];
  assign d_pc_plus_8[27] = pc_plus_4[27];
  assign d_pc_plus_8[26] = pc_plus_4[26];
  assign d_pc_plus_8[25] = pc_plus_4[25];
  assign d_pc_plus_8[24] = pc_plus_4[24];
  assign d_pc_plus_8[23] = pc_plus_4[23];
  assign d_pc_plus_8[22] = pc_plus_4[22];
  assign d_pc_plus_8[21] = pc_plus_4[21];
  assign d_pc_plus_8[20] = pc_plus_4[20];
  assign d_pc_plus_8[19] = pc_plus_4[19];
  assign d_pc_plus_8[18] = pc_plus_4[18];
  assign d_pc_plus_8[17] = pc_plus_4[17];
  assign d_pc_plus_8[16] = pc_plus_4[16];
  assign d_pc_plus_8[15] = pc_plus_4[15];
  assign d_pc_plus_8[14] = pc_plus_4[14];
  assign d_pc_plus_8[13] = pc_plus_4[13];
  assign d_pc_plus_8[12] = pc_plus_4[12];
  assign d_pc_plus_8[11] = pc_plus_4[11];
  assign d_pc_plus_8[10] = pc_plus_4[10];
  assign d_pc_plus_8[9] = pc_plus_4[9];
  assign d_pc_plus_8[8] = pc_plus_4[8];
  assign d_pc_plus_8[7] = pc_plus_4[7];
  assign d_pc_plus_8[6] = pc_plus_4[6];
  assign d_pc_plus_8[5] = pc_plus_4[5];
  assign d_pc_plus_8[4] = pc_plus_4[4];
  assign d_pc_plus_8[3] = pc_plus_4[3];
  assign d_pc_plus_8[2] = pc_plus_4[2];
  assign d_pc_plus_8[1] = pc_plus_4[1];
  assign d_pc_plus_8[0] = pc_plus_4[0];

  FD2 \pc_val_reg[0]  ( .D(n140), .CP(clk), .CD(n139), .Q(pc[0]), .QN(n106) );
  FD2 \pc_val_reg[31]  ( .D(n138), .CP(clk), .CD(n139), .Q(pc[31]) );
  FD2 \pc_val_reg[1]  ( .D(n137), .CP(clk), .CD(n139), .Q(pc[1]), .QN(n107) );
  FD2 \pc_val_reg[2]  ( .D(n136), .CP(clk), .CD(n139), .Q(pc[2]) );
  FD2 \pc_val_reg[3]  ( .D(n135), .CP(clk), .CD(n139), .Q(pc[3]) );
  FD2 \pc_val_reg[4]  ( .D(n134), .CP(clk), .CD(n139), .Q(pc[4]), .QN(n47) );
  FD2 \pc_val_reg[5]  ( .D(n133), .CP(clk), .CD(n139), .Q(pc[5]) );
  FD2 \pc_val_reg[6]  ( .D(n132), .CP(clk), .CD(n139), .Q(pc[6]) );
  FD2 \pc_val_reg[7]  ( .D(n131), .CP(clk), .CD(n139), .Q(pc[7]) );
  FD2 \pc_val_reg[8]  ( .D(n130), .CP(clk), .CD(n139), .Q(pc[8]) );
  FD2 \pc_val_reg[9]  ( .D(n129), .CP(clk), .CD(n139), .Q(pc[9]) );
  FD2 \pc_val_reg[10]  ( .D(n128), .CP(clk), .CD(n139), .Q(pc[10]) );
  FD2 \pc_val_reg[11]  ( .D(n127), .CP(clk), .CD(n139), .Q(pc[11]) );
  FD2 \pc_val_reg[12]  ( .D(n126), .CP(clk), .CD(n139), .Q(pc[12]) );
  FD2 \pc_val_reg[13]  ( .D(n125), .CP(clk), .CD(n139), .Q(pc[13]) );
  FD2 \pc_val_reg[14]  ( .D(n124), .CP(clk), .CD(n139), .QN(n97) );
  FD2 \pc_val_reg[15]  ( .D(n123), .CP(clk), .CD(n139), .Q(pc[15]) );
  FD2 \pc_val_reg[16]  ( .D(n122), .CP(clk), .CD(n139), .Q(pc[16]) );
  FD2 \pc_val_reg[17]  ( .D(n121), .CP(clk), .CD(n139), .QN(n87) );
  FD2 \pc_val_reg[18]  ( .D(n120), .CP(clk), .CD(n139), .Q(pc[18]) );
  FD2 \pc_val_reg[19]  ( .D(n119), .CP(clk), .CD(n139), .Q(pc[19]) );
  FD2 \pc_val_reg[20]  ( .D(n118), .CP(clk), .CD(n139), .Q(pc[20]) );
  FD2 \pc_val_reg[21]  ( .D(n117), .CP(clk), .CD(n139), .QN(n89) );
  FD2 \pc_val_reg[22]  ( .D(n116), .CP(clk), .CD(n139), .Q(pc[22]) );
  FD2 \pc_val_reg[23]  ( .D(n115), .CP(clk), .CD(n139), .Q(pc[23]) );
  FD2 \pc_val_reg[24]  ( .D(n114), .CP(clk), .CD(n139), .Q(pc[24]) );
  FD2 \pc_val_reg[25]  ( .D(n113), .CP(clk), .CD(n139), .Q(pc[25]) );
  FD2 \pc_val_reg[26]  ( .D(n112), .CP(clk), .CD(n139), .Q(pc[26]) );
  FD2 \pc_val_reg[27]  ( .D(n111), .CP(clk), .CD(n139), .Q(pc[27]) );
  FD2 \pc_val_reg[28]  ( .D(n110), .CP(clk), .CD(n139), .Q(pc[28]) );
  FD2 \pc_val_reg[29]  ( .D(n109), .CP(clk), .CD(n139), .Q(pc[29]) );
  FD2 \pc_val_reg[30]  ( .D(n108), .CP(clk), .CD(n139), .Q(pc[30]) );
  pc_DW01_add_2 add_26 ( .A(pc), .B(fd_br_signext_sl2), .CI(1'b0), .SUM(br_loc) );
  pc_DW01_add_3 r295 ( .A(pc), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(pc_plus_4) );
  NR2I U3 ( .A(n4), .B(n5), .Z(n3) );
  ND2I U6 ( .A(n10), .B(n11), .Z(n4) );
  AN2I U7 ( .A(br_loc[9]), .B(n9), .Z(n5) );
  NR2I U8 ( .A(n7), .B(n8), .Z(n6) );
  ND2I U9 ( .A(n38), .B(n39), .Z(n7) );
  AN2I U10 ( .A(br_loc[8]), .B(n27), .Z(n8) );
  AN2I U11 ( .A(n92), .B(n143), .Z(n9) );
  ND2I U12 ( .A(fwd_gpr_rd_data1[9]), .B(n96), .Z(n10) );
  ND2I U13 ( .A(pc[9]), .B(d_stall), .Z(n11) );
  AN2I U14 ( .A(n12), .B(n13), .Z(n202) );
  ND2I U15 ( .A(fwd_gpr_rd_data1[11]), .B(n96), .Z(n12) );
  ND2I U16 ( .A(pc[11]), .B(d_stall), .Z(n13) );
  AN2I U17 ( .A(n14), .B(n15), .Z(n162) );
  ND2I U18 ( .A(fwd_gpr_rd_data1[24]), .B(n102), .Z(n14) );
  ND2I U19 ( .A(pc[24]), .B(d_stall), .Z(n15) );
  IVI U20 ( .A(n91), .Z(n16) );
  IVI U21 ( .A(n142), .Z(n17) );
  IVI U22 ( .A(n142), .Z(n232) );
  IVI U23 ( .A(d_stall), .Z(n46) );
  AN2I U24 ( .A(n205), .B(n206), .Z(n18) );
  AN2I U25 ( .A(n218), .B(n217), .Z(n19) );
  AN2I U26 ( .A(n210), .B(n211), .Z(n20) );
  AN2I U27 ( .A(fwd_gpr_rd_data1[2]), .B(n96), .Z(n21) );
  AN2I U28 ( .A(pc[2]), .B(d_stall), .Z(n22) );
  NR2I U29 ( .A(n21), .B(n22), .Z(n225) );
  AN2I U30 ( .A(fwd_gpr_rd_data1[3]), .B(n102), .Z(n23) );
  AN2I U31 ( .A(pc[3]), .B(d_stall), .Z(n24) );
  NR2I U32 ( .A(n23), .B(n24), .Z(n222) );
  ND2I U33 ( .A(n216), .B(n19), .Z(n133) );
  AO2 U34 ( .A(fwd_gpr_rd_data1[5]), .B(n100), .C(pc[5]), .D(d_stall), .Z(n216) );
  AN2I U35 ( .A(n25), .B(n26), .Z(n221) );
  ND2I U36 ( .A(fd_Inst_25_0[2]), .B(n104), .Z(n25) );
  ND2I U37 ( .A(pc_plus_4[4]), .B(n198), .Z(n26) );
  AN2I U38 ( .A(n92), .B(n143), .Z(n27) );
  IVI U39 ( .A(n152), .Z(n28) );
  B4I U40 ( .A(n152), .Z(n198) );
  ND2I U41 ( .A(n162), .B(n163), .Z(n29) );
  ND2I U42 ( .A(n164), .B(n30), .Z(n114) );
  IVI U43 ( .A(n29), .Z(n30) );
  IVI U44 ( .A(n142), .Z(n31) );
  AN2I U45 ( .A(fd_Inst_25_0[21]), .B(n105), .Z(n32) );
  AN2I U46 ( .A(pc_plus_4[23]), .B(n198), .Z(n33) );
  NR2I U47 ( .A(n32), .B(n33), .Z(n167) );
  AO2P U48 ( .A(fd_Inst_25_0[3]), .B(n104), .C(pc_plus_4[5]), .D(n31), .Z(n218) );
  AO2P U49 ( .A(fd_Inst_25_0[1]), .B(n104), .C(pc_plus_4[3]), .D(n31), .Z(n224) );
  ND2I U50 ( .A(n212), .B(n20), .Z(n131) );
  ND2I U51 ( .A(fd_Inst_25_0[5]), .B(n104), .Z(n34) );
  ND2I U52 ( .A(pc_plus_4[7]), .B(n66), .Z(n35) );
  AN2I U53 ( .A(n34), .B(n35), .Z(n212) );
  ND2I U54 ( .A(n208), .B(n3), .Z(n129) );
  ND2I U55 ( .A(fd_Inst_25_0[7]), .B(n104), .Z(n36) );
  ND2I U56 ( .A(pc_plus_4[9]), .B(n66), .Z(n37) );
  AN2I U57 ( .A(n36), .B(n37), .Z(n208) );
  AO2P U58 ( .A(fwd_gpr_rd_data1[6]), .B(n71), .C(pc[6]), .D(d_stall), .Z(n213) );
  ND2I U59 ( .A(fwd_gpr_rd_data1[8]), .B(n101), .Z(n38) );
  ND2I U60 ( .A(pc[8]), .B(d_stall), .Z(n39) );
  ND2I U61 ( .A(fwd_gpr_rd_data1[12]), .B(n71), .Z(n40) );
  ND2I U62 ( .A(pc[12]), .B(d_stall), .Z(n41) );
  AN2I U63 ( .A(n40), .B(n41), .Z(n199) );
  ND2I U64 ( .A(n202), .B(n203), .Z(n42) );
  ND2I U65 ( .A(n204), .B(n43), .Z(n127) );
  IVI U66 ( .A(n42), .Z(n43) );
  ND2I U67 ( .A(n221), .B(n220), .Z(n44) );
  ND2I U68 ( .A(n219), .B(n45), .Z(n134) );
  IVI U69 ( .A(n44), .Z(n45) );
  EO1 U70 ( .A(fwd_gpr_rd_data1[4]), .B(n16), .C(n47), .D(n46), .Z(n219) );
  IVI U71 ( .A(n152), .Z(n48) );
  AN2I U72 ( .A(fd_Inst_25_0[24]), .B(n104), .Z(n49) );
  AN2I U73 ( .A(pc_plus_4[26]), .B(n198), .Z(n50) );
  NR2I U74 ( .A(n49), .B(n50), .Z(n158) );
  AN2I U75 ( .A(fd_Inst_25_0[11]), .B(n105), .Z(n51) );
  AN2I U76 ( .A(pc_plus_4[13]), .B(n232), .Z(n52) );
  NR2I U77 ( .A(n51), .B(n52), .Z(n197) );
  B4I U78 ( .A(n150), .Z(n105) );
  AO2P U79 ( .A(fd_Inst_25_0[0]), .B(n104), .C(pc_plus_4[2]), .D(n28), .Z(n227) );
  IVI U80 ( .A(n88), .Z(n53) );
  ND2I U81 ( .A(n213), .B(n214), .Z(n54) );
  ND2I U82 ( .A(n215), .B(n55), .Z(n132) );
  IVI U83 ( .A(n54), .Z(n55) );
  ND2I U84 ( .A(n209), .B(n6), .Z(n130) );
  ND2I U85 ( .A(n207), .B(n18), .Z(n128) );
  ND2I U86 ( .A(fd_Inst_25_0[8]), .B(n104), .Z(n56) );
  ND2I U87 ( .A(pc_plus_4[10]), .B(n48), .Z(n57) );
  AN2I U88 ( .A(n56), .B(n57), .Z(n207) );
  B4I U89 ( .A(n150), .Z(n104) );
  ND2I U90 ( .A(n199), .B(n200), .Z(n58) );
  ND2I U91 ( .A(n201), .B(n59), .Z(n126) );
  IVI U92 ( .A(n58), .Z(n59) );
  ND2I U93 ( .A(fd_Inst_25_0[10]), .B(n105), .Z(n60) );
  ND2I U94 ( .A(pc_plus_4[12]), .B(n48), .Z(n61) );
  AN2I U95 ( .A(n60), .B(n61), .Z(n201) );
  ND2I U96 ( .A(n186), .B(n187), .Z(n62) );
  ND2I U97 ( .A(n188), .B(n63), .Z(n122) );
  IVI U98 ( .A(n62), .Z(n63) );
  ND2I U99 ( .A(n180), .B(n181), .Z(n64) );
  ND2I U100 ( .A(n182), .B(n65), .Z(n120) );
  IVI U101 ( .A(n64), .Z(n65) );
  IVI U102 ( .A(n142), .Z(n66) );
  AN2I U103 ( .A(fd_Inst_25_0[22]), .B(n105), .Z(n67) );
  AN2I U104 ( .A(pc_plus_4[24]), .B(n17), .Z(n68) );
  NR2I U105 ( .A(n67), .B(n68), .Z(n164) );
  IVI U106 ( .A(n89), .Z(pc[21]) );
  IVI U107 ( .A(n87), .Z(pc[17]) );
  IVI U108 ( .A(n97), .Z(pc[14]) );
  AN2I U109 ( .A(n143), .B(n103), .Z(n69) );
  OR2I U110 ( .A(n103), .B(n233), .Z(n70) );
  AO3 U111 ( .A(n106), .B(n46), .C(n231), .D(n230), .Z(n140) );
  AO3 U112 ( .A(n107), .B(n46), .C(n229), .D(n228), .Z(n137) );
  IVI U113 ( .A(n88), .Z(n71) );
  AN2I U114 ( .A(n194), .B(n193), .Z(n72) );
  AN2I U115 ( .A(n185), .B(n184), .Z(n73) );
  AN2I U116 ( .A(n176), .B(n175), .Z(n74) );
  AN2I U117 ( .A(n170), .B(n169), .Z(n75) );
  AN2I U118 ( .A(n161), .B(n160), .Z(n76) );
  AN2I U119 ( .A(n155), .B(n154), .Z(n77) );
  AN2I U120 ( .A(n191), .B(n190), .Z(n78) );
  AN2I U121 ( .A(n177), .B(n178), .Z(n79) );
  AN2I U122 ( .A(n173), .B(n172), .Z(n80) );
  AN2I U123 ( .A(n167), .B(n166), .Z(n81) );
  AN2I U124 ( .A(n158), .B(n157), .Z(n82) );
  AO2 U125 ( .A(fwd_gpr_rd_data1[14]), .B(n16), .C(pc[14]), .D(d_stall), .Z(
        n192) );
  AO2 U126 ( .A(fwd_gpr_rd_data1[17]), .B(n99), .C(pc[17]), .D(d_stall), .Z(
        n183) );
  AO2 U127 ( .A(fwd_gpr_rd_data1[21]), .B(n99), .C(pc[21]), .D(d_stall), .Z(
        n171) );
  AN2I U128 ( .A(n92), .B(n143), .Z(n86) );
  ND2I U129 ( .A(n183), .B(n73), .Z(n121) );
  AO2P U130 ( .A(fwd_gpr_rd_data1[18]), .B(n99), .C(pc[18]), .D(d_stall), .Z(
        n180) );
  AO2P U131 ( .A(fwd_gpr_rd_data1[13]), .B(n99), .C(pc[13]), .D(d_stall), .Z(
        n195) );
  AO2P U132 ( .A(fwd_gpr_rd_data1[16]), .B(n101), .C(pc[16]), .D(d_stall), .Z(
        n186) );
  ND2I U133 ( .A(n179), .B(n79), .Z(n119) );
  IVI U134 ( .A(n90), .Z(n88) );
  ND2I U135 ( .A(n171), .B(n80), .Z(n117) );
  ND2I U136 ( .A(n165), .B(n81), .Z(n115) );
  ND2I U137 ( .A(n159), .B(n76), .Z(n113) );
  NR2I U138 ( .A(branch), .B(n70), .Z(n90) );
  ND2P U139 ( .A(n141), .B(n46), .Z(n233) );
  ND2I U140 ( .A(n156), .B(n82), .Z(n112) );
  IVI U141 ( .A(n90), .Z(n91) );
  AO2P U142 ( .A(pc_plus_4[0]), .B(n28), .C(br_loc[0]), .D(n86), .Z(n230) );
  AO2P U143 ( .A(pc_plus_4[1]), .B(n28), .C(br_loc[1]), .D(n86), .Z(n228) );
  IVI U144 ( .A(n151), .Z(n92) );
  IVI U145 ( .A(n86), .Z(n93) );
  IVI U146 ( .A(n93), .Z(n94) );
  IVI U147 ( .A(n93), .Z(n95) );
  IVI U148 ( .A(n88), .Z(n96) );
  ND2I U149 ( .A(n192), .B(n72), .Z(n124) );
  ND2I U150 ( .A(n189), .B(n78), .Z(n123) );
  ND2I U151 ( .A(n174), .B(n74), .Z(n118) );
  ND2I U152 ( .A(n168), .B(n75), .Z(n116) );
  ND2I U153 ( .A(n153), .B(n77), .Z(n111) );
  AN2I U154 ( .A(n92), .B(n143), .Z(n98) );
  IVI U155 ( .A(jump_reg), .Z(n103) );
  IVI U156 ( .A(n88), .Z(n99) );
  IVI U157 ( .A(n91), .Z(n100) );
  IVI U158 ( .A(n91), .Z(n101) );
  IVI U159 ( .A(n91), .Z(n102) );
  IVI U160 ( .A(rst), .Z(n139) );
  IVI U161 ( .A(jump), .Z(n141) );
  IVI U162 ( .A(n233), .Z(n143) );
  IVI U163 ( .A(branch), .Z(n151) );
  ND2I U164 ( .A(n69), .B(n151), .Z(n142) );
  AO2 U165 ( .A(pc_plus_4[30]), .B(n66), .C(br_loc[30]), .D(n27), .Z(n145) );
  AO2 U166 ( .A(fwd_gpr_rd_data1[30]), .B(n53), .C(pc[30]), .D(n233), .Z(n144)
         );
  ND2I U167 ( .A(n145), .B(n144), .Z(n108) );
  AO2 U168 ( .A(pc_plus_4[29]), .B(n66), .C(br_loc[29]), .D(n27), .Z(n147) );
  AO2 U169 ( .A(fwd_gpr_rd_data1[29]), .B(n100), .C(pc[29]), .D(n233), .Z(n146) );
  ND2I U170 ( .A(n147), .B(n146), .Z(n109) );
  AO2 U171 ( .A(pc_plus_4[28]), .B(n31), .C(br_loc[28]), .D(n9), .Z(n149) );
  AO2 U172 ( .A(fwd_gpr_rd_data1[28]), .B(n99), .C(pc[28]), .D(n233), .Z(n148)
         );
  ND2I U173 ( .A(n149), .B(n148), .Z(n110) );
  ND2I U174 ( .A(jump), .B(n46), .Z(n150) );
  ND2I U175 ( .A(n69), .B(n151), .Z(n152) );
  AO2 U176 ( .A(fd_Inst_25_0[25]), .B(n105), .C(pc_plus_4[27]), .D(n232), .Z(
        n155) );
  ND2I U177 ( .A(br_loc[27]), .B(n27), .Z(n154) );
  AO2 U178 ( .A(fwd_gpr_rd_data1[27]), .B(n53), .C(pc[27]), .D(d_stall), .Z(
        n153) );
  ND2I U179 ( .A(br_loc[26]), .B(n98), .Z(n157) );
  AO2 U180 ( .A(fwd_gpr_rd_data1[26]), .B(n53), .C(pc[26]), .D(d_stall), .Z(
        n156) );
  AO2 U181 ( .A(fd_Inst_25_0[23]), .B(n105), .C(pc_plus_4[25]), .D(n232), .Z(
        n161) );
  ND2I U182 ( .A(br_loc[25]), .B(n9), .Z(n160) );
  AO2 U183 ( .A(fwd_gpr_rd_data1[25]), .B(n100), .C(pc[25]), .D(d_stall), .Z(
        n159) );
  ND2I U184 ( .A(br_loc[24]), .B(n95), .Z(n163) );
  ND2I U185 ( .A(br_loc[23]), .B(n9), .Z(n166) );
  AO2 U186 ( .A(fwd_gpr_rd_data1[23]), .B(n100), .C(pc[23]), .D(d_stall), .Z(
        n165) );
  AO2 U187 ( .A(fd_Inst_25_0[20]), .B(n104), .C(pc_plus_4[22]), .D(n17), .Z(
        n170) );
  ND2I U188 ( .A(br_loc[22]), .B(n9), .Z(n169) );
  AO2 U189 ( .A(fwd_gpr_rd_data1[22]), .B(n53), .C(pc[22]), .D(d_stall), .Z(
        n168) );
  AO2 U190 ( .A(fd_Inst_25_0[19]), .B(n105), .C(pc_plus_4[21]), .D(n198), .Z(
        n173) );
  ND2I U191 ( .A(br_loc[21]), .B(n27), .Z(n172) );
  AO2 U192 ( .A(fd_Inst_25_0[18]), .B(n104), .C(pc_plus_4[20]), .D(n17), .Z(
        n176) );
  ND2I U193 ( .A(br_loc[20]), .B(n98), .Z(n175) );
  AO2 U194 ( .A(fwd_gpr_rd_data1[20]), .B(n71), .C(pc[20]), .D(d_stall), .Z(
        n174) );
  AO2 U195 ( .A(fd_Inst_25_0[17]), .B(n105), .C(pc_plus_4[19]), .D(n31), .Z(
        n179) );
  ND2I U196 ( .A(br_loc[19]), .B(n98), .Z(n178) );
  AO2 U197 ( .A(fwd_gpr_rd_data1[19]), .B(n16), .C(pc[19]), .D(d_stall), .Z(
        n177) );
  AO2 U198 ( .A(fd_Inst_25_0[16]), .B(n105), .C(pc_plus_4[18]), .D(n66), .Z(
        n182) );
  ND2I U199 ( .A(br_loc[18]), .B(n94), .Z(n181) );
  AO2 U200 ( .A(fd_Inst_25_0[15]), .B(n105), .C(pc_plus_4[17]), .D(n198), .Z(
        n185) );
  ND2I U201 ( .A(br_loc[17]), .B(n9), .Z(n184) );
  AO2 U202 ( .A(fd_Inst_25_0[14]), .B(n105), .C(pc_plus_4[16]), .D(n48), .Z(
        n188) );
  ND2I U203 ( .A(br_loc[16]), .B(n95), .Z(n187) );
  AO2 U204 ( .A(fd_Inst_25_0[13]), .B(n105), .C(pc_plus_4[15]), .D(n198), .Z(
        n191) );
  ND2I U205 ( .A(br_loc[15]), .B(n98), .Z(n190) );
  AO2 U206 ( .A(fwd_gpr_rd_data1[15]), .B(n53), .C(pc[15]), .D(d_stall), .Z(
        n189) );
  AO2 U207 ( .A(fd_Inst_25_0[12]), .B(n105), .C(pc_plus_4[14]), .D(n198), .Z(
        n194) );
  ND2I U208 ( .A(br_loc[14]), .B(n27), .Z(n193) );
  ND2I U209 ( .A(br_loc[13]), .B(n27), .Z(n196) );
  ND3 U210 ( .A(n197), .B(n196), .C(n195), .Z(n125) );
  ND2I U211 ( .A(br_loc[12]), .B(n95), .Z(n200) );
  AO2 U212 ( .A(fd_Inst_25_0[9]), .B(n105), .C(pc_plus_4[11]), .D(n48), .Z(
        n204) );
  ND2I U213 ( .A(br_loc[11]), .B(n94), .Z(n203) );
  ND2I U214 ( .A(br_loc[10]), .B(n98), .Z(n206) );
  AO2 U215 ( .A(fwd_gpr_rd_data1[10]), .B(n102), .C(pc[10]), .D(d_stall), .Z(
        n205) );
  AO2 U216 ( .A(fd_Inst_25_0[6]), .B(n104), .C(pc_plus_4[8]), .D(n48), .Z(n209) );
  ND2I U217 ( .A(br_loc[7]), .B(n9), .Z(n211) );
  AO2 U218 ( .A(fwd_gpr_rd_data1[7]), .B(n101), .C(pc[7]), .D(d_stall), .Z(
        n210) );
  AO2 U219 ( .A(fd_Inst_25_0[4]), .B(n104), .C(pc_plus_4[6]), .D(n48), .Z(n215) );
  ND2I U220 ( .A(br_loc[6]), .B(n98), .Z(n214) );
  ND2I U221 ( .A(br_loc[5]), .B(n27), .Z(n217) );
  ND2I U222 ( .A(br_loc[4]), .B(n94), .Z(n220) );
  ND2I U223 ( .A(br_loc[3]), .B(n9), .Z(n223) );
  ND3 U224 ( .A(n224), .B(n223), .C(n222), .Z(n135) );
  ND2I U225 ( .A(br_loc[2]), .B(n98), .Z(n226) );
  ND3 U226 ( .A(n227), .B(n226), .C(n225), .Z(n136) );
  ND2I U227 ( .A(fwd_gpr_rd_data1[1]), .B(n71), .Z(n229) );
  ND2I U228 ( .A(fwd_gpr_rd_data1[0]), .B(n53), .Z(n231) );
  AO2 U229 ( .A(pc_plus_4[31]), .B(n66), .C(br_loc[31]), .D(n98), .Z(n235) );
  AO2 U230 ( .A(fwd_gpr_rd_data1[31]), .B(n100), .C(pc[31]), .D(n233), .Z(n234) );
  ND2I U231 ( .A(n235), .B(n234), .Z(n138) );
endmodule


module control_unit_DW01_cmp6_3 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n34,
         n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n51,
         n54, n55, n56, n58, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n87,
         n90, n94, n95, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192;

  ND2I U5 ( .A(n8), .B(n5), .Z(n4) );
  NR2I U6 ( .A(n7), .B(n6), .Z(n5) );
  ENI U7 ( .A(A[31]), .B(n64), .Z(n6) );
  ENI U8 ( .A(A[30]), .B(n65), .Z(n7) );
  NR2I U9 ( .A(n10), .B(n9), .Z(n8) );
  ENI U10 ( .A(A[29]), .B(n66), .Z(n9) );
  ENI U11 ( .A(A[28]), .B(n67), .Z(n10) );
  ND2I U12 ( .A(n15), .B(n12), .Z(n11) );
  NR2I U13 ( .A(n14), .B(n13), .Z(n12) );
  ENI U14 ( .A(n68), .B(A[27]), .Z(n13) );
  ENI U15 ( .A(A[26]), .B(n69), .Z(n14) );
  NR2I U16 ( .A(n17), .B(n16), .Z(n15) );
  ENI U17 ( .A(n70), .B(A[25]), .Z(n16) );
  ENI U18 ( .A(n71), .B(A[24]), .Z(n17) );
  NR2I U21 ( .A(n22), .B(n21), .Z(n20) );
  ENI U22 ( .A(n72), .B(A[23]), .Z(n21) );
  ENI U23 ( .A(A[22]), .B(n73), .Z(n22) );
  NR2I U24 ( .A(n25), .B(n24), .Z(n23) );
  ENI U25 ( .A(n74), .B(A[21]), .Z(n24) );
  ENI U26 ( .A(A[20]), .B(n75), .Z(n25) );
  NR2I U28 ( .A(n29), .B(n28), .Z(n27) );
  ENI U29 ( .A(n76), .B(A[19]), .Z(n28) );
  ENI U30 ( .A(A[18]), .B(n77), .Z(n29) );
  NR2I U31 ( .A(n32), .B(n31), .Z(n30) );
  ENI U32 ( .A(A[17]), .B(n78), .Z(n31) );
  ENI U33 ( .A(n79), .B(A[16]), .Z(n32) );
  NR2I U37 ( .A(n38), .B(n37), .Z(n36) );
  ENI U38 ( .A(n80), .B(A[15]), .Z(n37) );
  NR2I U40 ( .A(n41), .B(n40), .Z(n39) );
  ENI U41 ( .A(n82), .B(A[13]), .Z(n40) );
  ENI U42 ( .A(A[12]), .B(n83), .Z(n41) );
  NR2I U44 ( .A(n45), .B(n44), .Z(n43) );
  ENI U45 ( .A(n84), .B(A[11]), .Z(n44) );
  NR2I U47 ( .A(n48), .B(n47), .Z(n46) );
  ENI U49 ( .A(n87), .B(A[8]), .Z(n48) );
  NR2I U55 ( .A(n56), .B(n55), .Z(n54) );
  ENI U56 ( .A(n90), .B(A[5]), .Z(n55) );
  ENI U63 ( .A(A[1]), .B(n94), .Z(n62) );
  ENI U64 ( .A(A[0]), .B(n95), .Z(n63) );
  ENI U100 ( .A(A[3]), .B(B[3]), .Z(n167) );
  IVI U101 ( .A(B[9]), .Z(n168) );
  ENI U102 ( .A(A[9]), .B(n168), .Z(n47) );
  ENI U103 ( .A(B[7]), .B(A[7]), .Z(n169) );
  AN2I U104 ( .A(n170), .B(n171), .Z(n3) );
  IVI U105 ( .A(n4), .Z(n170) );
  IVI U106 ( .A(n11), .Z(n171) );
  AN2I U107 ( .A(n172), .B(n173), .Z(n34) );
  IVI U108 ( .A(n192), .Z(n172) );
  IVI U109 ( .A(n191), .Z(n173) );
  AN2I U110 ( .A(n174), .B(n175), .Z(n61) );
  IVI U111 ( .A(n63), .Z(n174) );
  IVI U112 ( .A(n62), .Z(n175) );
  IVI U113 ( .A(n177), .Z(n45) );
  IVI U114 ( .A(n178), .Z(n176) );
  ENI U115 ( .A(A[10]), .B(B[10]), .Z(n177) );
  ND2I U116 ( .A(n176), .B(n179), .Z(n180) );
  ND2I U117 ( .A(n178), .B(B[4]), .Z(n181) );
  ND2I U118 ( .A(n180), .B(n181), .Z(n56) );
  IVI U119 ( .A(A[4]), .Z(n178) );
  IVI U120 ( .A(B[4]), .Z(n179) );
  ND2I U121 ( .A(n185), .B(n186), .Z(NE) );
  AN2I U122 ( .A(n183), .B(n169), .Z(n51) );
  ENI U123 ( .A(A[6]), .B(B[6]), .Z(n183) );
  AN2I U124 ( .A(n184), .B(n167), .Z(n58) );
  ENI U125 ( .A(A[2]), .B(B[2]), .Z(n184) );
  AN2I U126 ( .A(n185), .B(n186), .Z(EQ) );
  AN2I U127 ( .A(n49), .B(n34), .Z(n185) );
  AN2I U128 ( .A(n18), .B(n3), .Z(n186) );
  NR2I U129 ( .A(n187), .B(n188), .Z(n18) );
  ND2I U130 ( .A(n30), .B(n27), .Z(n187) );
  ND2I U131 ( .A(n23), .B(n20), .Z(n188) );
  NR2I U132 ( .A(n189), .B(n190), .Z(n49) );
  ND2I U133 ( .A(n61), .B(n58), .Z(n189) );
  ND2I U134 ( .A(n54), .B(n51), .Z(n190) );
  ND2I U135 ( .A(n46), .B(n43), .Z(n191) );
  ND2I U136 ( .A(n39), .B(n36), .Z(n192) );
  EOI U137 ( .A(A[14]), .B(B[14]), .Z(n38) );
  IVI U138 ( .A(B[0]), .Z(n95) );
  IVI U139 ( .A(B[1]), .Z(n94) );
  IVI U140 ( .A(B[5]), .Z(n90) );
  IVI U141 ( .A(B[8]), .Z(n87) );
  IVI U142 ( .A(B[11]), .Z(n84) );
  IVI U143 ( .A(B[12]), .Z(n83) );
  IVI U144 ( .A(B[13]), .Z(n82) );
  IVI U145 ( .A(B[15]), .Z(n80) );
  IVI U146 ( .A(B[16]), .Z(n79) );
  IVI U147 ( .A(B[17]), .Z(n78) );
  IVI U148 ( .A(B[18]), .Z(n77) );
  IVI U149 ( .A(B[19]), .Z(n76) );
  IVI U150 ( .A(B[20]), .Z(n75) );
  IVI U151 ( .A(B[21]), .Z(n74) );
  IVI U152 ( .A(B[22]), .Z(n73) );
  IVI U153 ( .A(B[23]), .Z(n72) );
  IVI U154 ( .A(B[24]), .Z(n71) );
  IVI U155 ( .A(B[25]), .Z(n70) );
  IVI U156 ( .A(B[26]), .Z(n69) );
  IVI U157 ( .A(B[27]), .Z(n68) );
  IVI U158 ( .A(B[28]), .Z(n67) );
  IVI U159 ( .A(B[29]), .Z(n66) );
  IVI U160 ( .A(B[30]), .Z(n65) );
  IVI U161 ( .A(B[31]), .Z(n64) );
endmodule


module control_unit ( mw_opcode, mw_funct, mw_rs, mw_rt, mw_rd, xm_opcode, 
        dx_opcode, dx_funct, fd_opcode, fd_funct, fwd_gpr_rd_data1, 
        fwd_gpr_rd_data2, w_RegWrite, w_RegDest, w_MemtoReg, w_isJAL, 
        m_MemRead, m_MemWrite, m_isJAL, m_RegDest, x_ALUSrc, x_isSLL_SRL, 
        x_ALU_Control, d_PCSrc1, d_PCSrc2, d_PCSrc3, d_isSLL_SRL );
  input [5:0] mw_opcode;
  input [5:0] mw_funct;
  input [4:0] mw_rs;
  input [4:0] mw_rt;
  input [4:0] mw_rd;
  input [5:0] xm_opcode;
  input [5:0] dx_opcode;
  input [5:0] dx_funct;
  input [5:0] fd_opcode;
  input [5:0] fd_funct;
  input [31:0] fwd_gpr_rd_data1;
  input [31:0] fwd_gpr_rd_data2;
  output [2:0] x_ALU_Control;
  output w_RegWrite, w_RegDest, w_MemtoReg, w_isJAL, m_MemRead, m_MemWrite,
         m_isJAL, m_RegDest, x_ALUSrc, x_isSLL_SRL, d_PCSrc1, d_PCSrc2,
         d_PCSrc3, d_isSLL_SRL;
  wire   N67, N68, n65, n1, n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123;

  NR2I U44 ( .A(n10), .B(n31), .Z(n65) );
  control_unit_DW01_cmp6_3 r294 ( .A(fwd_gpr_rd_data1), .B(fwd_gpr_rd_data2), 
        .TC(1'b0), .EQ(N67), .NE(N68) );
  AN2I U3 ( .A(n105), .B(n104), .Z(n1) );
  AN2I U4 ( .A(n96), .B(n95), .Z(n2) );
  AN2I U5 ( .A(n97), .B(n2), .Z(n3) );
  ND6P U6 ( .A(n20), .B(n21), .C(n22), .D(n23), .E(n95), .F(n96), .Z(n24) );
  IVDA U7 ( .A(n22), .Y(n4), .Z(n6) );
  AN2I U8 ( .A(n73), .B(n90), .Z(n7) );
  AN3 U9 ( .A(n105), .B(n108), .C(n103), .Z(n8) );
  IVI U10 ( .A(n23), .Z(n9) );
  IVI U11 ( .A(n20), .Z(n10) );
  IVI U12 ( .A(n15), .Z(n11) );
  IVI U13 ( .A(n14), .Z(n12) );
  AO3P U14 ( .A(dx_opcode[0]), .B(n93), .C(n92), .D(n91), .Z(x_ALU_Control[2])
         );
  ND4P U15 ( .A(n53), .B(n61), .C(n56), .D(n47), .Z(n51) );
  AN2I U16 ( .A(n13), .B(n1), .Z(w_isJAL) );
  IVI U17 ( .A(n106), .Z(n13) );
  ND6 U18 ( .A(n14), .B(n15), .C(n25), .D(n16), .E(n17), .F(n18), .Z(n19) );
  IVI U19 ( .A(mw_opcode[4]), .Z(n14) );
  IVI U20 ( .A(mw_opcode[2]), .Z(n15) );
  IVI U21 ( .A(mw_opcode[3]), .Z(n16) );
  IVI U22 ( .A(mw_opcode[5]), .Z(n17) );
  IVI U23 ( .A(mw_opcode[0]), .Z(n18) );
  IVI U24 ( .A(n19), .Z(w_RegDest) );
  IVI U25 ( .A(xm_opcode[2]), .Z(n20) );
  IVI U26 ( .A(xm_opcode[5]), .Z(n21) );
  IVI U27 ( .A(xm_opcode[1]), .Z(n22) );
  IVI U28 ( .A(xm_opcode[0]), .Z(n23) );
  IVI U29 ( .A(n24), .Z(m_RegDest) );
  IVI U30 ( .A(mw_opcode[1]), .Z(n25) );
  IVI U31 ( .A(n25), .Z(n26) );
  AN2I U32 ( .A(n52), .B(n55), .Z(n47) );
  IVI U33 ( .A(n108), .Z(n27) );
  IVI U34 ( .A(n104), .Z(n28) );
  IVI U35 ( .A(n103), .Z(n29) );
  IVI U36 ( .A(n109), .Z(n30) );
  IVI U37 ( .A(n95), .Z(n31) );
  IVI U38 ( .A(fd_opcode[0]), .Z(n32) );
  AN2I U39 ( .A(n40), .B(n33), .Z(m_isJAL) );
  NR2I U40 ( .A(n99), .B(n6), .Z(n33) );
  IVI U41 ( .A(n21), .Z(n34) );
  IVI U42 ( .A(n96), .Z(n35) );
  ND2I U43 ( .A(n97), .B(n2), .Z(n99) );
  NR2I U45 ( .A(fd_opcode[2]), .B(fd_opcode[4]), .Z(n36) );
  NR3P U46 ( .A(n51), .B(n50), .C(n37), .Z(d_isSLL_SRL) );
  IVI U47 ( .A(n36), .Z(n37) );
  NR6 U48 ( .A(n12), .B(n28), .C(n39), .D(n29), .E(n27), .F(n30), .Z(n38) );
  IVI U49 ( .A(n112), .Z(n39) );
  AO3P U50 ( .A(N67), .B(fd_opcode[0]), .C(n62), .D(n61), .Z(n63) );
  NR2I U51 ( .A(n98), .B(n34), .Z(n40) );
  AN3P U52 ( .A(n42), .B(n72), .C(n82), .Z(n41) );
  IVI U53 ( .A(n78), .Z(n43) );
  NR2I U54 ( .A(n80), .B(n43), .Z(n42) );
  AN3 U55 ( .A(n27), .B(n105), .C(n104), .Z(n44) );
  AN2I U56 ( .A(n46), .B(dx_opcode[2]), .Z(n45) );
  AN3 U57 ( .A(dx_opcode[3]), .B(n71), .C(n78), .Z(n46) );
  ND4P U58 ( .A(n49), .B(n58), .C(n48), .D(n32), .Z(n50) );
  IVI U59 ( .A(fd_opcode[1]), .Z(n61) );
  IVI U60 ( .A(fd_funct[4]), .Z(n53) );
  IVI U61 ( .A(fd_opcode[3]), .Z(n56) );
  IVI U62 ( .A(fd_funct[0]), .Z(n49) );
  IVI U63 ( .A(fd_funct[3]), .Z(n58) );
  IVI U64 ( .A(fd_funct[2]), .Z(n48) );
  NR2I U65 ( .A(fd_funct[2]), .B(fd_funct[0]), .Z(n54) );
  IVI U66 ( .A(fd_funct[5]), .Z(n52) );
  ND4 U67 ( .A(n54), .B(n53), .C(n32), .D(n52), .Z(n60) );
  IVI U68 ( .A(fd_opcode[4]), .Z(n57) );
  IVI U69 ( .A(fd_opcode[5]), .Z(n55) );
  ND3 U70 ( .A(n57), .B(n56), .C(n55), .Z(n66) );
  OR3 U71 ( .A(fd_funct[1]), .B(n58), .C(n66), .Z(n59) );
  NR4 U72 ( .A(n60), .B(n59), .C(fd_opcode[1]), .D(fd_opcode[2]), .Z(d_PCSrc3)
         );
  NR2I U73 ( .A(N68), .B(n32), .Z(n64) );
  IVI U74 ( .A(fd_opcode[2]), .Z(n67) );
  NR2I U75 ( .A(n66), .B(n67), .Z(n62) );
  NR2I U76 ( .A(n64), .B(n63), .Z(d_PCSrc2) );
  IVI U77 ( .A(n66), .Z(n68) );
  AN3 U78 ( .A(fd_opcode[1]), .B(n68), .C(n67), .Z(d_PCSrc1) );
  IVI U79 ( .A(dx_opcode[5]), .Z(n71) );
  IVI U80 ( .A(dx_opcode[3]), .Z(n70) );
  IVI U81 ( .A(dx_opcode[1]), .Z(n69) );
  ND3 U82 ( .A(n71), .B(n70), .C(n69), .Z(n80) );
  IVI U83 ( .A(dx_opcode[4]), .Z(n78) );
  IVI U84 ( .A(dx_opcode[0]), .Z(n72) );
  IVI U85 ( .A(dx_opcode[2]), .Z(n82) );
  IVI U86 ( .A(dx_funct[4]), .Z(n73) );
  IVI U87 ( .A(dx_funct[3]), .Z(n90) );
  ND4 U88 ( .A(dx_funct[2]), .B(dx_funct[5]), .C(n41), .D(n7), .Z(n84) );
  ND2I U89 ( .A(n45), .B(n72), .Z(n77) );
  IVI U90 ( .A(dx_funct[0]), .Z(n83) );
  IVI U91 ( .A(dx_funct[2]), .Z(n74) );
  ND4 U92 ( .A(n41), .B(n83), .C(n74), .D(n73), .Z(n75) );
  IVI U93 ( .A(n75), .Z(n89) );
  IVI U94 ( .A(dx_funct[5]), .Z(n76) );
  ND3 U95 ( .A(n89), .B(n90), .C(n76), .Z(n94) );
  AO3 U96 ( .A(dx_funct[0]), .B(n84), .C(n77), .D(n94), .Z(x_ALU_Control[0])
         );
  ND2I U97 ( .A(dx_funct[5]), .B(n78), .Z(n79) );
  IVI U98 ( .A(dx_funct[1]), .Z(n85) );
  NR4 U99 ( .A(dx_opcode[0]), .B(n80), .C(n79), .D(n85), .Z(n81) );
  ND4 U100 ( .A(n82), .B(n83), .C(n7), .D(n81), .Z(n91) );
  EOI U101 ( .A(dx_opcode[0]), .B(dx_opcode[1]), .Z(n87) );
  AO7 U102 ( .A(n84), .B(n83), .C(n94), .Z(n86) );
  AO2 U103 ( .A(n45), .B(n87), .C(n86), .D(n85), .Z(n88) );
  ND2I U104 ( .A(n91), .B(n88), .Z(x_ALU_Control[1]) );
  ND2I U105 ( .A(dx_opcode[1]), .B(n46), .Z(n93) );
  AO3 U106 ( .A(dx_funct[5]), .B(n90), .C(dx_funct[1]), .D(n89), .Z(n92) );
  IVI U107 ( .A(n94), .Z(x_isSLL_SRL) );
  AO6 U108 ( .A(dx_opcode[2]), .B(n42), .C(n41), .Z(x_ALUSrc) );
  IVI U109 ( .A(n10), .Z(n97) );
  IVI U110 ( .A(xm_opcode[3]), .Z(n96) );
  IVI U111 ( .A(xm_opcode[4]), .Z(n95) );
  IVI U112 ( .A(n9), .Z(n98) );
  EOI U113 ( .A(n4), .B(n98), .Z(n100) );
  AN4 U114 ( .A(n65), .B(n34), .C(n35), .D(n100), .Z(m_MemWrite) );
  AN3 U115 ( .A(n34), .B(n3), .C(n100), .Z(m_MemRead) );
  IVI U116 ( .A(mw_opcode[3]), .Z(n103) );
  IVI U117 ( .A(mw_opcode[5]), .Z(n108) );
  ND2I U118 ( .A(n26), .B(n108), .Z(n101) );
  NR2I U119 ( .A(n109), .B(n101), .Z(n102) );
  ND2I U120 ( .A(n103), .B(n102), .Z(n106) );
  IVI U121 ( .A(n12), .Z(n105) );
  IVI U122 ( .A(n11), .Z(n104) );
  IVI U123 ( .A(n26), .Z(n112) );
  EOI U124 ( .A(n30), .B(n112), .Z(n107) );
  AN3 U125 ( .A(n44), .B(n103), .C(n107), .Z(w_MemtoReg) );
  ND2I U126 ( .A(n28), .B(n8), .Z(n111) );
  IVI U127 ( .A(mw_opcode[0]), .Z(n109) );
  ND3 U128 ( .A(n8), .B(n109), .C(n104), .Z(n110) );
  MUX21L U129 ( .A(n111), .B(n110), .S(n39), .Z(n123) );
  ND3 U130 ( .A(n29), .B(n44), .C(n112), .Z(n114) );
  ND3 U131 ( .A(n39), .B(n29), .C(n44), .Z(n113) );
  MUX21L U132 ( .A(n114), .B(n113), .S(n30), .Z(n122) );
  NR4 U133 ( .A(mw_rd[3]), .B(mw_rd[2]), .C(mw_rd[1]), .D(mw_rd[0]), .Z(n116)
         );
  NR4 U134 ( .A(mw_rt[2]), .B(mw_rt[1]), .C(mw_rt[0]), .D(mw_rd[4]), .Z(n115)
         );
  ND2I U135 ( .A(n116), .B(n115), .Z(n117) );
  NR8 U136 ( .A(n117), .B(mw_rs[4]), .C(mw_rs[3]), .D(mw_rs[2]), .E(mw_rs[1]), 
        .F(mw_rs[0]), .G(mw_rt[4]), .H(mw_rt[3]), .Z(n121) );
  OR3 U137 ( .A(mw_funct[4]), .B(mw_funct[2]), .C(mw_funct[5]), .Z(n119) );
  ND2I U138 ( .A(mw_funct[3]), .B(n38), .Z(n118) );
  NR4 U139 ( .A(n119), .B(n118), .C(mw_funct[1]), .D(mw_funct[0]), .Z(n120) );
  NR4 U140 ( .A(n123), .B(n122), .C(n121), .D(n120), .Z(w_RegWrite) );
endmodule


module mux_2x1_DATA_WIDTH5_0 ( ip1, ip0, sel, out );
  input [4:0] ip1;
  input [4:0] ip0;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n11;

  IVI U1 ( .A(n2), .Z(n1) );
  EON1P U2 ( .A(n11), .B(n1), .C(ip1[4]), .D(n3), .Z(out[4]) );
  IVI U3 ( .A(ip0[2]), .Z(n8) );
  IVI U4 ( .A(ip0[4]), .Z(n11) );
  IVI U5 ( .A(ip1[2]), .Z(n7) );
  IVI U6 ( .A(ip1[3]), .Z(n4) );
  IVI U7 ( .A(sel), .Z(n2) );
  IVI U8 ( .A(n2), .Z(n3) );
  MUX21H U9 ( .A(ip1[0]), .B(ip0[0]), .S(n5), .Z(out[0]) );
  EON1 U10 ( .A(n4), .B(n9), .C(ip0[3]), .D(n5), .Z(out[3]) );
  IVI U11 ( .A(sel), .Z(n5) );
  MUX21L U12 ( .A(n7), .B(n8), .S(n9), .Z(out[2]) );
  IVI U13 ( .A(sel), .Z(n9) );
  MUX21H U14 ( .A(ip0[1]), .B(ip1[1]), .S(sel), .Z(out[1]) );
endmodule


module mux_2x1_DATA_WIDTH5_4 ( ip1, ip0, sel, out );
  input [4:0] ip1;
  input [4:0] ip0;
  output [4:0] out;
  input sel;
  wire   n1, n2, n5, n6, n7, n8, n9, n10, n11, n12;

  ND2I U1 ( .A(ip1[2]), .B(sel), .Z(n1) );
  ND2I U2 ( .A(ip0[2]), .B(n7), .Z(n2) );
  AN2I U3 ( .A(n1), .B(n2), .Z(n11) );
  ND2I U4 ( .A(n5), .B(n6), .Z(out[0]) );
  ND2I U5 ( .A(n8), .B(n9), .Z(out[4]) );
  ND2I U6 ( .A(ip1[0]), .B(sel), .Z(n5) );
  ND2I U7 ( .A(ip0[0]), .B(n7), .Z(n6) );
  IVI U8 ( .A(sel), .Z(n7) );
  ND2I U9 ( .A(ip0[4]), .B(n7), .Z(n8) );
  ND2I U10 ( .A(ip1[4]), .B(sel), .Z(n9) );
  IVI U11 ( .A(n10), .Z(out[1]) );
  IVI U12 ( .A(n11), .Z(out[2]) );
  IVI U13 ( .A(n12), .Z(out[3]) );
  AO2P U14 ( .A(ip1[1]), .B(sel), .C(ip0[1]), .D(n7), .Z(n10) );
  AO2P U15 ( .A(ip0[3]), .B(n7), .C(ip1[3]), .D(sel), .Z(n12) );
endmodule


module mux_2x1_DATA_WIDTH5_3 ( ip1, ip0, sel, out );
  input [4:0] ip1;
  input [4:0] ip0;
  output [4:0] out;
  input sel;
  wire   n1, n2, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n22, n23;

  IVI U1 ( .A(ip0[3]), .Z(n1) );
  IVI U2 ( .A(ip1[3]), .Z(n2) );
  MUX21L U3 ( .A(n1), .B(n2), .S(sel), .Z(out[3]) );
  AN2I U4 ( .A(n5), .B(n6), .Z(out[2]) );
  ND2I U5 ( .A(n22), .B(n4), .Z(n5) );
  ND2I U6 ( .A(n21), .B(n23), .Z(n6) );
  IVI U7 ( .A(n23), .Z(n4) );
  IVI U8 ( .A(ip0[2]), .Z(n21) );
  IVI U9 ( .A(ip1[2]), .Z(n22) );
  IVI U10 ( .A(ip0[1]), .Z(n11) );
  IVI U11 ( .A(ip1[1]), .Z(n12) );
  AN2I U12 ( .A(n9), .B(n10), .Z(out[4]) );
  ND2I U13 ( .A(n13), .B(n8), .Z(n9) );
  ND2I U14 ( .A(n14), .B(n15), .Z(n10) );
  IVI U15 ( .A(n15), .Z(n8) );
  IVI U16 ( .A(ip1[4]), .Z(n13) );
  IVI U17 ( .A(ip0[4]), .Z(n14) );
  MUX21L U18 ( .A(n11), .B(n12), .S(sel), .Z(out[1]) );
  IVI U19 ( .A(sel), .Z(n15) );
  AN2I U20 ( .A(n17), .B(n18), .Z(out[0]) );
  ND2I U21 ( .A(n19), .B(n23), .Z(n17) );
  ND2I U22 ( .A(n20), .B(n8), .Z(n18) );
  IVI U23 ( .A(ip0[0]), .Z(n19) );
  IVI U24 ( .A(ip1[0]), .Z(n20) );
  IVI U25 ( .A(sel), .Z(n23) );
endmodule


module mux_2x1_DATA_WIDTH5_2 ( ip1, ip0, sel, out );
  input [4:0] ip1;
  input [4:0] ip0;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  AN2I U1 ( .A(ip1[4]), .B(n12), .Z(n1) );
  AN2I U2 ( .A(ip1[2]), .B(n12), .Z(n2) );
  IVI U3 ( .A(n15), .Z(n3) );
  B3IP U4 ( .A(sel), .Z1(n15), .Z2(n17) );
  ND2I U5 ( .A(ip1[4]), .B(n16), .Z(n4) );
  IVI U6 ( .A(n17), .Z(n5) );
  IVI U7 ( .A(n5), .Z(n6) );
  ND2I U8 ( .A(ip1[2]), .B(n16), .Z(n7) );
  ND2I U9 ( .A(n16), .B(n21), .Z(n8) );
  ND2I U10 ( .A(n14), .B(n21), .Z(n9) );
  AN2I U11 ( .A(n8), .B(n9), .Z(out[3]) );
  ND2I U12 ( .A(n16), .B(n20), .Z(n10) );
  ND2I U13 ( .A(n13), .B(n20), .Z(n11) );
  AN2I U14 ( .A(n10), .B(n11), .Z(out[1]) );
  IVI U15 ( .A(ip0[3]), .Z(n14) );
  IVI U16 ( .A(n15), .Z(n12) );
  IVI U17 ( .A(n15), .Z(n16) );
  IVI U18 ( .A(ip0[1]), .Z(n13) );
  EO1P U19 ( .A(n17), .B(n4), .C(ip0[4]), .D(n1), .Z(out[4]) );
  EO1P U20 ( .A(n17), .B(n7), .C(ip0[2]), .D(n2), .Z(out[2]) );
  EO1P U21 ( .A(n6), .B(n19), .C(ip0[0]), .D(n18), .Z(out[0]) );
  ND2I U22 ( .A(ip1[0]), .B(n3), .Z(n19) );
  IVI U23 ( .A(n19), .Z(n18) );
  ND2I U24 ( .A(ip1[1]), .B(n17), .Z(n20) );
  ND2I U25 ( .A(ip1[3]), .B(n17), .Z(n21) );
endmodule


module mux_2x1_DATA_WIDTH32_8 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4;

  IVAP U1 ( .A(n4), .Z(n1) );
  IVAP U2 ( .A(n4), .Z(n2) );
  IVI U3 ( .A(n4), .Z(n3) );
  IVI U4 ( .A(sel), .Z(n4) );
  MUX21H U5 ( .A(ip0[0]), .B(ip1[0]), .S(n3), .Z(out[0]) );
  MUX21H U6 ( .A(ip0[1]), .B(ip1[1]), .S(n3), .Z(out[1]) );
  MUX21H U7 ( .A(ip0[2]), .B(ip1[2]), .S(n3), .Z(out[2]) );
  MUX21H U8 ( .A(ip0[3]), .B(ip1[3]), .S(n3), .Z(out[3]) );
  MUX21H U9 ( .A(ip0[4]), .B(ip1[4]), .S(n2), .Z(out[4]) );
  MUX21H U10 ( .A(ip0[5]), .B(ip1[5]), .S(n2), .Z(out[5]) );
  MUX21H U11 ( .A(ip0[6]), .B(ip1[6]), .S(n2), .Z(out[6]) );
  MUX21H U12 ( .A(ip0[7]), .B(ip1[7]), .S(n2), .Z(out[7]) );
  MUX21H U13 ( .A(ip0[8]), .B(ip1[8]), .S(n2), .Z(out[8]) );
  MUX21H U14 ( .A(ip0[9]), .B(ip1[9]), .S(n2), .Z(out[9]) );
  MUX21H U15 ( .A(ip0[10]), .B(ip1[10]), .S(n2), .Z(out[10]) );
  MUX21H U16 ( .A(ip0[11]), .B(ip1[11]), .S(n2), .Z(out[11]) );
  MUX21H U17 ( .A(ip0[12]), .B(ip1[12]), .S(n2), .Z(out[12]) );
  MUX21H U18 ( .A(ip0[13]), .B(ip1[13]), .S(n2), .Z(out[13]) );
  MUX21H U19 ( .A(ip0[14]), .B(ip1[14]), .S(n2), .Z(out[14]) );
  MUX21H U20 ( .A(ip0[15]), .B(ip1[15]), .S(n2), .Z(out[15]) );
  MUX21H U21 ( .A(ip0[16]), .B(ip1[16]), .S(n2), .Z(out[16]) );
  MUX21H U22 ( .A(ip0[17]), .B(ip1[17]), .S(n2), .Z(out[17]) );
  MUX21H U23 ( .A(ip0[18]), .B(ip1[18]), .S(n1), .Z(out[18]) );
  MUX21H U24 ( .A(ip0[19]), .B(ip1[19]), .S(n1), .Z(out[19]) );
  MUX21H U25 ( .A(ip0[20]), .B(ip1[20]), .S(n1), .Z(out[20]) );
  MUX21H U26 ( .A(ip0[21]), .B(ip1[21]), .S(n1), .Z(out[21]) );
  MUX21H U27 ( .A(ip0[22]), .B(ip1[22]), .S(n1), .Z(out[22]) );
  MUX21H U28 ( .A(ip0[23]), .B(ip1[23]), .S(n1), .Z(out[23]) );
  MUX21H U29 ( .A(ip0[24]), .B(ip1[24]), .S(n1), .Z(out[24]) );
  MUX21H U30 ( .A(ip0[25]), .B(ip1[25]), .S(n1), .Z(out[25]) );
  MUX21H U31 ( .A(ip0[26]), .B(ip1[26]), .S(n1), .Z(out[26]) );
  MUX21H U32 ( .A(ip0[27]), .B(ip1[27]), .S(n1), .Z(out[27]) );
  MUX21H U33 ( .A(ip0[28]), .B(ip1[28]), .S(n1), .Z(out[28]) );
  MUX21H U34 ( .A(ip0[29]), .B(ip1[29]), .S(n1), .Z(out[29]) );
  MUX21H U35 ( .A(ip0[30]), .B(ip1[30]), .S(n1), .Z(out[30]) );
  MUX21H U36 ( .A(ip0[31]), .B(ip1[31]), .S(n1), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_7 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3;

  B5IP U1 ( .A(n3), .Z(n1) );
  B5IP U2 ( .A(n3), .Z(n2) );
  IVI U3 ( .A(sel), .Z(n3) );
  MUX21H U4 ( .A(ip0[0]), .B(ip1[0]), .S(n1), .Z(out[0]) );
  MUX21H U5 ( .A(ip0[1]), .B(ip1[1]), .S(n1), .Z(out[1]) );
  MUX21H U6 ( .A(ip0[2]), .B(ip1[2]), .S(n2), .Z(out[2]) );
  MUX21H U7 ( .A(ip0[3]), .B(ip1[3]), .S(n2), .Z(out[3]) );
  MUX21H U8 ( .A(ip0[4]), .B(ip1[4]), .S(n2), .Z(out[4]) );
  MUX21H U9 ( .A(ip0[5]), .B(ip1[5]), .S(n2), .Z(out[5]) );
  MUX21H U10 ( .A(ip0[6]), .B(ip1[6]), .S(n2), .Z(out[6]) );
  MUX21H U11 ( .A(ip0[7]), .B(ip1[7]), .S(n2), .Z(out[7]) );
  MUX21H U12 ( .A(ip0[8]), .B(ip1[8]), .S(n2), .Z(out[8]) );
  MUX21H U13 ( .A(ip0[9]), .B(ip1[9]), .S(n2), .Z(out[9]) );
  MUX21H U14 ( .A(ip0[10]), .B(ip1[10]), .S(n2), .Z(out[10]) );
  MUX21H U15 ( .A(ip0[11]), .B(ip1[11]), .S(n2), .Z(out[11]) );
  MUX21H U16 ( .A(ip0[12]), .B(ip1[12]), .S(n2), .Z(out[12]) );
  MUX21H U17 ( .A(ip0[13]), .B(ip1[13]), .S(n2), .Z(out[13]) );
  MUX21H U18 ( .A(ip0[14]), .B(ip1[14]), .S(n2), .Z(out[14]) );
  MUX21H U19 ( .A(ip0[15]), .B(ip1[15]), .S(n2), .Z(out[15]) );
  MUX21H U20 ( .A(ip0[16]), .B(ip1[16]), .S(n2), .Z(out[16]) );
  MUX21H U21 ( .A(ip0[17]), .B(ip1[17]), .S(n2), .Z(out[17]) );
  MUX21H U22 ( .A(ip0[18]), .B(ip1[18]), .S(n1), .Z(out[18]) );
  MUX21H U23 ( .A(ip0[19]), .B(ip1[19]), .S(n1), .Z(out[19]) );
  MUX21H U24 ( .A(ip0[20]), .B(ip1[20]), .S(n1), .Z(out[20]) );
  MUX21H U25 ( .A(ip0[21]), .B(ip1[21]), .S(n1), .Z(out[21]) );
  MUX21H U26 ( .A(ip0[22]), .B(ip1[22]), .S(n1), .Z(out[22]) );
  MUX21H U27 ( .A(ip0[23]), .B(ip1[23]), .S(n1), .Z(out[23]) );
  MUX21H U28 ( .A(ip0[24]), .B(ip1[24]), .S(n1), .Z(out[24]) );
  MUX21H U29 ( .A(ip0[25]), .B(ip1[25]), .S(n1), .Z(out[25]) );
  MUX21H U30 ( .A(ip0[26]), .B(ip1[26]), .S(n1), .Z(out[26]) );
  MUX21H U31 ( .A(ip0[27]), .B(ip1[27]), .S(n1), .Z(out[27]) );
  MUX21H U32 ( .A(ip0[28]), .B(ip1[28]), .S(n1), .Z(out[28]) );
  MUX21H U33 ( .A(ip0[29]), .B(ip1[29]), .S(n1), .Z(out[29]) );
  MUX21H U34 ( .A(ip0[30]), .B(ip1[30]), .S(n1), .Z(out[30]) );
  MUX21H U35 ( .A(ip0[31]), .B(ip1[31]), .S(n1), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH5_1 ( ip1, ip0, sel, out );
  input [4:0] ip1;
  input [4:0] ip0;
  output [4:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  MUX21HP U1 ( .A(ip0[3]), .B(ip1[3]), .S(n5), .Z(out[3]) );
  MUX21HP U2 ( .A(ip0[4]), .B(ip1[4]), .S(n5), .Z(out[4]) );
  IVI U3 ( .A(sel), .Z(n1) );
  IVI U4 ( .A(n1), .Z(n2) );
  IVI U5 ( .A(n4), .Z(n3) );
  IVI U6 ( .A(sel), .Z(n4) );
  IVI U7 ( .A(n4), .Z(n5) );
  ND2I U8 ( .A(ip1[0]), .B(sel), .Z(n7) );
  ND2I U9 ( .A(ip0[0]), .B(n1), .Z(n6) );
  ND2I U10 ( .A(n7), .B(n6), .Z(out[0]) );
  ND2I U11 ( .A(ip1[1]), .B(n3), .Z(n9) );
  ND2I U12 ( .A(ip0[1]), .B(n4), .Z(n8) );
  ND2I U13 ( .A(n9), .B(n8), .Z(out[1]) );
  MUX21H U14 ( .A(ip0[2]), .B(ip1[2]), .S(n2), .Z(out[2]) );
endmodule


module gpr ( clk, RegWrite, rd_addr1, rd_addr2, wr_addr, wr_data, rd_data1, 
        rd_data2 );
  input [4:0] rd_addr1;
  input [4:0] rd_addr2;
  input [4:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_data1;
  output [31:0] rd_data2;
  input clk, RegWrite;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, \gpr[1][31] ,
         \gpr[1][30] , \gpr[1][29] , \gpr[1][28] , \gpr[1][27] , \gpr[1][26] ,
         \gpr[1][25] , \gpr[1][24] , \gpr[1][23] , \gpr[1][22] , \gpr[1][21] ,
         \gpr[1][20] , \gpr[1][19] , \gpr[1][18] , \gpr[1][17] , \gpr[1][16] ,
         \gpr[1][15] , \gpr[1][14] , \gpr[1][13] , \gpr[1][12] , \gpr[1][11] ,
         \gpr[1][10] , \gpr[1][9] , \gpr[1][8] , \gpr[1][7] , \gpr[1][6] ,
         \gpr[1][5] , \gpr[1][4] , \gpr[1][3] , \gpr[1][2] , \gpr[1][1] ,
         \gpr[1][0] , \gpr[2][31] , \gpr[2][30] , \gpr[2][29] , \gpr[2][28] ,
         \gpr[2][27] , \gpr[2][26] , \gpr[2][25] , \gpr[2][24] , \gpr[2][23] ,
         \gpr[2][22] , \gpr[2][21] , \gpr[2][20] , \gpr[2][19] , \gpr[2][18] ,
         \gpr[2][17] , \gpr[2][16] , \gpr[2][15] , \gpr[2][14] , \gpr[2][13] ,
         \gpr[2][12] , \gpr[2][11] , \gpr[2][10] , \gpr[2][9] , \gpr[2][8] ,
         \gpr[2][7] , \gpr[2][6] , \gpr[2][5] , \gpr[2][4] , \gpr[2][3] ,
         \gpr[2][2] , \gpr[2][1] , \gpr[2][0] , \gpr[3][31] , \gpr[3][30] ,
         \gpr[3][29] , \gpr[3][28] , \gpr[3][27] , \gpr[3][26] , \gpr[3][25] ,
         \gpr[3][24] , \gpr[3][23] , \gpr[3][22] , \gpr[3][21] , \gpr[3][20] ,
         \gpr[3][19] , \gpr[3][18] , \gpr[3][17] , \gpr[3][16] , \gpr[3][15] ,
         \gpr[3][14] , \gpr[3][13] , \gpr[3][12] , \gpr[3][11] , \gpr[3][10] ,
         \gpr[3][9] , \gpr[3][8] , \gpr[3][7] , \gpr[3][6] , \gpr[3][5] ,
         \gpr[3][4] , \gpr[3][3] , \gpr[3][2] , \gpr[3][1] , \gpr[3][0] ,
         \gpr[4][31] , \gpr[4][30] , \gpr[4][29] , \gpr[4][28] , \gpr[4][27] ,
         \gpr[4][26] , \gpr[4][25] , \gpr[4][24] , \gpr[4][23] , \gpr[4][22] ,
         \gpr[4][21] , \gpr[4][20] , \gpr[4][19] , \gpr[4][18] , \gpr[4][17] ,
         \gpr[4][16] , \gpr[4][15] , \gpr[4][14] , \gpr[4][13] , \gpr[4][12] ,
         \gpr[4][11] , \gpr[4][10] , \gpr[4][9] , \gpr[4][8] , \gpr[4][7] ,
         \gpr[4][6] , \gpr[4][5] , \gpr[4][4] , \gpr[4][3] , \gpr[4][2] ,
         \gpr[4][1] , \gpr[4][0] , \gpr[5][31] , \gpr[5][30] , \gpr[5][29] ,
         \gpr[5][28] , \gpr[5][27] , \gpr[5][26] , \gpr[5][25] , \gpr[5][24] ,
         \gpr[5][23] , \gpr[5][22] , \gpr[5][21] , \gpr[5][20] , \gpr[5][19] ,
         \gpr[5][18] , \gpr[5][17] , \gpr[5][16] , \gpr[5][15] , \gpr[5][14] ,
         \gpr[5][13] , \gpr[5][12] , \gpr[5][11] , \gpr[5][10] , \gpr[5][9] ,
         \gpr[5][8] , \gpr[5][7] , \gpr[5][6] , \gpr[5][5] , \gpr[5][4] ,
         \gpr[5][3] , \gpr[5][2] , \gpr[5][1] , \gpr[5][0] , \gpr[6][31] ,
         \gpr[6][30] , \gpr[6][29] , \gpr[6][28] , \gpr[6][27] , \gpr[6][26] ,
         \gpr[6][25] , \gpr[6][24] , \gpr[6][23] , \gpr[6][22] , \gpr[6][21] ,
         \gpr[6][20] , \gpr[6][19] , \gpr[6][18] , \gpr[6][17] , \gpr[6][16] ,
         \gpr[6][15] , \gpr[6][14] , \gpr[6][13] , \gpr[6][12] , \gpr[6][11] ,
         \gpr[6][10] , \gpr[6][9] , \gpr[6][8] , \gpr[6][7] , \gpr[6][6] ,
         \gpr[6][5] , \gpr[6][4] , \gpr[6][3] , \gpr[6][2] , \gpr[6][1] ,
         \gpr[6][0] , \gpr[7][31] , \gpr[7][30] , \gpr[7][29] , \gpr[7][28] ,
         \gpr[7][27] , \gpr[7][26] , \gpr[7][25] , \gpr[7][24] , \gpr[7][23] ,
         \gpr[7][22] , \gpr[7][21] , \gpr[7][20] , \gpr[7][19] , \gpr[7][18] ,
         \gpr[7][17] , \gpr[7][16] , \gpr[7][15] , \gpr[7][14] , \gpr[7][13] ,
         \gpr[7][12] , \gpr[7][11] , \gpr[7][10] , \gpr[7][9] , \gpr[7][8] ,
         \gpr[7][7] , \gpr[7][6] , \gpr[7][5] , \gpr[7][4] , \gpr[7][3] ,
         \gpr[7][2] , \gpr[7][1] , \gpr[7][0] , \gpr[8][31] , \gpr[8][30] ,
         \gpr[8][29] , \gpr[8][28] , \gpr[8][27] , \gpr[8][26] , \gpr[8][25] ,
         \gpr[8][24] , \gpr[8][23] , \gpr[8][22] , \gpr[8][21] , \gpr[8][20] ,
         \gpr[8][19] , \gpr[8][18] , \gpr[8][17] , \gpr[8][16] , \gpr[8][15] ,
         \gpr[8][14] , \gpr[8][13] , \gpr[8][12] , \gpr[8][11] , \gpr[8][10] ,
         \gpr[8][9] , \gpr[8][8] , \gpr[8][7] , \gpr[8][6] , \gpr[8][5] ,
         \gpr[8][4] , \gpr[8][3] , \gpr[8][2] , \gpr[8][1] , \gpr[8][0] ,
         \gpr[9][31] , \gpr[9][30] , \gpr[9][29] , \gpr[9][28] , \gpr[9][27] ,
         \gpr[9][26] , \gpr[9][25] , \gpr[9][24] , \gpr[9][23] , \gpr[9][22] ,
         \gpr[9][21] , \gpr[9][20] , \gpr[9][19] , \gpr[9][18] , \gpr[9][17] ,
         \gpr[9][16] , \gpr[9][15] , \gpr[9][14] , \gpr[9][13] , \gpr[9][12] ,
         \gpr[9][11] , \gpr[9][10] , \gpr[9][9] , \gpr[9][8] , \gpr[9][7] ,
         \gpr[9][6] , \gpr[9][5] , \gpr[9][4] , \gpr[9][3] , \gpr[9][2] ,
         \gpr[9][1] , \gpr[9][0] , \gpr[10][31] , \gpr[10][30] , \gpr[10][29] ,
         \gpr[10][28] , \gpr[10][27] , \gpr[10][26] , \gpr[10][25] ,
         \gpr[10][24] , \gpr[10][23] , \gpr[10][22] , \gpr[10][21] ,
         \gpr[10][20] , \gpr[10][19] , \gpr[10][18] , \gpr[10][17] ,
         \gpr[10][16] , \gpr[10][15] , \gpr[10][14] , \gpr[10][13] ,
         \gpr[10][12] , \gpr[10][11] , \gpr[10][10] , \gpr[10][9] ,
         \gpr[10][8] , \gpr[10][7] , \gpr[10][6] , \gpr[10][5] , \gpr[10][4] ,
         \gpr[10][3] , \gpr[10][2] , \gpr[10][1] , \gpr[10][0] , \gpr[11][31] ,
         \gpr[11][30] , \gpr[11][29] , \gpr[11][28] , \gpr[11][27] ,
         \gpr[11][26] , \gpr[11][25] , \gpr[11][24] , \gpr[11][23] ,
         \gpr[11][22] , \gpr[11][21] , \gpr[11][20] , \gpr[11][19] ,
         \gpr[11][18] , \gpr[11][17] , \gpr[11][16] , \gpr[11][15] ,
         \gpr[11][14] , \gpr[11][13] , \gpr[11][12] , \gpr[11][11] ,
         \gpr[11][10] , \gpr[11][9] , \gpr[11][8] , \gpr[11][7] , \gpr[11][6] ,
         \gpr[11][5] , \gpr[11][4] , \gpr[11][3] , \gpr[11][2] , \gpr[11][1] ,
         \gpr[11][0] , \gpr[12][31] , \gpr[12][30] , \gpr[12][29] ,
         \gpr[12][28] , \gpr[12][27] , \gpr[12][26] , \gpr[12][25] ,
         \gpr[12][24] , \gpr[12][23] , \gpr[12][22] , \gpr[12][21] ,
         \gpr[12][20] , \gpr[12][19] , \gpr[12][18] , \gpr[12][17] ,
         \gpr[12][16] , \gpr[12][15] , \gpr[12][14] , \gpr[12][13] ,
         \gpr[12][12] , \gpr[12][11] , \gpr[12][10] , \gpr[12][9] ,
         \gpr[12][8] , \gpr[12][7] , \gpr[12][6] , \gpr[12][5] , \gpr[12][4] ,
         \gpr[12][3] , \gpr[12][2] , \gpr[12][1] , \gpr[12][0] , \gpr[13][31] ,
         \gpr[13][30] , \gpr[13][29] , \gpr[13][28] , \gpr[13][27] ,
         \gpr[13][26] , \gpr[13][25] , \gpr[13][24] , \gpr[13][23] ,
         \gpr[13][22] , \gpr[13][21] , \gpr[13][20] , \gpr[13][19] ,
         \gpr[13][18] , \gpr[13][17] , \gpr[13][16] , \gpr[13][15] ,
         \gpr[13][14] , \gpr[13][13] , \gpr[13][12] , \gpr[13][11] ,
         \gpr[13][10] , \gpr[13][9] , \gpr[13][8] , \gpr[13][7] , \gpr[13][6] ,
         \gpr[13][5] , \gpr[13][4] , \gpr[13][3] , \gpr[13][2] , \gpr[13][1] ,
         \gpr[13][0] , \gpr[14][31] , \gpr[14][30] , \gpr[14][29] ,
         \gpr[14][28] , \gpr[14][27] , \gpr[14][26] , \gpr[14][25] ,
         \gpr[14][24] , \gpr[14][23] , \gpr[14][22] , \gpr[14][21] ,
         \gpr[14][20] , \gpr[14][19] , \gpr[14][18] , \gpr[14][17] ,
         \gpr[14][16] , \gpr[14][15] , \gpr[14][14] , \gpr[14][13] ,
         \gpr[14][12] , \gpr[14][11] , \gpr[14][10] , \gpr[14][9] ,
         \gpr[14][8] , \gpr[14][7] , \gpr[14][6] , \gpr[14][5] , \gpr[14][4] ,
         \gpr[14][3] , \gpr[14][2] , \gpr[14][1] , \gpr[14][0] , \gpr[15][31] ,
         \gpr[15][30] , \gpr[15][29] , \gpr[15][28] , \gpr[15][27] ,
         \gpr[15][26] , \gpr[15][25] , \gpr[15][24] , \gpr[15][23] ,
         \gpr[15][22] , \gpr[15][21] , \gpr[15][20] , \gpr[15][19] ,
         \gpr[15][18] , \gpr[15][17] , \gpr[15][16] , \gpr[15][15] ,
         \gpr[15][14] , \gpr[15][13] , \gpr[15][12] , \gpr[15][11] ,
         \gpr[15][10] , \gpr[15][9] , \gpr[15][8] , \gpr[15][7] , \gpr[15][6] ,
         \gpr[15][5] , \gpr[15][4] , \gpr[15][3] , \gpr[15][2] , \gpr[15][1] ,
         \gpr[15][0] , \gpr[16][31] , \gpr[16][30] , \gpr[16][29] ,
         \gpr[16][28] , \gpr[16][27] , \gpr[16][26] , \gpr[16][25] ,
         \gpr[16][24] , \gpr[16][23] , \gpr[16][22] , \gpr[16][21] ,
         \gpr[16][20] , \gpr[16][19] , \gpr[16][18] , \gpr[16][17] ,
         \gpr[16][16] , \gpr[16][15] , \gpr[16][14] , \gpr[16][13] ,
         \gpr[16][12] , \gpr[16][11] , \gpr[16][10] , \gpr[16][9] ,
         \gpr[16][8] , \gpr[16][7] , \gpr[16][6] , \gpr[16][5] , \gpr[16][4] ,
         \gpr[16][3] , \gpr[16][2] , \gpr[16][1] , \gpr[16][0] , \gpr[17][31] ,
         \gpr[17][30] , \gpr[17][29] , \gpr[17][28] , \gpr[17][27] ,
         \gpr[17][26] , \gpr[17][25] , \gpr[17][24] , \gpr[17][23] ,
         \gpr[17][22] , \gpr[17][21] , \gpr[17][20] , \gpr[17][19] ,
         \gpr[17][18] , \gpr[17][17] , \gpr[17][16] , \gpr[17][15] ,
         \gpr[17][14] , \gpr[17][13] , \gpr[17][12] , \gpr[17][11] ,
         \gpr[17][10] , \gpr[17][9] , \gpr[17][8] , \gpr[17][7] , \gpr[17][6] ,
         \gpr[17][5] , \gpr[17][4] , \gpr[17][3] , \gpr[17][2] , \gpr[17][1] ,
         \gpr[17][0] , \gpr[18][31] , \gpr[18][30] , \gpr[18][29] ,
         \gpr[18][28] , \gpr[18][27] , \gpr[18][26] , \gpr[18][25] ,
         \gpr[18][24] , \gpr[18][23] , \gpr[18][22] , \gpr[18][21] ,
         \gpr[18][20] , \gpr[18][19] , \gpr[18][18] , \gpr[18][17] ,
         \gpr[18][16] , \gpr[18][15] , \gpr[18][14] , \gpr[18][13] ,
         \gpr[18][12] , \gpr[18][11] , \gpr[18][10] , \gpr[18][9] ,
         \gpr[18][8] , \gpr[18][7] , \gpr[18][6] , \gpr[18][5] , \gpr[18][4] ,
         \gpr[18][3] , \gpr[18][2] , \gpr[18][1] , \gpr[18][0] , \gpr[19][31] ,
         \gpr[19][30] , \gpr[19][29] , \gpr[19][28] , \gpr[19][27] ,
         \gpr[19][26] , \gpr[19][25] , \gpr[19][24] , \gpr[19][23] ,
         \gpr[19][22] , \gpr[19][21] , \gpr[19][20] , \gpr[19][19] ,
         \gpr[19][18] , \gpr[19][17] , \gpr[19][16] , \gpr[19][15] ,
         \gpr[19][14] , \gpr[19][13] , \gpr[19][12] , \gpr[19][11] ,
         \gpr[19][10] , \gpr[19][9] , \gpr[19][8] , \gpr[19][7] , \gpr[19][6] ,
         \gpr[19][5] , \gpr[19][4] , \gpr[19][3] , \gpr[19][2] , \gpr[19][1] ,
         \gpr[19][0] , \gpr[20][31] , \gpr[20][30] , \gpr[20][29] ,
         \gpr[20][28] , \gpr[20][27] , \gpr[20][26] , \gpr[20][25] ,
         \gpr[20][24] , \gpr[20][23] , \gpr[20][22] , \gpr[20][21] ,
         \gpr[20][20] , \gpr[20][19] , \gpr[20][18] , \gpr[20][17] ,
         \gpr[20][16] , \gpr[20][15] , \gpr[20][14] , \gpr[20][13] ,
         \gpr[20][12] , \gpr[20][11] , \gpr[20][10] , \gpr[20][9] ,
         \gpr[20][8] , \gpr[20][7] , \gpr[20][6] , \gpr[20][5] , \gpr[20][4] ,
         \gpr[20][3] , \gpr[20][2] , \gpr[20][1] , \gpr[20][0] , \gpr[21][31] ,
         \gpr[21][30] , \gpr[21][29] , \gpr[21][28] , \gpr[21][27] ,
         \gpr[21][26] , \gpr[21][25] , \gpr[21][24] , \gpr[21][23] ,
         \gpr[21][22] , \gpr[21][21] , \gpr[21][20] , \gpr[21][19] ,
         \gpr[21][18] , \gpr[21][17] , \gpr[21][16] , \gpr[21][15] ,
         \gpr[21][14] , \gpr[21][13] , \gpr[21][12] , \gpr[21][11] ,
         \gpr[21][10] , \gpr[21][9] , \gpr[21][8] , \gpr[21][7] , \gpr[21][6] ,
         \gpr[21][5] , \gpr[21][4] , \gpr[21][3] , \gpr[21][2] , \gpr[21][1] ,
         \gpr[21][0] , \gpr[22][31] , \gpr[22][30] , \gpr[22][29] ,
         \gpr[22][28] , \gpr[22][27] , \gpr[22][26] , \gpr[22][25] ,
         \gpr[22][24] , \gpr[22][23] , \gpr[22][22] , \gpr[22][21] ,
         \gpr[22][20] , \gpr[22][19] , \gpr[22][18] , \gpr[22][17] ,
         \gpr[22][16] , \gpr[22][15] , \gpr[22][14] , \gpr[22][13] ,
         \gpr[22][12] , \gpr[22][11] , \gpr[22][10] , \gpr[22][9] ,
         \gpr[22][8] , \gpr[22][7] , \gpr[22][6] , \gpr[22][5] , \gpr[22][4] ,
         \gpr[22][3] , \gpr[22][2] , \gpr[22][1] , \gpr[22][0] , \gpr[23][31] ,
         \gpr[23][30] , \gpr[23][29] , \gpr[23][28] , \gpr[23][27] ,
         \gpr[23][26] , \gpr[23][25] , \gpr[23][24] , \gpr[23][23] ,
         \gpr[23][22] , \gpr[23][21] , \gpr[23][20] , \gpr[23][19] ,
         \gpr[23][18] , \gpr[23][17] , \gpr[23][16] , \gpr[23][15] ,
         \gpr[23][14] , \gpr[23][13] , \gpr[23][12] , \gpr[23][11] ,
         \gpr[23][10] , \gpr[23][9] , \gpr[23][8] , \gpr[23][7] , \gpr[23][6] ,
         \gpr[23][5] , \gpr[23][4] , \gpr[23][3] , \gpr[23][2] , \gpr[23][1] ,
         \gpr[23][0] , \gpr[24][31] , \gpr[24][30] , \gpr[24][29] ,
         \gpr[24][28] , \gpr[24][27] , \gpr[24][26] , \gpr[24][25] ,
         \gpr[24][24] , \gpr[24][23] , \gpr[24][22] , \gpr[24][21] ,
         \gpr[24][20] , \gpr[24][19] , \gpr[24][18] , \gpr[24][17] ,
         \gpr[24][16] , \gpr[24][15] , \gpr[24][14] , \gpr[24][13] ,
         \gpr[24][12] , \gpr[24][11] , \gpr[24][10] , \gpr[24][9] ,
         \gpr[24][8] , \gpr[24][7] , \gpr[24][6] , \gpr[24][5] , \gpr[24][4] ,
         \gpr[24][3] , \gpr[24][2] , \gpr[24][1] , \gpr[24][0] , \gpr[25][31] ,
         \gpr[25][30] , \gpr[25][29] , \gpr[25][28] , \gpr[25][27] ,
         \gpr[25][26] , \gpr[25][25] , \gpr[25][24] , \gpr[25][23] ,
         \gpr[25][22] , \gpr[25][21] , \gpr[25][20] , \gpr[25][19] ,
         \gpr[25][18] , \gpr[25][17] , \gpr[25][16] , \gpr[25][15] ,
         \gpr[25][14] , \gpr[25][13] , \gpr[25][12] , \gpr[25][11] ,
         \gpr[25][10] , \gpr[25][9] , \gpr[25][8] , \gpr[25][7] , \gpr[25][6] ,
         \gpr[25][5] , \gpr[25][4] , \gpr[25][3] , \gpr[25][2] , \gpr[25][1] ,
         \gpr[25][0] , \gpr[26][31] , \gpr[26][30] , \gpr[26][29] ,
         \gpr[26][28] , \gpr[26][27] , \gpr[26][26] , \gpr[26][25] ,
         \gpr[26][24] , \gpr[26][23] , \gpr[26][22] , \gpr[26][21] ,
         \gpr[26][20] , \gpr[26][19] , \gpr[26][18] , \gpr[26][17] ,
         \gpr[26][16] , \gpr[26][15] , \gpr[26][14] , \gpr[26][13] ,
         \gpr[26][12] , \gpr[26][11] , \gpr[26][10] , \gpr[26][9] ,
         \gpr[26][8] , \gpr[26][7] , \gpr[26][6] , \gpr[26][5] , \gpr[26][4] ,
         \gpr[26][3] , \gpr[26][2] , \gpr[26][1] , \gpr[26][0] , \gpr[27][31] ,
         \gpr[27][30] , \gpr[27][29] , \gpr[27][28] , \gpr[27][27] ,
         \gpr[27][26] , \gpr[27][25] , \gpr[27][24] , \gpr[27][23] ,
         \gpr[27][22] , \gpr[27][21] , \gpr[27][20] , \gpr[27][19] ,
         \gpr[27][18] , \gpr[27][17] , \gpr[27][16] , \gpr[27][15] ,
         \gpr[27][14] , \gpr[27][13] , \gpr[27][12] , \gpr[27][11] ,
         \gpr[27][10] , \gpr[27][9] , \gpr[27][8] , \gpr[27][7] , \gpr[27][6] ,
         \gpr[27][5] , \gpr[27][4] , \gpr[27][3] , \gpr[27][2] , \gpr[27][1] ,
         \gpr[27][0] , \gpr[28][31] , \gpr[28][30] , \gpr[28][29] ,
         \gpr[28][28] , \gpr[28][27] , \gpr[28][26] , \gpr[28][25] ,
         \gpr[28][24] , \gpr[28][23] , \gpr[28][22] , \gpr[28][21] ,
         \gpr[28][20] , \gpr[28][19] , \gpr[28][18] , \gpr[28][17] ,
         \gpr[28][16] , \gpr[28][15] , \gpr[28][14] , \gpr[28][13] ,
         \gpr[28][12] , \gpr[28][11] , \gpr[28][10] , \gpr[28][9] ,
         \gpr[28][8] , \gpr[28][7] , \gpr[28][6] , \gpr[28][5] , \gpr[28][4] ,
         \gpr[28][3] , \gpr[28][2] , \gpr[28][1] , \gpr[28][0] , \gpr[29][31] ,
         \gpr[29][30] , \gpr[29][29] , \gpr[29][28] , \gpr[29][27] ,
         \gpr[29][26] , \gpr[29][25] , \gpr[29][24] , \gpr[29][23] ,
         \gpr[29][22] , \gpr[29][21] , \gpr[29][20] , \gpr[29][19] ,
         \gpr[29][18] , \gpr[29][17] , \gpr[29][16] , \gpr[29][15] ,
         \gpr[29][14] , \gpr[29][13] , \gpr[29][12] , \gpr[29][11] ,
         \gpr[29][10] , \gpr[29][9] , \gpr[29][8] , \gpr[29][7] , \gpr[29][6] ,
         \gpr[29][5] , \gpr[29][4] , \gpr[29][3] , \gpr[29][2] , \gpr[29][1] ,
         \gpr[29][0] , \gpr[30][31] , \gpr[30][30] , \gpr[30][29] ,
         \gpr[30][28] , \gpr[30][27] , \gpr[30][26] , \gpr[30][25] ,
         \gpr[30][24] , \gpr[30][23] , \gpr[30][22] , \gpr[30][21] ,
         \gpr[30][20] , \gpr[30][19] , \gpr[30][18] , \gpr[30][17] ,
         \gpr[30][16] , \gpr[30][15] , \gpr[30][14] , \gpr[30][13] ,
         \gpr[30][12] , \gpr[30][11] , \gpr[30][10] , \gpr[30][9] ,
         \gpr[30][8] , \gpr[30][7] , \gpr[30][6] , \gpr[30][5] , \gpr[30][4] ,
         \gpr[30][3] , \gpr[30][2] , \gpr[30][1] , \gpr[30][0] , \gpr[31][31] ,
         \gpr[31][30] , \gpr[31][29] , \gpr[31][28] , \gpr[31][27] ,
         \gpr[31][26] , \gpr[31][25] , \gpr[31][24] , \gpr[31][23] ,
         \gpr[31][22] , \gpr[31][21] , \gpr[31][20] , \gpr[31][19] ,
         \gpr[31][18] , \gpr[31][17] , \gpr[31][16] , \gpr[31][15] ,
         \gpr[31][14] , \gpr[31][13] , \gpr[31][12] , \gpr[31][11] ,
         \gpr[31][10] , \gpr[31][9] , \gpr[31][8] , \gpr[31][7] , \gpr[31][6] ,
         \gpr[31][5] , \gpr[31][4] , \gpr[31][3] , \gpr[31][2] , \gpr[31][1] ,
         \gpr[31][0] , N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475;
  assign N13 = rd_addr1[0];
  assign N14 = rd_addr1[1];
  assign N15 = rd_addr1[2];
  assign N16 = rd_addr1[3];
  assign N17 = rd_addr1[4];
  assign N18 = rd_addr2[0];
  assign N19 = rd_addr2[1];
  assign N20 = rd_addr2[2];
  assign N21 = rd_addr2[3];
  assign N22 = rd_addr2[4];

  FD1 \gpr_reg[1][31]  ( .D(n1139), .CP(clk), .Q(\gpr[1][31] ), .QN(n6) );
  FD1 \gpr_reg[1][30]  ( .D(n1138), .CP(clk), .Q(\gpr[1][30] ), .QN(n7) );
  FD1 \gpr_reg[1][29]  ( .D(n1137), .CP(clk), .Q(\gpr[1][29] ), .QN(n8) );
  FD1 \gpr_reg[1][28]  ( .D(n1136), .CP(clk), .Q(\gpr[1][28] ), .QN(n9) );
  FD1 \gpr_reg[1][27]  ( .D(n1135), .CP(clk), .Q(\gpr[1][27] ), .QN(n10) );
  FD1 \gpr_reg[1][26]  ( .D(n1134), .CP(clk), .Q(\gpr[1][26] ), .QN(n1189) );
  FD1 \gpr_reg[1][25]  ( .D(n1133), .CP(clk), .Q(\gpr[1][25] ), .QN(n11) );
  FD1 \gpr_reg[1][24]  ( .D(n1132), .CP(clk), .Q(\gpr[1][24] ), .QN(n12) );
  FD1 \gpr_reg[1][23]  ( .D(n1131), .CP(clk), .Q(\gpr[1][23] ), .QN(n13) );
  FD1 \gpr_reg[1][22]  ( .D(n1130), .CP(clk), .Q(\gpr[1][22] ), .QN(n1188) );
  FD1 \gpr_reg[1][21]  ( .D(n1129), .CP(clk), .Q(\gpr[1][21] ), .QN(n14) );
  FD1 \gpr_reg[1][20]  ( .D(n1128), .CP(clk), .Q(\gpr[1][20] ), .QN(n1187) );
  FD1 \gpr_reg[1][19]  ( .D(n1127), .CP(clk), .Q(\gpr[1][19] ), .QN(n15) );
  FD1 \gpr_reg[1][18]  ( .D(n1126), .CP(clk), .Q(\gpr[1][18] ), .QN(n1186) );
  FD1 \gpr_reg[1][17]  ( .D(n1125), .CP(clk), .Q(\gpr[1][17] ), .QN(n16) );
  FD1 \gpr_reg[1][16]  ( .D(n1124), .CP(clk), .Q(\gpr[1][16] ), .QN(n17) );
  FD1 \gpr_reg[1][15]  ( .D(n1123), .CP(clk), .Q(\gpr[1][15] ), .QN(n18) );
  FD1 \gpr_reg[1][14]  ( .D(n1122), .CP(clk), .Q(\gpr[1][14] ), .QN(n1185) );
  FD1 \gpr_reg[1][13]  ( .D(n1121), .CP(clk), .Q(\gpr[1][13] ), .QN(n19) );
  FD1 \gpr_reg[1][12]  ( .D(n1120), .CP(clk), .Q(\gpr[1][12] ), .QN(n1184) );
  FD1 \gpr_reg[1][11]  ( .D(n1119), .CP(clk), .Q(\gpr[1][11] ), .QN(n3) );
  FD1 \gpr_reg[1][10]  ( .D(n1118), .CP(clk), .Q(\gpr[1][10] ), .QN(n1183) );
  FD1 \gpr_reg[1][9]  ( .D(n1117), .CP(clk), .Q(\gpr[1][9] ), .QN(n1182) );
  FD1 \gpr_reg[1][8]  ( .D(n1116), .CP(clk), .Q(\gpr[1][8] ), .QN(n4) );
  FD1 \gpr_reg[1][7]  ( .D(n1115), .CP(clk), .Q(\gpr[1][7] ), .QN(n1181) );
  FD1 \gpr_reg[1][5]  ( .D(n1113), .CP(clk), .Q(\gpr[1][5] ), .QN(n5) );
  FD1 \gpr_reg[1][3]  ( .D(n1111), .CP(clk), .Q(\gpr[1][3] ), .QN(n1180) );
  FD1 \gpr_reg[1][2]  ( .D(n1110), .CP(clk), .Q(\gpr[1][2] ), .QN(n142) );
  FD1 \gpr_reg[1][1]  ( .D(n1109), .CP(clk), .Q(\gpr[1][1] ), .QN(n1160) );
  FD1 \gpr_reg[1][0]  ( .D(n1108), .CP(clk), .Q(\gpr[1][0] ), .QN(n1159) );
  FD1 \gpr_reg[2][31]  ( .D(n1107), .CP(clk), .Q(\gpr[2][31] ), .QN(n1218) );
  FD1 \gpr_reg[2][30]  ( .D(n1106), .CP(clk), .Q(\gpr[2][30] ), .QN(n1217) );
  FD1 \gpr_reg[2][29]  ( .D(n1105), .CP(clk), .Q(\gpr[2][29] ), .QN(n1216) );
  FD1 \gpr_reg[2][28]  ( .D(n1104), .CP(clk), .Q(\gpr[2][28] ), .QN(n1215) );
  FD1 \gpr_reg[2][27]  ( .D(n1103), .CP(clk), .Q(\gpr[2][27] ), .QN(n1214) );
  FD1 \gpr_reg[2][26]  ( .D(n1102), .CP(clk), .Q(\gpr[2][26] ), .QN(n1213) );
  FD1 \gpr_reg[2][25]  ( .D(n1101), .CP(clk), .Q(\gpr[2][25] ), .QN(n1212) );
  FD1 \gpr_reg[2][24]  ( .D(n1100), .CP(clk), .Q(\gpr[2][24] ), .QN(n1211) );
  FD1 \gpr_reg[2][23]  ( .D(n1099), .CP(clk), .Q(\gpr[2][23] ), .QN(n1210) );
  FD1 \gpr_reg[2][22]  ( .D(n1098), .CP(clk), .Q(\gpr[2][22] ), .QN(n1209) );
  FD1 \gpr_reg[2][21]  ( .D(n1097), .CP(clk), .Q(\gpr[2][21] ), .QN(n1208) );
  FD1 \gpr_reg[2][20]  ( .D(n1096), .CP(clk), .Q(\gpr[2][20] ), .QN(n1207) );
  FD1 \gpr_reg[2][19]  ( .D(n1095), .CP(clk), .Q(\gpr[2][19] ), .QN(n1206) );
  FD1 \gpr_reg[2][18]  ( .D(n1094), .CP(clk), .Q(\gpr[2][18] ), .QN(n1205) );
  FD1 \gpr_reg[2][17]  ( .D(n1093), .CP(clk), .Q(\gpr[2][17] ), .QN(n1204) );
  FD1 \gpr_reg[2][16]  ( .D(n1092), .CP(clk), .Q(\gpr[2][16] ), .QN(n1203) );
  FD1 \gpr_reg[2][15]  ( .D(n1091), .CP(clk), .Q(\gpr[2][15] ), .QN(n1202) );
  FD1 \gpr_reg[2][14]  ( .D(n1090), .CP(clk), .Q(\gpr[2][14] ), .QN(n1201) );
  FD1 \gpr_reg[2][13]  ( .D(n1089), .CP(clk), .Q(\gpr[2][13] ), .QN(n1200) );
  FD1 \gpr_reg[2][12]  ( .D(n1088), .CP(clk), .Q(\gpr[2][12] ), .QN(n1199) );
  FD1 \gpr_reg[2][11]  ( .D(n1087), .CP(clk), .Q(\gpr[2][11] ), .QN(n1198) );
  FD1 \gpr_reg[2][10]  ( .D(n1086), .CP(clk), .Q(\gpr[2][10] ), .QN(n1197) );
  FD1 \gpr_reg[2][9]  ( .D(n1085), .CP(clk), .Q(\gpr[2][9] ), .QN(n1196) );
  FD1 \gpr_reg[2][8]  ( .D(n1084), .CP(clk), .Q(\gpr[2][8] ), .QN(n1195) );
  FD1 \gpr_reg[2][7]  ( .D(n1083), .CP(clk), .Q(\gpr[2][7] ), .QN(n1194) );
  FD1 \gpr_reg[2][6]  ( .D(n1082), .CP(clk), .Q(\gpr[2][6] ), .QN(n1193) );
  FD1 \gpr_reg[2][5]  ( .D(n1081), .CP(clk), .Q(\gpr[2][5] ), .QN(n1192) );
  FD1 \gpr_reg[2][4]  ( .D(n1080), .CP(clk), .Q(\gpr[2][4] ), .QN(n1191) );
  FD1 \gpr_reg[2][3]  ( .D(n1079), .CP(clk), .Q(\gpr[2][3] ), .QN(n1190) );
  FD1 \gpr_reg[2][2]  ( .D(n1078), .CP(clk), .Q(\gpr[2][2] ), .QN(n140) );
  FD1 \gpr_reg[2][1]  ( .D(n1077), .CP(clk), .Q(\gpr[2][1] ), .QN(n1140) );
  FD1 \gpr_reg[2][0]  ( .D(n1076), .CP(clk), .Q(\gpr[2][0] ), .QN(n147) );
  FD1 \gpr_reg[3][31]  ( .D(n1075), .CP(clk), .Q(\gpr[3][31] ), .QN(n1247) );
  FD1 \gpr_reg[3][30]  ( .D(n1074), .CP(clk), .Q(\gpr[3][30] ), .QN(n1246) );
  FD1 \gpr_reg[3][29]  ( .D(n1073), .CP(clk), .Q(\gpr[3][29] ), .QN(n1245) );
  FD1 \gpr_reg[3][28]  ( .D(n1072), .CP(clk), .Q(\gpr[3][28] ), .QN(n1244) );
  FD1 \gpr_reg[3][27]  ( .D(n1071), .CP(clk), .Q(\gpr[3][27] ), .QN(n1243) );
  FD1 \gpr_reg[3][26]  ( .D(n1070), .CP(clk), .Q(\gpr[3][26] ), .QN(n1242) );
  FD1 \gpr_reg[3][25]  ( .D(n1069), .CP(clk), .Q(\gpr[3][25] ), .QN(n1241) );
  FD1 \gpr_reg[3][24]  ( .D(n1068), .CP(clk), .Q(\gpr[3][24] ), .QN(n1240) );
  FD1 \gpr_reg[3][23]  ( .D(n1067), .CP(clk), .Q(\gpr[3][23] ), .QN(n1239) );
  FD1 \gpr_reg[3][22]  ( .D(n1066), .CP(clk), .Q(\gpr[3][22] ), .QN(n1238) );
  FD1 \gpr_reg[3][21]  ( .D(n1065), .CP(clk), .Q(\gpr[3][21] ), .QN(n1237) );
  FD1 \gpr_reg[3][20]  ( .D(n1064), .CP(clk), .Q(\gpr[3][20] ), .QN(n1236) );
  FD1 \gpr_reg[3][19]  ( .D(n1063), .CP(clk), .Q(\gpr[3][19] ), .QN(n1235) );
  FD1 \gpr_reg[3][18]  ( .D(n1062), .CP(clk), .Q(\gpr[3][18] ), .QN(n1234) );
  FD1 \gpr_reg[3][17]  ( .D(n1061), .CP(clk), .Q(\gpr[3][17] ), .QN(n1233) );
  FD1 \gpr_reg[3][16]  ( .D(n1060), .CP(clk), .Q(\gpr[3][16] ), .QN(n1232) );
  FD1 \gpr_reg[3][15]  ( .D(n1059), .CP(clk), .Q(\gpr[3][15] ), .QN(n1231) );
  FD1 \gpr_reg[3][14]  ( .D(n1058), .CP(clk), .Q(\gpr[3][14] ), .QN(n1230) );
  FD1 \gpr_reg[3][13]  ( .D(n1057), .CP(clk), .Q(\gpr[3][13] ), .QN(n1229) );
  FD1 \gpr_reg[3][12]  ( .D(n1056), .CP(clk), .Q(\gpr[3][12] ), .QN(n1228) );
  FD1 \gpr_reg[3][11]  ( .D(n1055), .CP(clk), .Q(\gpr[3][11] ), .QN(n1227) );
  FD1 \gpr_reg[3][10]  ( .D(n1054), .CP(clk), .Q(\gpr[3][10] ), .QN(n1226) );
  FD1 \gpr_reg[3][9]  ( .D(n1053), .CP(clk), .Q(\gpr[3][9] ), .QN(n1225) );
  FD1 \gpr_reg[3][8]  ( .D(n1052), .CP(clk), .Q(\gpr[3][8] ), .QN(n1224) );
  FD1 \gpr_reg[3][7]  ( .D(n1051), .CP(clk), .Q(\gpr[3][7] ), .QN(n1223) );
  FD1 \gpr_reg[3][6]  ( .D(n1050), .CP(clk), .Q(\gpr[3][6] ), .QN(n1222) );
  FD1 \gpr_reg[3][5]  ( .D(n1049), .CP(clk), .Q(\gpr[3][5] ), .QN(n1221) );
  FD1 \gpr_reg[3][4]  ( .D(n1048), .CP(clk), .Q(\gpr[3][4] ), .QN(n1220) );
  FD1 \gpr_reg[3][3]  ( .D(n1047), .CP(clk), .Q(\gpr[3][3] ), .QN(n1219) );
  FD1 \gpr_reg[3][2]  ( .D(n1046), .CP(clk), .Q(\gpr[3][2] ), .QN(n71) );
  FD1 \gpr_reg[3][1]  ( .D(n1045), .CP(clk), .Q(\gpr[3][1] ), .QN(n82) );
  FD1 \gpr_reg[3][0]  ( .D(n1044), .CP(clk), .Q(\gpr[3][0] ), .QN(n81) );
  FD1 \gpr_reg[4][31]  ( .D(n1043), .CP(clk), .Q(\gpr[4][31] ), .QN(n1176) );
  FD1 \gpr_reg[4][30]  ( .D(n1042), .CP(clk), .Q(\gpr[4][30] ), .QN(n1175) );
  FD1 \gpr_reg[4][29]  ( .D(n1041), .CP(clk), .Q(\gpr[4][29] ), .QN(n1174) );
  FD1 \gpr_reg[4][28]  ( .D(n1040), .CP(clk), .Q(\gpr[4][28] ), .QN(n1173) );
  FD1 \gpr_reg[4][27]  ( .D(n1039), .CP(clk), .Q(\gpr[4][27] ), .QN(n1172) );
  FD1 \gpr_reg[4][26]  ( .D(n1038), .CP(clk), .Q(\gpr[4][26] ), .QN(n1152) );
  FD1 \gpr_reg[4][25]  ( .D(n1037), .CP(clk), .Q(\gpr[4][25] ), .QN(n1171) );
  FD1 \gpr_reg[4][24]  ( .D(n1036), .CP(clk), .Q(\gpr[4][24] ), .QN(n1170) );
  FD1 \gpr_reg[4][23]  ( .D(n1035), .CP(clk), .Q(\gpr[4][23] ), .QN(n1151) );
  FD1 \gpr_reg[4][22]  ( .D(n1034), .CP(clk), .Q(\gpr[4][22] ), .QN(n1169) );
  FD1 \gpr_reg[4][21]  ( .D(n1033), .CP(clk), .Q(\gpr[4][21] ), .QN(n1150) );
  FD1 \gpr_reg[4][20]  ( .D(n1032), .CP(clk), .Q(\gpr[4][20] ), .QN(n1168) );
  FD1 \gpr_reg[4][19]  ( .D(n1031), .CP(clk), .Q(\gpr[4][19] ), .QN(n1149) );
  FD1 \gpr_reg[4][18]  ( .D(n1030), .CP(clk), .Q(\gpr[4][18] ), .QN(n1167) );
  FD1 \gpr_reg[4][17]  ( .D(n1029), .CP(clk), .Q(\gpr[4][17] ), .QN(n1166) );
  FD1 \gpr_reg[4][16]  ( .D(n1028), .CP(clk), .Q(\gpr[4][16] ), .QN(n1148) );
  FD1 \gpr_reg[4][15]  ( .D(n1027), .CP(clk), .Q(\gpr[4][15] ), .QN(n1147) );
  FD1 \gpr_reg[4][14]  ( .D(n1026), .CP(clk), .Q(\gpr[4][14] ), .QN(n1146) );
  FD1 \gpr_reg[4][13]  ( .D(n1025), .CP(clk), .Q(\gpr[4][13] ), .QN(n1145) );
  FD1 \gpr_reg[4][12]  ( .D(n1024), .CP(clk), .Q(\gpr[4][12] ), .QN(n1165) );
  FD1 \gpr_reg[4][11]  ( .D(n1023), .CP(clk), .Q(\gpr[4][11] ), .QN(n1164) );
  FD1 \gpr_reg[4][10]  ( .D(n1022), .CP(clk), .Q(\gpr[4][10] ), .QN(n1144) );
  FD1 \gpr_reg[4][9]  ( .D(n1021), .CP(clk), .Q(\gpr[4][9] ), .QN(n1143) );
  FD1 \gpr_reg[4][8]  ( .D(n1020), .CP(clk), .Q(\gpr[4][8] ), .QN(n1142) );
  FD1 \gpr_reg[4][7]  ( .D(n1019), .CP(clk), .Q(\gpr[4][7] ), .QN(n1163) );
  FD1 \gpr_reg[4][6]  ( .D(n1018), .CP(clk), .Q(\gpr[4][6] ), .QN(n1162) );
  FD1 \gpr_reg[4][5]  ( .D(n1017), .CP(clk), .Q(\gpr[4][5] ), .QN(n1141) );
  FD1 \gpr_reg[4][4]  ( .D(n1016), .CP(clk), .Q(\gpr[4][4] ), .QN(n141) );
  FD1 \gpr_reg[4][3]  ( .D(n1015), .CP(clk), .Q(\gpr[4][3] ), .QN(n1161) );
  FD1 \gpr_reg[4][2]  ( .D(n1014), .CP(clk), .Q(\gpr[4][2] ), .QN(n60) );
  FD1 \gpr_reg[4][1]  ( .D(n1013), .CP(clk), .Q(\gpr[4][1] ), .QN(n78) );
  FD1 \gpr_reg[4][0]  ( .D(n1012), .CP(clk), .Q(\gpr[4][0] ), .QN(n77) );
  FD1 \gpr_reg[5][31]  ( .D(n1011), .CP(clk), .Q(\gpr[5][31] ), .QN(n113) );
  FD1 \gpr_reg[5][30]  ( .D(n1010), .CP(clk), .Q(\gpr[5][30] ), .QN(n112) );
  FD1 \gpr_reg[5][29]  ( .D(n1009), .CP(clk), .Q(\gpr[5][29] ), .QN(n111) );
  FD1 \gpr_reg[5][28]  ( .D(n1008), .CP(clk), .Q(\gpr[5][28] ), .QN(n110) );
  FD1 \gpr_reg[5][27]  ( .D(n1007), .CP(clk), .Q(\gpr[5][27] ), .QN(n109) );
  FD1 \gpr_reg[5][26]  ( .D(n1006), .CP(clk), .Q(\gpr[5][26] ), .QN(n91) );
  FD1 \gpr_reg[5][25]  ( .D(n1005), .CP(clk), .Q(\gpr[5][25] ), .QN(n108) );
  FD1 \gpr_reg[5][24]  ( .D(n1004), .CP(clk), .Q(\gpr[5][24] ), .QN(n107) );
  FD1 \gpr_reg[5][23]  ( .D(n1003), .CP(clk), .Q(\gpr[5][23] ), .QN(n90) );
  FD1 \gpr_reg[5][22]  ( .D(n1002), .CP(clk), .Q(\gpr[5][22] ), .QN(n106) );
  FD1 \gpr_reg[5][21]  ( .D(n1001), .CP(clk), .Q(\gpr[5][21] ), .QN(n89) );
  FD1 \gpr_reg[5][20]  ( .D(n1000), .CP(clk), .Q(\gpr[5][20] ), .QN(n105) );
  FD1 \gpr_reg[5][19]  ( .D(n999), .CP(clk), .Q(\gpr[5][19] ), .QN(n88) );
  FD1 \gpr_reg[5][18]  ( .D(n998), .CP(clk), .Q(\gpr[5][18] ), .QN(n104) );
  FD1 \gpr_reg[5][17]  ( .D(n997), .CP(clk), .Q(\gpr[5][17] ), .QN(n103) );
  FD1 \gpr_reg[5][16]  ( .D(n996), .CP(clk), .Q(\gpr[5][16] ), .QN(n87) );
  FD1 \gpr_reg[5][15]  ( .D(n995), .CP(clk), .Q(\gpr[5][15] ), .QN(n102) );
  FD1 \gpr_reg[5][14]  ( .D(n994), .CP(clk), .Q(\gpr[5][14] ), .QN(n86) );
  FD1 \gpr_reg[5][13]  ( .D(n993), .CP(clk), .Q(\gpr[5][13] ), .QN(n85) );
  FD1 \gpr_reg[5][12]  ( .D(n992), .CP(clk), .Q(\gpr[5][12] ), .QN(n101) );
  FD1 \gpr_reg[5][11]  ( .D(n991), .CP(clk), .Q(\gpr[5][11] ), .QN(n100) );
  FD1 \gpr_reg[5][10]  ( .D(n990), .CP(clk), .Q(\gpr[5][10] ), .QN(n99) );
  FD1 \gpr_reg[5][9]  ( .D(n989), .CP(clk), .Q(\gpr[5][9] ), .QN(n84) );
  FD1 \gpr_reg[5][8]  ( .D(n988), .CP(clk), .Q(\gpr[5][8] ), .QN(n98) );
  FD1 \gpr_reg[5][7]  ( .D(n987), .CP(clk), .Q(\gpr[5][7] ), .QN(n97) );
  FD1 \gpr_reg[5][6]  ( .D(n986), .CP(clk), .Q(\gpr[5][6] ), .QN(n96) );
  FD1 \gpr_reg[5][5]  ( .D(n985), .CP(clk), .Q(\gpr[5][5] ), .QN(n83) );
  FD1 \gpr_reg[5][4]  ( .D(n984), .CP(clk), .Q(\gpr[5][4] ), .QN(n72) );
  FD1 \gpr_reg[5][3]  ( .D(n983), .CP(clk), .Q(\gpr[5][3] ), .QN(n95) );
  FD1 \gpr_reg[5][2]  ( .D(n982), .CP(clk), .Q(\gpr[5][2] ), .QN(n129) );
  FD1 \gpr_reg[5][1]  ( .D(n981), .CP(clk), .Q(\gpr[5][1] ), .QN(n144) );
  FD1 \gpr_reg[5][0]  ( .D(n980), .CP(clk), .Q(\gpr[5][0] ), .QN(n143) );
  FD1 \gpr_reg[6][31]  ( .D(n979), .CP(clk), .Q(\gpr[6][31] ), .QN(n1278) );
  FD1 \gpr_reg[6][30]  ( .D(n978), .CP(clk), .Q(\gpr[6][30] ), .QN(n1277) );
  FD1 \gpr_reg[6][29]  ( .D(n977), .CP(clk), .Q(\gpr[6][29] ), .QN(n1276) );
  FD1 \gpr_reg[6][28]  ( .D(n976), .CP(clk), .Q(\gpr[6][28] ), .QN(n1275) );
  FD1 \gpr_reg[6][27]  ( .D(n975), .CP(clk), .Q(\gpr[6][27] ), .QN(n1274) );
  FD1 \gpr_reg[6][26]  ( .D(n974), .CP(clk), .Q(\gpr[6][26] ), .QN(n1273) );
  FD1 \gpr_reg[6][25]  ( .D(n973), .CP(clk), .Q(\gpr[6][25] ), .QN(n1272) );
  FD1 \gpr_reg[6][24]  ( .D(n972), .CP(clk), .Q(\gpr[6][24] ), .QN(n1271) );
  FD1 \gpr_reg[6][23]  ( .D(n971), .CP(clk), .Q(\gpr[6][23] ), .QN(n1270) );
  FD1 \gpr_reg[6][22]  ( .D(n970), .CP(clk), .Q(\gpr[6][22] ), .QN(n1269) );
  FD1 \gpr_reg[6][21]  ( .D(n969), .CP(clk), .Q(\gpr[6][21] ), .QN(n1268) );
  FD1 \gpr_reg[6][20]  ( .D(n968), .CP(clk), .Q(\gpr[6][20] ), .QN(n1267) );
  FD1 \gpr_reg[6][19]  ( .D(n967), .CP(clk), .Q(\gpr[6][19] ), .QN(n1266) );
  FD1 \gpr_reg[6][18]  ( .D(n966), .CP(clk), .Q(\gpr[6][18] ), .QN(n1265) );
  FD1 \gpr_reg[6][17]  ( .D(n965), .CP(clk), .Q(\gpr[6][17] ), .QN(n1264) );
  FD1 \gpr_reg[6][16]  ( .D(n964), .CP(clk), .Q(\gpr[6][16] ), .QN(n1263) );
  FD1 \gpr_reg[6][15]  ( .D(n963), .CP(clk), .Q(\gpr[6][15] ), .QN(n1262) );
  FD1 \gpr_reg[6][14]  ( .D(n962), .CP(clk), .Q(\gpr[6][14] ), .QN(n1261) );
  FD1 \gpr_reg[6][13]  ( .D(n961), .CP(clk), .Q(\gpr[6][13] ), .QN(n1260) );
  FD1 \gpr_reg[6][12]  ( .D(n960), .CP(clk), .Q(\gpr[6][12] ), .QN(n1259) );
  FD1 \gpr_reg[6][11]  ( .D(n959), .CP(clk), .Q(\gpr[6][11] ), .QN(n1258) );
  FD1 \gpr_reg[6][10]  ( .D(n958), .CP(clk), .Q(\gpr[6][10] ), .QN(n1257) );
  FD1 \gpr_reg[6][9]  ( .D(n957), .CP(clk), .Q(\gpr[6][9] ), .QN(n1256) );
  FD1 \gpr_reg[6][8]  ( .D(n956), .CP(clk), .Q(\gpr[6][8] ), .QN(n1255) );
  FD1 \gpr_reg[6][7]  ( .D(n955), .CP(clk), .Q(\gpr[6][7] ), .QN(n1178) );
  FD1 \gpr_reg[6][6]  ( .D(n954), .CP(clk), .Q(\gpr[6][6] ), .QN(n1254) );
  FD1 \gpr_reg[6][5]  ( .D(n953), .CP(clk), .Q(\gpr[6][5] ), .QN(n1253) );
  FD1 \gpr_reg[6][4]  ( .D(n952), .CP(clk), .Q(\gpr[6][4] ), .QN(n1252) );
  FD1 \gpr_reg[6][3]  ( .D(n951), .CP(clk), .Q(\gpr[6][3] ), .QN(n1251) );
  FD1 \gpr_reg[6][2]  ( .D(n950), .CP(clk), .Q(\gpr[6][2] ), .QN(n1250) );
  FD1 \gpr_reg[6][1]  ( .D(n949), .CP(clk), .Q(\gpr[6][1] ), .QN(n1249) );
  FD1 \gpr_reg[6][0]  ( .D(n948), .CP(clk), .Q(\gpr[6][0] ), .QN(n1248) );
  FD1 \gpr_reg[7][31]  ( .D(n947), .CP(clk), .Q(\gpr[7][31] ), .QN(n1309) );
  FD1 \gpr_reg[7][30]  ( .D(n946), .CP(clk), .Q(\gpr[7][30] ), .QN(n1308) );
  FD1 \gpr_reg[7][29]  ( .D(n945), .CP(clk), .Q(\gpr[7][29] ), .QN(n1307) );
  FD1 \gpr_reg[7][28]  ( .D(n944), .CP(clk), .Q(\gpr[7][28] ), .QN(n1306) );
  FD1 \gpr_reg[7][27]  ( .D(n943), .CP(clk), .Q(\gpr[7][27] ), .QN(n1305) );
  FD1 \gpr_reg[7][26]  ( .D(n942), .CP(clk), .Q(\gpr[7][26] ), .QN(n1304) );
  FD1 \gpr_reg[7][25]  ( .D(n941), .CP(clk), .Q(\gpr[7][25] ), .QN(n1303) );
  FD1 \gpr_reg[7][24]  ( .D(n940), .CP(clk), .Q(\gpr[7][24] ), .QN(n1302) );
  FD1 \gpr_reg[7][23]  ( .D(n939), .CP(clk), .Q(\gpr[7][23] ), .QN(n1301) );
  FD1 \gpr_reg[7][22]  ( .D(n938), .CP(clk), .Q(\gpr[7][22] ), .QN(n1300) );
  FD1 \gpr_reg[7][21]  ( .D(n937), .CP(clk), .Q(\gpr[7][21] ), .QN(n1299) );
  FD1 \gpr_reg[7][20]  ( .D(n936), .CP(clk), .Q(\gpr[7][20] ), .QN(n1298) );
  FD1 \gpr_reg[7][19]  ( .D(n935), .CP(clk), .Q(\gpr[7][19] ), .QN(n1297) );
  FD1 \gpr_reg[7][18]  ( .D(n934), .CP(clk), .Q(\gpr[7][18] ), .QN(n1296) );
  FD1 \gpr_reg[7][17]  ( .D(n933), .CP(clk), .Q(\gpr[7][17] ), .QN(n1295) );
  FD1 \gpr_reg[7][16]  ( .D(n932), .CP(clk), .Q(\gpr[7][16] ), .QN(n1294) );
  FD1 \gpr_reg[7][15]  ( .D(n931), .CP(clk), .Q(\gpr[7][15] ), .QN(n1293) );
  FD1 \gpr_reg[7][14]  ( .D(n930), .CP(clk), .Q(\gpr[7][14] ), .QN(n1292) );
  FD1 \gpr_reg[7][13]  ( .D(n929), .CP(clk), .Q(\gpr[7][13] ), .QN(n1291) );
  FD1 \gpr_reg[7][12]  ( .D(n928), .CP(clk), .Q(\gpr[7][12] ), .QN(n1290) );
  FD1 \gpr_reg[7][11]  ( .D(n927), .CP(clk), .Q(\gpr[7][11] ), .QN(n1289) );
  FD1 \gpr_reg[7][10]  ( .D(n926), .CP(clk), .Q(\gpr[7][10] ), .QN(n1288) );
  FD1 \gpr_reg[7][9]  ( .D(n925), .CP(clk), .Q(\gpr[7][9] ), .QN(n1287) );
  FD1 \gpr_reg[7][8]  ( .D(n924), .CP(clk), .Q(\gpr[7][8] ), .QN(n1286) );
  FD1 \gpr_reg[7][7]  ( .D(n923), .CP(clk), .Q(\gpr[7][7] ), .QN(n114) );
  FD1 \gpr_reg[7][6]  ( .D(n922), .CP(clk), .Q(\gpr[7][6] ), .QN(n1285) );
  FD1 \gpr_reg[7][5]  ( .D(n921), .CP(clk), .Q(\gpr[7][5] ), .QN(n1284) );
  FD1 \gpr_reg[7][4]  ( .D(n920), .CP(clk), .Q(\gpr[7][4] ), .QN(n1283) );
  FD1 \gpr_reg[7][3]  ( .D(n919), .CP(clk), .Q(\gpr[7][3] ), .QN(n1282) );
  FD1 \gpr_reg[7][2]  ( .D(n918), .CP(clk), .Q(\gpr[7][2] ), .QN(n1281) );
  FD1 \gpr_reg[7][1]  ( .D(n917), .CP(clk), .Q(\gpr[7][1] ), .QN(n1280) );
  FD1 \gpr_reg[7][0]  ( .D(n916), .CP(clk), .Q(\gpr[7][0] ), .QN(n1279) );
  FD1 \gpr_reg[8][31]  ( .D(n915), .CP(clk), .Q(\gpr[8][31] ), .QN(n1337) );
  FD1 \gpr_reg[8][30]  ( .D(n914), .CP(clk), .Q(\gpr[8][30] ), .QN(n1336) );
  FD1 \gpr_reg[8][29]  ( .D(n913), .CP(clk), .Q(\gpr[8][29] ), .QN(n1335) );
  FD1 \gpr_reg[8][28]  ( .D(n912), .CP(clk), .Q(\gpr[8][28] ), .QN(n1334) );
  FD1 \gpr_reg[8][27]  ( .D(n911), .CP(clk), .Q(\gpr[8][27] ), .QN(n1333) );
  FD1 \gpr_reg[8][26]  ( .D(n910), .CP(clk), .Q(\gpr[8][26] ), .QN(n1332) );
  FD1 \gpr_reg[8][25]  ( .D(n909), .CP(clk), .Q(\gpr[8][25] ), .QN(n1331) );
  FD1 \gpr_reg[8][24]  ( .D(n908), .CP(clk), .Q(\gpr[8][24] ), .QN(n1330) );
  FD1 \gpr_reg[8][23]  ( .D(n907), .CP(clk), .Q(\gpr[8][23] ), .QN(n1329) );
  FD1 \gpr_reg[8][22]  ( .D(n906), .CP(clk), .Q(\gpr[8][22] ), .QN(n1328) );
  FD1 \gpr_reg[8][21]  ( .D(n905), .CP(clk), .Q(\gpr[8][21] ), .QN(n1327) );
  FD1 \gpr_reg[8][20]  ( .D(n904), .CP(clk), .Q(\gpr[8][20] ), .QN(n1326) );
  FD1 \gpr_reg[8][19]  ( .D(n903), .CP(clk), .Q(\gpr[8][19] ), .QN(n1325) );
  FD1 \gpr_reg[8][18]  ( .D(n902), .CP(clk), .Q(\gpr[8][18] ), .QN(n1324) );
  FD1 \gpr_reg[8][17]  ( .D(n901), .CP(clk), .Q(\gpr[8][17] ), .QN(n1323) );
  FD1 \gpr_reg[8][16]  ( .D(n900), .CP(clk), .Q(\gpr[8][16] ), .QN(n1322) );
  FD1 \gpr_reg[8][15]  ( .D(n899), .CP(clk), .Q(\gpr[8][15] ), .QN(n1321) );
  FD1 \gpr_reg[8][14]  ( .D(n898), .CP(clk), .Q(\gpr[8][14] ), .QN(n1320) );
  FD1 \gpr_reg[8][13]  ( .D(n897), .CP(clk), .Q(\gpr[8][13] ), .QN(n1319) );
  FD1 \gpr_reg[8][12]  ( .D(n896), .CP(clk), .Q(\gpr[8][12] ), .QN(n1318) );
  FD1 \gpr_reg[8][11]  ( .D(n895), .CP(clk), .Q(\gpr[8][11] ), .QN(n1317) );
  FD1 \gpr_reg[8][10]  ( .D(n894), .CP(clk), .Q(\gpr[8][10] ), .QN(n1316) );
  FD1 \gpr_reg[8][9]  ( .D(n893), .CP(clk), .Q(\gpr[8][9] ), .QN(n1315) );
  FD1 \gpr_reg[8][8]  ( .D(n892), .CP(clk), .Q(\gpr[8][8] ), .QN(n1314) );
  FD1 \gpr_reg[8][7]  ( .D(n891), .CP(clk), .Q(\gpr[8][7] ), .QN(n1313) );
  FD1 \gpr_reg[8][5]  ( .D(n889), .CP(clk), .Q(\gpr[8][5] ), .QN(n1312) );
  FD1 \gpr_reg[8][4]  ( .D(n888), .CP(clk), .Q(\gpr[8][4] ), .QN(n1311) );
  FD1 \gpr_reg[8][3]  ( .D(n887), .CP(clk), .Q(\gpr[8][3] ), .QN(n1310) );
  FD1 \gpr_reg[8][2]  ( .D(n886), .CP(clk), .Q(\gpr[8][2] ), .QN(n61) );
  FD1 \gpr_reg[8][1]  ( .D(n885), .CP(clk), .Q(\gpr[8][1] ), .QN(n80) );
  FD1 \gpr_reg[8][0]  ( .D(n884), .CP(clk), .Q(\gpr[8][0] ), .QN(n79) );
  FD1 \gpr_reg[9][31]  ( .D(n883), .CP(clk), .Q(\gpr[9][31] ), .QN(n1362) );
  FD1 \gpr_reg[9][30]  ( .D(n882), .CP(clk), .Q(\gpr[9][30] ), .QN(n1361) );
  FD1 \gpr_reg[9][29]  ( .D(n881), .CP(clk), .Q(\gpr[9][29] ), .QN(n1360) );
  FD1 \gpr_reg[9][28]  ( .D(n880), .CP(clk), .Q(\gpr[9][28] ), .QN(n1359) );
  FD1 \gpr_reg[9][27]  ( .D(n879), .CP(clk), .Q(\gpr[9][27] ), .QN(n1358) );
  FD1 \gpr_reg[9][26]  ( .D(n878), .CP(clk), .Q(\gpr[9][26] ), .QN(n1357) );
  FD1 \gpr_reg[9][25]  ( .D(n877), .CP(clk), .Q(\gpr[9][25] ), .QN(n1356) );
  FD1 \gpr_reg[9][24]  ( .D(n876), .CP(clk), .Q(\gpr[9][24] ), .QN(n1355) );
  FD1 \gpr_reg[9][23]  ( .D(n875), .CP(clk), .Q(\gpr[9][23] ), .QN(n1354) );
  FD1 \gpr_reg[9][22]  ( .D(n874), .CP(clk), .Q(\gpr[9][22] ), .QN(n1353) );
  FD1 \gpr_reg[9][21]  ( .D(n873), .CP(clk), .Q(\gpr[9][21] ), .QN(n1352) );
  FD1 \gpr_reg[9][20]  ( .D(n872), .CP(clk), .Q(\gpr[9][20] ), .QN(n1351) );
  FD1 \gpr_reg[9][19]  ( .D(n871), .CP(clk), .Q(\gpr[9][19] ), .QN(n1350) );
  FD1 \gpr_reg[9][18]  ( .D(n870), .CP(clk), .Q(\gpr[9][18] ), .QN(n1349) );
  FD1 \gpr_reg[9][17]  ( .D(n869), .CP(clk), .Q(\gpr[9][17] ), .QN(n1348) );
  FD1 \gpr_reg[9][16]  ( .D(n868), .CP(clk), .Q(\gpr[9][16] ), .QN(n1347) );
  FD1 \gpr_reg[9][15]  ( .D(n867), .CP(clk), .Q(\gpr[9][15] ), .QN(n1346) );
  FD1 \gpr_reg[9][14]  ( .D(n866), .CP(clk), .Q(\gpr[9][14] ), .QN(n1345) );
  FD1 \gpr_reg[9][13]  ( .D(n865), .CP(clk), .Q(\gpr[9][13] ), .QN(n1344) );
  FD1 \gpr_reg[9][12]  ( .D(n864), .CP(clk), .Q(\gpr[9][12] ), .QN(n1343) );
  FD1 \gpr_reg[9][11]  ( .D(n863), .CP(clk), .Q(\gpr[9][11] ), .QN(n1342) );
  FD1 \gpr_reg[9][10]  ( .D(n862), .CP(clk), .Q(\gpr[9][10] ), .QN(n1341) );
  FD1 \gpr_reg[9][8]  ( .D(n860), .CP(clk), .Q(\gpr[9][8] ), .QN(n1340) );
  FD1 \gpr_reg[9][7]  ( .D(n859), .CP(clk), .Q(\gpr[9][7] ), .QN(n1339) );
  FD1 \gpr_reg[9][3]  ( .D(n855), .CP(clk), .Q(\gpr[9][3] ), .QN(n1338) );
  FD1 \gpr_reg[9][2]  ( .D(n854), .CP(clk), .Q(\gpr[9][2] ), .QN(n130) );
  FD1 \gpr_reg[9][1]  ( .D(n853), .CP(clk), .Q(\gpr[9][1] ), .QN(n146) );
  FD1 \gpr_reg[9][0]  ( .D(n852), .CP(clk), .Q(\gpr[9][0] ), .QN(n145) );
  FD1 \gpr_reg[10][31]  ( .D(n851), .CP(clk), .Q(\gpr[10][31] ), .QN(n1393) );
  FD1 \gpr_reg[10][30]  ( .D(n850), .CP(clk), .Q(\gpr[10][30] ), .QN(n1392) );
  FD1 \gpr_reg[10][29]  ( .D(n849), .CP(clk), .Q(\gpr[10][29] ), .QN(n1391) );
  FD1 \gpr_reg[10][28]  ( .D(n848), .CP(clk), .Q(\gpr[10][28] ), .QN(n1390) );
  FD1 \gpr_reg[10][27]  ( .D(n847), .CP(clk), .Q(\gpr[10][27] ), .QN(n1389) );
  FD1 \gpr_reg[10][26]  ( .D(n846), .CP(clk), .Q(\gpr[10][26] ), .QN(n1388) );
  FD1 \gpr_reg[10][25]  ( .D(n845), .CP(clk), .Q(\gpr[10][25] ), .QN(n1387) );
  FD1 \gpr_reg[10][24]  ( .D(n844), .CP(clk), .Q(\gpr[10][24] ), .QN(n1386) );
  FD1 \gpr_reg[10][23]  ( .D(n843), .CP(clk), .Q(\gpr[10][23] ), .QN(n1385) );
  FD1 \gpr_reg[10][22]  ( .D(n842), .CP(clk), .Q(\gpr[10][22] ), .QN(n1384) );
  FD1 \gpr_reg[10][21]  ( .D(n841), .CP(clk), .Q(\gpr[10][21] ), .QN(n1383) );
  FD1 \gpr_reg[10][20]  ( .D(n840), .CP(clk), .Q(\gpr[10][20] ), .QN(n1382) );
  FD1 \gpr_reg[10][19]  ( .D(n839), .CP(clk), .Q(\gpr[10][19] ), .QN(n1381) );
  FD1 \gpr_reg[10][18]  ( .D(n838), .CP(clk), .Q(\gpr[10][18] ), .QN(n1380) );
  FD1 \gpr_reg[10][17]  ( .D(n837), .CP(clk), .Q(\gpr[10][17] ), .QN(n1379) );
  FD1 \gpr_reg[10][16]  ( .D(n836), .CP(clk), .Q(\gpr[10][16] ), .QN(n1378) );
  FD1 \gpr_reg[10][15]  ( .D(n835), .CP(clk), .Q(\gpr[10][15] ), .QN(n1377) );
  FD1 \gpr_reg[10][14]  ( .D(n834), .CP(clk), .Q(\gpr[10][14] ), .QN(n1376) );
  FD1 \gpr_reg[10][13]  ( .D(n833), .CP(clk), .Q(\gpr[10][13] ), .QN(n1375) );
  FD1 \gpr_reg[10][12]  ( .D(n832), .CP(clk), .Q(\gpr[10][12] ), .QN(n1374) );
  FD1 \gpr_reg[10][11]  ( .D(n831), .CP(clk), .Q(\gpr[10][11] ), .QN(n1373) );
  FD1 \gpr_reg[10][10]  ( .D(n830), .CP(clk), .Q(\gpr[10][10] ), .QN(n1372) );
  FD1 \gpr_reg[10][9]  ( .D(n829), .CP(clk), .Q(\gpr[10][9] ), .QN(n1371) );
  FD1 \gpr_reg[10][8]  ( .D(n828), .CP(clk), .Q(\gpr[10][8] ), .QN(n1370) );
  FD1 \gpr_reg[10][7]  ( .D(n827), .CP(clk), .Q(\gpr[10][7] ), .QN(n1369) );
  FD1 \gpr_reg[10][5]  ( .D(n825), .CP(clk), .Q(\gpr[10][5] ), .QN(n1368) );
  FD1 \gpr_reg[10][4]  ( .D(n824), .CP(clk), .Q(\gpr[10][4] ), .QN(n1367) );
  FD1 \gpr_reg[10][3]  ( .D(n823), .CP(clk), .Q(\gpr[10][3] ), .QN(n1366) );
  FD1 \gpr_reg[10][2]  ( .D(n822), .CP(clk), .Q(\gpr[10][2] ), .QN(n1365) );
  FD1 \gpr_reg[10][1]  ( .D(n821), .CP(clk), .Q(\gpr[10][1] ), .QN(n1364) );
  FD1 \gpr_reg[10][0]  ( .D(n820), .CP(clk), .Q(\gpr[10][0] ), .QN(n1363) );
  FD1 \gpr_reg[11][31]  ( .D(n819), .CP(clk), .Q(\gpr[11][31] ), .QN(n1424) );
  FD1 \gpr_reg[11][30]  ( .D(n818), .CP(clk), .Q(\gpr[11][30] ), .QN(n1423) );
  FD1 \gpr_reg[11][29]  ( .D(n817), .CP(clk), .Q(\gpr[11][29] ), .QN(n1422) );
  FD1 \gpr_reg[11][28]  ( .D(n816), .CP(clk), .Q(\gpr[11][28] ), .QN(n1421) );
  FD1 \gpr_reg[11][27]  ( .D(n815), .CP(clk), .Q(\gpr[11][27] ), .QN(n1420) );
  FD1 \gpr_reg[11][26]  ( .D(n814), .CP(clk), .Q(\gpr[11][26] ), .QN(n1419) );
  FD1 \gpr_reg[11][25]  ( .D(n813), .CP(clk), .Q(\gpr[11][25] ), .QN(n1418) );
  FD1 \gpr_reg[11][24]  ( .D(n812), .CP(clk), .Q(\gpr[11][24] ), .QN(n1417) );
  FD1 \gpr_reg[11][23]  ( .D(n811), .CP(clk), .Q(\gpr[11][23] ), .QN(n1416) );
  FD1 \gpr_reg[11][22]  ( .D(n810), .CP(clk), .Q(\gpr[11][22] ), .QN(n1415) );
  FD1 \gpr_reg[11][21]  ( .D(n809), .CP(clk), .Q(\gpr[11][21] ), .QN(n1414) );
  FD1 \gpr_reg[11][20]  ( .D(n808), .CP(clk), .Q(\gpr[11][20] ), .QN(n1413) );
  FD1 \gpr_reg[11][19]  ( .D(n807), .CP(clk), .Q(\gpr[11][19] ), .QN(n1412) );
  FD1 \gpr_reg[11][18]  ( .D(n806), .CP(clk), .Q(\gpr[11][18] ), .QN(n1411) );
  FD1 \gpr_reg[11][17]  ( .D(n805), .CP(clk), .Q(\gpr[11][17] ), .QN(n1410) );
  FD1 \gpr_reg[11][16]  ( .D(n804), .CP(clk), .Q(\gpr[11][16] ), .QN(n1409) );
  FD1 \gpr_reg[11][15]  ( .D(n803), .CP(clk), .Q(\gpr[11][15] ), .QN(n1408) );
  FD1 \gpr_reg[11][14]  ( .D(n802), .CP(clk), .Q(\gpr[11][14] ), .QN(n1407) );
  FD1 \gpr_reg[11][13]  ( .D(n801), .CP(clk), .Q(\gpr[11][13] ), .QN(n1406) );
  FD1 \gpr_reg[11][12]  ( .D(n800), .CP(clk), .Q(\gpr[11][12] ), .QN(n1405) );
  FD1 \gpr_reg[11][11]  ( .D(n799), .CP(clk), .Q(\gpr[11][11] ), .QN(n1404) );
  FD1 \gpr_reg[11][10]  ( .D(n798), .CP(clk), .Q(\gpr[11][10] ), .QN(n1403) );
  FD1 \gpr_reg[11][9]  ( .D(n797), .CP(clk), .Q(\gpr[11][9] ), .QN(n1402) );
  FD1 \gpr_reg[11][8]  ( .D(n796), .CP(clk), .Q(\gpr[11][8] ), .QN(n1401) );
  FD1 \gpr_reg[11][7]  ( .D(n795), .CP(clk), .Q(\gpr[11][7] ), .QN(n1400) );
  FD1 \gpr_reg[11][5]  ( .D(n793), .CP(clk), .Q(\gpr[11][5] ), .QN(n1399) );
  FD1 \gpr_reg[11][4]  ( .D(n792), .CP(clk), .Q(\gpr[11][4] ), .QN(n1398) );
  FD1 \gpr_reg[11][3]  ( .D(n791), .CP(clk), .Q(\gpr[11][3] ), .QN(n1397) );
  FD1 \gpr_reg[11][2]  ( .D(n790), .CP(clk), .Q(\gpr[11][2] ), .QN(n1396) );
  FD1 \gpr_reg[11][1]  ( .D(n789), .CP(clk), .Q(\gpr[11][1] ), .QN(n1395) );
  FD1 \gpr_reg[11][0]  ( .D(n788), .CP(clk), .Q(\gpr[11][0] ), .QN(n1394) );
  FD1 \gpr_reg[12][31]  ( .D(n787), .CP(clk), .Q(\gpr[12][31] ), .QN(n1455) );
  FD1 \gpr_reg[12][30]  ( .D(n786), .CP(clk), .Q(\gpr[12][30] ), .QN(n1454) );
  FD1 \gpr_reg[12][29]  ( .D(n785), .CP(clk), .Q(\gpr[12][29] ), .QN(n1453) );
  FD1 \gpr_reg[12][28]  ( .D(n784), .CP(clk), .Q(\gpr[12][28] ), .QN(n1452) );
  FD1 \gpr_reg[12][27]  ( .D(n783), .CP(clk), .Q(\gpr[12][27] ), .QN(n1451) );
  FD1 \gpr_reg[12][26]  ( .D(n782), .CP(clk), .Q(\gpr[12][26] ), .QN(n1450) );
  FD1 \gpr_reg[12][25]  ( .D(n781), .CP(clk), .Q(\gpr[12][25] ), .QN(n1449) );
  FD1 \gpr_reg[12][24]  ( .D(n780), .CP(clk), .Q(\gpr[12][24] ), .QN(n1448) );
  FD1 \gpr_reg[12][23]  ( .D(n779), .CP(clk), .Q(\gpr[12][23] ), .QN(n1447) );
  FD1 \gpr_reg[12][22]  ( .D(n778), .CP(clk), .Q(\gpr[12][22] ), .QN(n1446) );
  FD1 \gpr_reg[12][21]  ( .D(n777), .CP(clk), .Q(\gpr[12][21] ), .QN(n1445) );
  FD1 \gpr_reg[12][20]  ( .D(n776), .CP(clk), .Q(\gpr[12][20] ), .QN(n1444) );
  FD1 \gpr_reg[12][19]  ( .D(n775), .CP(clk), .Q(\gpr[12][19] ), .QN(n1443) );
  FD1 \gpr_reg[12][18]  ( .D(n774), .CP(clk), .Q(\gpr[12][18] ), .QN(n1442) );
  FD1 \gpr_reg[12][17]  ( .D(n773), .CP(clk), .Q(\gpr[12][17] ), .QN(n1441) );
  FD1 \gpr_reg[12][16]  ( .D(n772), .CP(clk), .Q(\gpr[12][16] ), .QN(n1440) );
  FD1 \gpr_reg[12][15]  ( .D(n771), .CP(clk), .Q(\gpr[12][15] ), .QN(n1439) );
  FD1 \gpr_reg[12][14]  ( .D(n770), .CP(clk), .Q(\gpr[12][14] ), .QN(n1438) );
  FD1 \gpr_reg[12][13]  ( .D(n769), .CP(clk), .Q(\gpr[12][13] ), .QN(n1437) );
  FD1 \gpr_reg[12][12]  ( .D(n768), .CP(clk), .Q(\gpr[12][12] ), .QN(n1436) );
  FD1 \gpr_reg[12][11]  ( .D(n767), .CP(clk), .Q(\gpr[12][11] ), .QN(n1435) );
  FD1 \gpr_reg[12][10]  ( .D(n766), .CP(clk), .Q(\gpr[12][10] ), .QN(n1434) );
  FD1 \gpr_reg[12][9]  ( .D(n765), .CP(clk), .Q(\gpr[12][9] ), .QN(n1433) );
  FD1 \gpr_reg[12][8]  ( .D(n764), .CP(clk), .Q(\gpr[12][8] ), .QN(n1432) );
  FD1 \gpr_reg[12][7]  ( .D(n763), .CP(clk), .Q(\gpr[12][7] ), .QN(n1431) );
  FD1 \gpr_reg[12][5]  ( .D(n761), .CP(clk), .Q(\gpr[12][5] ), .QN(n1430) );
  FD1 \gpr_reg[12][4]  ( .D(n760), .CP(clk), .Q(\gpr[12][4] ), .QN(n1429) );
  FD1 \gpr_reg[12][3]  ( .D(n759), .CP(clk), .Q(\gpr[12][3] ), .QN(n1428) );
  FD1 \gpr_reg[12][2]  ( .D(n758), .CP(clk), .Q(\gpr[12][2] ), .QN(n1427) );
  FD1 \gpr_reg[12][1]  ( .D(n757), .CP(clk), .Q(\gpr[12][1] ), .QN(n1426) );
  FD1 \gpr_reg[12][0]  ( .D(n756), .CP(clk), .Q(\gpr[12][0] ), .QN(n1425) );
  FD1 \gpr_reg[13][31]  ( .D(n755), .CP(clk), .Q(\gpr[13][31] ), .QN(n1486) );
  FD1 \gpr_reg[13][30]  ( .D(n754), .CP(clk), .Q(\gpr[13][30] ), .QN(n1485) );
  FD1 \gpr_reg[13][29]  ( .D(n753), .CP(clk), .Q(\gpr[13][29] ), .QN(n1484) );
  FD1 \gpr_reg[13][28]  ( .D(n752), .CP(clk), .Q(\gpr[13][28] ), .QN(n1483) );
  FD1 \gpr_reg[13][27]  ( .D(n751), .CP(clk), .Q(\gpr[13][27] ), .QN(n1482) );
  FD1 \gpr_reg[13][26]  ( .D(n750), .CP(clk), .Q(\gpr[13][26] ), .QN(n1481) );
  FD1 \gpr_reg[13][25]  ( .D(n749), .CP(clk), .Q(\gpr[13][25] ), .QN(n1480) );
  FD1 \gpr_reg[13][24]  ( .D(n748), .CP(clk), .Q(\gpr[13][24] ), .QN(n1479) );
  FD1 \gpr_reg[13][23]  ( .D(n747), .CP(clk), .Q(\gpr[13][23] ), .QN(n1478) );
  FD1 \gpr_reg[13][22]  ( .D(n746), .CP(clk), .Q(\gpr[13][22] ), .QN(n1477) );
  FD1 \gpr_reg[13][21]  ( .D(n745), .CP(clk), .Q(\gpr[13][21] ), .QN(n1476) );
  FD1 \gpr_reg[13][20]  ( .D(n744), .CP(clk), .Q(\gpr[13][20] ), .QN(n1475) );
  FD1 \gpr_reg[13][19]  ( .D(n743), .CP(clk), .Q(\gpr[13][19] ), .QN(n1474) );
  FD1 \gpr_reg[13][18]  ( .D(n742), .CP(clk), .Q(\gpr[13][18] ), .QN(n1473) );
  FD1 \gpr_reg[13][17]  ( .D(n741), .CP(clk), .Q(\gpr[13][17] ), .QN(n1472) );
  FD1 \gpr_reg[13][16]  ( .D(n740), .CP(clk), .Q(\gpr[13][16] ), .QN(n1471) );
  FD1 \gpr_reg[13][15]  ( .D(n739), .CP(clk), .Q(\gpr[13][15] ), .QN(n1470) );
  FD1 \gpr_reg[13][14]  ( .D(n738), .CP(clk), .Q(\gpr[13][14] ), .QN(n1469) );
  FD1 \gpr_reg[13][13]  ( .D(n737), .CP(clk), .Q(\gpr[13][13] ), .QN(n1468) );
  FD1 \gpr_reg[13][12]  ( .D(n736), .CP(clk), .Q(\gpr[13][12] ), .QN(n1467) );
  FD1 \gpr_reg[13][11]  ( .D(n735), .CP(clk), .Q(\gpr[13][11] ), .QN(n1466) );
  FD1 \gpr_reg[13][10]  ( .D(n734), .CP(clk), .Q(\gpr[13][10] ), .QN(n1465) );
  FD1 \gpr_reg[13][9]  ( .D(n733), .CP(clk), .Q(\gpr[13][9] ), .QN(n1464) );
  FD1 \gpr_reg[13][8]  ( .D(n732), .CP(clk), .Q(\gpr[13][8] ), .QN(n1463) );
  FD1 \gpr_reg[13][7]  ( .D(n731), .CP(clk), .Q(\gpr[13][7] ), .QN(n1462) );
  FD1 \gpr_reg[13][5]  ( .D(n729), .CP(clk), .Q(\gpr[13][5] ), .QN(n1461) );
  FD1 \gpr_reg[13][4]  ( .D(n728), .CP(clk), .Q(\gpr[13][4] ), .QN(n1460) );
  FD1 \gpr_reg[13][3]  ( .D(n727), .CP(clk), .Q(\gpr[13][3] ), .QN(n1459) );
  FD1 \gpr_reg[13][2]  ( .D(n726), .CP(clk), .Q(\gpr[13][2] ), .QN(n1458) );
  FD1 \gpr_reg[13][1]  ( .D(n725), .CP(clk), .Q(\gpr[13][1] ), .QN(n1457) );
  FD1 \gpr_reg[13][0]  ( .D(n724), .CP(clk), .Q(\gpr[13][0] ), .QN(n1456) );
  FD1 \gpr_reg[14][31]  ( .D(n723), .CP(clk), .Q(\gpr[14][31] ), .QN(n1514) );
  FD1 \gpr_reg[14][30]  ( .D(n722), .CP(clk), .Q(\gpr[14][30] ), .QN(n1513) );
  FD1 \gpr_reg[14][29]  ( .D(n721), .CP(clk), .Q(\gpr[14][29] ), .QN(n1512) );
  FD1 \gpr_reg[14][28]  ( .D(n720), .CP(clk), .Q(\gpr[14][28] ), .QN(n1511) );
  FD1 \gpr_reg[14][27]  ( .D(n719), .CP(clk), .Q(\gpr[14][27] ), .QN(n1510) );
  FD1 \gpr_reg[14][26]  ( .D(n718), .CP(clk), .Q(\gpr[14][26] ), .QN(n1509) );
  FD1 \gpr_reg[14][25]  ( .D(n717), .CP(clk), .Q(\gpr[14][25] ), .QN(n1508) );
  FD1 \gpr_reg[14][24]  ( .D(n716), .CP(clk), .Q(\gpr[14][24] ), .QN(n1507) );
  FD1 \gpr_reg[14][23]  ( .D(n715), .CP(clk), .Q(\gpr[14][23] ), .QN(n1506) );
  FD1 \gpr_reg[14][22]  ( .D(n714), .CP(clk), .Q(\gpr[14][22] ), .QN(n1505) );
  FD1 \gpr_reg[14][21]  ( .D(n713), .CP(clk), .Q(\gpr[14][21] ), .QN(n1504) );
  FD1 \gpr_reg[14][20]  ( .D(n712), .CP(clk), .Q(\gpr[14][20] ), .QN(n1503) );
  FD1 \gpr_reg[14][19]  ( .D(n711), .CP(clk), .Q(\gpr[14][19] ), .QN(n1502) );
  FD1 \gpr_reg[14][18]  ( .D(n710), .CP(clk), .Q(\gpr[14][18] ), .QN(n1501) );
  FD1 \gpr_reg[14][17]  ( .D(n709), .CP(clk), .Q(\gpr[14][17] ), .QN(n1500) );
  FD1 \gpr_reg[14][16]  ( .D(n708), .CP(clk), .Q(\gpr[14][16] ), .QN(n1499) );
  FD1 \gpr_reg[14][15]  ( .D(n707), .CP(clk), .Q(\gpr[14][15] ), .QN(n1498) );
  FD1 \gpr_reg[14][14]  ( .D(n706), .CP(clk), .Q(\gpr[14][14] ), .QN(n1497) );
  FD1 \gpr_reg[14][13]  ( .D(n705), .CP(clk), .Q(\gpr[14][13] ), .QN(n1496) );
  FD1 \gpr_reg[14][12]  ( .D(n704), .CP(clk), .Q(\gpr[14][12] ), .QN(n1495) );
  FD1 \gpr_reg[14][11]  ( .D(n703), .CP(clk), .Q(\gpr[14][11] ), .QN(n1494) );
  FD1 \gpr_reg[14][10]  ( .D(n702), .CP(clk), .Q(\gpr[14][10] ), .QN(n1493) );
  FD1 \gpr_reg[14][9]  ( .D(n701), .CP(clk), .Q(\gpr[14][9] ), .QN(n1492) );
  FD1 \gpr_reg[14][8]  ( .D(n700), .CP(clk), .Q(\gpr[14][8] ), .QN(n1491) );
  FD1 \gpr_reg[14][7]  ( .D(n699), .CP(clk), .Q(\gpr[14][7] ), .QN(n1490) );
  FD1 \gpr_reg[14][5]  ( .D(n697), .CP(clk), .Q(\gpr[14][5] ), .QN(n1489) );
  FD1 \gpr_reg[14][4]  ( .D(n696), .CP(clk), .Q(\gpr[14][4] ), .QN(n1488) );
  FD1 \gpr_reg[14][3]  ( .D(n695), .CP(clk), .Q(\gpr[14][3] ), .QN(n1487) );
  FD1 \gpr_reg[14][2]  ( .D(n694), .CP(clk), .Q(\gpr[14][2] ), .QN(n138) );
  FD1 \gpr_reg[14][1]  ( .D(n693), .CP(clk), .Q(\gpr[14][1] ), .QN(n135) );
  FD1 \gpr_reg[14][0]  ( .D(n692), .CP(clk), .Q(\gpr[14][0] ), .QN(n132) );
  FD1 \gpr_reg[15][31]  ( .D(n691), .CP(clk), .Q(\gpr[15][31] ), .QN(n1542) );
  FD1 \gpr_reg[15][30]  ( .D(n690), .CP(clk), .Q(\gpr[15][30] ), .QN(n1541) );
  FD1 \gpr_reg[15][29]  ( .D(n689), .CP(clk), .Q(\gpr[15][29] ), .QN(n1540) );
  FD1 \gpr_reg[15][28]  ( .D(n688), .CP(clk), .Q(\gpr[15][28] ), .QN(n1539) );
  FD1 \gpr_reg[15][27]  ( .D(n687), .CP(clk), .Q(\gpr[15][27] ), .QN(n1538) );
  FD1 \gpr_reg[15][26]  ( .D(n686), .CP(clk), .Q(\gpr[15][26] ), .QN(n1537) );
  FD1 \gpr_reg[15][25]  ( .D(n685), .CP(clk), .Q(\gpr[15][25] ), .QN(n1536) );
  FD1 \gpr_reg[15][24]  ( .D(n684), .CP(clk), .Q(\gpr[15][24] ), .QN(n1535) );
  FD1 \gpr_reg[15][23]  ( .D(n683), .CP(clk), .Q(\gpr[15][23] ), .QN(n1534) );
  FD1 \gpr_reg[15][22]  ( .D(n682), .CP(clk), .Q(\gpr[15][22] ), .QN(n1533) );
  FD1 \gpr_reg[15][21]  ( .D(n681), .CP(clk), .Q(\gpr[15][21] ), .QN(n1532) );
  FD1 \gpr_reg[15][20]  ( .D(n680), .CP(clk), .Q(\gpr[15][20] ), .QN(n1531) );
  FD1 \gpr_reg[15][19]  ( .D(n679), .CP(clk), .Q(\gpr[15][19] ), .QN(n1530) );
  FD1 \gpr_reg[15][18]  ( .D(n678), .CP(clk), .Q(\gpr[15][18] ), .QN(n1529) );
  FD1 \gpr_reg[15][17]  ( .D(n677), .CP(clk), .Q(\gpr[15][17] ), .QN(n1528) );
  FD1 \gpr_reg[15][16]  ( .D(n676), .CP(clk), .Q(\gpr[15][16] ), .QN(n1527) );
  FD1 \gpr_reg[15][15]  ( .D(n675), .CP(clk), .Q(\gpr[15][15] ), .QN(n1526) );
  FD1 \gpr_reg[15][14]  ( .D(n674), .CP(clk), .Q(\gpr[15][14] ), .QN(n1525) );
  FD1 \gpr_reg[15][13]  ( .D(n673), .CP(clk), .Q(\gpr[15][13] ), .QN(n1524) );
  FD1 \gpr_reg[15][12]  ( .D(n672), .CP(clk), .Q(\gpr[15][12] ), .QN(n1523) );
  FD1 \gpr_reg[15][11]  ( .D(n671), .CP(clk), .Q(\gpr[15][11] ), .QN(n1522) );
  FD1 \gpr_reg[15][10]  ( .D(n670), .CP(clk), .Q(\gpr[15][10] ), .QN(n1521) );
  FD1 \gpr_reg[15][9]  ( .D(n669), .CP(clk), .Q(\gpr[15][9] ), .QN(n1520) );
  FD1 \gpr_reg[15][8]  ( .D(n668), .CP(clk), .Q(\gpr[15][8] ), .QN(n1519) );
  FD1 \gpr_reg[15][7]  ( .D(n667), .CP(clk), .Q(\gpr[15][7] ), .QN(n1518) );
  FD1 \gpr_reg[15][5]  ( .D(n665), .CP(clk), .Q(\gpr[15][5] ), .QN(n1517) );
  FD1 \gpr_reg[15][4]  ( .D(n664), .CP(clk), .Q(\gpr[15][4] ), .QN(n1516) );
  FD1 \gpr_reg[15][3]  ( .D(n663), .CP(clk), .Q(\gpr[15][3] ), .QN(n1515) );
  FD1 \gpr_reg[15][2]  ( .D(n662), .CP(clk), .Q(\gpr[15][2] ), .QN(n69) );
  FD1 \gpr_reg[15][1]  ( .D(n661), .CP(clk), .Q(\gpr[15][1] ), .QN(n66) );
  FD1 \gpr_reg[15][0]  ( .D(n660), .CP(clk), .Q(\gpr[15][0] ), .QN(n63) );
  FD1 \gpr_reg[16][31]  ( .D(n659), .CP(clk), .Q(\gpr[16][31] ), .QN(n1574) );
  FD1 \gpr_reg[16][30]  ( .D(n658), .CP(clk), .Q(\gpr[16][30] ), .QN(n1573) );
  FD1 \gpr_reg[16][29]  ( .D(n657), .CP(clk), .Q(\gpr[16][29] ), .QN(n1572) );
  FD1 \gpr_reg[16][28]  ( .D(n656), .CP(clk), .Q(\gpr[16][28] ), .QN(n1571) );
  FD1 \gpr_reg[16][27]  ( .D(n655), .CP(clk), .Q(\gpr[16][27] ), .QN(n1570) );
  FD1 \gpr_reg[16][26]  ( .D(n654), .CP(clk), .Q(\gpr[16][26] ), .QN(n1569) );
  FD1 \gpr_reg[16][25]  ( .D(n653), .CP(clk), .Q(\gpr[16][25] ), .QN(n1568) );
  FD1 \gpr_reg[16][24]  ( .D(n652), .CP(clk), .Q(\gpr[16][24] ), .QN(n1567) );
  FD1 \gpr_reg[16][23]  ( .D(n651), .CP(clk), .Q(\gpr[16][23] ), .QN(n1566) );
  FD1 \gpr_reg[16][22]  ( .D(n650), .CP(clk), .Q(\gpr[16][22] ), .QN(n1565) );
  FD1 \gpr_reg[16][21]  ( .D(n649), .CP(clk), .Q(\gpr[16][21] ), .QN(n1564) );
  FD1 \gpr_reg[16][20]  ( .D(n648), .CP(clk), .Q(\gpr[16][20] ), .QN(n1563) );
  FD1 \gpr_reg[16][19]  ( .D(n647), .CP(clk), .Q(\gpr[16][19] ), .QN(n1562) );
  FD1 \gpr_reg[16][18]  ( .D(n646), .CP(clk), .Q(\gpr[16][18] ), .QN(n1561) );
  FD1 \gpr_reg[16][17]  ( .D(n645), .CP(clk), .Q(\gpr[16][17] ), .QN(n1560) );
  FD1 \gpr_reg[16][16]  ( .D(n644), .CP(clk), .Q(\gpr[16][16] ), .QN(n1559) );
  FD1 \gpr_reg[16][15]  ( .D(n643), .CP(clk), .Q(\gpr[16][15] ), .QN(n1558) );
  FD1 \gpr_reg[16][14]  ( .D(n642), .CP(clk), .Q(\gpr[16][14] ), .QN(n1557) );
  FD1 \gpr_reg[16][13]  ( .D(n641), .CP(clk), .Q(\gpr[16][13] ), .QN(n1556) );
  FD1 \gpr_reg[16][12]  ( .D(n640), .CP(clk), .Q(\gpr[16][12] ), .QN(n1555) );
  FD1 \gpr_reg[16][11]  ( .D(n639), .CP(clk), .Q(\gpr[16][11] ), .QN(n1554) );
  FD1 \gpr_reg[16][10]  ( .D(n638), .CP(clk), .Q(\gpr[16][10] ), .QN(n1553) );
  FD1 \gpr_reg[16][9]  ( .D(n637), .CP(clk), .Q(\gpr[16][9] ), .QN(n1552) );
  FD1 \gpr_reg[16][8]  ( .D(n636), .CP(clk), .Q(\gpr[16][8] ), .QN(n1551) );
  FD1 \gpr_reg[16][7]  ( .D(n635), .CP(clk), .Q(\gpr[16][7] ), .QN(n1550) );
  FD1 \gpr_reg[16][6]  ( .D(n634), .CP(clk), .Q(\gpr[16][6] ), .QN(n1549) );
  FD1 \gpr_reg[16][5]  ( .D(n633), .CP(clk), .Q(\gpr[16][5] ), .QN(n1548) );
  FD1 \gpr_reg[16][4]  ( .D(n632), .CP(clk), .Q(\gpr[16][4] ), .QN(n1547) );
  FD1 \gpr_reg[16][3]  ( .D(n631), .CP(clk), .Q(\gpr[16][3] ), .QN(n1546) );
  FD1 \gpr_reg[16][2]  ( .D(n630), .CP(clk), .Q(\gpr[16][2] ), .QN(n1545) );
  FD1 \gpr_reg[16][1]  ( .D(n629), .CP(clk), .Q(\gpr[16][1] ), .QN(n1544) );
  FD1 \gpr_reg[16][0]  ( .D(n628), .CP(clk), .Q(\gpr[16][0] ), .QN(n1543) );
  FD1 \gpr_reg[17][31]  ( .D(n627), .CP(clk), .Q(\gpr[17][31] ), .QN(n1605) );
  FD1 \gpr_reg[17][30]  ( .D(n626), .CP(clk), .Q(\gpr[17][30] ), .QN(n1604) );
  FD1 \gpr_reg[17][29]  ( .D(n625), .CP(clk), .Q(\gpr[17][29] ), .QN(n1603) );
  FD1 \gpr_reg[17][28]  ( .D(n624), .CP(clk), .Q(\gpr[17][28] ), .QN(n1602) );
  FD1 \gpr_reg[17][27]  ( .D(n623), .CP(clk), .Q(\gpr[17][27] ), .QN(n1601) );
  FD1 \gpr_reg[17][26]  ( .D(n622), .CP(clk), .Q(\gpr[17][26] ), .QN(n1600) );
  FD1 \gpr_reg[17][25]  ( .D(n621), .CP(clk), .Q(\gpr[17][25] ), .QN(n1599) );
  FD1 \gpr_reg[17][24]  ( .D(n620), .CP(clk), .Q(\gpr[17][24] ), .QN(n1598) );
  FD1 \gpr_reg[17][23]  ( .D(n619), .CP(clk), .Q(\gpr[17][23] ), .QN(n1597) );
  FD1 \gpr_reg[17][22]  ( .D(n618), .CP(clk), .Q(\gpr[17][22] ), .QN(n1596) );
  FD1 \gpr_reg[17][21]  ( .D(n617), .CP(clk), .Q(\gpr[17][21] ), .QN(n1595) );
  FD1 \gpr_reg[17][20]  ( .D(n616), .CP(clk), .Q(\gpr[17][20] ), .QN(n1594) );
  FD1 \gpr_reg[17][19]  ( .D(n615), .CP(clk), .Q(\gpr[17][19] ), .QN(n1593) );
  FD1 \gpr_reg[17][18]  ( .D(n614), .CP(clk), .Q(\gpr[17][18] ), .QN(n1592) );
  FD1 \gpr_reg[17][17]  ( .D(n613), .CP(clk), .Q(\gpr[17][17] ), .QN(n1591) );
  FD1 \gpr_reg[17][16]  ( .D(n612), .CP(clk), .Q(\gpr[17][16] ), .QN(n1590) );
  FD1 \gpr_reg[17][15]  ( .D(n611), .CP(clk), .Q(\gpr[17][15] ), .QN(n1589) );
  FD1 \gpr_reg[17][14]  ( .D(n610), .CP(clk), .Q(\gpr[17][14] ), .QN(n1588) );
  FD1 \gpr_reg[17][13]  ( .D(n609), .CP(clk), .Q(\gpr[17][13] ), .QN(n1587) );
  FD1 \gpr_reg[17][12]  ( .D(n608), .CP(clk), .Q(\gpr[17][12] ), .QN(n1586) );
  FD1 \gpr_reg[17][11]  ( .D(n607), .CP(clk), .Q(\gpr[17][11] ), .QN(n1585) );
  FD1 \gpr_reg[17][10]  ( .D(n606), .CP(clk), .Q(\gpr[17][10] ), .QN(n1584) );
  FD1 \gpr_reg[17][8]  ( .D(n604), .CP(clk), .Q(\gpr[17][8] ), .QN(n1583) );
  FD1 \gpr_reg[17][7]  ( .D(n603), .CP(clk), .Q(\gpr[17][7] ), .QN(n1582) );
  FD1 \gpr_reg[17][6]  ( .D(n602), .CP(clk), .Q(\gpr[17][6] ), .QN(n1581) );
  FD1 \gpr_reg[17][5]  ( .D(n601), .CP(clk), .Q(\gpr[17][5] ), .QN(n1580) );
  FD1 \gpr_reg[17][4]  ( .D(n600), .CP(clk), .Q(\gpr[17][4] ), .QN(n1579) );
  FD1 \gpr_reg[17][3]  ( .D(n599), .CP(clk), .Q(\gpr[17][3] ), .QN(n1578) );
  FD1 \gpr_reg[17][2]  ( .D(n598), .CP(clk), .Q(\gpr[17][2] ), .QN(n1577) );
  FD1 \gpr_reg[17][1]  ( .D(n597), .CP(clk), .Q(\gpr[17][1] ), .QN(n1576) );
  FD1 \gpr_reg[17][0]  ( .D(n596), .CP(clk), .Q(\gpr[17][0] ), .QN(n1575) );
  FD1 \gpr_reg[18][31]  ( .D(n595), .CP(clk), .Q(\gpr[18][31] ), .QN(n1634) );
  FD1 \gpr_reg[18][30]  ( .D(n594), .CP(clk), .Q(\gpr[18][30] ), .QN(n1633) );
  FD1 \gpr_reg[18][29]  ( .D(n593), .CP(clk), .Q(\gpr[18][29] ), .QN(n1632) );
  FD1 \gpr_reg[18][28]  ( .D(n592), .CP(clk), .Q(\gpr[18][28] ), .QN(n1631) );
  FD1 \gpr_reg[18][27]  ( .D(n591), .CP(clk), .Q(\gpr[18][27] ), .QN(n1630) );
  FD1 \gpr_reg[18][26]  ( .D(n590), .CP(clk), .Q(\gpr[18][26] ), .QN(n1629) );
  FD1 \gpr_reg[18][25]  ( .D(n589), .CP(clk), .Q(\gpr[18][25] ), .QN(n1628) );
  FD1 \gpr_reg[18][24]  ( .D(n588), .CP(clk), .Q(\gpr[18][24] ), .QN(n1627) );
  FD1 \gpr_reg[18][23]  ( .D(n587), .CP(clk), .Q(\gpr[18][23] ), .QN(n1626) );
  FD1 \gpr_reg[18][22]  ( .D(n586), .CP(clk), .Q(\gpr[18][22] ), .QN(n1625) );
  FD1 \gpr_reg[18][21]  ( .D(n585), .CP(clk), .Q(\gpr[18][21] ), .QN(n1624) );
  FD1 \gpr_reg[18][20]  ( .D(n584), .CP(clk), .Q(\gpr[18][20] ), .QN(n1623) );
  FD1 \gpr_reg[18][19]  ( .D(n583), .CP(clk), .Q(\gpr[18][19] ), .QN(n1622) );
  FD1 \gpr_reg[18][18]  ( .D(n582), .CP(clk), .Q(\gpr[18][18] ), .QN(n1621) );
  FD1 \gpr_reg[18][17]  ( .D(n581), .CP(clk), .Q(\gpr[18][17] ), .QN(n1620) );
  FD1 \gpr_reg[18][16]  ( .D(n580), .CP(clk), .Q(\gpr[18][16] ), .QN(n1619) );
  FD1 \gpr_reg[18][15]  ( .D(n579), .CP(clk), .Q(\gpr[18][15] ), .QN(n1618) );
  FD1 \gpr_reg[18][14]  ( .D(n578), .CP(clk), .Q(\gpr[18][14] ), .QN(n1617) );
  FD1 \gpr_reg[18][13]  ( .D(n577), .CP(clk), .Q(\gpr[18][13] ), .QN(n1616) );
  FD1 \gpr_reg[18][12]  ( .D(n576), .CP(clk), .Q(\gpr[18][12] ), .QN(n1615) );
  FD1 \gpr_reg[18][11]  ( .D(n575), .CP(clk), .Q(\gpr[18][11] ), .QN(n1614) );
  FD1 \gpr_reg[18][10]  ( .D(n574), .CP(clk), .Q(\gpr[18][10] ), .QN(n1613) );
  FD1 \gpr_reg[18][9]  ( .D(n573), .CP(clk), .Q(\gpr[18][9] ), .QN(n1612) );
  FD1 \gpr_reg[18][8]  ( .D(n572), .CP(clk), .Q(\gpr[18][8] ), .QN(n1611) );
  FD1 \gpr_reg[18][7]  ( .D(n571), .CP(clk), .Q(\gpr[18][7] ), .QN(n1610) );
  FD1 \gpr_reg[18][6]  ( .D(n570), .CP(clk), .Q(\gpr[18][6] ), .QN(n1609) );
  FD1 \gpr_reg[18][5]  ( .D(n569), .CP(clk), .Q(\gpr[18][5] ), .QN(n1608) );
  FD1 \gpr_reg[18][4]  ( .D(n568), .CP(clk), .Q(\gpr[18][4] ), .QN(n1607) );
  FD1 \gpr_reg[18][3]  ( .D(n567), .CP(clk), .Q(\gpr[18][3] ), .QN(n1606) );
  FD1 \gpr_reg[18][2]  ( .D(n566), .CP(clk), .Q(\gpr[18][2] ), .QN(n139) );
  FD1 \gpr_reg[18][1]  ( .D(n565), .CP(clk), .Q(\gpr[18][1] ), .QN(n136) );
  FD1 \gpr_reg[18][0]  ( .D(n564), .CP(clk), .Q(\gpr[18][0] ), .QN(n133) );
  FD1 \gpr_reg[19][31]  ( .D(n563), .CP(clk), .Q(\gpr[19][31] ), .QN(n1663) );
  FD1 \gpr_reg[19][30]  ( .D(n562), .CP(clk), .Q(\gpr[19][30] ), .QN(n1662) );
  FD1 \gpr_reg[19][29]  ( .D(n561), .CP(clk), .Q(\gpr[19][29] ), .QN(n1661) );
  FD1 \gpr_reg[19][28]  ( .D(n560), .CP(clk), .Q(\gpr[19][28] ), .QN(n1660) );
  FD1 \gpr_reg[19][27]  ( .D(n559), .CP(clk), .Q(\gpr[19][27] ), .QN(n1659) );
  FD1 \gpr_reg[19][26]  ( .D(n558), .CP(clk), .Q(\gpr[19][26] ), .QN(n1658) );
  FD1 \gpr_reg[19][25]  ( .D(n557), .CP(clk), .Q(\gpr[19][25] ), .QN(n1657) );
  FD1 \gpr_reg[19][24]  ( .D(n556), .CP(clk), .Q(\gpr[19][24] ), .QN(n1656) );
  FD1 \gpr_reg[19][23]  ( .D(n555), .CP(clk), .Q(\gpr[19][23] ), .QN(n1655) );
  FD1 \gpr_reg[19][22]  ( .D(n554), .CP(clk), .Q(\gpr[19][22] ), .QN(n1654) );
  FD1 \gpr_reg[19][21]  ( .D(n553), .CP(clk), .Q(\gpr[19][21] ), .QN(n1653) );
  FD1 \gpr_reg[19][20]  ( .D(n552), .CP(clk), .Q(\gpr[19][20] ), .QN(n1652) );
  FD1 \gpr_reg[19][19]  ( .D(n551), .CP(clk), .Q(\gpr[19][19] ), .QN(n1651) );
  FD1 \gpr_reg[19][18]  ( .D(n550), .CP(clk), .Q(\gpr[19][18] ), .QN(n1650) );
  FD1 \gpr_reg[19][17]  ( .D(n549), .CP(clk), .Q(\gpr[19][17] ), .QN(n1649) );
  FD1 \gpr_reg[19][16]  ( .D(n548), .CP(clk), .Q(\gpr[19][16] ), .QN(n1648) );
  FD1 \gpr_reg[19][15]  ( .D(n547), .CP(clk), .Q(\gpr[19][15] ), .QN(n1647) );
  FD1 \gpr_reg[19][14]  ( .D(n546), .CP(clk), .Q(\gpr[19][14] ), .QN(n1646) );
  FD1 \gpr_reg[19][13]  ( .D(n545), .CP(clk), .Q(\gpr[19][13] ), .QN(n1645) );
  FD1 \gpr_reg[19][12]  ( .D(n544), .CP(clk), .Q(\gpr[19][12] ), .QN(n1644) );
  FD1 \gpr_reg[19][11]  ( .D(n543), .CP(clk), .Q(\gpr[19][11] ), .QN(n1643) );
  FD1 \gpr_reg[19][10]  ( .D(n542), .CP(clk), .Q(\gpr[19][10] ), .QN(n1642) );
  FD1 \gpr_reg[19][9]  ( .D(n541), .CP(clk), .Q(\gpr[19][9] ), .QN(n1641) );
  FD1 \gpr_reg[19][8]  ( .D(n540), .CP(clk), .Q(\gpr[19][8] ), .QN(n1640) );
  FD1 \gpr_reg[19][7]  ( .D(n539), .CP(clk), .Q(\gpr[19][7] ), .QN(n1639) );
  FD1 \gpr_reg[19][6]  ( .D(n538), .CP(clk), .Q(\gpr[19][6] ), .QN(n1638) );
  FD1 \gpr_reg[19][5]  ( .D(n537), .CP(clk), .Q(\gpr[19][5] ), .QN(n1637) );
  FD1 \gpr_reg[19][4]  ( .D(n536), .CP(clk), .Q(\gpr[19][4] ), .QN(n1636) );
  FD1 \gpr_reg[19][3]  ( .D(n535), .CP(clk), .Q(\gpr[19][3] ), .QN(n1635) );
  FD1 \gpr_reg[19][2]  ( .D(n534), .CP(clk), .Q(\gpr[19][2] ), .QN(n70) );
  FD1 \gpr_reg[19][1]  ( .D(n533), .CP(clk), .Q(\gpr[19][1] ), .QN(n67) );
  FD1 \gpr_reg[19][0]  ( .D(n532), .CP(clk), .Q(\gpr[19][0] ), .QN(n64) );
  FD1 \gpr_reg[20][31]  ( .D(n531), .CP(clk), .Q(\gpr[20][31] ), .QN(n1691) );
  FD1 \gpr_reg[20][30]  ( .D(n530), .CP(clk), .Q(\gpr[20][30] ), .QN(n1690) );
  FD1 \gpr_reg[20][29]  ( .D(n529), .CP(clk), .Q(\gpr[20][29] ), .QN(n1689) );
  FD1 \gpr_reg[20][28]  ( .D(n528), .CP(clk), .Q(\gpr[20][28] ), .QN(n1688) );
  FD1 \gpr_reg[20][27]  ( .D(n527), .CP(clk), .Q(\gpr[20][27] ), .QN(n1687) );
  FD1 \gpr_reg[20][26]  ( .D(n526), .CP(clk), .Q(\gpr[20][26] ), .QN(n1686) );
  FD1 \gpr_reg[20][25]  ( .D(n525), .CP(clk), .Q(\gpr[20][25] ), .QN(n1685) );
  FD1 \gpr_reg[20][24]  ( .D(n524), .CP(clk), .Q(\gpr[20][24] ), .QN(n1684) );
  FD1 \gpr_reg[20][23]  ( .D(n523), .CP(clk), .Q(\gpr[20][23] ), .QN(n1683) );
  FD1 \gpr_reg[20][22]  ( .D(n522), .CP(clk), .Q(\gpr[20][22] ), .QN(n1682) );
  FD1 \gpr_reg[20][21]  ( .D(n521), .CP(clk), .Q(\gpr[20][21] ), .QN(n1681) );
  FD1 \gpr_reg[20][20]  ( .D(n520), .CP(clk), .Q(\gpr[20][20] ), .QN(n1680) );
  FD1 \gpr_reg[20][19]  ( .D(n519), .CP(clk), .Q(\gpr[20][19] ), .QN(n1679) );
  FD1 \gpr_reg[20][18]  ( .D(n518), .CP(clk), .Q(\gpr[20][18] ), .QN(n1678) );
  FD1 \gpr_reg[20][17]  ( .D(n517), .CP(clk), .Q(\gpr[20][17] ), .QN(n1677) );
  FD1 \gpr_reg[20][16]  ( .D(n516), .CP(clk), .Q(\gpr[20][16] ), .QN(n1676) );
  FD1 \gpr_reg[20][15]  ( .D(n515), .CP(clk), .Q(\gpr[20][15] ), .QN(n1675) );
  FD1 \gpr_reg[20][14]  ( .D(n514), .CP(clk), .Q(\gpr[20][14] ), .QN(n1674) );
  FD1 \gpr_reg[20][13]  ( .D(n513), .CP(clk), .Q(\gpr[20][13] ), .QN(n1673) );
  FD1 \gpr_reg[20][12]  ( .D(n512), .CP(clk), .Q(\gpr[20][12] ), .QN(n1672) );
  FD1 \gpr_reg[20][11]  ( .D(n511), .CP(clk), .Q(\gpr[20][11] ), .QN(n1671) );
  FD1 \gpr_reg[20][10]  ( .D(n510), .CP(clk), .Q(\gpr[20][10] ), .QN(n1670) );
  FD1 \gpr_reg[20][9]  ( .D(n509), .CP(clk), .Q(\gpr[20][9] ), .QN(n1669) );
  FD1 \gpr_reg[20][8]  ( .D(n508), .CP(clk), .Q(\gpr[20][8] ), .QN(n1668) );
  FD1 \gpr_reg[20][7]  ( .D(n507), .CP(clk), .Q(\gpr[20][7] ), .QN(n1667) );
  FD1 \gpr_reg[20][6]  ( .D(n506), .CP(clk), .Q(\gpr[20][6] ), .QN(n1666) );
  FD1 \gpr_reg[20][5]  ( .D(n505), .CP(clk), .Q(\gpr[20][5] ), .QN(n1665) );
  FD1 \gpr_reg[20][3]  ( .D(n503), .CP(clk), .Q(\gpr[20][3] ), .QN(n1664) );
  FD1 \gpr_reg[20][2]  ( .D(n502), .CP(clk), .Q(\gpr[20][2] ), .QN(n55) );
  FD1 \gpr_reg[20][1]  ( .D(n501), .CP(clk), .Q(\gpr[20][1] ), .QN(n54) );
  FD1 \gpr_reg[20][0]  ( .D(n500), .CP(clk), .Q(\gpr[20][0] ), .QN(n59) );
  FD1 \gpr_reg[21][31]  ( .D(n499), .CP(clk), .Q(\gpr[21][31] ), .QN(n1720) );
  FD1 \gpr_reg[21][30]  ( .D(n498), .CP(clk), .Q(\gpr[21][30] ), .QN(n1719) );
  FD1 \gpr_reg[21][29]  ( .D(n497), .CP(clk), .Q(\gpr[21][29] ), .QN(n1718) );
  FD1 \gpr_reg[21][28]  ( .D(n496), .CP(clk), .Q(\gpr[21][28] ), .QN(n1717) );
  FD1 \gpr_reg[21][27]  ( .D(n495), .CP(clk), .Q(\gpr[21][27] ), .QN(n1716) );
  FD1 \gpr_reg[21][26]  ( .D(n494), .CP(clk), .Q(\gpr[21][26] ), .QN(n1715) );
  FD1 \gpr_reg[21][25]  ( .D(n493), .CP(clk), .Q(\gpr[21][25] ), .QN(n1714) );
  FD1 \gpr_reg[21][24]  ( .D(n492), .CP(clk), .Q(\gpr[21][24] ), .QN(n1713) );
  FD1 \gpr_reg[21][23]  ( .D(n491), .CP(clk), .Q(\gpr[21][23] ), .QN(n1712) );
  FD1 \gpr_reg[21][22]  ( .D(n490), .CP(clk), .Q(\gpr[21][22] ), .QN(n1711) );
  FD1 \gpr_reg[21][21]  ( .D(n489), .CP(clk), .Q(\gpr[21][21] ), .QN(n1710) );
  FD1 \gpr_reg[21][20]  ( .D(n488), .CP(clk), .Q(\gpr[21][20] ), .QN(n1709) );
  FD1 \gpr_reg[21][19]  ( .D(n487), .CP(clk), .Q(\gpr[21][19] ), .QN(n1708) );
  FD1 \gpr_reg[21][18]  ( .D(n486), .CP(clk), .Q(\gpr[21][18] ), .QN(n1707) );
  FD1 \gpr_reg[21][17]  ( .D(n485), .CP(clk), .Q(\gpr[21][17] ), .QN(n1706) );
  FD1 \gpr_reg[21][16]  ( .D(n484), .CP(clk), .Q(\gpr[21][16] ), .QN(n1705) );
  FD1 \gpr_reg[21][15]  ( .D(n483), .CP(clk), .Q(\gpr[21][15] ), .QN(n1704) );
  FD1 \gpr_reg[21][14]  ( .D(n482), .CP(clk), .Q(\gpr[21][14] ), .QN(n1703) );
  FD1 \gpr_reg[21][13]  ( .D(n481), .CP(clk), .Q(\gpr[21][13] ), .QN(n1702) );
  FD1 \gpr_reg[21][12]  ( .D(n480), .CP(clk), .Q(\gpr[21][12] ), .QN(n1701) );
  FD1 \gpr_reg[21][11]  ( .D(n479), .CP(clk), .Q(\gpr[21][11] ), .QN(n1700) );
  FD1 \gpr_reg[21][10]  ( .D(n478), .CP(clk), .Q(\gpr[21][10] ), .QN(n1699) );
  FD1 \gpr_reg[21][9]  ( .D(n477), .CP(clk), .Q(\gpr[21][9] ), .QN(n1698) );
  FD1 \gpr_reg[21][8]  ( .D(n476), .CP(clk), .Q(\gpr[21][8] ), .QN(n1697) );
  FD1 \gpr_reg[21][7]  ( .D(n475), .CP(clk), .Q(\gpr[21][7] ), .QN(n1696) );
  FD1 \gpr_reg[21][6]  ( .D(n474), .CP(clk), .Q(\gpr[21][6] ), .QN(n1695) );
  FD1 \gpr_reg[21][5]  ( .D(n473), .CP(clk), .Q(\gpr[21][5] ), .QN(n1694) );
  FD1 \gpr_reg[21][4]  ( .D(n472), .CP(clk), .Q(\gpr[21][4] ), .QN(n1693) );
  FD1 \gpr_reg[21][3]  ( .D(n471), .CP(clk), .Q(\gpr[21][3] ), .QN(n1692) );
  FD1 \gpr_reg[21][2]  ( .D(n470), .CP(clk), .Q(\gpr[21][2] ), .QN(n124) );
  FD1 \gpr_reg[21][1]  ( .D(n469), .CP(clk), .Q(\gpr[21][1] ), .QN(n123) );
  FD1 \gpr_reg[21][0]  ( .D(n468), .CP(clk), .Q(\gpr[21][0] ), .QN(n128) );
  FD1 \gpr_reg[22][31]  ( .D(n467), .CP(clk), .Q(\gpr[22][31] ), .QN(n1751) );
  FD1 \gpr_reg[22][30]  ( .D(n466), .CP(clk), .Q(\gpr[22][30] ), .QN(n1750) );
  FD1 \gpr_reg[22][29]  ( .D(n465), .CP(clk), .Q(\gpr[22][29] ), .QN(n1749) );
  FD1 \gpr_reg[22][28]  ( .D(n464), .CP(clk), .Q(\gpr[22][28] ), .QN(n1748) );
  FD1 \gpr_reg[22][27]  ( .D(n463), .CP(clk), .Q(\gpr[22][27] ), .QN(n1747) );
  FD1 \gpr_reg[22][26]  ( .D(n462), .CP(clk), .Q(\gpr[22][26] ), .QN(n1746) );
  FD1 \gpr_reg[22][25]  ( .D(n461), .CP(clk), .Q(\gpr[22][25] ), .QN(n1745) );
  FD1 \gpr_reg[22][24]  ( .D(n460), .CP(clk), .Q(\gpr[22][24] ), .QN(n1744) );
  FD1 \gpr_reg[22][23]  ( .D(n459), .CP(clk), .Q(\gpr[22][23] ), .QN(n1743) );
  FD1 \gpr_reg[22][22]  ( .D(n458), .CP(clk), .Q(\gpr[22][22] ), .QN(n1742) );
  FD1 \gpr_reg[22][21]  ( .D(n457), .CP(clk), .Q(\gpr[22][21] ), .QN(n1741) );
  FD1 \gpr_reg[22][20]  ( .D(n456), .CP(clk), .Q(\gpr[22][20] ), .QN(n1740) );
  FD1 \gpr_reg[22][19]  ( .D(n455), .CP(clk), .Q(\gpr[22][19] ), .QN(n1739) );
  FD1 \gpr_reg[22][18]  ( .D(n454), .CP(clk), .Q(\gpr[22][18] ), .QN(n1738) );
  FD1 \gpr_reg[22][17]  ( .D(n453), .CP(clk), .Q(\gpr[22][17] ), .QN(n1737) );
  FD1 \gpr_reg[22][16]  ( .D(n452), .CP(clk), .Q(\gpr[22][16] ), .QN(n1736) );
  FD1 \gpr_reg[22][15]  ( .D(n451), .CP(clk), .Q(\gpr[22][15] ), .QN(n1735) );
  FD1 \gpr_reg[22][14]  ( .D(n450), .CP(clk), .Q(\gpr[22][14] ), .QN(n1734) );
  FD1 \gpr_reg[22][13]  ( .D(n449), .CP(clk), .Q(\gpr[22][13] ), .QN(n1733) );
  FD1 \gpr_reg[22][12]  ( .D(n448), .CP(clk), .Q(\gpr[22][12] ), .QN(n1732) );
  FD1 \gpr_reg[22][11]  ( .D(n447), .CP(clk), .Q(\gpr[22][11] ), .QN(n1731) );
  FD1 \gpr_reg[22][10]  ( .D(n446), .CP(clk), .Q(\gpr[22][10] ), .QN(n1730) );
  FD1 \gpr_reg[22][9]  ( .D(n445), .CP(clk), .Q(\gpr[22][9] ), .QN(n1729) );
  FD1 \gpr_reg[22][8]  ( .D(n444), .CP(clk), .Q(\gpr[22][8] ), .QN(n1728) );
  FD1 \gpr_reg[22][7]  ( .D(n443), .CP(clk), .Q(\gpr[22][7] ), .QN(n1727) );
  FD1 \gpr_reg[22][6]  ( .D(n442), .CP(clk), .Q(\gpr[22][6] ), .QN(n1726) );
  FD1 \gpr_reg[22][5]  ( .D(n441), .CP(clk), .Q(\gpr[22][5] ), .QN(n1725) );
  FD1 \gpr_reg[22][4]  ( .D(n440), .CP(clk), .Q(\gpr[22][4] ), .QN(n1724) );
  FD1 \gpr_reg[22][3]  ( .D(n439), .CP(clk), .Q(\gpr[22][3] ), .QN(n1723) );
  FD1 \gpr_reg[22][1]  ( .D(n437), .CP(clk), .Q(\gpr[22][1] ), .QN(n1722) );
  FD1 \gpr_reg[22][0]  ( .D(n436), .CP(clk), .Q(\gpr[22][0] ), .QN(n1721) );
  FD1 \gpr_reg[23][31]  ( .D(n435), .CP(clk), .Q(\gpr[23][31] ), .QN(n1782) );
  FD1 \gpr_reg[23][30]  ( .D(n434), .CP(clk), .Q(\gpr[23][30] ), .QN(n1781) );
  FD1 \gpr_reg[23][29]  ( .D(n433), .CP(clk), .Q(\gpr[23][29] ), .QN(n1780) );
  FD1 \gpr_reg[23][28]  ( .D(n432), .CP(clk), .Q(\gpr[23][28] ), .QN(n1779) );
  FD1 \gpr_reg[23][27]  ( .D(n431), .CP(clk), .Q(\gpr[23][27] ), .QN(n1778) );
  FD1 \gpr_reg[23][26]  ( .D(n430), .CP(clk), .Q(\gpr[23][26] ), .QN(n1777) );
  FD1 \gpr_reg[23][25]  ( .D(n429), .CP(clk), .Q(\gpr[23][25] ), .QN(n1776) );
  FD1 \gpr_reg[23][24]  ( .D(n428), .CP(clk), .Q(\gpr[23][24] ), .QN(n1775) );
  FD1 \gpr_reg[23][23]  ( .D(n427), .CP(clk), .Q(\gpr[23][23] ), .QN(n1774) );
  FD1 \gpr_reg[23][22]  ( .D(n426), .CP(clk), .Q(\gpr[23][22] ), .QN(n1773) );
  FD1 \gpr_reg[23][21]  ( .D(n425), .CP(clk), .Q(\gpr[23][21] ), .QN(n1772) );
  FD1 \gpr_reg[23][20]  ( .D(n424), .CP(clk), .Q(\gpr[23][20] ), .QN(n1771) );
  FD1 \gpr_reg[23][19]  ( .D(n423), .CP(clk), .Q(\gpr[23][19] ), .QN(n1770) );
  FD1 \gpr_reg[23][18]  ( .D(n422), .CP(clk), .Q(\gpr[23][18] ), .QN(n1769) );
  FD1 \gpr_reg[23][17]  ( .D(n421), .CP(clk), .Q(\gpr[23][17] ), .QN(n1768) );
  FD1 \gpr_reg[23][16]  ( .D(n420), .CP(clk), .Q(\gpr[23][16] ), .QN(n1767) );
  FD1 \gpr_reg[23][15]  ( .D(n419), .CP(clk), .Q(\gpr[23][15] ), .QN(n1766) );
  FD1 \gpr_reg[23][14]  ( .D(n418), .CP(clk), .Q(\gpr[23][14] ), .QN(n1765) );
  FD1 \gpr_reg[23][13]  ( .D(n417), .CP(clk), .Q(\gpr[23][13] ), .QN(n1764) );
  FD1 \gpr_reg[23][12]  ( .D(n416), .CP(clk), .Q(\gpr[23][12] ), .QN(n1763) );
  FD1 \gpr_reg[23][11]  ( .D(n415), .CP(clk), .Q(\gpr[23][11] ), .QN(n1762) );
  FD1 \gpr_reg[23][10]  ( .D(n414), .CP(clk), .Q(\gpr[23][10] ), .QN(n1761) );
  FD1 \gpr_reg[23][9]  ( .D(n413), .CP(clk), .Q(\gpr[23][9] ), .QN(n1760) );
  FD1 \gpr_reg[23][8]  ( .D(n412), .CP(clk), .Q(\gpr[23][8] ), .QN(n1759) );
  FD1 \gpr_reg[23][7]  ( .D(n411), .CP(clk), .Q(\gpr[23][7] ), .QN(n1758) );
  FD1 \gpr_reg[23][6]  ( .D(n410), .CP(clk), .Q(\gpr[23][6] ), .QN(n1757) );
  FD1 \gpr_reg[23][5]  ( .D(n409), .CP(clk), .Q(\gpr[23][5] ), .QN(n1756) );
  FD1 \gpr_reg[23][4]  ( .D(n408), .CP(clk), .Q(\gpr[23][4] ), .QN(n1755) );
  FD1 \gpr_reg[23][3]  ( .D(n407), .CP(clk), .Q(\gpr[23][3] ), .QN(n1754) );
  FD1 \gpr_reg[23][1]  ( .D(n405), .CP(clk), .Q(\gpr[23][1] ), .QN(n1753) );
  FD1 \gpr_reg[23][0]  ( .D(n404), .CP(clk), .Q(\gpr[23][0] ), .QN(n1752) );
  FD1 \gpr_reg[24][31]  ( .D(n403), .CP(clk), .Q(\gpr[24][31] ), .QN(n1811) );
  FD1 \gpr_reg[24][30]  ( .D(n402), .CP(clk), .Q(\gpr[24][30] ), .QN(n1810) );
  FD1 \gpr_reg[24][29]  ( .D(n401), .CP(clk), .Q(\gpr[24][29] ), .QN(n1809) );
  FD1 \gpr_reg[24][28]  ( .D(n400), .CP(clk), .Q(\gpr[24][28] ), .QN(n1808) );
  FD1 \gpr_reg[24][27]  ( .D(n399), .CP(clk), .Q(\gpr[24][27] ), .QN(n1807) );
  FD1 \gpr_reg[24][26]  ( .D(n398), .CP(clk), .Q(\gpr[24][26] ), .QN(n1806) );
  FD1 \gpr_reg[24][25]  ( .D(n397), .CP(clk), .Q(\gpr[24][25] ), .QN(n1805) );
  FD1 \gpr_reg[24][24]  ( .D(n396), .CP(clk), .Q(\gpr[24][24] ), .QN(n1804) );
  FD1 \gpr_reg[24][23]  ( .D(n395), .CP(clk), .Q(\gpr[24][23] ), .QN(n1803) );
  FD1 \gpr_reg[24][22]  ( .D(n394), .CP(clk), .Q(\gpr[24][22] ), .QN(n1802) );
  FD1 \gpr_reg[24][21]  ( .D(n393), .CP(clk), .Q(\gpr[24][21] ), .QN(n1801) );
  FD1 \gpr_reg[24][20]  ( .D(n392), .CP(clk), .Q(\gpr[24][20] ), .QN(n1800) );
  FD1 \gpr_reg[24][19]  ( .D(n391), .CP(clk), .Q(\gpr[24][19] ), .QN(n1799) );
  FD1 \gpr_reg[24][18]  ( .D(n390), .CP(clk), .Q(\gpr[24][18] ), .QN(n1798) );
  FD1 \gpr_reg[24][17]  ( .D(n389), .CP(clk), .Q(\gpr[24][17] ), .QN(n1797) );
  FD1 \gpr_reg[24][16]  ( .D(n388), .CP(clk), .Q(\gpr[24][16] ), .QN(n1796) );
  FD1 \gpr_reg[24][15]  ( .D(n387), .CP(clk), .Q(\gpr[24][15] ), .QN(n1795) );
  FD1 \gpr_reg[24][14]  ( .D(n386), .CP(clk), .Q(\gpr[24][14] ), .QN(n1794) );
  FD1 \gpr_reg[24][13]  ( .D(n385), .CP(clk), .Q(\gpr[24][13] ), .QN(n1793) );
  FD1 \gpr_reg[24][12]  ( .D(n384), .CP(clk), .Q(\gpr[24][12] ), .QN(n1792) );
  FD1 \gpr_reg[24][11]  ( .D(n383), .CP(clk), .Q(\gpr[24][11] ), .QN(n1791) );
  FD1 \gpr_reg[24][10]  ( .D(n382), .CP(clk), .Q(\gpr[24][10] ), .QN(n1790) );
  FD1 \gpr_reg[24][9]  ( .D(n381), .CP(clk), .Q(\gpr[24][9] ), .QN(n1789) );
  FD1 \gpr_reg[24][8]  ( .D(n380), .CP(clk), .Q(\gpr[24][8] ), .QN(n1788) );
  FD1 \gpr_reg[24][7]  ( .D(n379), .CP(clk), .Q(\gpr[24][7] ), .QN(n1787) );
  FD1 \gpr_reg[24][6]  ( .D(n378), .CP(clk), .Q(\gpr[24][6] ), .QN(n1786) );
  FD1 \gpr_reg[24][5]  ( .D(n377), .CP(clk), .Q(\gpr[24][5] ), .QN(n1785) );
  FD1 \gpr_reg[24][4]  ( .D(n376), .CP(clk), .Q(\gpr[24][4] ), .QN(n1784) );
  FD1 \gpr_reg[24][3]  ( .D(n375), .CP(clk), .Q(\gpr[24][3] ), .QN(n1783) );
  FD1 \gpr_reg[24][2]  ( .D(n374), .CP(clk), .Q(\gpr[24][2] ), .QN(n58) );
  FD1 \gpr_reg[24][1]  ( .D(n373), .CP(clk), .Q(\gpr[24][1] ), .QN(n57) );
  FD1 \gpr_reg[24][0]  ( .D(n372), .CP(clk), .Q(\gpr[24][0] ), .QN(n56) );
  FD1 \gpr_reg[25][31]  ( .D(n371), .CP(clk), .Q(\gpr[25][31] ), .QN(n1838) );
  FD1 \gpr_reg[25][30]  ( .D(n370), .CP(clk), .Q(\gpr[25][30] ), .QN(n1837) );
  FD1 \gpr_reg[25][29]  ( .D(n369), .CP(clk), .Q(\gpr[25][29] ), .QN(n1836) );
  FD1 \gpr_reg[25][28]  ( .D(n368), .CP(clk), .Q(\gpr[25][28] ), .QN(n1835) );
  FD1 \gpr_reg[25][27]  ( .D(n367), .CP(clk), .Q(\gpr[25][27] ), .QN(n1834) );
  FD1 \gpr_reg[25][26]  ( .D(n366), .CP(clk), .Q(\gpr[25][26] ), .QN(n1833) );
  FD1 \gpr_reg[25][25]  ( .D(n365), .CP(clk), .Q(\gpr[25][25] ), .QN(n1832) );
  FD1 \gpr_reg[25][24]  ( .D(n364), .CP(clk), .Q(\gpr[25][24] ), .QN(n1831) );
  FD1 \gpr_reg[25][23]  ( .D(n363), .CP(clk), .Q(\gpr[25][23] ), .QN(n1830) );
  FD1 \gpr_reg[25][22]  ( .D(n362), .CP(clk), .Q(\gpr[25][22] ), .QN(n1829) );
  FD1 \gpr_reg[25][21]  ( .D(n361), .CP(clk), .Q(\gpr[25][21] ), .QN(n1828) );
  FD1 \gpr_reg[25][20]  ( .D(n360), .CP(clk), .Q(\gpr[25][20] ), .QN(n1827) );
  FD1 \gpr_reg[25][19]  ( .D(n359), .CP(clk), .Q(\gpr[25][19] ), .QN(n1826) );
  FD1 \gpr_reg[25][18]  ( .D(n358), .CP(clk), .Q(\gpr[25][18] ), .QN(n1825) );
  FD1 \gpr_reg[25][17]  ( .D(n357), .CP(clk), .Q(\gpr[25][17] ), .QN(n1824) );
  FD1 \gpr_reg[25][16]  ( .D(n356), .CP(clk), .Q(\gpr[25][16] ), .QN(n1823) );
  FD1 \gpr_reg[25][15]  ( .D(n355), .CP(clk), .Q(\gpr[25][15] ), .QN(n1822) );
  FD1 \gpr_reg[25][14]  ( .D(n354), .CP(clk), .Q(\gpr[25][14] ), .QN(n1821) );
  FD1 \gpr_reg[25][13]  ( .D(n353), .CP(clk), .Q(\gpr[25][13] ), .QN(n1820) );
  FD1 \gpr_reg[25][12]  ( .D(n352), .CP(clk), .Q(\gpr[25][12] ), .QN(n1819) );
  FD1 \gpr_reg[25][11]  ( .D(n351), .CP(clk), .Q(\gpr[25][11] ), .QN(n1818) );
  FD1 \gpr_reg[25][10]  ( .D(n350), .CP(clk), .Q(\gpr[25][10] ), .QN(n1817) );
  FD1 \gpr_reg[25][8]  ( .D(n348), .CP(clk), .Q(\gpr[25][8] ), .QN(n1816) );
  FD1 \gpr_reg[25][7]  ( .D(n347), .CP(clk), .Q(\gpr[25][7] ), .QN(n1815) );
  FD1 \gpr_reg[25][6]  ( .D(n346), .CP(clk), .Q(\gpr[25][6] ), .QN(n1814) );
  FD1 \gpr_reg[25][4]  ( .D(n344), .CP(clk), .Q(\gpr[25][4] ), .QN(n1813) );
  FD1 \gpr_reg[25][3]  ( .D(n343), .CP(clk), .Q(\gpr[25][3] ), .QN(n1812) );
  FD1 \gpr_reg[25][2]  ( .D(n342), .CP(clk), .Q(\gpr[25][2] ), .QN(n127) );
  FD1 \gpr_reg[25][1]  ( .D(n341), .CP(clk), .Q(\gpr[25][1] ), .QN(n126) );
  FD1 \gpr_reg[25][0]  ( .D(n340), .CP(clk), .Q(\gpr[25][0] ), .QN(n125) );
  FD1 \gpr_reg[26][31]  ( .D(n339), .CP(clk), .Q(\gpr[26][31] ), .QN(n1869) );
  FD1 \gpr_reg[26][30]  ( .D(n338), .CP(clk), .Q(\gpr[26][30] ), .QN(n1868) );
  FD1 \gpr_reg[26][29]  ( .D(n337), .CP(clk), .Q(\gpr[26][29] ), .QN(n1867) );
  FD1 \gpr_reg[26][28]  ( .D(n336), .CP(clk), .Q(\gpr[26][28] ), .QN(n1866) );
  FD1 \gpr_reg[26][27]  ( .D(n335), .CP(clk), .Q(\gpr[26][27] ), .QN(n1865) );
  FD1 \gpr_reg[26][26]  ( .D(n334), .CP(clk), .Q(\gpr[26][26] ), .QN(n1864) );
  FD1 \gpr_reg[26][25]  ( .D(n333), .CP(clk), .Q(\gpr[26][25] ), .QN(n1863) );
  FD1 \gpr_reg[26][24]  ( .D(n332), .CP(clk), .Q(\gpr[26][24] ), .QN(n1862) );
  FD1 \gpr_reg[26][23]  ( .D(n331), .CP(clk), .Q(\gpr[26][23] ), .QN(n1861) );
  FD1 \gpr_reg[26][22]  ( .D(n330), .CP(clk), .Q(\gpr[26][22] ), .QN(n1860) );
  FD1 \gpr_reg[26][21]  ( .D(n329), .CP(clk), .Q(\gpr[26][21] ), .QN(n1859) );
  FD1 \gpr_reg[26][20]  ( .D(n328), .CP(clk), .Q(\gpr[26][20] ), .QN(n1858) );
  FD1 \gpr_reg[26][19]  ( .D(n327), .CP(clk), .Q(\gpr[26][19] ), .QN(n1857) );
  FD1 \gpr_reg[26][18]  ( .D(n326), .CP(clk), .Q(\gpr[26][18] ), .QN(n1856) );
  FD1 \gpr_reg[26][17]  ( .D(n325), .CP(clk), .Q(\gpr[26][17] ), .QN(n1855) );
  FD1 \gpr_reg[26][16]  ( .D(n324), .CP(clk), .Q(\gpr[26][16] ), .QN(n1854) );
  FD1 \gpr_reg[26][15]  ( .D(n323), .CP(clk), .Q(\gpr[26][15] ), .QN(n1853) );
  FD1 \gpr_reg[26][14]  ( .D(n322), .CP(clk), .Q(\gpr[26][14] ), .QN(n1852) );
  FD1 \gpr_reg[26][13]  ( .D(n321), .CP(clk), .Q(\gpr[26][13] ), .QN(n1851) );
  FD1 \gpr_reg[26][12]  ( .D(n320), .CP(clk), .Q(\gpr[26][12] ), .QN(n1850) );
  FD1 \gpr_reg[26][11]  ( .D(n319), .CP(clk), .Q(\gpr[26][11] ), .QN(n1849) );
  FD1 \gpr_reg[26][10]  ( .D(n318), .CP(clk), .Q(\gpr[26][10] ), .QN(n1848) );
  FD1 \gpr_reg[26][9]  ( .D(n317), .CP(clk), .Q(\gpr[26][9] ), .QN(n1847) );
  FD1 \gpr_reg[26][8]  ( .D(n316), .CP(clk), .Q(\gpr[26][8] ), .QN(n1846) );
  FD1 \gpr_reg[26][7]  ( .D(n315), .CP(clk), .Q(\gpr[26][7] ), .QN(n1845) );
  FD1 \gpr_reg[26][6]  ( .D(n314), .CP(clk), .Q(\gpr[26][6] ), .QN(n1844) );
  FD1 \gpr_reg[26][5]  ( .D(n313), .CP(clk), .Q(\gpr[26][5] ), .QN(n1843) );
  FD1 \gpr_reg[26][4]  ( .D(n312), .CP(clk), .Q(\gpr[26][4] ), .QN(n1842) );
  FD1 \gpr_reg[26][3]  ( .D(n311), .CP(clk), .Q(\gpr[26][3] ), .QN(n1841) );
  FD1 \gpr_reg[26][1]  ( .D(n309), .CP(clk), .Q(\gpr[26][1] ), .QN(n1840) );
  FD1 \gpr_reg[26][0]  ( .D(n308), .CP(clk), .Q(\gpr[26][0] ), .QN(n1839) );
  FD1 \gpr_reg[27][31]  ( .D(n307), .CP(clk), .Q(\gpr[27][31] ), .QN(n1900) );
  FD1 \gpr_reg[27][30]  ( .D(n306), .CP(clk), .Q(\gpr[27][30] ), .QN(n1899) );
  FD1 \gpr_reg[27][29]  ( .D(n305), .CP(clk), .Q(\gpr[27][29] ), .QN(n1898) );
  FD1 \gpr_reg[27][28]  ( .D(n304), .CP(clk), .Q(\gpr[27][28] ), .QN(n1897) );
  FD1 \gpr_reg[27][27]  ( .D(n303), .CP(clk), .Q(\gpr[27][27] ), .QN(n1896) );
  FD1 \gpr_reg[27][26]  ( .D(n302), .CP(clk), .Q(\gpr[27][26] ), .QN(n1895) );
  FD1 \gpr_reg[27][25]  ( .D(n301), .CP(clk), .Q(\gpr[27][25] ), .QN(n1894) );
  FD1 \gpr_reg[27][24]  ( .D(n300), .CP(clk), .Q(\gpr[27][24] ), .QN(n1893) );
  FD1 \gpr_reg[27][23]  ( .D(n299), .CP(clk), .Q(\gpr[27][23] ), .QN(n1892) );
  FD1 \gpr_reg[27][22]  ( .D(n298), .CP(clk), .Q(\gpr[27][22] ), .QN(n1891) );
  FD1 \gpr_reg[27][21]  ( .D(n297), .CP(clk), .Q(\gpr[27][21] ), .QN(n1890) );
  FD1 \gpr_reg[27][20]  ( .D(n296), .CP(clk), .Q(\gpr[27][20] ), .QN(n1889) );
  FD1 \gpr_reg[27][19]  ( .D(n295), .CP(clk), .Q(\gpr[27][19] ), .QN(n1888) );
  FD1 \gpr_reg[27][18]  ( .D(n294), .CP(clk), .Q(\gpr[27][18] ), .QN(n1887) );
  FD1 \gpr_reg[27][17]  ( .D(n293), .CP(clk), .Q(\gpr[27][17] ), .QN(n1886) );
  FD1 \gpr_reg[27][16]  ( .D(n292), .CP(clk), .Q(\gpr[27][16] ), .QN(n1885) );
  FD1 \gpr_reg[27][15]  ( .D(n291), .CP(clk), .Q(\gpr[27][15] ), .QN(n1884) );
  FD1 \gpr_reg[27][14]  ( .D(n290), .CP(clk), .Q(\gpr[27][14] ), .QN(n1883) );
  FD1 \gpr_reg[27][13]  ( .D(n289), .CP(clk), .Q(\gpr[27][13] ), .QN(n1882) );
  FD1 \gpr_reg[27][12]  ( .D(n288), .CP(clk), .Q(\gpr[27][12] ), .QN(n1881) );
  FD1 \gpr_reg[27][11]  ( .D(n287), .CP(clk), .Q(\gpr[27][11] ), .QN(n1880) );
  FD1 \gpr_reg[27][10]  ( .D(n286), .CP(clk), .Q(\gpr[27][10] ), .QN(n1879) );
  FD1 \gpr_reg[27][9]  ( .D(n285), .CP(clk), .Q(\gpr[27][9] ), .QN(n1878) );
  FD1 \gpr_reg[27][8]  ( .D(n284), .CP(clk), .Q(\gpr[27][8] ), .QN(n1877) );
  FD1 \gpr_reg[27][7]  ( .D(n283), .CP(clk), .Q(\gpr[27][7] ), .QN(n1876) );
  FD1 \gpr_reg[27][6]  ( .D(n282), .CP(clk), .Q(\gpr[27][6] ), .QN(n1875) );
  FD1 \gpr_reg[27][5]  ( .D(n281), .CP(clk), .Q(\gpr[27][5] ), .QN(n1874) );
  FD1 \gpr_reg[27][4]  ( .D(n280), .CP(clk), .Q(\gpr[27][4] ), .QN(n1873) );
  FD1 \gpr_reg[27][3]  ( .D(n279), .CP(clk), .Q(\gpr[27][3] ), .QN(n1872) );
  FD1 \gpr_reg[27][2]  ( .D(n278), .CP(clk), .Q(\gpr[27][2] ), .QN(n2092) );
  FD1 \gpr_reg[27][1]  ( .D(n277), .CP(clk), .Q(\gpr[27][1] ), .QN(n1871) );
  FD1 \gpr_reg[27][0]  ( .D(n276), .CP(clk), .Q(\gpr[27][0] ), .QN(n1870) );
  FD1 \gpr_reg[28][31]  ( .D(n275), .CP(clk), .Q(\gpr[28][31] ), .QN(n1931) );
  FD1 \gpr_reg[28][30]  ( .D(n274), .CP(clk), .Q(\gpr[28][30] ), .QN(n1930) );
  FD1 \gpr_reg[28][29]  ( .D(n273), .CP(clk), .Q(\gpr[28][29] ), .QN(n1929) );
  FD1 \gpr_reg[28][28]  ( .D(n272), .CP(clk), .Q(\gpr[28][28] ), .QN(n1928) );
  FD1 \gpr_reg[28][27]  ( .D(n271), .CP(clk), .Q(\gpr[28][27] ), .QN(n1927) );
  FD1 \gpr_reg[28][26]  ( .D(n270), .CP(clk), .Q(\gpr[28][26] ), .QN(n1926) );
  FD1 \gpr_reg[28][25]  ( .D(n269), .CP(clk), .Q(\gpr[28][25] ), .QN(n1925) );
  FD1 \gpr_reg[28][24]  ( .D(n268), .CP(clk), .Q(\gpr[28][24] ), .QN(n1924) );
  FD1 \gpr_reg[28][23]  ( .D(n267), .CP(clk), .Q(\gpr[28][23] ), .QN(n1923) );
  FD1 \gpr_reg[28][22]  ( .D(n266), .CP(clk), .Q(\gpr[28][22] ), .QN(n1922) );
  FD1 \gpr_reg[28][21]  ( .D(n265), .CP(clk), .Q(\gpr[28][21] ), .QN(n1921) );
  FD1 \gpr_reg[28][20]  ( .D(n264), .CP(clk), .Q(\gpr[28][20] ), .QN(n1920) );
  FD1 \gpr_reg[28][19]  ( .D(n263), .CP(clk), .Q(\gpr[28][19] ), .QN(n1919) );
  FD1 \gpr_reg[28][18]  ( .D(n262), .CP(clk), .Q(\gpr[28][18] ), .QN(n1918) );
  FD1 \gpr_reg[28][17]  ( .D(n261), .CP(clk), .Q(\gpr[28][17] ), .QN(n1917) );
  FD1 \gpr_reg[28][16]  ( .D(n260), .CP(clk), .Q(\gpr[28][16] ), .QN(n1916) );
  FD1 \gpr_reg[28][15]  ( .D(n259), .CP(clk), .Q(\gpr[28][15] ), .QN(n1915) );
  FD1 \gpr_reg[28][13]  ( .D(n257), .CP(clk), .Q(\gpr[28][13] ), .QN(n1914) );
  FD1 \gpr_reg[28][12]  ( .D(n256), .CP(clk), .Q(\gpr[28][12] ), .QN(n1913) );
  FD1 \gpr_reg[28][11]  ( .D(n255), .CP(clk), .Q(\gpr[28][11] ), .QN(n1912) );
  FD1 \gpr_reg[28][10]  ( .D(n254), .CP(clk), .Q(\gpr[28][10] ), .QN(n1911) );
  FD1 \gpr_reg[28][9]  ( .D(n253), .CP(clk), .Q(\gpr[28][9] ), .QN(n1910) );
  FD1 \gpr_reg[28][8]  ( .D(n252), .CP(clk), .Q(\gpr[28][8] ), .QN(n1909) );
  FD1 \gpr_reg[28][7]  ( .D(n251), .CP(clk), .Q(\gpr[28][7] ), .QN(n1908) );
  FD1 \gpr_reg[28][6]  ( .D(n250), .CP(clk), .Q(\gpr[28][6] ), .QN(n1907) );
  FD1 \gpr_reg[28][5]  ( .D(n249), .CP(clk), .Q(\gpr[28][5] ), .QN(n1906) );
  FD1 \gpr_reg[28][4]  ( .D(n248), .CP(clk), .Q(\gpr[28][4] ), .QN(n1905) );
  FD1 \gpr_reg[28][3]  ( .D(n247), .CP(clk), .Q(\gpr[28][3] ), .QN(n1904) );
  FD1 \gpr_reg[28][2]  ( .D(n246), .CP(clk), .Q(\gpr[28][2] ), .QN(n1903) );
  FD1 \gpr_reg[28][1]  ( .D(n245), .CP(clk), .Q(\gpr[28][1] ), .QN(n1902) );
  FD1 \gpr_reg[28][0]  ( .D(n244), .CP(clk), .Q(\gpr[28][0] ), .QN(n1901) );
  FD1 \gpr_reg[29][31]  ( .D(n243), .CP(clk), .Q(\gpr[29][31] ), .QN(n1963) );
  FD1 \gpr_reg[29][30]  ( .D(n242), .CP(clk), .Q(\gpr[29][30] ), .QN(n1962) );
  FD1 \gpr_reg[29][29]  ( .D(n241), .CP(clk), .Q(\gpr[29][29] ), .QN(n1961) );
  FD1 \gpr_reg[29][28]  ( .D(n240), .CP(clk), .Q(\gpr[29][28] ), .QN(n1960) );
  FD1 \gpr_reg[29][27]  ( .D(n239), .CP(clk), .Q(\gpr[29][27] ), .QN(n1959) );
  FD1 \gpr_reg[29][26]  ( .D(n238), .CP(clk), .Q(\gpr[29][26] ), .QN(n1958) );
  FD1 \gpr_reg[29][25]  ( .D(n237), .CP(clk), .Q(\gpr[29][25] ), .QN(n1957) );
  FD1 \gpr_reg[29][24]  ( .D(n236), .CP(clk), .Q(\gpr[29][24] ), .QN(n1956) );
  FD1 \gpr_reg[29][23]  ( .D(n235), .CP(clk), .Q(\gpr[29][23] ), .QN(n1955) );
  FD1 \gpr_reg[29][22]  ( .D(n234), .CP(clk), .Q(\gpr[29][22] ), .QN(n1954) );
  FD1 \gpr_reg[29][21]  ( .D(n233), .CP(clk), .Q(\gpr[29][21] ), .QN(n1953) );
  FD1 \gpr_reg[29][20]  ( .D(n232), .CP(clk), .Q(\gpr[29][20] ), .QN(n1952) );
  FD1 \gpr_reg[29][19]  ( .D(n231), .CP(clk), .Q(\gpr[29][19] ), .QN(n1951) );
  FD1 \gpr_reg[29][18]  ( .D(n230), .CP(clk), .Q(\gpr[29][18] ), .QN(n1950) );
  FD1 \gpr_reg[29][17]  ( .D(n229), .CP(clk), .Q(\gpr[29][17] ), .QN(n1949) );
  FD1 \gpr_reg[29][16]  ( .D(n228), .CP(clk), .Q(\gpr[29][16] ), .QN(n1948) );
  FD1 \gpr_reg[29][15]  ( .D(n227), .CP(clk), .Q(\gpr[29][15] ), .QN(n1947) );
  FD1 \gpr_reg[29][14]  ( .D(n226), .CP(clk), .Q(\gpr[29][14] ), .QN(n1946) );
  FD1 \gpr_reg[29][13]  ( .D(n225), .CP(clk), .Q(\gpr[29][13] ), .QN(n1945) );
  FD1 \gpr_reg[29][12]  ( .D(n224), .CP(clk), .Q(\gpr[29][12] ), .QN(n1944) );
  FD1 \gpr_reg[29][11]  ( .D(n223), .CP(clk), .Q(\gpr[29][11] ), .QN(n1943) );
  FD1 \gpr_reg[29][10]  ( .D(n222), .CP(clk), .Q(\gpr[29][10] ), .QN(n1942) );
  FD1 \gpr_reg[29][9]  ( .D(n221), .CP(clk), .Q(\gpr[29][9] ), .QN(n1941) );
  FD1 \gpr_reg[29][8]  ( .D(n220), .CP(clk), .Q(\gpr[29][8] ), .QN(n1940) );
  FD1 \gpr_reg[29][7]  ( .D(n219), .CP(clk), .Q(\gpr[29][7] ), .QN(n1939) );
  FD1 \gpr_reg[29][6]  ( .D(n218), .CP(clk), .Q(\gpr[29][6] ), .QN(n1938) );
  FD1 \gpr_reg[29][5]  ( .D(n217), .CP(clk), .Q(\gpr[29][5] ), .QN(n1937) );
  FD1 \gpr_reg[29][4]  ( .D(n216), .CP(clk), .Q(\gpr[29][4] ), .QN(n1936) );
  FD1 \gpr_reg[29][3]  ( .D(n215), .CP(clk), .Q(\gpr[29][3] ), .QN(n1935) );
  FD1 \gpr_reg[29][2]  ( .D(n214), .CP(clk), .Q(\gpr[29][2] ), .QN(n1934) );
  FD1 \gpr_reg[29][1]  ( .D(n213), .CP(clk), .Q(\gpr[29][1] ), .QN(n1933) );
  FD1 \gpr_reg[29][0]  ( .D(n212), .CP(clk), .Q(\gpr[29][0] ), .QN(n1932) );
  FD1 \gpr_reg[30][31]  ( .D(n211), .CP(clk), .Q(\gpr[30][31] ), .QN(n1988) );
  FD1 \gpr_reg[30][30]  ( .D(n210), .CP(clk), .Q(\gpr[30][30] ), .QN(n1987) );
  FD1 \gpr_reg[30][29]  ( .D(n209), .CP(clk), .Q(\gpr[30][29] ), .QN(n1986) );
  FD1 \gpr_reg[30][28]  ( .D(n208), .CP(clk), .Q(\gpr[30][28] ), .QN(n1985) );
  FD1 \gpr_reg[30][27]  ( .D(n207), .CP(clk), .Q(\gpr[30][27] ), .QN(n1984) );
  FD1 \gpr_reg[30][26]  ( .D(n206), .CP(clk), .Q(\gpr[30][26] ), .QN(n1983) );
  FD1 \gpr_reg[30][25]  ( .D(n205), .CP(clk), .Q(\gpr[30][25] ), .QN(n1982) );
  FD1 \gpr_reg[30][24]  ( .D(n204), .CP(clk), .Q(\gpr[30][24] ), .QN(n1981) );
  FD1 \gpr_reg[30][23]  ( .D(n203), .CP(clk), .Q(\gpr[30][23] ), .QN(n1980) );
  FD1 \gpr_reg[30][22]  ( .D(n202), .CP(clk), .Q(\gpr[30][22] ), .QN(n1979) );
  FD1 \gpr_reg[30][21]  ( .D(n201), .CP(clk), .Q(\gpr[30][21] ), .QN(n1978) );
  FD1 \gpr_reg[30][20]  ( .D(n200), .CP(clk), .Q(\gpr[30][20] ), .QN(n1977) );
  FD1 \gpr_reg[30][19]  ( .D(n199), .CP(clk), .Q(\gpr[30][19] ), .QN(n1976) );
  FD1 \gpr_reg[30][18]  ( .D(n198), .CP(clk), .Q(\gpr[30][18] ), .QN(n1975) );
  FD1 \gpr_reg[30][17]  ( .D(n197), .CP(clk), .Q(\gpr[30][17] ), .QN(n1974) );
  FD1 \gpr_reg[30][16]  ( .D(n196), .CP(clk), .Q(\gpr[30][16] ), .QN(n1973) );
  FD1 \gpr_reg[30][15]  ( .D(n195), .CP(clk), .Q(\gpr[30][15] ), .QN(n1972) );
  FD1 \gpr_reg[30][13]  ( .D(n193), .CP(clk), .Q(\gpr[30][13] ), .QN(n1971) );
  FD1 \gpr_reg[30][12]  ( .D(n192), .CP(clk), .Q(\gpr[30][12] ), .QN(n1970) );
  FD1 \gpr_reg[30][11]  ( .D(n191), .CP(clk), .Q(\gpr[30][11] ), .QN(n1969) );
  FD1 \gpr_reg[30][10]  ( .D(n190), .CP(clk), .Q(\gpr[30][10] ), .QN(n1968) );
  FD1 \gpr_reg[30][8]  ( .D(n188), .CP(clk), .Q(\gpr[30][8] ), .QN(n1967) );
  FD1 \gpr_reg[30][6]  ( .D(n186), .CP(clk), .Q(\gpr[30][6] ), .QN(n1966) );
  FD1 \gpr_reg[30][5]  ( .D(n185), .CP(clk), .Q(\gpr[30][5] ), .QN(n1965) );
  FD1 \gpr_reg[30][3]  ( .D(n183), .CP(clk), .Q(\gpr[30][3] ), .QN(n1964) );
  FD1 \gpr_reg[30][2]  ( .D(n182), .CP(clk), .Q(\gpr[30][2] ), .QN(n137) );
  FD1 \gpr_reg[30][1]  ( .D(n181), .CP(clk), .Q(\gpr[30][1] ), .QN(n134) );
  FD1 \gpr_reg[30][0]  ( .D(n180), .CP(clk), .Q(\gpr[30][0] ), .QN(n131) );
  FD1 \gpr_reg[31][31]  ( .D(n179), .CP(clk), .Q(\gpr[31][31] ), .QN(n2017) );
  FD1 \gpr_reg[31][30]  ( .D(n178), .CP(clk), .Q(\gpr[31][30] ), .QN(n2016) );
  FD1 \gpr_reg[31][29]  ( .D(n177), .CP(clk), .Q(\gpr[31][29] ), .QN(n2015) );
  FD1 \gpr_reg[31][28]  ( .D(n176), .CP(clk), .Q(\gpr[31][28] ), .QN(n2014) );
  FD1 \gpr_reg[31][27]  ( .D(n175), .CP(clk), .Q(\gpr[31][27] ), .QN(n2013) );
  FD1 \gpr_reg[31][26]  ( .D(n174), .CP(clk), .Q(\gpr[31][26] ), .QN(n2012) );
  FD1 \gpr_reg[31][25]  ( .D(n173), .CP(clk), .Q(\gpr[31][25] ), .QN(n2011) );
  FD1 \gpr_reg[31][24]  ( .D(n172), .CP(clk), .Q(\gpr[31][24] ), .QN(n2010) );
  FD1 \gpr_reg[31][23]  ( .D(n171), .CP(clk), .Q(\gpr[31][23] ), .QN(n2009) );
  FD1 \gpr_reg[31][22]  ( .D(n170), .CP(clk), .Q(\gpr[31][22] ), .QN(n2008) );
  FD1 \gpr_reg[31][21]  ( .D(n169), .CP(clk), .Q(\gpr[31][21] ), .QN(n2007) );
  FD1 \gpr_reg[31][20]  ( .D(n168), .CP(clk), .Q(\gpr[31][20] ), .QN(n2006) );
  FD1 \gpr_reg[31][19]  ( .D(n167), .CP(clk), .Q(\gpr[31][19] ), .QN(n2005) );
  FD1 \gpr_reg[31][18]  ( .D(n166), .CP(clk), .Q(\gpr[31][18] ), .QN(n2004) );
  FD1 \gpr_reg[31][17]  ( .D(n165), .CP(clk), .Q(\gpr[31][17] ), .QN(n2003) );
  FD1 \gpr_reg[31][16]  ( .D(n164), .CP(clk), .Q(\gpr[31][16] ), .QN(n2002) );
  FD1 \gpr_reg[31][15]  ( .D(n163), .CP(clk), .Q(\gpr[31][15] ), .QN(n2001) );
  FD1 \gpr_reg[31][14]  ( .D(n162), .CP(clk), .Q(\gpr[31][14] ), .QN(n2000) );
  FD1 \gpr_reg[31][13]  ( .D(n161), .CP(clk), .Q(\gpr[31][13] ), .QN(n1999) );
  FD1 \gpr_reg[31][12]  ( .D(n160), .CP(clk), .Q(\gpr[31][12] ), .QN(n1998) );
  FD1 \gpr_reg[31][11]  ( .D(n159), .CP(clk), .Q(\gpr[31][11] ), .QN(n1997) );
  FD1 \gpr_reg[31][10]  ( .D(n158), .CP(clk), .Q(\gpr[31][10] ), .QN(n1996) );
  FD1 \gpr_reg[31][9]  ( .D(n157), .CP(clk), .Q(\gpr[31][9] ), .QN(n1995) );
  FD1 \gpr_reg[31][8]  ( .D(n156), .CP(clk), .Q(\gpr[31][8] ), .QN(n1994) );
  FD1 \gpr_reg[31][7]  ( .D(n155), .CP(clk), .Q(\gpr[31][7] ), .QN(n1993) );
  FD1 \gpr_reg[31][6]  ( .D(n154), .CP(clk), .Q(\gpr[31][6] ), .QN(n1992) );
  FD1 \gpr_reg[31][5]  ( .D(n153), .CP(clk), .Q(\gpr[31][5] ), .QN(n1991) );
  FD1 \gpr_reg[31][4]  ( .D(n152), .CP(clk), .Q(\gpr[31][4] ), .QN(n1990) );
  FD1 \gpr_reg[31][3]  ( .D(n151), .CP(clk), .Q(\gpr[31][3] ), .QN(n1989) );
  FD1 \gpr_reg[31][2]  ( .D(n150), .CP(clk), .Q(\gpr[31][2] ), .QN(n68) );
  FD1 \gpr_reg[31][1]  ( .D(n149), .CP(clk), .Q(\gpr[31][1] ), .QN(n65) );
  FD1 \gpr_reg[31][0]  ( .D(n148), .CP(clk), .Q(\gpr[31][0] ), .QN(n62) );
  FD1 \gpr_reg[1][6]  ( .D(n1114), .CP(clk), .Q(\gpr[1][6] ), .QN(n3217) );
  FD1 \gpr_reg[1][4]  ( .D(n1112), .CP(clk), .Q(\gpr[1][4] ), .QN(n3216) );
  FD1 \gpr_reg[8][6]  ( .D(n890), .CP(clk), .Q(\gpr[8][6] ), .QN(n3225) );
  FD1 \gpr_reg[15][6]  ( .D(n666), .CP(clk), .Q(\gpr[15][6] ), .QN(n3247) );
  FD1 \gpr_reg[14][6]  ( .D(n698), .CP(clk), .Q(\gpr[14][6] ), .QN(n3245) );
  FD1 \gpr_reg[13][6]  ( .D(n730), .CP(clk), .Q(\gpr[13][6] ), .QN(n3242) );
  FD1 \gpr_reg[12][6]  ( .D(n762), .CP(clk), .Q(\gpr[12][6] ), .QN(n3239) );
  FD1 \gpr_reg[11][6]  ( .D(n794), .CP(clk), .Q(\gpr[11][6] ), .QN(n3236) );
  FD1 \gpr_reg[10][6]  ( .D(n826), .CP(clk), .Q(\gpr[10][6] ), .QN(n3233) );
  FD1 \gpr_reg[9][6]  ( .D(n858), .CP(clk), .Q(\gpr[9][6] ), .QN(n3229) );
  FD1 \gpr_reg[9][4]  ( .D(n856), .CP(clk), .Q(\gpr[9][4] ), .QN(n3227) );
  FD1 \gpr_reg[9][5]  ( .D(n857), .CP(clk), .Q(\gpr[9][5] ), .QN(n3228) );
  FD1 \gpr_reg[9][9]  ( .D(n861), .CP(clk), .Q(\gpr[9][9] ), .QN(n3230) );
  FD1 \gpr_reg[17][9]  ( .D(n605), .CP(clk), .Q(\gpr[17][9] ), .QN(n3250) );
  FD1 \gpr_reg[20][4]  ( .D(n504), .CP(clk), .Q(\gpr[20][4] ), .QN(n3254) );
  FD1 \gpr_reg[25][5]  ( .D(n345), .CP(clk), .Q(\gpr[25][5] ), .QN(n3261) );
  FD1 \gpr_reg[25][9]  ( .D(n349), .CP(clk), .Q(\gpr[25][9] ), .QN(n3262) );
  FD1 \gpr_reg[28][14]  ( .D(n258), .CP(clk), .Q(\gpr[28][14] ), .QN(n3267) );
  FD1 \gpr_reg[30][4]  ( .D(n184), .CP(clk), .Q(\gpr[30][4] ), .QN(n3270) );
  FD1 \gpr_reg[30][7]  ( .D(n187), .CP(clk), .Q(\gpr[30][7] ), .QN(n3271) );
  FD1 \gpr_reg[30][9]  ( .D(n189), .CP(clk), .Q(\gpr[30][9] ), .QN(n3272) );
  FD1 \gpr_reg[30][14]  ( .D(n194), .CP(clk), .Q(\gpr[30][14] ), .QN(n3273) );
  FD1 \gpr_reg[23][2]  ( .D(n406), .CP(clk), .Q(\gpr[23][2] ), .QN(n3259) );
  FD1 \gpr_reg[22][2]  ( .D(n438), .CP(clk), .Q(\gpr[22][2] ), .QN(n3257) );
  FD1 \gpr_reg[26][2]  ( .D(n310), .CP(clk), .Q(\gpr[26][2] ), .QN(n3264) );
  B5IP U4 ( .A(n2081), .Z(n3161) );
  IVI U5 ( .A(n2092), .Z(n34) );
  IVI U6 ( .A(n3264), .Z(n33) );
  IVI U7 ( .A(n3257), .Z(n35) );
  ND4 U8 ( .A(n3637), .B(n3636), .C(n3635), .D(n2061), .Z(n3647) );
  ND4 U9 ( .A(n3520), .B(n3519), .C(n3518), .D(n2063), .Z(n3530) );
  AO4 U10 ( .A(n3341), .B(n4455), .C(n3340), .D(n4459), .Z(n3342) );
  IVI U11 ( .A(n3206), .Z(n3213) );
  B3IP U12 ( .A(n2026), .Z1(n1), .Z2(n2) );
  IVI U13 ( .A(n3214), .Z(n3208) );
  IVI U14 ( .A(n3214), .Z(n3209) );
  IVI U15 ( .A(n48), .Z(n3134) );
  IVDAP U16 ( .A(n2052), .Y(n2057), .Z(n2058) );
  B2IP U17 ( .A(n2995), .Z1(n20), .Z2(n21) );
  IVI U18 ( .A(n3214), .Z(n3210) );
  B2IP U19 ( .A(n2946), .Z1(n22), .Z2(n23) );
  B2IP U20 ( .A(n2947), .Z1(n24), .Z2(n25) );
  IVI U21 ( .A(n24), .Z(n2970) );
  ND2I U22 ( .A(n2064), .B(n26), .Z(n116) );
  AN2I U23 ( .A(n3392), .B(n3211), .Z(n26) );
  IVI U24 ( .A(n1), .Z(n27) );
  MUX21LP U25 ( .A(n3394), .B(n3393), .S(n2072), .Z(n3395) );
  MUX21LP U26 ( .A(n3432), .B(n3431), .S(n2072), .Z(n3433) );
  MUX21LP U27 ( .A(n3438), .B(n3437), .S(n2072), .Z(n3439) );
  MUX21LP U28 ( .A(n3435), .B(n3434), .S(n2072), .Z(n3436) );
  B5IP U29 ( .A(n2070), .Z(n2072) );
  MUX31LP U30 ( .D0(\gpr[13][2] ), .D1(\gpr[12][2] ), .D2(n3338), .A(n2027), 
        .B(n2), .Z(n3341) );
  AN2I U31 ( .A(n2093), .B(n3335), .Z(n28) );
  AN2I U32 ( .A(n2079), .B(n3334), .Z(n29) );
  NR2I U33 ( .A(n28), .B(n29), .Z(n3336) );
  IVI U34 ( .A(n3282), .Z(n2093) );
  IVI U35 ( .A(n3421), .Z(n30) );
  ND2I U36 ( .A(n31), .B(n32), .Z(n2024) );
  AN4 U37 ( .A(n3408), .B(n3407), .C(n3406), .D(n2059), .Z(n31) );
  NR2I U38 ( .A(n3417), .B(n30), .Z(n32) );
  MUX21L U39 ( .A(n33), .B(n34), .S(n3148), .Z(n3333) );
  MUX21L U40 ( .A(n35), .B(\gpr[23][2] ), .S(n2031), .Z(n3332) );
  MUX31LP U41 ( .D0(n127), .D1(n58), .D2(n3333), .A(n2043), .B(n27), .Z(n3334)
         );
  IVI U42 ( .A(N14), .Z(n36) );
  IVI U43 ( .A(N14), .Z(n37) );
  IVI U44 ( .A(N14), .Z(n3202) );
  IVI U45 ( .A(n3203), .Z(n2070) );
  B5I U46 ( .A(n3203), .Z(n3201) );
  MUX21L U47 ( .A(n3398), .B(n3397), .S(n3194), .Z(n3399) );
  MUX21L U48 ( .A(n3552), .B(n3551), .S(n3192), .Z(n3553) );
  MUX21L U49 ( .A(n4403), .B(n4402), .S(n3195), .Z(n4404) );
  ND4 U50 ( .A(n3831), .B(n3830), .C(n3829), .D(n2059), .Z(n3841) );
  IVI U51 ( .A(n3212), .Z(n3211) );
  B2IP U52 ( .A(n2980), .Z1(n38), .Z2(n39) );
  IVDAP U53 ( .A(n2945), .Y(n40), .Z(n41) );
  B2IP U54 ( .A(n2995), .Z1(n42), .Z2(n43) );
  B2IP U55 ( .A(n2980), .Z1(n44), .Z2(n45) );
  B2IP U56 ( .A(n2947), .Z1(n46), .Z2(n47) );
  AN2I U57 ( .A(n3276), .B(n3275), .Z(n48) );
  AN2I U58 ( .A(n2106), .B(n1179), .Z(n49) );
  B2IP U59 ( .A(n40), .Z1(n50), .Z2(n51) );
  B2IP U60 ( .A(N21), .Z1(n52), .Z2(n53) );
  B2IP U61 ( .A(n2102), .Z1(n73), .Z2(n74) );
  B2IP U62 ( .A(n49), .Z1(n75), .Z2(n76) );
  ND2P U63 ( .A(n3220), .B(n1179), .Z(n92) );
  ND2I U64 ( .A(n2103), .B(n1177), .Z(n93) );
  ND2I U65 ( .A(n1177), .B(n2105), .Z(n94) );
  AN2I U66 ( .A(N17), .B(N16), .Z(n115) );
  AN2I U67 ( .A(n4248), .B(n2062), .Z(n117) );
  OR2I U68 ( .A(n2065), .B(n3777), .Z(n118) );
  IVI U69 ( .A(N18), .Z(n2945) );
  B2IP U70 ( .A(n2995), .Z1(n119), .Z2(n120) );
  B2IP U71 ( .A(N22), .Z1(n121), .Z2(n122) );
  ND2I U72 ( .A(n3220), .B(n2112), .Z(n1153) );
  ND2I U73 ( .A(n3220), .B(n2109), .Z(n1154) );
  ND2I U74 ( .A(n3220), .B(n2111), .Z(n1155) );
  ND2I U75 ( .A(n3220), .B(n2108), .Z(n1156) );
  ND2I U76 ( .A(n3220), .B(n2110), .Z(n1157) );
  ND2I U77 ( .A(n3220), .B(n2104), .Z(n1158) );
  AN3P U78 ( .A(n3224), .B(n3223), .C(n3222), .Z(n1177) );
  AN2I U79 ( .A(wr_addr[0]), .B(n3219), .Z(n1179) );
  IVI U80 ( .A(n2029), .Z(n2018) );
  IVI U81 ( .A(n2018), .Z(n2019) );
  B4I U82 ( .A(n2039), .Z(n3170) );
  MUX31LP U83 ( .D0(n126), .D1(n57), .D2(n3310), .A(n2019), .B(n2083), .Z(
        n3311) );
  B4IP U84 ( .A(n3185), .Z(n3178) );
  B5IP U85 ( .A(n2044), .Z(n3167) );
  B4IP U86 ( .A(n37), .Z(n3191) );
  IVI U87 ( .A(n3152), .Z(n2020) );
  MUX21L U88 ( .A(n3821), .B(n3820), .S(n2), .Z(n3822) );
  B4IP U89 ( .A(n3201), .Z(n3196) );
  B5IP U90 ( .A(n3187), .Z(n3157) );
  B5IP U91 ( .A(n3186), .Z(n3166) );
  IVI U92 ( .A(n3182), .Z(n3181) );
  IVI U93 ( .A(n3182), .Z(n3168) );
  B4IP U94 ( .A(n2085), .Z(n3179) );
  IVI U95 ( .A(n2091), .Z(n2021) );
  B4IP U96 ( .A(n2082), .Z(n3162) );
  IVI U97 ( .A(n2084), .Z(n2048) );
  B4I U98 ( .A(n2084), .Z(n3171) );
  B4IP U99 ( .A(n3188), .Z(n3155) );
  MUX31LP U100 ( .D0(n77), .D1(n143), .D2(n3277), .A(n3167), .B(n3197), .Z(
        n3278) );
  B4IP U101 ( .A(n2044), .Z(n3169) );
  MUX21LP U102 ( .A(n4008), .B(n4007), .S(n3199), .Z(n4009) );
  B5IP U103 ( .A(n36), .Z(n3197) );
  ND4P U104 ( .A(n3870), .B(n3869), .C(n3868), .D(n2065), .Z(n3880) );
  IVI U105 ( .A(n3202), .Z(n3194) );
  MUX21LP U106 ( .A(n3594), .B(n3593), .S(n3192), .Z(n3595) );
  MUX21LP U107 ( .A(n3591), .B(n3590), .S(n3192), .Z(n3592) );
  MUX21LP U108 ( .A(n3588), .B(n3587), .S(n3192), .Z(n3589) );
  IVI U109 ( .A(n3284), .Z(n2022) );
  IVI U110 ( .A(n3284), .Z(n2074) );
  ND4P U111 ( .A(n4143), .B(n4142), .C(n4141), .D(n2057), .Z(n4153) );
  B4I U112 ( .A(n3189), .Z(n2034) );
  ND4P U113 ( .A(n4221), .B(n4220), .C(n4219), .D(n2061), .Z(n4231) );
  ND4P U114 ( .A(n4335), .B(n4334), .C(n4333), .D(n2059), .Z(n4345) );
  MUX21L U115 ( .A(n4364), .B(n4363), .S(n3196), .Z(n4365) );
  MUX21L U116 ( .A(n4367), .B(n4366), .S(n3196), .Z(n4368) );
  MUX21L U117 ( .A(n4370), .B(n4369), .S(n3196), .Z(n4371) );
  IVI U118 ( .A(n3152), .Z(n2023) );
  B4IP U119 ( .A(n2087), .Z(n3174) );
  MUX31LP U120 ( .D0(n61), .D1(n130), .D2(n3330), .A(n2041), .B(n3198), .Z(
        n3344) );
  AN2I U121 ( .A(n2024), .B(n2025), .Z(rd_data1[4]) );
  AN2I U122 ( .A(n116), .B(n3422), .Z(n2025) );
  IVI U123 ( .A(n36), .Z(n2026) );
  B4IP U124 ( .A(n2030), .Z(n3195) );
  IVI U125 ( .A(n2037), .Z(n2027) );
  IVI U126 ( .A(n2020), .Z(n2028) );
  IVI U127 ( .A(n3149), .Z(n2029) );
  AO4P U128 ( .A(n3295), .B(n4455), .C(n3294), .D(n4459), .Z(n3296) );
  MUX21LP U129 ( .A(n4133), .B(n4132), .S(n3191), .Z(n4134) );
  ND4P U130 ( .A(n3754), .B(n3753), .C(n3752), .D(n2057), .Z(n3764) );
  IVI U131 ( .A(n3151), .Z(n2031) );
  ND4P U132 ( .A(n4182), .B(n4181), .C(n4180), .D(n2055), .Z(n4192) );
  B5IP U133 ( .A(n3202), .Z(n3192) );
  MUX21LP U134 ( .A(n3891), .B(n3890), .S(n3200), .Z(n3892) );
  MUX21LP U135 ( .A(n3930), .B(n3929), .S(n3200), .Z(n3931) );
  MUX21LP U136 ( .A(n3882), .B(n3881), .S(n3200), .Z(n3883) );
  MUX21LP U137 ( .A(n3934), .B(n3933), .S(n3200), .Z(n3935) );
  MUX21LP U138 ( .A(n3852), .B(n3851), .S(n3200), .Z(n3853) );
  MUX21LP U139 ( .A(n3856), .B(n3855), .S(n3200), .Z(n3857) );
  MUX21LP U140 ( .A(n3875), .B(n3874), .S(n3200), .Z(n3876) );
  MUX21LP U141 ( .A(n3872), .B(n3871), .S(n3200), .Z(n3873) );
  MUX21LP U142 ( .A(n3006), .B(n3283), .S(n2083), .Z(n3287) );
  B4IP U143 ( .A(n3183), .Z(n3176) );
  MUX31LP U144 ( .D0(\gpr[29][2] ), .D1(\gpr[28][2] ), .D2(n3331), .A(n2067), 
        .B(n3197), .Z(n3337) );
  B5IP U145 ( .A(n3186), .Z(n3164) );
  ND4P U146 ( .A(n4258), .B(n4259), .C(n4260), .D(n4451), .Z(n4270) );
  AO1P U147 ( .A(n4274), .B(n4275), .C(n117), .D(n4276), .Z(rd_data1[26]) );
  ND2I U148 ( .A(n2032), .B(n118), .Z(n2033) );
  IVI U149 ( .A(n3811), .Z(n2032) );
  IVI U150 ( .A(n2033), .Z(rd_data1[14]) );
  B4IP U151 ( .A(n2028), .Z(n3165) );
  IVI U152 ( .A(n2039), .Z(n2035) );
  IVI U153 ( .A(n2091), .Z(n3172) );
  IVI U154 ( .A(n3184), .Z(n2036) );
  IVI U155 ( .A(n2091), .Z(n2037) );
  IVI U156 ( .A(n2029), .Z(n2038) );
  IVI U157 ( .A(n2020), .Z(n2039) );
  IVI U158 ( .A(n2023), .Z(n2091) );
  IVI U159 ( .A(n2100), .Z(n2040) );
  IVI U160 ( .A(n2020), .Z(n2100) );
  IVI U161 ( .A(n3189), .Z(n2041) );
  IVI U162 ( .A(n3150), .Z(n2042) );
  IVI U163 ( .A(n2070), .Z(n2049) );
  IVI U164 ( .A(n3150), .Z(n2043) );
  IVI U165 ( .A(n3150), .Z(n2044) );
  B4IP U166 ( .A(n2067), .Z(n3158) );
  ND2I U167 ( .A(n115), .B(n3213), .Z(n2045) );
  ND2I U168 ( .A(n115), .B(n3213), .Z(n2046) );
  ND2I U169 ( .A(n3205), .B(n3293), .Z(n2047) );
  AO4P U170 ( .A(n3318), .B(n4455), .C(n3317), .D(n4459), .Z(n3319) );
  IVI U171 ( .A(n3202), .Z(n2050) );
  B3IP U172 ( .A(n3190), .Z1(n2030), .Z2(n2083) );
  IVI U173 ( .A(n4451), .Z(n2051) );
  IVI U174 ( .A(n4451), .Z(n2052) );
  IVI U175 ( .A(n4451), .Z(n2053) );
  IVI U176 ( .A(n4451), .Z(n2054) );
  B3IP U177 ( .A(n2051), .Z1(n2055), .Z2(n2056) );
  B3IP U178 ( .A(n2052), .Z1(n2059), .Z2(n2060) );
  B3IP U179 ( .A(n2053), .Z1(n2061), .Z2(n2062) );
  B3IP U180 ( .A(n2054), .Z1(n2063), .Z2(n2064) );
  B3IP U181 ( .A(n2054), .Z1(n2065), .Z2(n2066) );
  IVI U182 ( .A(n2023), .Z(n2067) );
  B4IP U183 ( .A(n2090), .Z(n3177) );
  IVI U184 ( .A(n2029), .Z(n2068) );
  ND2I U185 ( .A(n115), .B(n3205), .Z(n4447) );
  IVI U186 ( .A(n3148), .Z(n2069) );
  IVI U187 ( .A(n2043), .Z(n2071) );
  IVI U188 ( .A(n3203), .Z(n2073) );
  OR2P U189 ( .A(n3207), .B(N17), .Z(n4455) );
  IVI U190 ( .A(n2046), .Z(n2075) );
  IVI U191 ( .A(n2045), .Z(n2076) );
  IVI U192 ( .A(n2046), .Z(n2077) );
  IVI U193 ( .A(n2045), .Z(n2078) );
  IVI U194 ( .A(n2046), .Z(n2079) );
  IVI U195 ( .A(n2045), .Z(n2080) );
  IVI U196 ( .A(n2031), .Z(n2081) );
  IVI U197 ( .A(n2031), .Z(n2082) );
  IVI U198 ( .A(n3204), .Z(n3190) );
  IVI U199 ( .A(n2089), .Z(n2084) );
  IVI U200 ( .A(n3149), .Z(n2085) );
  IVI U201 ( .A(n3148), .Z(n2086) );
  IVI U202 ( .A(n2023), .Z(n2087) );
  B4I U203 ( .A(n3184), .Z(n2088) );
  MUX31LP U204 ( .D0(\gpr[16][2] ), .D1(\gpr[17][2] ), .D2(n3339), .A(n2021), 
        .B(n3191), .Z(n3340) );
  B5IP U205 ( .A(n2069), .Z(n3159) );
  MUX31LP U206 ( .D0(\gpr[16][0] ), .D1(\gpr[17][0] ), .D2(n3292), .A(n3158), 
        .B(n2050), .Z(n3294) );
  IVI U207 ( .A(n3151), .Z(n2089) );
  ND4P U208 ( .A(n3676), .B(n3675), .C(n3674), .D(n2065), .Z(n3686) );
  MUX21LP U209 ( .A(n3833), .B(n3832), .S(n3192), .Z(n3834) );
  B4IP U210 ( .A(n2042), .Z(n3153) );
  ND4P U211 ( .A(n4104), .B(n4103), .C(n4102), .D(n2061), .Z(n4114) );
  IVI U212 ( .A(n4447), .Z(n3135) );
  ND4P U213 ( .A(n4374), .B(n4373), .C(n4372), .D(n2063), .Z(n4384) );
  IVI U214 ( .A(n2020), .Z(n2090) );
  ND4P U215 ( .A(n4454), .B(n4453), .C(n4452), .D(n2061), .Z(n4466) );
  MUX31LP U216 ( .D0(\gpr[16][1] ), .D1(\gpr[17][1] ), .D2(n3316), .A(n2068), 
        .B(n3192), .Z(n3317) );
  IVI U217 ( .A(n2047), .Z(n2094) );
  IVI U218 ( .A(n3282), .Z(n2095) );
  IVI U219 ( .A(n2047), .Z(n2096) );
  IVI U220 ( .A(n2047), .Z(n2097) );
  IVI U221 ( .A(n3282), .Z(n2098) );
  IVI U222 ( .A(n3282), .Z(n2099) );
  ND4P U223 ( .A(n4413), .B(n4412), .C(n4411), .D(n2061), .Z(n4423) );
  B4IP U224 ( .A(n2100), .Z(n2101) );
  IVI U225 ( .A(n3152), .Z(n3149) );
  AO3P U226 ( .A(n3314), .B(n4447), .C(n2055), .D(n3313), .Z(n3320) );
  MUX21LP U227 ( .A(n3363), .B(n3362), .S(n2072), .Z(n3364) );
  AO2P U228 ( .A(n2094), .B(n3287), .C(n2078), .D(n3286), .Z(n3288) );
  AO3P U229 ( .A(n3289), .B(n4447), .C(n2061), .D(n3288), .Z(n3297) );
  AO2P U230 ( .A(n2095), .B(n3312), .C(n2080), .D(n3311), .Z(n3313) );
  AO3P U231 ( .A(n3337), .B(n4447), .C(n2055), .D(n3336), .Z(n3343) );
  MUX31LP U232 ( .D0(n78), .D1(n144), .D2(n3305), .A(n3174), .B(n3192), .Z(
        n3306) );
  MUX31LP U233 ( .D0(n79), .D1(n145), .D2(n3280), .A(n2088), .B(n3191), .Z(
        n3298) );
  MUX31LP U234 ( .D0(n80), .D1(n146), .D2(n3307), .A(n3159), .B(n3198), .Z(
        n3321) );
  MUX31LP U235 ( .D0(\gpr[12][1] ), .D1(\gpr[13][1] ), .D2(n3315), .A(n3173), 
        .B(n2049), .Z(n3318) );
  MUX31LP U236 ( .D0(\gpr[12][0] ), .D1(\gpr[13][0] ), .D2(n3290), .A(n2041), 
        .B(n2050), .Z(n3295) );
  MUX31LP U237 ( .D0(\gpr[28][1] ), .D1(\gpr[29][1] ), .D2(n3308), .A(n3164), 
        .B(n3193), .Z(n3314) );
  MUX31LP U238 ( .D0(\gpr[28][0] ), .D1(\gpr[29][0] ), .D2(n3281), .A(n2068), 
        .B(n2), .Z(n3289) );
  MUX31LP U239 ( .D0(n56), .D1(n125), .D2(n3285), .A(n3172), .B(n2083), .Z(
        n3286) );
  MUX31LP U240 ( .D0(n54), .D1(n123), .D2(n3309), .A(n2037), .B(n3194), .Z(
        n3312) );
  AN3P U241 ( .A(wr_addr[3]), .B(RegWrite), .C(n3221), .Z(n2106) );
  IVAP U242 ( .A(n50), .Z(n2953) );
  B5IP U243 ( .A(n20), .Z(n2999) );
  IVI U244 ( .A(n2948), .Z(n2977) );
  MUX31LP U245 ( .D0(n55), .D1(n124), .D2(n3332), .A(n3172), .B(n3194), .Z(
        n3335) );
  IVAP U246 ( .A(n2948), .Z(n2979) );
  IVAP U247 ( .A(n2950), .Z(n2963) );
  IVI U248 ( .A(n2951), .Z(n2956) );
  IVI U249 ( .A(n2948), .Z(n2978) );
  IVI U250 ( .A(n2949), .Z(n2967) );
  IVI U251 ( .A(n41), .Z(n2976) );
  IVI U252 ( .A(n41), .Z(n2973) );
  IVI U253 ( .A(n41), .Z(n2959) );
  ND4 U254 ( .A(n3559), .B(n3558), .C(n3557), .D(n2065), .Z(n3569) );
  ND4 U255 ( .A(n4026), .B(n4025), .C(n4024), .D(n2055), .Z(n4036) );
  ND4 U256 ( .A(n4065), .B(n4064), .C(n4063), .D(n2055), .Z(n4075) );
  ND4 U257 ( .A(n3987), .B(n3986), .C(n3985), .D(n2063), .Z(n3997) );
  ND4 U258 ( .A(n3948), .B(n3947), .C(n3946), .D(n2055), .Z(n3958) );
  ND4 U259 ( .A(n3909), .B(n3908), .C(n3907), .D(n2061), .Z(n3919) );
  B4IP U260 ( .A(n2086), .Z(n3173) );
  IVI U261 ( .A(n41), .Z(n2958) );
  IVI U262 ( .A(n41), .Z(n2957) );
  IVI U263 ( .A(n2951), .Z(n2954) );
  IVI U264 ( .A(n2949), .Z(n2965) );
  IVI U265 ( .A(n2950), .Z(n2962) );
  IVI U266 ( .A(n41), .Z(n2975) );
  IVI U267 ( .A(n2949), .Z(n2974) );
  IVI U268 ( .A(n41), .Z(n2972) );
  IVI U269 ( .A(n2949), .Z(n2966) );
  IVI U270 ( .A(n2950), .Z(n2964) );
  IVI U271 ( .A(n41), .Z(n2971) );
  IVI U272 ( .A(n2951), .Z(n2955) );
  B4IP U273 ( .A(n44), .Z(n2987) );
  IVI U274 ( .A(n119), .Z(n2996) );
  IVI U275 ( .A(n3256), .Z(n3063) );
  IVI U276 ( .A(n3256), .Z(n3062) );
  IVI U277 ( .A(n93), .Z(n3045) );
  IVI U278 ( .A(n93), .Z(n3044) );
  IVI U279 ( .A(n3274), .Z(n3131) );
  IVI U280 ( .A(n3274), .Z(n3130) );
  IVI U281 ( .A(n3269), .Z(n3087) );
  IVI U282 ( .A(n3269), .Z(n3086) );
  IVI U283 ( .A(n3268), .Z(n3084) );
  IVI U284 ( .A(n3268), .Z(n3083) );
  IVI U285 ( .A(n3266), .Z(n3081) );
  IVI U286 ( .A(n3266), .Z(n3080) );
  IVI U287 ( .A(n3265), .Z(n3078) );
  IVI U288 ( .A(n3265), .Z(n3077) );
  IVI U289 ( .A(n3263), .Z(n3075) );
  IVI U290 ( .A(n3263), .Z(n3074) );
  IVI U291 ( .A(n3260), .Z(n3072) );
  IVI U292 ( .A(n3260), .Z(n3071) );
  IVI U293 ( .A(n94), .Z(n3069) );
  IVI U294 ( .A(n94), .Z(n3068) );
  IVI U295 ( .A(n3258), .Z(n3066) );
  IVI U296 ( .A(n3258), .Z(n3065) );
  IVI U297 ( .A(n3255), .Z(n3060) );
  IVI U298 ( .A(n3255), .Z(n3059) );
  IVI U299 ( .A(n3253), .Z(n3057) );
  IVI U300 ( .A(n3253), .Z(n3056) );
  IVI U301 ( .A(n3252), .Z(n3054) );
  IVI U302 ( .A(n3252), .Z(n3053) );
  IVI U303 ( .A(n3251), .Z(n3051) );
  IVI U304 ( .A(n3251), .Z(n3050) );
  IVI U305 ( .A(n3249), .Z(n3048) );
  IVI U306 ( .A(n3249), .Z(n3047) );
  IVI U307 ( .A(n92), .Z(n3026) );
  IVI U308 ( .A(n92), .Z(n3025) );
  IVI U309 ( .A(n1158), .Z(n3023) );
  IVI U310 ( .A(n1158), .Z(n3022) );
  IVI U311 ( .A(n1157), .Z(n3020) );
  IVI U312 ( .A(n1157), .Z(n3019) );
  IVI U313 ( .A(n1156), .Z(n3017) );
  IVI U314 ( .A(n1156), .Z(n3016) );
  IVI U315 ( .A(n1155), .Z(n3014) );
  IVI U316 ( .A(n1155), .Z(n3013) );
  IVI U317 ( .A(n1154), .Z(n3011) );
  IVI U318 ( .A(n1154), .Z(n3010) );
  IVI U319 ( .A(n1153), .Z(n3008) );
  IVI U320 ( .A(n1153), .Z(n3007) );
  ND4P U321 ( .A(n3370), .B(n3369), .C(n3368), .D(n2061), .Z(n3380) );
  ND4P U322 ( .A(n3481), .B(n3480), .C(n3479), .D(n2063), .Z(n3491) );
  ND4P U323 ( .A(n3793), .B(n3792), .C(n3791), .D(n2057), .Z(n3803) );
  ND4P U324 ( .A(n3442), .B(n3441), .C(n3440), .D(n2065), .Z(n3452) );
  ND4P U325 ( .A(n3598), .B(n3597), .C(n3596), .D(n2059), .Z(n3608) );
  MUX31LP U326 ( .D0(n2115), .D1(n2116), .D2(n2117), .A(n2983), .B(n21), .Z(
        n2114) );
  MUX21LP U327 ( .A(n2119), .B(n2120), .S(n2983), .Z(n2118) );
  MUX31LP U328 ( .D0(n2271), .D1(n2272), .D2(n2273), .A(n2985), .B(n21), .Z(
        n2270) );
  MUX21LP U329 ( .A(n2275), .B(n2276), .S(n2986), .Z(n2274) );
  MUX31LP U330 ( .D0(n2479), .D1(n2480), .D2(n2481), .A(n39), .B(n2999), .Z(
        n2478) );
  MUX21LP U331 ( .A(n2483), .B(n2484), .S(n45), .Z(n2482) );
  MUX31LP U332 ( .D0(n2713), .D1(n2714), .D2(n2715), .A(n2990), .B(n2999), .Z(
        n2712) );
  MUX21LP U333 ( .A(n2717), .B(n2718), .S(n2990), .Z(n2716) );
  MUX31LP U334 ( .D0(n2921), .D1(n2922), .D2(n2923), .A(n2991), .B(n2997), .Z(
        n2920) );
  MUX31LP U335 ( .D0(n2895), .D1(n2896), .D2(n2897), .A(n2983), .B(n120), .Z(
        n2894) );
  MUX21LP U336 ( .A(n2899), .B(n2900), .S(n2983), .Z(n2898) );
  MUX31LP U337 ( .D0(n2869), .D1(n2870), .D2(n2871), .A(n39), .B(n2997), .Z(
        n2868) );
  MUX21LP U338 ( .A(n2873), .B(n2874), .S(n2983), .Z(n2872) );
  IVI U339 ( .A(wr_data[0]), .Z(n3089) );
  IVI U340 ( .A(wr_data[1]), .Z(n3091) );
  IVI U341 ( .A(wr_data[2]), .Z(n3093) );
  IVI U342 ( .A(wr_data[3]), .Z(n3095) );
  IVI U343 ( .A(wr_data[0]), .Z(n3090) );
  IVI U344 ( .A(wr_data[1]), .Z(n3092) );
  IVI U345 ( .A(wr_data[2]), .Z(n3094) );
  IVI U346 ( .A(wr_data[3]), .Z(n3096) );
  MUX31LP U347 ( .D0(\gpr[28][10] ), .D1(\gpr[29][10] ), .D2(n2373), .A(n2956), 
        .B(n2992), .Z(n2377) );
  MUX31LP U348 ( .D0(\gpr[28][9] ), .D1(\gpr[29][9] ), .D2(n2347), .A(n2954), 
        .B(n2992), .Z(n2351) );
  MUX31LP U349 ( .D0(\gpr[28][6] ), .D1(\gpr[29][6] ), .D2(n2269), .A(n2967), 
        .B(n2992), .Z(n2273) );
  MUX31LP U350 ( .D0(\gpr[28][4] ), .D1(\gpr[29][4] ), .D2(n2217), .A(n2965), 
        .B(n2991), .Z(n2221) );
  MUX31LP U351 ( .D0(\gpr[28][2] ), .D1(\gpr[29][2] ), .D2(n2165), .A(n2963), 
        .B(n2991), .Z(n2169) );
  MUX31LP U352 ( .D0(\gpr[28][1] ), .D1(\gpr[29][1] ), .D2(n2139), .A(n2962), 
        .B(n2991), .Z(n2143) );
  MUX31LP U353 ( .D0(\gpr[28][12] ), .D1(\gpr[29][12] ), .D2(n2425), .A(n2958), 
        .B(n2992), .Z(n2429) );
  MUX31LP U354 ( .D0(\gpr[28][13] ), .D1(\gpr[29][13] ), .D2(n2451), .A(n2959), 
        .B(n2992), .Z(n2455) );
  MUX31LP U355 ( .D0(\gpr[28][21] ), .D1(\gpr[29][21] ), .D2(n2659), .A(n2977), 
        .B(n2993), .Z(n2663) );
  MUX31LP U356 ( .D0(\gpr[28][20] ), .D1(\gpr[29][20] ), .D2(n2633), .A(n2976), 
        .B(n2993), .Z(n2637) );
  MUX31LP U357 ( .D0(\gpr[28][22] ), .D1(\gpr[29][22] ), .D2(n2685), .A(n2978), 
        .B(n2993), .Z(n2689) );
  MUX31LP U358 ( .D0(\gpr[28][19] ), .D1(\gpr[29][19] ), .D2(n2607), .A(n2975), 
        .B(n2993), .Z(n2611) );
  MUX31LP U359 ( .D0(\gpr[28][18] ), .D1(\gpr[29][18] ), .D2(n2581), .A(n2974), 
        .B(n2992), .Z(n2585) );
  MUX31LP U360 ( .D0(\gpr[28][17] ), .D1(\gpr[29][17] ), .D2(n2555), .A(n2973), 
        .B(n2992), .Z(n2559) );
  MUX31LP U361 ( .D0(\gpr[28][16] ), .D1(\gpr[29][16] ), .D2(n2529), .A(n2972), 
        .B(n2992), .Z(n2533) );
  MUX31LP U362 ( .D0(\gpr[28][15] ), .D1(\gpr[29][15] ), .D2(n2503), .A(n2971), 
        .B(n2992), .Z(n2507) );
  MUX31LP U363 ( .D0(\gpr[28][11] ), .D1(\gpr[29][11] ), .D2(n2399), .A(n2957), 
        .B(n2992), .Z(n2403) );
  MUX31LP U364 ( .D0(\gpr[28][8] ), .D1(\gpr[29][8] ), .D2(n2321), .A(n2954), 
        .B(n2992), .Z(n2325) );
  MUX31LP U365 ( .D0(\gpr[28][7] ), .D1(\gpr[29][7] ), .D2(n2295), .A(n51), 
        .B(n2992), .Z(n2299) );
  MUX31LP U366 ( .D0(\gpr[28][5] ), .D1(\gpr[29][5] ), .D2(n2243), .A(n2966), 
        .B(n2991), .Z(n2247) );
  MUX31LP U367 ( .D0(\gpr[28][3] ), .D1(\gpr[29][3] ), .D2(n2191), .A(n2964), 
        .B(n2991), .Z(n2195) );
  B5IP U368 ( .A(n2069), .Z(n3156) );
  B5IP U369 ( .A(n2042), .Z(n3154) );
  B5IP U370 ( .A(n3187), .Z(n3160) );
  B5IP U371 ( .A(n2081), .Z(n3163) );
  B5IP U372 ( .A(n3183), .Z(n3175) );
  B5IP U373 ( .A(n3182), .Z(n3180) );
  B5IP U374 ( .A(n46), .Z(n2969) );
  B5IP U375 ( .A(n46), .Z(n2968) );
  B5IP U376 ( .A(n22), .Z(n2960) );
  B5IP U377 ( .A(n22), .Z(n2961) );
  B5IP U378 ( .A(n44), .Z(n2988) );
  B5IP U379 ( .A(n38), .Z(n2986) );
  B5IP U380 ( .A(n44), .Z(n2989) );
  IVI U381 ( .A(n2981), .Z(n2993) );
  IVI U382 ( .A(n2981), .Z(n2992) );
  IVI U383 ( .A(n50), .Z(n2952) );
  IVI U384 ( .A(n3149), .Z(n3189) );
  IVI U385 ( .A(n2089), .Z(n3184) );
  IVI U386 ( .A(n3279), .Z(n3146) );
  B5IP U387 ( .A(n52), .Z(n3001) );
  B5IP U388 ( .A(n52), .Z(n3003) );
  B5IP U389 ( .A(n52), .Z(n3002) );
  B5IP U390 ( .A(n75), .Z(n3042) );
  B5IP U391 ( .A(n3244), .Z(n3040) );
  B5IP U392 ( .A(n3241), .Z(n3038) );
  B5IP U393 ( .A(n3238), .Z(n3036) );
  B5IP U394 ( .A(n3235), .Z(n3034) );
  B5IP U395 ( .A(n3232), .Z(n3032) );
  B5IP U396 ( .A(n3226), .Z(n3030) );
  B5IP U397 ( .A(n73), .Z(n3028) );
  AN2I U398 ( .A(n2106), .B(n1177), .Z(n2102) );
  AN2I U399 ( .A(n2107), .B(n3248), .Z(n2103) );
  AN2I U400 ( .A(n3219), .B(n3222), .Z(n2104) );
  ND4 U401 ( .A(n4296), .B(n4295), .C(n4294), .D(n2055), .Z(n4306) );
  ND4 U402 ( .A(n3715), .B(n3714), .C(n3713), .D(n2063), .Z(n3725) );
  MUX31L U403 ( .D0(n2141), .D1(n2142), .D2(n2143), .A(n2984), .B(n21), .Z(
        n2140) );
  MUX31L U404 ( .D0(n2427), .D1(n2428), .D2(n2429), .A(n45), .B(n21), .Z(n2426) );
  MUX31L U405 ( .D0(n2453), .D1(n2454), .D2(n2455), .A(n45), .B(n2999), .Z(
        n2452) );
  MUX31L U406 ( .D0(n2661), .D1(n2662), .D2(n2663), .A(n45), .B(n2999), .Z(
        n2660) );
  MUX31L U407 ( .D0(n2635), .D1(n2636), .D2(n2637), .A(n45), .B(n2999), .Z(
        n2634) );
  MUX31L U408 ( .D0(n2401), .D1(n2402), .D2(n2403), .A(n2987), .B(n21), .Z(
        n2400) );
  MUX31L U409 ( .D0(n2375), .D1(n2376), .D2(n2377), .A(n2987), .B(n21), .Z(
        n2374) );
  MUX31L U410 ( .D0(n2557), .D1(n2558), .D2(n2559), .A(n2989), .B(n2999), .Z(
        n2556) );
  MUX31L U411 ( .D0(n2531), .D1(n2532), .D2(n2533), .A(n2988), .B(n2999), .Z(
        n2530) );
  MUX31L U412 ( .D0(n2583), .D1(n2584), .D2(n2585), .A(n2989), .B(n2999), .Z(
        n2582) );
  MUX31L U413 ( .D0(n2219), .D1(n2220), .D2(n2221), .A(n2985), .B(n21), .Z(
        n2218) );
  MUX31L U414 ( .D0(n2193), .D1(n2194), .D2(n2195), .A(n2984), .B(n21), .Z(
        n2192) );
  MUX31L U415 ( .D0(n2167), .D1(n2168), .D2(n2169), .A(n2984), .B(n21), .Z(
        n2166) );
  MUX31L U416 ( .D0(n2297), .D1(n2298), .D2(n2299), .A(n2986), .B(n21), .Z(
        n2296) );
  MUX31L U417 ( .D0(n2245), .D1(n2246), .D2(n2247), .A(n2985), .B(n21), .Z(
        n2244) );
  MUX31L U418 ( .D0(n2609), .D1(n2610), .D2(n2611), .A(n2989), .B(n2999), .Z(
        n2608) );
  MUX31L U419 ( .D0(n2505), .D1(n2506), .D2(n2507), .A(n2988), .B(n2999), .Z(
        n2504) );
  MUX31L U420 ( .D0(n2323), .D1(n2324), .D2(n2325), .A(n2986), .B(n21), .Z(
        n2322) );
  MUX31L U421 ( .D0(n2687), .D1(n2688), .D2(n2689), .A(n45), .B(n2999), .Z(
        n2686) );
  MUX31L U422 ( .D0(n2349), .D1(n2350), .D2(n2351), .A(n2987), .B(n21), .Z(
        n2348) );
  NR3 U423 ( .A(N20), .B(n2991), .C(n47), .Z(n3276) );
  AN2I U424 ( .A(wr_addr[3]), .B(n2107), .Z(n2105) );
  AN2I U425 ( .A(wr_addr[4]), .B(RegWrite), .Z(n2107) );
  AN3 U426 ( .A(wr_addr[2]), .B(n3224), .C(n3222), .Z(n2108) );
  AN3 U427 ( .A(wr_addr[1]), .B(n3223), .C(n3222), .Z(n2109) );
  AN3 U428 ( .A(wr_addr[0]), .B(wr_addr[2]), .C(n3224), .Z(n2110) );
  AN3 U429 ( .A(wr_addr[0]), .B(wr_addr[1]), .C(n3223), .Z(n2111) );
  AN3 U430 ( .A(wr_addr[0]), .B(n3224), .C(n3223), .Z(n2112) );
  IVAP U431 ( .A(wr_data[4]), .Z(n3097) );
  IVAP U432 ( .A(wr_data[5]), .Z(n3099) );
  IVAP U433 ( .A(wr_data[6]), .Z(n3100) );
  IVAP U434 ( .A(wr_data[7]), .Z(n3101) );
  IVAP U435 ( .A(wr_data[8]), .Z(n3102) );
  IVAP U436 ( .A(wr_data[9]), .Z(n3103) );
  IVAP U437 ( .A(wr_data[10]), .Z(n3104) );
  IVAP U438 ( .A(wr_data[11]), .Z(n3105) );
  IVAP U439 ( .A(wr_data[12]), .Z(n3106) );
  IVAP U440 ( .A(wr_data[13]), .Z(n3107) );
  IVAP U441 ( .A(wr_data[14]), .Z(n3108) );
  IVAP U442 ( .A(wr_data[15]), .Z(n3110) );
  IVAP U443 ( .A(wr_data[16]), .Z(n3111) );
  IVAP U444 ( .A(wr_data[17]), .Z(n3113) );
  IVAP U445 ( .A(wr_data[18]), .Z(n3114) );
  IVAP U446 ( .A(wr_data[19]), .Z(n3115) );
  IVAP U447 ( .A(wr_data[20]), .Z(n3116) );
  IVAP U448 ( .A(wr_data[21]), .Z(n3117) );
  IVAP U449 ( .A(wr_data[22]), .Z(n3118) );
  IVAP U450 ( .A(wr_data[23]), .Z(n3121) );
  IVAP U451 ( .A(wr_data[24]), .Z(n3122) );
  IVAP U452 ( .A(wr_data[25]), .Z(n3123) );
  IVAP U453 ( .A(wr_data[26]), .Z(n3124) );
  IVAP U454 ( .A(wr_data[27]), .Z(n3125) );
  IVAP U455 ( .A(wr_data[28]), .Z(n3126) );
  IVAP U456 ( .A(wr_data[29]), .Z(n3127) );
  IVAP U457 ( .A(wr_data[30]), .Z(n3129) );
  IVAP U458 ( .A(wr_data[31]), .Z(n3133) );
  IVAP U459 ( .A(wr_data[4]), .Z(n3098) );
  IVAP U460 ( .A(wr_data[14]), .Z(n3109) );
  IVAP U461 ( .A(wr_data[16]), .Z(n3112) );
  IVAP U462 ( .A(wr_data[22]), .Z(n3119) );
  IVAP U463 ( .A(wr_data[29]), .Z(n3128) );
  MUX31L U464 ( .D0(n60), .D1(n129), .D2(n3328), .A(n3177), .B(n3194), .Z(
        n3329) );
  MUX31L U465 ( .D0(\gpr[28][24] ), .D1(\gpr[29][24] ), .D2(n2737), .A(n2968), 
        .B(n2993), .Z(n2741) );
  MUX31L U466 ( .D0(\gpr[28][28] ), .D1(\gpr[29][28] ), .D2(n2841), .A(n51), 
        .B(n2993), .Z(n2845) );
  MUX31L U467 ( .D0(\gpr[28][27] ), .D1(\gpr[29][27] ), .D2(n2815), .A(n25), 
        .B(n2993), .Z(n2819) );
  MUX31L U468 ( .D0(\gpr[28][26] ), .D1(\gpr[29][26] ), .D2(n2789), .A(n51), 
        .B(n2993), .Z(n2793) );
  MUX31L U469 ( .D0(\gpr[28][0] ), .D1(\gpr[29][0] ), .D2(n2113), .A(n2961), 
        .B(n2991), .Z(n2117) );
  MUX31L U470 ( .D0(\gpr[28][31] ), .D1(\gpr[29][31] ), .D2(n2919), .A(n25), 
        .B(n2993), .Z(n2923) );
  MUX31L U471 ( .D0(\gpr[28][30] ), .D1(\gpr[29][30] ), .D2(n2893), .A(n25), 
        .B(n2993), .Z(n2897) );
  MUX31L U472 ( .D0(\gpr[28][29] ), .D1(\gpr[29][29] ), .D2(n2867), .A(n2970), 
        .B(n2993), .Z(n2871) );
  MUX31L U473 ( .D0(\gpr[28][25] ), .D1(\gpr[29][25] ), .D2(n2763), .A(n2969), 
        .B(n2993), .Z(n2767) );
  MUX31L U474 ( .D0(\gpr[28][23] ), .D1(\gpr[29][23] ), .D2(n2711), .A(n2979), 
        .B(n2993), .Z(n2715) );
  MUX31L U475 ( .D0(\gpr[28][14] ), .D1(\gpr[29][14] ), .D2(n2477), .A(n2960), 
        .B(n2992), .Z(n2481) );
  MUX21H U476 ( .A(\gpr[30][0] ), .B(\gpr[31][0] ), .S(n2979), .Z(n2113) );
  MUX21L U477 ( .A(n2122), .B(n2123), .S(n2983), .Z(n2121) );
  MUX21L U478 ( .A(n2125), .B(n2126), .S(n2983), .Z(n2124) );
  MUX21L U479 ( .A(n2128), .B(n2129), .S(n2983), .Z(n2127) );
  MUX21L U480 ( .A(n2131), .B(n2132), .S(n2984), .Z(n2130) );
  MUX21L U481 ( .A(n2134), .B(n2135), .S(n2984), .Z(n2133) );
  MUX31LP U482 ( .D0(n2136), .D1(n2137), .D2(n2138), .A(n3000), .B(n3004), .Z(
        N120) );
  MUX21H U483 ( .A(\gpr[30][1] ), .B(\gpr[31][1] ), .S(n2960), .Z(n2139) );
  MUX21L U484 ( .A(n2145), .B(n2146), .S(n2984), .Z(n2144) );
  MUX21L U485 ( .A(n2148), .B(n2149), .S(n2984), .Z(n2147) );
  MUX21L U486 ( .A(n2151), .B(n2152), .S(n2984), .Z(n2150) );
  MUX21L U487 ( .A(n2154), .B(n2155), .S(n2984), .Z(n2153) );
  MUX21L U488 ( .A(n2157), .B(n2158), .S(n2984), .Z(n2156) );
  MUX21L U489 ( .A(n2160), .B(n2161), .S(n2984), .Z(n2159) );
  MUX31LP U490 ( .D0(n2162), .D1(n2163), .D2(n2164), .A(n3000), .B(n3004), .Z(
        N119) );
  MUX21H U491 ( .A(\gpr[30][2] ), .B(\gpr[31][2] ), .S(n2960), .Z(n2165) );
  MUX21L U492 ( .A(n2171), .B(n2172), .S(n2984), .Z(n2170) );
  MUX21L U493 ( .A(n2174), .B(n2175), .S(n2984), .Z(n2173) );
  MUX21L U494 ( .A(n2177), .B(n2178), .S(n2984), .Z(n2176) );
  MUX21L U495 ( .A(n2180), .B(n2181), .S(n2984), .Z(n2179) );
  MUX21L U496 ( .A(n2183), .B(n2184), .S(n2984), .Z(n2182) );
  MUX21L U497 ( .A(n2186), .B(n2187), .S(n2984), .Z(n2185) );
  MUX31LP U498 ( .D0(n2188), .D1(n2189), .D2(n2190), .A(n3000), .B(n3004), .Z(
        N118) );
  MUX21H U499 ( .A(\gpr[30][3] ), .B(\gpr[31][3] ), .S(n2960), .Z(n2191) );
  MUX21L U500 ( .A(n2197), .B(n2198), .S(n2984), .Z(n2196) );
  MUX21L U501 ( .A(n2200), .B(n2201), .S(n2984), .Z(n2199) );
  MUX21L U502 ( .A(n2203), .B(n2204), .S(n2985), .Z(n2202) );
  MUX21L U503 ( .A(n2206), .B(n2207), .S(n2985), .Z(n2205) );
  MUX21L U504 ( .A(n2209), .B(n2210), .S(n2985), .Z(n2208) );
  MUX21L U505 ( .A(n2212), .B(n2213), .S(n2985), .Z(n2211) );
  MUX31LP U506 ( .D0(n2214), .D1(n2215), .D2(n2216), .A(n3001), .B(n3004), .Z(
        N117) );
  MUX21H U507 ( .A(\gpr[30][4] ), .B(\gpr[31][4] ), .S(n2960), .Z(n2217) );
  MUX21L U508 ( .A(n2223), .B(n2224), .S(n2985), .Z(n2222) );
  MUX21L U509 ( .A(n2226), .B(n2227), .S(n2985), .Z(n2225) );
  MUX21L U510 ( .A(n2229), .B(n2230), .S(n2985), .Z(n2228) );
  MUX21L U511 ( .A(n2232), .B(n2233), .S(n2985), .Z(n2231) );
  MUX21L U512 ( .A(n2235), .B(n2236), .S(n2985), .Z(n2234) );
  MUX21L U513 ( .A(n2238), .B(n2239), .S(n2985), .Z(n2237) );
  MUX31LP U514 ( .D0(n2240), .D1(n2241), .D2(n2242), .A(n3001), .B(n3004), .Z(
        N116) );
  MUX21H U515 ( .A(\gpr[30][5] ), .B(\gpr[31][5] ), .S(n2960), .Z(n2243) );
  MUX21L U516 ( .A(n2249), .B(n2250), .S(n2985), .Z(n2248) );
  MUX21L U517 ( .A(n2252), .B(n2253), .S(n2985), .Z(n2251) );
  MUX21L U518 ( .A(n2255), .B(n2256), .S(n2985), .Z(n2254) );
  MUX21L U519 ( .A(n2258), .B(n2259), .S(n2985), .Z(n2257) );
  MUX21L U520 ( .A(n2261), .B(n2262), .S(n2985), .Z(n2260) );
  MUX21L U521 ( .A(n2264), .B(n2265), .S(n2985), .Z(n2263) );
  MUX31LP U522 ( .D0(n2266), .D1(n2267), .D2(n2268), .A(n3001), .B(n3004), .Z(
        N115) );
  MUX21H U523 ( .A(\gpr[30][6] ), .B(\gpr[31][6] ), .S(n2960), .Z(n2269) );
  MUX21L U524 ( .A(n2278), .B(n2279), .S(n2986), .Z(n2277) );
  MUX21L U525 ( .A(n2281), .B(n2282), .S(n2986), .Z(n2280) );
  MUX21L U526 ( .A(n2284), .B(n2285), .S(n2986), .Z(n2283) );
  MUX21L U527 ( .A(n2287), .B(n2288), .S(n2986), .Z(n2286) );
  MUX21L U528 ( .A(n2290), .B(n2291), .S(n2986), .Z(n2289) );
  MUX31LP U529 ( .D0(n2292), .D1(n2293), .D2(n2294), .A(n3001), .B(n3004), .Z(
        N114) );
  MUX21H U530 ( .A(\gpr[30][7] ), .B(\gpr[31][7] ), .S(n2960), .Z(n2295) );
  MUX21L U531 ( .A(n2301), .B(n2302), .S(n2986), .Z(n2300) );
  MUX21L U532 ( .A(n2304), .B(n2305), .S(n2986), .Z(n2303) );
  MUX21L U533 ( .A(n2307), .B(n2308), .S(n2986), .Z(n2306) );
  MUX21L U534 ( .A(n2310), .B(n2311), .S(n2986), .Z(n2309) );
  MUX21L U535 ( .A(n2313), .B(n2314), .S(n2986), .Z(n2312) );
  MUX21L U536 ( .A(n2316), .B(n2317), .S(n2986), .Z(n2315) );
  MUX31LP U537 ( .D0(n2318), .D1(n2319), .D2(n2320), .A(n3001), .B(n3004), .Z(
        N113) );
  MUX21H U538 ( .A(\gpr[30][8] ), .B(\gpr[31][8] ), .S(n2960), .Z(n2321) );
  MUX21L U539 ( .A(n2327), .B(n2328), .S(n2986), .Z(n2326) );
  MUX21L U540 ( .A(n2330), .B(n2331), .S(n2986), .Z(n2329) );
  MUX21L U541 ( .A(n2333), .B(n2334), .S(n2986), .Z(n2332) );
  MUX21L U542 ( .A(n2336), .B(n2337), .S(n2986), .Z(n2335) );
  MUX21L U543 ( .A(n2339), .B(n2340), .S(n2986), .Z(n2338) );
  MUX21L U544 ( .A(n2342), .B(n2343), .S(n2987), .Z(n2341) );
  MUX31LP U545 ( .D0(n2344), .D1(n2345), .D2(n2346), .A(n3001), .B(n3004), .Z(
        N112) );
  MUX21H U546 ( .A(\gpr[30][9] ), .B(\gpr[31][9] ), .S(n23), .Z(n2347) );
  MUX21L U547 ( .A(n2353), .B(n2354), .S(n2987), .Z(n2352) );
  MUX21L U548 ( .A(n2356), .B(n2357), .S(n2987), .Z(n2355) );
  MUX21L U549 ( .A(n2359), .B(n2360), .S(n2987), .Z(n2358) );
  MUX21L U550 ( .A(n2362), .B(n2363), .S(n2987), .Z(n2361) );
  MUX21L U551 ( .A(n2365), .B(n2366), .S(n2987), .Z(n2364) );
  MUX21L U552 ( .A(n2368), .B(n2369), .S(n2987), .Z(n2367) );
  MUX31LP U553 ( .D0(n2370), .D1(n2371), .D2(n2372), .A(n3001), .B(n3004), .Z(
        N111) );
  MUX21H U554 ( .A(\gpr[30][10] ), .B(\gpr[31][10] ), .S(n23), .Z(n2373) );
  MUX21L U555 ( .A(n2379), .B(n2380), .S(n2987), .Z(n2378) );
  MUX21L U556 ( .A(n2382), .B(n2383), .S(n2987), .Z(n2381) );
  MUX21L U557 ( .A(n2385), .B(n2386), .S(n2987), .Z(n2384) );
  MUX21L U558 ( .A(n2388), .B(n2389), .S(n2987), .Z(n2387) );
  MUX21L U559 ( .A(n2391), .B(n2392), .S(n2987), .Z(n2390) );
  MUX21L U560 ( .A(n2394), .B(n2395), .S(n2987), .Z(n2393) );
  MUX31LP U561 ( .D0(n2396), .D1(n2397), .D2(n2398), .A(n3001), .B(n3004), .Z(
        N110) );
  MUX21H U562 ( .A(\gpr[30][11] ), .B(\gpr[31][11] ), .S(n23), .Z(n2399) );
  MUX21L U563 ( .A(n2405), .B(n2406), .S(n2987), .Z(n2404) );
  MUX21L U564 ( .A(n2408), .B(n2409), .S(n2987), .Z(n2407) );
  MUX21L U565 ( .A(n2411), .B(n2412), .S(n2987), .Z(n2410) );
  MUX21L U566 ( .A(n2414), .B(n2415), .S(n45), .Z(n2413) );
  MUX21L U567 ( .A(n2417), .B(n2418), .S(n2986), .Z(n2416) );
  MUX21L U568 ( .A(n2420), .B(n2421), .S(n39), .Z(n2419) );
  MUX31LP U569 ( .D0(n2422), .D1(n2423), .D2(n2424), .A(n3001), .B(n3004), .Z(
        N109) );
  MUX21H U570 ( .A(\gpr[30][12] ), .B(\gpr[31][12] ), .S(n23), .Z(n2425) );
  MUX21L U571 ( .A(n2431), .B(n2432), .S(n39), .Z(n2430) );
  MUX21L U572 ( .A(n2434), .B(n2435), .S(n45), .Z(n2433) );
  MUX21L U573 ( .A(n2437), .B(n2438), .S(n39), .Z(n2436) );
  MUX21L U574 ( .A(n2440), .B(n2441), .S(n45), .Z(n2439) );
  MUX21L U575 ( .A(n2443), .B(n2444), .S(n39), .Z(n2442) );
  MUX21L U576 ( .A(n2446), .B(n2447), .S(n45), .Z(n2445) );
  MUX31LP U577 ( .D0(n2448), .D1(n2449), .D2(n2450), .A(n3001), .B(n3004), .Z(
        N108) );
  MUX21H U578 ( .A(\gpr[30][13] ), .B(\gpr[31][13] ), .S(n23), .Z(n2451) );
  MUX21L U579 ( .A(n2457), .B(n2458), .S(n45), .Z(n2456) );
  MUX21L U580 ( .A(n2460), .B(n2461), .S(n2990), .Z(n2459) );
  MUX21L U581 ( .A(n2463), .B(n2464), .S(n2990), .Z(n2462) );
  MUX21L U582 ( .A(n2466), .B(n2467), .S(n45), .Z(n2465) );
  MUX21L U583 ( .A(n2469), .B(n2470), .S(n2990), .Z(n2468) );
  MUX21L U584 ( .A(n2472), .B(n2473), .S(n39), .Z(n2471) );
  MUX31LP U585 ( .D0(n2474), .D1(n2475), .D2(n2476), .A(n3001), .B(n122), .Z(
        N107) );
  MUX21H U586 ( .A(\gpr[30][14] ), .B(\gpr[31][14] ), .S(n23), .Z(n2477) );
  MUX21L U587 ( .A(n2486), .B(n2487), .S(n2988), .Z(n2485) );
  MUX21L U588 ( .A(n2489), .B(n2490), .S(n2988), .Z(n2488) );
  MUX21L U589 ( .A(n2492), .B(n2493), .S(n2988), .Z(n2491) );
  MUX21L U590 ( .A(n2495), .B(n2496), .S(n2988), .Z(n2494) );
  MUX21L U591 ( .A(n2498), .B(n2499), .S(n2988), .Z(n2497) );
  MUX31LP U592 ( .D0(n2500), .D1(n2501), .D2(n2502), .A(n3001), .B(n122), .Z(
        N106) );
  MUX21H U593 ( .A(\gpr[30][15] ), .B(\gpr[31][15] ), .S(n23), .Z(n2503) );
  MUX21L U594 ( .A(n2509), .B(n2510), .S(n2988), .Z(n2508) );
  MUX21L U595 ( .A(n2512), .B(n2513), .S(n2988), .Z(n2511) );
  MUX21L U596 ( .A(n2515), .B(n2516), .S(n2988), .Z(n2514) );
  MUX21L U597 ( .A(n2518), .B(n2519), .S(n2988), .Z(n2517) );
  MUX21L U598 ( .A(n2521), .B(n2522), .S(n2988), .Z(n2520) );
  MUX21L U599 ( .A(n2524), .B(n2525), .S(n2988), .Z(n2523) );
  MUX31LP U600 ( .D0(n2526), .D1(n2527), .D2(n2528), .A(n3001), .B(n122), .Z(
        N105) );
  MUX21H U601 ( .A(\gpr[30][16] ), .B(\gpr[31][16] ), .S(n23), .Z(n2529) );
  MUX21L U602 ( .A(n2535), .B(n2536), .S(n2988), .Z(n2534) );
  MUX21L U603 ( .A(n2538), .B(n2539), .S(n2988), .Z(n2537) );
  MUX21L U604 ( .A(n2541), .B(n2542), .S(n2988), .Z(n2540) );
  MUX21L U605 ( .A(n2544), .B(n2545), .S(n2988), .Z(n2543) );
  MUX21L U606 ( .A(n2547), .B(n2548), .S(n2988), .Z(n2546) );
  MUX21L U607 ( .A(n2550), .B(n2551), .S(n2988), .Z(n2549) );
  MUX31LP U608 ( .D0(n2552), .D1(n2553), .D2(n2554), .A(n3001), .B(n122), .Z(
        N104) );
  MUX21H U609 ( .A(\gpr[30][17] ), .B(\gpr[31][17] ), .S(n23), .Z(n2555) );
  MUX21L U610 ( .A(n2561), .B(n2562), .S(n2989), .Z(n2560) );
  MUX21L U611 ( .A(n2564), .B(n2565), .S(n2989), .Z(n2563) );
  MUX21L U612 ( .A(n2567), .B(n2568), .S(n2989), .Z(n2566) );
  MUX21L U613 ( .A(n2570), .B(n2571), .S(n2989), .Z(n2569) );
  MUX21L U614 ( .A(n2573), .B(n2574), .S(n2989), .Z(n2572) );
  MUX21L U615 ( .A(n2576), .B(n2577), .S(n2989), .Z(n2575) );
  MUX31LP U616 ( .D0(n2578), .D1(n2579), .D2(n2580), .A(n3001), .B(n122), .Z(
        N103) );
  MUX21H U617 ( .A(\gpr[30][18] ), .B(\gpr[31][18] ), .S(n23), .Z(n2581) );
  MUX21L U618 ( .A(n2587), .B(n2588), .S(n2989), .Z(n2586) );
  MUX21L U619 ( .A(n2590), .B(n2591), .S(n2989), .Z(n2589) );
  MUX21L U620 ( .A(n2593), .B(n2594), .S(n2989), .Z(n2592) );
  MUX21L U621 ( .A(n2596), .B(n2597), .S(n2989), .Z(n2595) );
  MUX21L U622 ( .A(n2599), .B(n2600), .S(n2989), .Z(n2598) );
  MUX21L U623 ( .A(n2602), .B(n2603), .S(n2989), .Z(n2601) );
  MUX31LP U624 ( .D0(n2604), .D1(n2605), .D2(n2606), .A(n3001), .B(n122), .Z(
        N102) );
  MUX21H U625 ( .A(\gpr[30][19] ), .B(\gpr[31][19] ), .S(n23), .Z(n2607) );
  MUX21L U626 ( .A(n2613), .B(n2614), .S(n2989), .Z(n2612) );
  MUX21L U627 ( .A(n2616), .B(n2617), .S(n2989), .Z(n2615) );
  MUX21L U628 ( .A(n2619), .B(n2620), .S(n2989), .Z(n2618) );
  MUX21L U629 ( .A(n2622), .B(n2623), .S(n2989), .Z(n2621) );
  MUX21L U630 ( .A(n2625), .B(n2626), .S(n45), .Z(n2624) );
  MUX21L U631 ( .A(n2628), .B(n2629), .S(n45), .Z(n2627) );
  MUX31LP U632 ( .D0(n2630), .D1(n2631), .D2(n2632), .A(n3001), .B(n122), .Z(
        N101) );
  MUX21H U633 ( .A(\gpr[30][20] ), .B(\gpr[31][20] ), .S(n23), .Z(n2633) );
  MUX21L U634 ( .A(n2639), .B(n2640), .S(n45), .Z(n2638) );
  MUX21L U635 ( .A(n2642), .B(n2643), .S(n45), .Z(n2641) );
  MUX21L U636 ( .A(n2645), .B(n2646), .S(n45), .Z(n2644) );
  MUX21L U637 ( .A(n2648), .B(n2649), .S(n45), .Z(n2647) );
  MUX21L U638 ( .A(n2651), .B(n2652), .S(n45), .Z(n2650) );
  MUX21L U639 ( .A(n2654), .B(n2655), .S(n45), .Z(n2653) );
  MUX31LP U640 ( .D0(n2656), .D1(n2657), .D2(n2658), .A(n3001), .B(n122), .Z(
        N100) );
  MUX21H U641 ( .A(\gpr[30][21] ), .B(\gpr[31][21] ), .S(n23), .Z(n2659) );
  MUX21L U642 ( .A(n2665), .B(n2666), .S(n45), .Z(n2664) );
  MUX21L U643 ( .A(n2668), .B(n2669), .S(n45), .Z(n2667) );
  MUX21L U644 ( .A(n2671), .B(n2672), .S(n45), .Z(n2670) );
  MUX21L U645 ( .A(n2674), .B(n2675), .S(n45), .Z(n2673) );
  MUX21L U646 ( .A(n2677), .B(n2678), .S(n45), .Z(n2676) );
  MUX21L U647 ( .A(n2680), .B(n2681), .S(n45), .Z(n2679) );
  MUX31LP U648 ( .D0(n2682), .D1(n2683), .D2(n2684), .A(n3001), .B(n122), .Z(
        N99) );
  MUX21H U649 ( .A(\gpr[30][22] ), .B(\gpr[31][22] ), .S(n23), .Z(n2685) );
  MUX21L U650 ( .A(n2691), .B(n2692), .S(n45), .Z(n2690) );
  MUX21L U651 ( .A(n2694), .B(n2695), .S(n45), .Z(n2693) );
  MUX21L U652 ( .A(n2697), .B(n2698), .S(n2990), .Z(n2696) );
  MUX21L U653 ( .A(n2700), .B(n2701), .S(n2990), .Z(n2699) );
  MUX21L U654 ( .A(n2703), .B(n2704), .S(n2990), .Z(n2702) );
  MUX21L U655 ( .A(n2706), .B(n2707), .S(n2990), .Z(n2705) );
  MUX31LP U656 ( .D0(n2708), .D1(n2709), .D2(n2710), .A(n53), .B(n122), .Z(N98) );
  MUX21H U657 ( .A(\gpr[30][23] ), .B(\gpr[31][23] ), .S(n2961), .Z(n2711) );
  MUX21L U658 ( .A(n2720), .B(n2721), .S(n2990), .Z(n2719) );
  MUX21L U659 ( .A(n2723), .B(n2724), .S(n2990), .Z(n2722) );
  MUX21L U660 ( .A(n2726), .B(n2727), .S(n2990), .Z(n2725) );
  MUX21L U661 ( .A(n2729), .B(n2730), .S(n2990), .Z(n2728) );
  MUX21L U662 ( .A(n2732), .B(n2733), .S(n2990), .Z(n2731) );
  MUX31LP U663 ( .D0(n2734), .D1(n2735), .D2(n2736), .A(n53), .B(n122), .Z(N97) );
  MUX21H U664 ( .A(\gpr[30][24] ), .B(\gpr[31][24] ), .S(n2961), .Z(n2737) );
  MUX31LP U665 ( .D0(n2739), .D1(n2740), .D2(n2741), .A(n2990), .B(n2999), .Z(
        n2738) );
  MUX21L U666 ( .A(n2743), .B(n2744), .S(n2990), .Z(n2742) );
  MUX21L U667 ( .A(n2746), .B(n2747), .S(n2990), .Z(n2745) );
  MUX21L U668 ( .A(n2749), .B(n2750), .S(n2990), .Z(n2748) );
  MUX21L U669 ( .A(n2752), .B(n2753), .S(n2990), .Z(n2751) );
  MUX21L U670 ( .A(n2755), .B(n2756), .S(n2990), .Z(n2754) );
  MUX21L U671 ( .A(n2758), .B(n2759), .S(n2990), .Z(n2757) );
  MUX31LP U672 ( .D0(n2760), .D1(n2761), .D2(n2762), .A(n53), .B(n122), .Z(N96) );
  MUX21H U673 ( .A(\gpr[30][25] ), .B(\gpr[31][25] ), .S(n2961), .Z(n2763) );
  MUX31LP U674 ( .D0(n2765), .D1(n2766), .D2(n2767), .A(n2990), .B(n2999), .Z(
        n2764) );
  MUX21L U675 ( .A(n2769), .B(n2770), .S(n39), .Z(n2768) );
  MUX21L U676 ( .A(n2772), .B(n2773), .S(n39), .Z(n2771) );
  MUX21L U677 ( .A(n2775), .B(n2776), .S(n39), .Z(n2774) );
  MUX21L U678 ( .A(n2778), .B(n2779), .S(n39), .Z(n2777) );
  MUX21L U679 ( .A(n2781), .B(n2782), .S(n39), .Z(n2780) );
  MUX21L U680 ( .A(n2784), .B(n2785), .S(n39), .Z(n2783) );
  MUX31LP U681 ( .D0(n2786), .D1(n2787), .D2(n2788), .A(n53), .B(n122), .Z(N95) );
  MUX21H U682 ( .A(\gpr[30][26] ), .B(\gpr[31][26] ), .S(n2961), .Z(n2789) );
  MUX31LP U683 ( .D0(n2791), .D1(n2792), .D2(n2793), .A(n39), .B(n2997), .Z(
        n2790) );
  MUX21L U684 ( .A(n2795), .B(n2796), .S(n39), .Z(n2794) );
  MUX21L U685 ( .A(n2798), .B(n2799), .S(n39), .Z(n2797) );
  MUX21L U686 ( .A(n2801), .B(n2802), .S(n39), .Z(n2800) );
  MUX21L U687 ( .A(n2804), .B(n2805), .S(n39), .Z(n2803) );
  MUX21L U688 ( .A(n2807), .B(n2808), .S(n39), .Z(n2806) );
  MUX21L U689 ( .A(n2810), .B(n2811), .S(n39), .Z(n2809) );
  MUX31LP U690 ( .D0(n2812), .D1(n2813), .D2(n2814), .A(n53), .B(n3004), .Z(
        N94) );
  MUX21H U691 ( .A(\gpr[30][27] ), .B(\gpr[31][27] ), .S(n2961), .Z(n2815) );
  MUX31LP U692 ( .D0(n2817), .D1(n2818), .D2(n2819), .A(n39), .B(n120), .Z(
        n2816) );
  MUX21L U693 ( .A(n2821), .B(n2822), .S(n39), .Z(n2820) );
  MUX21L U694 ( .A(n2824), .B(n2825), .S(n39), .Z(n2823) );
  MUX21L U695 ( .A(n2827), .B(n2828), .S(n39), .Z(n2826) );
  MUX21L U696 ( .A(n2830), .B(n2831), .S(n39), .Z(n2829) );
  MUX21L U697 ( .A(n2833), .B(n2834), .S(n39), .Z(n2832) );
  MUX21L U698 ( .A(n2836), .B(n2837), .S(n2984), .Z(n2835) );
  MUX31LP U699 ( .D0(n2838), .D1(n2839), .D2(n2840), .A(n53), .B(n122), .Z(N93) );
  MUX21H U700 ( .A(\gpr[30][28] ), .B(\gpr[31][28] ), .S(n2961), .Z(n2841) );
  MUX31LP U701 ( .D0(n2843), .D1(n2844), .D2(n2845), .A(n2990), .B(n120), .Z(
        n2842) );
  MUX21L U702 ( .A(n2847), .B(n2848), .S(n39), .Z(n2846) );
  MUX21L U703 ( .A(n2850), .B(n2851), .S(n2990), .Z(n2849) );
  MUX21L U704 ( .A(n2853), .B(n2854), .S(n2983), .Z(n2852) );
  MUX21L U705 ( .A(n2856), .B(n2857), .S(n39), .Z(n2855) );
  MUX21L U706 ( .A(n2859), .B(n2860), .S(n2990), .Z(n2858) );
  MUX21L U707 ( .A(n2862), .B(n2863), .S(n39), .Z(n2861) );
  MUX31LP U708 ( .D0(n2864), .D1(n2865), .D2(n2866), .A(n53), .B(n122), .Z(N92) );
  MUX21H U709 ( .A(\gpr[30][29] ), .B(\gpr[31][29] ), .S(n2961), .Z(n2867) );
  MUX21L U710 ( .A(n2876), .B(n2877), .S(n39), .Z(n2875) );
  MUX21L U711 ( .A(n2879), .B(n2880), .S(n2990), .Z(n2878) );
  MUX21L U712 ( .A(n2882), .B(n2883), .S(n2984), .Z(n2881) );
  MUX21L U713 ( .A(n2885), .B(n2886), .S(n39), .Z(n2884) );
  MUX21L U714 ( .A(n2888), .B(n2889), .S(n2990), .Z(n2887) );
  MUX31LP U715 ( .D0(n2890), .D1(n2891), .D2(n2892), .A(n53), .B(n3004), .Z(
        N91) );
  MUX21H U716 ( .A(\gpr[30][30] ), .B(\gpr[31][30] ), .S(n2961), .Z(n2893) );
  MUX21L U717 ( .A(n2902), .B(n2903), .S(n2990), .Z(n2901) );
  MUX21L U718 ( .A(n2905), .B(n2906), .S(n2983), .Z(n2904) );
  MUX21L U719 ( .A(n2908), .B(n2909), .S(n2991), .Z(n2907) );
  MUX21L U720 ( .A(n2911), .B(n2912), .S(n2991), .Z(n2910) );
  MUX21L U721 ( .A(n2914), .B(n2915), .S(n2991), .Z(n2913) );
  MUX31LP U722 ( .D0(n2916), .D1(n2917), .D2(n2918), .A(n53), .B(n3004), .Z(
        N90) );
  MUX21H U723 ( .A(\gpr[30][31] ), .B(\gpr[31][31] ), .S(n2961), .Z(n2919) );
  MUX21L U724 ( .A(n2925), .B(n2926), .S(n2991), .Z(n2924) );
  MUX21L U725 ( .A(n2928), .B(n2929), .S(n2991), .Z(n2927) );
  MUX21L U726 ( .A(n2931), .B(n2932), .S(n2991), .Z(n2930) );
  MUX21L U727 ( .A(n2934), .B(n2935), .S(n2991), .Z(n2933) );
  MUX21L U728 ( .A(n2937), .B(n2938), .S(n2991), .Z(n2936) );
  MUX21L U729 ( .A(n2940), .B(n2941), .S(n2991), .Z(n2939) );
  MUX31LP U730 ( .D0(n2942), .D1(n2943), .D2(n2944), .A(n53), .B(n122), .Z(N89) );
  MUX21L U731 ( .A(\gpr[26][0] ), .B(\gpr[27][0] ), .S(n2961), .Z(n2116) );
  MUX21L U732 ( .A(\gpr[24][0] ), .B(\gpr[25][0] ), .S(n2961), .Z(n2115) );
  MUX21L U733 ( .A(\gpr[22][0] ), .B(\gpr[23][0] ), .S(n2961), .Z(n2120) );
  MUX21L U734 ( .A(\gpr[20][0] ), .B(\gpr[21][0] ), .S(n2961), .Z(n2119) );
  MUX21L U735 ( .A(\gpr[18][0] ), .B(\gpr[19][0] ), .S(n2962), .Z(n2123) );
  MUX21L U736 ( .A(\gpr[16][0] ), .B(\gpr[17][0] ), .S(n2962), .Z(n2122) );
  MUX31LP U737 ( .D0(n2121), .D1(n2118), .D2(n2114), .A(n120), .B(n53), .Z(
        n2138) );
  MUX21L U738 ( .A(\gpr[14][0] ), .B(\gpr[15][0] ), .S(n2962), .Z(n2126) );
  MUX21L U739 ( .A(\gpr[12][0] ), .B(\gpr[13][0] ), .S(n2962), .Z(n2125) );
  MUX21L U740 ( .A(\gpr[10][0] ), .B(\gpr[11][0] ), .S(n2962), .Z(n2129) );
  MUX21L U741 ( .A(\gpr[8][0] ), .B(\gpr[9][0] ), .S(n2962), .Z(n2128) );
  MUX21L U742 ( .A(n2127), .B(n2124), .S(n120), .Z(n2137) );
  MUX21L U743 ( .A(\gpr[6][0] ), .B(\gpr[7][0] ), .S(n2962), .Z(n2132) );
  MUX21L U744 ( .A(\gpr[4][0] ), .B(\gpr[5][0] ), .S(n2962), .Z(n2131) );
  MUX21L U745 ( .A(\gpr[2][0] ), .B(\gpr[3][0] ), .S(n2962), .Z(n2135) );
  ND2I U746 ( .A(n2952), .B(\gpr[1][0] ), .Z(n2134) );
  MUX21L U747 ( .A(n2133), .B(n2130), .S(n2997), .Z(n2136) );
  MUX21L U748 ( .A(\gpr[26][1] ), .B(\gpr[27][1] ), .S(n2962), .Z(n2142) );
  MUX21L U749 ( .A(\gpr[24][1] ), .B(\gpr[25][1] ), .S(n2962), .Z(n2141) );
  MUX21L U750 ( .A(\gpr[22][1] ), .B(\gpr[23][1] ), .S(n2962), .Z(n2146) );
  MUX21L U751 ( .A(\gpr[20][1] ), .B(\gpr[21][1] ), .S(n2962), .Z(n2145) );
  MUX21L U752 ( .A(\gpr[18][1] ), .B(\gpr[19][1] ), .S(n2963), .Z(n2149) );
  MUX21L U753 ( .A(\gpr[16][1] ), .B(\gpr[17][1] ), .S(n2963), .Z(n2148) );
  MUX31LP U754 ( .D0(n2147), .D1(n2144), .D2(n2140), .A(n2997), .B(n53), .Z(
        n2164) );
  MUX21L U755 ( .A(\gpr[14][1] ), .B(\gpr[15][1] ), .S(n2963), .Z(n2152) );
  MUX21L U756 ( .A(\gpr[12][1] ), .B(\gpr[13][1] ), .S(n2963), .Z(n2151) );
  MUX21L U757 ( .A(\gpr[10][1] ), .B(\gpr[11][1] ), .S(n2963), .Z(n2155) );
  MUX21L U758 ( .A(\gpr[8][1] ), .B(\gpr[9][1] ), .S(n2963), .Z(n2154) );
  MUX21L U759 ( .A(n2153), .B(n2150), .S(n120), .Z(n2163) );
  MUX21L U760 ( .A(\gpr[6][1] ), .B(\gpr[7][1] ), .S(n2963), .Z(n2158) );
  MUX21L U761 ( .A(\gpr[4][1] ), .B(\gpr[5][1] ), .S(n2963), .Z(n2157) );
  MUX21L U762 ( .A(\gpr[2][1] ), .B(\gpr[3][1] ), .S(n2963), .Z(n2161) );
  ND2I U763 ( .A(\gpr[1][1] ), .B(n51), .Z(n2160) );
  MUX21L U764 ( .A(n2159), .B(n2156), .S(n2997), .Z(n2162) );
  MUX21L U765 ( .A(\gpr[26][2] ), .B(\gpr[27][2] ), .S(n2963), .Z(n2168) );
  MUX21L U766 ( .A(\gpr[24][2] ), .B(\gpr[25][2] ), .S(n2963), .Z(n2167) );
  MUX21L U767 ( .A(\gpr[22][2] ), .B(\gpr[23][2] ), .S(n2963), .Z(n2172) );
  MUX21L U768 ( .A(\gpr[20][2] ), .B(\gpr[21][2] ), .S(n2964), .Z(n2171) );
  MUX21L U769 ( .A(\gpr[18][2] ), .B(\gpr[19][2] ), .S(n2964), .Z(n2175) );
  MUX21L U770 ( .A(\gpr[16][2] ), .B(\gpr[17][2] ), .S(n2964), .Z(n2174) );
  MUX31LP U771 ( .D0(n2173), .D1(n2170), .D2(n2166), .A(n2997), .B(n53), .Z(
        n2190) );
  MUX21L U772 ( .A(\gpr[14][2] ), .B(\gpr[15][2] ), .S(n2964), .Z(n2178) );
  MUX21L U773 ( .A(\gpr[12][2] ), .B(\gpr[13][2] ), .S(n2964), .Z(n2177) );
  MUX21L U774 ( .A(\gpr[10][2] ), .B(\gpr[11][2] ), .S(n2964), .Z(n2181) );
  MUX21L U775 ( .A(\gpr[8][2] ), .B(\gpr[9][2] ), .S(n2964), .Z(n2180) );
  MUX21L U776 ( .A(n2179), .B(n2176), .S(n120), .Z(n2189) );
  MUX21L U777 ( .A(\gpr[6][2] ), .B(\gpr[7][2] ), .S(n2964), .Z(n2184) );
  MUX21L U778 ( .A(\gpr[4][2] ), .B(\gpr[5][2] ), .S(n2964), .Z(n2183) );
  MUX21L U779 ( .A(\gpr[2][2] ), .B(\gpr[3][2] ), .S(n2964), .Z(n2187) );
  ND2I U780 ( .A(\gpr[1][2] ), .B(n51), .Z(n2186) );
  MUX21L U781 ( .A(n2185), .B(n2182), .S(n2997), .Z(n2188) );
  MUX21L U782 ( .A(\gpr[26][3] ), .B(\gpr[27][3] ), .S(n2964), .Z(n2194) );
  MUX21L U783 ( .A(\gpr[24][3] ), .B(\gpr[25][3] ), .S(n2964), .Z(n2193) );
  MUX21L U784 ( .A(\gpr[22][3] ), .B(\gpr[23][3] ), .S(n2964), .Z(n2198) );
  MUX21L U785 ( .A(\gpr[20][3] ), .B(\gpr[21][3] ), .S(n2965), .Z(n2197) );
  MUX21L U786 ( .A(\gpr[18][3] ), .B(\gpr[19][3] ), .S(n2965), .Z(n2201) );
  MUX21L U787 ( .A(\gpr[16][3] ), .B(\gpr[17][3] ), .S(n2965), .Z(n2200) );
  MUX31LP U788 ( .D0(n2199), .D1(n2196), .D2(n2192), .A(n120), .B(n53), .Z(
        n2216) );
  MUX21L U789 ( .A(\gpr[14][3] ), .B(\gpr[15][3] ), .S(n2965), .Z(n2204) );
  MUX21L U790 ( .A(\gpr[12][3] ), .B(\gpr[13][3] ), .S(n2965), .Z(n2203) );
  MUX21L U791 ( .A(\gpr[10][3] ), .B(\gpr[11][3] ), .S(n2965), .Z(n2207) );
  MUX21L U792 ( .A(\gpr[8][3] ), .B(\gpr[9][3] ), .S(n2965), .Z(n2206) );
  MUX21L U793 ( .A(n2205), .B(n2202), .S(n2998), .Z(n2215) );
  MUX21L U794 ( .A(\gpr[6][3] ), .B(\gpr[7][3] ), .S(n2965), .Z(n2210) );
  MUX21L U795 ( .A(\gpr[4][3] ), .B(\gpr[5][3] ), .S(n2965), .Z(n2209) );
  MUX21L U796 ( .A(\gpr[2][3] ), .B(\gpr[3][3] ), .S(n2965), .Z(n2213) );
  ND2I U797 ( .A(\gpr[1][3] ), .B(n51), .Z(n2212) );
  MUX21L U798 ( .A(n2211), .B(n2208), .S(n2998), .Z(n2214) );
  MUX21L U799 ( .A(\gpr[26][4] ), .B(\gpr[27][4] ), .S(n2965), .Z(n2220) );
  MUX21L U800 ( .A(\gpr[24][4] ), .B(\gpr[25][4] ), .S(n2965), .Z(n2219) );
  MUX21L U801 ( .A(\gpr[22][4] ), .B(\gpr[23][4] ), .S(n2965), .Z(n2224) );
  MUX21L U802 ( .A(\gpr[20][4] ), .B(\gpr[21][4] ), .S(n2966), .Z(n2223) );
  MUX21L U803 ( .A(\gpr[18][4] ), .B(\gpr[19][4] ), .S(n2966), .Z(n2227) );
  MUX21L U804 ( .A(\gpr[16][4] ), .B(\gpr[17][4] ), .S(n2966), .Z(n2226) );
  MUX31LP U805 ( .D0(n2225), .D1(n2222), .D2(n2218), .A(n2998), .B(n53), .Z(
        n2242) );
  MUX21L U806 ( .A(\gpr[14][4] ), .B(\gpr[15][4] ), .S(n2966), .Z(n2230) );
  MUX21L U807 ( .A(\gpr[12][4] ), .B(\gpr[13][4] ), .S(n2966), .Z(n2229) );
  MUX21L U808 ( .A(\gpr[10][4] ), .B(\gpr[11][4] ), .S(n2966), .Z(n2233) );
  MUX21L U809 ( .A(\gpr[8][4] ), .B(\gpr[9][4] ), .S(n2966), .Z(n2232) );
  MUX21L U810 ( .A(n2231), .B(n2228), .S(n2998), .Z(n2241) );
  MUX21L U811 ( .A(\gpr[6][4] ), .B(\gpr[7][4] ), .S(n2966), .Z(n2236) );
  MUX21L U812 ( .A(\gpr[4][4] ), .B(\gpr[5][4] ), .S(n2966), .Z(n2235) );
  MUX21L U813 ( .A(\gpr[2][4] ), .B(\gpr[3][4] ), .S(n2966), .Z(n2239) );
  ND2I U814 ( .A(\gpr[1][4] ), .B(n51), .Z(n2238) );
  MUX21L U815 ( .A(n2237), .B(n2234), .S(n2998), .Z(n2240) );
  MUX21L U816 ( .A(\gpr[26][5] ), .B(\gpr[27][5] ), .S(n2966), .Z(n2246) );
  MUX21L U817 ( .A(\gpr[24][5] ), .B(\gpr[25][5] ), .S(n2966), .Z(n2245) );
  MUX21L U818 ( .A(\gpr[22][5] ), .B(\gpr[23][5] ), .S(n2966), .Z(n2250) );
  MUX21L U819 ( .A(\gpr[20][5] ), .B(\gpr[21][5] ), .S(n2967), .Z(n2249) );
  MUX21L U820 ( .A(\gpr[18][5] ), .B(\gpr[19][5] ), .S(n2967), .Z(n2253) );
  MUX21L U821 ( .A(\gpr[16][5] ), .B(\gpr[17][5] ), .S(n2967), .Z(n2252) );
  MUX31LP U822 ( .D0(n2251), .D1(n2248), .D2(n2244), .A(n2998), .B(n53), .Z(
        n2268) );
  MUX21L U823 ( .A(\gpr[14][5] ), .B(\gpr[15][5] ), .S(n2967), .Z(n2256) );
  MUX21L U824 ( .A(\gpr[12][5] ), .B(\gpr[13][5] ), .S(n2967), .Z(n2255) );
  MUX21L U825 ( .A(\gpr[10][5] ), .B(\gpr[11][5] ), .S(n2967), .Z(n2259) );
  MUX21L U826 ( .A(\gpr[8][5] ), .B(\gpr[9][5] ), .S(n2967), .Z(n2258) );
  MUX21L U827 ( .A(n2257), .B(n2254), .S(n2998), .Z(n2267) );
  MUX21L U828 ( .A(\gpr[6][5] ), .B(\gpr[7][5] ), .S(n2967), .Z(n2262) );
  MUX21L U829 ( .A(\gpr[4][5] ), .B(\gpr[5][5] ), .S(n2967), .Z(n2261) );
  MUX21L U830 ( .A(\gpr[2][5] ), .B(\gpr[3][5] ), .S(n2967), .Z(n2265) );
  ND2I U831 ( .A(\gpr[1][5] ), .B(n2952), .Z(n2264) );
  MUX21L U832 ( .A(n2263), .B(n2260), .S(n2998), .Z(n2266) );
  MUX21L U833 ( .A(\gpr[26][6] ), .B(\gpr[27][6] ), .S(n2967), .Z(n2272) );
  MUX21L U834 ( .A(\gpr[24][6] ), .B(\gpr[25][6] ), .S(n2967), .Z(n2271) );
  MUX21L U835 ( .A(\gpr[22][6] ), .B(\gpr[23][6] ), .S(n2967), .Z(n2276) );
  MUX21L U836 ( .A(\gpr[20][6] ), .B(\gpr[21][6] ), .S(n47), .Z(n2275) );
  MUX21L U837 ( .A(\gpr[18][6] ), .B(\gpr[19][6] ), .S(n47), .Z(n2279) );
  MUX21L U838 ( .A(\gpr[16][6] ), .B(\gpr[17][6] ), .S(n47), .Z(n2278) );
  MUX31LP U839 ( .D0(n2277), .D1(n2274), .D2(n2270), .A(n2998), .B(n3002), .Z(
        n2294) );
  MUX21L U840 ( .A(\gpr[14][6] ), .B(\gpr[15][6] ), .S(n47), .Z(n2282) );
  MUX21L U841 ( .A(\gpr[12][6] ), .B(\gpr[13][6] ), .S(n2963), .Z(n2281) );
  MUX21L U842 ( .A(\gpr[10][6] ), .B(\gpr[11][6] ), .S(n2955), .Z(n2285) );
  MUX21L U843 ( .A(\gpr[8][6] ), .B(\gpr[9][6] ), .S(n51), .Z(n2284) );
  MUX21L U844 ( .A(n2283), .B(n2280), .S(n2998), .Z(n2293) );
  MUX21L U845 ( .A(\gpr[6][6] ), .B(\gpr[7][6] ), .S(n2953), .Z(n2288) );
  MUX21L U846 ( .A(\gpr[4][6] ), .B(\gpr[5][6] ), .S(n51), .Z(n2287) );
  MUX21L U847 ( .A(\gpr[2][6] ), .B(\gpr[3][6] ), .S(n2955), .Z(n2291) );
  ND2I U848 ( .A(\gpr[1][6] ), .B(n2952), .Z(n2290) );
  MUX21L U849 ( .A(n2289), .B(n2286), .S(n2998), .Z(n2292) );
  MUX21L U850 ( .A(\gpr[26][7] ), .B(\gpr[27][7] ), .S(n2953), .Z(n2298) );
  MUX21L U851 ( .A(\gpr[24][7] ), .B(\gpr[25][7] ), .S(n51), .Z(n2297) );
  MUX21L U852 ( .A(\gpr[22][7] ), .B(\gpr[23][7] ), .S(n2953), .Z(n2302) );
  MUX21L U853 ( .A(\gpr[20][7] ), .B(\gpr[21][7] ), .S(n2953), .Z(n2301) );
  MUX21L U854 ( .A(\gpr[18][7] ), .B(\gpr[19][7] ), .S(n2955), .Z(n2305) );
  MUX21L U855 ( .A(\gpr[16][7] ), .B(\gpr[17][7] ), .S(n2953), .Z(n2304) );
  MUX31LP U856 ( .D0(n2303), .D1(n2300), .D2(n2296), .A(n2998), .B(n3002), .Z(
        n2320) );
  MUX21L U857 ( .A(\gpr[14][7] ), .B(\gpr[15][7] ), .S(n2953), .Z(n2308) );
  MUX21L U858 ( .A(\gpr[12][7] ), .B(\gpr[13][7] ), .S(n2953), .Z(n2307) );
  MUX21L U859 ( .A(\gpr[10][7] ), .B(\gpr[11][7] ), .S(n2953), .Z(n2311) );
  MUX21L U860 ( .A(\gpr[8][7] ), .B(\gpr[9][7] ), .S(n2954), .Z(n2310) );
  MUX21L U861 ( .A(n2309), .B(n2306), .S(n2998), .Z(n2319) );
  MUX21L U862 ( .A(\gpr[6][7] ), .B(\gpr[7][7] ), .S(n2953), .Z(n2314) );
  MUX21L U863 ( .A(\gpr[4][7] ), .B(\gpr[5][7] ), .S(n2954), .Z(n2313) );
  MUX21L U864 ( .A(\gpr[2][7] ), .B(\gpr[3][7] ), .S(n2953), .Z(n2317) );
  ND2I U865 ( .A(\gpr[1][7] ), .B(n51), .Z(n2316) );
  MUX21L U866 ( .A(n2315), .B(n2312), .S(n2998), .Z(n2318) );
  MUX21L U867 ( .A(\gpr[26][8] ), .B(\gpr[27][8] ), .S(n2954), .Z(n2324) );
  MUX21L U868 ( .A(\gpr[24][8] ), .B(\gpr[25][8] ), .S(n2953), .Z(n2323) );
  MUX21L U869 ( .A(\gpr[22][8] ), .B(\gpr[23][8] ), .S(n2953), .Z(n2328) );
  MUX21L U870 ( .A(\gpr[20][8] ), .B(\gpr[21][8] ), .S(n2954), .Z(n2327) );
  MUX21L U871 ( .A(\gpr[18][8] ), .B(\gpr[19][8] ), .S(n2953), .Z(n2331) );
  MUX21L U872 ( .A(\gpr[16][8] ), .B(\gpr[17][8] ), .S(n2953), .Z(n2330) );
  MUX31LP U873 ( .D0(n2329), .D1(n2326), .D2(n2322), .A(n2998), .B(n3002), .Z(
        n2346) );
  MUX21L U874 ( .A(\gpr[14][8] ), .B(\gpr[15][8] ), .S(n2954), .Z(n2334) );
  MUX21L U875 ( .A(\gpr[12][8] ), .B(\gpr[13][8] ), .S(n2954), .Z(n2333) );
  MUX21L U876 ( .A(\gpr[10][8] ), .B(\gpr[11][8] ), .S(n2954), .Z(n2337) );
  MUX21L U877 ( .A(\gpr[8][8] ), .B(\gpr[9][8] ), .S(n2954), .Z(n2336) );
  MUX21L U878 ( .A(n2335), .B(n2332), .S(n2998), .Z(n2345) );
  MUX21L U879 ( .A(\gpr[6][8] ), .B(\gpr[7][8] ), .S(n2954), .Z(n2340) );
  MUX21L U880 ( .A(\gpr[4][8] ), .B(\gpr[5][8] ), .S(n2954), .Z(n2339) );
  MUX21L U881 ( .A(\gpr[2][8] ), .B(\gpr[3][8] ), .S(n2954), .Z(n2343) );
  ND2I U882 ( .A(\gpr[1][8] ), .B(n51), .Z(n2342) );
  MUX21L U883 ( .A(n2341), .B(n2338), .S(n2998), .Z(n2344) );
  MUX21L U884 ( .A(\gpr[26][9] ), .B(\gpr[27][9] ), .S(n2955), .Z(n2350) );
  MUX21L U885 ( .A(\gpr[24][9] ), .B(\gpr[25][9] ), .S(n2954), .Z(n2349) );
  MUX21L U886 ( .A(\gpr[22][9] ), .B(\gpr[23][9] ), .S(n2955), .Z(n2354) );
  MUX21L U887 ( .A(\gpr[20][9] ), .B(\gpr[21][9] ), .S(n2955), .Z(n2353) );
  MUX21L U888 ( .A(\gpr[18][9] ), .B(\gpr[19][9] ), .S(n2955), .Z(n2357) );
  MUX21L U889 ( .A(\gpr[16][9] ), .B(\gpr[17][9] ), .S(n2955), .Z(n2356) );
  MUX31LP U890 ( .D0(n2355), .D1(n2352), .D2(n2348), .A(n2998), .B(n3002), .Z(
        n2372) );
  MUX21L U891 ( .A(\gpr[14][9] ), .B(\gpr[15][9] ), .S(n2955), .Z(n2360) );
  MUX21L U892 ( .A(\gpr[12][9] ), .B(\gpr[13][9] ), .S(n2955), .Z(n2359) );
  MUX21L U893 ( .A(\gpr[10][9] ), .B(\gpr[11][9] ), .S(n2955), .Z(n2363) );
  MUX21L U894 ( .A(\gpr[8][9] ), .B(\gpr[9][9] ), .S(n2955), .Z(n2362) );
  MUX21L U895 ( .A(n2361), .B(n2358), .S(n2998), .Z(n2371) );
  MUX21L U896 ( .A(\gpr[6][9] ), .B(\gpr[7][9] ), .S(n2955), .Z(n2366) );
  MUX21L U897 ( .A(\gpr[4][9] ), .B(\gpr[5][9] ), .S(n2955), .Z(n2365) );
  MUX21L U898 ( .A(\gpr[2][9] ), .B(\gpr[3][9] ), .S(n2956), .Z(n2369) );
  ND2I U899 ( .A(\gpr[1][9] ), .B(n51), .Z(n2368) );
  MUX21L U900 ( .A(n2367), .B(n2364), .S(n43), .Z(n2370) );
  MUX21L U901 ( .A(\gpr[26][10] ), .B(\gpr[27][10] ), .S(n2956), .Z(n2376) );
  MUX21L U902 ( .A(\gpr[24][10] ), .B(\gpr[25][10] ), .S(n2956), .Z(n2375) );
  MUX21L U903 ( .A(\gpr[22][10] ), .B(\gpr[23][10] ), .S(n2956), .Z(n2380) );
  MUX21L U904 ( .A(\gpr[20][10] ), .B(\gpr[21][10] ), .S(n2956), .Z(n2379) );
  MUX21L U905 ( .A(\gpr[18][10] ), .B(\gpr[19][10] ), .S(n2956), .Z(n2383) );
  MUX21L U906 ( .A(\gpr[16][10] ), .B(\gpr[17][10] ), .S(n2956), .Z(n2382) );
  MUX31LP U907 ( .D0(n2381), .D1(n2378), .D2(n2374), .A(n43), .B(n3002), .Z(
        n2398) );
  MUX21L U908 ( .A(\gpr[14][10] ), .B(\gpr[15][10] ), .S(n2956), .Z(n2386) );
  MUX21L U909 ( .A(\gpr[12][10] ), .B(\gpr[13][10] ), .S(n2956), .Z(n2385) );
  MUX21L U910 ( .A(\gpr[10][10] ), .B(\gpr[11][10] ), .S(n2956), .Z(n2389) );
  MUX21L U911 ( .A(\gpr[8][10] ), .B(\gpr[9][10] ), .S(n2956), .Z(n2388) );
  MUX21L U912 ( .A(n2387), .B(n2384), .S(n43), .Z(n2397) );
  MUX21L U913 ( .A(\gpr[6][10] ), .B(\gpr[7][10] ), .S(n2956), .Z(n2392) );
  MUX21L U914 ( .A(\gpr[4][10] ), .B(\gpr[5][10] ), .S(n2957), .Z(n2391) );
  MUX21L U915 ( .A(\gpr[2][10] ), .B(\gpr[3][10] ), .S(n2957), .Z(n2395) );
  ND2I U916 ( .A(\gpr[1][10] ), .B(n51), .Z(n2394) );
  MUX21L U917 ( .A(n2393), .B(n2390), .S(n43), .Z(n2396) );
  MUX21L U918 ( .A(\gpr[26][11] ), .B(\gpr[27][11] ), .S(n2957), .Z(n2402) );
  MUX21L U919 ( .A(\gpr[24][11] ), .B(\gpr[25][11] ), .S(n2957), .Z(n2401) );
  MUX21L U920 ( .A(\gpr[22][11] ), .B(\gpr[23][11] ), .S(n2957), .Z(n2406) );
  MUX21L U921 ( .A(\gpr[20][11] ), .B(\gpr[21][11] ), .S(n2957), .Z(n2405) );
  MUX21L U922 ( .A(\gpr[18][11] ), .B(\gpr[19][11] ), .S(n2957), .Z(n2409) );
  MUX21L U923 ( .A(\gpr[16][11] ), .B(\gpr[17][11] ), .S(n2957), .Z(n2408) );
  MUX31LP U924 ( .D0(n2407), .D1(n2404), .D2(n2400), .A(n43), .B(n3002), .Z(
        n2424) );
  MUX21L U925 ( .A(\gpr[14][11] ), .B(\gpr[15][11] ), .S(n2957), .Z(n2412) );
  MUX21L U926 ( .A(\gpr[12][11] ), .B(\gpr[13][11] ), .S(n2957), .Z(n2411) );
  MUX21L U927 ( .A(\gpr[10][11] ), .B(\gpr[11][11] ), .S(n2957), .Z(n2415) );
  MUX21L U928 ( .A(\gpr[8][11] ), .B(\gpr[9][11] ), .S(n2957), .Z(n2414) );
  MUX21L U929 ( .A(n2413), .B(n2410), .S(n43), .Z(n2423) );
  MUX21L U930 ( .A(\gpr[6][11] ), .B(\gpr[7][11] ), .S(n2957), .Z(n2418) );
  MUX21L U931 ( .A(\gpr[4][11] ), .B(\gpr[5][11] ), .S(n2958), .Z(n2417) );
  MUX21L U932 ( .A(\gpr[2][11] ), .B(\gpr[3][11] ), .S(n2958), .Z(n2421) );
  ND2I U933 ( .A(\gpr[1][11] ), .B(n51), .Z(n2420) );
  MUX21L U934 ( .A(n2419), .B(n2416), .S(n43), .Z(n2422) );
  MUX21L U935 ( .A(\gpr[26][12] ), .B(\gpr[27][12] ), .S(n2958), .Z(n2428) );
  MUX21L U936 ( .A(\gpr[24][12] ), .B(\gpr[25][12] ), .S(n2958), .Z(n2427) );
  MUX21L U937 ( .A(\gpr[22][12] ), .B(\gpr[23][12] ), .S(n2958), .Z(n2432) );
  MUX21L U938 ( .A(\gpr[20][12] ), .B(\gpr[21][12] ), .S(n2958), .Z(n2431) );
  MUX21L U939 ( .A(\gpr[18][12] ), .B(\gpr[19][12] ), .S(n2958), .Z(n2435) );
  MUX21L U940 ( .A(\gpr[16][12] ), .B(\gpr[17][12] ), .S(n2958), .Z(n2434) );
  MUX31LP U941 ( .D0(n2433), .D1(n2430), .D2(n2426), .A(n43), .B(n3002), .Z(
        n2450) );
  MUX21L U942 ( .A(\gpr[14][12] ), .B(\gpr[15][12] ), .S(n2958), .Z(n2438) );
  MUX21L U943 ( .A(\gpr[12][12] ), .B(\gpr[13][12] ), .S(n2958), .Z(n2437) );
  MUX21L U944 ( .A(\gpr[10][12] ), .B(\gpr[11][12] ), .S(n2958), .Z(n2441) );
  MUX21L U945 ( .A(\gpr[8][12] ), .B(\gpr[9][12] ), .S(n2958), .Z(n2440) );
  MUX21L U946 ( .A(n2439), .B(n2436), .S(n43), .Z(n2449) );
  MUX21L U947 ( .A(\gpr[6][12] ), .B(\gpr[7][12] ), .S(n2958), .Z(n2444) );
  MUX21L U948 ( .A(\gpr[4][12] ), .B(\gpr[5][12] ), .S(n2959), .Z(n2443) );
  MUX21L U949 ( .A(\gpr[2][12] ), .B(\gpr[3][12] ), .S(n2959), .Z(n2447) );
  ND2I U950 ( .A(\gpr[1][12] ), .B(n2952), .Z(n2446) );
  MUX21L U951 ( .A(n2445), .B(n2442), .S(n43), .Z(n2448) );
  MUX21L U952 ( .A(\gpr[26][13] ), .B(\gpr[27][13] ), .S(n2959), .Z(n2454) );
  MUX21L U953 ( .A(\gpr[24][13] ), .B(\gpr[25][13] ), .S(n2959), .Z(n2453) );
  MUX21L U954 ( .A(\gpr[22][13] ), .B(\gpr[23][13] ), .S(n2959), .Z(n2458) );
  MUX21L U955 ( .A(\gpr[20][13] ), .B(\gpr[21][13] ), .S(n2959), .Z(n2457) );
  MUX21L U956 ( .A(\gpr[18][13] ), .B(\gpr[19][13] ), .S(n2959), .Z(n2461) );
  MUX21L U957 ( .A(\gpr[16][13] ), .B(\gpr[17][13] ), .S(n2959), .Z(n2460) );
  MUX31LP U958 ( .D0(n2459), .D1(n2456), .D2(n2452), .A(n43), .B(n3002), .Z(
        n2476) );
  MUX21L U959 ( .A(\gpr[14][13] ), .B(\gpr[15][13] ), .S(n2959), .Z(n2464) );
  MUX21L U960 ( .A(\gpr[12][13] ), .B(\gpr[13][13] ), .S(n2959), .Z(n2463) );
  MUX21L U961 ( .A(\gpr[10][13] ), .B(\gpr[11][13] ), .S(n2959), .Z(n2467) );
  MUX21L U962 ( .A(\gpr[8][13] ), .B(\gpr[9][13] ), .S(n2959), .Z(n2466) );
  MUX21L U963 ( .A(n2465), .B(n2462), .S(n43), .Z(n2475) );
  MUX21L U964 ( .A(\gpr[6][13] ), .B(\gpr[7][13] ), .S(n2959), .Z(n2470) );
  MUX21L U965 ( .A(\gpr[4][13] ), .B(\gpr[5][13] ), .S(n2960), .Z(n2469) );
  MUX21L U966 ( .A(\gpr[2][13] ), .B(\gpr[3][13] ), .S(n2960), .Z(n2473) );
  ND2I U967 ( .A(\gpr[1][13] ), .B(n2952), .Z(n2472) );
  MUX21L U968 ( .A(n2471), .B(n2468), .S(n43), .Z(n2474) );
  MUX21L U969 ( .A(\gpr[26][14] ), .B(\gpr[27][14] ), .S(n2960), .Z(n2480) );
  MUX21L U970 ( .A(\gpr[24][14] ), .B(\gpr[25][14] ), .S(n2960), .Z(n2479) );
  MUX21L U971 ( .A(\gpr[22][14] ), .B(\gpr[23][14] ), .S(n2960), .Z(n2484) );
  MUX21L U972 ( .A(\gpr[20][14] ), .B(\gpr[21][14] ), .S(n2956), .Z(n2483) );
  MUX21L U973 ( .A(\gpr[18][14] ), .B(\gpr[19][14] ), .S(n2971), .Z(n2487) );
  MUX21L U974 ( .A(\gpr[16][14] ), .B(\gpr[17][14] ), .S(n2971), .Z(n2486) );
  MUX31LP U975 ( .D0(n2485), .D1(n2482), .D2(n2478), .A(n43), .B(n3002), .Z(
        n2502) );
  MUX21L U976 ( .A(\gpr[14][14] ), .B(\gpr[15][14] ), .S(n2971), .Z(n2490) );
  MUX21L U977 ( .A(\gpr[12][14] ), .B(\gpr[13][14] ), .S(n2971), .Z(n2489) );
  MUX21L U978 ( .A(\gpr[10][14] ), .B(\gpr[11][14] ), .S(n2971), .Z(n2493) );
  MUX21L U979 ( .A(\gpr[8][14] ), .B(\gpr[9][14] ), .S(n2971), .Z(n2492) );
  MUX21L U980 ( .A(n2491), .B(n2488), .S(n43), .Z(n2501) );
  MUX21L U981 ( .A(\gpr[6][14] ), .B(\gpr[7][14] ), .S(n2971), .Z(n2496) );
  MUX21L U982 ( .A(\gpr[4][14] ), .B(\gpr[5][14] ), .S(n2971), .Z(n2495) );
  MUX21L U983 ( .A(\gpr[2][14] ), .B(\gpr[3][14] ), .S(n2971), .Z(n2499) );
  ND2I U984 ( .A(\gpr[1][14] ), .B(n2952), .Z(n2498) );
  MUX21L U985 ( .A(n2497), .B(n2494), .S(n43), .Z(n2500) );
  MUX21L U986 ( .A(\gpr[26][15] ), .B(\gpr[27][15] ), .S(n2971), .Z(n2506) );
  MUX21L U987 ( .A(\gpr[24][15] ), .B(\gpr[25][15] ), .S(n2971), .Z(n2505) );
  MUX21L U988 ( .A(\gpr[22][15] ), .B(\gpr[23][15] ), .S(n2972), .Z(n2510) );
  MUX21L U989 ( .A(\gpr[20][15] ), .B(\gpr[21][15] ), .S(n2972), .Z(n2509) );
  MUX21L U990 ( .A(\gpr[18][15] ), .B(\gpr[19][15] ), .S(n2972), .Z(n2513) );
  MUX21L U991 ( .A(\gpr[16][15] ), .B(\gpr[17][15] ), .S(n2972), .Z(n2512) );
  MUX31LP U992 ( .D0(n2511), .D1(n2508), .D2(n2504), .A(n43), .B(n3002), .Z(
        n2528) );
  MUX21L U993 ( .A(\gpr[14][15] ), .B(\gpr[15][15] ), .S(n2972), .Z(n2516) );
  MUX21L U994 ( .A(\gpr[12][15] ), .B(\gpr[13][15] ), .S(n2972), .Z(n2515) );
  MUX21L U995 ( .A(\gpr[10][15] ), .B(\gpr[11][15] ), .S(n2972), .Z(n2519) );
  MUX21L U996 ( .A(\gpr[8][15] ), .B(\gpr[9][15] ), .S(n2972), .Z(n2518) );
  MUX21L U997 ( .A(n2517), .B(n2514), .S(n43), .Z(n2527) );
  MUX21L U998 ( .A(\gpr[6][15] ), .B(\gpr[7][15] ), .S(n2972), .Z(n2522) );
  MUX21L U999 ( .A(\gpr[4][15] ), .B(\gpr[5][15] ), .S(n2972), .Z(n2521) );
  MUX21L U1000 ( .A(\gpr[2][15] ), .B(\gpr[3][15] ), .S(n2972), .Z(n2525) );
  ND2I U1001 ( .A(\gpr[1][15] ), .B(n2952), .Z(n2524) );
  MUX21L U1002 ( .A(n2523), .B(n2520), .S(n43), .Z(n2526) );
  MUX21L U1003 ( .A(\gpr[26][16] ), .B(\gpr[27][16] ), .S(n2972), .Z(n2532) );
  MUX21L U1004 ( .A(\gpr[24][16] ), .B(\gpr[25][16] ), .S(n2972), .Z(n2531) );
  MUX21L U1005 ( .A(\gpr[22][16] ), .B(\gpr[23][16] ), .S(n2973), .Z(n2536) );
  MUX21L U1006 ( .A(\gpr[20][16] ), .B(\gpr[21][16] ), .S(n2973), .Z(n2535) );
  MUX21L U1007 ( .A(\gpr[18][16] ), .B(\gpr[19][16] ), .S(n2973), .Z(n2539) );
  MUX21L U1008 ( .A(\gpr[16][16] ), .B(\gpr[17][16] ), .S(n2973), .Z(n2538) );
  MUX31LP U1009 ( .D0(n2537), .D1(n2534), .D2(n2530), .A(n120), .B(n3002), .Z(
        n2554) );
  MUX21L U1010 ( .A(\gpr[14][16] ), .B(\gpr[15][16] ), .S(n2973), .Z(n2542) );
  MUX21L U1011 ( .A(\gpr[12][16] ), .B(\gpr[13][16] ), .S(n2973), .Z(n2541) );
  MUX21L U1012 ( .A(\gpr[10][16] ), .B(\gpr[11][16] ), .S(n2973), .Z(n2545) );
  MUX21L U1013 ( .A(\gpr[8][16] ), .B(\gpr[9][16] ), .S(n2973), .Z(n2544) );
  MUX21L U1014 ( .A(n2543), .B(n2540), .S(n120), .Z(n2553) );
  MUX21L U1015 ( .A(\gpr[6][16] ), .B(\gpr[7][16] ), .S(n2973), .Z(n2548) );
  MUX21L U1016 ( .A(\gpr[4][16] ), .B(\gpr[5][16] ), .S(n2973), .Z(n2547) );
  MUX21L U1017 ( .A(\gpr[2][16] ), .B(\gpr[3][16] ), .S(n2973), .Z(n2551) );
  ND2I U1018 ( .A(\gpr[1][16] ), .B(n2952), .Z(n2550) );
  MUX21L U1019 ( .A(n2549), .B(n2546), .S(n120), .Z(n2552) );
  MUX21L U1020 ( .A(\gpr[26][17] ), .B(\gpr[27][17] ), .S(n2973), .Z(n2558) );
  MUX21L U1021 ( .A(\gpr[24][17] ), .B(\gpr[25][17] ), .S(n2973), .Z(n2557) );
  MUX21L U1022 ( .A(\gpr[22][17] ), .B(\gpr[23][17] ), .S(n2974), .Z(n2562) );
  MUX21L U1023 ( .A(\gpr[20][17] ), .B(\gpr[21][17] ), .S(n2974), .Z(n2561) );
  MUX21L U1024 ( .A(\gpr[18][17] ), .B(\gpr[19][17] ), .S(n2974), .Z(n2565) );
  MUX21L U1025 ( .A(\gpr[16][17] ), .B(\gpr[17][17] ), .S(n2974), .Z(n2564) );
  MUX31LP U1026 ( .D0(n2563), .D1(n2560), .D2(n2556), .A(n120), .B(n3002), .Z(
        n2580) );
  MUX21L U1027 ( .A(\gpr[14][17] ), .B(\gpr[15][17] ), .S(n2974), .Z(n2568) );
  MUX21L U1028 ( .A(\gpr[12][17] ), .B(\gpr[13][17] ), .S(n2974), .Z(n2567) );
  MUX21L U1029 ( .A(\gpr[10][17] ), .B(\gpr[11][17] ), .S(n2974), .Z(n2571) );
  MUX21L U1030 ( .A(\gpr[8][17] ), .B(\gpr[9][17] ), .S(n2974), .Z(n2570) );
  MUX21L U1031 ( .A(n2569), .B(n2566), .S(n120), .Z(n2579) );
  MUX21L U1032 ( .A(\gpr[6][17] ), .B(\gpr[7][17] ), .S(n2974), .Z(n2574) );
  MUX21L U1033 ( .A(\gpr[4][17] ), .B(\gpr[5][17] ), .S(n2974), .Z(n2573) );
  MUX21L U1034 ( .A(\gpr[2][17] ), .B(\gpr[3][17] ), .S(n2974), .Z(n2577) );
  ND2I U1035 ( .A(\gpr[1][17] ), .B(n51), .Z(n2576) );
  MUX21L U1036 ( .A(n2575), .B(n2572), .S(n120), .Z(n2578) );
  MUX21L U1037 ( .A(\gpr[26][18] ), .B(\gpr[27][18] ), .S(n2974), .Z(n2584) );
  MUX21L U1038 ( .A(\gpr[24][18] ), .B(\gpr[25][18] ), .S(n2974), .Z(n2583) );
  MUX21L U1039 ( .A(\gpr[22][18] ), .B(\gpr[23][18] ), .S(n2975), .Z(n2588) );
  MUX21L U1040 ( .A(\gpr[20][18] ), .B(\gpr[21][18] ), .S(n2975), .Z(n2587) );
  MUX21L U1041 ( .A(\gpr[18][18] ), .B(\gpr[19][18] ), .S(n2975), .Z(n2591) );
  MUX21L U1042 ( .A(\gpr[16][18] ), .B(\gpr[17][18] ), .S(n2975), .Z(n2590) );
  MUX31LP U1043 ( .D0(n2589), .D1(n2586), .D2(n2582), .A(n120), .B(n3002), .Z(
        n2606) );
  MUX21L U1044 ( .A(\gpr[14][18] ), .B(\gpr[15][18] ), .S(n2975), .Z(n2594) );
  MUX21L U1045 ( .A(\gpr[12][18] ), .B(\gpr[13][18] ), .S(n2975), .Z(n2593) );
  MUX21L U1046 ( .A(\gpr[10][18] ), .B(\gpr[11][18] ), .S(n2975), .Z(n2597) );
  MUX21L U1047 ( .A(\gpr[8][18] ), .B(\gpr[9][18] ), .S(n2975), .Z(n2596) );
  MUX21L U1048 ( .A(n2595), .B(n2592), .S(n120), .Z(n2605) );
  MUX21L U1049 ( .A(\gpr[6][18] ), .B(\gpr[7][18] ), .S(n2975), .Z(n2600) );
  MUX21L U1050 ( .A(\gpr[4][18] ), .B(\gpr[5][18] ), .S(n2975), .Z(n2599) );
  MUX21L U1051 ( .A(\gpr[2][18] ), .B(\gpr[3][18] ), .S(n2975), .Z(n2603) );
  ND2I U1052 ( .A(\gpr[1][18] ), .B(n51), .Z(n2602) );
  MUX21L U1053 ( .A(n2601), .B(n2598), .S(n120), .Z(n2604) );
  MUX21L U1054 ( .A(\gpr[26][19] ), .B(\gpr[27][19] ), .S(n2975), .Z(n2610) );
  MUX21L U1055 ( .A(\gpr[24][19] ), .B(\gpr[25][19] ), .S(n2976), .Z(n2609) );
  MUX21L U1056 ( .A(\gpr[22][19] ), .B(\gpr[23][19] ), .S(n2976), .Z(n2614) );
  MUX21L U1057 ( .A(\gpr[20][19] ), .B(\gpr[21][19] ), .S(n2976), .Z(n2613) );
  MUX21L U1058 ( .A(\gpr[18][19] ), .B(\gpr[19][19] ), .S(n2976), .Z(n2617) );
  MUX21L U1059 ( .A(\gpr[16][19] ), .B(\gpr[17][19] ), .S(n2976), .Z(n2616) );
  MUX31LP U1060 ( .D0(n2615), .D1(n2612), .D2(n2608), .A(n120), .B(n3003), .Z(
        n2632) );
  MUX21L U1061 ( .A(\gpr[14][19] ), .B(\gpr[15][19] ), .S(n2976), .Z(n2620) );
  MUX21L U1062 ( .A(\gpr[12][19] ), .B(\gpr[13][19] ), .S(n2976), .Z(n2619) );
  MUX21L U1063 ( .A(\gpr[10][19] ), .B(\gpr[11][19] ), .S(n2976), .Z(n2623) );
  MUX21L U1064 ( .A(\gpr[8][19] ), .B(\gpr[9][19] ), .S(n2976), .Z(n2622) );
  MUX21L U1065 ( .A(n2621), .B(n2618), .S(n120), .Z(n2631) );
  MUX21L U1066 ( .A(\gpr[6][19] ), .B(\gpr[7][19] ), .S(n2976), .Z(n2626) );
  MUX21L U1067 ( .A(\gpr[4][19] ), .B(\gpr[5][19] ), .S(n2976), .Z(n2625) );
  MUX21L U1068 ( .A(\gpr[2][19] ), .B(\gpr[3][19] ), .S(n2976), .Z(n2629) );
  ND2I U1069 ( .A(\gpr[1][19] ), .B(n51), .Z(n2628) );
  MUX21L U1070 ( .A(n2627), .B(n2624), .S(n120), .Z(n2630) );
  MUX21L U1071 ( .A(\gpr[26][20] ), .B(\gpr[27][20] ), .S(n2976), .Z(n2636) );
  MUX21L U1072 ( .A(\gpr[24][20] ), .B(\gpr[25][20] ), .S(n2977), .Z(n2635) );
  MUX21L U1073 ( .A(\gpr[22][20] ), .B(\gpr[23][20] ), .S(n2977), .Z(n2640) );
  MUX21L U1074 ( .A(\gpr[20][20] ), .B(\gpr[21][20] ), .S(n2977), .Z(n2639) );
  MUX21L U1075 ( .A(\gpr[18][20] ), .B(\gpr[19][20] ), .S(n2977), .Z(n2643) );
  MUX21L U1076 ( .A(\gpr[16][20] ), .B(\gpr[17][20] ), .S(n2977), .Z(n2642) );
  MUX31LP U1077 ( .D0(n2641), .D1(n2638), .D2(n2634), .A(n120), .B(n3003), .Z(
        n2658) );
  MUX21L U1078 ( .A(\gpr[14][20] ), .B(\gpr[15][20] ), .S(n2977), .Z(n2646) );
  MUX21L U1079 ( .A(\gpr[12][20] ), .B(\gpr[13][20] ), .S(n2977), .Z(n2645) );
  MUX21L U1080 ( .A(\gpr[10][20] ), .B(\gpr[11][20] ), .S(n2977), .Z(n2649) );
  MUX21L U1081 ( .A(\gpr[8][20] ), .B(\gpr[9][20] ), .S(n2977), .Z(n2648) );
  MUX21L U1082 ( .A(n2647), .B(n2644), .S(n120), .Z(n2657) );
  MUX21L U1083 ( .A(\gpr[6][20] ), .B(\gpr[7][20] ), .S(n2977), .Z(n2652) );
  MUX21L U1084 ( .A(\gpr[4][20] ), .B(\gpr[5][20] ), .S(n2977), .Z(n2651) );
  MUX21L U1085 ( .A(\gpr[2][20] ), .B(\gpr[3][20] ), .S(n2977), .Z(n2655) );
  ND2I U1086 ( .A(\gpr[1][20] ), .B(n2952), .Z(n2654) );
  MUX21L U1087 ( .A(n2653), .B(n2650), .S(n120), .Z(n2656) );
  MUX21L U1088 ( .A(\gpr[26][21] ), .B(\gpr[27][21] ), .S(n2977), .Z(n2662) );
  MUX21L U1089 ( .A(\gpr[24][21] ), .B(\gpr[25][21] ), .S(n2978), .Z(n2661) );
  MUX21L U1090 ( .A(\gpr[22][21] ), .B(\gpr[23][21] ), .S(n2978), .Z(n2666) );
  MUX21L U1091 ( .A(\gpr[20][21] ), .B(\gpr[21][21] ), .S(n2978), .Z(n2665) );
  MUX21L U1092 ( .A(\gpr[18][21] ), .B(\gpr[19][21] ), .S(n2978), .Z(n2669) );
  MUX21L U1093 ( .A(\gpr[16][21] ), .B(\gpr[17][21] ), .S(n2978), .Z(n2668) );
  MUX31LP U1094 ( .D0(n2667), .D1(n2664), .D2(n2660), .A(n120), .B(n3003), .Z(
        n2684) );
  MUX21L U1095 ( .A(\gpr[14][21] ), .B(\gpr[15][21] ), .S(n2978), .Z(n2672) );
  MUX21L U1096 ( .A(\gpr[12][21] ), .B(\gpr[13][21] ), .S(n2978), .Z(n2671) );
  MUX21L U1097 ( .A(\gpr[10][21] ), .B(\gpr[11][21] ), .S(n2978), .Z(n2675) );
  MUX21L U1098 ( .A(\gpr[8][21] ), .B(\gpr[9][21] ), .S(n2978), .Z(n2674) );
  MUX21L U1099 ( .A(n2673), .B(n2670), .S(n120), .Z(n2683) );
  MUX21L U1100 ( .A(\gpr[6][21] ), .B(\gpr[7][21] ), .S(n2978), .Z(n2678) );
  MUX21L U1101 ( .A(\gpr[4][21] ), .B(\gpr[5][21] ), .S(n2978), .Z(n2677) );
  MUX21L U1102 ( .A(\gpr[2][21] ), .B(\gpr[3][21] ), .S(n2978), .Z(n2681) );
  ND2I U1103 ( .A(\gpr[1][21] ), .B(n2952), .Z(n2680) );
  MUX21L U1104 ( .A(n2679), .B(n2676), .S(n120), .Z(n2682) );
  MUX21L U1105 ( .A(\gpr[26][22] ), .B(\gpr[27][22] ), .S(n2978), .Z(n2688) );
  MUX21L U1106 ( .A(\gpr[24][22] ), .B(\gpr[25][22] ), .S(n2979), .Z(n2687) );
  MUX21L U1107 ( .A(\gpr[22][22] ), .B(\gpr[23][22] ), .S(n2979), .Z(n2692) );
  MUX21L U1108 ( .A(\gpr[20][22] ), .B(\gpr[21][22] ), .S(n2979), .Z(n2691) );
  MUX21L U1109 ( .A(\gpr[18][22] ), .B(\gpr[19][22] ), .S(n2979), .Z(n2695) );
  MUX21L U1110 ( .A(\gpr[16][22] ), .B(\gpr[17][22] ), .S(n2979), .Z(n2694) );
  MUX31LP U1111 ( .D0(n2693), .D1(n2690), .D2(n2686), .A(n120), .B(n3003), .Z(
        n2710) );
  MUX21L U1112 ( .A(\gpr[14][22] ), .B(\gpr[15][22] ), .S(n2979), .Z(n2698) );
  MUX21L U1113 ( .A(\gpr[12][22] ), .B(\gpr[13][22] ), .S(n2979), .Z(n2697) );
  MUX21L U1114 ( .A(\gpr[10][22] ), .B(\gpr[11][22] ), .S(n2979), .Z(n2701) );
  MUX21L U1115 ( .A(\gpr[8][22] ), .B(\gpr[9][22] ), .S(n2979), .Z(n2700) );
  MUX21L U1116 ( .A(n2699), .B(n2696), .S(n2997), .Z(n2709) );
  MUX21L U1117 ( .A(\gpr[6][22] ), .B(\gpr[7][22] ), .S(n2979), .Z(n2704) );
  MUX21L U1118 ( .A(\gpr[4][22] ), .B(\gpr[5][22] ), .S(n2979), .Z(n2703) );
  MUX21L U1119 ( .A(\gpr[2][22] ), .B(\gpr[3][22] ), .S(n2979), .Z(n2707) );
  ND2I U1120 ( .A(\gpr[1][22] ), .B(n2952), .Z(n2706) );
  MUX21L U1121 ( .A(n2705), .B(n2702), .S(n2997), .Z(n2708) );
  MUX21L U1122 ( .A(\gpr[26][23] ), .B(\gpr[27][23] ), .S(n2975), .Z(n2714) );
  MUX21L U1123 ( .A(\gpr[24][23] ), .B(\gpr[25][23] ), .S(n47), .Z(n2713) );
  MUX21L U1124 ( .A(\gpr[22][23] ), .B(\gpr[23][23] ), .S(n47), .Z(n2718) );
  MUX21L U1125 ( .A(\gpr[20][23] ), .B(\gpr[21][23] ), .S(n47), .Z(n2717) );
  MUX21L U1126 ( .A(\gpr[18][23] ), .B(\gpr[19][23] ), .S(n47), .Z(n2721) );
  MUX21L U1127 ( .A(\gpr[16][23] ), .B(\gpr[17][23] ), .S(n47), .Z(n2720) );
  MUX31LP U1128 ( .D0(n2719), .D1(n2716), .D2(n2712), .A(n2997), .B(n3003), 
        .Z(n2736) );
  MUX21L U1129 ( .A(\gpr[14][23] ), .B(\gpr[15][23] ), .S(n47), .Z(n2724) );
  MUX21L U1130 ( .A(\gpr[12][23] ), .B(\gpr[13][23] ), .S(n47), .Z(n2723) );
  MUX21L U1131 ( .A(\gpr[10][23] ), .B(\gpr[11][23] ), .S(n47), .Z(n2727) );
  MUX21L U1132 ( .A(\gpr[8][23] ), .B(\gpr[9][23] ), .S(n47), .Z(n2726) );
  MUX21L U1133 ( .A(n2725), .B(n2722), .S(n2997), .Z(n2735) );
  MUX21L U1134 ( .A(\gpr[6][23] ), .B(\gpr[7][23] ), .S(n47), .Z(n2730) );
  MUX21L U1135 ( .A(\gpr[4][23] ), .B(\gpr[5][23] ), .S(n2968), .Z(n2729) );
  MUX21L U1136 ( .A(\gpr[2][23] ), .B(\gpr[3][23] ), .S(n2968), .Z(n2733) );
  ND2I U1137 ( .A(\gpr[1][23] ), .B(n51), .Z(n2732) );
  MUX21L U1138 ( .A(n2731), .B(n2728), .S(n2997), .Z(n2734) );
  MUX21L U1139 ( .A(\gpr[26][24] ), .B(\gpr[27][24] ), .S(n2968), .Z(n2740) );
  MUX21L U1140 ( .A(\gpr[24][24] ), .B(\gpr[25][24] ), .S(n2968), .Z(n2739) );
  MUX21L U1141 ( .A(\gpr[22][24] ), .B(\gpr[23][24] ), .S(n2968), .Z(n2744) );
  MUX21L U1142 ( .A(\gpr[20][24] ), .B(\gpr[21][24] ), .S(n2968), .Z(n2743) );
  MUX21L U1143 ( .A(\gpr[18][24] ), .B(\gpr[19][24] ), .S(n2968), .Z(n2747) );
  MUX21L U1144 ( .A(\gpr[16][24] ), .B(\gpr[17][24] ), .S(n2968), .Z(n2746) );
  MUX31LP U1145 ( .D0(n2745), .D1(n2742), .D2(n2738), .A(n2997), .B(n3003), 
        .Z(n2762) );
  MUX21L U1146 ( .A(\gpr[14][24] ), .B(\gpr[15][24] ), .S(n2968), .Z(n2750) );
  MUX21L U1147 ( .A(\gpr[12][24] ), .B(\gpr[13][24] ), .S(n2968), .Z(n2749) );
  MUX21L U1148 ( .A(\gpr[10][24] ), .B(\gpr[11][24] ), .S(n2968), .Z(n2753) );
  MUX21L U1149 ( .A(\gpr[8][24] ), .B(\gpr[9][24] ), .S(n2968), .Z(n2752) );
  MUX21L U1150 ( .A(n2751), .B(n2748), .S(n2997), .Z(n2761) );
  MUX21L U1151 ( .A(\gpr[6][24] ), .B(\gpr[7][24] ), .S(n2968), .Z(n2756) );
  MUX21L U1152 ( .A(\gpr[4][24] ), .B(\gpr[5][24] ), .S(n2969), .Z(n2755) );
  MUX21L U1153 ( .A(\gpr[2][24] ), .B(\gpr[3][24] ), .S(n2969), .Z(n2759) );
  ND2I U1154 ( .A(\gpr[1][24] ), .B(n2952), .Z(n2758) );
  MUX21L U1155 ( .A(n2757), .B(n2754), .S(n2997), .Z(n2760) );
  MUX21L U1156 ( .A(\gpr[26][25] ), .B(\gpr[27][25] ), .S(n2969), .Z(n2766) );
  MUX21L U1157 ( .A(\gpr[24][25] ), .B(\gpr[25][25] ), .S(n2969), .Z(n2765) );
  MUX21L U1158 ( .A(\gpr[22][25] ), .B(\gpr[23][25] ), .S(n2969), .Z(n2770) );
  MUX21L U1159 ( .A(\gpr[20][25] ), .B(\gpr[21][25] ), .S(n2969), .Z(n2769) );
  MUX21L U1160 ( .A(\gpr[18][25] ), .B(\gpr[19][25] ), .S(n2969), .Z(n2773) );
  MUX21L U1161 ( .A(\gpr[16][25] ), .B(\gpr[17][25] ), .S(n2969), .Z(n2772) );
  MUX31LP U1162 ( .D0(n2771), .D1(n2768), .D2(n2764), .A(n2997), .B(n3003), 
        .Z(n2788) );
  MUX21L U1163 ( .A(\gpr[14][25] ), .B(\gpr[15][25] ), .S(n2969), .Z(n2776) );
  MUX21L U1164 ( .A(\gpr[12][25] ), .B(\gpr[13][25] ), .S(n2969), .Z(n2775) );
  MUX21L U1165 ( .A(\gpr[10][25] ), .B(\gpr[11][25] ), .S(n2969), .Z(n2779) );
  MUX21L U1166 ( .A(\gpr[8][25] ), .B(\gpr[9][25] ), .S(n2969), .Z(n2778) );
  MUX21L U1167 ( .A(n2777), .B(n2774), .S(n2997), .Z(n2787) );
  MUX21L U1168 ( .A(\gpr[6][25] ), .B(\gpr[7][25] ), .S(n2969), .Z(n2782) );
  MUX21L U1169 ( .A(\gpr[4][25] ), .B(\gpr[5][25] ), .S(n2952), .Z(n2781) );
  MUX21L U1170 ( .A(\gpr[2][25] ), .B(\gpr[3][25] ), .S(n47), .Z(n2785) );
  ND2I U1171 ( .A(\gpr[1][25] ), .B(n51), .Z(n2784) );
  MUX21L U1172 ( .A(n2783), .B(n2780), .S(n2997), .Z(n2786) );
  MUX21L U1173 ( .A(\gpr[26][26] ), .B(\gpr[27][26] ), .S(n2957), .Z(n2792) );
  MUX21L U1174 ( .A(\gpr[24][26] ), .B(\gpr[25][26] ), .S(n2959), .Z(n2791) );
  MUX21L U1175 ( .A(\gpr[22][26] ), .B(\gpr[23][26] ), .S(n2974), .Z(n2796) );
  MUX21L U1176 ( .A(\gpr[20][26] ), .B(\gpr[21][26] ), .S(n2963), .Z(n2795) );
  MUX21L U1177 ( .A(\gpr[18][26] ), .B(\gpr[19][26] ), .S(n2953), .Z(n2799) );
  MUX21L U1178 ( .A(\gpr[16][26] ), .B(\gpr[17][26] ), .S(n47), .Z(n2798) );
  MUX31LP U1179 ( .D0(n2797), .D1(n2794), .D2(n2790), .A(n2997), .B(n3003), 
        .Z(n2814) );
  MUX21L U1180 ( .A(\gpr[14][26] ), .B(\gpr[15][26] ), .S(n2969), .Z(n2802) );
  MUX21L U1181 ( .A(\gpr[12][26] ), .B(\gpr[13][26] ), .S(n2975), .Z(n2801) );
  MUX21L U1182 ( .A(\gpr[10][26] ), .B(\gpr[11][26] ), .S(n2972), .Z(n2805) );
  MUX21L U1183 ( .A(\gpr[8][26] ), .B(\gpr[9][26] ), .S(n2966), .Z(n2804) );
  MUX21L U1184 ( .A(n2803), .B(n2800), .S(n2997), .Z(n2813) );
  MUX21L U1185 ( .A(\gpr[6][26] ), .B(\gpr[7][26] ), .S(n2967), .Z(n2808) );
  MUX21L U1186 ( .A(\gpr[4][26] ), .B(\gpr[5][26] ), .S(n2974), .Z(n2807) );
  MUX21L U1187 ( .A(\gpr[2][26] ), .B(\gpr[3][26] ), .S(n47), .Z(n2811) );
  ND2I U1188 ( .A(\gpr[1][26] ), .B(n51), .Z(n2810) );
  MUX21L U1189 ( .A(n2809), .B(n2806), .S(n2997), .Z(n2812) );
  MUX21L U1190 ( .A(\gpr[26][27] ), .B(\gpr[27][27] ), .S(n2955), .Z(n2818) );
  MUX21L U1191 ( .A(\gpr[24][27] ), .B(\gpr[25][27] ), .S(n2956), .Z(n2817) );
  MUX21L U1192 ( .A(\gpr[22][27] ), .B(\gpr[23][27] ), .S(n2969), .Z(n2822) );
  MUX21L U1193 ( .A(\gpr[20][27] ), .B(\gpr[21][27] ), .S(n47), .Z(n2821) );
  MUX21L U1194 ( .A(\gpr[18][27] ), .B(\gpr[19][27] ), .S(n2969), .Z(n2825) );
  MUX21L U1195 ( .A(\gpr[16][27] ), .B(\gpr[17][27] ), .S(n51), .Z(n2824) );
  MUX31LP U1196 ( .D0(n2823), .D1(n2820), .D2(n2816), .A(n2997), .B(n3003), 
        .Z(n2840) );
  MUX21L U1197 ( .A(\gpr[14][27] ), .B(\gpr[15][27] ), .S(n2963), .Z(n2828) );
  MUX21L U1198 ( .A(\gpr[12][27] ), .B(\gpr[13][27] ), .S(n2953), .Z(n2827) );
  MUX21L U1199 ( .A(\gpr[10][27] ), .B(\gpr[11][27] ), .S(n2976), .Z(n2831) );
  MUX21L U1200 ( .A(\gpr[8][27] ), .B(\gpr[9][27] ), .S(n2973), .Z(n2830) );
  MUX21L U1201 ( .A(n2829), .B(n2826), .S(n2997), .Z(n2839) );
  MUX21L U1202 ( .A(\gpr[6][27] ), .B(\gpr[7][27] ), .S(n51), .Z(n2834) );
  MUX21L U1203 ( .A(\gpr[4][27] ), .B(\gpr[5][27] ), .S(n2966), .Z(n2833) );
  MUX21L U1204 ( .A(\gpr[2][27] ), .B(\gpr[3][27] ), .S(n2967), .Z(n2837) );
  ND2I U1205 ( .A(\gpr[1][27] ), .B(n51), .Z(n2836) );
  MUX21L U1206 ( .A(n2835), .B(n2832), .S(n2997), .Z(n2838) );
  MUX21L U1207 ( .A(\gpr[26][28] ), .B(\gpr[27][28] ), .S(n51), .Z(n2844) );
  MUX21L U1208 ( .A(\gpr[24][28] ), .B(\gpr[25][28] ), .S(n2963), .Z(n2843) );
  MUX21L U1209 ( .A(\gpr[22][28] ), .B(\gpr[23][28] ), .S(n2952), .Z(n2848) );
  MUX21L U1210 ( .A(\gpr[20][28] ), .B(\gpr[21][28] ), .S(n2952), .Z(n2847) );
  MUX21L U1211 ( .A(\gpr[18][28] ), .B(\gpr[19][28] ), .S(n51), .Z(n2851) );
  MUX21L U1212 ( .A(\gpr[16][28] ), .B(\gpr[17][28] ), .S(n2952), .Z(n2850) );
  MUX31LP U1213 ( .D0(n2849), .D1(n2846), .D2(n2842), .A(n2997), .B(n3003), 
        .Z(n2866) );
  MUX21L U1214 ( .A(\gpr[14][28] ), .B(\gpr[15][28] ), .S(n2952), .Z(n2854) );
  MUX21L U1215 ( .A(\gpr[12][28] ), .B(\gpr[13][28] ), .S(n2970), .Z(n2853) );
  MUX21L U1216 ( .A(\gpr[10][28] ), .B(\gpr[11][28] ), .S(n47), .Z(n2857) );
  MUX21L U1217 ( .A(\gpr[8][28] ), .B(\gpr[9][28] ), .S(n51), .Z(n2856) );
  MUX21L U1218 ( .A(n2855), .B(n2852), .S(n2997), .Z(n2865) );
  MUX21L U1219 ( .A(\gpr[6][28] ), .B(\gpr[7][28] ), .S(n2970), .Z(n2860) );
  MUX21L U1220 ( .A(\gpr[4][28] ), .B(\gpr[5][28] ), .S(n2970), .Z(n2859) );
  MUX21L U1221 ( .A(\gpr[2][28] ), .B(\gpr[3][28] ), .S(n2970), .Z(n2863) );
  ND2I U1222 ( .A(\gpr[1][28] ), .B(n2952), .Z(n2862) );
  MUX21L U1223 ( .A(n2861), .B(n2858), .S(n2996), .Z(n2864) );
  MUX21L U1224 ( .A(\gpr[26][29] ), .B(\gpr[27][29] ), .S(n2970), .Z(n2870) );
  MUX21L U1225 ( .A(\gpr[24][29] ), .B(\gpr[25][29] ), .S(n2970), .Z(n2869) );
  MUX21L U1226 ( .A(\gpr[22][29] ), .B(\gpr[23][29] ), .S(n2970), .Z(n2874) );
  MUX21L U1227 ( .A(\gpr[20][29] ), .B(\gpr[21][29] ), .S(n2970), .Z(n2873) );
  MUX21L U1228 ( .A(\gpr[18][29] ), .B(\gpr[19][29] ), .S(n2970), .Z(n2877) );
  MUX21L U1229 ( .A(\gpr[16][29] ), .B(\gpr[17][29] ), .S(n2970), .Z(n2876) );
  MUX31LP U1230 ( .D0(n2875), .D1(n2872), .D2(n2868), .A(n2996), .B(n3003), 
        .Z(n2892) );
  MUX21L U1231 ( .A(\gpr[14][29] ), .B(\gpr[15][29] ), .S(n2970), .Z(n2880) );
  MUX21L U1232 ( .A(\gpr[12][29] ), .B(\gpr[13][29] ), .S(n2970), .Z(n2879) );
  MUX21L U1233 ( .A(\gpr[10][29] ), .B(\gpr[11][29] ), .S(n2970), .Z(n2883) );
  MUX21L U1234 ( .A(\gpr[8][29] ), .B(\gpr[9][29] ), .S(n2970), .Z(n2882) );
  MUX21L U1235 ( .A(n2881), .B(n2878), .S(n2996), .Z(n2891) );
  MUX21L U1236 ( .A(\gpr[6][29] ), .B(\gpr[7][29] ), .S(n25), .Z(n2886) );
  MUX21L U1237 ( .A(\gpr[4][29] ), .B(\gpr[5][29] ), .S(n25), .Z(n2885) );
  MUX21L U1238 ( .A(\gpr[2][29] ), .B(\gpr[3][29] ), .S(n25), .Z(n2889) );
  ND2I U1239 ( .A(\gpr[1][29] ), .B(n2952), .Z(n2888) );
  MUX21L U1240 ( .A(n2887), .B(n2884), .S(n2996), .Z(n2890) );
  MUX21L U1241 ( .A(\gpr[26][30] ), .B(\gpr[27][30] ), .S(n25), .Z(n2896) );
  MUX21L U1242 ( .A(\gpr[24][30] ), .B(\gpr[25][30] ), .S(n25), .Z(n2895) );
  MUX21L U1243 ( .A(\gpr[22][30] ), .B(\gpr[23][30] ), .S(n25), .Z(n2900) );
  MUX21L U1244 ( .A(\gpr[20][30] ), .B(\gpr[21][30] ), .S(n25), .Z(n2899) );
  MUX21L U1245 ( .A(\gpr[18][30] ), .B(\gpr[19][30] ), .S(n25), .Z(n2903) );
  MUX21L U1246 ( .A(\gpr[16][30] ), .B(\gpr[17][30] ), .S(n25), .Z(n2902) );
  MUX31LP U1247 ( .D0(n2901), .D1(n2898), .D2(n2894), .A(n2996), .B(n3003), 
        .Z(n2918) );
  MUX21L U1248 ( .A(\gpr[14][30] ), .B(\gpr[15][30] ), .S(n25), .Z(n2906) );
  MUX21L U1249 ( .A(\gpr[12][30] ), .B(\gpr[13][30] ), .S(n25), .Z(n2905) );
  MUX21L U1250 ( .A(\gpr[10][30] ), .B(\gpr[11][30] ), .S(n25), .Z(n2909) );
  MUX21L U1251 ( .A(\gpr[8][30] ), .B(\gpr[9][30] ), .S(n25), .Z(n2908) );
  MUX21L U1252 ( .A(n2907), .B(n2904), .S(n2996), .Z(n2917) );
  MUX21L U1253 ( .A(\gpr[6][30] ), .B(\gpr[7][30] ), .S(n2967), .Z(n2912) );
  MUX21L U1254 ( .A(\gpr[4][30] ), .B(\gpr[5][30] ), .S(n2970), .Z(n2911) );
  MUX21L U1255 ( .A(\gpr[2][30] ), .B(\gpr[3][30] ), .S(n47), .Z(n2915) );
  ND2I U1256 ( .A(\gpr[1][30] ), .B(n2952), .Z(n2914) );
  MUX21L U1257 ( .A(n2913), .B(n2910), .S(n2996), .Z(n2916) );
  MUX21L U1258 ( .A(\gpr[26][31] ), .B(\gpr[27][31] ), .S(n47), .Z(n2922) );
  MUX21L U1259 ( .A(\gpr[24][31] ), .B(\gpr[25][31] ), .S(n47), .Z(n2921) );
  MUX21L U1260 ( .A(\gpr[22][31] ), .B(\gpr[23][31] ), .S(n47), .Z(n2926) );
  MUX21L U1261 ( .A(\gpr[20][31] ), .B(\gpr[21][31] ), .S(n47), .Z(n2925) );
  MUX21L U1262 ( .A(\gpr[18][31] ), .B(\gpr[19][31] ), .S(n47), .Z(n2929) );
  MUX21L U1263 ( .A(\gpr[16][31] ), .B(\gpr[17][31] ), .S(n47), .Z(n2928) );
  MUX31LP U1264 ( .D0(n2927), .D1(n2924), .D2(n2920), .A(n2996), .B(n3003), 
        .Z(n2944) );
  MUX21L U1265 ( .A(\gpr[14][31] ), .B(\gpr[15][31] ), .S(n2963), .Z(n2932) );
  MUX21L U1266 ( .A(\gpr[12][31] ), .B(\gpr[13][31] ), .S(n47), .Z(n2931) );
  MUX21L U1267 ( .A(\gpr[10][31] ), .B(\gpr[11][31] ), .S(n2952), .Z(n2935) );
  MUX21L U1268 ( .A(\gpr[8][31] ), .B(\gpr[9][31] ), .S(n2963), .Z(n2934) );
  MUX21L U1269 ( .A(n2933), .B(n2930), .S(n2996), .Z(n2943) );
  MUX21L U1270 ( .A(\gpr[6][31] ), .B(\gpr[7][31] ), .S(n2971), .Z(n2938) );
  MUX21L U1271 ( .A(\gpr[4][31] ), .B(\gpr[5][31] ), .S(n2971), .Z(n2937) );
  MUX21L U1272 ( .A(\gpr[2][31] ), .B(\gpr[3][31] ), .S(n2958), .Z(n2941) );
  ND2I U1273 ( .A(\gpr[1][31] ), .B(n2952), .Z(n2940) );
  MUX21L U1274 ( .A(n2939), .B(n2936), .S(n2996), .Z(n2942) );
  IVI U1275 ( .A(n2945), .Z(n2946) );
  IVI U1276 ( .A(n2945), .Z(n2947) );
  IVI U1277 ( .A(n40), .Z(n2948) );
  IVI U1278 ( .A(n2946), .Z(n2949) );
  IVI U1279 ( .A(n2946), .Z(n2950) );
  IVI U1280 ( .A(n2947), .Z(n2951) );
  IVI U1281 ( .A(n3147), .Z(n2980) );
  IVI U1282 ( .A(n2980), .Z(n2981) );
  IVI U1283 ( .A(n2980), .Z(n2982) );
  IVI U1284 ( .A(n2982), .Z(n2983) );
  IVI U1285 ( .A(N20), .Z(n2994) );
  IVI U1286 ( .A(n2994), .Z(n2995) );
  IVI U1287 ( .A(n52), .Z(n3000) );
  B4IP U1288 ( .A(n2982), .Z(n2984) );
  B4IP U1289 ( .A(n2982), .Z(n2985) );
  B4IP U1290 ( .A(n38), .Z(n2990) );
  B4IP U1291 ( .A(n2981), .Z(n2991) );
  B4IP U1292 ( .A(n119), .Z(n2997) );
  B4IP U1293 ( .A(n42), .Z(n2998) );
  B4IP U1294 ( .A(n121), .Z(n3004) );
  IVI U1295 ( .A(n2100), .Z(n3005) );
  MUX21H U1296 ( .A(n128), .B(n59), .S(n2084), .Z(n3006) );
  B4IP U1297 ( .A(n3279), .Z(n3145) );
  B4IP U1298 ( .A(n2030), .Z(n3193) );
  B4IP U1299 ( .A(n3201), .Z(n3198) );
  B4IP U1300 ( .A(n1), .Z(n3199) );
  B4IP U1301 ( .A(n2073), .Z(n3200) );
  IVI U1302 ( .A(n1153), .Z(n3009) );
  IVI U1303 ( .A(n1154), .Z(n3012) );
  IVI U1304 ( .A(n1155), .Z(n3015) );
  IVI U1305 ( .A(n1156), .Z(n3018) );
  IVI U1306 ( .A(n1157), .Z(n3021) );
  IVI U1307 ( .A(n1158), .Z(n3024) );
  IVI U1308 ( .A(n92), .Z(n3027) );
  IVI U1309 ( .A(n73), .Z(n3029) );
  IVI U1310 ( .A(n3226), .Z(n3031) );
  IVI U1311 ( .A(n3232), .Z(n3033) );
  IVI U1312 ( .A(n3235), .Z(n3035) );
  IVI U1313 ( .A(n3238), .Z(n3037) );
  IVI U1314 ( .A(n3241), .Z(n3039) );
  IVI U1315 ( .A(n3244), .Z(n3041) );
  IVI U1316 ( .A(n75), .Z(n3043) );
  IVI U1317 ( .A(n93), .Z(n3046) );
  IVI U1318 ( .A(n3249), .Z(n3049) );
  IVI U1319 ( .A(n3251), .Z(n3052) );
  IVI U1320 ( .A(n3252), .Z(n3055) );
  IVI U1321 ( .A(n3253), .Z(n3058) );
  IVI U1322 ( .A(n3255), .Z(n3061) );
  IVI U1323 ( .A(n3256), .Z(n3064) );
  IVI U1324 ( .A(n3258), .Z(n3067) );
  IVI U1325 ( .A(n94), .Z(n3070) );
  IVI U1326 ( .A(n3260), .Z(n3073) );
  IVI U1327 ( .A(n3263), .Z(n3076) );
  IVI U1328 ( .A(n3265), .Z(n3079) );
  IVI U1329 ( .A(n3266), .Z(n3082) );
  IVI U1330 ( .A(n3268), .Z(n3085) );
  IVI U1331 ( .A(n3269), .Z(n3088) );
  IVI U1332 ( .A(wr_data[22]), .Z(n3120) );
  IVI U1333 ( .A(n3274), .Z(n3132) );
  IVI U1334 ( .A(n4447), .Z(n3136) );
  IVI U1335 ( .A(n4447), .Z(n3137) );
  IVI U1336 ( .A(n4447), .Z(n3138) );
  IVI U1337 ( .A(n4455), .Z(n3139) );
  IVI U1338 ( .A(n4455), .Z(n3140) );
  IVI U1339 ( .A(n4455), .Z(n3141) );
  IVI U1340 ( .A(n4459), .Z(n3142) );
  IVI U1341 ( .A(n4459), .Z(n3143) );
  IVI U1342 ( .A(n4459), .Z(n3144) );
  IVI U1343 ( .A(N19), .Z(n3147) );
  IVI U1344 ( .A(n3152), .Z(n3148) );
  IVI U1345 ( .A(n3151), .Z(n3150) );
  IVI U1346 ( .A(N13), .Z(n3151) );
  IVI U1347 ( .A(N13), .Z(n3152) );
  IVI U1348 ( .A(n3148), .Z(n3182) );
  IVI U1349 ( .A(n2089), .Z(n3183) );
  IVI U1350 ( .A(n2089), .Z(n3185) );
  IVI U1351 ( .A(n2031), .Z(n3186) );
  IVI U1352 ( .A(n3150), .Z(n3187) );
  IVI U1353 ( .A(n2089), .Z(n3188) );
  IVI U1354 ( .A(n3204), .Z(n3203) );
  IVI U1355 ( .A(N14), .Z(n3204) );
  IVI U1356 ( .A(n3207), .Z(n3205) );
  IVI U1357 ( .A(n3207), .Z(n3206) );
  IVI U1358 ( .A(N15), .Z(n3207) );
  IVI U1359 ( .A(n3205), .Z(n3212) );
  IVI U1360 ( .A(n3205), .Z(n3214) );
  IVI U1361 ( .A(wr_addr[3]), .Z(n3248) );
  IVI U1362 ( .A(wr_addr[4]), .Z(n3221) );
  ND3 U1363 ( .A(RegWrite), .B(n3248), .C(n3221), .Z(n3215) );
  IVI U1364 ( .A(n3215), .Z(n3220) );
  IVI U1365 ( .A(wr_addr[1]), .Z(n3224) );
  IVI U1366 ( .A(wr_addr[2]), .Z(n3223) );
  MUX21L U1367 ( .A(n1159), .B(n3089), .S(n3009), .Z(n1108) );
  MUX21L U1368 ( .A(n1160), .B(n3091), .S(n3009), .Z(n1109) );
  MUX21L U1369 ( .A(n142), .B(n3093), .S(n3009), .Z(n1110) );
  MUX21L U1370 ( .A(n1180), .B(n3095), .S(n3009), .Z(n1111) );
  MUX21L U1371 ( .A(n3216), .B(n3098), .S(n3008), .Z(n1112) );
  MUX21L U1372 ( .A(n5), .B(n3099), .S(n3008), .Z(n1113) );
  MUX21L U1373 ( .A(n3217), .B(n3100), .S(n3008), .Z(n1114) );
  MUX21L U1374 ( .A(n1181), .B(n3101), .S(n3008), .Z(n1115) );
  MUX21L U1375 ( .A(n4), .B(n3102), .S(n3008), .Z(n1116) );
  MUX21L U1376 ( .A(n1182), .B(n3103), .S(n3008), .Z(n1117) );
  MUX21L U1377 ( .A(n1183), .B(n3104), .S(n3008), .Z(n1118) );
  MUX21L U1378 ( .A(n3), .B(n3105), .S(n3008), .Z(n1119) );
  MUX21L U1379 ( .A(n1184), .B(n3106), .S(n3008), .Z(n1120) );
  MUX21L U1380 ( .A(n19), .B(n3107), .S(n3008), .Z(n1121) );
  MUX21L U1381 ( .A(n1185), .B(n3108), .S(n3008), .Z(n1122) );
  MUX21L U1382 ( .A(n18), .B(n3110), .S(n3008), .Z(n1123) );
  MUX21L U1383 ( .A(n17), .B(n3112), .S(n3008), .Z(n1124) );
  MUX21L U1384 ( .A(n16), .B(n3113), .S(n3008), .Z(n1125) );
  MUX21L U1385 ( .A(n1186), .B(n3114), .S(n3007), .Z(n1126) );
  MUX21L U1386 ( .A(n15), .B(n3115), .S(n3007), .Z(n1127) );
  MUX21L U1387 ( .A(n1187), .B(n3116), .S(n3007), .Z(n1128) );
  MUX21L U1388 ( .A(n14), .B(n3117), .S(n3007), .Z(n1129) );
  MUX21L U1389 ( .A(n1188), .B(n3120), .S(n3007), .Z(n1130) );
  MUX21L U1390 ( .A(n13), .B(n3121), .S(n3007), .Z(n1131) );
  MUX21L U1391 ( .A(n12), .B(n3122), .S(n3007), .Z(n1132) );
  MUX21L U1392 ( .A(n11), .B(n3123), .S(n3007), .Z(n1133) );
  MUX21L U1393 ( .A(n1189), .B(n3124), .S(n3007), .Z(n1134) );
  MUX21L U1394 ( .A(n10), .B(n3125), .S(n3007), .Z(n1135) );
  MUX21L U1395 ( .A(n9), .B(n3126), .S(n3007), .Z(n1136) );
  MUX21L U1396 ( .A(n8), .B(n3127), .S(n3007), .Z(n1137) );
  MUX21L U1397 ( .A(n7), .B(n3129), .S(n3007), .Z(n1138) );
  MUX21L U1398 ( .A(n6), .B(n3133), .S(n3007), .Z(n1139) );
  IVI U1399 ( .A(wr_addr[0]), .Z(n3222) );
  MUX21L U1400 ( .A(n147), .B(n3090), .S(n3012), .Z(n1076) );
  MUX21L U1401 ( .A(n1140), .B(n3092), .S(n3012), .Z(n1077) );
  MUX21L U1402 ( .A(n140), .B(n3094), .S(n3012), .Z(n1078) );
  MUX21L U1403 ( .A(n1190), .B(n3096), .S(n3012), .Z(n1079) );
  MUX21L U1404 ( .A(n1191), .B(n3097), .S(n3011), .Z(n1080) );
  MUX21L U1405 ( .A(n1192), .B(n3099), .S(n3011), .Z(n1081) );
  MUX21L U1406 ( .A(n1193), .B(n3100), .S(n3011), .Z(n1082) );
  MUX21L U1407 ( .A(n1194), .B(n3101), .S(n3011), .Z(n1083) );
  MUX21L U1408 ( .A(n1195), .B(n3102), .S(n3011), .Z(n1084) );
  MUX21L U1409 ( .A(n1196), .B(n3103), .S(n3011), .Z(n1085) );
  MUX21L U1410 ( .A(n1197), .B(n3104), .S(n3011), .Z(n1086) );
  MUX21L U1411 ( .A(n1198), .B(n3105), .S(n3011), .Z(n1087) );
  MUX21L U1412 ( .A(n1199), .B(n3106), .S(n3011), .Z(n1088) );
  MUX21L U1413 ( .A(n1200), .B(n3107), .S(n3011), .Z(n1089) );
  MUX21L U1414 ( .A(n1201), .B(n3109), .S(n3011), .Z(n1090) );
  MUX21L U1415 ( .A(n1202), .B(n3110), .S(n3011), .Z(n1091) );
  MUX21L U1416 ( .A(n1203), .B(n3111), .S(n3011), .Z(n1092) );
  MUX21L U1417 ( .A(n1204), .B(n3113), .S(n3011), .Z(n1093) );
  MUX21L U1418 ( .A(n1205), .B(n3114), .S(n3010), .Z(n1094) );
  MUX21L U1419 ( .A(n1206), .B(n3115), .S(n3010), .Z(n1095) );
  MUX21L U1420 ( .A(n1207), .B(n3116), .S(n3010), .Z(n1096) );
  MUX21L U1421 ( .A(n1208), .B(n3117), .S(n3010), .Z(n1097) );
  MUX21L U1422 ( .A(n1209), .B(n3120), .S(n3010), .Z(n1098) );
  MUX21L U1423 ( .A(n1210), .B(n3121), .S(n3010), .Z(n1099) );
  MUX21L U1424 ( .A(n1211), .B(n3122), .S(n3010), .Z(n1100) );
  MUX21L U1425 ( .A(n1212), .B(n3123), .S(n3010), .Z(n1101) );
  MUX21L U1426 ( .A(n1213), .B(n3124), .S(n3010), .Z(n1102) );
  MUX21L U1427 ( .A(n1214), .B(n3125), .S(n3010), .Z(n1103) );
  MUX21L U1428 ( .A(n1215), .B(n3126), .S(n3010), .Z(n1104) );
  MUX21L U1429 ( .A(n1216), .B(n3128), .S(n3010), .Z(n1105) );
  MUX21L U1430 ( .A(n1217), .B(n3129), .S(n3010), .Z(n1106) );
  MUX21L U1431 ( .A(n1218), .B(n3133), .S(n3010), .Z(n1107) );
  MUX21L U1432 ( .A(n81), .B(n3089), .S(n3015), .Z(n1044) );
  MUX21L U1433 ( .A(n82), .B(n3091), .S(n3015), .Z(n1045) );
  MUX21L U1434 ( .A(n71), .B(n3093), .S(n3015), .Z(n1046) );
  MUX21L U1435 ( .A(n1219), .B(n3095), .S(n3015), .Z(n1047) );
  MUX21L U1436 ( .A(n1220), .B(n3098), .S(n3014), .Z(n1048) );
  MUX21L U1437 ( .A(n1221), .B(n3099), .S(n3014), .Z(n1049) );
  MUX21L U1438 ( .A(n1222), .B(n3100), .S(n3014), .Z(n1050) );
  MUX21L U1439 ( .A(n1223), .B(n3101), .S(n3014), .Z(n1051) );
  MUX21L U1440 ( .A(n1224), .B(n3102), .S(n3014), .Z(n1052) );
  MUX21L U1441 ( .A(n1225), .B(n3103), .S(n3014), .Z(n1053) );
  MUX21L U1442 ( .A(n1226), .B(n3104), .S(n3014), .Z(n1054) );
  MUX21L U1443 ( .A(n1227), .B(n3105), .S(n3014), .Z(n1055) );
  MUX21L U1444 ( .A(n1228), .B(n3106), .S(n3014), .Z(n1056) );
  MUX21L U1445 ( .A(n1229), .B(n3107), .S(n3014), .Z(n1057) );
  MUX21L U1446 ( .A(n1230), .B(n3108), .S(n3014), .Z(n1058) );
  MUX21L U1447 ( .A(n1231), .B(n3110), .S(n3014), .Z(n1059) );
  MUX21L U1448 ( .A(n1232), .B(n3112), .S(n3014), .Z(n1060) );
  MUX21L U1449 ( .A(n1233), .B(n3113), .S(n3014), .Z(n1061) );
  MUX21L U1450 ( .A(n1234), .B(n3114), .S(n3013), .Z(n1062) );
  MUX21L U1451 ( .A(n1235), .B(n3115), .S(n3013), .Z(n1063) );
  MUX21L U1452 ( .A(n1236), .B(n3116), .S(n3013), .Z(n1064) );
  MUX21L U1453 ( .A(n1237), .B(n3117), .S(n3013), .Z(n1065) );
  MUX21L U1454 ( .A(n1238), .B(n3120), .S(n3013), .Z(n1066) );
  MUX21L U1455 ( .A(n1239), .B(n3121), .S(n3013), .Z(n1067) );
  MUX21L U1456 ( .A(n1240), .B(n3122), .S(n3013), .Z(n1068) );
  MUX21L U1457 ( .A(n1241), .B(n3123), .S(n3013), .Z(n1069) );
  MUX21L U1458 ( .A(n1242), .B(n3124), .S(n3013), .Z(n1070) );
  MUX21L U1459 ( .A(n1243), .B(n3125), .S(n3013), .Z(n1071) );
  MUX21L U1460 ( .A(n1244), .B(n3126), .S(n3013), .Z(n1072) );
  MUX21L U1461 ( .A(n1245), .B(n3127), .S(n3013), .Z(n1073) );
  MUX21L U1462 ( .A(n1246), .B(n3129), .S(n3013), .Z(n1074) );
  MUX21L U1463 ( .A(n1247), .B(n3133), .S(n3013), .Z(n1075) );
  MUX21L U1464 ( .A(n77), .B(n3090), .S(n3018), .Z(n1012) );
  MUX21L U1465 ( .A(n78), .B(n3092), .S(n3018), .Z(n1013) );
  MUX21L U1466 ( .A(n60), .B(n3094), .S(n3018), .Z(n1014) );
  MUX21L U1467 ( .A(n1161), .B(n3096), .S(n3018), .Z(n1015) );
  MUX21L U1468 ( .A(n141), .B(n3098), .S(n3017), .Z(n1016) );
  MUX21L U1469 ( .A(n1141), .B(n3099), .S(n3017), .Z(n1017) );
  MUX21L U1470 ( .A(n1162), .B(n3100), .S(n3017), .Z(n1018) );
  MUX21L U1471 ( .A(n1163), .B(n3101), .S(n3017), .Z(n1019) );
  MUX21L U1472 ( .A(n1142), .B(n3102), .S(n3017), .Z(n1020) );
  MUX21L U1473 ( .A(n1143), .B(n3103), .S(n3017), .Z(n1021) );
  MUX21L U1474 ( .A(n1144), .B(n3104), .S(n3017), .Z(n1022) );
  MUX21L U1475 ( .A(n1164), .B(n3105), .S(n3017), .Z(n1023) );
  MUX21L U1476 ( .A(n1165), .B(n3106), .S(n3017), .Z(n1024) );
  MUX21L U1477 ( .A(n1145), .B(n3107), .S(n3017), .Z(n1025) );
  MUX21L U1478 ( .A(n1146), .B(n3109), .S(n3017), .Z(n1026) );
  MUX21L U1479 ( .A(n1147), .B(n3110), .S(n3017), .Z(n1027) );
  MUX21L U1480 ( .A(n1148), .B(n3112), .S(n3017), .Z(n1028) );
  MUX21L U1481 ( .A(n1166), .B(n3113), .S(n3017), .Z(n1029) );
  MUX21L U1482 ( .A(n1167), .B(n3114), .S(n3016), .Z(n1030) );
  MUX21L U1483 ( .A(n1149), .B(n3115), .S(n3016), .Z(n1031) );
  MUX21L U1484 ( .A(n1168), .B(n3116), .S(n3016), .Z(n1032) );
  MUX21L U1485 ( .A(n1150), .B(n3117), .S(n3016), .Z(n1033) );
  MUX21L U1486 ( .A(n1169), .B(n3119), .S(n3016), .Z(n1034) );
  MUX21L U1487 ( .A(n1151), .B(n3121), .S(n3016), .Z(n1035) );
  MUX21L U1488 ( .A(n1170), .B(n3122), .S(n3016), .Z(n1036) );
  MUX21L U1489 ( .A(n1171), .B(n3123), .S(n3016), .Z(n1037) );
  MUX21L U1490 ( .A(n1152), .B(n3124), .S(n3016), .Z(n1038) );
  MUX21L U1491 ( .A(n1172), .B(n3125), .S(n3016), .Z(n1039) );
  MUX21L U1492 ( .A(n1173), .B(n3126), .S(n3016), .Z(n1040) );
  MUX21L U1493 ( .A(n1174), .B(n3128), .S(n3016), .Z(n1041) );
  MUX21L U1494 ( .A(n1175), .B(n3129), .S(n3016), .Z(n1042) );
  MUX21L U1495 ( .A(n1176), .B(n3133), .S(n3016), .Z(n1043) );
  MUX21L U1496 ( .A(n143), .B(n3090), .S(n3021), .Z(n980) );
  MUX21L U1497 ( .A(n144), .B(n3092), .S(n3021), .Z(n981) );
  MUX21L U1498 ( .A(n129), .B(n3094), .S(n3021), .Z(n982) );
  MUX21L U1499 ( .A(n95), .B(n3096), .S(n3021), .Z(n983) );
  MUX21L U1500 ( .A(n72), .B(n3098), .S(n3020), .Z(n984) );
  MUX21L U1501 ( .A(n83), .B(n3099), .S(n3020), .Z(n985) );
  MUX21L U1502 ( .A(n96), .B(n3100), .S(n3020), .Z(n986) );
  MUX21L U1503 ( .A(n97), .B(n3101), .S(n3020), .Z(n987) );
  MUX21L U1504 ( .A(n98), .B(n3102), .S(n3020), .Z(n988) );
  MUX21L U1505 ( .A(n84), .B(n3103), .S(n3020), .Z(n989) );
  MUX21L U1506 ( .A(n99), .B(n3104), .S(n3020), .Z(n990) );
  MUX21L U1507 ( .A(n100), .B(n3105), .S(n3020), .Z(n991) );
  MUX21L U1508 ( .A(n101), .B(n3106), .S(n3020), .Z(n992) );
  MUX21L U1509 ( .A(n85), .B(n3107), .S(n3020), .Z(n993) );
  MUX21L U1510 ( .A(n86), .B(n3109), .S(n3020), .Z(n994) );
  MUX21L U1511 ( .A(n102), .B(n3110), .S(n3020), .Z(n995) );
  MUX21L U1512 ( .A(n87), .B(n3112), .S(n3020), .Z(n996) );
  MUX21L U1513 ( .A(n103), .B(n3113), .S(n3020), .Z(n997) );
  MUX21L U1514 ( .A(n104), .B(n3114), .S(n3019), .Z(n998) );
  MUX21L U1515 ( .A(n88), .B(n3115), .S(n3019), .Z(n999) );
  MUX21L U1516 ( .A(n105), .B(n3116), .S(n3019), .Z(n1000) );
  MUX21L U1517 ( .A(n89), .B(n3117), .S(n3019), .Z(n1001) );
  MUX21L U1518 ( .A(n106), .B(n3119), .S(n3019), .Z(n1002) );
  MUX21L U1519 ( .A(n90), .B(n3121), .S(n3019), .Z(n1003) );
  MUX21L U1520 ( .A(n107), .B(n3122), .S(n3019), .Z(n1004) );
  MUX21L U1521 ( .A(n108), .B(n3123), .S(n3019), .Z(n1005) );
  MUX21L U1522 ( .A(n91), .B(n3124), .S(n3019), .Z(n1006) );
  MUX21L U1523 ( .A(n109), .B(n3125), .S(n3019), .Z(n1007) );
  MUX21L U1524 ( .A(n110), .B(n3126), .S(n3019), .Z(n1008) );
  MUX21L U1525 ( .A(n111), .B(n3128), .S(n3019), .Z(n1009) );
  MUX21L U1526 ( .A(n112), .B(n3129), .S(n3019), .Z(n1010) );
  MUX21L U1527 ( .A(n113), .B(n3133), .S(n3019), .Z(n1011) );
  ND2I U1528 ( .A(wr_addr[2]), .B(wr_addr[1]), .Z(n3218) );
  IVI U1529 ( .A(n3218), .Z(n3219) );
  MUX21L U1530 ( .A(n1248), .B(n3090), .S(n3024), .Z(n948) );
  MUX21L U1531 ( .A(n1249), .B(n3092), .S(n3024), .Z(n949) );
  MUX21L U1532 ( .A(n1250), .B(n3094), .S(n3024), .Z(n950) );
  MUX21L U1533 ( .A(n1251), .B(n3096), .S(n3024), .Z(n951) );
  MUX21L U1534 ( .A(n1252), .B(n3098), .S(n3023), .Z(n952) );
  MUX21L U1535 ( .A(n1253), .B(n3099), .S(n3023), .Z(n953) );
  MUX21L U1536 ( .A(n1254), .B(n3100), .S(n3023), .Z(n954) );
  MUX21L U1537 ( .A(n1178), .B(n3101), .S(n3023), .Z(n955) );
  MUX21L U1538 ( .A(n1255), .B(n3102), .S(n3023), .Z(n956) );
  MUX21L U1539 ( .A(n1256), .B(n3103), .S(n3023), .Z(n957) );
  MUX21L U1540 ( .A(n1257), .B(n3104), .S(n3023), .Z(n958) );
  MUX21L U1541 ( .A(n1258), .B(n3105), .S(n3023), .Z(n959) );
  MUX21L U1542 ( .A(n1259), .B(n3106), .S(n3023), .Z(n960) );
  MUX21L U1543 ( .A(n1260), .B(n3107), .S(n3023), .Z(n961) );
  MUX21L U1544 ( .A(n1261), .B(n3109), .S(n3023), .Z(n962) );
  MUX21L U1545 ( .A(n1262), .B(n3110), .S(n3023), .Z(n963) );
  MUX21L U1546 ( .A(n1263), .B(n3112), .S(n3023), .Z(n964) );
  MUX21L U1547 ( .A(n1264), .B(n3113), .S(n3023), .Z(n965) );
  MUX21L U1548 ( .A(n1265), .B(n3114), .S(n3022), .Z(n966) );
  MUX21L U1549 ( .A(n1266), .B(n3115), .S(n3022), .Z(n967) );
  MUX21L U1550 ( .A(n1267), .B(n3116), .S(n3022), .Z(n968) );
  MUX21L U1551 ( .A(n1268), .B(n3117), .S(n3022), .Z(n969) );
  MUX21L U1552 ( .A(n1269), .B(n3119), .S(n3022), .Z(n970) );
  MUX21L U1553 ( .A(n1270), .B(n3121), .S(n3022), .Z(n971) );
  MUX21L U1554 ( .A(n1271), .B(n3122), .S(n3022), .Z(n972) );
  MUX21L U1555 ( .A(n1272), .B(n3123), .S(n3022), .Z(n973) );
  MUX21L U1556 ( .A(n1273), .B(n3124), .S(n3022), .Z(n974) );
  MUX21L U1557 ( .A(n1274), .B(n3125), .S(n3022), .Z(n975) );
  MUX21L U1558 ( .A(n1275), .B(n3126), .S(n3022), .Z(n976) );
  MUX21L U1559 ( .A(n1276), .B(n3128), .S(n3022), .Z(n977) );
  MUX21L U1560 ( .A(n1277), .B(n3129), .S(n3022), .Z(n978) );
  MUX21L U1561 ( .A(n1278), .B(n3133), .S(n3022), .Z(n979) );
  MUX21L U1562 ( .A(n1279), .B(n3090), .S(n3027), .Z(n916) );
  MUX21L U1563 ( .A(n1280), .B(n3092), .S(n3027), .Z(n917) );
  MUX21L U1564 ( .A(n1281), .B(n3094), .S(n3027), .Z(n918) );
  MUX21L U1565 ( .A(n1282), .B(n3096), .S(n3027), .Z(n919) );
  MUX21L U1566 ( .A(n1283), .B(n3098), .S(n3026), .Z(n920) );
  MUX21L U1567 ( .A(n1284), .B(n3099), .S(n3026), .Z(n921) );
  MUX21L U1568 ( .A(n1285), .B(n3100), .S(n3026), .Z(n922) );
  MUX21L U1569 ( .A(n114), .B(n3101), .S(n3026), .Z(n923) );
  MUX21L U1570 ( .A(n1286), .B(n3102), .S(n3026), .Z(n924) );
  MUX21L U1571 ( .A(n1287), .B(n3103), .S(n3026), .Z(n925) );
  MUX21L U1572 ( .A(n1288), .B(n3104), .S(n3026), .Z(n926) );
  MUX21L U1573 ( .A(n1289), .B(n3105), .S(n3026), .Z(n927) );
  MUX21L U1574 ( .A(n1290), .B(n3106), .S(n3026), .Z(n928) );
  MUX21L U1575 ( .A(n1291), .B(n3107), .S(n3026), .Z(n929) );
  MUX21L U1576 ( .A(n1292), .B(n3109), .S(n3026), .Z(n930) );
  MUX21L U1577 ( .A(n1293), .B(n3110), .S(n3026), .Z(n931) );
  MUX21L U1578 ( .A(n1294), .B(n3112), .S(n3026), .Z(n932) );
  MUX21L U1579 ( .A(n1295), .B(n3113), .S(n3026), .Z(n933) );
  MUX21L U1580 ( .A(n1296), .B(n3114), .S(n3025), .Z(n934) );
  MUX21L U1581 ( .A(n1297), .B(n3115), .S(n3025), .Z(n935) );
  MUX21L U1582 ( .A(n1298), .B(n3116), .S(n3025), .Z(n936) );
  MUX21L U1583 ( .A(n1299), .B(n3117), .S(n3025), .Z(n937) );
  MUX21L U1584 ( .A(n1300), .B(n3119), .S(n3025), .Z(n938) );
  MUX21L U1585 ( .A(n1301), .B(n3121), .S(n3025), .Z(n939) );
  MUX21L U1586 ( .A(n1302), .B(n3122), .S(n3025), .Z(n940) );
  MUX21L U1587 ( .A(n1303), .B(n3123), .S(n3025), .Z(n941) );
  MUX21L U1588 ( .A(n1304), .B(n3124), .S(n3025), .Z(n942) );
  MUX21L U1589 ( .A(n1305), .B(n3125), .S(n3025), .Z(n943) );
  MUX21L U1590 ( .A(n1306), .B(n3126), .S(n3025), .Z(n944) );
  MUX21L U1591 ( .A(n1307), .B(n3128), .S(n3025), .Z(n945) );
  MUX21L U1592 ( .A(n1308), .B(n3129), .S(n3025), .Z(n946) );
  MUX21L U1593 ( .A(n1309), .B(n3133), .S(n3025), .Z(n947) );
  MUX21L U1594 ( .A(n79), .B(n3090), .S(n3029), .Z(n884) );
  MUX21L U1595 ( .A(n80), .B(n3092), .S(n3029), .Z(n885) );
  MUX21L U1596 ( .A(n61), .B(n3094), .S(n3029), .Z(n886) );
  MUX21L U1597 ( .A(n1310), .B(n3096), .S(n3029), .Z(n887) );
  MUX21L U1598 ( .A(n1311), .B(n3098), .S(n3028), .Z(n888) );
  MUX21L U1599 ( .A(n1312), .B(n3099), .S(n3028), .Z(n889) );
  MUX21L U1600 ( .A(n3225), .B(n3100), .S(n3028), .Z(n890) );
  MUX21L U1601 ( .A(n1313), .B(n3101), .S(n3028), .Z(n891) );
  MUX21L U1602 ( .A(n1314), .B(n3102), .S(n3028), .Z(n892) );
  MUX21L U1603 ( .A(n1315), .B(n3103), .S(n3028), .Z(n893) );
  MUX21L U1604 ( .A(n1316), .B(n3104), .S(n3028), .Z(n894) );
  MUX21L U1605 ( .A(n1317), .B(n3105), .S(n3028), .Z(n895) );
  MUX21L U1606 ( .A(n1318), .B(n3106), .S(n3028), .Z(n896) );
  MUX21L U1607 ( .A(n1319), .B(n3107), .S(n3028), .Z(n897) );
  MUX21L U1608 ( .A(n1320), .B(n3109), .S(n3028), .Z(n898) );
  MUX21L U1609 ( .A(n1321), .B(n3110), .S(n3028), .Z(n899) );
  MUX21L U1610 ( .A(n1322), .B(n3112), .S(n3028), .Z(n900) );
  MUX21L U1611 ( .A(n1323), .B(n3113), .S(n3028), .Z(n901) );
  MUX21L U1612 ( .A(n1324), .B(n3114), .S(n74), .Z(n902) );
  MUX21L U1613 ( .A(n1325), .B(n3115), .S(n74), .Z(n903) );
  MUX21L U1614 ( .A(n1326), .B(n3116), .S(n74), .Z(n904) );
  MUX21L U1615 ( .A(n1327), .B(n3117), .S(n74), .Z(n905) );
  MUX21L U1616 ( .A(n1328), .B(n3119), .S(n74), .Z(n906) );
  MUX21L U1617 ( .A(n1329), .B(n3121), .S(n74), .Z(n907) );
  MUX21L U1618 ( .A(n1330), .B(n3122), .S(n74), .Z(n908) );
  MUX21L U1619 ( .A(n1331), .B(n3123), .S(n74), .Z(n909) );
  MUX21L U1620 ( .A(n1332), .B(n3124), .S(n74), .Z(n910) );
  MUX21L U1621 ( .A(n1333), .B(n3125), .S(n74), .Z(n911) );
  MUX21L U1622 ( .A(n1334), .B(n3126), .S(n74), .Z(n912) );
  MUX21L U1623 ( .A(n1335), .B(n3128), .S(n74), .Z(n913) );
  MUX21L U1624 ( .A(n1336), .B(n3129), .S(n74), .Z(n914) );
  MUX21L U1625 ( .A(n1337), .B(n3133), .S(n74), .Z(n915) );
  ND2I U1626 ( .A(n2106), .B(n2112), .Z(n3226) );
  IVI U1627 ( .A(n3226), .Z(n3231) );
  MUX21L U1628 ( .A(n145), .B(n3090), .S(n3031), .Z(n852) );
  MUX21L U1629 ( .A(n146), .B(n3092), .S(n3031), .Z(n853) );
  MUX21L U1630 ( .A(n130), .B(n3094), .S(n3031), .Z(n854) );
  MUX21L U1631 ( .A(n1338), .B(n3096), .S(n3031), .Z(n855) );
  MUX21L U1632 ( .A(n3227), .B(n3098), .S(n3030), .Z(n856) );
  MUX21L U1633 ( .A(n3228), .B(n3099), .S(n3030), .Z(n857) );
  MUX21L U1634 ( .A(n3229), .B(n3100), .S(n3030), .Z(n858) );
  MUX21L U1635 ( .A(n1339), .B(n3101), .S(n3030), .Z(n859) );
  MUX21L U1636 ( .A(n1340), .B(n3102), .S(n3030), .Z(n860) );
  MUX21L U1637 ( .A(n3230), .B(n3103), .S(n3030), .Z(n861) );
  MUX21L U1638 ( .A(n1341), .B(n3104), .S(n3030), .Z(n862) );
  MUX21L U1639 ( .A(n1342), .B(n3105), .S(n3030), .Z(n863) );
  MUX21L U1640 ( .A(n1343), .B(n3106), .S(n3030), .Z(n864) );
  MUX21L U1641 ( .A(n1344), .B(n3107), .S(n3030), .Z(n865) );
  MUX21L U1642 ( .A(n1345), .B(n3109), .S(n3030), .Z(n866) );
  MUX21L U1643 ( .A(n1346), .B(n3110), .S(n3030), .Z(n867) );
  MUX21L U1644 ( .A(n1347), .B(n3112), .S(n3030), .Z(n868) );
  MUX21L U1645 ( .A(n1348), .B(n3113), .S(n3030), .Z(n869) );
  MUX21L U1646 ( .A(n1349), .B(n3114), .S(n3231), .Z(n870) );
  MUX21L U1647 ( .A(n1350), .B(n3115), .S(n3030), .Z(n871) );
  MUX21L U1648 ( .A(n1351), .B(n3116), .S(n3030), .Z(n872) );
  MUX21L U1649 ( .A(n1352), .B(n3117), .S(n3031), .Z(n873) );
  MUX21L U1650 ( .A(n1353), .B(n3119), .S(n3231), .Z(n874) );
  MUX21L U1651 ( .A(n1354), .B(n3121), .S(n3031), .Z(n875) );
  MUX21L U1652 ( .A(n1355), .B(n3122), .S(n3231), .Z(n876) );
  MUX21L U1653 ( .A(n1356), .B(n3123), .S(n3031), .Z(n877) );
  MUX21L U1654 ( .A(n1357), .B(n3124), .S(n3231), .Z(n878) );
  MUX21L U1655 ( .A(n1358), .B(n3125), .S(n3031), .Z(n879) );
  MUX21L U1656 ( .A(n1359), .B(n3126), .S(n3231), .Z(n880) );
  MUX21L U1657 ( .A(n1360), .B(n3128), .S(n3231), .Z(n881) );
  MUX21L U1658 ( .A(n1361), .B(n3129), .S(n3231), .Z(n882) );
  MUX21L U1659 ( .A(n1362), .B(n3133), .S(n3231), .Z(n883) );
  ND2I U1660 ( .A(n2106), .B(n2109), .Z(n3232) );
  IVI U1661 ( .A(n3232), .Z(n3234) );
  MUX21L U1662 ( .A(n1363), .B(n3090), .S(n3033), .Z(n820) );
  MUX21L U1663 ( .A(n1364), .B(n3092), .S(n3033), .Z(n821) );
  MUX21L U1664 ( .A(n1365), .B(n3094), .S(n3033), .Z(n822) );
  MUX21L U1665 ( .A(n1366), .B(n3096), .S(n3033), .Z(n823) );
  MUX21L U1666 ( .A(n1367), .B(n3098), .S(n3032), .Z(n824) );
  MUX21L U1667 ( .A(n1368), .B(n3099), .S(n3032), .Z(n825) );
  MUX21L U1668 ( .A(n3233), .B(n3100), .S(n3032), .Z(n826) );
  MUX21L U1669 ( .A(n1369), .B(n3101), .S(n3032), .Z(n827) );
  MUX21L U1670 ( .A(n1370), .B(n3102), .S(n3032), .Z(n828) );
  MUX21L U1671 ( .A(n1371), .B(n3103), .S(n3032), .Z(n829) );
  MUX21L U1672 ( .A(n1372), .B(n3104), .S(n3032), .Z(n830) );
  MUX21L U1673 ( .A(n1373), .B(n3105), .S(n3032), .Z(n831) );
  MUX21L U1674 ( .A(n1374), .B(n3106), .S(n3032), .Z(n832) );
  MUX21L U1675 ( .A(n1375), .B(n3107), .S(n3032), .Z(n833) );
  MUX21L U1676 ( .A(n1376), .B(n3109), .S(n3032), .Z(n834) );
  MUX21L U1677 ( .A(n1377), .B(n3110), .S(n3032), .Z(n835) );
  MUX21L U1678 ( .A(n1378), .B(n3112), .S(n3032), .Z(n836) );
  MUX21L U1679 ( .A(n1379), .B(n3113), .S(n3032), .Z(n837) );
  MUX21L U1680 ( .A(n1380), .B(n3114), .S(n3234), .Z(n838) );
  MUX21L U1681 ( .A(n1381), .B(n3115), .S(n3032), .Z(n839) );
  MUX21L U1682 ( .A(n1382), .B(n3116), .S(n3032), .Z(n840) );
  MUX21L U1683 ( .A(n1383), .B(n3117), .S(n3033), .Z(n841) );
  MUX21L U1684 ( .A(n1384), .B(n3119), .S(n3234), .Z(n842) );
  MUX21L U1685 ( .A(n1385), .B(n3121), .S(n3033), .Z(n843) );
  MUX21L U1686 ( .A(n1386), .B(n3122), .S(n3234), .Z(n844) );
  MUX21L U1687 ( .A(n1387), .B(n3123), .S(n3033), .Z(n845) );
  MUX21L U1688 ( .A(n1388), .B(n3124), .S(n3234), .Z(n846) );
  MUX21L U1689 ( .A(n1389), .B(n3125), .S(n3033), .Z(n847) );
  MUX21L U1690 ( .A(n1390), .B(n3126), .S(n3234), .Z(n848) );
  MUX21L U1691 ( .A(n1391), .B(n3128), .S(n3234), .Z(n849) );
  MUX21L U1692 ( .A(n1392), .B(n3129), .S(n3234), .Z(n850) );
  MUX21L U1693 ( .A(n1393), .B(n3133), .S(n3234), .Z(n851) );
  ND2I U1694 ( .A(n2106), .B(n2111), .Z(n3235) );
  IVI U1695 ( .A(n3235), .Z(n3237) );
  MUX21L U1696 ( .A(n1394), .B(n3090), .S(n3035), .Z(n788) );
  MUX21L U1697 ( .A(n1395), .B(n3092), .S(n3035), .Z(n789) );
  MUX21L U1698 ( .A(n1396), .B(n3094), .S(n3035), .Z(n790) );
  MUX21L U1699 ( .A(n1397), .B(n3096), .S(n3035), .Z(n791) );
  MUX21L U1700 ( .A(n1398), .B(n3098), .S(n3034), .Z(n792) );
  MUX21L U1701 ( .A(n1399), .B(n3099), .S(n3034), .Z(n793) );
  MUX21L U1702 ( .A(n3236), .B(n3100), .S(n3034), .Z(n794) );
  MUX21L U1703 ( .A(n1400), .B(n3101), .S(n3034), .Z(n795) );
  MUX21L U1704 ( .A(n1401), .B(n3102), .S(n3034), .Z(n796) );
  MUX21L U1705 ( .A(n1402), .B(n3103), .S(n3034), .Z(n797) );
  MUX21L U1706 ( .A(n1403), .B(n3104), .S(n3034), .Z(n798) );
  MUX21L U1707 ( .A(n1404), .B(n3105), .S(n3034), .Z(n799) );
  MUX21L U1708 ( .A(n1405), .B(n3106), .S(n3034), .Z(n800) );
  MUX21L U1709 ( .A(n1406), .B(n3107), .S(n3034), .Z(n801) );
  MUX21L U1710 ( .A(n1407), .B(n3109), .S(n3034), .Z(n802) );
  MUX21L U1711 ( .A(n1408), .B(n3110), .S(n3034), .Z(n803) );
  MUX21L U1712 ( .A(n1409), .B(n3112), .S(n3034), .Z(n804) );
  MUX21L U1713 ( .A(n1410), .B(n3113), .S(n3034), .Z(n805) );
  MUX21L U1714 ( .A(n1411), .B(n3114), .S(n3237), .Z(n806) );
  MUX21L U1715 ( .A(n1412), .B(n3115), .S(n3034), .Z(n807) );
  MUX21L U1716 ( .A(n1413), .B(n3116), .S(n3034), .Z(n808) );
  MUX21L U1717 ( .A(n1414), .B(n3117), .S(n3035), .Z(n809) );
  MUX21L U1718 ( .A(n1415), .B(n3119), .S(n3237), .Z(n810) );
  MUX21L U1719 ( .A(n1416), .B(n3121), .S(n3035), .Z(n811) );
  MUX21L U1720 ( .A(n1417), .B(n3122), .S(n3237), .Z(n812) );
  MUX21L U1721 ( .A(n1418), .B(n3123), .S(n3035), .Z(n813) );
  MUX21L U1722 ( .A(n1419), .B(n3124), .S(n3237), .Z(n814) );
  MUX21L U1723 ( .A(n1420), .B(n3125), .S(n3035), .Z(n815) );
  MUX21L U1724 ( .A(n1421), .B(n3126), .S(n3237), .Z(n816) );
  MUX21L U1725 ( .A(n1422), .B(n3128), .S(n3237), .Z(n817) );
  MUX21L U1726 ( .A(n1423), .B(n3129), .S(n3237), .Z(n818) );
  MUX21L U1727 ( .A(n1424), .B(n3133), .S(n3237), .Z(n819) );
  ND2I U1728 ( .A(n2106), .B(n2108), .Z(n3238) );
  IVI U1729 ( .A(n3238), .Z(n3240) );
  MUX21L U1730 ( .A(n1425), .B(n3090), .S(n3037), .Z(n756) );
  MUX21L U1731 ( .A(n1426), .B(n3092), .S(n3037), .Z(n757) );
  MUX21L U1732 ( .A(n1427), .B(n3094), .S(n3037), .Z(n758) );
  MUX21L U1733 ( .A(n1428), .B(n3096), .S(n3037), .Z(n759) );
  MUX21L U1734 ( .A(n1429), .B(n3098), .S(n3036), .Z(n760) );
  MUX21L U1735 ( .A(n1430), .B(n3099), .S(n3036), .Z(n761) );
  MUX21L U1736 ( .A(n3239), .B(n3100), .S(n3036), .Z(n762) );
  MUX21L U1737 ( .A(n1431), .B(n3101), .S(n3036), .Z(n763) );
  MUX21L U1738 ( .A(n1432), .B(n3102), .S(n3036), .Z(n764) );
  MUX21L U1739 ( .A(n1433), .B(n3103), .S(n3036), .Z(n765) );
  MUX21L U1740 ( .A(n1434), .B(n3104), .S(n3036), .Z(n766) );
  MUX21L U1741 ( .A(n1435), .B(n3105), .S(n3036), .Z(n767) );
  MUX21L U1742 ( .A(n1436), .B(n3106), .S(n3036), .Z(n768) );
  MUX21L U1743 ( .A(n1437), .B(n3107), .S(n3036), .Z(n769) );
  MUX21L U1744 ( .A(n1438), .B(n3109), .S(n3036), .Z(n770) );
  MUX21L U1745 ( .A(n1439), .B(n3110), .S(n3036), .Z(n771) );
  MUX21L U1746 ( .A(n1440), .B(n3112), .S(n3036), .Z(n772) );
  MUX21L U1747 ( .A(n1441), .B(n3113), .S(n3036), .Z(n773) );
  MUX21L U1748 ( .A(n1442), .B(n3114), .S(n3240), .Z(n774) );
  MUX21L U1749 ( .A(n1443), .B(n3115), .S(n3036), .Z(n775) );
  MUX21L U1750 ( .A(n1444), .B(n3116), .S(n3036), .Z(n776) );
  MUX21L U1751 ( .A(n1445), .B(n3117), .S(n3037), .Z(n777) );
  MUX21L U1752 ( .A(n1446), .B(n3119), .S(n3240), .Z(n778) );
  MUX21L U1753 ( .A(n1447), .B(n3121), .S(n3037), .Z(n779) );
  MUX21L U1754 ( .A(n1448), .B(n3122), .S(n3240), .Z(n780) );
  MUX21L U1755 ( .A(n1449), .B(n3123), .S(n3037), .Z(n781) );
  MUX21L U1756 ( .A(n1450), .B(n3124), .S(n3240), .Z(n782) );
  MUX21L U1757 ( .A(n1451), .B(n3125), .S(n3037), .Z(n783) );
  MUX21L U1758 ( .A(n1452), .B(n3126), .S(n3240), .Z(n784) );
  MUX21L U1759 ( .A(n1453), .B(n3128), .S(n3240), .Z(n785) );
  MUX21L U1760 ( .A(n1454), .B(n3129), .S(n3240), .Z(n786) );
  MUX21L U1761 ( .A(n1455), .B(n3133), .S(n3240), .Z(n787) );
  ND2I U1762 ( .A(n2106), .B(n2110), .Z(n3241) );
  IVI U1763 ( .A(n3241), .Z(n3243) );
  MUX21L U1764 ( .A(n1456), .B(n3090), .S(n3039), .Z(n724) );
  MUX21L U1765 ( .A(n1457), .B(n3092), .S(n3039), .Z(n725) );
  MUX21L U1766 ( .A(n1458), .B(n3094), .S(n3039), .Z(n726) );
  MUX21L U1767 ( .A(n1459), .B(n3096), .S(n3039), .Z(n727) );
  MUX21L U1768 ( .A(n1460), .B(n3098), .S(n3038), .Z(n728) );
  MUX21L U1769 ( .A(n1461), .B(n3099), .S(n3038), .Z(n729) );
  MUX21L U1770 ( .A(n3242), .B(n3100), .S(n3038), .Z(n730) );
  MUX21L U1771 ( .A(n1462), .B(n3101), .S(n3038), .Z(n731) );
  MUX21L U1772 ( .A(n1463), .B(n3102), .S(n3038), .Z(n732) );
  MUX21L U1773 ( .A(n1464), .B(n3103), .S(n3038), .Z(n733) );
  MUX21L U1774 ( .A(n1465), .B(n3104), .S(n3038), .Z(n734) );
  MUX21L U1775 ( .A(n1466), .B(n3105), .S(n3038), .Z(n735) );
  MUX21L U1776 ( .A(n1467), .B(n3106), .S(n3038), .Z(n736) );
  MUX21L U1777 ( .A(n1468), .B(n3107), .S(n3038), .Z(n737) );
  MUX21L U1778 ( .A(n1469), .B(n3109), .S(n3038), .Z(n738) );
  MUX21L U1779 ( .A(n1470), .B(n3110), .S(n3038), .Z(n739) );
  MUX21L U1780 ( .A(n1471), .B(n3112), .S(n3038), .Z(n740) );
  MUX21L U1781 ( .A(n1472), .B(n3113), .S(n3038), .Z(n741) );
  MUX21L U1782 ( .A(n1473), .B(n3114), .S(n3243), .Z(n742) );
  MUX21L U1783 ( .A(n1474), .B(n3115), .S(n3038), .Z(n743) );
  MUX21L U1784 ( .A(n1475), .B(n3116), .S(n3038), .Z(n744) );
  MUX21L U1785 ( .A(n1476), .B(n3117), .S(n3039), .Z(n745) );
  MUX21L U1786 ( .A(n1477), .B(n3119), .S(n3243), .Z(n746) );
  MUX21L U1787 ( .A(n1478), .B(n3121), .S(n3039), .Z(n747) );
  MUX21L U1788 ( .A(n1479), .B(n3122), .S(n3243), .Z(n748) );
  MUX21L U1789 ( .A(n1480), .B(n3123), .S(n3039), .Z(n749) );
  MUX21L U1790 ( .A(n1481), .B(n3124), .S(n3243), .Z(n750) );
  MUX21L U1791 ( .A(n1482), .B(n3125), .S(n3039), .Z(n751) );
  MUX21L U1792 ( .A(n1483), .B(n3126), .S(n3243), .Z(n752) );
  MUX21L U1793 ( .A(n1484), .B(n3128), .S(n3243), .Z(n753) );
  MUX21L U1794 ( .A(n1485), .B(n3129), .S(n3243), .Z(n754) );
  MUX21L U1795 ( .A(n1486), .B(n3133), .S(n3243), .Z(n755) );
  ND2I U1796 ( .A(n2106), .B(n2104), .Z(n3244) );
  IVI U1797 ( .A(n3244), .Z(n3246) );
  MUX21L U1798 ( .A(n132), .B(n3090), .S(n3041), .Z(n692) );
  MUX21L U1799 ( .A(n135), .B(n3092), .S(n3041), .Z(n693) );
  MUX21L U1800 ( .A(n138), .B(n3094), .S(n3041), .Z(n694) );
  MUX21L U1801 ( .A(n1487), .B(n3096), .S(n3041), .Z(n695) );
  MUX21L U1802 ( .A(n1488), .B(n3098), .S(n3040), .Z(n696) );
  MUX21L U1803 ( .A(n1489), .B(n3099), .S(n3040), .Z(n697) );
  MUX21L U1804 ( .A(n3245), .B(n3100), .S(n3040), .Z(n698) );
  MUX21L U1805 ( .A(n1490), .B(n3101), .S(n3040), .Z(n699) );
  MUX21L U1806 ( .A(n1491), .B(n3102), .S(n3040), .Z(n700) );
  MUX21L U1807 ( .A(n1492), .B(n3103), .S(n3040), .Z(n701) );
  MUX21L U1808 ( .A(n1493), .B(n3104), .S(n3040), .Z(n702) );
  MUX21L U1809 ( .A(n1494), .B(n3105), .S(n3040), .Z(n703) );
  MUX21L U1810 ( .A(n1495), .B(n3106), .S(n3040), .Z(n704) );
  MUX21L U1811 ( .A(n1496), .B(n3107), .S(n3040), .Z(n705) );
  MUX21L U1812 ( .A(n1497), .B(n3109), .S(n3040), .Z(n706) );
  MUX21L U1813 ( .A(n1498), .B(n3110), .S(n3040), .Z(n707) );
  MUX21L U1814 ( .A(n1499), .B(n3112), .S(n3040), .Z(n708) );
  MUX21L U1815 ( .A(n1500), .B(n3113), .S(n3040), .Z(n709) );
  MUX21L U1816 ( .A(n1501), .B(n3114), .S(n3246), .Z(n710) );
  MUX21L U1817 ( .A(n1502), .B(n3115), .S(n3040), .Z(n711) );
  MUX21L U1818 ( .A(n1503), .B(n3116), .S(n3040), .Z(n712) );
  MUX21L U1819 ( .A(n1504), .B(n3117), .S(n3041), .Z(n713) );
  MUX21L U1820 ( .A(n1505), .B(n3119), .S(n3246), .Z(n714) );
  MUX21L U1821 ( .A(n1506), .B(n3121), .S(n3041), .Z(n715) );
  MUX21L U1822 ( .A(n1507), .B(n3122), .S(n3246), .Z(n716) );
  MUX21L U1823 ( .A(n1508), .B(n3123), .S(n3041), .Z(n717) );
  MUX21L U1824 ( .A(n1509), .B(n3124), .S(n3246), .Z(n718) );
  MUX21L U1825 ( .A(n1510), .B(n3125), .S(n3041), .Z(n719) );
  MUX21L U1826 ( .A(n1511), .B(n3126), .S(n3246), .Z(n720) );
  MUX21L U1827 ( .A(n1512), .B(n3128), .S(n3246), .Z(n721) );
  MUX21L U1828 ( .A(n1513), .B(n3129), .S(n3246), .Z(n722) );
  MUX21L U1829 ( .A(n1514), .B(n3133), .S(n3246), .Z(n723) );
  MUX21L U1830 ( .A(n63), .B(n3090), .S(n3043), .Z(n660) );
  MUX21L U1831 ( .A(n66), .B(n3092), .S(n3043), .Z(n661) );
  MUX21L U1832 ( .A(n69), .B(n3094), .S(n3043), .Z(n662) );
  MUX21L U1833 ( .A(n1515), .B(n3096), .S(n3043), .Z(n663) );
  MUX21L U1834 ( .A(n1516), .B(n3098), .S(n3042), .Z(n664) );
  MUX21L U1835 ( .A(n1517), .B(n3099), .S(n3042), .Z(n665) );
  MUX21L U1836 ( .A(n3247), .B(n3100), .S(n3042), .Z(n666) );
  MUX21L U1837 ( .A(n1518), .B(n3101), .S(n3042), .Z(n667) );
  MUX21L U1838 ( .A(n1519), .B(n3102), .S(n3042), .Z(n668) );
  MUX21L U1839 ( .A(n1520), .B(n3103), .S(n3042), .Z(n669) );
  MUX21L U1840 ( .A(n1521), .B(n3104), .S(n3042), .Z(n670) );
  MUX21L U1841 ( .A(n1522), .B(n3105), .S(n3042), .Z(n671) );
  MUX21L U1842 ( .A(n1523), .B(n3106), .S(n3042), .Z(n672) );
  MUX21L U1843 ( .A(n1524), .B(n3107), .S(n3042), .Z(n673) );
  MUX21L U1844 ( .A(n1525), .B(n3109), .S(n3042), .Z(n674) );
  MUX21L U1845 ( .A(n1526), .B(n3110), .S(n3042), .Z(n675) );
  MUX21L U1846 ( .A(n1527), .B(n3112), .S(n3042), .Z(n676) );
  MUX21L U1847 ( .A(n1528), .B(n3113), .S(n3042), .Z(n677) );
  MUX21L U1848 ( .A(n1529), .B(n3114), .S(n76), .Z(n678) );
  MUX21L U1849 ( .A(n1530), .B(n3115), .S(n76), .Z(n679) );
  MUX21L U1850 ( .A(n1531), .B(n3116), .S(n76), .Z(n680) );
  MUX21L U1851 ( .A(n1532), .B(n3117), .S(n76), .Z(n681) );
  MUX21L U1852 ( .A(n1533), .B(n3119), .S(n76), .Z(n682) );
  MUX21L U1853 ( .A(n1534), .B(n3121), .S(n76), .Z(n683) );
  MUX21L U1854 ( .A(n1535), .B(n3122), .S(n76), .Z(n684) );
  MUX21L U1855 ( .A(n1536), .B(n3123), .S(n76), .Z(n685) );
  MUX21L U1856 ( .A(n1537), .B(n3124), .S(n76), .Z(n686) );
  MUX21L U1857 ( .A(n1538), .B(n3125), .S(n76), .Z(n687) );
  MUX21L U1858 ( .A(n1539), .B(n3126), .S(n76), .Z(n688) );
  MUX21L U1859 ( .A(n1540), .B(n3128), .S(n76), .Z(n689) );
  MUX21L U1860 ( .A(n1541), .B(n3129), .S(n76), .Z(n690) );
  MUX21L U1861 ( .A(n1542), .B(n3133), .S(n76), .Z(n691) );
  MUX21L U1862 ( .A(n1543), .B(n3090), .S(n3046), .Z(n628) );
  MUX21L U1863 ( .A(n1544), .B(n3092), .S(n3046), .Z(n629) );
  MUX21L U1864 ( .A(n1545), .B(n3094), .S(n3046), .Z(n630) );
  MUX21L U1865 ( .A(n1546), .B(n3096), .S(n3046), .Z(n631) );
  MUX21L U1866 ( .A(n1547), .B(n3098), .S(n3045), .Z(n632) );
  MUX21L U1867 ( .A(n1548), .B(n3099), .S(n3045), .Z(n633) );
  MUX21L U1868 ( .A(n1549), .B(n3100), .S(n3045), .Z(n634) );
  MUX21L U1869 ( .A(n1550), .B(n3101), .S(n3045), .Z(n635) );
  MUX21L U1870 ( .A(n1551), .B(n3102), .S(n3045), .Z(n636) );
  MUX21L U1871 ( .A(n1552), .B(n3103), .S(n3045), .Z(n637) );
  MUX21L U1872 ( .A(n1553), .B(n3104), .S(n3045), .Z(n638) );
  MUX21L U1873 ( .A(n1554), .B(n3105), .S(n3045), .Z(n639) );
  MUX21L U1874 ( .A(n1555), .B(n3106), .S(n3045), .Z(n640) );
  MUX21L U1875 ( .A(n1556), .B(n3107), .S(n3045), .Z(n641) );
  MUX21L U1876 ( .A(n1557), .B(n3109), .S(n3045), .Z(n642) );
  MUX21L U1877 ( .A(n1558), .B(n3110), .S(n3045), .Z(n643) );
  MUX21L U1878 ( .A(n1559), .B(n3112), .S(n3045), .Z(n644) );
  MUX21L U1879 ( .A(n1560), .B(n3113), .S(n3045), .Z(n645) );
  MUX21L U1880 ( .A(n1561), .B(n3114), .S(n3044), .Z(n646) );
  MUX21L U1881 ( .A(n1562), .B(n3115), .S(n3044), .Z(n647) );
  MUX21L U1882 ( .A(n1563), .B(n3116), .S(n3044), .Z(n648) );
  MUX21L U1883 ( .A(n1564), .B(n3117), .S(n3044), .Z(n649) );
  MUX21L U1884 ( .A(n1565), .B(n3119), .S(n3044), .Z(n650) );
  MUX21L U1885 ( .A(n1566), .B(n3121), .S(n3044), .Z(n651) );
  MUX21L U1886 ( .A(n1567), .B(n3122), .S(n3044), .Z(n652) );
  MUX21L U1887 ( .A(n1568), .B(n3123), .S(n3044), .Z(n653) );
  MUX21L U1888 ( .A(n1569), .B(n3124), .S(n3044), .Z(n654) );
  MUX21L U1889 ( .A(n1570), .B(n3125), .S(n3044), .Z(n655) );
  MUX21L U1890 ( .A(n1571), .B(n3126), .S(n3044), .Z(n656) );
  MUX21L U1891 ( .A(n1572), .B(n3128), .S(n3044), .Z(n657) );
  MUX21L U1892 ( .A(n1573), .B(n3129), .S(n3044), .Z(n658) );
  MUX21L U1893 ( .A(n1574), .B(n3133), .S(n3044), .Z(n659) );
  ND2I U1894 ( .A(n2103), .B(n2112), .Z(n3249) );
  MUX21L U1895 ( .A(n1575), .B(n3090), .S(n3049), .Z(n596) );
  MUX21L U1896 ( .A(n1576), .B(n3092), .S(n3049), .Z(n597) );
  MUX21L U1897 ( .A(n1577), .B(n3094), .S(n3049), .Z(n598) );
  MUX21L U1898 ( .A(n1578), .B(n3096), .S(n3049), .Z(n599) );
  MUX21L U1899 ( .A(n1579), .B(n3098), .S(n3048), .Z(n600) );
  MUX21L U1900 ( .A(n1580), .B(n3099), .S(n3048), .Z(n601) );
  MUX21L U1901 ( .A(n1581), .B(n3100), .S(n3048), .Z(n602) );
  MUX21L U1902 ( .A(n1582), .B(n3101), .S(n3048), .Z(n603) );
  MUX21L U1903 ( .A(n1583), .B(n3102), .S(n3048), .Z(n604) );
  MUX21L U1904 ( .A(n3250), .B(n3103), .S(n3048), .Z(n605) );
  MUX21L U1905 ( .A(n1584), .B(n3104), .S(n3048), .Z(n606) );
  MUX21L U1906 ( .A(n1585), .B(n3105), .S(n3048), .Z(n607) );
  MUX21L U1907 ( .A(n1586), .B(n3106), .S(n3048), .Z(n608) );
  MUX21L U1908 ( .A(n1587), .B(n3107), .S(n3048), .Z(n609) );
  MUX21L U1909 ( .A(n1588), .B(n3109), .S(n3048), .Z(n610) );
  MUX21L U1910 ( .A(n1589), .B(n3110), .S(n3048), .Z(n611) );
  MUX21L U1911 ( .A(n1590), .B(n3112), .S(n3048), .Z(n612) );
  MUX21L U1912 ( .A(n1591), .B(n3113), .S(n3048), .Z(n613) );
  MUX21L U1913 ( .A(n1592), .B(n3114), .S(n3047), .Z(n614) );
  MUX21L U1914 ( .A(n1593), .B(n3115), .S(n3047), .Z(n615) );
  MUX21L U1915 ( .A(n1594), .B(n3116), .S(n3047), .Z(n616) );
  MUX21L U1916 ( .A(n1595), .B(n3117), .S(n3047), .Z(n617) );
  MUX21L U1917 ( .A(n1596), .B(n3119), .S(n3047), .Z(n618) );
  MUX21L U1918 ( .A(n1597), .B(n3121), .S(n3047), .Z(n619) );
  MUX21L U1919 ( .A(n1598), .B(n3122), .S(n3047), .Z(n620) );
  MUX21L U1920 ( .A(n1599), .B(n3123), .S(n3047), .Z(n621) );
  MUX21L U1921 ( .A(n1600), .B(n3124), .S(n3047), .Z(n622) );
  MUX21L U1922 ( .A(n1601), .B(n3125), .S(n3047), .Z(n623) );
  MUX21L U1923 ( .A(n1602), .B(n3126), .S(n3047), .Z(n624) );
  MUX21L U1924 ( .A(n1603), .B(n3128), .S(n3047), .Z(n625) );
  MUX21L U1925 ( .A(n1604), .B(n3129), .S(n3047), .Z(n626) );
  MUX21L U1926 ( .A(n1605), .B(n3133), .S(n3047), .Z(n627) );
  ND2I U1927 ( .A(n2103), .B(n2109), .Z(n3251) );
  MUX21L U1928 ( .A(n133), .B(n3089), .S(n3052), .Z(n564) );
  MUX21L U1929 ( .A(n136), .B(n3091), .S(n3052), .Z(n565) );
  MUX21L U1930 ( .A(n139), .B(n3093), .S(n3052), .Z(n566) );
  MUX21L U1931 ( .A(n1606), .B(n3095), .S(n3052), .Z(n567) );
  MUX21L U1932 ( .A(n1607), .B(n3097), .S(n3051), .Z(n568) );
  MUX21L U1933 ( .A(n1608), .B(n3099), .S(n3051), .Z(n569) );
  MUX21L U1934 ( .A(n1609), .B(n3100), .S(n3051), .Z(n570) );
  MUX21L U1935 ( .A(n1610), .B(n3101), .S(n3051), .Z(n571) );
  MUX21L U1936 ( .A(n1611), .B(n3102), .S(n3051), .Z(n572) );
  MUX21L U1937 ( .A(n1612), .B(n3103), .S(n3051), .Z(n573) );
  MUX21L U1938 ( .A(n1613), .B(n3104), .S(n3051), .Z(n574) );
  MUX21L U1939 ( .A(n1614), .B(n3105), .S(n3051), .Z(n575) );
  MUX21L U1940 ( .A(n1615), .B(n3106), .S(n3051), .Z(n576) );
  MUX21L U1941 ( .A(n1616), .B(n3107), .S(n3051), .Z(n577) );
  MUX21L U1942 ( .A(n1617), .B(n3108), .S(n3051), .Z(n578) );
  MUX21L U1943 ( .A(n1618), .B(n3110), .S(n3051), .Z(n579) );
  MUX21L U1944 ( .A(n1619), .B(n3111), .S(n3051), .Z(n580) );
  MUX21L U1945 ( .A(n1620), .B(n3113), .S(n3051), .Z(n581) );
  MUX21L U1946 ( .A(n1621), .B(n3114), .S(n3050), .Z(n582) );
  MUX21L U1947 ( .A(n1622), .B(n3115), .S(n3050), .Z(n583) );
  MUX21L U1948 ( .A(n1623), .B(n3116), .S(n3050), .Z(n584) );
  MUX21L U1949 ( .A(n1624), .B(n3117), .S(n3050), .Z(n585) );
  MUX21L U1950 ( .A(n1625), .B(n3118), .S(n3050), .Z(n586) );
  MUX21L U1951 ( .A(n1626), .B(n3121), .S(n3050), .Z(n587) );
  MUX21L U1952 ( .A(n1627), .B(n3122), .S(n3050), .Z(n588) );
  MUX21L U1953 ( .A(n1628), .B(n3123), .S(n3050), .Z(n589) );
  MUX21L U1954 ( .A(n1629), .B(n3124), .S(n3050), .Z(n590) );
  MUX21L U1955 ( .A(n1630), .B(n3125), .S(n3050), .Z(n591) );
  MUX21L U1956 ( .A(n1631), .B(n3126), .S(n3050), .Z(n592) );
  MUX21L U1957 ( .A(n1632), .B(n3127), .S(n3050), .Z(n593) );
  MUX21L U1958 ( .A(n1633), .B(n3129), .S(n3050), .Z(n594) );
  MUX21L U1959 ( .A(n1634), .B(n3133), .S(n3050), .Z(n595) );
  ND2I U1960 ( .A(n2103), .B(n2111), .Z(n3252) );
  MUX21L U1961 ( .A(n64), .B(n3089), .S(n3055), .Z(n532) );
  MUX21L U1962 ( .A(n67), .B(n3091), .S(n3055), .Z(n533) );
  MUX21L U1963 ( .A(n70), .B(n3093), .S(n3055), .Z(n534) );
  MUX21L U1964 ( .A(n1635), .B(n3095), .S(n3055), .Z(n535) );
  MUX21L U1965 ( .A(n1636), .B(n3097), .S(n3054), .Z(n536) );
  MUX21L U1966 ( .A(n1637), .B(n3099), .S(n3054), .Z(n537) );
  MUX21L U1967 ( .A(n1638), .B(n3100), .S(n3054), .Z(n538) );
  MUX21L U1968 ( .A(n1639), .B(n3101), .S(n3054), .Z(n539) );
  MUX21L U1969 ( .A(n1640), .B(n3102), .S(n3054), .Z(n540) );
  MUX21L U1970 ( .A(n1641), .B(n3103), .S(n3054), .Z(n541) );
  MUX21L U1971 ( .A(n1642), .B(n3104), .S(n3054), .Z(n542) );
  MUX21L U1972 ( .A(n1643), .B(n3105), .S(n3054), .Z(n543) );
  MUX21L U1973 ( .A(n1644), .B(n3106), .S(n3054), .Z(n544) );
  MUX21L U1974 ( .A(n1645), .B(n3107), .S(n3054), .Z(n545) );
  MUX21L U1975 ( .A(n1646), .B(n3108), .S(n3054), .Z(n546) );
  MUX21L U1976 ( .A(n1647), .B(n3110), .S(n3054), .Z(n547) );
  MUX21L U1977 ( .A(n1648), .B(n3111), .S(n3054), .Z(n548) );
  MUX21L U1978 ( .A(n1649), .B(n3113), .S(n3054), .Z(n549) );
  MUX21L U1979 ( .A(n1650), .B(n3114), .S(n3053), .Z(n550) );
  MUX21L U1980 ( .A(n1651), .B(n3115), .S(n3053), .Z(n551) );
  MUX21L U1981 ( .A(n1652), .B(n3116), .S(n3053), .Z(n552) );
  MUX21L U1982 ( .A(n1653), .B(n3117), .S(n3053), .Z(n553) );
  MUX21L U1983 ( .A(n1654), .B(n3118), .S(n3053), .Z(n554) );
  MUX21L U1984 ( .A(n1655), .B(n3121), .S(n3053), .Z(n555) );
  MUX21L U1985 ( .A(n1656), .B(n3122), .S(n3053), .Z(n556) );
  MUX21L U1986 ( .A(n1657), .B(n3123), .S(n3053), .Z(n557) );
  MUX21L U1987 ( .A(n1658), .B(n3124), .S(n3053), .Z(n558) );
  MUX21L U1988 ( .A(n1659), .B(n3125), .S(n3053), .Z(n559) );
  MUX21L U1989 ( .A(n1660), .B(n3126), .S(n3053), .Z(n560) );
  MUX21L U1990 ( .A(n1661), .B(n3127), .S(n3053), .Z(n561) );
  MUX21L U1991 ( .A(n1662), .B(n3129), .S(n3053), .Z(n562) );
  MUX21L U1992 ( .A(n1663), .B(n3133), .S(n3053), .Z(n563) );
  ND2I U1993 ( .A(n2103), .B(n2108), .Z(n3253) );
  MUX21L U1994 ( .A(n59), .B(n3089), .S(n3058), .Z(n500) );
  MUX21L U1995 ( .A(n54), .B(n3091), .S(n3058), .Z(n501) );
  MUX21L U1996 ( .A(n55), .B(n3093), .S(n3058), .Z(n502) );
  MUX21L U1997 ( .A(n1664), .B(n3095), .S(n3058), .Z(n503) );
  MUX21L U1998 ( .A(n3254), .B(n3097), .S(n3057), .Z(n504) );
  MUX21L U1999 ( .A(n1665), .B(n3099), .S(n3057), .Z(n505) );
  MUX21L U2000 ( .A(n1666), .B(n3100), .S(n3057), .Z(n506) );
  MUX21L U2001 ( .A(n1667), .B(n3101), .S(n3057), .Z(n507) );
  MUX21L U2002 ( .A(n1668), .B(n3102), .S(n3057), .Z(n508) );
  MUX21L U2003 ( .A(n1669), .B(n3103), .S(n3057), .Z(n509) );
  MUX21L U2004 ( .A(n1670), .B(n3104), .S(n3057), .Z(n510) );
  MUX21L U2005 ( .A(n1671), .B(n3105), .S(n3057), .Z(n511) );
  MUX21L U2006 ( .A(n1672), .B(n3106), .S(n3057), .Z(n512) );
  MUX21L U2007 ( .A(n1673), .B(n3107), .S(n3057), .Z(n513) );
  MUX21L U2008 ( .A(n1674), .B(n3108), .S(n3057), .Z(n514) );
  MUX21L U2009 ( .A(n1675), .B(n3110), .S(n3057), .Z(n515) );
  MUX21L U2010 ( .A(n1676), .B(n3111), .S(n3057), .Z(n516) );
  MUX21L U2011 ( .A(n1677), .B(n3113), .S(n3057), .Z(n517) );
  MUX21L U2012 ( .A(n1678), .B(n3114), .S(n3056), .Z(n518) );
  MUX21L U2013 ( .A(n1679), .B(n3115), .S(n3056), .Z(n519) );
  MUX21L U2014 ( .A(n1680), .B(n3116), .S(n3056), .Z(n520) );
  MUX21L U2015 ( .A(n1681), .B(n3117), .S(n3056), .Z(n521) );
  MUX21L U2016 ( .A(n1682), .B(n3118), .S(n3056), .Z(n522) );
  MUX21L U2017 ( .A(n1683), .B(n3121), .S(n3056), .Z(n523) );
  MUX21L U2018 ( .A(n1684), .B(n3122), .S(n3056), .Z(n524) );
  MUX21L U2019 ( .A(n1685), .B(n3123), .S(n3056), .Z(n525) );
  MUX21L U2020 ( .A(n1686), .B(n3124), .S(n3056), .Z(n526) );
  MUX21L U2021 ( .A(n1687), .B(n3125), .S(n3056), .Z(n527) );
  MUX21L U2022 ( .A(n1688), .B(n3126), .S(n3056), .Z(n528) );
  MUX21L U2023 ( .A(n1689), .B(n3127), .S(n3056), .Z(n529) );
  MUX21L U2024 ( .A(n1690), .B(n3129), .S(n3056), .Z(n530) );
  MUX21L U2025 ( .A(n1691), .B(n3133), .S(n3056), .Z(n531) );
  ND2I U2026 ( .A(n2103), .B(n2110), .Z(n3255) );
  MUX21L U2027 ( .A(n128), .B(n3089), .S(n3061), .Z(n468) );
  MUX21L U2028 ( .A(n123), .B(n3091), .S(n3061), .Z(n469) );
  MUX21L U2029 ( .A(n124), .B(n3093), .S(n3061), .Z(n470) );
  MUX21L U2030 ( .A(n1692), .B(n3095), .S(n3061), .Z(n471) );
  MUX21L U2031 ( .A(n1693), .B(n3097), .S(n3060), .Z(n472) );
  MUX21L U2032 ( .A(n1694), .B(n3099), .S(n3060), .Z(n473) );
  MUX21L U2033 ( .A(n1695), .B(n3100), .S(n3060), .Z(n474) );
  MUX21L U2034 ( .A(n1696), .B(n3101), .S(n3060), .Z(n475) );
  MUX21L U2035 ( .A(n1697), .B(n3102), .S(n3060), .Z(n476) );
  MUX21L U2036 ( .A(n1698), .B(n3103), .S(n3060), .Z(n477) );
  MUX21L U2037 ( .A(n1699), .B(n3104), .S(n3060), .Z(n478) );
  MUX21L U2038 ( .A(n1700), .B(n3105), .S(n3060), .Z(n479) );
  MUX21L U2039 ( .A(n1701), .B(n3106), .S(n3060), .Z(n480) );
  MUX21L U2040 ( .A(n1702), .B(n3107), .S(n3060), .Z(n481) );
  MUX21L U2041 ( .A(n1703), .B(n3108), .S(n3060), .Z(n482) );
  MUX21L U2042 ( .A(n1704), .B(n3110), .S(n3060), .Z(n483) );
  MUX21L U2043 ( .A(n1705), .B(n3111), .S(n3060), .Z(n484) );
  MUX21L U2044 ( .A(n1706), .B(n3113), .S(n3060), .Z(n485) );
  MUX21L U2045 ( .A(n1707), .B(n3114), .S(n3059), .Z(n486) );
  MUX21L U2046 ( .A(n1708), .B(n3115), .S(n3059), .Z(n487) );
  MUX21L U2047 ( .A(n1709), .B(n3116), .S(n3059), .Z(n488) );
  MUX21L U2048 ( .A(n1710), .B(n3117), .S(n3059), .Z(n489) );
  MUX21L U2049 ( .A(n1711), .B(n3118), .S(n3059), .Z(n490) );
  MUX21L U2050 ( .A(n1712), .B(n3121), .S(n3059), .Z(n491) );
  MUX21L U2051 ( .A(n1713), .B(n3122), .S(n3059), .Z(n492) );
  MUX21L U2052 ( .A(n1714), .B(n3123), .S(n3059), .Z(n493) );
  MUX21L U2053 ( .A(n1715), .B(n3124), .S(n3059), .Z(n494) );
  MUX21L U2054 ( .A(n1716), .B(n3125), .S(n3059), .Z(n495) );
  MUX21L U2055 ( .A(n1717), .B(n3126), .S(n3059), .Z(n496) );
  MUX21L U2056 ( .A(n1718), .B(n3127), .S(n3059), .Z(n497) );
  MUX21L U2057 ( .A(n1719), .B(n3129), .S(n3059), .Z(n498) );
  MUX21L U2058 ( .A(n1720), .B(n3133), .S(n3059), .Z(n499) );
  ND2I U2059 ( .A(n2103), .B(n2104), .Z(n3256) );
  MUX21L U2060 ( .A(n1721), .B(n3089), .S(n3064), .Z(n436) );
  MUX21L U2061 ( .A(n1722), .B(n3091), .S(n3064), .Z(n437) );
  MUX21L U2062 ( .A(n3257), .B(n3093), .S(n3064), .Z(n438) );
  MUX21L U2063 ( .A(n1723), .B(n3095), .S(n3064), .Z(n439) );
  MUX21L U2064 ( .A(n1724), .B(n3097), .S(n3063), .Z(n440) );
  MUX21L U2065 ( .A(n1725), .B(n3099), .S(n3063), .Z(n441) );
  MUX21L U2066 ( .A(n1726), .B(n3100), .S(n3063), .Z(n442) );
  MUX21L U2067 ( .A(n1727), .B(n3101), .S(n3063), .Z(n443) );
  MUX21L U2068 ( .A(n1728), .B(n3102), .S(n3063), .Z(n444) );
  MUX21L U2069 ( .A(n1729), .B(n3103), .S(n3063), .Z(n445) );
  MUX21L U2070 ( .A(n1730), .B(n3104), .S(n3063), .Z(n446) );
  MUX21L U2071 ( .A(n1731), .B(n3105), .S(n3063), .Z(n447) );
  MUX21L U2072 ( .A(n1732), .B(n3106), .S(n3063), .Z(n448) );
  MUX21L U2073 ( .A(n1733), .B(n3107), .S(n3063), .Z(n449) );
  MUX21L U2074 ( .A(n1734), .B(n3108), .S(n3063), .Z(n450) );
  MUX21L U2075 ( .A(n1735), .B(n3110), .S(n3063), .Z(n451) );
  MUX21L U2076 ( .A(n1736), .B(n3111), .S(n3063), .Z(n452) );
  MUX21L U2077 ( .A(n1737), .B(n3113), .S(n3063), .Z(n453) );
  MUX21L U2078 ( .A(n1738), .B(n3114), .S(n3062), .Z(n454) );
  MUX21L U2079 ( .A(n1739), .B(n3115), .S(n3062), .Z(n455) );
  MUX21L U2080 ( .A(n1740), .B(n3116), .S(n3062), .Z(n456) );
  MUX21L U2081 ( .A(n1741), .B(n3117), .S(n3062), .Z(n457) );
  MUX21L U2082 ( .A(n1742), .B(n3118), .S(n3062), .Z(n458) );
  MUX21L U2083 ( .A(n1743), .B(n3121), .S(n3062), .Z(n459) );
  MUX21L U2084 ( .A(n1744), .B(n3122), .S(n3062), .Z(n460) );
  MUX21L U2085 ( .A(n1745), .B(n3123), .S(n3062), .Z(n461) );
  MUX21L U2086 ( .A(n1746), .B(n3124), .S(n3062), .Z(n462) );
  MUX21L U2087 ( .A(n1747), .B(n3125), .S(n3062), .Z(n463) );
  MUX21L U2088 ( .A(n1748), .B(n3126), .S(n3062), .Z(n464) );
  MUX21L U2089 ( .A(n1749), .B(n3127), .S(n3062), .Z(n465) );
  MUX21L U2090 ( .A(n1750), .B(n3129), .S(n3062), .Z(n466) );
  MUX21L U2091 ( .A(n1751), .B(n3133), .S(n3062), .Z(n467) );
  ND2I U2092 ( .A(n2103), .B(n1179), .Z(n3258) );
  MUX21L U2093 ( .A(n1752), .B(n3089), .S(n3067), .Z(n404) );
  MUX21L U2094 ( .A(n1753), .B(n3091), .S(n3067), .Z(n405) );
  MUX21L U2095 ( .A(n3259), .B(n3093), .S(n3067), .Z(n406) );
  MUX21L U2096 ( .A(n1754), .B(n3095), .S(n3067), .Z(n407) );
  MUX21L U2097 ( .A(n1755), .B(n3097), .S(n3066), .Z(n408) );
  MUX21L U2098 ( .A(n1756), .B(n3099), .S(n3066), .Z(n409) );
  MUX21L U2099 ( .A(n1757), .B(n3100), .S(n3066), .Z(n410) );
  MUX21L U2100 ( .A(n1758), .B(n3101), .S(n3066), .Z(n411) );
  MUX21L U2101 ( .A(n1759), .B(n3102), .S(n3066), .Z(n412) );
  MUX21L U2102 ( .A(n1760), .B(n3103), .S(n3066), .Z(n413) );
  MUX21L U2103 ( .A(n1761), .B(n3104), .S(n3066), .Z(n414) );
  MUX21L U2104 ( .A(n1762), .B(n3105), .S(n3066), .Z(n415) );
  MUX21L U2105 ( .A(n1763), .B(n3106), .S(n3066), .Z(n416) );
  MUX21L U2106 ( .A(n1764), .B(n3107), .S(n3066), .Z(n417) );
  MUX21L U2107 ( .A(n1765), .B(n3108), .S(n3066), .Z(n418) );
  MUX21L U2108 ( .A(n1766), .B(n3110), .S(n3066), .Z(n419) );
  MUX21L U2109 ( .A(n1767), .B(n3111), .S(n3066), .Z(n420) );
  MUX21L U2110 ( .A(n1768), .B(n3113), .S(n3066), .Z(n421) );
  MUX21L U2111 ( .A(n1769), .B(n3114), .S(n3065), .Z(n422) );
  MUX21L U2112 ( .A(n1770), .B(n3115), .S(n3065), .Z(n423) );
  MUX21L U2113 ( .A(n1771), .B(n3116), .S(n3065), .Z(n424) );
  MUX21L U2114 ( .A(n1772), .B(n3117), .S(n3065), .Z(n425) );
  MUX21L U2115 ( .A(n1773), .B(n3118), .S(n3065), .Z(n426) );
  MUX21L U2116 ( .A(n1774), .B(n3121), .S(n3065), .Z(n427) );
  MUX21L U2117 ( .A(n1775), .B(n3122), .S(n3065), .Z(n428) );
  MUX21L U2118 ( .A(n1776), .B(n3123), .S(n3065), .Z(n429) );
  MUX21L U2119 ( .A(n1777), .B(n3124), .S(n3065), .Z(n430) );
  MUX21L U2120 ( .A(n1778), .B(n3125), .S(n3065), .Z(n431) );
  MUX21L U2121 ( .A(n1779), .B(n3126), .S(n3065), .Z(n432) );
  MUX21L U2122 ( .A(n1780), .B(n3127), .S(n3065), .Z(n433) );
  MUX21L U2123 ( .A(n1781), .B(n3129), .S(n3065), .Z(n434) );
  MUX21L U2124 ( .A(n1782), .B(n3133), .S(n3065), .Z(n435) );
  MUX21L U2125 ( .A(n56), .B(n3089), .S(n3070), .Z(n372) );
  MUX21L U2126 ( .A(n57), .B(n3091), .S(n3070), .Z(n373) );
  MUX21L U2127 ( .A(n58), .B(n3093), .S(n3070), .Z(n374) );
  MUX21L U2128 ( .A(n1783), .B(n3095), .S(n3070), .Z(n375) );
  MUX21L U2129 ( .A(n1784), .B(n3097), .S(n3069), .Z(n376) );
  MUX21L U2130 ( .A(n1785), .B(n3099), .S(n3069), .Z(n377) );
  MUX21L U2131 ( .A(n1786), .B(n3100), .S(n3069), .Z(n378) );
  MUX21L U2132 ( .A(n1787), .B(n3101), .S(n3069), .Z(n379) );
  MUX21L U2133 ( .A(n1788), .B(n3102), .S(n3069), .Z(n380) );
  MUX21L U2134 ( .A(n1789), .B(n3103), .S(n3069), .Z(n381) );
  MUX21L U2135 ( .A(n1790), .B(n3104), .S(n3069), .Z(n382) );
  MUX21L U2136 ( .A(n1791), .B(n3105), .S(n3069), .Z(n383) );
  MUX21L U2137 ( .A(n1792), .B(n3106), .S(n3069), .Z(n384) );
  MUX21L U2138 ( .A(n1793), .B(n3107), .S(n3069), .Z(n385) );
  MUX21L U2139 ( .A(n1794), .B(n3108), .S(n3069), .Z(n386) );
  MUX21L U2140 ( .A(n1795), .B(n3110), .S(n3069), .Z(n387) );
  MUX21L U2141 ( .A(n1796), .B(n3111), .S(n3069), .Z(n388) );
  MUX21L U2142 ( .A(n1797), .B(n3113), .S(n3069), .Z(n389) );
  MUX21L U2143 ( .A(n1798), .B(n3114), .S(n3068), .Z(n390) );
  MUX21L U2144 ( .A(n1799), .B(n3115), .S(n3068), .Z(n391) );
  MUX21L U2145 ( .A(n1800), .B(n3116), .S(n3068), .Z(n392) );
  MUX21L U2146 ( .A(n1801), .B(n3117), .S(n3068), .Z(n393) );
  MUX21L U2147 ( .A(n1802), .B(n3118), .S(n3068), .Z(n394) );
  MUX21L U2148 ( .A(n1803), .B(n3121), .S(n3068), .Z(n395) );
  MUX21L U2149 ( .A(n1804), .B(n3122), .S(n3068), .Z(n396) );
  MUX21L U2150 ( .A(n1805), .B(n3123), .S(n3068), .Z(n397) );
  MUX21L U2151 ( .A(n1806), .B(n3124), .S(n3068), .Z(n398) );
  MUX21L U2152 ( .A(n1807), .B(n3125), .S(n3068), .Z(n399) );
  MUX21L U2153 ( .A(n1808), .B(n3126), .S(n3068), .Z(n400) );
  MUX21L U2154 ( .A(n1809), .B(n3127), .S(n3068), .Z(n401) );
  MUX21L U2155 ( .A(n1810), .B(n3129), .S(n3068), .Z(n402) );
  MUX21L U2156 ( .A(n1811), .B(n3133), .S(n3068), .Z(n403) );
  ND2I U2157 ( .A(n2112), .B(n2105), .Z(n3260) );
  MUX21L U2158 ( .A(n125), .B(n3089), .S(n3073), .Z(n340) );
  MUX21L U2159 ( .A(n126), .B(n3091), .S(n3073), .Z(n341) );
  MUX21L U2160 ( .A(n127), .B(n3093), .S(n3073), .Z(n342) );
  MUX21L U2161 ( .A(n1812), .B(n3095), .S(n3073), .Z(n343) );
  MUX21L U2162 ( .A(n1813), .B(n3097), .S(n3072), .Z(n344) );
  MUX21L U2163 ( .A(n3261), .B(n3099), .S(n3072), .Z(n345) );
  MUX21L U2164 ( .A(n1814), .B(n3100), .S(n3072), .Z(n346) );
  MUX21L U2165 ( .A(n1815), .B(n3101), .S(n3072), .Z(n347) );
  MUX21L U2166 ( .A(n1816), .B(n3102), .S(n3072), .Z(n348) );
  MUX21L U2167 ( .A(n3262), .B(n3103), .S(n3072), .Z(n349) );
  MUX21L U2168 ( .A(n1817), .B(n3104), .S(n3072), .Z(n350) );
  MUX21L U2169 ( .A(n1818), .B(n3105), .S(n3072), .Z(n351) );
  MUX21L U2170 ( .A(n1819), .B(n3106), .S(n3072), .Z(n352) );
  MUX21L U2171 ( .A(n1820), .B(n3107), .S(n3072), .Z(n353) );
  MUX21L U2172 ( .A(n1821), .B(n3108), .S(n3072), .Z(n354) );
  MUX21L U2173 ( .A(n1822), .B(n3110), .S(n3072), .Z(n355) );
  MUX21L U2174 ( .A(n1823), .B(n3111), .S(n3072), .Z(n356) );
  MUX21L U2175 ( .A(n1824), .B(n3113), .S(n3072), .Z(n357) );
  MUX21L U2176 ( .A(n1825), .B(n3114), .S(n3071), .Z(n358) );
  MUX21L U2177 ( .A(n1826), .B(n3115), .S(n3071), .Z(n359) );
  MUX21L U2178 ( .A(n1827), .B(n3116), .S(n3071), .Z(n360) );
  MUX21L U2179 ( .A(n1828), .B(n3117), .S(n3071), .Z(n361) );
  MUX21L U2180 ( .A(n1829), .B(n3118), .S(n3071), .Z(n362) );
  MUX21L U2181 ( .A(n1830), .B(n3121), .S(n3071), .Z(n363) );
  MUX21L U2182 ( .A(n1831), .B(n3122), .S(n3071), .Z(n364) );
  MUX21L U2183 ( .A(n1832), .B(n3123), .S(n3071), .Z(n365) );
  MUX21L U2184 ( .A(n1833), .B(n3124), .S(n3071), .Z(n366) );
  MUX21L U2185 ( .A(n1834), .B(n3125), .S(n3071), .Z(n367) );
  MUX21L U2186 ( .A(n1835), .B(n3126), .S(n3071), .Z(n368) );
  MUX21L U2187 ( .A(n1836), .B(n3127), .S(n3071), .Z(n369) );
  MUX21L U2188 ( .A(n1837), .B(n3129), .S(n3071), .Z(n370) );
  MUX21L U2189 ( .A(n1838), .B(n3133), .S(n3071), .Z(n371) );
  ND2I U2190 ( .A(n2109), .B(n2105), .Z(n3263) );
  MUX21L U2191 ( .A(n1839), .B(n3089), .S(n3076), .Z(n308) );
  MUX21L U2192 ( .A(n1840), .B(n3091), .S(n3076), .Z(n309) );
  MUX21L U2193 ( .A(n3264), .B(n3093), .S(n3076), .Z(n310) );
  MUX21L U2194 ( .A(n1841), .B(n3095), .S(n3076), .Z(n311) );
  MUX21L U2195 ( .A(n1842), .B(n3097), .S(n3075), .Z(n312) );
  MUX21L U2196 ( .A(n1843), .B(n3099), .S(n3075), .Z(n313) );
  MUX21L U2197 ( .A(n1844), .B(n3100), .S(n3075), .Z(n314) );
  MUX21L U2198 ( .A(n1845), .B(n3101), .S(n3075), .Z(n315) );
  MUX21L U2199 ( .A(n1846), .B(n3102), .S(n3075), .Z(n316) );
  MUX21L U2200 ( .A(n1847), .B(n3103), .S(n3075), .Z(n317) );
  MUX21L U2201 ( .A(n1848), .B(n3104), .S(n3075), .Z(n318) );
  MUX21L U2202 ( .A(n1849), .B(n3105), .S(n3075), .Z(n319) );
  MUX21L U2203 ( .A(n1850), .B(n3106), .S(n3075), .Z(n320) );
  MUX21L U2204 ( .A(n1851), .B(n3107), .S(n3075), .Z(n321) );
  MUX21L U2205 ( .A(n1852), .B(n3108), .S(n3075), .Z(n322) );
  MUX21L U2206 ( .A(n1853), .B(n3110), .S(n3075), .Z(n323) );
  MUX21L U2207 ( .A(n1854), .B(n3111), .S(n3075), .Z(n324) );
  MUX21L U2208 ( .A(n1855), .B(n3113), .S(n3075), .Z(n325) );
  MUX21L U2209 ( .A(n1856), .B(n3114), .S(n3074), .Z(n326) );
  MUX21L U2210 ( .A(n1857), .B(n3115), .S(n3074), .Z(n327) );
  MUX21L U2211 ( .A(n1858), .B(n3116), .S(n3074), .Z(n328) );
  MUX21L U2212 ( .A(n1859), .B(n3117), .S(n3074), .Z(n329) );
  MUX21L U2213 ( .A(n1860), .B(n3118), .S(n3074), .Z(n330) );
  MUX21L U2214 ( .A(n1861), .B(n3121), .S(n3074), .Z(n331) );
  MUX21L U2215 ( .A(n1862), .B(n3122), .S(n3074), .Z(n332) );
  MUX21L U2216 ( .A(n1863), .B(n3123), .S(n3074), .Z(n333) );
  MUX21L U2217 ( .A(n1864), .B(n3124), .S(n3074), .Z(n334) );
  MUX21L U2218 ( .A(n1865), .B(n3125), .S(n3074), .Z(n335) );
  MUX21L U2219 ( .A(n1866), .B(n3126), .S(n3074), .Z(n336) );
  MUX21L U2220 ( .A(n1867), .B(n3127), .S(n3074), .Z(n337) );
  MUX21L U2221 ( .A(n1868), .B(n3129), .S(n3074), .Z(n338) );
  MUX21L U2222 ( .A(n1869), .B(n3133), .S(n3074), .Z(n339) );
  ND2I U2223 ( .A(n2111), .B(n2105), .Z(n3265) );
  MUX21L U2224 ( .A(n1870), .B(n3089), .S(n3079), .Z(n276) );
  MUX21L U2225 ( .A(n1871), .B(n3091), .S(n3079), .Z(n277) );
  MUX21L U2226 ( .A(n2092), .B(n3093), .S(n3079), .Z(n278) );
  MUX21L U2227 ( .A(n1872), .B(n3095), .S(n3079), .Z(n279) );
  MUX21L U2228 ( .A(n1873), .B(n3097), .S(n3078), .Z(n280) );
  MUX21L U2229 ( .A(n1874), .B(n3099), .S(n3078), .Z(n281) );
  MUX21L U2230 ( .A(n1875), .B(n3100), .S(n3078), .Z(n282) );
  MUX21L U2231 ( .A(n1876), .B(n3101), .S(n3078), .Z(n283) );
  MUX21L U2232 ( .A(n1877), .B(n3102), .S(n3078), .Z(n284) );
  MUX21L U2233 ( .A(n1878), .B(n3103), .S(n3078), .Z(n285) );
  MUX21L U2234 ( .A(n1879), .B(n3104), .S(n3078), .Z(n286) );
  MUX21L U2235 ( .A(n1880), .B(n3105), .S(n3078), .Z(n287) );
  MUX21L U2236 ( .A(n1881), .B(n3106), .S(n3078), .Z(n288) );
  MUX21L U2237 ( .A(n1882), .B(n3107), .S(n3078), .Z(n289) );
  MUX21L U2238 ( .A(n1883), .B(n3108), .S(n3078), .Z(n290) );
  MUX21L U2239 ( .A(n1884), .B(n3110), .S(n3078), .Z(n291) );
  MUX21L U2240 ( .A(n1885), .B(n3111), .S(n3078), .Z(n292) );
  MUX21L U2241 ( .A(n1886), .B(n3113), .S(n3078), .Z(n293) );
  MUX21L U2242 ( .A(n1887), .B(n3114), .S(n3077), .Z(n294) );
  MUX21L U2243 ( .A(n1888), .B(n3115), .S(n3077), .Z(n295) );
  MUX21L U2244 ( .A(n1889), .B(n3116), .S(n3077), .Z(n296) );
  MUX21L U2245 ( .A(n1890), .B(n3117), .S(n3077), .Z(n297) );
  MUX21L U2246 ( .A(n1891), .B(n3118), .S(n3077), .Z(n298) );
  MUX21L U2247 ( .A(n1892), .B(n3121), .S(n3077), .Z(n299) );
  MUX21L U2248 ( .A(n1893), .B(n3122), .S(n3077), .Z(n300) );
  MUX21L U2249 ( .A(n1894), .B(n3123), .S(n3077), .Z(n301) );
  MUX21L U2250 ( .A(n1895), .B(n3124), .S(n3077), .Z(n302) );
  MUX21L U2251 ( .A(n1896), .B(n3125), .S(n3077), .Z(n303) );
  MUX21L U2252 ( .A(n1897), .B(n3126), .S(n3077), .Z(n304) );
  MUX21L U2253 ( .A(n1898), .B(n3127), .S(n3077), .Z(n305) );
  MUX21L U2254 ( .A(n1899), .B(n3129), .S(n3077), .Z(n306) );
  MUX21L U2255 ( .A(n1900), .B(n3133), .S(n3077), .Z(n307) );
  ND2I U2256 ( .A(n2108), .B(n2105), .Z(n3266) );
  MUX21L U2257 ( .A(n1901), .B(n3089), .S(n3082), .Z(n244) );
  MUX21L U2258 ( .A(n1902), .B(n3091), .S(n3082), .Z(n245) );
  MUX21L U2259 ( .A(n1903), .B(n3093), .S(n3082), .Z(n246) );
  MUX21L U2260 ( .A(n1904), .B(n3095), .S(n3082), .Z(n247) );
  MUX21L U2261 ( .A(n1905), .B(n3097), .S(n3081), .Z(n248) );
  MUX21L U2262 ( .A(n1906), .B(n3099), .S(n3081), .Z(n249) );
  MUX21L U2263 ( .A(n1907), .B(n3100), .S(n3081), .Z(n250) );
  MUX21L U2264 ( .A(n1908), .B(n3101), .S(n3081), .Z(n251) );
  MUX21L U2265 ( .A(n1909), .B(n3102), .S(n3081), .Z(n252) );
  MUX21L U2266 ( .A(n1910), .B(n3103), .S(n3081), .Z(n253) );
  MUX21L U2267 ( .A(n1911), .B(n3104), .S(n3081), .Z(n254) );
  MUX21L U2268 ( .A(n1912), .B(n3105), .S(n3081), .Z(n255) );
  MUX21L U2269 ( .A(n1913), .B(n3106), .S(n3081), .Z(n256) );
  MUX21L U2270 ( .A(n1914), .B(n3107), .S(n3081), .Z(n257) );
  MUX21L U2271 ( .A(n3267), .B(n3108), .S(n3081), .Z(n258) );
  MUX21L U2272 ( .A(n1915), .B(n3110), .S(n3081), .Z(n259) );
  MUX21L U2273 ( .A(n1916), .B(n3111), .S(n3081), .Z(n260) );
  MUX21L U2274 ( .A(n1917), .B(n3113), .S(n3081), .Z(n261) );
  MUX21L U2275 ( .A(n1918), .B(n3114), .S(n3080), .Z(n262) );
  MUX21L U2276 ( .A(n1919), .B(n3115), .S(n3080), .Z(n263) );
  MUX21L U2277 ( .A(n1920), .B(n3116), .S(n3080), .Z(n264) );
  MUX21L U2278 ( .A(n1921), .B(n3117), .S(n3080), .Z(n265) );
  MUX21L U2279 ( .A(n1922), .B(n3118), .S(n3080), .Z(n266) );
  MUX21L U2280 ( .A(n1923), .B(n3121), .S(n3080), .Z(n267) );
  MUX21L U2281 ( .A(n1924), .B(n3122), .S(n3080), .Z(n268) );
  MUX21L U2282 ( .A(n1925), .B(n3123), .S(n3080), .Z(n269) );
  MUX21L U2283 ( .A(n1926), .B(n3124), .S(n3080), .Z(n270) );
  MUX21L U2284 ( .A(n1927), .B(n3125), .S(n3080), .Z(n271) );
  MUX21L U2285 ( .A(n1928), .B(n3126), .S(n3080), .Z(n272) );
  MUX21L U2286 ( .A(n1929), .B(n3127), .S(n3080), .Z(n273) );
  MUX21L U2287 ( .A(n1930), .B(n3129), .S(n3080), .Z(n274) );
  MUX21L U2288 ( .A(n1931), .B(n3133), .S(n3080), .Z(n275) );
  ND2I U2289 ( .A(n2110), .B(n2105), .Z(n3268) );
  MUX21L U2290 ( .A(n1932), .B(n3089), .S(n3085), .Z(n212) );
  MUX21L U2291 ( .A(n1933), .B(n3091), .S(n3085), .Z(n213) );
  MUX21L U2292 ( .A(n1934), .B(n3093), .S(n3085), .Z(n214) );
  MUX21L U2293 ( .A(n1935), .B(n3095), .S(n3085), .Z(n215) );
  MUX21L U2294 ( .A(n1936), .B(n3097), .S(n3084), .Z(n216) );
  MUX21L U2295 ( .A(n1937), .B(n3099), .S(n3084), .Z(n217) );
  MUX21L U2296 ( .A(n1938), .B(n3100), .S(n3084), .Z(n218) );
  MUX21L U2297 ( .A(n1939), .B(n3101), .S(n3084), .Z(n219) );
  MUX21L U2298 ( .A(n1940), .B(n3102), .S(n3084), .Z(n220) );
  MUX21L U2299 ( .A(n1941), .B(n3103), .S(n3084), .Z(n221) );
  MUX21L U2300 ( .A(n1942), .B(n3104), .S(n3084), .Z(n222) );
  MUX21L U2301 ( .A(n1943), .B(n3105), .S(n3084), .Z(n223) );
  MUX21L U2302 ( .A(n1944), .B(n3106), .S(n3084), .Z(n224) );
  MUX21L U2303 ( .A(n1945), .B(n3107), .S(n3084), .Z(n225) );
  MUX21L U2304 ( .A(n1946), .B(n3108), .S(n3084), .Z(n226) );
  MUX21L U2305 ( .A(n1947), .B(n3110), .S(n3084), .Z(n227) );
  MUX21L U2306 ( .A(n1948), .B(n3111), .S(n3084), .Z(n228) );
  MUX21L U2307 ( .A(n1949), .B(n3113), .S(n3084), .Z(n229) );
  MUX21L U2308 ( .A(n1950), .B(n3114), .S(n3083), .Z(n230) );
  MUX21L U2309 ( .A(n1951), .B(n3115), .S(n3083), .Z(n231) );
  MUX21L U2310 ( .A(n1952), .B(n3116), .S(n3083), .Z(n232) );
  MUX21L U2311 ( .A(n1953), .B(n3117), .S(n3083), .Z(n233) );
  MUX21L U2312 ( .A(n1954), .B(n3118), .S(n3083), .Z(n234) );
  MUX21L U2313 ( .A(n1955), .B(n3121), .S(n3083), .Z(n235) );
  MUX21L U2314 ( .A(n1956), .B(n3122), .S(n3083), .Z(n236) );
  MUX21L U2315 ( .A(n1957), .B(n3123), .S(n3083), .Z(n237) );
  MUX21L U2316 ( .A(n1958), .B(n3124), .S(n3083), .Z(n238) );
  MUX21L U2317 ( .A(n1959), .B(n3125), .S(n3083), .Z(n239) );
  MUX21L U2318 ( .A(n1960), .B(n3126), .S(n3083), .Z(n240) );
  MUX21L U2319 ( .A(n1961), .B(n3127), .S(n3083), .Z(n241) );
  MUX21L U2320 ( .A(n1962), .B(n3129), .S(n3083), .Z(n242) );
  MUX21L U2321 ( .A(n1963), .B(n3133), .S(n3083), .Z(n243) );
  ND2I U2322 ( .A(n2104), .B(n2105), .Z(n3269) );
  MUX21L U2323 ( .A(n131), .B(n3089), .S(n3088), .Z(n180) );
  MUX21L U2324 ( .A(n134), .B(n3091), .S(n3088), .Z(n181) );
  MUX21L U2325 ( .A(n137), .B(n3093), .S(n3088), .Z(n182) );
  MUX21L U2326 ( .A(n1964), .B(n3095), .S(n3088), .Z(n183) );
  MUX21L U2327 ( .A(n3270), .B(n3097), .S(n3087), .Z(n184) );
  MUX21L U2328 ( .A(n1965), .B(n3099), .S(n3087), .Z(n185) );
  MUX21L U2329 ( .A(n1966), .B(n3100), .S(n3087), .Z(n186) );
  MUX21L U2330 ( .A(n3271), .B(n3101), .S(n3087), .Z(n187) );
  MUX21L U2331 ( .A(n1967), .B(n3102), .S(n3087), .Z(n188) );
  MUX21L U2332 ( .A(n3272), .B(n3103), .S(n3087), .Z(n189) );
  MUX21L U2333 ( .A(n1968), .B(n3104), .S(n3087), .Z(n190) );
  MUX21L U2334 ( .A(n1969), .B(n3105), .S(n3087), .Z(n191) );
  MUX21L U2335 ( .A(n1970), .B(n3106), .S(n3087), .Z(n192) );
  MUX21L U2336 ( .A(n1971), .B(n3107), .S(n3087), .Z(n193) );
  MUX21L U2337 ( .A(n3273), .B(n3108), .S(n3087), .Z(n194) );
  MUX21L U2338 ( .A(n1972), .B(n3110), .S(n3087), .Z(n195) );
  MUX21L U2339 ( .A(n1973), .B(n3111), .S(n3087), .Z(n196) );
  MUX21L U2340 ( .A(n1974), .B(n3113), .S(n3087), .Z(n197) );
  MUX21L U2341 ( .A(n1975), .B(n3114), .S(n3086), .Z(n198) );
  MUX21L U2342 ( .A(n1976), .B(n3115), .S(n3086), .Z(n199) );
  MUX21L U2343 ( .A(n1977), .B(n3116), .S(n3086), .Z(n200) );
  MUX21L U2344 ( .A(n1978), .B(n3117), .S(n3086), .Z(n201) );
  MUX21L U2345 ( .A(n1979), .B(n3118), .S(n3086), .Z(n202) );
  MUX21L U2346 ( .A(n1980), .B(n3121), .S(n3086), .Z(n203) );
  MUX21L U2347 ( .A(n1981), .B(n3122), .S(n3086), .Z(n204) );
  MUX21L U2348 ( .A(n1982), .B(n3123), .S(n3086), .Z(n205) );
  MUX21L U2349 ( .A(n1983), .B(n3124), .S(n3086), .Z(n206) );
  MUX21L U2350 ( .A(n1984), .B(n3125), .S(n3086), .Z(n207) );
  MUX21L U2351 ( .A(n1985), .B(n3126), .S(n3086), .Z(n208) );
  MUX21L U2352 ( .A(n1986), .B(n3127), .S(n3086), .Z(n209) );
  MUX21L U2353 ( .A(n1987), .B(n3129), .S(n3086), .Z(n210) );
  MUX21L U2354 ( .A(n1988), .B(n3133), .S(n3086), .Z(n211) );
  ND2I U2355 ( .A(n1179), .B(n2105), .Z(n3274) );
  MUX21L U2356 ( .A(n62), .B(n3089), .S(n3132), .Z(n148) );
  MUX21L U2357 ( .A(n65), .B(n3091), .S(n3132), .Z(n149) );
  MUX21L U2358 ( .A(n68), .B(n3093), .S(n3132), .Z(n150) );
  MUX21L U2359 ( .A(n1989), .B(n3095), .S(n3132), .Z(n151) );
  MUX21L U2360 ( .A(n1990), .B(n3097), .S(n3131), .Z(n152) );
  MUX21L U2361 ( .A(n1991), .B(n3099), .S(n3131), .Z(n153) );
  MUX21L U2362 ( .A(n1992), .B(n3100), .S(n3131), .Z(n154) );
  MUX21L U2363 ( .A(n1993), .B(n3101), .S(n3131), .Z(n155) );
  MUX21L U2364 ( .A(n1994), .B(n3102), .S(n3131), .Z(n156) );
  MUX21L U2365 ( .A(n1995), .B(n3103), .S(n3131), .Z(n157) );
  MUX21L U2366 ( .A(n1996), .B(n3104), .S(n3131), .Z(n158) );
  MUX21L U2367 ( .A(n1997), .B(n3105), .S(n3131), .Z(n159) );
  MUX21L U2368 ( .A(n1998), .B(n3106), .S(n3131), .Z(n160) );
  MUX21L U2369 ( .A(n1999), .B(n3107), .S(n3131), .Z(n161) );
  MUX21L U2370 ( .A(n2000), .B(n3108), .S(n3131), .Z(n162) );
  MUX21L U2371 ( .A(n2001), .B(n3110), .S(n3131), .Z(n163) );
  MUX21L U2372 ( .A(n2002), .B(n3111), .S(n3131), .Z(n164) );
  MUX21L U2373 ( .A(n2003), .B(n3113), .S(n3131), .Z(n165) );
  MUX21L U2374 ( .A(n2004), .B(n3114), .S(n3130), .Z(n166) );
  MUX21L U2375 ( .A(n2005), .B(n3115), .S(n3130), .Z(n167) );
  MUX21L U2376 ( .A(n2006), .B(n3116), .S(n3130), .Z(n168) );
  MUX21L U2377 ( .A(n2007), .B(n3117), .S(n3130), .Z(n169) );
  MUX21L U2378 ( .A(n2008), .B(n3118), .S(n3130), .Z(n170) );
  MUX21L U2379 ( .A(n2009), .B(n3121), .S(n3130), .Z(n171) );
  MUX21L U2380 ( .A(n2010), .B(n3122), .S(n3130), .Z(n172) );
  MUX21L U2381 ( .A(n2011), .B(n3123), .S(n3130), .Z(n173) );
  MUX21L U2382 ( .A(n2012), .B(n3124), .S(n3130), .Z(n174) );
  MUX21L U2383 ( .A(n2013), .B(n3125), .S(n3130), .Z(n175) );
  MUX21L U2384 ( .A(n2014), .B(n3126), .S(n3130), .Z(n176) );
  MUX21L U2385 ( .A(n2015), .B(n3127), .S(n3130), .Z(n177) );
  MUX21L U2386 ( .A(n2016), .B(n3129), .S(n3130), .Z(n178) );
  MUX21L U2387 ( .A(n2017), .B(n3133), .S(n3130), .Z(n179) );
  NR2I U2388 ( .A(N21), .B(N22), .Z(n3275) );
  AN2I U2389 ( .A(N120), .B(n3134), .Z(rd_data2[0]) );
  AN2I U2390 ( .A(N119), .B(n3134), .Z(rd_data2[1]) );
  AN2I U2391 ( .A(N118), .B(n3134), .Z(rd_data2[2]) );
  AN2I U2392 ( .A(N117), .B(n3134), .Z(rd_data2[3]) );
  AN2I U2393 ( .A(N116), .B(n3134), .Z(rd_data2[4]) );
  AN2I U2394 ( .A(N115), .B(n3134), .Z(rd_data2[5]) );
  AN2I U2395 ( .A(N114), .B(n3134), .Z(rd_data2[6]) );
  AN2I U2396 ( .A(N113), .B(n3134), .Z(rd_data2[7]) );
  AN2I U2397 ( .A(N112), .B(n3134), .Z(rd_data2[8]) );
  AN2I U2398 ( .A(N111), .B(n3134), .Z(rd_data2[9]) );
  AN2I U2399 ( .A(N110), .B(n3134), .Z(rd_data2[10]) );
  AN2I U2400 ( .A(N109), .B(n3134), .Z(rd_data2[11]) );
  AN2I U2401 ( .A(N108), .B(n3134), .Z(rd_data2[12]) );
  AN2I U2402 ( .A(N107), .B(n3134), .Z(rd_data2[13]) );
  AN2I U2403 ( .A(N106), .B(n3134), .Z(rd_data2[14]) );
  AN2I U2404 ( .A(N105), .B(n3134), .Z(rd_data2[15]) );
  AN2I U2405 ( .A(N104), .B(n3134), .Z(rd_data2[16]) );
  AN2I U2406 ( .A(N103), .B(n3134), .Z(rd_data2[17]) );
  AN2I U2407 ( .A(N102), .B(n3134), .Z(rd_data2[18]) );
  AN2I U2408 ( .A(N101), .B(n3134), .Z(rd_data2[19]) );
  AN2I U2409 ( .A(N100), .B(n3134), .Z(rd_data2[20]) );
  AN2I U2410 ( .A(N99), .B(n3134), .Z(rd_data2[21]) );
  AN2I U2411 ( .A(N98), .B(n3134), .Z(rd_data2[22]) );
  AN2I U2412 ( .A(N97), .B(n3134), .Z(rd_data2[23]) );
  AN2I U2413 ( .A(N96), .B(n3134), .Z(rd_data2[24]) );
  AN2I U2414 ( .A(N95), .B(n3134), .Z(rd_data2[25]) );
  AN2I U2415 ( .A(N94), .B(n3134), .Z(rd_data2[26]) );
  AN2I U2416 ( .A(N93), .B(n3134), .Z(rd_data2[27]) );
  AN2I U2417 ( .A(N92), .B(n3134), .Z(rd_data2[28]) );
  AN2I U2418 ( .A(N91), .B(n3134), .Z(rd_data2[29]) );
  AN2I U2419 ( .A(N90), .B(n3134), .Z(rd_data2[30]) );
  AN2I U2420 ( .A(N89), .B(n3134), .Z(rd_data2[31]) );
  MUX21L U2421 ( .A(\gpr[6][0] ), .B(\gpr[7][0] ), .S(n3153), .Z(n3277) );
  NR2I U2422 ( .A(n3214), .B(n3278), .Z(n3304) );
  IVI U2423 ( .A(N16), .Z(n3293) );
  IVI U2424 ( .A(N17), .Z(n3291) );
  ND2I U2425 ( .A(n3293), .B(n3291), .Z(n4451) );
  ND2I U2426 ( .A(n3212), .B(n3291), .Z(n3279) );
  MUX21L U2427 ( .A(\gpr[10][0] ), .B(\gpr[11][0] ), .S(n2088), .Z(n3280) );
  MUX21L U2428 ( .A(n131), .B(n62), .S(n2071), .Z(n3281) );
  ND2I U2429 ( .A(n3206), .B(n3293), .Z(n3282) );
  MUX21L U2430 ( .A(\gpr[22][0] ), .B(\gpr[23][0] ), .S(n2037), .Z(n3283) );
  ND2I U2431 ( .A(n115), .B(n3213), .Z(n3284) );
  MUX21L U2432 ( .A(\gpr[26][0] ), .B(\gpr[27][0] ), .S(n2034), .Z(n3285) );
  MUX21L U2433 ( .A(n132), .B(n63), .S(n3172), .Z(n3290) );
  MUX21L U2434 ( .A(n133), .B(n64), .S(n3170), .Z(n3292) );
  ND2I U2435 ( .A(n3293), .B(n3213), .Z(n4459) );
  AO1P U2436 ( .A(n3145), .B(n3298), .C(n3297), .D(n3296), .Z(n3303) );
  NR2I U2437 ( .A(n2082), .B(n1159), .Z(n3300) );
  MUX21L U2438 ( .A(n147), .B(n81), .S(n3174), .Z(n3299) );
  MUX21L U2439 ( .A(n3300), .B(n3299), .S(n3195), .Z(n3301) );
  AN3 U2440 ( .A(n3301), .B(n2060), .C(n3213), .Z(n3302) );
  AO1P U2441 ( .A(n3304), .B(n2060), .C(n3303), .D(n3302), .Z(rd_data1[0]) );
  MUX21L U2442 ( .A(\gpr[6][1] ), .B(\gpr[7][1] ), .S(n3180), .Z(n3305) );
  NR2I U2443 ( .A(n3214), .B(n3306), .Z(n3327) );
  MUX21L U2444 ( .A(\gpr[10][1] ), .B(\gpr[11][1] ), .S(n3180), .Z(n3307) );
  MUX21L U2445 ( .A(n134), .B(n65), .S(n2021), .Z(n3308) );
  MUX21L U2446 ( .A(\gpr[22][1] ), .B(\gpr[23][1] ), .S(n2038), .Z(n3309) );
  MUX21L U2447 ( .A(\gpr[26][1] ), .B(\gpr[27][1] ), .S(n2018), .Z(n3310) );
  MUX21L U2448 ( .A(n135), .B(n66), .S(n2034), .Z(n3315) );
  MUX21L U2449 ( .A(n136), .B(n67), .S(n3170), .Z(n3316) );
  AO1P U2450 ( .A(n3145), .B(n3321), .C(n3320), .D(n3319), .Z(n3326) );
  NR2I U2451 ( .A(n3188), .B(n1160), .Z(n3323) );
  MUX21L U2452 ( .A(n1140), .B(n82), .S(n3174), .Z(n3322) );
  MUX21L U2453 ( .A(n3323), .B(n3322), .S(n3195), .Z(n3324) );
  AN3 U2454 ( .A(n3324), .B(n2056), .C(n3214), .Z(n3325) );
  AO1P U2455 ( .A(n3327), .B(n2064), .C(n3326), .D(n3325), .Z(rd_data1[1]) );
  MUX21L U2456 ( .A(\gpr[6][2] ), .B(\gpr[7][2] ), .S(n3169), .Z(n3328) );
  NR2I U2457 ( .A(n3214), .B(n3329), .Z(n3350) );
  MUX21L U2458 ( .A(\gpr[10][2] ), .B(\gpr[11][2] ), .S(n3173), .Z(n3330) );
  MUX21L U2459 ( .A(n137), .B(n68), .S(n2041), .Z(n3331) );
  MUX21L U2460 ( .A(n138), .B(n69), .S(n2034), .Z(n3338) );
  MUX21L U2461 ( .A(n139), .B(n70), .S(n2038), .Z(n3339) );
  AO1P U2462 ( .A(n3145), .B(n3344), .C(n3343), .D(n3342), .Z(n3349) );
  NR2I U2463 ( .A(n2028), .B(n142), .Z(n3346) );
  MUX21L U2464 ( .A(n140), .B(n71), .S(n3176), .Z(n3345) );
  MUX21L U2465 ( .A(n3346), .B(n3345), .S(n3195), .Z(n3347) );
  AN3 U2466 ( .A(n3347), .B(n2062), .C(n3214), .Z(n3348) );
  AO1P U2467 ( .A(n3350), .B(n2060), .C(n3349), .D(n3348), .Z(rd_data1[2]) );
  MUX21L U2468 ( .A(n1161), .B(n95), .S(n3162), .Z(n3352) );
  MUX21L U2469 ( .A(n1251), .B(n1282), .S(n3171), .Z(n3351) );
  MUX21L U2470 ( .A(n3352), .B(n3351), .S(n3195), .Z(n3353) );
  ND2I U2471 ( .A(n3353), .B(n3210), .Z(n3354) );
  NR2I U2472 ( .A(n2055), .B(n3354), .Z(n3389) );
  ND2I U2473 ( .A(\gpr[1][3] ), .B(n2040), .Z(n3356) );
  MUX21L U2474 ( .A(\gpr[2][3] ), .B(\gpr[3][3] ), .S(n2036), .Z(n3355) );
  MUX21L U2475 ( .A(n3356), .B(n3355), .S(n3195), .Z(n3357) );
  NR2I U2476 ( .A(n3357), .B(n3210), .Z(n3358) );
  ND2I U2477 ( .A(n3358), .B(n2064), .Z(n3387) );
  MUX21L U2478 ( .A(\gpr[20][3] ), .B(\gpr[21][3] ), .S(n3175), .Z(n3360) );
  MUX21L U2479 ( .A(\gpr[22][3] ), .B(\gpr[23][3] ), .S(n3178), .Z(n3359) );
  MUX21L U2480 ( .A(n3360), .B(n3359), .S(n2072), .Z(n3361) );
  ND2I U2481 ( .A(n2098), .B(n3361), .Z(n3370) );
  MUX21L U2482 ( .A(\gpr[24][3] ), .B(\gpr[25][3] ), .S(n3180), .Z(n3363) );
  MUX21L U2483 ( .A(\gpr[26][3] ), .B(\gpr[27][3] ), .S(n3169), .Z(n3362) );
  ND2I U2484 ( .A(n2078), .B(n3364), .Z(n3369) );
  MUX21L U2485 ( .A(\gpr[28][3] ), .B(\gpr[29][3] ), .S(n3005), .Z(n3366) );
  MUX21L U2486 ( .A(\gpr[30][3] ), .B(\gpr[31][3] ), .S(n3180), .Z(n3365) );
  MUX21L U2487 ( .A(n3366), .B(n3365), .S(n2072), .Z(n3367) );
  ND2I U2488 ( .A(n3138), .B(n3367), .Z(n3368) );
  MUX21L U2489 ( .A(\gpr[12][3] ), .B(\gpr[13][3] ), .S(n3167), .Z(n3372) );
  MUX21L U2490 ( .A(\gpr[14][3] ), .B(\gpr[15][3] ), .S(n3005), .Z(n3371) );
  MUX21L U2491 ( .A(n3372), .B(n3371), .S(n2049), .Z(n3373) );
  ND2I U2492 ( .A(n3139), .B(n3373), .Z(n3378) );
  MUX21L U2493 ( .A(\gpr[16][3] ), .B(\gpr[17][3] ), .S(n3171), .Z(n3375) );
  MUX21L U2494 ( .A(\gpr[18][3] ), .B(\gpr[19][3] ), .S(n3180), .Z(n3374) );
  MUX21L U2495 ( .A(n3375), .B(n3374), .S(n2049), .Z(n3376) );
  ND2I U2496 ( .A(n3142), .B(n3376), .Z(n3377) );
  ND2I U2497 ( .A(n3378), .B(n3377), .Z(n3379) );
  NR2I U2498 ( .A(n3380), .B(n3379), .Z(n3385) );
  MUX21L U2499 ( .A(\gpr[8][3] ), .B(\gpr[9][3] ), .S(n3167), .Z(n3382) );
  MUX21L U2500 ( .A(\gpr[10][3] ), .B(\gpr[11][3] ), .S(n2071), .Z(n3381) );
  MUX21L U2501 ( .A(n3382), .B(n3381), .S(n2050), .Z(n3383) );
  ND2I U2502 ( .A(n3145), .B(n3383), .Z(n3384) );
  ND2I U2503 ( .A(n3385), .B(n3384), .Z(n3386) );
  ND2I U2504 ( .A(n3387), .B(n3386), .Z(n3388) );
  NR2I U2505 ( .A(n3389), .B(n3388), .Z(rd_data1[3]) );
  MUX21L U2506 ( .A(n141), .B(n72), .S(n3169), .Z(n3391) );
  MUX21L U2507 ( .A(n1252), .B(n1283), .S(n2048), .Z(n3390) );
  MUX21L U2508 ( .A(n3391), .B(n3390), .S(n2049), .Z(n3392) );
  ND2I U2509 ( .A(\gpr[1][4] ), .B(n3180), .Z(n3394) );
  MUX21L U2510 ( .A(\gpr[2][4] ), .B(\gpr[3][4] ), .S(n3169), .Z(n3393) );
  NR2I U2511 ( .A(n3395), .B(n3211), .Z(n3396) );
  ND2I U2512 ( .A(n3396), .B(n2056), .Z(n3422) );
  MUX21L U2513 ( .A(\gpr[20][4] ), .B(\gpr[21][4] ), .S(n3170), .Z(n3398) );
  MUX21L U2514 ( .A(\gpr[22][4] ), .B(\gpr[23][4] ), .S(n2035), .Z(n3397) );
  ND2I U2515 ( .A(n2096), .B(n3399), .Z(n3408) );
  MUX21L U2516 ( .A(\gpr[24][4] ), .B(\gpr[25][4] ), .S(n2035), .Z(n3401) );
  MUX21L U2517 ( .A(\gpr[26][4] ), .B(\gpr[27][4] ), .S(n2035), .Z(n3400) );
  MUX21L U2518 ( .A(n3401), .B(n3400), .S(n3194), .Z(n3402) );
  ND2I U2519 ( .A(n2076), .B(n3402), .Z(n3407) );
  MUX21L U2520 ( .A(\gpr[28][4] ), .B(\gpr[29][4] ), .S(n3170), .Z(n3404) );
  MUX21L U2521 ( .A(\gpr[30][4] ), .B(\gpr[31][4] ), .S(n3170), .Z(n3403) );
  MUX21L U2522 ( .A(n3404), .B(n3403), .S(n2072), .Z(n3405) );
  ND2I U2523 ( .A(n3136), .B(n3405), .Z(n3406) );
  MUX21L U2524 ( .A(\gpr[12][4] ), .B(\gpr[13][4] ), .S(n3177), .Z(n3410) );
  MUX21L U2525 ( .A(\gpr[14][4] ), .B(\gpr[15][4] ), .S(n3177), .Z(n3409) );
  MUX21L U2526 ( .A(n3410), .B(n3409), .S(n2072), .Z(n3411) );
  ND2I U2527 ( .A(n3139), .B(n3411), .Z(n3416) );
  MUX21L U2528 ( .A(\gpr[16][4] ), .B(\gpr[17][4] ), .S(n3176), .Z(n3413) );
  MUX21L U2529 ( .A(\gpr[18][4] ), .B(\gpr[19][4] ), .S(n3177), .Z(n3412) );
  MUX21L U2530 ( .A(n3413), .B(n3412), .S(n2072), .Z(n3414) );
  ND2I U2531 ( .A(n3142), .B(n3414), .Z(n3415) );
  ND2I U2532 ( .A(n3416), .B(n3415), .Z(n3417) );
  MUX21L U2533 ( .A(\gpr[8][4] ), .B(\gpr[9][4] ), .S(n3176), .Z(n3419) );
  MUX21L U2534 ( .A(\gpr[10][4] ), .B(\gpr[11][4] ), .S(n3177), .Z(n3418) );
  MUX21L U2535 ( .A(n3419), .B(n3418), .S(n2049), .Z(n3420) );
  ND2I U2536 ( .A(n3145), .B(n3420), .Z(n3421) );
  MUX21L U2537 ( .A(n1141), .B(n83), .S(n3177), .Z(n3424) );
  MUX21L U2538 ( .A(n1253), .B(n1284), .S(n3176), .Z(n3423) );
  MUX21L U2539 ( .A(n3424), .B(n3423), .S(n2050), .Z(n3425) );
  ND2I U2540 ( .A(n3425), .B(n3208), .Z(n3426) );
  NR2I U2541 ( .A(n2061), .B(n3426), .Z(n3461) );
  ND2I U2542 ( .A(\gpr[1][5] ), .B(n3168), .Z(n3428) );
  MUX21L U2543 ( .A(\gpr[2][5] ), .B(\gpr[3][5] ), .S(n3005), .Z(n3427) );
  MUX21L U2544 ( .A(n3428), .B(n3427), .S(n2049), .Z(n3429) );
  NR2I U2545 ( .A(n3429), .B(n3208), .Z(n3430) );
  ND2I U2546 ( .A(n3430), .B(n2060), .Z(n3459) );
  MUX21L U2547 ( .A(\gpr[20][5] ), .B(\gpr[21][5] ), .S(n3169), .Z(n3432) );
  MUX21L U2548 ( .A(\gpr[22][5] ), .B(\gpr[23][5] ), .S(n2048), .Z(n3431) );
  ND2I U2549 ( .A(n2095), .B(n3433), .Z(n3442) );
  MUX21L U2550 ( .A(\gpr[24][5] ), .B(\gpr[25][5] ), .S(n3169), .Z(n3435) );
  MUX21L U2551 ( .A(\gpr[26][5] ), .B(\gpr[27][5] ), .S(n3181), .Z(n3434) );
  ND2I U2552 ( .A(n2080), .B(n3436), .Z(n3441) );
  MUX21L U2553 ( .A(\gpr[28][5] ), .B(\gpr[29][5] ), .S(n3169), .Z(n3438) );
  MUX21L U2554 ( .A(\gpr[30][5] ), .B(\gpr[31][5] ), .S(n2048), .Z(n3437) );
  ND2I U2555 ( .A(n3137), .B(n3439), .Z(n3440) );
  MUX21L U2556 ( .A(\gpr[12][5] ), .B(\gpr[13][5] ), .S(n3167), .Z(n3444) );
  MUX21L U2557 ( .A(\gpr[14][5] ), .B(\gpr[15][5] ), .S(n3179), .Z(n3443) );
  MUX21L U2558 ( .A(n3444), .B(n3443), .S(n3193), .Z(n3445) );
  ND2I U2559 ( .A(n3139), .B(n3445), .Z(n3450) );
  MUX21L U2560 ( .A(\gpr[16][5] ), .B(\gpr[17][5] ), .S(n3167), .Z(n3447) );
  MUX21L U2561 ( .A(\gpr[18][5] ), .B(\gpr[19][5] ), .S(n2071), .Z(n3446) );
  MUX21L U2562 ( .A(n3447), .B(n3446), .S(n3193), .Z(n3448) );
  ND2I U2563 ( .A(n3142), .B(n3448), .Z(n3449) );
  ND2I U2564 ( .A(n3450), .B(n3449), .Z(n3451) );
  NR2I U2565 ( .A(n3452), .B(n3451), .Z(n3457) );
  MUX21L U2566 ( .A(\gpr[8][5] ), .B(\gpr[9][5] ), .S(n3167), .Z(n3454) );
  MUX21L U2567 ( .A(\gpr[10][5] ), .B(\gpr[11][5] ), .S(n3179), .Z(n3453) );
  MUX21L U2568 ( .A(n3454), .B(n3453), .S(n3193), .Z(n3455) );
  ND2I U2569 ( .A(n3145), .B(n3455), .Z(n3456) );
  ND2I U2570 ( .A(n3457), .B(n3456), .Z(n3458) );
  ND2I U2571 ( .A(n3459), .B(n3458), .Z(n3460) );
  NR2I U2572 ( .A(n3461), .B(n3460), .Z(rd_data1[5]) );
  MUX21L U2573 ( .A(n1162), .B(n96), .S(n2071), .Z(n3463) );
  MUX21L U2574 ( .A(n1254), .B(n1285), .S(n3171), .Z(n3462) );
  MUX21L U2575 ( .A(n3463), .B(n3462), .S(n3193), .Z(n3464) );
  ND2I U2576 ( .A(n3464), .B(n3208), .Z(n3465) );
  NR2I U2577 ( .A(n2061), .B(n3465), .Z(n3500) );
  ND2I U2578 ( .A(\gpr[1][6] ), .B(n3178), .Z(n3467) );
  MUX21L U2579 ( .A(\gpr[2][6] ), .B(\gpr[3][6] ), .S(n3167), .Z(n3466) );
  MUX21L U2580 ( .A(n3467), .B(n3466), .S(n3193), .Z(n3468) );
  NR2I U2581 ( .A(n3468), .B(n3208), .Z(n3469) );
  ND2I U2582 ( .A(n3469), .B(n2062), .Z(n3498) );
  MUX21L U2583 ( .A(\gpr[20][6] ), .B(\gpr[21][6] ), .S(n3171), .Z(n3471) );
  MUX21L U2584 ( .A(\gpr[22][6] ), .B(\gpr[23][6] ), .S(n2041), .Z(n3470) );
  MUX21L U2585 ( .A(n3471), .B(n3470), .S(n3193), .Z(n3472) );
  ND2I U2586 ( .A(n2093), .B(n3472), .Z(n3481) );
  MUX21L U2587 ( .A(\gpr[24][6] ), .B(\gpr[25][6] ), .S(n3171), .Z(n3474) );
  MUX21L U2588 ( .A(\gpr[26][6] ), .B(\gpr[27][6] ), .S(n3171), .Z(n3473) );
  MUX21L U2589 ( .A(n3474), .B(n3473), .S(n3193), .Z(n3475) );
  ND2I U2590 ( .A(n2078), .B(n3475), .Z(n3480) );
  MUX21L U2591 ( .A(\gpr[28][6] ), .B(\gpr[29][6] ), .S(n3171), .Z(n3477) );
  MUX21L U2592 ( .A(\gpr[30][6] ), .B(\gpr[31][6] ), .S(n3179), .Z(n3476) );
  MUX21L U2593 ( .A(n3477), .B(n3476), .S(n3193), .Z(n3478) );
  ND2I U2594 ( .A(n3137), .B(n3478), .Z(n3479) );
  MUX21L U2595 ( .A(\gpr[12][6] ), .B(\gpr[13][6] ), .S(n3171), .Z(n3483) );
  MUX21L U2596 ( .A(\gpr[14][6] ), .B(\gpr[15][6] ), .S(n3179), .Z(n3482) );
  MUX21L U2597 ( .A(n3483), .B(n3482), .S(n3193), .Z(n3484) );
  ND2I U2598 ( .A(n3139), .B(n3484), .Z(n3489) );
  MUX21L U2599 ( .A(\gpr[16][6] ), .B(\gpr[17][6] ), .S(n3180), .Z(n3486) );
  MUX21L U2600 ( .A(\gpr[18][6] ), .B(\gpr[19][6] ), .S(n3167), .Z(n3485) );
  MUX21L U2601 ( .A(n3486), .B(n3485), .S(n3193), .Z(n3487) );
  ND2I U2602 ( .A(n3142), .B(n3487), .Z(n3488) );
  ND2I U2603 ( .A(n3489), .B(n3488), .Z(n3490) );
  NR2I U2604 ( .A(n3491), .B(n3490), .Z(n3496) );
  MUX21L U2605 ( .A(\gpr[8][6] ), .B(\gpr[9][6] ), .S(n3168), .Z(n3493) );
  MUX21L U2606 ( .A(\gpr[10][6] ), .B(\gpr[11][6] ), .S(n2071), .Z(n3492) );
  MUX21L U2607 ( .A(n3493), .B(n3492), .S(n3193), .Z(n3494) );
  ND2I U2608 ( .A(n3145), .B(n3494), .Z(n3495) );
  ND2I U2609 ( .A(n3496), .B(n3495), .Z(n3497) );
  ND2I U2610 ( .A(n3498), .B(n3497), .Z(n3499) );
  NR2I U2611 ( .A(n3500), .B(n3499), .Z(rd_data1[6]) );
  MUX21L U2612 ( .A(n1163), .B(n97), .S(n3167), .Z(n3502) );
  MUX21L U2613 ( .A(n1178), .B(n114), .S(n3167), .Z(n3501) );
  MUX21L U2614 ( .A(n3502), .B(n3501), .S(n3193), .Z(n3503) );
  ND2I U2615 ( .A(n3503), .B(n3208), .Z(n3504) );
  NR2I U2616 ( .A(n2065), .B(n3504), .Z(n3539) );
  ND2I U2617 ( .A(\gpr[1][7] ), .B(n3179), .Z(n3506) );
  MUX21L U2618 ( .A(\gpr[2][7] ), .B(\gpr[3][7] ), .S(n3167), .Z(n3505) );
  MUX21L U2619 ( .A(n3506), .B(n3505), .S(n3193), .Z(n3507) );
  NR2I U2620 ( .A(n3507), .B(n3208), .Z(n3508) );
  ND2I U2621 ( .A(n3508), .B(n2066), .Z(n3537) );
  MUX21L U2622 ( .A(\gpr[20][7] ), .B(\gpr[21][7] ), .S(n3167), .Z(n3510) );
  MUX21L U2623 ( .A(\gpr[22][7] ), .B(\gpr[23][7] ), .S(n2041), .Z(n3509) );
  MUX21L U2624 ( .A(n3510), .B(n3509), .S(n3193), .Z(n3511) );
  ND2I U2625 ( .A(n2099), .B(n3511), .Z(n3520) );
  MUX21L U2626 ( .A(\gpr[24][7] ), .B(\gpr[25][7] ), .S(n3005), .Z(n3513) );
  MUX21L U2627 ( .A(\gpr[26][7] ), .B(\gpr[27][7] ), .S(n3180), .Z(n3512) );
  MUX21L U2628 ( .A(n3513), .B(n3512), .S(n3193), .Z(n3514) );
  ND2I U2629 ( .A(n2075), .B(n3514), .Z(n3519) );
  MUX21L U2630 ( .A(\gpr[28][7] ), .B(\gpr[29][7] ), .S(n3169), .Z(n3516) );
  MUX21L U2631 ( .A(\gpr[30][7] ), .B(\gpr[31][7] ), .S(n3169), .Z(n3515) );
  MUX21L U2632 ( .A(n3516), .B(n3515), .S(n3193), .Z(n3517) );
  ND2I U2633 ( .A(n3135), .B(n3517), .Z(n3518) );
  MUX21L U2634 ( .A(\gpr[12][7] ), .B(\gpr[13][7] ), .S(n2071), .Z(n3522) );
  MUX21L U2635 ( .A(\gpr[14][7] ), .B(\gpr[15][7] ), .S(n3167), .Z(n3521) );
  MUX21L U2636 ( .A(n3522), .B(n3521), .S(n3193), .Z(n3523) );
  ND2I U2637 ( .A(n3139), .B(n3523), .Z(n3528) );
  MUX21L U2638 ( .A(\gpr[16][7] ), .B(\gpr[17][7] ), .S(n3171), .Z(n3525) );
  MUX21L U2639 ( .A(\gpr[18][7] ), .B(\gpr[19][7] ), .S(n3180), .Z(n3524) );
  MUX21L U2640 ( .A(n3525), .B(n3524), .S(n3193), .Z(n3526) );
  ND2I U2641 ( .A(n3142), .B(n3526), .Z(n3527) );
  ND2I U2642 ( .A(n3528), .B(n3527), .Z(n3529) );
  NR2I U2643 ( .A(n3530), .B(n3529), .Z(n3535) );
  MUX21L U2644 ( .A(\gpr[8][7] ), .B(\gpr[9][7] ), .S(n3167), .Z(n3532) );
  MUX21L U2645 ( .A(\gpr[10][7] ), .B(\gpr[11][7] ), .S(n3178), .Z(n3531) );
  MUX21L U2646 ( .A(n3532), .B(n3531), .S(n3193), .Z(n3533) );
  ND2I U2647 ( .A(n3145), .B(n3533), .Z(n3534) );
  ND2I U2648 ( .A(n3535), .B(n3534), .Z(n3536) );
  ND2I U2649 ( .A(n3537), .B(n3536), .Z(n3538) );
  NR2I U2650 ( .A(n3539), .B(n3538), .Z(rd_data1[7]) );
  MUX21L U2651 ( .A(n1142), .B(n98), .S(n3178), .Z(n3541) );
  MUX21L U2652 ( .A(n1255), .B(n1286), .S(n3166), .Z(n3540) );
  MUX21L U2653 ( .A(n3541), .B(n3540), .S(n3195), .Z(n3542) );
  ND2I U2654 ( .A(n3542), .B(n3208), .Z(n3543) );
  NR2I U2655 ( .A(n2061), .B(n3543), .Z(n3578) );
  ND2I U2656 ( .A(\gpr[1][8] ), .B(n2040), .Z(n3545) );
  MUX21L U2657 ( .A(\gpr[2][8] ), .B(\gpr[3][8] ), .S(n3178), .Z(n3544) );
  MUX21L U2658 ( .A(n3545), .B(n3544), .S(n3192), .Z(n3546) );
  NR2I U2659 ( .A(n3546), .B(n3208), .Z(n3547) );
  ND2I U2660 ( .A(n3547), .B(n2060), .Z(n3576) );
  MUX21L U2661 ( .A(\gpr[20][8] ), .B(\gpr[21][8] ), .S(n2101), .Z(n3549) );
  MUX21L U2662 ( .A(\gpr[22][8] ), .B(\gpr[23][8] ), .S(n2048), .Z(n3548) );
  MUX21L U2663 ( .A(n3549), .B(n3548), .S(n3192), .Z(n3550) );
  ND2I U2664 ( .A(n2094), .B(n3550), .Z(n3559) );
  MUX21L U2665 ( .A(\gpr[24][8] ), .B(\gpr[25][8] ), .S(n2021), .Z(n3552) );
  MUX21L U2666 ( .A(\gpr[26][8] ), .B(\gpr[27][8] ), .S(n2036), .Z(n3551) );
  ND2I U2667 ( .A(n2077), .B(n3553), .Z(n3558) );
  MUX21L U2668 ( .A(\gpr[28][8] ), .B(\gpr[29][8] ), .S(n3168), .Z(n3555) );
  MUX21L U2669 ( .A(\gpr[30][8] ), .B(\gpr[31][8] ), .S(n3181), .Z(n3554) );
  MUX21L U2670 ( .A(n3555), .B(n3554), .S(n3192), .Z(n3556) );
  ND2I U2671 ( .A(n3135), .B(n3556), .Z(n3557) );
  MUX21L U2672 ( .A(\gpr[12][8] ), .B(\gpr[13][8] ), .S(n3156), .Z(n3561) );
  MUX21L U2673 ( .A(\gpr[14][8] ), .B(\gpr[15][8] ), .S(n3159), .Z(n3560) );
  MUX21L U2674 ( .A(n3561), .B(n3560), .S(n3192), .Z(n3562) );
  ND2I U2675 ( .A(n3139), .B(n3562), .Z(n3567) );
  MUX21L U2676 ( .A(\gpr[16][8] ), .B(\gpr[17][8] ), .S(n3180), .Z(n3564) );
  MUX21L U2677 ( .A(\gpr[18][8] ), .B(\gpr[19][8] ), .S(n3180), .Z(n3563) );
  MUX21L U2678 ( .A(n3564), .B(n3563), .S(n3192), .Z(n3565) );
  ND2I U2679 ( .A(n3142), .B(n3565), .Z(n3566) );
  ND2I U2680 ( .A(n3567), .B(n3566), .Z(n3568) );
  NR2I U2681 ( .A(n3569), .B(n3568), .Z(n3574) );
  MUX21L U2682 ( .A(\gpr[8][8] ), .B(\gpr[9][8] ), .S(n3180), .Z(n3571) );
  MUX21L U2683 ( .A(\gpr[10][8] ), .B(\gpr[11][8] ), .S(n3178), .Z(n3570) );
  MUX21L U2684 ( .A(n3571), .B(n3570), .S(n3192), .Z(n3572) );
  ND2I U2685 ( .A(n3145), .B(n3572), .Z(n3573) );
  ND2I U2686 ( .A(n3574), .B(n3573), .Z(n3575) );
  ND2I U2687 ( .A(n3576), .B(n3575), .Z(n3577) );
  NR2I U2688 ( .A(n3578), .B(n3577), .Z(rd_data1[8]) );
  MUX21L U2689 ( .A(n1143), .B(n84), .S(n3180), .Z(n3580) );
  MUX21L U2690 ( .A(n1256), .B(n1287), .S(n3168), .Z(n3579) );
  MUX21L U2691 ( .A(n3580), .B(n3579), .S(n3192), .Z(n3581) );
  ND2I U2692 ( .A(n3581), .B(n3208), .Z(n3582) );
  NR2I U2693 ( .A(n2065), .B(n3582), .Z(n3617) );
  ND2I U2694 ( .A(\gpr[1][9] ), .B(n3178), .Z(n3584) );
  MUX21L U2695 ( .A(\gpr[2][9] ), .B(\gpr[3][9] ), .S(n3168), .Z(n3583) );
  MUX21L U2696 ( .A(n3584), .B(n3583), .S(n3192), .Z(n3585) );
  NR2I U2697 ( .A(n3585), .B(n3208), .Z(n3586) );
  ND2I U2698 ( .A(n3586), .B(n2062), .Z(n3615) );
  MUX21L U2699 ( .A(\gpr[20][9] ), .B(\gpr[21][9] ), .S(n3179), .Z(n3588) );
  MUX21L U2700 ( .A(\gpr[22][9] ), .B(\gpr[23][9] ), .S(n3179), .Z(n3587) );
  ND2I U2701 ( .A(n2097), .B(n3589), .Z(n3598) );
  MUX21L U2702 ( .A(\gpr[24][9] ), .B(\gpr[25][9] ), .S(n3179), .Z(n3591) );
  MUX21L U2703 ( .A(\gpr[26][9] ), .B(\gpr[27][9] ), .S(n3179), .Z(n3590) );
  ND2I U2704 ( .A(n2077), .B(n3592), .Z(n3597) );
  MUX21L U2705 ( .A(\gpr[28][9] ), .B(\gpr[29][9] ), .S(n3179), .Z(n3594) );
  MUX21L U2706 ( .A(\gpr[30][9] ), .B(\gpr[31][9] ), .S(n2034), .Z(n3593) );
  ND2I U2707 ( .A(n3136), .B(n3595), .Z(n3596) );
  MUX21L U2708 ( .A(\gpr[12][9] ), .B(\gpr[13][9] ), .S(n2021), .Z(n3600) );
  MUX21L U2709 ( .A(\gpr[14][9] ), .B(\gpr[15][9] ), .S(n3158), .Z(n3599) );
  MUX21L U2710 ( .A(n3600), .B(n3599), .S(n3192), .Z(n3601) );
  ND2I U2711 ( .A(n3139), .B(n3601), .Z(n3606) );
  MUX21L U2712 ( .A(\gpr[16][9] ), .B(\gpr[17][9] ), .S(n3181), .Z(n3603) );
  MUX21L U2713 ( .A(\gpr[18][9] ), .B(\gpr[19][9] ), .S(n3181), .Z(n3602) );
  MUX21L U2714 ( .A(n3603), .B(n3602), .S(n3192), .Z(n3604) );
  ND2I U2715 ( .A(n3142), .B(n3604), .Z(n3605) );
  ND2I U2716 ( .A(n3606), .B(n3605), .Z(n3607) );
  NR2I U2717 ( .A(n3608), .B(n3607), .Z(n3613) );
  MUX21L U2718 ( .A(\gpr[8][9] ), .B(\gpr[9][9] ), .S(n3176), .Z(n3610) );
  MUX21L U2719 ( .A(\gpr[10][9] ), .B(\gpr[11][9] ), .S(n3168), .Z(n3609) );
  MUX21L U2720 ( .A(n3610), .B(n3609), .S(n3192), .Z(n3611) );
  ND2I U2721 ( .A(n3145), .B(n3611), .Z(n3612) );
  ND2I U2722 ( .A(n3613), .B(n3612), .Z(n3614) );
  ND2I U2723 ( .A(n3615), .B(n3614), .Z(n3616) );
  NR2I U2724 ( .A(n3617), .B(n3616), .Z(rd_data1[9]) );
  MUX21L U2725 ( .A(n1144), .B(n99), .S(n3178), .Z(n3619) );
  MUX21L U2726 ( .A(n1257), .B(n1288), .S(n3178), .Z(n3618) );
  MUX21L U2727 ( .A(n3619), .B(n3618), .S(n2072), .Z(n3620) );
  ND2I U2728 ( .A(n3620), .B(n3208), .Z(n3621) );
  NR2I U2729 ( .A(n2063), .B(n3621), .Z(n3656) );
  ND2I U2730 ( .A(\gpr[1][10] ), .B(n3168), .Z(n3623) );
  MUX21L U2731 ( .A(\gpr[2][10] ), .B(\gpr[3][10] ), .S(n3178), .Z(n3622) );
  MUX21L U2732 ( .A(n3623), .B(n3622), .S(n3192), .Z(n3624) );
  NR2I U2733 ( .A(n3624), .B(n3209), .Z(n3625) );
  ND2I U2734 ( .A(n3625), .B(n2066), .Z(n3654) );
  MUX21L U2735 ( .A(\gpr[20][10] ), .B(\gpr[21][10] ), .S(n3179), .Z(n3627) );
  MUX21L U2736 ( .A(\gpr[22][10] ), .B(\gpr[23][10] ), .S(n3179), .Z(n3626) );
  MUX21L U2737 ( .A(n3627), .B(n3626), .S(n3192), .Z(n3628) );
  ND2I U2738 ( .A(n2098), .B(n3628), .Z(n3637) );
  MUX21L U2739 ( .A(\gpr[24][10] ), .B(\gpr[25][10] ), .S(n3170), .Z(n3630) );
  MUX21L U2740 ( .A(\gpr[26][10] ), .B(\gpr[27][10] ), .S(n3179), .Z(n3629) );
  MUX21L U2741 ( .A(n3630), .B(n3629), .S(n3191), .Z(n3631) );
  ND2I U2742 ( .A(n2076), .B(n3631), .Z(n3636) );
  MUX21L U2743 ( .A(\gpr[28][10] ), .B(\gpr[29][10] ), .S(n3179), .Z(n3633) );
  MUX21L U2744 ( .A(\gpr[30][10] ), .B(\gpr[31][10] ), .S(n3179), .Z(n3632) );
  MUX21L U2745 ( .A(n3633), .B(n3632), .S(n3191), .Z(n3634) );
  ND2I U2746 ( .A(n3136), .B(n3634), .Z(n3635) );
  MUX21L U2747 ( .A(\gpr[12][10] ), .B(\gpr[13][10] ), .S(n3180), .Z(n3639) );
  MUX21L U2748 ( .A(\gpr[14][10] ), .B(\gpr[15][10] ), .S(n3177), .Z(n3638) );
  MUX21L U2749 ( .A(n3639), .B(n3638), .S(n3191), .Z(n3640) );
  ND2I U2750 ( .A(n3139), .B(n3640), .Z(n3645) );
  MUX21L U2751 ( .A(\gpr[16][10] ), .B(\gpr[17][10] ), .S(n3157), .Z(n3642) );
  MUX21L U2752 ( .A(\gpr[18][10] ), .B(\gpr[19][10] ), .S(n3176), .Z(n3641) );
  MUX21L U2753 ( .A(n3642), .B(n3641), .S(n3191), .Z(n3643) );
  ND2I U2754 ( .A(n3142), .B(n3643), .Z(n3644) );
  ND2I U2755 ( .A(n3645), .B(n3644), .Z(n3646) );
  NR2I U2756 ( .A(n3647), .B(n3646), .Z(n3652) );
  MUX21L U2757 ( .A(\gpr[8][10] ), .B(\gpr[9][10] ), .S(n3177), .Z(n3649) );
  MUX21L U2758 ( .A(\gpr[10][10] ), .B(\gpr[11][10] ), .S(n3177), .Z(n3648) );
  MUX21L U2759 ( .A(n3649), .B(n3648), .S(n3191), .Z(n3650) );
  ND2I U2760 ( .A(n3145), .B(n3650), .Z(n3651) );
  ND2I U2761 ( .A(n3652), .B(n3651), .Z(n3653) );
  ND2I U2762 ( .A(n3654), .B(n3653), .Z(n3655) );
  NR2I U2763 ( .A(n3656), .B(n3655), .Z(rd_data1[10]) );
  MUX21L U2764 ( .A(n1164), .B(n100), .S(n3176), .Z(n3658) );
  MUX21L U2765 ( .A(n1258), .B(n1289), .S(n3177), .Z(n3657) );
  MUX21L U2766 ( .A(n3658), .B(n3657), .S(n3191), .Z(n3659) );
  ND2I U2767 ( .A(n3659), .B(n3209), .Z(n3660) );
  NR2I U2768 ( .A(n2063), .B(n3660), .Z(n3695) );
  ND2I U2769 ( .A(\gpr[1][11] ), .B(n3180), .Z(n3662) );
  MUX21L U2770 ( .A(\gpr[2][11] ), .B(\gpr[3][11] ), .S(n3177), .Z(n3661) );
  MUX21L U2771 ( .A(n3662), .B(n3661), .S(n3191), .Z(n3663) );
  NR2I U2772 ( .A(n3663), .B(n3209), .Z(n3664) );
  ND2I U2773 ( .A(n3664), .B(n2066), .Z(n3693) );
  MUX21L U2774 ( .A(\gpr[20][11] ), .B(\gpr[21][11] ), .S(n3177), .Z(n3666) );
  MUX21L U2775 ( .A(\gpr[22][11] ), .B(\gpr[23][11] ), .S(n2021), .Z(n3665) );
  MUX21L U2776 ( .A(n3666), .B(n3665), .S(n3191), .Z(n3667) );
  ND2I U2777 ( .A(n2095), .B(n3667), .Z(n3676) );
  MUX21L U2778 ( .A(\gpr[24][11] ), .B(\gpr[25][11] ), .S(n3176), .Z(n3669) );
  MUX21L U2779 ( .A(\gpr[26][11] ), .B(\gpr[27][11] ), .S(n3177), .Z(n3668) );
  MUX21L U2780 ( .A(n3669), .B(n3668), .S(n3191), .Z(n3670) );
  ND2I U2781 ( .A(n2077), .B(n3670), .Z(n3675) );
  MUX21L U2782 ( .A(\gpr[28][11] ), .B(\gpr[29][11] ), .S(n3177), .Z(n3672) );
  MUX21L U2783 ( .A(\gpr[30][11] ), .B(\gpr[31][11] ), .S(n3176), .Z(n3671) );
  MUX21L U2784 ( .A(n3672), .B(n3671), .S(n3191), .Z(n3673) );
  ND2I U2785 ( .A(n3135), .B(n3673), .Z(n3674) );
  MUX21L U2786 ( .A(\gpr[12][11] ), .B(\gpr[13][11] ), .S(n3177), .Z(n3678) );
  MUX21L U2787 ( .A(\gpr[14][11] ), .B(\gpr[15][11] ), .S(n3176), .Z(n3677) );
  MUX21L U2788 ( .A(n3678), .B(n3677), .S(n3191), .Z(n3679) );
  ND2I U2789 ( .A(n3139), .B(n3679), .Z(n3684) );
  MUX21L U2790 ( .A(\gpr[16][11] ), .B(\gpr[17][11] ), .S(n3177), .Z(n3681) );
  MUX21L U2791 ( .A(\gpr[18][11] ), .B(\gpr[19][11] ), .S(n3177), .Z(n3680) );
  MUX21L U2792 ( .A(n3681), .B(n3680), .S(n3191), .Z(n3682) );
  ND2I U2793 ( .A(n3142), .B(n3682), .Z(n3683) );
  ND2I U2794 ( .A(n3684), .B(n3683), .Z(n3685) );
  NR2I U2795 ( .A(n3686), .B(n3685), .Z(n3691) );
  MUX21L U2796 ( .A(\gpr[8][11] ), .B(\gpr[9][11] ), .S(n3177), .Z(n3688) );
  MUX21L U2797 ( .A(\gpr[10][11] ), .B(\gpr[11][11] ), .S(n3177), .Z(n3687) );
  MUX21L U2798 ( .A(n3688), .B(n3687), .S(n3191), .Z(n3689) );
  ND2I U2799 ( .A(n3145), .B(n3689), .Z(n3690) );
  ND2I U2800 ( .A(n3691), .B(n3690), .Z(n3692) );
  ND2I U2801 ( .A(n3693), .B(n3692), .Z(n3694) );
  NR2I U2802 ( .A(n3695), .B(n3694), .Z(rd_data1[11]) );
  MUX21L U2803 ( .A(n1165), .B(n101), .S(n3177), .Z(n3697) );
  MUX21L U2804 ( .A(n1259), .B(n1290), .S(n3176), .Z(n3696) );
  MUX21L U2805 ( .A(n3697), .B(n3696), .S(n3191), .Z(n3698) );
  ND2I U2806 ( .A(n3698), .B(n3209), .Z(n3699) );
  NR2I U2807 ( .A(n2055), .B(n3699), .Z(n3734) );
  ND2I U2808 ( .A(\gpr[1][12] ), .B(n3178), .Z(n3701) );
  MUX21L U2809 ( .A(\gpr[2][12] ), .B(\gpr[3][12] ), .S(n3176), .Z(n3700) );
  MUX21L U2810 ( .A(n3701), .B(n3700), .S(n3191), .Z(n3702) );
  NR2I U2811 ( .A(n3702), .B(n3209), .Z(n3703) );
  ND2I U2812 ( .A(n3703), .B(n2066), .Z(n3732) );
  MUX21L U2813 ( .A(\gpr[20][12] ), .B(\gpr[21][12] ), .S(n3177), .Z(n3705) );
  MUX21L U2814 ( .A(\gpr[22][12] ), .B(\gpr[23][12] ), .S(n3175), .Z(n3704) );
  MUX21L U2815 ( .A(n3705), .B(n3704), .S(n3191), .Z(n3706) );
  ND2I U2816 ( .A(n2095), .B(n3706), .Z(n3715) );
  MUX21L U2817 ( .A(\gpr[24][12] ), .B(\gpr[25][12] ), .S(n3175), .Z(n3708) );
  MUX21L U2818 ( .A(\gpr[26][12] ), .B(\gpr[27][12] ), .S(n3175), .Z(n3707) );
  MUX21L U2819 ( .A(n3708), .B(n3707), .S(n3191), .Z(n3709) );
  ND2I U2820 ( .A(n2022), .B(n3709), .Z(n3714) );
  MUX21L U2821 ( .A(\gpr[28][12] ), .B(\gpr[29][12] ), .S(n3175), .Z(n3711) );
  MUX21L U2822 ( .A(\gpr[30][12] ), .B(\gpr[31][12] ), .S(n3175), .Z(n3710) );
  MUX21L U2823 ( .A(n3711), .B(n3710), .S(n3191), .Z(n3712) );
  ND2I U2824 ( .A(n3138), .B(n3712), .Z(n3713) );
  MUX21L U2825 ( .A(\gpr[12][12] ), .B(\gpr[13][12] ), .S(n3175), .Z(n3717) );
  MUX21L U2826 ( .A(\gpr[14][12] ), .B(\gpr[15][12] ), .S(n3175), .Z(n3716) );
  MUX21L U2827 ( .A(n3717), .B(n3716), .S(n3191), .Z(n3718) );
  ND2I U2828 ( .A(n3140), .B(n3718), .Z(n3723) );
  MUX21L U2829 ( .A(\gpr[16][12] ), .B(\gpr[17][12] ), .S(n3175), .Z(n3720) );
  MUX21L U2830 ( .A(\gpr[18][12] ), .B(\gpr[19][12] ), .S(n3175), .Z(n3719) );
  MUX21L U2831 ( .A(n3720), .B(n3719), .S(n3193), .Z(n3721) );
  ND2I U2832 ( .A(n3143), .B(n3721), .Z(n3722) );
  ND2I U2833 ( .A(n3723), .B(n3722), .Z(n3724) );
  NR2I U2834 ( .A(n3725), .B(n3724), .Z(n3730) );
  MUX21L U2835 ( .A(\gpr[8][12] ), .B(\gpr[9][12] ), .S(n2036), .Z(n3727) );
  MUX21L U2836 ( .A(\gpr[10][12] ), .B(\gpr[11][12] ), .S(n2036), .Z(n3726) );
  MUX21L U2837 ( .A(n3727), .B(n3726), .S(n2), .Z(n3728) );
  ND2I U2838 ( .A(n3145), .B(n3728), .Z(n3729) );
  ND2I U2839 ( .A(n3730), .B(n3729), .Z(n3731) );
  ND2I U2840 ( .A(n3732), .B(n3731), .Z(n3733) );
  NR2I U2841 ( .A(n3734), .B(n3733), .Z(rd_data1[12]) );
  MUX21L U2842 ( .A(n1145), .B(n85), .S(n2036), .Z(n3736) );
  MUX21L U2843 ( .A(n1260), .B(n1291), .S(n2036), .Z(n3735) );
  MUX21L U2844 ( .A(n3736), .B(n3735), .S(n2050), .Z(n3737) );
  ND2I U2845 ( .A(n3737), .B(n3209), .Z(n3738) );
  NR2I U2846 ( .A(n2063), .B(n3738), .Z(n3773) );
  ND2I U2847 ( .A(\gpr[1][13] ), .B(n3180), .Z(n3740) );
  MUX21L U2848 ( .A(\gpr[2][13] ), .B(\gpr[3][13] ), .S(n3175), .Z(n3739) );
  MUX21L U2849 ( .A(n3740), .B(n3739), .S(n3193), .Z(n3741) );
  NR2I U2850 ( .A(n3741), .B(n3209), .Z(n3742) );
  ND2I U2851 ( .A(n3742), .B(n2062), .Z(n3771) );
  MUX21L U2852 ( .A(\gpr[20][13] ), .B(\gpr[21][13] ), .S(n3179), .Z(n3744) );
  MUX21L U2853 ( .A(\gpr[22][13] ), .B(\gpr[23][13] ), .S(n2088), .Z(n3743) );
  MUX21L U2854 ( .A(n3744), .B(n3743), .S(n2083), .Z(n3745) );
  ND2I U2855 ( .A(n2093), .B(n3745), .Z(n3754) );
  MUX21L U2856 ( .A(\gpr[24][13] ), .B(\gpr[25][13] ), .S(n3179), .Z(n3747) );
  MUX21L U2857 ( .A(\gpr[26][13] ), .B(\gpr[27][13] ), .S(n2088), .Z(n3746) );
  MUX21L U2858 ( .A(n3747), .B(n3746), .S(n2083), .Z(n3748) );
  ND2I U2859 ( .A(n2075), .B(n3748), .Z(n3753) );
  MUX21L U2860 ( .A(\gpr[28][13] ), .B(\gpr[29][13] ), .S(n2088), .Z(n3750) );
  MUX21L U2861 ( .A(\gpr[30][13] ), .B(\gpr[31][13] ), .S(n2088), .Z(n3749) );
  MUX21L U2862 ( .A(n3750), .B(n3749), .S(n2083), .Z(n3751) );
  ND2I U2863 ( .A(n3135), .B(n3751), .Z(n3752) );
  MUX21L U2864 ( .A(\gpr[12][13] ), .B(\gpr[13][13] ), .S(n2036), .Z(n3756) );
  MUX21L U2865 ( .A(\gpr[14][13] ), .B(\gpr[15][13] ), .S(n3174), .Z(n3755) );
  MUX21L U2866 ( .A(n3756), .B(n3755), .S(n2050), .Z(n3757) );
  ND2I U2867 ( .A(n3140), .B(n3757), .Z(n3762) );
  MUX21L U2868 ( .A(\gpr[16][13] ), .B(\gpr[17][13] ), .S(n3174), .Z(n3759) );
  MUX21L U2869 ( .A(\gpr[18][13] ), .B(\gpr[19][13] ), .S(n3174), .Z(n3758) );
  MUX21L U2870 ( .A(n3759), .B(n3758), .S(n3196), .Z(n3760) );
  ND2I U2871 ( .A(n3143), .B(n3760), .Z(n3761) );
  ND2I U2872 ( .A(n3762), .B(n3761), .Z(n3763) );
  NR2I U2873 ( .A(n3764), .B(n3763), .Z(n3769) );
  MUX21L U2874 ( .A(\gpr[8][13] ), .B(\gpr[9][13] ), .S(n3174), .Z(n3766) );
  MUX21L U2875 ( .A(\gpr[10][13] ), .B(\gpr[11][13] ), .S(n3174), .Z(n3765) );
  MUX21L U2876 ( .A(n3766), .B(n3765), .S(n3196), .Z(n3767) );
  ND2I U2877 ( .A(n3145), .B(n3767), .Z(n3768) );
  ND2I U2878 ( .A(n3769), .B(n3768), .Z(n3770) );
  ND2I U2879 ( .A(n3771), .B(n3770), .Z(n3772) );
  NR2I U2880 ( .A(n3773), .B(n3772), .Z(rd_data1[13]) );
  MUX21L U2881 ( .A(n1146), .B(n86), .S(n3174), .Z(n3775) );
  MUX21L U2882 ( .A(n1261), .B(n1292), .S(n3174), .Z(n3774) );
  MUX21L U2883 ( .A(n3775), .B(n3774), .S(n3196), .Z(n3776) );
  ND2I U2884 ( .A(n3776), .B(n3209), .Z(n3777) );
  ND2I U2885 ( .A(\gpr[1][14] ), .B(n3180), .Z(n3779) );
  MUX21L U2886 ( .A(\gpr[2][14] ), .B(\gpr[3][14] ), .S(n3173), .Z(n3778) );
  MUX21L U2887 ( .A(n3779), .B(n3778), .S(n3192), .Z(n3780) );
  NR2I U2888 ( .A(n3780), .B(n3209), .Z(n3781) );
  ND2I U2889 ( .A(n3781), .B(n2058), .Z(n3810) );
  MUX21L U2890 ( .A(\gpr[20][14] ), .B(\gpr[21][14] ), .S(n3173), .Z(n3783) );
  MUX21L U2891 ( .A(\gpr[22][14] ), .B(\gpr[23][14] ), .S(n3173), .Z(n3782) );
  MUX21L U2892 ( .A(n3783), .B(n3782), .S(n2050), .Z(n3784) );
  ND2I U2893 ( .A(n2099), .B(n3784), .Z(n3793) );
  MUX21L U2894 ( .A(\gpr[24][14] ), .B(\gpr[25][14] ), .S(n3173), .Z(n3786) );
  MUX21L U2895 ( .A(\gpr[26][14] ), .B(\gpr[27][14] ), .S(n3173), .Z(n3785) );
  MUX21L U2896 ( .A(n3786), .B(n3785), .S(n2050), .Z(n3787) );
  ND2I U2897 ( .A(n2074), .B(n3787), .Z(n3792) );
  MUX21L U2898 ( .A(\gpr[28][14] ), .B(\gpr[29][14] ), .S(n3173), .Z(n3789) );
  MUX21L U2899 ( .A(\gpr[30][14] ), .B(\gpr[31][14] ), .S(n3173), .Z(n3788) );
  MUX21L U2900 ( .A(n3789), .B(n3788), .S(n2050), .Z(n3790) );
  ND2I U2901 ( .A(n3136), .B(n3790), .Z(n3791) );
  MUX21L U2902 ( .A(\gpr[12][14] ), .B(\gpr[13][14] ), .S(n3173), .Z(n3795) );
  MUX21L U2903 ( .A(\gpr[14][14] ), .B(\gpr[15][14] ), .S(n3173), .Z(n3794) );
  MUX21L U2904 ( .A(n3795), .B(n3794), .S(n3196), .Z(n3796) );
  ND2I U2905 ( .A(n3140), .B(n3796), .Z(n3801) );
  MUX21L U2906 ( .A(\gpr[16][14] ), .B(\gpr[17][14] ), .S(n3173), .Z(n3798) );
  MUX21L U2907 ( .A(\gpr[18][14] ), .B(\gpr[19][14] ), .S(n3173), .Z(n3797) );
  MUX21L U2908 ( .A(n3798), .B(n3797), .S(n3196), .Z(n3799) );
  ND2I U2909 ( .A(n3143), .B(n3799), .Z(n3800) );
  ND2I U2910 ( .A(n3801), .B(n3800), .Z(n3802) );
  NR2I U2911 ( .A(n3803), .B(n3802), .Z(n3808) );
  MUX21L U2912 ( .A(\gpr[8][14] ), .B(\gpr[9][14] ), .S(n3173), .Z(n3805) );
  MUX21L U2913 ( .A(\gpr[10][14] ), .B(\gpr[11][14] ), .S(n3173), .Z(n3804) );
  MUX21L U2914 ( .A(n3805), .B(n3804), .S(n3191), .Z(n3806) );
  ND2I U2915 ( .A(n3145), .B(n3806), .Z(n3807) );
  ND2I U2916 ( .A(n3808), .B(n3807), .Z(n3809) );
  ND2I U2917 ( .A(n3810), .B(n3809), .Z(n3811) );
  MUX21L U2918 ( .A(n1147), .B(n102), .S(n3173), .Z(n3813) );
  MUX21L U2919 ( .A(n1262), .B(n1293), .S(n3005), .Z(n3812) );
  MUX21L U2920 ( .A(n3813), .B(n3812), .S(n3200), .Z(n3814) );
  ND2I U2921 ( .A(n3814), .B(n3210), .Z(n3815) );
  NR2I U2922 ( .A(n2061), .B(n3815), .Z(n3850) );
  ND2I U2923 ( .A(\gpr[1][15] ), .B(n2048), .Z(n3817) );
  MUX21L U2924 ( .A(\gpr[2][15] ), .B(\gpr[3][15] ), .S(n2071), .Z(n3816) );
  MUX21L U2925 ( .A(n3817), .B(n3816), .S(n2049), .Z(n3818) );
  NR2I U2926 ( .A(n3818), .B(n3210), .Z(n3819) );
  ND2I U2927 ( .A(n3819), .B(n2066), .Z(n3848) );
  MUX21L U2928 ( .A(\gpr[20][15] ), .B(\gpr[21][15] ), .S(n3162), .Z(n3821) );
  MUX21L U2929 ( .A(\gpr[22][15] ), .B(\gpr[23][15] ), .S(n3161), .Z(n3820) );
  ND2I U2930 ( .A(n2094), .B(n3822), .Z(n3831) );
  MUX21L U2931 ( .A(\gpr[24][15] ), .B(\gpr[25][15] ), .S(n3162), .Z(n3824) );
  MUX21L U2932 ( .A(\gpr[26][15] ), .B(\gpr[27][15] ), .S(n2088), .Z(n3823) );
  MUX21L U2933 ( .A(n3824), .B(n3823), .S(n2050), .Z(n3825) );
  ND2I U2934 ( .A(n2022), .B(n3825), .Z(n3830) );
  MUX21L U2935 ( .A(\gpr[28][15] ), .B(\gpr[29][15] ), .S(n2088), .Z(n3827) );
  MUX21L U2936 ( .A(\gpr[30][15] ), .B(\gpr[31][15] ), .S(n3176), .Z(n3826) );
  MUX21L U2937 ( .A(n3827), .B(n3826), .S(n3192), .Z(n3828) );
  ND2I U2938 ( .A(n3135), .B(n3828), .Z(n3829) );
  MUX21L U2939 ( .A(\gpr[12][15] ), .B(\gpr[13][15] ), .S(n3159), .Z(n3833) );
  MUX21L U2940 ( .A(\gpr[14][15] ), .B(\gpr[15][15] ), .S(n3174), .Z(n3832) );
  ND2I U2941 ( .A(n3140), .B(n3834), .Z(n3839) );
  MUX21L U2942 ( .A(\gpr[16][15] ), .B(\gpr[17][15] ), .S(n3159), .Z(n3836) );
  MUX21L U2943 ( .A(\gpr[18][15] ), .B(\gpr[19][15] ), .S(n3174), .Z(n3835) );
  MUX21L U2944 ( .A(n3836), .B(n3835), .S(n2), .Z(n3837) );
  ND2I U2945 ( .A(n3143), .B(n3837), .Z(n3838) );
  ND2I U2946 ( .A(n3839), .B(n3838), .Z(n3840) );
  NR2I U2947 ( .A(n3841), .B(n3840), .Z(n3846) );
  MUX21L U2948 ( .A(\gpr[8][15] ), .B(\gpr[9][15] ), .S(n3174), .Z(n3843) );
  MUX21L U2949 ( .A(\gpr[10][15] ), .B(\gpr[11][15] ), .S(n3159), .Z(n3842) );
  MUX21L U2950 ( .A(n3843), .B(n3842), .S(n3192), .Z(n3844) );
  ND2I U2951 ( .A(n3145), .B(n3844), .Z(n3845) );
  ND2I U2952 ( .A(n3846), .B(n3845), .Z(n3847) );
  ND2I U2953 ( .A(n3848), .B(n3847), .Z(n3849) );
  NR2I U2954 ( .A(n3850), .B(n3849), .Z(rd_data1[15]) );
  MUX21L U2955 ( .A(n1148), .B(n87), .S(n3174), .Z(n3852) );
  MUX21L U2956 ( .A(n1263), .B(n1294), .S(n3159), .Z(n3851) );
  ND2I U2957 ( .A(n3853), .B(n3210), .Z(n3854) );
  NR2I U2958 ( .A(n2057), .B(n3854), .Z(n3889) );
  ND2I U2959 ( .A(\gpr[1][16] ), .B(n3180), .Z(n3856) );
  MUX21L U2960 ( .A(\gpr[2][16] ), .B(\gpr[3][16] ), .S(n3159), .Z(n3855) );
  NR2I U2961 ( .A(n3857), .B(n3210), .Z(n3858) );
  ND2I U2962 ( .A(n3858), .B(n2064), .Z(n3887) );
  MUX21L U2963 ( .A(\gpr[20][16] ), .B(\gpr[21][16] ), .S(n3160), .Z(n3860) );
  MUX21L U2964 ( .A(\gpr[22][16] ), .B(\gpr[23][16] ), .S(n3160), .Z(n3859) );
  MUX21L U2965 ( .A(n3860), .B(n3859), .S(n3200), .Z(n3861) );
  ND2I U2966 ( .A(n2095), .B(n3861), .Z(n3870) );
  MUX21L U2967 ( .A(\gpr[24][16] ), .B(\gpr[25][16] ), .S(n3160), .Z(n3863) );
  MUX21L U2968 ( .A(\gpr[26][16] ), .B(\gpr[27][16] ), .S(n3160), .Z(n3862) );
  MUX21L U2969 ( .A(n3863), .B(n3862), .S(n3200), .Z(n3864) );
  ND2I U2970 ( .A(n2076), .B(n3864), .Z(n3869) );
  MUX21L U2971 ( .A(\gpr[28][16] ), .B(\gpr[29][16] ), .S(n3160), .Z(n3866) );
  MUX21L U2972 ( .A(\gpr[30][16] ), .B(\gpr[31][16] ), .S(n3160), .Z(n3865) );
  MUX21L U2973 ( .A(n3866), .B(n3865), .S(n3200), .Z(n3867) );
  ND2I U2974 ( .A(n3137), .B(n3867), .Z(n3868) );
  MUX21L U2975 ( .A(\gpr[12][16] ), .B(\gpr[13][16] ), .S(n3159), .Z(n3872) );
  MUX21L U2976 ( .A(\gpr[14][16] ), .B(\gpr[15][16] ), .S(n3174), .Z(n3871) );
  ND2I U2977 ( .A(n3140), .B(n3873), .Z(n3878) );
  MUX21L U2978 ( .A(\gpr[16][16] ), .B(\gpr[17][16] ), .S(n3159), .Z(n3875) );
  MUX21L U2979 ( .A(\gpr[18][16] ), .B(\gpr[19][16] ), .S(n3155), .Z(n3874) );
  ND2I U2980 ( .A(n3143), .B(n3876), .Z(n3877) );
  ND2I U2981 ( .A(n3878), .B(n3877), .Z(n3879) );
  NR2I U2982 ( .A(n3880), .B(n3879), .Z(n3885) );
  MUX21L U2983 ( .A(\gpr[8][16] ), .B(\gpr[9][16] ), .S(n3174), .Z(n3882) );
  MUX21L U2984 ( .A(\gpr[10][16] ), .B(\gpr[11][16] ), .S(n3159), .Z(n3881) );
  ND2I U2985 ( .A(n3145), .B(n3883), .Z(n3884) );
  ND2I U2986 ( .A(n3885), .B(n3884), .Z(n3886) );
  ND2I U2987 ( .A(n3887), .B(n3886), .Z(n3888) );
  NR2I U2988 ( .A(n3889), .B(n3888), .Z(rd_data1[16]) );
  MUX21L U2989 ( .A(n1166), .B(n103), .S(n3174), .Z(n3891) );
  MUX21L U2990 ( .A(n1264), .B(n1295), .S(n3159), .Z(n3890) );
  ND2I U2991 ( .A(n3892), .B(n3210), .Z(n3893) );
  NR2I U2992 ( .A(n2065), .B(n3893), .Z(n3928) );
  ND2I U2993 ( .A(\gpr[1][17] ), .B(n3178), .Z(n3895) );
  MUX21L U2994 ( .A(\gpr[2][17] ), .B(\gpr[3][17] ), .S(n3159), .Z(n3894) );
  MUX21L U2995 ( .A(n3895), .B(n3894), .S(n3200), .Z(n3896) );
  NR2I U2996 ( .A(n3896), .B(n3210), .Z(n3897) );
  ND2I U2997 ( .A(n3897), .B(n2062), .Z(n3926) );
  MUX21L U2998 ( .A(\gpr[20][17] ), .B(\gpr[21][17] ), .S(n3157), .Z(n3899) );
  MUX21L U2999 ( .A(\gpr[22][17] ), .B(\gpr[23][17] ), .S(n3157), .Z(n3898) );
  MUX21L U3000 ( .A(n3899), .B(n3898), .S(n3200), .Z(n3900) );
  ND2I U3001 ( .A(n2096), .B(n3900), .Z(n3909) );
  MUX21L U3002 ( .A(\gpr[24][17] ), .B(\gpr[25][17] ), .S(n3157), .Z(n3902) );
  MUX21L U3003 ( .A(\gpr[26][17] ), .B(\gpr[27][17] ), .S(n3157), .Z(n3901) );
  MUX21L U3004 ( .A(n3902), .B(n3901), .S(n3200), .Z(n3903) );
  ND2I U3005 ( .A(n2077), .B(n3903), .Z(n3908) );
  MUX21L U3006 ( .A(\gpr[28][17] ), .B(\gpr[29][17] ), .S(n3157), .Z(n3905) );
  MUX21L U3007 ( .A(\gpr[30][17] ), .B(\gpr[31][17] ), .S(n3157), .Z(n3904) );
  MUX21L U3008 ( .A(n3905), .B(n3904), .S(n3200), .Z(n3906) );
  ND2I U3009 ( .A(n3138), .B(n3906), .Z(n3907) );
  MUX21L U3010 ( .A(\gpr[12][17] ), .B(\gpr[13][17] ), .S(n3159), .Z(n3911) );
  MUX21L U3011 ( .A(\gpr[14][17] ), .B(\gpr[15][17] ), .S(n3174), .Z(n3910) );
  MUX21L U3012 ( .A(n3911), .B(n3910), .S(n3200), .Z(n3912) );
  ND2I U3013 ( .A(n3140), .B(n3912), .Z(n3917) );
  MUX21L U3014 ( .A(\gpr[16][17] ), .B(\gpr[17][17] ), .S(n3159), .Z(n3914) );
  MUX21L U3015 ( .A(\gpr[18][17] ), .B(\gpr[19][17] ), .S(n3174), .Z(n3913) );
  MUX21L U3016 ( .A(n3914), .B(n3913), .S(n3200), .Z(n3915) );
  ND2I U3017 ( .A(n3143), .B(n3915), .Z(n3916) );
  ND2I U3018 ( .A(n3917), .B(n3916), .Z(n3918) );
  NR2I U3019 ( .A(n3919), .B(n3918), .Z(n3924) );
  MUX21L U3020 ( .A(\gpr[8][17] ), .B(\gpr[9][17] ), .S(n3174), .Z(n3921) );
  MUX21L U3021 ( .A(\gpr[10][17] ), .B(\gpr[11][17] ), .S(n3159), .Z(n3920) );
  MUX21L U3022 ( .A(n3921), .B(n3920), .S(n3200), .Z(n3922) );
  ND2I U3023 ( .A(n3145), .B(n3922), .Z(n3923) );
  ND2I U3024 ( .A(n3924), .B(n3923), .Z(n3925) );
  ND2I U3025 ( .A(n3926), .B(n3925), .Z(n3927) );
  NR2I U3026 ( .A(n3928), .B(n3927), .Z(rd_data1[17]) );
  MUX21L U3027 ( .A(n1167), .B(n104), .S(n3174), .Z(n3930) );
  MUX21L U3028 ( .A(n1265), .B(n1296), .S(n3159), .Z(n3929) );
  ND2I U3029 ( .A(n3931), .B(n3210), .Z(n3932) );
  NR2I U3030 ( .A(n2065), .B(n3932), .Z(n3967) );
  ND2I U3031 ( .A(\gpr[1][18] ), .B(n3178), .Z(n3934) );
  MUX21L U3032 ( .A(\gpr[2][18] ), .B(\gpr[3][18] ), .S(n3174), .Z(n3933) );
  NR2I U3033 ( .A(n3935), .B(n3210), .Z(n3936) );
  ND2I U3034 ( .A(n3936), .B(n2058), .Z(n3965) );
  MUX21L U3035 ( .A(\gpr[20][18] ), .B(\gpr[21][18] ), .S(n3160), .Z(n3938) );
  MUX21L U3036 ( .A(\gpr[22][18] ), .B(\gpr[23][18] ), .S(n3158), .Z(n3937) );
  MUX21L U3037 ( .A(n3938), .B(n3937), .S(n3200), .Z(n3939) );
  ND2I U3038 ( .A(n2097), .B(n3939), .Z(n3948) );
  MUX21L U3039 ( .A(\gpr[24][18] ), .B(\gpr[25][18] ), .S(n3158), .Z(n3941) );
  MUX21L U3040 ( .A(\gpr[26][18] ), .B(\gpr[27][18] ), .S(n3158), .Z(n3940) );
  MUX21L U3041 ( .A(n3941), .B(n3940), .S(n3199), .Z(n3942) );
  ND2I U3042 ( .A(n2022), .B(n3942), .Z(n3947) );
  MUX21L U3043 ( .A(\gpr[28][18] ), .B(\gpr[29][18] ), .S(n3158), .Z(n3944) );
  MUX21L U3044 ( .A(\gpr[30][18] ), .B(\gpr[31][18] ), .S(n3158), .Z(n3943) );
  MUX21L U3045 ( .A(n3944), .B(n3943), .S(n3199), .Z(n3945) );
  ND2I U3046 ( .A(n3135), .B(n3945), .Z(n3946) );
  MUX21L U3047 ( .A(\gpr[12][18] ), .B(\gpr[13][18] ), .S(n3158), .Z(n3950) );
  MUX21L U3048 ( .A(\gpr[14][18] ), .B(\gpr[15][18] ), .S(n3158), .Z(n3949) );
  MUX21L U3049 ( .A(n3950), .B(n3949), .S(n3199), .Z(n3951) );
  ND2I U3050 ( .A(n3140), .B(n3951), .Z(n3956) );
  MUX21L U3051 ( .A(\gpr[16][18] ), .B(\gpr[17][18] ), .S(n3158), .Z(n3953) );
  MUX21L U3052 ( .A(\gpr[18][18] ), .B(\gpr[19][18] ), .S(n3158), .Z(n3952) );
  MUX21L U3053 ( .A(n3953), .B(n3952), .S(n3199), .Z(n3954) );
  ND2I U3054 ( .A(n3143), .B(n3954), .Z(n3955) );
  ND2I U3055 ( .A(n3956), .B(n3955), .Z(n3957) );
  NR2I U3056 ( .A(n3958), .B(n3957), .Z(n3963) );
  MUX21L U3057 ( .A(\gpr[8][18] ), .B(\gpr[9][18] ), .S(n3158), .Z(n3960) );
  MUX21L U3058 ( .A(\gpr[10][18] ), .B(\gpr[11][18] ), .S(n3158), .Z(n3959) );
  MUX21L U3059 ( .A(n3960), .B(n3959), .S(n3199), .Z(n3961) );
  ND2I U3060 ( .A(n3145), .B(n3961), .Z(n3962) );
  ND2I U3061 ( .A(n3963), .B(n3962), .Z(n3964) );
  ND2I U3062 ( .A(n3965), .B(n3964), .Z(n3966) );
  NR2I U3063 ( .A(n3967), .B(n3966), .Z(rd_data1[18]) );
  MUX21L U3064 ( .A(n1149), .B(n88), .S(n3158), .Z(n3969) );
  MUX21L U3065 ( .A(n1266), .B(n1297), .S(n3158), .Z(n3968) );
  MUX21L U3066 ( .A(n3969), .B(n3968), .S(n3199), .Z(n3970) );
  ND2I U3067 ( .A(n3970), .B(n3210), .Z(n3971) );
  NR2I U3068 ( .A(n2059), .B(n3971), .Z(n4006) );
  ND2I U3069 ( .A(\gpr[1][19] ), .B(n2041), .Z(n3973) );
  MUX21L U3070 ( .A(\gpr[2][19] ), .B(\gpr[3][19] ), .S(n3158), .Z(n3972) );
  MUX21L U3071 ( .A(n3973), .B(n3972), .S(n3199), .Z(n3974) );
  NR2I U3072 ( .A(n3974), .B(n3210), .Z(n3975) );
  ND2I U3073 ( .A(n3975), .B(n2060), .Z(n4004) );
  MUX21L U3074 ( .A(\gpr[20][19] ), .B(\gpr[21][19] ), .S(n3160), .Z(n3977) );
  MUX21L U3075 ( .A(\gpr[22][19] ), .B(\gpr[23][19] ), .S(n3160), .Z(n3976) );
  MUX21L U3076 ( .A(n3977), .B(n3976), .S(n3199), .Z(n3978) );
  ND2I U3077 ( .A(n2098), .B(n3978), .Z(n3987) );
  MUX21L U3078 ( .A(\gpr[24][19] ), .B(\gpr[25][19] ), .S(n3160), .Z(n3980) );
  MUX21L U3079 ( .A(\gpr[26][19] ), .B(\gpr[27][19] ), .S(n3160), .Z(n3979) );
  MUX21L U3080 ( .A(n3980), .B(n3979), .S(n3199), .Z(n3981) );
  ND2I U3081 ( .A(n2022), .B(n3981), .Z(n3986) );
  MUX21L U3082 ( .A(\gpr[28][19] ), .B(\gpr[29][19] ), .S(n3160), .Z(n3983) );
  MUX21L U3083 ( .A(\gpr[30][19] ), .B(\gpr[31][19] ), .S(n3160), .Z(n3982) );
  MUX21L U3084 ( .A(n3983), .B(n3982), .S(n3199), .Z(n3984) );
  ND2I U3085 ( .A(n3137), .B(n3984), .Z(n3985) );
  MUX21L U3086 ( .A(\gpr[12][19] ), .B(\gpr[13][19] ), .S(n3157), .Z(n3989) );
  MUX21L U3087 ( .A(\gpr[14][19] ), .B(\gpr[15][19] ), .S(n3157), .Z(n3988) );
  MUX21L U3088 ( .A(n3989), .B(n3988), .S(n3199), .Z(n3990) );
  ND2I U3089 ( .A(n3140), .B(n3990), .Z(n3995) );
  MUX21L U3090 ( .A(\gpr[16][19] ), .B(\gpr[17][19] ), .S(n3157), .Z(n3992) );
  MUX21L U3091 ( .A(\gpr[18][19] ), .B(\gpr[19][19] ), .S(n3157), .Z(n3991) );
  MUX21L U3092 ( .A(n3992), .B(n3991), .S(n3199), .Z(n3993) );
  ND2I U3093 ( .A(n3143), .B(n3993), .Z(n3994) );
  ND2I U3094 ( .A(n3995), .B(n3994), .Z(n3996) );
  NR2I U3095 ( .A(n3997), .B(n3996), .Z(n4002) );
  MUX21L U3096 ( .A(\gpr[8][19] ), .B(\gpr[9][19] ), .S(n3157), .Z(n3999) );
  MUX21L U3097 ( .A(\gpr[10][19] ), .B(\gpr[11][19] ), .S(n3157), .Z(n3998) );
  MUX21L U3098 ( .A(n3999), .B(n3998), .S(n3199), .Z(n4000) );
  ND2I U3099 ( .A(n3145), .B(n4000), .Z(n4001) );
  ND2I U3100 ( .A(n4002), .B(n4001), .Z(n4003) );
  ND2I U3101 ( .A(n4004), .B(n4003), .Z(n4005) );
  NR2I U3102 ( .A(n4006), .B(n4005), .Z(rd_data1[19]) );
  MUX21L U3103 ( .A(n1168), .B(n105), .S(n3157), .Z(n4008) );
  MUX21L U3104 ( .A(n1267), .B(n1298), .S(n3156), .Z(n4007) );
  ND2I U3105 ( .A(n4009), .B(n3209), .Z(n4010) );
  NR2I U3106 ( .A(n2055), .B(n4010), .Z(n4045) );
  ND2I U3107 ( .A(\gpr[1][20] ), .B(n3178), .Z(n4012) );
  MUX21L U3108 ( .A(\gpr[2][20] ), .B(\gpr[3][20] ), .S(n3156), .Z(n4011) );
  MUX21L U3109 ( .A(n4012), .B(n4011), .S(n3199), .Z(n4013) );
  NR2I U3110 ( .A(n4013), .B(n3210), .Z(n4014) );
  ND2I U3111 ( .A(n4014), .B(n2066), .Z(n4043) );
  MUX21L U3112 ( .A(\gpr[20][20] ), .B(\gpr[21][20] ), .S(n3156), .Z(n4016) );
  MUX21L U3113 ( .A(\gpr[22][20] ), .B(\gpr[23][20] ), .S(n3156), .Z(n4015) );
  MUX21L U3114 ( .A(n4016), .B(n4015), .S(n3199), .Z(n4017) );
  ND2I U3115 ( .A(n2096), .B(n4017), .Z(n4026) );
  MUX21L U3116 ( .A(\gpr[24][20] ), .B(\gpr[25][20] ), .S(n3156), .Z(n4019) );
  MUX21L U3117 ( .A(\gpr[26][20] ), .B(\gpr[27][20] ), .S(n3156), .Z(n4018) );
  MUX21L U3118 ( .A(n4019), .B(n4018), .S(n3199), .Z(n4020) );
  ND2I U3119 ( .A(n2022), .B(n4020), .Z(n4025) );
  MUX21L U3120 ( .A(\gpr[28][20] ), .B(\gpr[29][20] ), .S(n3156), .Z(n4022) );
  MUX21L U3121 ( .A(\gpr[30][20] ), .B(\gpr[31][20] ), .S(n3156), .Z(n4021) );
  MUX21L U3122 ( .A(n4022), .B(n4021), .S(n3199), .Z(n4023) );
  ND2I U3123 ( .A(n3138), .B(n4023), .Z(n4024) );
  MUX21L U3124 ( .A(\gpr[12][20] ), .B(\gpr[13][20] ), .S(n3156), .Z(n4028) );
  MUX21L U3125 ( .A(\gpr[14][20] ), .B(\gpr[15][20] ), .S(n3156), .Z(n4027) );
  MUX21L U3126 ( .A(n4028), .B(n4027), .S(n3199), .Z(n4029) );
  ND2I U3127 ( .A(n3140), .B(n4029), .Z(n4034) );
  MUX21L U3128 ( .A(\gpr[16][20] ), .B(\gpr[17][20] ), .S(n3156), .Z(n4031) );
  MUX21L U3129 ( .A(\gpr[18][20] ), .B(\gpr[19][20] ), .S(n3156), .Z(n4030) );
  MUX21L U3130 ( .A(n4031), .B(n4030), .S(n3198), .Z(n4032) );
  ND2I U3131 ( .A(n3143), .B(n4032), .Z(n4033) );
  ND2I U3132 ( .A(n4034), .B(n4033), .Z(n4035) );
  NR2I U3133 ( .A(n4036), .B(n4035), .Z(n4041) );
  MUX21L U3134 ( .A(\gpr[8][20] ), .B(\gpr[9][20] ), .S(n3156), .Z(n4038) );
  MUX21L U3135 ( .A(\gpr[10][20] ), .B(\gpr[11][20] ), .S(n3156), .Z(n4037) );
  MUX21L U3136 ( .A(n4038), .B(n4037), .S(n3198), .Z(n4039) );
  ND2I U3137 ( .A(n3145), .B(n4039), .Z(n4040) );
  ND2I U3138 ( .A(n4041), .B(n4040), .Z(n4042) );
  ND2I U3139 ( .A(n4043), .B(n4042), .Z(n4044) );
  NR2I U3140 ( .A(n4045), .B(n4044), .Z(rd_data1[20]) );
  MUX21L U3141 ( .A(n1150), .B(n89), .S(n3155), .Z(n4047) );
  MUX21L U3142 ( .A(n1268), .B(n1299), .S(n3155), .Z(n4046) );
  MUX21L U3143 ( .A(n4047), .B(n4046), .S(n3198), .Z(n4048) );
  ND2I U3144 ( .A(n4048), .B(n3208), .Z(n4049) );
  NR2I U3145 ( .A(n2055), .B(n4049), .Z(n4084) );
  ND2I U3146 ( .A(\gpr[1][21] ), .B(n3180), .Z(n4051) );
  MUX21L U3147 ( .A(\gpr[2][21] ), .B(\gpr[3][21] ), .S(n3155), .Z(n4050) );
  MUX21L U3148 ( .A(n4051), .B(n4050), .S(n3198), .Z(n4052) );
  NR2I U3149 ( .A(n4052), .B(n3210), .Z(n4053) );
  ND2I U3150 ( .A(n4053), .B(n2066), .Z(n4082) );
  MUX21L U3151 ( .A(\gpr[20][21] ), .B(\gpr[21][21] ), .S(n3154), .Z(n4055) );
  MUX21L U3152 ( .A(\gpr[22][21] ), .B(\gpr[23][21] ), .S(n3154), .Z(n4054) );
  MUX21L U3153 ( .A(n4055), .B(n4054), .S(n3191), .Z(n4056) );
  ND2I U3154 ( .A(n2096), .B(n4056), .Z(n4065) );
  MUX21L U3155 ( .A(\gpr[24][21] ), .B(\gpr[25][21] ), .S(n3154), .Z(n4058) );
  MUX21L U3156 ( .A(\gpr[26][21] ), .B(\gpr[27][21] ), .S(n3154), .Z(n4057) );
  MUX21L U3157 ( .A(n4058), .B(n4057), .S(n3191), .Z(n4059) );
  ND2I U3158 ( .A(n2076), .B(n4059), .Z(n4064) );
  MUX21L U3159 ( .A(\gpr[28][21] ), .B(\gpr[29][21] ), .S(n3154), .Z(n4061) );
  MUX21L U3160 ( .A(\gpr[30][21] ), .B(\gpr[31][21] ), .S(n3154), .Z(n4060) );
  MUX21L U3161 ( .A(n4061), .B(n4060), .S(n3191), .Z(n4062) );
  ND2I U3162 ( .A(n3137), .B(n4062), .Z(n4063) );
  MUX21L U3163 ( .A(\gpr[12][21] ), .B(\gpr[13][21] ), .S(n3155), .Z(n4067) );
  MUX21L U3164 ( .A(\gpr[14][21] ), .B(\gpr[15][21] ), .S(n3155), .Z(n4066) );
  MUX21L U3165 ( .A(n4067), .B(n4066), .S(n3198), .Z(n4068) );
  ND2I U3166 ( .A(n3141), .B(n4068), .Z(n4073) );
  MUX21L U3167 ( .A(\gpr[16][21] ), .B(\gpr[17][21] ), .S(n3155), .Z(n4070) );
  MUX21L U3168 ( .A(\gpr[18][21] ), .B(\gpr[19][21] ), .S(n3155), .Z(n4069) );
  MUX21L U3169 ( .A(n4070), .B(n4069), .S(n3198), .Z(n4071) );
  ND2I U3170 ( .A(n3144), .B(n4071), .Z(n4072) );
  ND2I U3171 ( .A(n4073), .B(n4072), .Z(n4074) );
  NR2I U3172 ( .A(n4075), .B(n4074), .Z(n4080) );
  MUX21L U3173 ( .A(\gpr[8][21] ), .B(\gpr[9][21] ), .S(n3155), .Z(n4077) );
  MUX21L U3174 ( .A(\gpr[10][21] ), .B(\gpr[11][21] ), .S(n3155), .Z(n4076) );
  MUX21L U3175 ( .A(n4077), .B(n4076), .S(n3198), .Z(n4078) );
  ND2I U3176 ( .A(n3146), .B(n4078), .Z(n4079) );
  ND2I U3177 ( .A(n4080), .B(n4079), .Z(n4081) );
  ND2I U3178 ( .A(n4082), .B(n4081), .Z(n4083) );
  NR2I U3179 ( .A(n4084), .B(n4083), .Z(rd_data1[21]) );
  MUX21L U3180 ( .A(n1169), .B(n106), .S(n3155), .Z(n4086) );
  MUX21L U3181 ( .A(n1269), .B(n1300), .S(n3155), .Z(n4085) );
  MUX21L U3182 ( .A(n4086), .B(n4085), .S(n3198), .Z(n4087) );
  ND2I U3183 ( .A(n4087), .B(n3210), .Z(n4088) );
  NR2I U3184 ( .A(n2061), .B(n4088), .Z(n4123) );
  ND2I U3185 ( .A(\gpr[1][22] ), .B(n2040), .Z(n4090) );
  MUX21L U3186 ( .A(\gpr[2][22] ), .B(\gpr[3][22] ), .S(n3155), .Z(n4089) );
  MUX21L U3187 ( .A(n4090), .B(n4089), .S(n3198), .Z(n4091) );
  NR2I U3188 ( .A(n4091), .B(n3209), .Z(n4092) );
  ND2I U3189 ( .A(n4092), .B(n2064), .Z(n4121) );
  MUX21L U3190 ( .A(\gpr[20][22] ), .B(\gpr[21][22] ), .S(n3154), .Z(n4094) );
  MUX21L U3191 ( .A(\gpr[22][22] ), .B(\gpr[23][22] ), .S(n3154), .Z(n4093) );
  MUX21L U3192 ( .A(n4094), .B(n4093), .S(n3196), .Z(n4095) );
  ND2I U3193 ( .A(n2097), .B(n4095), .Z(n4104) );
  MUX21L U3194 ( .A(\gpr[24][22] ), .B(\gpr[25][22] ), .S(n3154), .Z(n4097) );
  MUX21L U3195 ( .A(\gpr[26][22] ), .B(\gpr[27][22] ), .S(n3154), .Z(n4096) );
  MUX21L U3196 ( .A(n4097), .B(n4096), .S(n3194), .Z(n4098) );
  ND2I U3197 ( .A(n2074), .B(n4098), .Z(n4103) );
  MUX21L U3198 ( .A(\gpr[28][22] ), .B(\gpr[29][22] ), .S(n3154), .Z(n4100) );
  MUX21L U3199 ( .A(\gpr[30][22] ), .B(\gpr[31][22] ), .S(n3155), .Z(n4099) );
  MUX21L U3200 ( .A(n4100), .B(n4099), .S(n3191), .Z(n4101) );
  ND2I U3201 ( .A(n3138), .B(n4101), .Z(n4102) );
  MUX21L U3202 ( .A(\gpr[12][22] ), .B(\gpr[13][22] ), .S(n3155), .Z(n4106) );
  MUX21L U3203 ( .A(\gpr[14][22] ), .B(\gpr[15][22] ), .S(n3155), .Z(n4105) );
  MUX21L U3204 ( .A(n4106), .B(n4105), .S(n3198), .Z(n4107) );
  ND2I U3205 ( .A(n3141), .B(n4107), .Z(n4112) );
  MUX21L U3206 ( .A(\gpr[16][22] ), .B(\gpr[17][22] ), .S(n3155), .Z(n4109) );
  MUX21L U3207 ( .A(\gpr[18][22] ), .B(\gpr[19][22] ), .S(n3155), .Z(n4108) );
  MUX21L U3208 ( .A(n4109), .B(n4108), .S(n3198), .Z(n4110) );
  ND2I U3209 ( .A(n3144), .B(n4110), .Z(n4111) );
  ND2I U3210 ( .A(n4112), .B(n4111), .Z(n4113) );
  NR2I U3211 ( .A(n4114), .B(n4113), .Z(n4119) );
  MUX21L U3212 ( .A(\gpr[8][22] ), .B(\gpr[9][22] ), .S(n3153), .Z(n4116) );
  MUX21L U3213 ( .A(\gpr[10][22] ), .B(\gpr[11][22] ), .S(n3153), .Z(n4115) );
  MUX21L U3214 ( .A(n4116), .B(n4115), .S(n3198), .Z(n4117) );
  ND2I U3215 ( .A(n3146), .B(n4117), .Z(n4118) );
  ND2I U3216 ( .A(n4119), .B(n4118), .Z(n4120) );
  ND2I U3217 ( .A(n4121), .B(n4120), .Z(n4122) );
  NR2I U3218 ( .A(n4123), .B(n4122), .Z(rd_data1[22]) );
  MUX21L U3219 ( .A(n1151), .B(n90), .S(n3153), .Z(n4125) );
  MUX21L U3220 ( .A(n1270), .B(n1301), .S(n3153), .Z(n4124) );
  MUX21L U3221 ( .A(n4125), .B(n4124), .S(n3198), .Z(n4126) );
  ND2I U3222 ( .A(n4126), .B(n3209), .Z(n4127) );
  NR2I U3223 ( .A(n2061), .B(n4127), .Z(n4162) );
  ND2I U3224 ( .A(\gpr[1][23] ), .B(n2040), .Z(n4129) );
  MUX21L U3225 ( .A(\gpr[2][23] ), .B(\gpr[3][23] ), .S(n3153), .Z(n4128) );
  MUX21L U3226 ( .A(n4129), .B(n4128), .S(n3198), .Z(n4130) );
  NR2I U3227 ( .A(n4130), .B(n3210), .Z(n4131) );
  ND2I U3228 ( .A(n4131), .B(n2066), .Z(n4160) );
  MUX21L U3229 ( .A(\gpr[20][23] ), .B(\gpr[21][23] ), .S(n3153), .Z(n4133) );
  MUX21L U3230 ( .A(\gpr[22][23] ), .B(\gpr[23][23] ), .S(n3153), .Z(n4132) );
  ND2I U3231 ( .A(n2098), .B(n4134), .Z(n4143) );
  MUX21L U3232 ( .A(\gpr[24][23] ), .B(\gpr[25][23] ), .S(n3153), .Z(n4136) );
  MUX21L U3233 ( .A(\gpr[26][23] ), .B(\gpr[27][23] ), .S(n3153), .Z(n4135) );
  MUX21L U3234 ( .A(n4136), .B(n4135), .S(n3191), .Z(n4137) );
  ND2I U3235 ( .A(n2076), .B(n4137), .Z(n4142) );
  MUX21L U3236 ( .A(\gpr[28][23] ), .B(\gpr[29][23] ), .S(n3153), .Z(n4139) );
  MUX21L U3237 ( .A(\gpr[30][23] ), .B(\gpr[31][23] ), .S(n3153), .Z(n4138) );
  MUX21L U3238 ( .A(n4139), .B(n4138), .S(n3200), .Z(n4140) );
  ND2I U3239 ( .A(n3135), .B(n4140), .Z(n4141) );
  MUX21L U3240 ( .A(\gpr[12][23] ), .B(\gpr[13][23] ), .S(n3153), .Z(n4145) );
  MUX21L U3241 ( .A(\gpr[14][23] ), .B(\gpr[15][23] ), .S(n3153), .Z(n4144) );
  MUX21L U3242 ( .A(n4145), .B(n4144), .S(n3198), .Z(n4146) );
  ND2I U3243 ( .A(n3141), .B(n4146), .Z(n4151) );
  MUX21L U3244 ( .A(\gpr[16][23] ), .B(\gpr[17][23] ), .S(n3157), .Z(n4148) );
  MUX21L U3245 ( .A(\gpr[18][23] ), .B(\gpr[19][23] ), .S(n3166), .Z(n4147) );
  MUX21L U3246 ( .A(n4148), .B(n4147), .S(n3198), .Z(n4149) );
  ND2I U3247 ( .A(n3144), .B(n4149), .Z(n4150) );
  ND2I U3248 ( .A(n4151), .B(n4150), .Z(n4152) );
  NR2I U3249 ( .A(n4153), .B(n4152), .Z(n4158) );
  MUX21L U3250 ( .A(\gpr[8][23] ), .B(\gpr[9][23] ), .S(n3178), .Z(n4155) );
  MUX21L U3251 ( .A(\gpr[10][23] ), .B(\gpr[11][23] ), .S(n3166), .Z(n4154) );
  MUX21L U3252 ( .A(n4155), .B(n4154), .S(n3198), .Z(n4156) );
  ND2I U3253 ( .A(n3146), .B(n4156), .Z(n4157) );
  ND2I U3254 ( .A(n4158), .B(n4157), .Z(n4159) );
  ND2I U3255 ( .A(n4160), .B(n4159), .Z(n4161) );
  NR2I U3256 ( .A(n4162), .B(n4161), .Z(rd_data1[23]) );
  MUX21L U3257 ( .A(n1170), .B(n107), .S(n3178), .Z(n4164) );
  MUX21L U3258 ( .A(n1271), .B(n1302), .S(n3166), .Z(n4163) );
  MUX21L U3259 ( .A(n4164), .B(n4163), .S(n3198), .Z(n4165) );
  ND2I U3260 ( .A(n4165), .B(n3211), .Z(n4166) );
  NR2I U3261 ( .A(n2063), .B(n4166), .Z(n4201) );
  ND2I U3262 ( .A(\gpr[1][24] ), .B(n2021), .Z(n4168) );
  MUX21L U3263 ( .A(\gpr[2][24] ), .B(\gpr[3][24] ), .S(n3166), .Z(n4167) );
  MUX21L U3264 ( .A(n4168), .B(n4167), .S(n3198), .Z(n4169) );
  NR2I U3265 ( .A(n4169), .B(n3211), .Z(n4170) );
  ND2I U3266 ( .A(n4170), .B(n2058), .Z(n4199) );
  MUX21L U3267 ( .A(\gpr[20][24] ), .B(\gpr[21][24] ), .S(n3179), .Z(n4172) );
  MUX21L U3268 ( .A(\gpr[22][24] ), .B(\gpr[23][24] ), .S(n2040), .Z(n4171) );
  MUX21L U3269 ( .A(n4172), .B(n4171), .S(n2050), .Z(n4173) );
  ND2I U3270 ( .A(n2099), .B(n4173), .Z(n4182) );
  MUX21L U3271 ( .A(\gpr[24][24] ), .B(\gpr[25][24] ), .S(n2071), .Z(n4175) );
  MUX21L U3272 ( .A(\gpr[26][24] ), .B(\gpr[27][24] ), .S(n2101), .Z(n4174) );
  MUX21L U3273 ( .A(n4175), .B(n4174), .S(n3191), .Z(n4176) );
  ND2I U3274 ( .A(n2074), .B(n4176), .Z(n4181) );
  MUX21L U3275 ( .A(\gpr[28][24] ), .B(\gpr[29][24] ), .S(n2101), .Z(n4178) );
  MUX21L U3276 ( .A(\gpr[30][24] ), .B(\gpr[31][24] ), .S(n2101), .Z(n4177) );
  MUX21L U3277 ( .A(n4178), .B(n4177), .S(n3195), .Z(n4179) );
  ND2I U3278 ( .A(n3135), .B(n4179), .Z(n4180) );
  MUX21L U3279 ( .A(\gpr[12][24] ), .B(\gpr[13][24] ), .S(n3159), .Z(n4184) );
  MUX21L U3280 ( .A(\gpr[14][24] ), .B(\gpr[15][24] ), .S(n3166), .Z(n4183) );
  MUX21L U3281 ( .A(n4184), .B(n4183), .S(n3198), .Z(n4185) );
  ND2I U3282 ( .A(n3141), .B(n4185), .Z(n4190) );
  MUX21L U3283 ( .A(\gpr[16][24] ), .B(\gpr[17][24] ), .S(n3171), .Z(n4187) );
  MUX21L U3284 ( .A(\gpr[18][24] ), .B(\gpr[19][24] ), .S(n3166), .Z(n4186) );
  MUX21L U3285 ( .A(n4187), .B(n4186), .S(n3198), .Z(n4188) );
  ND2I U3286 ( .A(n3144), .B(n4188), .Z(n4189) );
  ND2I U3287 ( .A(n4190), .B(n4189), .Z(n4191) );
  NR2I U3288 ( .A(n4192), .B(n4191), .Z(n4197) );
  MUX21L U3289 ( .A(\gpr[8][24] ), .B(\gpr[9][24] ), .S(n3178), .Z(n4194) );
  MUX21L U3290 ( .A(\gpr[10][24] ), .B(\gpr[11][24] ), .S(n3166), .Z(n4193) );
  MUX21L U3291 ( .A(n4194), .B(n4193), .S(n3198), .Z(n4195) );
  ND2I U3292 ( .A(n3146), .B(n4195), .Z(n4196) );
  ND2I U3293 ( .A(n4197), .B(n4196), .Z(n4198) );
  ND2I U3294 ( .A(n4199), .B(n4198), .Z(n4200) );
  NR2I U3295 ( .A(n4201), .B(n4200), .Z(rd_data1[24]) );
  MUX21L U3296 ( .A(n1171), .B(n108), .S(n3178), .Z(n4203) );
  MUX21L U3297 ( .A(n1272), .B(n1303), .S(n3166), .Z(n4202) );
  MUX21L U3298 ( .A(n4203), .B(n4202), .S(n3198), .Z(n4204) );
  ND2I U3299 ( .A(n4204), .B(n3211), .Z(n4205) );
  NR2I U3300 ( .A(n2057), .B(n4205), .Z(n4240) );
  ND2I U3301 ( .A(\gpr[1][25] ), .B(n3168), .Z(n4207) );
  MUX21L U3302 ( .A(\gpr[2][25] ), .B(\gpr[3][25] ), .S(n3178), .Z(n4206) );
  MUX21L U3303 ( .A(n4207), .B(n4206), .S(n3198), .Z(n4208) );
  NR2I U3304 ( .A(n4208), .B(n3211), .Z(n4209) );
  ND2I U3305 ( .A(n4209), .B(n2056), .Z(n4238) );
  MUX21L U3306 ( .A(\gpr[20][25] ), .B(\gpr[21][25] ), .S(n2101), .Z(n4211) );
  MUX21L U3307 ( .A(\gpr[22][25] ), .B(\gpr[23][25] ), .S(n3162), .Z(n4210) );
  MUX21L U3308 ( .A(n4211), .B(n4210), .S(n3200), .Z(n4212) );
  ND2I U3309 ( .A(n2093), .B(n4212), .Z(n4221) );
  MUX21L U3310 ( .A(\gpr[24][25] ), .B(\gpr[25][25] ), .S(n2040), .Z(n4214) );
  MUX21L U3311 ( .A(\gpr[26][25] ), .B(\gpr[27][25] ), .S(n2088), .Z(n4213) );
  MUX21L U3312 ( .A(n4214), .B(n4213), .S(n3197), .Z(n4215) );
  ND2I U3313 ( .A(n2022), .B(n4215), .Z(n4220) );
  MUX21L U3314 ( .A(\gpr[28][25] ), .B(\gpr[29][25] ), .S(n2101), .Z(n4217) );
  MUX21L U3315 ( .A(\gpr[30][25] ), .B(\gpr[31][25] ), .S(n3158), .Z(n4216) );
  MUX21L U3316 ( .A(n4217), .B(n4216), .S(n3197), .Z(n4218) );
  ND2I U3317 ( .A(n3137), .B(n4218), .Z(n4219) );
  MUX21L U3318 ( .A(\gpr[12][25] ), .B(\gpr[13][25] ), .S(n3178), .Z(n4223) );
  MUX21L U3319 ( .A(\gpr[14][25] ), .B(\gpr[15][25] ), .S(n3166), .Z(n4222) );
  MUX21L U3320 ( .A(n4223), .B(n4222), .S(n3197), .Z(n4224) );
  ND2I U3321 ( .A(n3141), .B(n4224), .Z(n4229) );
  MUX21L U3322 ( .A(\gpr[16][25] ), .B(\gpr[17][25] ), .S(n3178), .Z(n4226) );
  MUX21L U3323 ( .A(\gpr[18][25] ), .B(\gpr[19][25] ), .S(n3166), .Z(n4225) );
  MUX21L U3324 ( .A(n4226), .B(n4225), .S(n3197), .Z(n4227) );
  ND2I U3325 ( .A(n3144), .B(n4227), .Z(n4228) );
  ND2I U3326 ( .A(n4229), .B(n4228), .Z(n4230) );
  NR2I U3327 ( .A(n4231), .B(n4230), .Z(n4236) );
  MUX21L U3328 ( .A(\gpr[8][25] ), .B(\gpr[9][25] ), .S(n3178), .Z(n4233) );
  MUX21L U3329 ( .A(\gpr[10][25] ), .B(\gpr[11][25] ), .S(n3166), .Z(n4232) );
  MUX21L U3330 ( .A(n4233), .B(n4232), .S(n3197), .Z(n4234) );
  ND2I U3331 ( .A(n3146), .B(n4234), .Z(n4235) );
  ND2I U3332 ( .A(n4236), .B(n4235), .Z(n4237) );
  ND2I U3333 ( .A(n4238), .B(n4237), .Z(n4239) );
  NR2I U3334 ( .A(n4240), .B(n4239), .Z(rd_data1[25]) );
  MUX21L U3335 ( .A(n1152), .B(n91), .S(n3157), .Z(n4242) );
  MUX21L U3336 ( .A(n1273), .B(n1304), .S(n3164), .Z(n4241) );
  MUX21L U3337 ( .A(n4242), .B(n4241), .S(n3197), .Z(n4243) );
  ND2I U3338 ( .A(n4243), .B(n3211), .Z(n4244) );
  NR2I U3339 ( .A(n2055), .B(n4244), .Z(n4276) );
  ND2I U3340 ( .A(\gpr[1][26] ), .B(n3168), .Z(n4246) );
  MUX21L U3341 ( .A(\gpr[2][26] ), .B(\gpr[3][26] ), .S(n3164), .Z(n4245) );
  MUX21L U3342 ( .A(n4246), .B(n4245), .S(n3197), .Z(n4247) );
  NR2I U3343 ( .A(n4247), .B(n3211), .Z(n4248) );
  MUX21L U3344 ( .A(\gpr[20][26] ), .B(\gpr[21][26] ), .S(n3164), .Z(n4250) );
  MUX21L U3345 ( .A(\gpr[22][26] ), .B(\gpr[23][26] ), .S(n3165), .Z(n4249) );
  MUX21L U3346 ( .A(n4250), .B(n4249), .S(n3197), .Z(n4251) );
  ND2I U3347 ( .A(n2094), .B(n4251), .Z(n4260) );
  MUX21L U3348 ( .A(\gpr[24][26] ), .B(\gpr[25][26] ), .S(n3164), .Z(n4253) );
  MUX21L U3349 ( .A(\gpr[26][26] ), .B(\gpr[27][26] ), .S(n3165), .Z(n4252) );
  MUX21L U3350 ( .A(n4253), .B(n4252), .S(n3197), .Z(n4254) );
  ND2I U3351 ( .A(n2075), .B(n4254), .Z(n4259) );
  MUX21L U3352 ( .A(\gpr[28][26] ), .B(\gpr[29][26] ), .S(n3164), .Z(n4256) );
  MUX21L U3353 ( .A(\gpr[30][26] ), .B(\gpr[31][26] ), .S(n3165), .Z(n4255) );
  MUX21L U3354 ( .A(n4256), .B(n4255), .S(n3197), .Z(n4257) );
  ND2I U3355 ( .A(n3138), .B(n4257), .Z(n4258) );
  MUX21L U3356 ( .A(\gpr[12][26] ), .B(\gpr[13][26] ), .S(n3164), .Z(n4262) );
  MUX21L U3357 ( .A(\gpr[14][26] ), .B(\gpr[15][26] ), .S(n3165), .Z(n4261) );
  MUX21L U3358 ( .A(n4262), .B(n4261), .S(n3197), .Z(n4263) );
  ND2I U3359 ( .A(n3141), .B(n4263), .Z(n4268) );
  MUX21L U3360 ( .A(\gpr[16][26] ), .B(\gpr[17][26] ), .S(n3164), .Z(n4265) );
  MUX21L U3361 ( .A(\gpr[18][26] ), .B(\gpr[19][26] ), .S(n3165), .Z(n4264) );
  MUX21L U3362 ( .A(n4265), .B(n4264), .S(n3197), .Z(n4266) );
  ND2I U3363 ( .A(n3144), .B(n4266), .Z(n4267) );
  ND2I U3364 ( .A(n4268), .B(n4267), .Z(n4269) );
  NR2I U3365 ( .A(n4270), .B(n4269), .Z(n4275) );
  MUX21L U3366 ( .A(\gpr[8][26] ), .B(\gpr[9][26] ), .S(n3165), .Z(n4272) );
  MUX21L U3367 ( .A(\gpr[10][26] ), .B(\gpr[11][26] ), .S(n3166), .Z(n4271) );
  MUX21L U3368 ( .A(n4272), .B(n4271), .S(n3197), .Z(n4273) );
  ND2I U3369 ( .A(n3146), .B(n4273), .Z(n4274) );
  MUX21L U3370 ( .A(n1172), .B(n109), .S(n3166), .Z(n4278) );
  MUX21L U3371 ( .A(n1274), .B(n1305), .S(n3165), .Z(n4277) );
  MUX21L U3372 ( .A(n4278), .B(n4277), .S(n3197), .Z(n4279) );
  ND2I U3373 ( .A(n4279), .B(n3211), .Z(n4280) );
  NR2I U3374 ( .A(n2065), .B(n4280), .Z(n4315) );
  ND2I U3375 ( .A(\gpr[1][27] ), .B(n3180), .Z(n4282) );
  MUX21L U3376 ( .A(\gpr[2][27] ), .B(\gpr[3][27] ), .S(n3166), .Z(n4281) );
  MUX21L U3377 ( .A(n4282), .B(n4281), .S(n3197), .Z(n4283) );
  NR2I U3378 ( .A(n4283), .B(n3211), .Z(n4284) );
  ND2I U3379 ( .A(n4284), .B(n2058), .Z(n4313) );
  MUX21L U3380 ( .A(\gpr[20][27] ), .B(\gpr[21][27] ), .S(n3164), .Z(n4286) );
  MUX21L U3381 ( .A(\gpr[22][27] ), .B(\gpr[23][27] ), .S(n3165), .Z(n4285) );
  MUX21L U3382 ( .A(n4286), .B(n4285), .S(n3197), .Z(n4287) );
  ND2I U3383 ( .A(n2097), .B(n4287), .Z(n4296) );
  MUX21L U3384 ( .A(\gpr[24][27] ), .B(\gpr[25][27] ), .S(n3164), .Z(n4289) );
  MUX21L U3385 ( .A(\gpr[26][27] ), .B(\gpr[27][27] ), .S(n3165), .Z(n4288) );
  MUX21L U3386 ( .A(n4289), .B(n4288), .S(n3197), .Z(n4290) );
  ND2I U3387 ( .A(n2074), .B(n4290), .Z(n4295) );
  MUX21L U3388 ( .A(\gpr[28][27] ), .B(\gpr[29][27] ), .S(n3164), .Z(n4292) );
  MUX21L U3389 ( .A(\gpr[30][27] ), .B(\gpr[31][27] ), .S(n3165), .Z(n4291) );
  MUX21L U3390 ( .A(n4292), .B(n4291), .S(n3197), .Z(n4293) );
  ND2I U3391 ( .A(n3135), .B(n4293), .Z(n4294) );
  MUX21L U3392 ( .A(\gpr[12][27] ), .B(\gpr[13][27] ), .S(n3166), .Z(n4298) );
  MUX21L U3393 ( .A(\gpr[14][27] ), .B(\gpr[15][27] ), .S(n3165), .Z(n4297) );
  MUX21L U3394 ( .A(n4298), .B(n4297), .S(n3197), .Z(n4299) );
  ND2I U3395 ( .A(n3141), .B(n4299), .Z(n4304) );
  MUX21L U3396 ( .A(\gpr[16][27] ), .B(\gpr[17][27] ), .S(n3166), .Z(n4301) );
  MUX21L U3397 ( .A(\gpr[18][27] ), .B(\gpr[19][27] ), .S(n3165), .Z(n4300) );
  MUX21L U3398 ( .A(n4301), .B(n4300), .S(n3196), .Z(n4302) );
  ND2I U3399 ( .A(n3144), .B(n4302), .Z(n4303) );
  ND2I U3400 ( .A(n4304), .B(n4303), .Z(n4305) );
  NR2I U3401 ( .A(n4306), .B(n4305), .Z(n4311) );
  MUX21L U3402 ( .A(\gpr[8][27] ), .B(\gpr[9][27] ), .S(n3165), .Z(n4308) );
  MUX21L U3403 ( .A(\gpr[10][27] ), .B(\gpr[11][27] ), .S(n3165), .Z(n4307) );
  MUX21L U3404 ( .A(n4308), .B(n4307), .S(n3196), .Z(n4309) );
  ND2I U3405 ( .A(n3146), .B(n4309), .Z(n4310) );
  ND2I U3406 ( .A(n4311), .B(n4310), .Z(n4312) );
  ND2I U3407 ( .A(n4313), .B(n4312), .Z(n4314) );
  NR2I U3408 ( .A(n4315), .B(n4314), .Z(rd_data1[27]) );
  MUX21L U3409 ( .A(n1173), .B(n110), .S(n3163), .Z(n4317) );
  MUX21L U3410 ( .A(n1275), .B(n1306), .S(n3163), .Z(n4316) );
  MUX21L U3411 ( .A(n4317), .B(n4316), .S(n3196), .Z(n4318) );
  ND2I U3412 ( .A(n4318), .B(n3211), .Z(n4319) );
  NR2I U3413 ( .A(n2061), .B(n4319), .Z(n4354) );
  ND2I U3414 ( .A(\gpr[1][28] ), .B(n3178), .Z(n4321) );
  MUX21L U3415 ( .A(\gpr[2][28] ), .B(\gpr[3][28] ), .S(n3163), .Z(n4320) );
  MUX21L U3416 ( .A(n4321), .B(n4320), .S(n3196), .Z(n4322) );
  NR2I U3417 ( .A(n4322), .B(n3209), .Z(n4323) );
  ND2I U3418 ( .A(n4323), .B(n2064), .Z(n4352) );
  MUX21L U3419 ( .A(\gpr[20][28] ), .B(\gpr[21][28] ), .S(n3163), .Z(n4325) );
  MUX21L U3420 ( .A(\gpr[22][28] ), .B(\gpr[23][28] ), .S(n3163), .Z(n4324) );
  MUX21L U3421 ( .A(n4325), .B(n4324), .S(n3196), .Z(n4326) );
  ND2I U3422 ( .A(n2099), .B(n4326), .Z(n4335) );
  MUX21L U3423 ( .A(\gpr[24][28] ), .B(\gpr[25][28] ), .S(n3163), .Z(n4328) );
  MUX21L U3424 ( .A(\gpr[26][28] ), .B(\gpr[27][28] ), .S(n3163), .Z(n4327) );
  MUX21L U3425 ( .A(n4328), .B(n4327), .S(n3196), .Z(n4329) );
  ND2I U3426 ( .A(n2077), .B(n4329), .Z(n4334) );
  MUX21L U3427 ( .A(\gpr[28][28] ), .B(\gpr[29][28] ), .S(n3163), .Z(n4331) );
  MUX21L U3428 ( .A(\gpr[30][28] ), .B(\gpr[31][28] ), .S(n3163), .Z(n4330) );
  MUX21L U3429 ( .A(n4331), .B(n4330), .S(n3196), .Z(n4332) );
  ND2I U3430 ( .A(n3137), .B(n4332), .Z(n4333) );
  MUX21L U3431 ( .A(\gpr[12][28] ), .B(\gpr[13][28] ), .S(n3163), .Z(n4337) );
  MUX21L U3432 ( .A(\gpr[14][28] ), .B(\gpr[15][28] ), .S(n3163), .Z(n4336) );
  MUX21L U3433 ( .A(n4337), .B(n4336), .S(n3196), .Z(n4338) );
  ND2I U3434 ( .A(n3141), .B(n4338), .Z(n4343) );
  MUX21L U3435 ( .A(\gpr[16][28] ), .B(\gpr[17][28] ), .S(n3163), .Z(n4340) );
  MUX21L U3436 ( .A(\gpr[18][28] ), .B(\gpr[19][28] ), .S(n3163), .Z(n4339) );
  MUX21L U3437 ( .A(n4340), .B(n4339), .S(n3196), .Z(n4341) );
  ND2I U3438 ( .A(n3144), .B(n4341), .Z(n4342) );
  ND2I U3439 ( .A(n4343), .B(n4342), .Z(n4344) );
  NR2I U3440 ( .A(n4345), .B(n4344), .Z(n4350) );
  MUX21L U3441 ( .A(\gpr[8][28] ), .B(\gpr[9][28] ), .S(n3163), .Z(n4347) );
  MUX21L U3442 ( .A(\gpr[10][28] ), .B(\gpr[11][28] ), .S(n2068), .Z(n4346) );
  MUX21L U3443 ( .A(n4347), .B(n4346), .S(n3196), .Z(n4348) );
  ND2I U3444 ( .A(n3146), .B(n4348), .Z(n4349) );
  ND2I U3445 ( .A(n4350), .B(n4349), .Z(n4351) );
  ND2I U3446 ( .A(n4352), .B(n4351), .Z(n4353) );
  NR2I U3447 ( .A(n4354), .B(n4353), .Z(rd_data1[28]) );
  MUX21L U3448 ( .A(n1174), .B(n111), .S(n2068), .Z(n4356) );
  MUX21L U3449 ( .A(n1276), .B(n1307), .S(n2068), .Z(n4355) );
  MUX21L U3450 ( .A(n4356), .B(n4355), .S(n3196), .Z(n4357) );
  ND2I U3451 ( .A(n4357), .B(n3208), .Z(n4358) );
  NR2I U3452 ( .A(n2059), .B(n4358), .Z(n4393) );
  ND2I U3453 ( .A(\gpr[1][29] ), .B(n3168), .Z(n4360) );
  MUX21L U3454 ( .A(\gpr[2][29] ), .B(\gpr[3][29] ), .S(n2068), .Z(n4359) );
  MUX21L U3455 ( .A(n4360), .B(n4359), .S(n3196), .Z(n4361) );
  NR2I U3456 ( .A(n4361), .B(n3208), .Z(n4362) );
  ND2I U3457 ( .A(n4362), .B(n2066), .Z(n4391) );
  MUX21L U3458 ( .A(\gpr[20][29] ), .B(\gpr[21][29] ), .S(n2101), .Z(n4364) );
  MUX21L U3459 ( .A(\gpr[22][29] ), .B(\gpr[23][29] ), .S(n2101), .Z(n4363) );
  ND2I U3460 ( .A(n2093), .B(n4365), .Z(n4374) );
  MUX21L U3461 ( .A(\gpr[24][29] ), .B(\gpr[25][29] ), .S(n2101), .Z(n4367) );
  MUX21L U3462 ( .A(\gpr[26][29] ), .B(\gpr[27][29] ), .S(n2101), .Z(n4366) );
  ND2I U3463 ( .A(n2080), .B(n4368), .Z(n4373) );
  MUX21L U3464 ( .A(\gpr[28][29] ), .B(\gpr[29][29] ), .S(n2101), .Z(n4370) );
  MUX21L U3465 ( .A(\gpr[30][29] ), .B(\gpr[31][29] ), .S(n2101), .Z(n4369) );
  ND2I U3466 ( .A(n3137), .B(n4371), .Z(n4372) );
  MUX21L U3467 ( .A(\gpr[12][29] ), .B(\gpr[13][29] ), .S(n2101), .Z(n4376) );
  MUX21L U3468 ( .A(\gpr[14][29] ), .B(\gpr[15][29] ), .S(n2068), .Z(n4375) );
  MUX21L U3469 ( .A(n4376), .B(n4375), .S(n3196), .Z(n4377) );
  ND2I U3470 ( .A(n3141), .B(n4377), .Z(n4382) );
  MUX21L U3471 ( .A(\gpr[16][29] ), .B(\gpr[17][29] ), .S(n2101), .Z(n4379) );
  MUX21L U3472 ( .A(\gpr[18][29] ), .B(\gpr[19][29] ), .S(n2101), .Z(n4378) );
  MUX21L U3473 ( .A(n4379), .B(n4378), .S(n3196), .Z(n4380) );
  ND2I U3474 ( .A(n3144), .B(n4380), .Z(n4381) );
  ND2I U3475 ( .A(n4382), .B(n4381), .Z(n4383) );
  NR2I U3476 ( .A(n4384), .B(n4383), .Z(n4389) );
  MUX21L U3477 ( .A(\gpr[8][29] ), .B(\gpr[9][29] ), .S(n3162), .Z(n4386) );
  MUX21L U3478 ( .A(\gpr[10][29] ), .B(\gpr[11][29] ), .S(n3162), .Z(n4385) );
  MUX21L U3479 ( .A(n4386), .B(n4385), .S(n3196), .Z(n4387) );
  ND2I U3480 ( .A(n3146), .B(n4387), .Z(n4388) );
  ND2I U3481 ( .A(n4389), .B(n4388), .Z(n4390) );
  ND2I U3482 ( .A(n4391), .B(n4390), .Z(n4392) );
  NR2I U3483 ( .A(n4393), .B(n4392), .Z(rd_data1[29]) );
  MUX21L U3484 ( .A(n1175), .B(n112), .S(n3162), .Z(n4395) );
  MUX21L U3485 ( .A(n1277), .B(n1308), .S(n3162), .Z(n4394) );
  MUX21L U3486 ( .A(n4395), .B(n4394), .S(n3196), .Z(n4396) );
  ND2I U3487 ( .A(n4396), .B(n3209), .Z(n4397) );
  NR2I U3488 ( .A(n2063), .B(n4397), .Z(n4432) );
  ND2I U3489 ( .A(\gpr[1][30] ), .B(n3179), .Z(n4399) );
  MUX21L U3490 ( .A(\gpr[2][30] ), .B(\gpr[3][30] ), .S(n3162), .Z(n4398) );
  MUX21L U3491 ( .A(n4399), .B(n4398), .S(n3195), .Z(n4400) );
  NR2I U3492 ( .A(n4400), .B(n3209), .Z(n4401) );
  ND2I U3493 ( .A(n4401), .B(n2062), .Z(n4430) );
  MUX21L U3494 ( .A(\gpr[20][30] ), .B(\gpr[21][30] ), .S(n3162), .Z(n4403) );
  MUX21L U3495 ( .A(\gpr[22][30] ), .B(\gpr[23][30] ), .S(n3162), .Z(n4402) );
  ND2I U3496 ( .A(n2096), .B(n4404), .Z(n4413) );
  MUX21L U3497 ( .A(\gpr[24][30] ), .B(\gpr[25][30] ), .S(n3162), .Z(n4406) );
  MUX21L U3498 ( .A(\gpr[26][30] ), .B(\gpr[27][30] ), .S(n3162), .Z(n4405) );
  MUX21L U3499 ( .A(n4406), .B(n4405), .S(n3195), .Z(n4407) );
  ND2I U3500 ( .A(n2074), .B(n4407), .Z(n4412) );
  MUX21L U3501 ( .A(\gpr[28][30] ), .B(\gpr[29][30] ), .S(n3162), .Z(n4409) );
  MUX21L U3502 ( .A(\gpr[30][30] ), .B(\gpr[31][30] ), .S(n3162), .Z(n4408) );
  MUX21L U3503 ( .A(n4409), .B(n4408), .S(n3195), .Z(n4410) );
  ND2I U3504 ( .A(n3138), .B(n4410), .Z(n4411) );
  MUX21L U3505 ( .A(\gpr[12][30] ), .B(\gpr[13][30] ), .S(n3162), .Z(n4415) );
  MUX21L U3506 ( .A(\gpr[14][30] ), .B(\gpr[15][30] ), .S(n3162), .Z(n4414) );
  MUX21L U3507 ( .A(n4415), .B(n4414), .S(n3195), .Z(n4416) );
  ND2I U3508 ( .A(n3140), .B(n4416), .Z(n4421) );
  MUX21L U3509 ( .A(\gpr[16][30] ), .B(\gpr[17][30] ), .S(n3162), .Z(n4418) );
  MUX21L U3510 ( .A(\gpr[18][30] ), .B(\gpr[19][30] ), .S(n3161), .Z(n4417) );
  MUX21L U3511 ( .A(n4418), .B(n4417), .S(n3195), .Z(n4419) );
  ND2I U3512 ( .A(n3143), .B(n4419), .Z(n4420) );
  ND2I U3513 ( .A(n4421), .B(n4420), .Z(n4422) );
  NR2I U3514 ( .A(n4423), .B(n4422), .Z(n4428) );
  MUX21L U3515 ( .A(\gpr[8][30] ), .B(\gpr[9][30] ), .S(n3161), .Z(n4425) );
  MUX21L U3516 ( .A(\gpr[10][30] ), .B(\gpr[11][30] ), .S(n3161), .Z(n4424) );
  MUX21L U3517 ( .A(n4425), .B(n4424), .S(n3195), .Z(n4426) );
  ND2I U3518 ( .A(n3146), .B(n4426), .Z(n4427) );
  ND2I U3519 ( .A(n4428), .B(n4427), .Z(n4429) );
  ND2I U3520 ( .A(n4430), .B(n4429), .Z(n4431) );
  NR2I U3521 ( .A(n4432), .B(n4431), .Z(rd_data1[30]) );
  MUX21L U3522 ( .A(n1176), .B(n113), .S(n3161), .Z(n4434) );
  MUX21L U3523 ( .A(n1278), .B(n1309), .S(n3161), .Z(n4433) );
  MUX21L U3524 ( .A(n4434), .B(n4433), .S(n3195), .Z(n4435) );
  ND2I U3525 ( .A(n4435), .B(n3208), .Z(n4436) );
  NR2I U3526 ( .A(n2065), .B(n4436), .Z(n4475) );
  ND2I U3527 ( .A(n2040), .B(\gpr[1][31] ), .Z(n4438) );
  MUX21L U3528 ( .A(\gpr[2][31] ), .B(\gpr[3][31] ), .S(n3161), .Z(n4437) );
  MUX21L U3529 ( .A(n4438), .B(n4437), .S(n3195), .Z(n4439) );
  NR2I U3530 ( .A(n4439), .B(n3208), .Z(n4440) );
  ND2I U3531 ( .A(n4440), .B(n2056), .Z(n4473) );
  MUX21L U3532 ( .A(\gpr[20][31] ), .B(\gpr[21][31] ), .S(n3161), .Z(n4442) );
  MUX21L U3533 ( .A(\gpr[22][31] ), .B(\gpr[23][31] ), .S(n3161), .Z(n4441) );
  MUX21L U3534 ( .A(n4442), .B(n4441), .S(n3195), .Z(n4443) );
  ND2I U3535 ( .A(n2094), .B(n4443), .Z(n4454) );
  MUX21L U3536 ( .A(\gpr[24][31] ), .B(\gpr[25][31] ), .S(n3161), .Z(n4445) );
  MUX21L U3537 ( .A(\gpr[26][31] ), .B(\gpr[27][31] ), .S(n3161), .Z(n4444) );
  MUX21L U3538 ( .A(n4445), .B(n4444), .S(n3195), .Z(n4446) );
  ND2I U3539 ( .A(n2075), .B(n4446), .Z(n4453) );
  MUX21L U3540 ( .A(\gpr[28][31] ), .B(\gpr[29][31] ), .S(n3161), .Z(n4449) );
  MUX21L U3541 ( .A(\gpr[30][31] ), .B(\gpr[31][31] ), .S(n3161), .Z(n4448) );
  MUX21L U3542 ( .A(n4449), .B(n4448), .S(n3195), .Z(n4450) );
  ND2I U3543 ( .A(n3135), .B(n4450), .Z(n4452) );
  MUX21L U3544 ( .A(\gpr[12][31] ), .B(\gpr[13][31] ), .S(n3161), .Z(n4457) );
  MUX21L U3545 ( .A(\gpr[14][31] ), .B(\gpr[15][31] ), .S(n3161), .Z(n4456) );
  MUX21L U3546 ( .A(n4457), .B(n4456), .S(n3195), .Z(n4458) );
  ND2I U3547 ( .A(n3140), .B(n4458), .Z(n4464) );
  MUX21L U3548 ( .A(\gpr[16][31] ), .B(\gpr[17][31] ), .S(n3159), .Z(n4461) );
  MUX21L U3549 ( .A(\gpr[18][31] ), .B(\gpr[19][31] ), .S(n3174), .Z(n4460) );
  MUX21L U3550 ( .A(n4461), .B(n4460), .S(n3198), .Z(n4462) );
  ND2I U3551 ( .A(n3143), .B(n4462), .Z(n4463) );
  ND2I U3552 ( .A(n4464), .B(n4463), .Z(n4465) );
  NR2I U3553 ( .A(n4466), .B(n4465), .Z(n4471) );
  MUX21L U3554 ( .A(\gpr[8][31] ), .B(\gpr[9][31] ), .S(n3165), .Z(n4468) );
  MUX21L U3555 ( .A(\gpr[10][31] ), .B(\gpr[11][31] ), .S(n3166), .Z(n4467) );
  MUX21L U3556 ( .A(n4468), .B(n4467), .S(n3191), .Z(n4469) );
  ND2I U3557 ( .A(n3146), .B(n4469), .Z(n4470) );
  ND2I U3558 ( .A(n4471), .B(n4470), .Z(n4472) );
  ND2I U3559 ( .A(n4473), .B(n4472), .Z(n4474) );
  NR2I U3560 ( .A(n4475), .B(n4474), .Z(rd_data1[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_6 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4;

  B5IP U1 ( .A(n4), .Z(n2) );
  IVI U2 ( .A(n4), .Z(n1) );
  IVI U3 ( .A(n4), .Z(n3) );
  IVI U4 ( .A(sel), .Z(n4) );
  MUX21H U5 ( .A(ip0[0]), .B(ip1[0]), .S(n3), .Z(out[0]) );
  MUX21H U6 ( .A(ip0[1]), .B(ip1[1]), .S(n3), .Z(out[1]) );
  MUX21H U7 ( .A(ip0[2]), .B(ip1[2]), .S(n3), .Z(out[2]) );
  MUX21H U8 ( .A(ip0[3]), .B(ip1[3]), .S(n3), .Z(out[3]) );
  MUX21H U9 ( .A(ip0[4]), .B(ip1[4]), .S(n2), .Z(out[4]) );
  MUX21H U10 ( .A(ip0[5]), .B(ip1[5]), .S(n2), .Z(out[5]) );
  MUX21H U11 ( .A(ip0[6]), .B(ip1[6]), .S(n2), .Z(out[6]) );
  MUX21H U12 ( .A(ip0[7]), .B(ip1[7]), .S(n2), .Z(out[7]) );
  MUX21H U13 ( .A(ip0[8]), .B(ip1[8]), .S(n2), .Z(out[8]) );
  MUX21H U14 ( .A(ip0[9]), .B(ip1[9]), .S(n2), .Z(out[9]) );
  MUX21H U15 ( .A(ip0[10]), .B(ip1[10]), .S(n2), .Z(out[10]) );
  MUX21H U16 ( .A(ip0[11]), .B(ip1[11]), .S(n2), .Z(out[11]) );
  MUX21H U17 ( .A(ip0[12]), .B(ip1[12]), .S(n2), .Z(out[12]) );
  MUX21H U18 ( .A(ip0[13]), .B(ip1[13]), .S(n2), .Z(out[13]) );
  MUX21H U19 ( .A(ip0[14]), .B(ip1[14]), .S(n2), .Z(out[14]) );
  MUX21H U20 ( .A(ip0[15]), .B(ip1[15]), .S(n2), .Z(out[15]) );
  MUX21H U21 ( .A(ip0[16]), .B(ip1[16]), .S(n2), .Z(out[16]) );
  MUX21H U22 ( .A(ip0[17]), .B(ip1[17]), .S(n2), .Z(out[17]) );
  MUX21H U23 ( .A(ip0[18]), .B(ip1[18]), .S(n1), .Z(out[18]) );
  MUX21H U24 ( .A(ip0[19]), .B(ip1[19]), .S(n1), .Z(out[19]) );
  MUX21H U25 ( .A(ip0[20]), .B(ip1[20]), .S(n1), .Z(out[20]) );
  MUX21H U26 ( .A(ip0[21]), .B(ip1[21]), .S(n1), .Z(out[21]) );
  MUX21H U27 ( .A(ip0[22]), .B(ip1[22]), .S(n1), .Z(out[22]) );
  MUX21H U28 ( .A(ip0[23]), .B(ip1[23]), .S(n1), .Z(out[23]) );
  MUX21H U29 ( .A(ip0[24]), .B(ip1[24]), .S(n1), .Z(out[24]) );
  MUX21H U30 ( .A(ip0[25]), .B(ip1[25]), .S(n1), .Z(out[25]) );
  MUX21H U31 ( .A(ip0[26]), .B(ip1[26]), .S(n1), .Z(out[26]) );
  MUX21H U32 ( .A(ip0[27]), .B(ip1[27]), .S(n1), .Z(out[27]) );
  MUX21H U33 ( .A(ip0[28]), .B(ip1[28]), .S(n1), .Z(out[28]) );
  MUX21H U34 ( .A(ip0[29]), .B(ip1[29]), .S(n1), .Z(out[29]) );
  MUX21H U35 ( .A(ip0[30]), .B(ip1[30]), .S(n1), .Z(out[30]) );
  MUX21H U36 ( .A(ip0[31]), .B(ip1[31]), .S(n1), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_5 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4;

  IVAP U1 ( .A(n4), .Z(n2) );
  IVAP U2 ( .A(n4), .Z(n1) );
  IVI U3 ( .A(n4), .Z(n3) );
  IVI U4 ( .A(sel), .Z(n4) );
  MUX21H U5 ( .A(ip0[0]), .B(ip1[0]), .S(n3), .Z(out[0]) );
  MUX21H U6 ( .A(ip0[1]), .B(ip1[1]), .S(n3), .Z(out[1]) );
  MUX21H U7 ( .A(ip0[2]), .B(ip1[2]), .S(n3), .Z(out[2]) );
  MUX21H U8 ( .A(ip0[3]), .B(ip1[3]), .S(n3), .Z(out[3]) );
  MUX21H U9 ( .A(ip0[4]), .B(ip1[4]), .S(n2), .Z(out[4]) );
  MUX21H U10 ( .A(ip0[5]), .B(ip1[5]), .S(n2), .Z(out[5]) );
  MUX21H U11 ( .A(ip0[6]), .B(ip1[6]), .S(n2), .Z(out[6]) );
  MUX21H U12 ( .A(ip0[7]), .B(ip1[7]), .S(n2), .Z(out[7]) );
  MUX21H U13 ( .A(ip0[8]), .B(ip1[8]), .S(n2), .Z(out[8]) );
  MUX21H U14 ( .A(ip0[9]), .B(ip1[9]), .S(n2), .Z(out[9]) );
  MUX21H U15 ( .A(ip0[10]), .B(ip1[10]), .S(n2), .Z(out[10]) );
  MUX21H U16 ( .A(ip0[11]), .B(ip1[11]), .S(n2), .Z(out[11]) );
  MUX21H U17 ( .A(ip0[12]), .B(ip1[12]), .S(n2), .Z(out[12]) );
  MUX21H U18 ( .A(ip0[13]), .B(ip1[13]), .S(n2), .Z(out[13]) );
  MUX21H U19 ( .A(ip0[14]), .B(ip1[14]), .S(n2), .Z(out[14]) );
  MUX21H U20 ( .A(ip0[15]), .B(ip1[15]), .S(n2), .Z(out[15]) );
  MUX21H U21 ( .A(ip0[16]), .B(ip1[16]), .S(n2), .Z(out[16]) );
  MUX21H U22 ( .A(ip0[17]), .B(ip1[17]), .S(n2), .Z(out[17]) );
  MUX21H U23 ( .A(ip0[18]), .B(ip1[18]), .S(n1), .Z(out[18]) );
  MUX21H U24 ( .A(ip0[19]), .B(ip1[19]), .S(n1), .Z(out[19]) );
  MUX21H U25 ( .A(ip0[20]), .B(ip1[20]), .S(n1), .Z(out[20]) );
  MUX21H U26 ( .A(ip0[21]), .B(ip1[21]), .S(n1), .Z(out[21]) );
  MUX21H U27 ( .A(ip0[22]), .B(ip1[22]), .S(n1), .Z(out[22]) );
  MUX21H U28 ( .A(ip0[23]), .B(ip1[23]), .S(n1), .Z(out[23]) );
  MUX21H U29 ( .A(ip0[24]), .B(ip1[24]), .S(n1), .Z(out[24]) );
  MUX21H U30 ( .A(ip0[25]), .B(ip1[25]), .S(n1), .Z(out[25]) );
  MUX21H U31 ( .A(ip0[26]), .B(ip1[26]), .S(n1), .Z(out[26]) );
  MUX21H U32 ( .A(ip0[27]), .B(ip1[27]), .S(n1), .Z(out[27]) );
  MUX21H U33 ( .A(ip0[28]), .B(ip1[28]), .S(n1), .Z(out[28]) );
  MUX21H U34 ( .A(ip0[29]), .B(ip1[29]), .S(n1), .Z(out[29]) );
  MUX21H U35 ( .A(ip0[30]), .B(ip1[30]), .S(n1), .Z(out[30]) );
  MUX21H U36 ( .A(ip0[31]), .B(ip1[31]), .S(n1), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_4 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33;

  IVI U1 ( .A(n9), .Z(n1) );
  EON1P U2 ( .A(n21), .B(n22), .C(ip1[1]), .D(n8), .Z(out[1]) );
  IVI U3 ( .A(n9), .Z(n29) );
  EON1 U4 ( .A(n17), .B(n22), .C(ip1[2]), .D(n8), .Z(out[2]) );
  IVI U5 ( .A(ip1[9]), .Z(n26) );
  IVI U6 ( .A(ip1[17]), .Z(n24) );
  IVI U7 ( .A(ip0[17]), .Z(n23) );
  IVI U8 ( .A(ip1[16]), .Z(n28) );
  IVI U9 ( .A(ip1[12]), .Z(n11) );
  IVI U10 ( .A(ip1[10]), .Z(n5) );
  IVI U11 ( .A(ip0[20]), .Z(n14) );
  IVI U12 ( .A(ip1[20]), .Z(n15) );
  IVI U13 ( .A(ip1[18]), .Z(n13) );
  IVI U14 ( .A(ip0[18]), .Z(n12) );
  IVI U15 ( .A(ip0[9]), .Z(n25) );
  IVI U16 ( .A(ip1[8]), .Z(n7) );
  IVI U17 ( .A(ip1[3]), .Z(n19) );
  IVI U18 ( .A(ip0[3]), .Z(n18) );
  IVI U19 ( .A(ip0[1]), .Z(n21) );
  IVI U20 ( .A(ip0[16]), .Z(n27) );
  IVI U21 ( .A(ip0[12]), .Z(n10) );
  IVI U22 ( .A(ip0[10]), .Z(n4) );
  IVI U23 ( .A(ip0[2]), .Z(n17) );
  IVI U24 ( .A(n9), .Z(n2) );
  AO2 U25 ( .A(ip0[0]), .B(n31), .C(ip1[0]), .D(n8), .Z(n32) );
  AO2 U26 ( .A(ip0[4]), .B(n31), .C(ip1[4]), .D(n8), .Z(n33) );
  IVI U27 ( .A(n31), .Z(n3) );
  MUX21L U28 ( .A(n4), .B(n5), .S(n1), .Z(out[10]) );
  EON1 U29 ( .A(n7), .B(n31), .C(ip0[8]), .D(n31), .Z(out[8]) );
  IVDAP U30 ( .A(sel), .Y(n31), .Z(n22) );
  B4IP U31 ( .A(n9), .Z(n30) );
  B3IP U32 ( .A(sel), .Z1(n9), .Z2(n8) );
  MUX21L U33 ( .A(n10), .B(n11), .S(n1), .Z(out[12]) );
  MUX21L U34 ( .A(n12), .B(n13), .S(n29), .Z(out[18]) );
  MUX21L U35 ( .A(n14), .B(n15), .S(n2), .Z(out[20]) );
  MUX21L U36 ( .A(n27), .B(n28), .S(n8), .Z(out[16]) );
  MUX21L U37 ( .A(n18), .B(n19), .S(n2), .Z(out[3]) );
  MUX21L U38 ( .A(n23), .B(n24), .S(n8), .Z(out[17]) );
  MUX21L U39 ( .A(n25), .B(n26), .S(n30), .Z(out[9]) );
  IVI U40 ( .A(n32), .Z(out[0]) );
  IVI U41 ( .A(n33), .Z(out[4]) );
  MUX21H U42 ( .A(ip0[5]), .B(ip1[5]), .S(n8), .Z(out[5]) );
  MUX21H U43 ( .A(ip0[6]), .B(ip1[6]), .S(n3), .Z(out[6]) );
  MUX21H U44 ( .A(ip0[7]), .B(ip1[7]), .S(n2), .Z(out[7]) );
  MUX21H U45 ( .A(ip0[11]), .B(ip1[11]), .S(n3), .Z(out[11]) );
  MUX21H U46 ( .A(ip0[13]), .B(ip1[13]), .S(n30), .Z(out[13]) );
  MUX21H U47 ( .A(ip0[14]), .B(ip1[14]), .S(n29), .Z(out[14]) );
  MUX21H U48 ( .A(ip0[15]), .B(ip1[15]), .S(n30), .Z(out[15]) );
  MUX21H U49 ( .A(ip0[19]), .B(ip1[19]), .S(n29), .Z(out[19]) );
  MUX21H U50 ( .A(ip0[21]), .B(ip1[21]), .S(n30), .Z(out[21]) );
  MUX21H U51 ( .A(ip0[22]), .B(ip1[22]), .S(n8), .Z(out[22]) );
  MUX21H U52 ( .A(ip0[23]), .B(ip1[23]), .S(n30), .Z(out[23]) );
  MUX21H U53 ( .A(ip0[24]), .B(ip1[24]), .S(n30), .Z(out[24]) );
  MUX21H U54 ( .A(ip0[25]), .B(ip1[25]), .S(n2), .Z(out[25]) );
  MUX21H U55 ( .A(ip0[26]), .B(ip1[26]), .S(n30), .Z(out[26]) );
  MUX21H U56 ( .A(ip0[27]), .B(ip1[27]), .S(n30), .Z(out[27]) );
  MUX21H U57 ( .A(ip0[28]), .B(ip1[28]), .S(n22), .Z(out[28]) );
  MUX21H U58 ( .A(ip0[29]), .B(ip1[29]), .S(n22), .Z(out[29]) );
  MUX21H U59 ( .A(ip0[30]), .B(ip1[30]), .S(n29), .Z(out[30]) );
  MUX21H U60 ( .A(ip0[31]), .B(ip1[31]), .S(n1), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_3 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30;

  AO2P U1 ( .A(ip0[4]), .B(n14), .C(ip1[4]), .D(n23), .Z(n30) );
  IVI U2 ( .A(n25), .Z(n1) );
  AO2P U3 ( .A(ip0[2]), .B(n14), .C(ip1[2]), .D(n23), .Z(n29) );
  IVI U4 ( .A(ip0[3]), .Z(n17) );
  IVI U5 ( .A(ip1[3]), .Z(n18) );
  IVI U6 ( .A(ip1[1]), .Z(n16) );
  IVI U7 ( .A(ip0[1]), .Z(n8) );
  IVI U8 ( .A(ip1[15]), .Z(n4) );
  IVI U9 ( .A(ip0[15]), .Z(n3) );
  IVI U10 ( .A(ip1[13]), .Z(n13) );
  IVI U11 ( .A(ip0[13]), .Z(n12) );
  IVI U12 ( .A(ip1[12]), .Z(n7) );
  IVI U13 ( .A(ip0[12]), .Z(n6) );
  IVI U14 ( .A(n25), .Z(n2) );
  MUX21H U15 ( .A(ip1[7]), .B(ip0[7]), .S(n14), .Z(out[7]) );
  MUX21L U16 ( .A(n3), .B(n4), .S(n19), .Z(out[15]) );
  IVI U17 ( .A(n26), .Z(n5) );
  IVI U18 ( .A(n27), .Z(n10) );
  MUX21L U19 ( .A(n6), .B(n7), .S(n10), .Z(out[12]) );
  AO4P U20 ( .A(n16), .B(n26), .C(n8), .D(n2), .Z(out[1]) );
  IVI U21 ( .A(n25), .Z(n20) );
  IVI U22 ( .A(n26), .Z(n9) );
  IVI U23 ( .A(n22), .Z(n11) );
  B3IP U24 ( .A(n11), .Z1(n14), .Z2(n19) );
  IVI U25 ( .A(n22), .Z(n21) );
  MUX21L U26 ( .A(n12), .B(n13), .S(n19), .Z(out[13]) );
  MUX21H U27 ( .A(ip1[20]), .B(ip0[20]), .S(n14), .Z(out[20]) );
  MUX21L U28 ( .A(n17), .B(n18), .S(n24), .Z(out[3]) );
  IVI U29 ( .A(n25), .Z(n24) );
  IVI U30 ( .A(n25), .Z(n23) );
  IVI U31 ( .A(sel), .Z(n25) );
  AO2P U32 ( .A(ip1[0]), .B(n1), .C(ip0[0]), .D(n27), .Z(n28) );
  IVI U33 ( .A(sel), .Z(n22) );
  IVI U34 ( .A(n21), .Z(n26) );
  IVI U35 ( .A(n21), .Z(n27) );
  IVI U36 ( .A(n28), .Z(out[0]) );
  IVI U37 ( .A(n29), .Z(out[2]) );
  IVI U38 ( .A(n30), .Z(out[4]) );
  MUX21H U39 ( .A(ip0[5]), .B(ip1[5]), .S(n23), .Z(out[5]) );
  MUX21H U40 ( .A(ip0[6]), .B(ip1[6]), .S(n20), .Z(out[6]) );
  MUX21H U41 ( .A(ip0[8]), .B(ip1[8]), .S(n2), .Z(out[8]) );
  MUX21H U42 ( .A(ip0[9]), .B(ip1[9]), .S(n9), .Z(out[9]) );
  MUX21H U43 ( .A(ip0[10]), .B(ip1[10]), .S(n23), .Z(out[10]) );
  MUX21H U44 ( .A(ip0[11]), .B(ip1[11]), .S(n5), .Z(out[11]) );
  MUX21H U45 ( .A(ip0[14]), .B(ip1[14]), .S(n2), .Z(out[14]) );
  MUX21H U46 ( .A(ip0[16]), .B(ip1[16]), .S(n20), .Z(out[16]) );
  MUX21H U47 ( .A(ip0[17]), .B(ip1[17]), .S(n19), .Z(out[17]) );
  MUX21H U48 ( .A(ip0[18]), .B(ip1[18]), .S(n19), .Z(out[18]) );
  MUX21H U49 ( .A(ip0[19]), .B(ip1[19]), .S(n24), .Z(out[19]) );
  MUX21H U50 ( .A(ip0[21]), .B(ip1[21]), .S(n19), .Z(out[21]) );
  MUX21H U51 ( .A(ip0[22]), .B(ip1[22]), .S(n9), .Z(out[22]) );
  MUX21H U52 ( .A(ip0[23]), .B(ip1[23]), .S(n20), .Z(out[23]) );
  MUX21H U53 ( .A(ip0[24]), .B(ip1[24]), .S(n24), .Z(out[24]) );
  MUX21H U54 ( .A(ip0[25]), .B(ip1[25]), .S(n24), .Z(out[25]) );
  MUX21H U55 ( .A(ip0[26]), .B(ip1[26]), .S(n19), .Z(out[26]) );
  MUX21H U56 ( .A(ip0[27]), .B(ip1[27]), .S(n19), .Z(out[27]) );
  MUX21H U57 ( .A(ip0[28]), .B(ip1[28]), .S(n5), .Z(out[28]) );
  MUX21H U58 ( .A(ip0[29]), .B(ip1[29]), .S(n2), .Z(out[29]) );
  MUX21H U59 ( .A(ip0[30]), .B(ip1[30]), .S(n20), .Z(out[30]) );
  MUX21H U60 ( .A(ip0[31]), .B(ip1[31]), .S(n10), .Z(out[31]) );
endmodule


module mux_2x1_DATA_WIDTH32_2 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n5, n6, n8, n9, n10, n11, n14, n15, n17, n18, n19, n20, n21,
         n22, n23, n24, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n37,
         n38, n39, n40, n41, n42, n44, n45, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73;

  B4I U1 ( .A(n61), .Z(out[5]) );
  IVDAP U2 ( .A(n51), .Y(n1), .Z(n2) );
  ND2I U3 ( .A(n26), .B(n27), .Z(out[27]) );
  ND2I U4 ( .A(n37), .B(n38), .Z(out[20]) );
  ND2I U5 ( .A(ip1[7]), .B(n11), .Z(n5) );
  ND2I U6 ( .A(ip0[7]), .B(n54), .Z(n6) );
  ND2I U7 ( .A(n5), .B(n6), .Z(out[7]) );
  ND2I U8 ( .A(ip1[2]), .B(n52), .Z(n8) );
  ND2I U9 ( .A(ip0[2]), .B(n56), .Z(n9) );
  AN2I U10 ( .A(n8), .B(n9), .Z(n59) );
  B4IP U11 ( .A(n59), .Z(out[2]) );
  ND2I U12 ( .A(n44), .B(n45), .Z(out[17]) );
  B3IP U13 ( .A(sel), .Z1(n10), .Z2(n11) );
  ND2I U14 ( .A(n28), .B(n29), .Z(out[3]) );
  ND2I U15 ( .A(n39), .B(n40), .Z(out[28]) );
  B4IP U16 ( .A(n60), .Z(out[4]) );
  ND2I U17 ( .A(ip1[18]), .B(n1), .Z(n14) );
  ND2I U18 ( .A(ip0[18]), .B(n53), .Z(n15) );
  ND2I U19 ( .A(n14), .B(n15), .Z(out[18]) );
  ND2I U20 ( .A(ip1[0]), .B(n52), .Z(n17) );
  ND2I U21 ( .A(ip0[0]), .B(n10), .Z(n18) );
  AN2I U22 ( .A(n17), .B(n18), .Z(n57) );
  B5IP U23 ( .A(n57), .Z(out[0]) );
  IVI U24 ( .A(n64), .Z(out[10]) );
  ND2I U25 ( .A(ip1[1]), .B(n52), .Z(n19) );
  ND2I U26 ( .A(ip0[1]), .B(n56), .Z(n20) );
  AN2I U27 ( .A(n19), .B(n20), .Z(n58) );
  B4IP U28 ( .A(n58), .Z(out[1]) );
  ND2I U29 ( .A(ip1[25]), .B(n11), .Z(n21) );
  ND2I U30 ( .A(ip0[25]), .B(n2), .Z(n22) );
  AN2I U31 ( .A(n21), .B(n22), .Z(n72) );
  B4IP U32 ( .A(n72), .Z(out[25]) );
  ND2I U33 ( .A(ip1[19]), .B(n52), .Z(n23) );
  ND2I U34 ( .A(ip0[19]), .B(n54), .Z(n24) );
  ND2I U35 ( .A(n23), .B(n24), .Z(out[19]) );
  B5I U36 ( .A(n70), .Z(out[22]) );
  ND2I U37 ( .A(ip1[27]), .B(n11), .Z(n26) );
  ND2I U38 ( .A(ip0[27]), .B(n2), .Z(n27) );
  ND2I U39 ( .A(ip1[3]), .B(n11), .Z(n28) );
  ND2I U40 ( .A(ip0[3]), .B(n56), .Z(n29) );
  ND2I U41 ( .A(ip1[4]), .B(n11), .Z(n30) );
  ND2I U42 ( .A(ip0[4]), .B(n53), .Z(n31) );
  AN2I U43 ( .A(n30), .B(n31), .Z(n60) );
  AO2P U44 ( .A(ip1[22]), .B(n11), .C(ip0[22]), .D(n56), .Z(n70) );
  AO2P U45 ( .A(ip1[26]), .B(n52), .C(ip0[26]), .D(n2), .Z(n73) );
  B5I U46 ( .A(n73), .Z(out[26]) );
  ND2I U47 ( .A(ip1[24]), .B(n1), .Z(n32) );
  ND2I U48 ( .A(ip0[24]), .B(n2), .Z(n33) );
  AN2I U49 ( .A(n32), .B(n33), .Z(n71) );
  B4IP U50 ( .A(n71), .Z(out[24]) );
  ND2I U51 ( .A(ip1[6]), .B(n11), .Z(n34) );
  ND2I U52 ( .A(ip0[6]), .B(n53), .Z(n35) );
  ND2I U53 ( .A(n34), .B(n35), .Z(out[6]) );
  ND2I U54 ( .A(ip1[20]), .B(n11), .Z(n37) );
  ND2I U55 ( .A(ip0[20]), .B(n56), .Z(n38) );
  B4I U56 ( .A(n67), .Z(out[13]) );
  ND2I U57 ( .A(ip1[28]), .B(n52), .Z(n39) );
  ND2I U58 ( .A(ip0[28]), .B(n2), .Z(n40) );
  B4IP U59 ( .A(n10), .Z(n52) );
  IVI U60 ( .A(n63), .Z(out[9]) );
  IVI U61 ( .A(n66), .Z(out[12]) );
  ND2I U62 ( .A(ip1[14]), .B(n11), .Z(n41) );
  ND2I U63 ( .A(ip0[14]), .B(n55), .Z(n42) );
  ND2P U64 ( .A(n41), .B(n42), .Z(out[14]) );
  AO2P U65 ( .A(ip1[21]), .B(n52), .C(ip0[21]), .D(n56), .Z(n69) );
  B5I U66 ( .A(n69), .Z(out[21]) );
  AO2P U67 ( .A(ip1[5]), .B(n52), .C(ip0[5]), .D(n53), .Z(n61) );
  AO2P U68 ( .A(ip1[12]), .B(n1), .C(ip0[12]), .D(n53), .Z(n66) );
  ND2I U69 ( .A(ip1[17]), .B(n52), .Z(n44) );
  ND2I U70 ( .A(ip0[17]), .B(n2), .Z(n45) );
  AO2P U71 ( .A(ip1[13]), .B(n52), .C(ip0[13]), .D(n55), .Z(n67) );
  IVI U72 ( .A(n68), .Z(out[16]) );
  AO2P U73 ( .A(ip1[10]), .B(n1), .C(ip0[10]), .D(n53), .Z(n64) );
  ND2I U74 ( .A(ip1[8]), .B(n11), .Z(n47) );
  ND2I U75 ( .A(ip0[8]), .B(n54), .Z(n48) );
  AN2I U76 ( .A(n47), .B(n48), .Z(n62) );
  B4IP U77 ( .A(n62), .Z(out[8]) );
  AO2P U78 ( .A(ip1[16]), .B(n11), .C(ip0[16]), .D(n55), .Z(n68) );
  MUX21LP U79 ( .A(ip1[30]), .B(ip0[30]), .S(n10), .Z(n49) );
  B4IP U80 ( .A(n49), .Z(out[30]) );
  MUX21HP U81 ( .A(ip0[23]), .B(ip1[23]), .S(n52), .Z(out[23]) );
  MUX21HP U82 ( .A(ip0[15]), .B(ip1[15]), .S(n52), .Z(out[15]) );
  MUX21HP U83 ( .A(ip0[31]), .B(ip1[31]), .S(n52), .Z(out[31]) );
  AO2P U84 ( .A(ip1[9]), .B(n11), .C(ip0[9]), .D(n54), .Z(n63) );
  MUX21HP U85 ( .A(ip0[29]), .B(ip1[29]), .S(n11), .Z(out[29]) );
  IVI U86 ( .A(sel), .Z(n51) );
  IVI U87 ( .A(n51), .Z(n50) );
  IVI U88 ( .A(sel), .Z(n53) );
  IVI U89 ( .A(n50), .Z(n54) );
  IVI U90 ( .A(n50), .Z(n55) );
  IVI U91 ( .A(n50), .Z(n56) );
  AO2 U92 ( .A(ip1[11]), .B(n1), .C(ip0[11]), .D(n53), .Z(n65) );
  IVI U93 ( .A(n65), .Z(out[11]) );
endmodule


module mux_2x1_DATA_WIDTH32_1 ( ip1, ip0, sel, out );
  input [31:0] ip1;
  input [31:0] ip0;
  output [31:0] out;
  input sel;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40;

  IVI U1 ( .A(n21), .Z(n1) );
  B5I U2 ( .A(sel), .Z(n17) );
  MUX21H U3 ( .A(ip0[29]), .B(ip1[29]), .S(n16), .Z(out[29]) );
  B3IP U4 ( .A(n15), .Z1(n2), .Z2(n4) );
  B5I U5 ( .A(n14), .Z(n20) );
  IVI U6 ( .A(n17), .Z(n8) );
  IVI U7 ( .A(ip0[0]), .Z(n13) );
  B5IP U8 ( .A(n10), .Z(out[30]) );
  IVI U9 ( .A(n7), .Z(out[19]) );
  AO2P U10 ( .A(ip1[12]), .B(n16), .C(ip0[12]), .D(n20), .Z(n35) );
  AO2P U11 ( .A(ip1[1]), .B(n16), .C(ip0[1]), .D(n18), .Z(n22) );
  ND2I U12 ( .A(n5), .B(n6), .Z(out[24]) );
  AO2P U13 ( .A(ip1[9]), .B(n8), .C(ip0[9]), .D(n2), .Z(n32) );
  AO2P U14 ( .A(ip1[4]), .B(n8), .C(ip0[4]), .D(n19), .Z(n27) );
  ND2I U15 ( .A(ip1[24]), .B(n16), .Z(n5) );
  ND2I U16 ( .A(ip0[24]), .B(n21), .Z(n6) );
  IVI U17 ( .A(n11), .Z(out[22]) );
  MUX21H U18 ( .A(ip0[25]), .B(ip1[25]), .S(n8), .Z(out[25]) );
  AO2P U19 ( .A(ip1[7]), .B(n8), .C(ip0[7]), .D(n2), .Z(n30) );
  AO2P U20 ( .A(ip1[6]), .B(n8), .C(ip0[6]), .D(n19), .Z(n29) );
  IVI U21 ( .A(n9), .Z(out[14]) );
  MUX21L U22 ( .A(ip0[14]), .B(ip1[14]), .S(n16), .Z(n9) );
  MUX21LP U23 ( .A(ip1[19]), .B(ip0[19]), .S(n19), .Z(n7) );
  AO2 U24 ( .A(ip1[5]), .B(n8), .C(ip0[5]), .D(n19), .Z(n28) );
  AO2 U25 ( .A(ip1[10]), .B(n8), .C(ip0[10]), .D(n20), .Z(n33) );
  MUX21HP U26 ( .A(ip0[27]), .B(ip1[27]), .S(n8), .Z(out[27]) );
  MUX21HP U27 ( .A(ip0[26]), .B(ip1[26]), .S(n16), .Z(out[26]) );
  AO2P U28 ( .A(ip1[13]), .B(n16), .C(ip0[13]), .D(n2), .Z(n36) );
  AO2P U29 ( .A(ip1[8]), .B(n16), .C(ip0[8]), .D(n2), .Z(n31) );
  IVI U30 ( .A(n29), .Z(out[6]) );
  MUX21H U31 ( .A(ip0[31]), .B(ip1[31]), .S(n4), .Z(out[31]) );
  AO2P U32 ( .A(ip1[17]), .B(n4), .C(ip0[17]), .D(n2), .Z(n38) );
  MUX21HP U33 ( .A(ip0[28]), .B(ip1[28]), .S(n4), .Z(out[28]) );
  IVI U34 ( .A(n40), .Z(out[20]) );
  IVI U35 ( .A(n28), .Z(out[5]) );
  MUX21LP U36 ( .A(ip0[30]), .B(ip1[30]), .S(n15), .Z(n10) );
  IVI U37 ( .A(n27), .Z(out[4]) );
  IVI U38 ( .A(n37), .Z(out[16]) );
  IVI U39 ( .A(n36), .Z(out[13]) );
  MUX21HP U40 ( .A(ip0[23]), .B(ip1[23]), .S(n16), .Z(out[23]) );
  MUX21LP U41 ( .A(ip0[22]), .B(ip1[22]), .S(n4), .Z(n11) );
  MUX21H U42 ( .A(ip0[15]), .B(ip1[15]), .S(n8), .Z(out[15]) );
  IVI U43 ( .A(n31), .Z(out[8]) );
  AO2P U44 ( .A(ip1[16]), .B(n4), .C(ip0[16]), .D(n2), .Z(n37) );
  IVI U45 ( .A(n35), .Z(out[12]) );
  EO1P U46 ( .A(n13), .B(n20), .C(ip1[0]), .D(n21), .Z(out[0]) );
  MUX21HP U47 ( .A(ip0[21]), .B(ip1[21]), .S(n8), .Z(out[21]) );
  IVI U48 ( .A(n30), .Z(out[7]) );
  AO2P U49 ( .A(ip1[20]), .B(n1), .C(ip0[20]), .D(n21), .Z(n40) );
  IVI U50 ( .A(n17), .Z(n14) );
  IVI U51 ( .A(n17), .Z(n15) );
  IVI U52 ( .A(n17), .Z(n16) );
  IVI U53 ( .A(n14), .Z(n18) );
  IVI U54 ( .A(n14), .Z(n19) );
  IVI U55 ( .A(n14), .Z(n21) );
  IVI U56 ( .A(n22), .Z(out[1]) );
  ND2I U57 ( .A(ip0[2]), .B(n18), .Z(n24) );
  ND2I U58 ( .A(ip1[2]), .B(n8), .Z(n23) );
  ND2I U59 ( .A(n24), .B(n23), .Z(out[2]) );
  ND2I U60 ( .A(ip0[3]), .B(n18), .Z(n26) );
  ND2I U61 ( .A(ip1[3]), .B(n15), .Z(n25) );
  ND2I U62 ( .A(n26), .B(n25), .Z(out[3]) );
  IVI U63 ( .A(n32), .Z(out[9]) );
  IVI U64 ( .A(n33), .Z(out[10]) );
  AO2 U65 ( .A(ip1[11]), .B(n8), .C(ip0[11]), .D(n20), .Z(n34) );
  IVI U66 ( .A(n34), .Z(out[11]) );
  IVI U67 ( .A(n38), .Z(out[17]) );
  AO2 U68 ( .A(ip1[18]), .B(n4), .C(ip0[18]), .D(n21), .Z(n39) );
  IVI U69 ( .A(n39), .Z(out[18]) );
endmodule


module alu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n4, n6, n8, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n26, n27, n28, n29, n30, n31, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n85, n86, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n145, n146, n149, n150,
         n151, n152, n153, n154, n155, n157, n158, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n197, n198, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n216, n217, n222, n223, n224, n225, n226, n228, n229, n230,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n260, n261, n262, n264, n267, n268, n269,
         n270, n271, n272, n273, n274, n277, n279, n280, n281, n384, n385,
         n386, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n450, n451, n452, n453,
         n454, n455, n456, n458, n459;

  EOI U16 ( .A(n26), .B(n17), .Z(n15) );
  EOI U17 ( .A(n17), .B(n27), .Z(n16) );
  ENI U18 ( .A(A[31]), .B(B[31]), .Z(n17) );
  ENI U24 ( .A(n36), .B(n454), .Z(n22) );
  ENI U25 ( .A(n37), .B(n454), .Z(n23) );
  NR2I U28 ( .A(A[30]), .B(B[30]), .Z(n26) );
  ND2I U29 ( .A(A[30]), .B(B[30]), .Z(n27) );
  ENI U41 ( .A(A[29]), .B(B[29]), .Z(n38) );
  NR2I U42 ( .A(A[29]), .B(B[29]), .Z(n39) );
  ND2I U43 ( .A(A[29]), .B(B[29]), .Z(n40) );
  EOI U47 ( .A(n54), .B(n45), .Z(n43) );
  EOI U48 ( .A(n55), .B(n45), .Z(n44) );
  ENI U49 ( .A(A[28]), .B(B[28]), .Z(n45) );
  NR2I U50 ( .A(A[28]), .B(B[28]), .Z(n46) );
  ND2I U51 ( .A(A[28]), .B(B[28]), .Z(n47) );
  EOI U61 ( .A(n407), .B(n60), .Z(n56) );
  EOI U62 ( .A(n60), .B(n69), .Z(n57) );
  ENI U65 ( .A(A[27]), .B(B[27]), .Z(n60) );
  NR2I U66 ( .A(A[27]), .B(B[27]), .Z(n61) );
  ND2I U67 ( .A(A[27]), .B(B[27]), .Z(n62) );
  EOI U72 ( .A(n73), .B(n67), .Z(n66) );
  ENI U73 ( .A(A[26]), .B(B[26]), .Z(n67) );
  NR2I U74 ( .A(A[26]), .B(B[26]), .Z(n68) );
  ND2I U75 ( .A(A[26]), .B(B[26]), .Z(n69) );
  EOI U81 ( .A(n85), .B(n78), .Z(n74) );
  EOI U82 ( .A(n78), .B(n86), .Z(n75) );
  ENI U85 ( .A(A[25]), .B(B[25]), .Z(n78) );
  NR2I U86 ( .A(A[25]), .B(B[25]), .Z(n79) );
  ND2I U87 ( .A(A[25]), .B(B[25]), .Z(n80) );
  ENI U89 ( .A(n431), .B(n393), .Z(n81) );
  ENI U90 ( .A(n432), .B(n393), .Z(n82) );
  NR2I U93 ( .A(A[24]), .B(B[24]), .Z(n85) );
  ND2I U94 ( .A(A[24]), .B(B[24]), .Z(n86) );
  EOI U106 ( .A(n109), .B(n101), .Z(n97) );
  EOI U107 ( .A(n101), .B(n110), .Z(n98) );
  ENI U110 ( .A(A[23]), .B(B[23]), .Z(n101) );
  NR2I U111 ( .A(A[23]), .B(B[23]), .Z(n102) );
  ND2I U112 ( .A(A[23]), .B(B[23]), .Z(n103) );
  EOI U117 ( .A(n114), .B(n108), .Z(n107) );
  ENI U118 ( .A(A[22]), .B(B[22]), .Z(n108) );
  NR2I U119 ( .A(A[22]), .B(B[22]), .Z(n109) );
  ND2I U120 ( .A(A[22]), .B(B[22]), .Z(n110) );
  EOI U126 ( .A(n126), .B(n119), .Z(n115) );
  EOI U127 ( .A(n119), .B(n127), .Z(n116) );
  ENI U130 ( .A(A[21]), .B(B[21]), .Z(n119) );
  NR2I U131 ( .A(A[21]), .B(B[21]), .Z(n120) );
  ND2I U132 ( .A(A[21]), .B(B[21]), .Z(n121) );
  ENI U134 ( .A(n128), .B(n392), .Z(n122) );
  ENI U135 ( .A(n129), .B(n392), .Z(n123) );
  ND2I U139 ( .A(A[20]), .B(B[20]), .Z(n127) );
  EOI U147 ( .A(n405), .B(n138), .Z(n134) );
  EOI U148 ( .A(n138), .B(n146), .Z(n135) );
  ENI U151 ( .A(A[19]), .B(B[19]), .Z(n138) );
  NR2I U152 ( .A(A[19]), .B(B[19]), .Z(n139) );
  ND2I U153 ( .A(A[19]), .B(B[19]), .Z(n140) );
  ENI U155 ( .A(n151), .B(n456), .Z(n141) );
  ENI U156 ( .A(n152), .B(n456), .Z(n142) );
  NR2I U159 ( .A(A[18]), .B(B[18]), .Z(n145) );
  ND2I U160 ( .A(A[18]), .B(B[18]), .Z(n146) );
  EOI U164 ( .A(n157), .B(n153), .Z(n149) );
  EOI U165 ( .A(n153), .B(n158), .Z(n150) );
  ENI U168 ( .A(A[17]), .B(B[17]), .Z(n153) );
  NR2I U169 ( .A(A[17]), .B(B[17]), .Z(n154) );
  ND2I U170 ( .A(A[17]), .B(B[17]), .Z(n155) );
  NR2I U173 ( .A(A[16]), .B(B[16]), .Z(n157) );
  ND2I U174 ( .A(A[16]), .B(B[16]), .Z(n158) );
  MUX21LP U176 ( .A(n163), .B(n162), .S(n232), .Z(n4) );
  EOI U185 ( .A(n172), .B(n180), .Z(n168) );
  EOI U186 ( .A(n172), .B(n181), .Z(n169) );
  EOI U189 ( .A(A[15]), .B(B[15]), .Z(n172) );
  NR2I U190 ( .A(A[15]), .B(B[15]), .Z(n173) );
  ND2I U191 ( .A(A[15]), .B(B[15]), .Z(n174) );
  ENI U197 ( .A(A[14]), .B(B[14]), .Z(n179) );
  NR2I U198 ( .A(A[14]), .B(B[14]), .Z(n180) );
  ND2I U199 ( .A(A[14]), .B(B[14]), .Z(n181) );
  EOI U205 ( .A(n418), .B(n190), .Z(n186) );
  EOI U206 ( .A(n190), .B(n198), .Z(n187) );
  ENI U209 ( .A(A[13]), .B(B[13]), .Z(n190) );
  NR2I U210 ( .A(A[13]), .B(B[13]), .Z(n191) );
  ND2I U211 ( .A(A[13]), .B(B[13]), .Z(n192) );
  ENI U213 ( .A(n421), .B(n391), .Z(n193) );
  ENI U214 ( .A(n200), .B(n391), .Z(n194) );
  NR2I U217 ( .A(A[12]), .B(B[12]), .Z(n197) );
  ND2I U218 ( .A(A[12]), .B(B[12]), .Z(n198) );
  EOI U226 ( .A(n416), .B(n209), .Z(n205) );
  EOI U227 ( .A(n209), .B(n217), .Z(n206) );
  ENI U230 ( .A(A[11]), .B(B[11]), .Z(n209) );
  NR2I U231 ( .A(A[11]), .B(B[11]), .Z(n210) );
  ND2I U232 ( .A(A[11]), .B(B[11]), .Z(n211) );
  ENI U234 ( .A(n435), .B(n390), .Z(n212) );
  ENI U235 ( .A(n385), .B(n390), .Z(n213) );
  NR2I U238 ( .A(A[10]), .B(B[10]), .Z(n216) );
  ND2I U239 ( .A(A[10]), .B(B[10]), .Z(n217) );
  ENI U247 ( .A(n437), .B(n396), .Z(n224) );
  NR2I U248 ( .A(A[9]), .B(B[9]), .Z(n225) );
  ND2I U249 ( .A(n437), .B(n396), .Z(n226) );
  NR2I U252 ( .A(A[8]), .B(B[8]), .Z(n228) );
  ND2I U253 ( .A(A[8]), .B(B[8]), .Z(n229) );
  MUX21LP U257 ( .A(n235), .B(n236), .S(n264), .Z(n232) );
  EOI U262 ( .A(n398), .B(n241), .Z(n237) );
  EOI U263 ( .A(n241), .B(n248), .Z(n238) );
  EOI U266 ( .A(A[7]), .B(B[7]), .Z(n241) );
  NR2I U267 ( .A(A[7]), .B(B[7]), .Z(n242) );
  ND2I U268 ( .A(A[7]), .B(B[7]), .Z(n243) );
  EOI U270 ( .A(n249), .B(n246), .Z(n244) );
  EOI U271 ( .A(n250), .B(n246), .Z(n245) );
  EOI U272 ( .A(A[6]), .B(B[6]), .Z(n246) );
  NR2I U273 ( .A(A[6]), .B(B[6]), .Z(n247) );
  ND2I U274 ( .A(A[6]), .B(B[6]), .Z(n248) );
  EOI U278 ( .A(n255), .B(n389), .Z(n251) );
  EOI U279 ( .A(n255), .B(n261), .Z(n252) );
  EOI U282 ( .A(A[5]), .B(B[5]), .Z(n255) );
  NR2I U283 ( .A(A[5]), .B(B[5]), .Z(n256) );
  ND2I U284 ( .A(A[5]), .B(B[5]), .Z(n257) );
  ENI U285 ( .A(n262), .B(n455), .Z(SUM[4]) );
  NR2I U288 ( .A(B[4]), .B(A[4]), .Z(n260) );
  ND2I U289 ( .A(B[4]), .B(A[4]), .Z(n261) );
  ENI U298 ( .A(B[3]), .B(A[3]), .Z(n269) );
  NR2I U299 ( .A(B[3]), .B(A[3]), .Z(n270) );
  ND2I U300 ( .A(B[3]), .B(A[3]), .Z(n271) );
  ENI U302 ( .A(B[2]), .B(A[2]), .Z(n272) );
  NR2I U303 ( .A(B[2]), .B(A[2]), .Z(n273) );
  ND2I U304 ( .A(B[2]), .B(A[2]), .Z(n274) );
  NR2I U310 ( .A(B[1]), .B(A[1]), .Z(n279) );
  ND2I U311 ( .A(n427), .B(A[1]), .Z(n280) );
  EOI U312 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  ND2I U313 ( .A(B[0]), .B(A[0]), .Z(n281) );
  IVI U317 ( .A(n452), .Z(n384) );
  MUX21L U318 ( .A(n137), .B(n136), .S(n151), .Z(n132) );
  B2I U319 ( .A(n223), .Z2(n385) );
  MUX21H U320 ( .A(n57), .B(n56), .S(n76), .Z(n386) );
  MUX21H U321 ( .A(n233), .B(n234), .S(n409), .Z(SUM[7]) );
  B3IP U322 ( .A(n4), .Z1(n444), .Z2(n459) );
  IVDAP U323 ( .A(A[9]), .Z(n437) );
  MUX21LP U324 ( .A(n39), .B(n40), .S(n47), .Z(n37) );
  IVI U325 ( .A(A[20]), .Z(n400) );
  IVI U326 ( .A(B[20]), .Z(n401) );
  MUX21H U327 ( .A(n57), .B(n56), .S(n77), .Z(n388) );
  NR2I U328 ( .A(n412), .B(A[4]), .Z(n389) );
  EOI U329 ( .A(A[10]), .B(B[10]), .Z(n390) );
  EOI U330 ( .A(A[12]), .B(B[12]), .Z(n391) );
  EOI U331 ( .A(A[20]), .B(B[20]), .Z(n392) );
  EOI U332 ( .A(A[24]), .B(B[24]), .Z(n393) );
  IVI U333 ( .A(n436), .Z(n394) );
  MUX21L U334 ( .A(n240), .B(n239), .S(n253), .Z(n235) );
  IVI U335 ( .A(B[9]), .Z(n395) );
  IVI U336 ( .A(n395), .Z(n396) );
  IVI U337 ( .A(n4), .Z(n397) );
  NR2I U338 ( .A(A[6]), .B(B[6]), .Z(n398) );
  MUX21L U339 ( .A(n139), .B(n140), .S(n146), .Z(n137) );
  MUX21LP U340 ( .A(n137), .B(n136), .S(n151), .Z(n399) );
  AN2I U341 ( .A(n400), .B(n401), .Z(n126) );
  NR2I U342 ( .A(A[21]), .B(B[21]), .Z(n402) );
  IVI U343 ( .A(n229), .Z(n403) );
  IVI U344 ( .A(n403), .Z(n404) );
  NR2I U345 ( .A(A[18]), .B(B[18]), .Z(n405) );
  ND2I U346 ( .A(B[0]), .B(A[0]), .Z(n406) );
  NR2I U347 ( .A(A[26]), .B(B[26]), .Z(n407) );
  NR2I U348 ( .A(A[25]), .B(B[25]), .Z(n408) );
  IVI U349 ( .A(n262), .Z(n409) );
  MUX21L U350 ( .A(n105), .B(n104), .S(n428), .Z(SUM[22]) );
  MUX21L U351 ( .A(n240), .B(n239), .S(n254), .Z(n236) );
  MUX21L U352 ( .A(n270), .B(n271), .S(n274), .Z(n268) );
  MUX21L U353 ( .A(n270), .B(n271), .S(n273), .Z(n267) );
  MUX21LP U354 ( .A(n166), .B(n167), .S(n204), .Z(n163) );
  MUX21LP U355 ( .A(n163), .B(n162), .S(n232), .Z(n410) );
  MUX21LP U356 ( .A(n166), .B(n167), .S(n203), .Z(n162) );
  IVI U357 ( .A(B[4]), .Z(n411) );
  IVI U358 ( .A(n411), .Z(n412) );
  NR2I U359 ( .A(A[17]), .B(B[17]), .Z(n413) );
  NR2I U360 ( .A(A[5]), .B(B[5]), .Z(n414) );
  NR2I U361 ( .A(A[13]), .B(B[13]), .Z(n415) );
  NR2I U362 ( .A(A[10]), .B(B[10]), .Z(n416) );
  NR2I U363 ( .A(B[2]), .B(A[2]), .Z(n417) );
  NR2I U364 ( .A(A[12]), .B(B[12]), .Z(n418) );
  IVI U365 ( .A(n277), .Z(n419) );
  IVI U366 ( .A(n419), .Z(n420) );
  MUX21LP U367 ( .A(n39), .B(n40), .S(n46), .Z(n36) );
  IVI U368 ( .A(n203), .Z(n421) );
  IVI U369 ( .A(n421), .Z(n422) );
  IVI U370 ( .A(n204), .Z(n423) );
  IVI U371 ( .A(n423), .Z(n424) );
  IVI U372 ( .A(n128), .Z(n425) );
  MUX21LP U373 ( .A(n173), .B(n174), .S(n180), .Z(n170) );
  MUX21LP U374 ( .A(n79), .B(n80), .S(n86), .Z(n77) );
  IVI U375 ( .A(B[1]), .Z(n426) );
  IVI U376 ( .A(n426), .Z(n427) );
  IVI U377 ( .A(n410), .Z(n428) );
  MUX21L U378 ( .A(n429), .B(n430), .S(n397), .Z(SUM[23]) );
  MUX21H U379 ( .A(n93), .B(n94), .S(n133), .Z(n429) );
  MUX21H U380 ( .A(n93), .B(n94), .S(n425), .Z(n430) );
  MUX21LP U381 ( .A(n256), .B(n257), .S(n261), .Z(n254) );
  MUX21LP U382 ( .A(n95), .B(n96), .S(n132), .Z(n431) );
  MUX21LP U383 ( .A(n95), .B(n96), .S(n133), .Z(n432) );
  NR2I U384 ( .A(A[11]), .B(B[11]), .Z(n433) );
  MUX21LP U385 ( .A(n59), .B(n58), .S(n76), .Z(n54) );
  MUX21LP U386 ( .A(n100), .B(n99), .S(n118), .Z(n96) );
  MUX21LP U387 ( .A(n171), .B(n170), .S(n188), .Z(n166) );
  MUX21LP U388 ( .A(n242), .B(n243), .S(n248), .Z(n240) );
  MUX21LP U389 ( .A(n137), .B(n136), .S(n152), .Z(n133) );
  MUX21LP U390 ( .A(n169), .B(n168), .S(n189), .Z(n165) );
  MUX21LP U391 ( .A(n171), .B(n170), .S(n189), .Z(n167) );
  MUX21LP U392 ( .A(n191), .B(n192), .S(n198), .Z(n189) );
  MUX21LP U393 ( .A(n210), .B(n211), .S(n217), .Z(n208) );
  MUX21LP U394 ( .A(n100), .B(n99), .S(n117), .Z(n95) );
  MUX21L U395 ( .A(n112), .B(n111), .S(n452), .Z(SUM[21]) );
  MUX21L U396 ( .A(n29), .B(n28), .S(n428), .Z(SUM[29]) );
  MUX21L U397 ( .A(n19), .B(n18), .S(n397), .Z(SUM[30]) );
  IVI U398 ( .A(n222), .Z(n434) );
  IVI U399 ( .A(n434), .Z(n435) );
  IVI U400 ( .A(n230), .Z(n436) );
  B3IP U401 ( .A(n410), .Z1(n452), .Z2(n458) );
  MUX21LP U402 ( .A(n242), .B(n243), .S(n247), .Z(n239) );
  MUX21LP U403 ( .A(n225), .B(n226), .S(n229), .Z(n223) );
  MUX21LP U404 ( .A(n95), .B(n96), .S(n133), .Z(n6) );
  MUX21LP U405 ( .A(n95), .B(n96), .S(n399), .Z(n8) );
  MUX21H U406 ( .A(n438), .B(n439), .S(n452), .Z(SUM[31]) );
  MUX21H U407 ( .A(n12), .B(n11), .S(n6), .Z(n438) );
  MUX21H U408 ( .A(n12), .B(n11), .S(n8), .Z(n439) );
  MUX21LP U409 ( .A(n208), .B(n207), .S(n222), .Z(n203) );
  MUX21LP U410 ( .A(n208), .B(n207), .S(n223), .Z(n204) );
  MUX21LP U411 ( .A(n59), .B(n58), .S(n77), .Z(n55) );
  MUX21H U412 ( .A(n440), .B(n441), .S(n444), .Z(SUM[25]) );
  MUX21H U413 ( .A(n75), .B(n74), .S(n6), .Z(n440) );
  MUX21H U414 ( .A(n75), .B(n74), .S(n8), .Z(n441) );
  MUX21LP U415 ( .A(n154), .B(n155), .S(n158), .Z(n152) );
  MUX21LP U416 ( .A(n413), .B(n155), .S(n157), .Z(n151) );
  MUX21LP U417 ( .A(n225), .B(n226), .S(n228), .Z(n222) );
  MUX21LP U418 ( .A(n414), .B(n257), .S(n260), .Z(n253) );
  MUX21LP U419 ( .A(n415), .B(n192), .S(n197), .Z(n188) );
  MUX21LP U420 ( .A(n402), .B(n121), .S(n127), .Z(n118) );
  MUX21LP U421 ( .A(n120), .B(n121), .S(n126), .Z(n117) );
  MUX21LP U422 ( .A(n408), .B(n80), .S(n85), .Z(n76) );
  MUX21LP U423 ( .A(n139), .B(n140), .S(n145), .Z(n136) );
  MUX21LP U424 ( .A(n102), .B(n103), .S(n109), .Z(n99) );
  MUX21LP U425 ( .A(n433), .B(n211), .S(n216), .Z(n207) );
  MUX21LP U426 ( .A(n61), .B(n62), .S(n69), .Z(n59) );
  MUX21LP U427 ( .A(n61), .B(n62), .S(n68), .Z(n58) );
  MUX21LP U428 ( .A(n16), .B(n15), .S(n36), .Z(n13) );
  MUX21LP U429 ( .A(n16), .B(n15), .S(n37), .Z(n14) );
  MUX21LP U430 ( .A(n268), .B(n267), .S(n277), .Z(n264) );
  MUX21LP U431 ( .A(n279), .B(n280), .S(n281), .Z(n277) );
  EOI U432 ( .A(n4), .B(n442), .Z(SUM[16]) );
  ENI U433 ( .A(A[16]), .B(B[16]), .Z(n442) );
  ENI U434 ( .A(n443), .B(n406), .Z(SUM[1]) );
  EOI U435 ( .A(A[1]), .B(n427), .Z(n443) );
  MUX21L U436 ( .A(n31), .B(n30), .S(n432), .Z(n29) );
  MUX21L U437 ( .A(n31), .B(n30), .S(n431), .Z(n28) );
  MUX21L U438 ( .A(n48), .B(n49), .S(n459), .Z(SUM[27]) );
  MUX21L U439 ( .A(n388), .B(n386), .S(n6), .Z(n49) );
  MUX21L U440 ( .A(n388), .B(n386), .S(n8), .Z(n48) );
  MUX21L U441 ( .A(n21), .B(n20), .S(n432), .Z(n19) );
  MUX21L U442 ( .A(n21), .B(n20), .S(n431), .Z(n18) );
  MUX21L U443 ( .A(n22), .B(n23), .S(n55), .Z(n21) );
  MUX21L U444 ( .A(n13), .B(n14), .S(n55), .Z(n12) );
  MUX21L U445 ( .A(n135), .B(n134), .S(n152), .Z(n131) );
  MUX21L U446 ( .A(n135), .B(n134), .S(n151), .Z(n130) );
  MUX21L U447 ( .A(n175), .B(n176), .S(n230), .Z(SUM[14]) );
  MUX21L U448 ( .A(n182), .B(n183), .S(n230), .Z(SUM[13]) );
  MUX21L U449 ( .A(n448), .B(n447), .S(n230), .Z(SUM[9]) );
  MUX21L U450 ( .A(n445), .B(n446), .S(n54), .Z(n30) );
  MUX21L U451 ( .A(n22), .B(n23), .S(n54), .Z(n20) );
  MUX21L U452 ( .A(n445), .B(n446), .S(n55), .Z(n31) );
  MUX21L U453 ( .A(n178), .B(n177), .S(n200), .Z(n176) );
  MUX21L U454 ( .A(n178), .B(n177), .S(n421), .Z(n175) );
  MUX21L U455 ( .A(n187), .B(n186), .S(n200), .Z(n183) );
  MUX21L U456 ( .A(n187), .B(n186), .S(n421), .Z(n182) );
  MUX21L U457 ( .A(n161), .B(n160), .S(n436), .Z(SUM[15]) );
  MUX21L U458 ( .A(n164), .B(n165), .S(n424), .Z(n161) );
  MUX21L U459 ( .A(n164), .B(n165), .S(n422), .Z(n160) );
  MUX21L U460 ( .A(n98), .B(n97), .S(n117), .Z(n93) );
  MUX21L U461 ( .A(n98), .B(n97), .S(n118), .Z(n94) );
  MUX21L U462 ( .A(n169), .B(n168), .S(n188), .Z(n164) );
  MUX21L U463 ( .A(n13), .B(n14), .S(n54), .Z(n11) );
  MUX21L U464 ( .A(n107), .B(n106), .S(n129), .Z(n105) );
  MUX21L U465 ( .A(n107), .B(n106), .S(n128), .Z(n104) );
  MUX21L U466 ( .A(n66), .B(n65), .S(n6), .Z(n64) );
  MUX21L U467 ( .A(n66), .B(n65), .S(n8), .Z(n63) );
  MUX21L U468 ( .A(n116), .B(n115), .S(n129), .Z(n112) );
  MUX21L U469 ( .A(n116), .B(n115), .S(n128), .Z(n111) );
  MUX21L U470 ( .A(n41), .B(n42), .S(n384), .Z(SUM[28]) );
  MUX21L U471 ( .A(n44), .B(n43), .S(n6), .Z(n42) );
  MUX21L U472 ( .A(n44), .B(n43), .S(n8), .Z(n41) );
  MUX21L U473 ( .A(n122), .B(n123), .S(n459), .Z(SUM[20]) );
  MUX21H U474 ( .A(n150), .B(n149), .S(n444), .Z(SUM[17]) );
  MUX21L U475 ( .A(n81), .B(n82), .S(n458), .Z(SUM[24]) );
  MUX21L U476 ( .A(n173), .B(n174), .S(n181), .Z(n171) );
  ENI U477 ( .A(n188), .B(n179), .Z(n177) );
  ENI U478 ( .A(n189), .B(n179), .Z(n178) );
  MUX21L U479 ( .A(n193), .B(n194), .S(n230), .Z(SUM[12]) );
  MUX21L U480 ( .A(n201), .B(n202), .S(n394), .Z(SUM[11]) );
  MUX21L U481 ( .A(n206), .B(n205), .S(n435), .Z(n201) );
  MUX21L U482 ( .A(n206), .B(n205), .S(n385), .Z(n202) );
  MUX21L U483 ( .A(n212), .B(n213), .S(n394), .Z(SUM[10]) );
  ENI U484 ( .A(n46), .B(n38), .Z(n445) );
  ENI U485 ( .A(n38), .B(n47), .Z(n446) );
  ENI U486 ( .A(n117), .B(n108), .Z(n106) );
  ENI U487 ( .A(n76), .B(n67), .Z(n65) );
  MUX21L U488 ( .A(n102), .B(n103), .S(n110), .Z(n100) );
  ENI U489 ( .A(n224), .B(n404), .Z(n447) );
  ENI U490 ( .A(n228), .B(n224), .Z(n448) );
  MUX21L U491 ( .A(n238), .B(n237), .S(n253), .Z(n233) );
  MUX21L U492 ( .A(n238), .B(n237), .S(n254), .Z(n234) );
  MUX21L U493 ( .A(n450), .B(n451), .S(n420), .Z(SUM[3]) );
  ENI U494 ( .A(n269), .B(n274), .Z(n450) );
  ENI U495 ( .A(n417), .B(n269), .Z(n451) );
  ENI U496 ( .A(n394), .B(n453), .Z(SUM[8]) );
  EOI U497 ( .A(A[8]), .B(B[8]), .Z(n453) );
  EOI U498 ( .A(A[30]), .B(B[30]), .Z(n454) );
  ENI U499 ( .A(n412), .B(A[4]), .Z(n455) );
  MUX21L U500 ( .A(n245), .B(n244), .S(n262), .Z(SUM[6]) );
  MUX21L U501 ( .A(n252), .B(n251), .S(n262), .Z(SUM[5]) );
  EOI U502 ( .A(A[18]), .B(B[18]), .Z(n456) );
  ENI U503 ( .A(n420), .B(n272), .Z(SUM[2]) );
  MUX21L U504 ( .A(n141), .B(n142), .S(n458), .Z(SUM[18]) );
  MUX21L U505 ( .A(n130), .B(n131), .S(n459), .Z(SUM[19]) );
  MUX21L U506 ( .A(n63), .B(n64), .S(n458), .Z(SUM[26]) );
  IVI U507 ( .A(n77), .Z(n73) );
  IVI U508 ( .A(n264), .Z(n262) );
  IVI U509 ( .A(n254), .Z(n250) );
  IVI U510 ( .A(n253), .Z(n249) );
  IVI U511 ( .A(n232), .Z(n230) );
  IVI U512 ( .A(n204), .Z(n200) );
  IVI U513 ( .A(n133), .Z(n129) );
  IVI U514 ( .A(n399), .Z(n128) );
  IVI U515 ( .A(n118), .Z(n114) );
endmodule


module alu_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n4, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n20, n21, n22,
         n23, n26, n27, n28, n29, n30, n31, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n74, n75, n76, n77, n78,
         n79, n80, n85, n86, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n110, n111, n112, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n145, n146, n151, n152, n153, n154, n155, n156, n157,
         n158, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n216, n217, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n260, n261, n262,
         n264, n267, n268, n269, n271, n272, n273, n274, n277, n278, n279,
         n280, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n312, n313, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n474, n475,
         n476, n477, n478, n480, n481, n482, n483, n484, n485, n486, n487;

  EOI U16 ( .A(n26), .B(n17), .Z(n15) );
  EOI U17 ( .A(n17), .B(n27), .Z(n16) );
  ENI U24 ( .A(n36), .B(n480), .Z(n22) );
  ENI U25 ( .A(n37), .B(n480), .Z(n23) );
  NR2I U28 ( .A(A[30]), .B(n283), .Z(n26) );
  ND2I U29 ( .A(A[30]), .B(n283), .Z(n27) );
  ENI U41 ( .A(n284), .B(A[29]), .Z(n38) );
  NR2I U42 ( .A(n284), .B(A[29]), .Z(n39) );
  ND2I U43 ( .A(n284), .B(A[29]), .Z(n40) );
  EOI U47 ( .A(n54), .B(n45), .Z(n43) );
  EOI U48 ( .A(n55), .B(n45), .Z(n44) );
  ENI U49 ( .A(n285), .B(A[28]), .Z(n45) );
  NR2I U50 ( .A(n285), .B(A[28]), .Z(n46) );
  ND2I U51 ( .A(n285), .B(A[28]), .Z(n47) );
  EOI U61 ( .A(n68), .B(n60), .Z(n56) );
  EOI U62 ( .A(n60), .B(n69), .Z(n57) );
  ENI U65 ( .A(A[27]), .B(n286), .Z(n60) );
  NR2I U66 ( .A(A[27]), .B(n286), .Z(n61) );
  ND2I U67 ( .A(A[27]), .B(n286), .Z(n62) );
  ENI U73 ( .A(n287), .B(A[26]), .Z(n67) );
  NR2I U74 ( .A(n287), .B(A[26]), .Z(n68) );
  ND2I U75 ( .A(n287), .B(A[26]), .Z(n69) );
  EOI U81 ( .A(n85), .B(n78), .Z(n74) );
  EOI U82 ( .A(n78), .B(n86), .Z(n75) );
  ENI U85 ( .A(A[25]), .B(n288), .Z(n78) );
  NR2I U86 ( .A(A[25]), .B(n288), .Z(n79) );
  ND2I U87 ( .A(A[25]), .B(n288), .Z(n80) );
  NR2I U93 ( .A(n289), .B(A[24]), .Z(n85) );
  ND2I U94 ( .A(n289), .B(A[24]), .Z(n86) );
  EOI U106 ( .A(n443), .B(n101), .Z(n97) );
  EOI U107 ( .A(n101), .B(n110), .Z(n98) );
  ENI U110 ( .A(A[23]), .B(n290), .Z(n101) );
  NR2I U111 ( .A(A[23]), .B(n290), .Z(n102) );
  ND2I U112 ( .A(A[23]), .B(n290), .Z(n103) );
  ENI U118 ( .A(A[22]), .B(n291), .Z(n108) );
  ND2I U120 ( .A(A[22]), .B(n291), .Z(n110) );
  EOI U126 ( .A(n455), .B(n119), .Z(n115) );
  EOI U127 ( .A(n119), .B(n127), .Z(n116) );
  ENI U130 ( .A(A[21]), .B(n292), .Z(n119) );
  NR2I U131 ( .A(A[21]), .B(n292), .Z(n120) );
  ND2I U132 ( .A(A[21]), .B(n292), .Z(n121) );
  ENI U134 ( .A(n128), .B(n482), .Z(n122) );
  ENI U135 ( .A(n129), .B(n482), .Z(n123) );
  ND2I U139 ( .A(n293), .B(A[20]), .Z(n127) );
  EOI U147 ( .A(n145), .B(n138), .Z(n134) );
  EOI U148 ( .A(n138), .B(n146), .Z(n135) );
  ENI U151 ( .A(A[19]), .B(n294), .Z(n138) );
  NR2I U152 ( .A(A[19]), .B(n294), .Z(n139) );
  ND2I U153 ( .A(A[19]), .B(n294), .Z(n140) );
  ENI U155 ( .A(n151), .B(n483), .Z(n141) );
  ENI U156 ( .A(n152), .B(n483), .Z(n142) );
  NR2I U159 ( .A(n295), .B(A[18]), .Z(n145) );
  ND2I U160 ( .A(n295), .B(A[18]), .Z(n146) );
  ENI U168 ( .A(A[17]), .B(n296), .Z(n153) );
  NR2I U169 ( .A(A[17]), .B(n296), .Z(n154) );
  ND2I U170 ( .A(A[17]), .B(n296), .Z(n155) );
  EOI U171 ( .A(n460), .B(n156), .Z(DIFF[16]) );
  ENI U172 ( .A(n297), .B(n463), .Z(n156) );
  ND2I U174 ( .A(n297), .B(n463), .Z(n158) );
  EOI U185 ( .A(n172), .B(n180), .Z(n168) );
  EOI U186 ( .A(n172), .B(n181), .Z(n169) );
  EOI U189 ( .A(A[15]), .B(n298), .Z(n172) );
  NR2I U190 ( .A(A[15]), .B(n298), .Z(n173) );
  ND2I U191 ( .A(A[15]), .B(n298), .Z(n174) );
  ENI U197 ( .A(A[14]), .B(n299), .Z(n179) );
  NR2I U198 ( .A(A[14]), .B(n299), .Z(n180) );
  ND2I U199 ( .A(A[14]), .B(n299), .Z(n181) );
  EOI U205 ( .A(n197), .B(n190), .Z(n186) );
  EOI U206 ( .A(n190), .B(n198), .Z(n187) );
  ENI U209 ( .A(A[13]), .B(n300), .Z(n190) );
  NR2I U210 ( .A(A[13]), .B(n300), .Z(n191) );
  ND2I U211 ( .A(A[13]), .B(n300), .Z(n192) );
  ENI U213 ( .A(n199), .B(n478), .Z(n193) );
  ENI U214 ( .A(n200), .B(n478), .Z(n194) );
  NR2I U217 ( .A(n301), .B(A[12]), .Z(n197) );
  ND2I U218 ( .A(n301), .B(A[12]), .Z(n198) );
  EOI U226 ( .A(n216), .B(n209), .Z(n205) );
  EOI U227 ( .A(n209), .B(n217), .Z(n206) );
  ENI U230 ( .A(A[11]), .B(n302), .Z(n209) );
  NR2I U231 ( .A(A[11]), .B(n302), .Z(n210) );
  ND2I U232 ( .A(A[11]), .B(n302), .Z(n211) );
  ENI U234 ( .A(n222), .B(n430), .Z(n212) );
  ENI U235 ( .A(n223), .B(n430), .Z(n213) );
  NR2I U238 ( .A(A[10]), .B(n303), .Z(n216) );
  ND2I U239 ( .A(A[10]), .B(n303), .Z(n217) );
  ENI U247 ( .A(n304), .B(A[9]), .Z(n224) );
  NR2I U248 ( .A(n304), .B(A[9]), .Z(n225) );
  ND2I U249 ( .A(n304), .B(A[9]), .Z(n226) );
  EOI U250 ( .A(n230), .B(n227), .Z(DIFF[8]) );
  ENI U251 ( .A(n305), .B(A[8]), .Z(n227) );
  NR2I U252 ( .A(n305), .B(A[8]), .Z(n228) );
  ND2I U253 ( .A(n305), .B(A[8]), .Z(n229) );
  EOI U262 ( .A(n241), .B(n247), .Z(n237) );
  EOI U263 ( .A(n241), .B(n248), .Z(n238) );
  EOI U266 ( .A(A[7]), .B(n306), .Z(n241) );
  NR2I U267 ( .A(A[7]), .B(n306), .Z(n242) );
  ND2I U268 ( .A(A[7]), .B(n306), .Z(n243) );
  EOI U270 ( .A(n249), .B(n246), .Z(n244) );
  EOI U271 ( .A(n250), .B(n246), .Z(n245) );
  EOI U272 ( .A(n307), .B(A[6]), .Z(n246) );
  NR2I U273 ( .A(n307), .B(A[6]), .Z(n247) );
  ND2I U274 ( .A(n307), .B(A[6]), .Z(n248) );
  EOI U278 ( .A(n260), .B(n255), .Z(n251) );
  EOI U279 ( .A(n255), .B(n261), .Z(n252) );
  EOI U282 ( .A(A[5]), .B(n308), .Z(n255) );
  NR2I U283 ( .A(A[5]), .B(n308), .Z(n256) );
  ND2I U284 ( .A(A[5]), .B(n308), .Z(n257) );
  NR2I U288 ( .A(n309), .B(A[4]), .Z(n260) );
  ND2I U289 ( .A(n309), .B(A[4]), .Z(n261) );
  ENI U298 ( .A(n487), .B(A[3]), .Z(n269) );
  ND2I U300 ( .A(n487), .B(A[3]), .Z(n271) );
  ENI U302 ( .A(n486), .B(A[2]), .Z(n272) );
  NR2I U303 ( .A(n486), .B(A[2]), .Z(n273) );
  ND2I U304 ( .A(n486), .B(A[2]), .Z(n274) );
  EOI U309 ( .A(n312), .B(A[1]), .Z(n278) );
  NR2I U310 ( .A(n312), .B(A[1]), .Z(n279) );
  ND2I U311 ( .A(n312), .B(A[1]), .Z(n280) );
  ENI U312 ( .A(A[0]), .B(n458), .Z(DIFF[0]) );
  MUX21LP U349 ( .A(n175), .B(n176), .S(n454), .Z(DIFF[14]) );
  NR2I U350 ( .A(A[5]), .B(n308), .Z(n416) );
  MUX21LP U351 ( .A(n236), .B(n235), .S(n421), .Z(n464) );
  MUX21LP U352 ( .A(n210), .B(n211), .S(n217), .Z(n208) );
  MUX21H U353 ( .A(n21), .B(n20), .S(n436), .Z(n417) );
  ND2I U354 ( .A(n268), .B(n418), .Z(n419) );
  ND2I U355 ( .A(n267), .B(n277), .Z(n420) );
  ND2I U356 ( .A(n419), .B(n420), .Z(n421) );
  IVI U357 ( .A(n277), .Z(n418) );
  MUX21LP U358 ( .A(n137), .B(n136), .S(n152), .Z(n422) );
  MUX21LP U359 ( .A(n459), .B(n226), .S(n228), .Z(n222) );
  B4I U360 ( .A(B[2]), .Z(n486) );
  MUX21H U361 ( .A(n75), .B(n74), .S(n449), .Z(n423) );
  EOI U362 ( .A(n436), .B(n481), .Z(n424) );
  MUX21H U363 ( .A(n57), .B(n56), .S(n76), .Z(n425) );
  MUX21H U364 ( .A(n21), .B(n20), .S(n6), .Z(n426) );
  MUX21H U365 ( .A(n75), .B(n74), .S(n436), .Z(n427) );
  EOI U366 ( .A(n449), .B(n481), .Z(n428) );
  MUX21H U367 ( .A(n57), .B(n56), .S(n77), .Z(n429) );
  EOI U368 ( .A(A[10]), .B(n303), .Z(n430) );
  ENI U369 ( .A(n228), .B(n224), .Z(n431) );
  MUX21L U370 ( .A(n433), .B(n434), .S(n262), .Z(DIFF[7]) );
  MUX21H U371 ( .A(n238), .B(n237), .S(n254), .Z(n433) );
  MUX21H U372 ( .A(n238), .B(n237), .S(n253), .Z(n434) );
  MUX21L U373 ( .A(n160), .B(n161), .S(n435), .Z(DIFF[15]) );
  IVI U374 ( .A(n464), .Z(n435) );
  MUX21LP U375 ( .A(n162), .B(n163), .S(n438), .Z(n460) );
  MUX21LP U376 ( .A(n95), .B(n96), .S(n132), .Z(n436) );
  MUX21L U377 ( .A(n95), .B(n96), .S(n132), .Z(n8) );
  MUX21LP U378 ( .A(n137), .B(n136), .S(n151), .Z(n132) );
  NR2I U379 ( .A(A[13]), .B(n300), .Z(n437) );
  MUX21LP U380 ( .A(n162), .B(n163), .S(n442), .Z(n4) );
  ND2I U381 ( .A(n440), .B(n441), .Z(n438) );
  B3IP U382 ( .A(n460), .Z1(n466), .Z2(n485) );
  MUX21LP U383 ( .A(n166), .B(n167), .S(n204), .Z(n163) );
  ND2I U384 ( .A(n235), .B(n439), .Z(n440) );
  ND2I U385 ( .A(n236), .B(n264), .Z(n441) );
  ND2I U386 ( .A(n440), .B(n441), .Z(n442) );
  IVI U387 ( .A(n264), .Z(n439) );
  MUX21LP U388 ( .A(n240), .B(n239), .S(n253), .Z(n235) );
  MUX21LP U389 ( .A(n240), .B(n239), .S(n254), .Z(n236) );
  MUX21LP U390 ( .A(n268), .B(n267), .S(n277), .Z(n264) );
  NR2I U391 ( .A(A[22]), .B(n291), .Z(n443) );
  MUX21LP U392 ( .A(n137), .B(n136), .S(n151), .Z(n444) );
  ND2I U393 ( .A(n31), .B(n445), .Z(n446) );
  ND2I U394 ( .A(n30), .B(n449), .Z(n447) );
  ND2I U395 ( .A(n446), .B(n447), .Z(n448) );
  IVI U396 ( .A(n6), .Z(n445) );
  IVI U397 ( .A(n448), .Z(n29) );
  MUX21LP U398 ( .A(n95), .B(n96), .S(n422), .Z(n449) );
  MUX21LP U399 ( .A(n191), .B(n192), .S(n198), .Z(n189) );
  MUX21LP U400 ( .A(n225), .B(n226), .S(n229), .Z(n223) );
  MUX21LP U401 ( .A(n166), .B(n167), .S(n203), .Z(n162) );
  MUX21LP U402 ( .A(n59), .B(n58), .S(n76), .Z(n54) );
  AN2I U403 ( .A(B[16]), .B(n462), .Z(n157) );
  MUX21LP U404 ( .A(n280), .B(n279), .S(n450), .Z(n277) );
  OR2I U405 ( .A(n313), .B(A[0]), .Z(n450) );
  B2I U406 ( .A(n4), .Z2(n484) );
  IVI U407 ( .A(n457), .Z(n451) );
  NR2I U408 ( .A(n451), .B(A[0]), .Z(n452) );
  IVI U409 ( .A(n464), .Z(n453) );
  IVI U410 ( .A(n464), .Z(n454) );
  IVI U411 ( .A(n464), .Z(n230) );
  MUX21LP U412 ( .A(n28), .B(n29), .S(n4), .Z(DIFF[29]) );
  NR2I U413 ( .A(n293), .B(A[20]), .Z(n455) );
  NR2I U414 ( .A(A[21]), .B(n292), .Z(n456) );
  IVI U415 ( .A(n313), .Z(n457) );
  IVI U416 ( .A(n457), .Z(n458) );
  NR2I U417 ( .A(n304), .B(A[9]), .Z(n459) );
  IVI U418 ( .A(B[0]), .Z(n313) );
  NR2I U419 ( .A(n487), .B(A[3]), .Z(n461) );
  IVI U420 ( .A(B[3]), .Z(n487) );
  IVI U421 ( .A(A[16]), .Z(n462) );
  IVI U422 ( .A(n462), .Z(n463) );
  MUX21LP U423 ( .A(n137), .B(n136), .S(n152), .Z(n133) );
  MUX21LP U424 ( .A(n100), .B(n99), .S(n118), .Z(n96) );
  MUX21LP U425 ( .A(n256), .B(n257), .S(n261), .Z(n254) );
  MUX21LP U426 ( .A(n100), .B(n99), .S(n117), .Z(n95) );
  IVI U427 ( .A(n418), .Z(n465) );
  MUX21LP U428 ( .A(n461), .B(n271), .S(n273), .Z(n267) );
  MUX21LP U429 ( .A(n461), .B(n271), .S(n274), .Z(n268) );
  MUX21L U430 ( .A(n242), .B(n243), .S(n247), .Z(n239) );
  MUX21L U431 ( .A(n16), .B(n15), .S(n36), .Z(n13) );
  MUX21LP U432 ( .A(n95), .B(n96), .S(n133), .Z(n6) );
  MUX21LP U433 ( .A(n208), .B(n207), .S(n223), .Z(n204) );
  MUX21LP U434 ( .A(n208), .B(n207), .S(n222), .Z(n203) );
  MUX21H U435 ( .A(n423), .B(n427), .S(n466), .Z(DIFF[25]) );
  MUX21LP U436 ( .A(n154), .B(n155), .S(n158), .Z(n152) );
  MUX21LP U437 ( .A(n154), .B(n155), .S(n157), .Z(n151) );
  MUX21LP U438 ( .A(n437), .B(n192), .S(n197), .Z(n188) );
  MUX21H U439 ( .A(n426), .B(n417), .S(n466), .Z(DIFF[30]) );
  MUX21H U440 ( .A(n428), .B(n424), .S(n466), .Z(DIFF[24]) );
  MUX21LP U441 ( .A(n120), .B(n121), .S(n127), .Z(n118) );
  MUX21LP U442 ( .A(n416), .B(n257), .S(n260), .Z(n253) );
  MUX21LP U443 ( .A(n456), .B(n121), .S(n455), .Z(n117) );
  MUX21LP U444 ( .A(n139), .B(n140), .S(n146), .Z(n137) );
  MUX21LP U445 ( .A(n139), .B(n140), .S(n145), .Z(n136) );
  MUX21LP U446 ( .A(n102), .B(n103), .S(n443), .Z(n99) );
  MUX21LP U447 ( .A(n210), .B(n211), .S(n216), .Z(n207) );
  MUX21LP U448 ( .A(n79), .B(n80), .S(n86), .Z(n77) );
  MUX21LP U449 ( .A(n79), .B(n80), .S(n85), .Z(n76) );
  MUX21LP U450 ( .A(n102), .B(n103), .S(n110), .Z(n100) );
  MUX21LP U451 ( .A(n61), .B(n62), .S(n69), .Z(n59) );
  MUX21LP U452 ( .A(n61), .B(n62), .S(n68), .Z(n58) );
  ENI U453 ( .A(n262), .B(n467), .Z(DIFF[4]) );
  ENI U454 ( .A(n309), .B(A[4]), .Z(n467) );
  MUX21L U455 ( .A(n31), .B(n30), .S(n8), .Z(n28) );
  MUX21L U456 ( .A(n12), .B(n11), .S(n436), .Z(n9) );
  MUX21L U457 ( .A(n429), .B(n425), .S(n436), .Z(n48) );
  MUX21L U458 ( .A(n12), .B(n11), .S(n6), .Z(n10) );
  MUX21L U459 ( .A(n429), .B(n425), .S(n449), .Z(n49) );
  MUX21H U460 ( .A(n93), .B(n94), .S(n444), .Z(n468) );
  MUX21H U461 ( .A(n93), .B(n94), .S(n422), .Z(n469) );
  MUX21L U462 ( .A(n171), .B(n170), .S(n189), .Z(n167) );
  MUX21L U463 ( .A(n171), .B(n170), .S(n188), .Z(n166) );
  MUX21L U464 ( .A(n178), .B(n177), .S(n199), .Z(n175) );
  MUX21L U465 ( .A(n182), .B(n183), .S(n435), .Z(DIFF[13]) );
  MUX21L U466 ( .A(n187), .B(n186), .S(n199), .Z(n182) );
  MUX21L U467 ( .A(n431), .B(n472), .S(n435), .Z(DIFF[9]) );
  MUX21L U468 ( .A(n201), .B(n202), .S(n454), .Z(DIFF[11]) );
  MUX21L U469 ( .A(n206), .B(n205), .S(n222), .Z(n201) );
  MUX21L U470 ( .A(n206), .B(n205), .S(n223), .Z(n202) );
  MUX21L U471 ( .A(n59), .B(n58), .S(n77), .Z(n55) );
  MUX21L U472 ( .A(n470), .B(n471), .S(n54), .Z(n30) );
  MUX21L U473 ( .A(n470), .B(n471), .S(n55), .Z(n31) );
  MUX21L U474 ( .A(n178), .B(n177), .S(n200), .Z(n176) );
  MUX21L U475 ( .A(n187), .B(n186), .S(n200), .Z(n183) );
  MUX21L U476 ( .A(n44), .B(n43), .S(n436), .Z(n41) );
  MUX21L U477 ( .A(n66), .B(n65), .S(n436), .Z(n63) );
  MUX21L U478 ( .A(n164), .B(n165), .S(n204), .Z(n161) );
  MUX21L U479 ( .A(n164), .B(n165), .S(n203), .Z(n160) );
  MUX21L U480 ( .A(n169), .B(n168), .S(n189), .Z(n165) );
  MUX21L U481 ( .A(n13), .B(n14), .S(n54), .Z(n11) );
  MUX21L U482 ( .A(n22), .B(n23), .S(n54), .Z(n20) );
  MUX21L U483 ( .A(n169), .B(n168), .S(n188), .Z(n164) );
  MUX21L U484 ( .A(n44), .B(n43), .S(n449), .Z(n42) );
  MUX21L U485 ( .A(n66), .B(n65), .S(n449), .Z(n64) );
  MUX21L U486 ( .A(n13), .B(n14), .S(n55), .Z(n12) );
  MUX21L U487 ( .A(n22), .B(n23), .S(n55), .Z(n21) );
  MUX21L U488 ( .A(n98), .B(n97), .S(n117), .Z(n93) );
  MUX21L U489 ( .A(n107), .B(n106), .S(n128), .Z(n104) );
  MUX21L U490 ( .A(n116), .B(n115), .S(n128), .Z(n111) );
  MUX21L U491 ( .A(n107), .B(n106), .S(n129), .Z(n105) );
  MUX21L U492 ( .A(n116), .B(n115), .S(n129), .Z(n112) );
  MUX21L U493 ( .A(n98), .B(n97), .S(n118), .Z(n94) );
  MUX21L U494 ( .A(n135), .B(n134), .S(n151), .Z(n130) );
  MUX21L U495 ( .A(n135), .B(n134), .S(n152), .Z(n131) );
  MUX21L U496 ( .A(n242), .B(n243), .S(n248), .Z(n240) );
  MUX21L U497 ( .A(n173), .B(n174), .S(n180), .Z(n170) );
  MUX21L U498 ( .A(n41), .B(n42), .S(n460), .Z(DIFF[28]) );
  MUX21L U499 ( .A(n122), .B(n123), .S(n484), .Z(DIFF[20]) );
  MUX21L U500 ( .A(n63), .B(n64), .S(n485), .Z(DIFF[26]) );
  MUX21L U501 ( .A(n468), .B(n469), .S(n485), .Z(DIFF[23]) );
  MUX21L U502 ( .A(n104), .B(n105), .S(n485), .Z(DIFF[22]) );
  MUX21L U503 ( .A(n111), .B(n112), .S(n460), .Z(DIFF[21]) );
  MUX21L U504 ( .A(n476), .B(n477), .S(n484), .Z(DIFF[17]) );
  MUX21L U505 ( .A(n9), .B(n10), .S(n460), .Z(DIFF[31]) );
  MUX21L U506 ( .A(n141), .B(n142), .S(n484), .Z(DIFF[18]) );
  MUX21L U507 ( .A(n48), .B(n49), .S(n460), .Z(DIFF[27]) );
  MUX21L U508 ( .A(n130), .B(n131), .S(n485), .Z(DIFF[19]) );
  MUX21L U509 ( .A(n193), .B(n194), .S(n453), .Z(DIFF[12]) );
  MUX21L U510 ( .A(n173), .B(n174), .S(n181), .Z(n171) );
  ENI U511 ( .A(n188), .B(n179), .Z(n177) );
  ENI U512 ( .A(n189), .B(n179), .Z(n178) );
  MUX21L U513 ( .A(n212), .B(n213), .S(n453), .Z(DIFF[10]) );
  ENI U514 ( .A(n46), .B(n38), .Z(n470) );
  ENI U515 ( .A(n38), .B(n47), .Z(n471) );
  MUX21L U516 ( .A(n16), .B(n15), .S(n37), .Z(n14) );
  ENI U517 ( .A(n224), .B(n229), .Z(n472) );
  MUX21L U518 ( .A(n39), .B(n40), .S(n46), .Z(n36) );
  MUX21L U519 ( .A(n39), .B(n40), .S(n47), .Z(n37) );
  ENI U520 ( .A(n76), .B(n67), .Z(n65) );
  ENI U521 ( .A(n117), .B(n108), .Z(n106) );
  ENI U522 ( .A(n77), .B(n67), .Z(n66) );
  ENI U523 ( .A(n118), .B(n108), .Z(n107) );
  MUX21L U524 ( .A(n474), .B(n475), .S(n465), .Z(DIFF[3]) );
  ENI U525 ( .A(n269), .B(n274), .Z(n474) );
  ENI U526 ( .A(n273), .B(n269), .Z(n475) );
  ENI U527 ( .A(n157), .B(n153), .Z(n476) );
  ENI U528 ( .A(n153), .B(n158), .Z(n477) );
  MUX21L U529 ( .A(n245), .B(n244), .S(n262), .Z(DIFF[6]) );
  MUX21L U530 ( .A(n252), .B(n251), .S(n262), .Z(DIFF[5]) );
  ENI U531 ( .A(n465), .B(n272), .Z(DIFF[2]) );
  EOI U532 ( .A(n301), .B(A[12]), .Z(n478) );
  EOI U533 ( .A(A[31]), .B(B[31]), .Z(n17) );
  ENI U534 ( .A(n278), .B(n452), .Z(DIFF[1]) );
  EOI U535 ( .A(A[30]), .B(n283), .Z(n480) );
  EOI U536 ( .A(n289), .B(A[24]), .Z(n481) );
  EOI U537 ( .A(n293), .B(A[20]), .Z(n482) );
  EOI U538 ( .A(n295), .B(A[18]), .Z(n483) );
  IVI U539 ( .A(B[1]), .Z(n312) );
  IVI U540 ( .A(B[4]), .Z(n309) );
  IVI U541 ( .A(B[5]), .Z(n308) );
  IVI U542 ( .A(B[6]), .Z(n307) );
  IVI U543 ( .A(B[7]), .Z(n306) );
  IVI U544 ( .A(B[8]), .Z(n305) );
  IVI U545 ( .A(B[9]), .Z(n304) );
  IVI U546 ( .A(B[10]), .Z(n303) );
  IVI U547 ( .A(B[11]), .Z(n302) );
  IVI U548 ( .A(B[12]), .Z(n301) );
  IVI U549 ( .A(B[13]), .Z(n300) );
  IVI U550 ( .A(B[14]), .Z(n299) );
  IVI U551 ( .A(B[15]), .Z(n298) );
  IVI U552 ( .A(B[16]), .Z(n297) );
  IVI U553 ( .A(B[17]), .Z(n296) );
  IVI U554 ( .A(B[18]), .Z(n295) );
  IVI U555 ( .A(B[19]), .Z(n294) );
  IVI U556 ( .A(B[20]), .Z(n293) );
  IVI U557 ( .A(B[21]), .Z(n292) );
  IVI U558 ( .A(B[22]), .Z(n291) );
  IVI U559 ( .A(B[23]), .Z(n290) );
  IVI U560 ( .A(B[24]), .Z(n289) );
  IVI U561 ( .A(B[25]), .Z(n288) );
  IVI U562 ( .A(B[26]), .Z(n287) );
  IVI U563 ( .A(B[27]), .Z(n286) );
  IVI U564 ( .A(B[28]), .Z(n285) );
  IVI U565 ( .A(B[29]), .Z(n284) );
  IVI U566 ( .A(B[30]), .Z(n283) );
  IVI U567 ( .A(n264), .Z(n262) );
  IVI U568 ( .A(n254), .Z(n250) );
  IVI U569 ( .A(n253), .Z(n249) );
  IVI U570 ( .A(n204), .Z(n200) );
  IVI U571 ( .A(n203), .Z(n199) );
  IVI U572 ( .A(n133), .Z(n129) );
  IVI U573 ( .A(n444), .Z(n128) );
endmodule


module alu_DW_cmp_1 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151;

  NR2I U10 ( .A(n151), .B(A[31]), .Z(n9) );
  ND2I U11 ( .A(n151), .B(A[31]), .Z(n10) );
  NR2I U12 ( .A(n150), .B(B[30]), .Z(n11) );
  ND2I U13 ( .A(n150), .B(B[30]), .Z(n12) );
  NR2I U16 ( .A(n149), .B(B[29]), .Z(n15) );
  ND2I U17 ( .A(n149), .B(B[29]), .Z(n16) );
  NR2I U18 ( .A(n148), .B(B[28]), .Z(n17) );
  ND2I U19 ( .A(n148), .B(B[28]), .Z(n18) );
  NR2I U24 ( .A(n147), .B(B[27]), .Z(n23) );
  ND2I U25 ( .A(n147), .B(B[27]), .Z(n24) );
  NR2I U26 ( .A(n146), .B(B[26]), .Z(n25) );
  ND2I U27 ( .A(n146), .B(B[26]), .Z(n26) );
  NR2I U30 ( .A(n145), .B(B[25]), .Z(n29) );
  ND2I U31 ( .A(n145), .B(B[25]), .Z(n30) );
  NR2I U32 ( .A(n144), .B(B[24]), .Z(n31) );
  ND2I U33 ( .A(n144), .B(B[24]), .Z(n32) );
  NR2I U40 ( .A(n143), .B(B[23]), .Z(n39) );
  ND2I U41 ( .A(n143), .B(B[23]), .Z(n40) );
  NR2I U42 ( .A(n142), .B(B[22]), .Z(n41) );
  ND2I U43 ( .A(n142), .B(B[22]), .Z(n42) );
  NR2I U46 ( .A(n141), .B(B[21]), .Z(n45) );
  ND2I U47 ( .A(n141), .B(B[21]), .Z(n46) );
  NR2I U48 ( .A(n140), .B(B[20]), .Z(n47) );
  ND2I U49 ( .A(n140), .B(B[20]), .Z(n48) );
  NR2I U54 ( .A(n139), .B(B[19]), .Z(n53) );
  ND2I U55 ( .A(n139), .B(B[19]), .Z(n54) );
  NR2I U56 ( .A(n138), .B(B[18]), .Z(n55) );
  ND2I U57 ( .A(n138), .B(B[18]), .Z(n56) );
  NR2I U60 ( .A(n137), .B(B[17]), .Z(n59) );
  ND2I U61 ( .A(n137), .B(B[17]), .Z(n60) );
  NR2I U62 ( .A(n136), .B(B[16]), .Z(n61) );
  ND2I U63 ( .A(n136), .B(B[16]), .Z(n62) );
  NR2I U71 ( .A(n135), .B(B[15]), .Z(n70) );
  ND2I U72 ( .A(n135), .B(B[15]), .Z(n71) );
  NR2I U73 ( .A(n134), .B(B[14]), .Z(n72) );
  ND2I U74 ( .A(n134), .B(B[14]), .Z(n73) );
  NR2I U77 ( .A(n133), .B(B[13]), .Z(n76) );
  ND2I U78 ( .A(n133), .B(B[13]), .Z(n77) );
  NR2I U79 ( .A(n132), .B(B[12]), .Z(n78) );
  ND2I U80 ( .A(n132), .B(B[12]), .Z(n79) );
  NR2I U85 ( .A(n131), .B(B[11]), .Z(n84) );
  ND2I U86 ( .A(n131), .B(B[11]), .Z(n85) );
  NR2I U87 ( .A(n130), .B(B[10]), .Z(n86) );
  ND2I U88 ( .A(n130), .B(B[10]), .Z(n87) );
  NR2I U91 ( .A(n129), .B(B[9]), .Z(n90) );
  ND2I U92 ( .A(n129), .B(B[9]), .Z(n91) );
  NR2I U93 ( .A(n128), .B(B[8]), .Z(n92) );
  ND2I U94 ( .A(n128), .B(B[8]), .Z(n93) );
  NR2I U100 ( .A(n127), .B(B[7]), .Z(n99) );
  ND2I U101 ( .A(n127), .B(B[7]), .Z(n100) );
  NR2I U102 ( .A(n126), .B(B[6]), .Z(n101) );
  ND2I U103 ( .A(n126), .B(B[6]), .Z(n102) );
  NR2I U106 ( .A(n125), .B(B[5]), .Z(n105) );
  ND2I U107 ( .A(n125), .B(B[5]), .Z(n106) );
  NR2I U108 ( .A(n124), .B(B[4]), .Z(n107) );
  ND2I U109 ( .A(n124), .B(B[4]), .Z(n108) );
  NR2I U113 ( .A(B[3]), .B(n123), .Z(n112) );
  ND2I U114 ( .A(B[3]), .B(n123), .Z(n113) );
  NR2I U115 ( .A(B[2]), .B(n122), .Z(n114) );
  ND2I U116 ( .A(B[2]), .B(n122), .Z(n115) );
  NR2I U118 ( .A(n121), .B(B[1]), .Z(n117) );
  ND2I U119 ( .A(n121), .B(B[1]), .Z(n118) );
  ND2I U120 ( .A(n120), .B(B[0]), .Z(n119) );
  MUX21L U765 ( .A(n65), .B(n64), .S(n94), .Z(n63) );
  IVI U766 ( .A(A[9]), .Z(n129) );
  MUX21LP U767 ( .A(n45), .B(n46), .S(n48), .Z(n44) );
  MUX21LP U768 ( .A(n45), .B(n46), .S(n47), .Z(n43) );
  MUX21L U769 ( .A(n1), .B(n2), .S(n63), .Z(GE_LT_GT_LE) );
  MUX21LP U770 ( .A(n4), .B(n3), .S(n33), .Z(n1) );
  MUX21LP U771 ( .A(n4), .B(n3), .S(n34), .Z(n2) );
  MUX21LP U772 ( .A(n23), .B(n24), .S(n25), .Z(n21) );
  MUX21LP U773 ( .A(n69), .B(n68), .S(n75), .Z(n67) );
  MUX21L U774 ( .A(n53), .B(n54), .S(n55), .Z(n51) );
  MUX21L U775 ( .A(n9), .B(n10), .S(n11), .Z(n7) );
  MUX21LP U776 ( .A(n69), .B(n68), .S(n74), .Z(n66) );
  MUX21L U777 ( .A(n112), .B(n113), .S(n114), .Z(n110) );
  MUX21L U778 ( .A(n112), .B(n113), .S(n115), .Z(n111) );
  MUX21L U779 ( .A(n95), .B(n96), .S(n109), .Z(n94) );
  MUX21L U780 ( .A(n98), .B(n97), .S(n104), .Z(n96) );
  MUX21L U781 ( .A(n98), .B(n97), .S(n103), .Z(n95) );
  MUX21L U782 ( .A(n111), .B(n110), .S(n116), .Z(n109) );
  MUX21L U783 ( .A(n117), .B(n118), .S(n119), .Z(n116) );
  MUX21L U784 ( .A(n66), .B(n67), .S(n80), .Z(n64) );
  MUX21L U785 ( .A(n83), .B(n82), .S(n88), .Z(n80) );
  MUX21L U786 ( .A(n90), .B(n91), .S(n92), .Z(n88) );
  MUX21L U787 ( .A(n105), .B(n106), .S(n107), .Z(n103) );
  MUX21L U788 ( .A(n35), .B(n36), .S(n49), .Z(n33) );
  MUX21L U789 ( .A(n52), .B(n51), .S(n57), .Z(n49) );
  MUX21L U790 ( .A(n59), .B(n60), .S(n61), .Z(n57) );
  MUX21L U791 ( .A(n66), .B(n67), .S(n81), .Z(n65) );
  MUX21L U792 ( .A(n83), .B(n82), .S(n89), .Z(n81) );
  MUX21L U793 ( .A(n90), .B(n91), .S(n93), .Z(n89) );
  MUX21L U794 ( .A(n70), .B(n71), .S(n72), .Z(n68) );
  MUX21L U795 ( .A(n39), .B(n40), .S(n41), .Z(n37) );
  MUX21L U796 ( .A(n70), .B(n71), .S(n73), .Z(n69) );
  MUX21L U797 ( .A(n76), .B(n77), .S(n78), .Z(n74) );
  MUX21L U798 ( .A(n76), .B(n77), .S(n79), .Z(n75) );
  MUX21L U799 ( .A(n84), .B(n85), .S(n86), .Z(n82) );
  MUX21L U800 ( .A(n84), .B(n85), .S(n87), .Z(n83) );
  MUX21L U801 ( .A(n53), .B(n54), .S(n56), .Z(n52) );
  MUX21L U802 ( .A(n38), .B(n37), .S(n43), .Z(n35) );
  MUX21L U803 ( .A(n23), .B(n24), .S(n26), .Z(n22) );
  MUX21L U804 ( .A(n38), .B(n37), .S(n44), .Z(n36) );
  MUX21L U805 ( .A(n39), .B(n40), .S(n42), .Z(n38) );
  MUX21L U806 ( .A(n99), .B(n100), .S(n101), .Z(n97) );
  MUX21L U807 ( .A(n99), .B(n100), .S(n102), .Z(n98) );
  MUX21L U808 ( .A(n5), .B(n6), .S(n19), .Z(n3) );
  MUX21L U809 ( .A(n22), .B(n21), .S(n27), .Z(n19) );
  MUX21L U810 ( .A(n29), .B(n30), .S(n31), .Z(n27) );
  MUX21L U811 ( .A(n5), .B(n6), .S(n20), .Z(n4) );
  MUX21L U812 ( .A(n22), .B(n21), .S(n28), .Z(n20) );
  MUX21L U813 ( .A(n29), .B(n30), .S(n32), .Z(n28) );
  MUX21L U814 ( .A(n8), .B(n7), .S(n13), .Z(n5) );
  MUX21L U815 ( .A(n15), .B(n16), .S(n17), .Z(n13) );
  MUX21L U816 ( .A(n8), .B(n7), .S(n14), .Z(n6) );
  MUX21L U817 ( .A(n15), .B(n16), .S(n18), .Z(n14) );
  MUX21L U818 ( .A(n105), .B(n106), .S(n108), .Z(n104) );
  MUX21L U819 ( .A(n35), .B(n36), .S(n50), .Z(n34) );
  MUX21L U820 ( .A(n52), .B(n51), .S(n58), .Z(n50) );
  MUX21L U821 ( .A(n59), .B(n60), .S(n62), .Z(n58) );
  MUX21L U822 ( .A(n9), .B(n10), .S(n12), .Z(n8) );
  IVI U823 ( .A(B[31]), .Z(n151) );
  IVI U824 ( .A(A[30]), .Z(n150) );
  IVI U825 ( .A(A[29]), .Z(n149) );
  IVI U826 ( .A(A[28]), .Z(n148) );
  IVI U827 ( .A(A[27]), .Z(n147) );
  IVI U828 ( .A(A[26]), .Z(n146) );
  IVI U829 ( .A(A[25]), .Z(n145) );
  IVI U830 ( .A(A[24]), .Z(n144) );
  IVI U831 ( .A(A[23]), .Z(n143) );
  IVI U832 ( .A(A[22]), .Z(n142) );
  IVI U833 ( .A(A[21]), .Z(n141) );
  IVI U834 ( .A(A[20]), .Z(n140) );
  IVI U835 ( .A(A[19]), .Z(n139) );
  IVI U836 ( .A(A[18]), .Z(n138) );
  IVI U837 ( .A(A[17]), .Z(n137) );
  IVI U838 ( .A(A[16]), .Z(n136) );
  IVI U839 ( .A(A[15]), .Z(n135) );
  IVI U840 ( .A(A[14]), .Z(n134) );
  IVI U841 ( .A(A[13]), .Z(n133) );
  IVI U842 ( .A(A[12]), .Z(n132) );
  IVI U843 ( .A(A[11]), .Z(n131) );
  IVI U844 ( .A(A[10]), .Z(n130) );
  IVI U845 ( .A(A[8]), .Z(n128) );
  IVI U846 ( .A(A[7]), .Z(n127) );
  IVI U847 ( .A(A[6]), .Z(n126) );
  IVI U848 ( .A(A[5]), .Z(n125) );
  IVI U849 ( .A(A[4]), .Z(n124) );
  IVI U850 ( .A(A[3]), .Z(n123) );
  IVI U851 ( .A(A[2]), .Z(n122) );
  IVI U852 ( .A(A[1]), .Z(n121) );
  IVI U853 ( .A(A[0]), .Z(n120) );
endmodule


module alu ( r1, r2, control, result );
  input [31:0] r1;
  input [31:0] r2;
  input [2:0] control;
  output [31:0] result;
  wire   N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N159, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080;

  alu_DW01_add_1 add_17 ( .A(r1), .B({n192, n116, n225, r2[28:26], n152, 
        r2[24:23], n127, n194, n189, n41, r2[18:16], n138, n299, n211, n298, 
        r2[11:8], n251, n147, n224, r2[4], n373, n343, n350, n348}), .CI(1'b0), 
        .SUM({N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31}) );
  alu_DW01_sub_1 sub_23 ( .A({r1[31:10], n103, r1[8:0]}), .B({n220, r2[30:16], 
        n138, r2[14:4], n373, n48, n266, n349}), .CI(1'b0), .DIFF({N223, N222, 
        N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, 
        N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, 
        N197, N196, N195, N194, N193, N192}) );
  alu_DW_cmp_1 lt_21 ( .A({r1[31:27], n209, r1[25:17], n50, r1[15:13], n260, 
        n106, n258, n103, r1[8], n107, r1[6:5], n226, r1[3:0]}), .B({n192, 
        r2[30], n217, r2[28:26], n152, r2[24:23], n127, n194, n189, n41, n166, 
        r2[17], n155, n138, r2[14], n211, n298, r2[11], n218, n23, n196, n251, 
        n147, n224, n227, n373, n343, n231, n161}), .TC(1'b1), .GE_LT(1'b1), 
        .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N159) );
  MUX21H U3 ( .A(r1[5]), .B(n257), .S(n123), .Z(n314) );
  IVI U4 ( .A(n802), .Z(n1) );
  IVI U5 ( .A(n1), .Z(n2) );
  IVI U6 ( .A(n513), .Z(n3) );
  IVI U7 ( .A(n3), .Z(n4) );
  NR2I U8 ( .A(n141), .B(n142), .Z(n5) );
  IVI U12 ( .A(n6), .Z(n7) );
  ND4P U13 ( .A(n840), .B(n878), .C(n915), .D(n157), .Z(n550) );
  IVI U14 ( .A(n212), .Z(n8) );
  ND2I U15 ( .A(n292), .B(n49), .Z(n9) );
  B4I U16 ( .A(n9), .Z(n121) );
  ND4 U17 ( .A(n611), .B(n610), .C(n609), .D(n608), .Z(result[8]) );
  IVI U18 ( .A(n570), .Z(n10) );
  IVI U19 ( .A(n902), .Z(n12) );
  IVI U20 ( .A(n12), .Z(n16) );
  IVI U21 ( .A(n335), .Z(n17) );
  IVI U22 ( .A(n17), .Z(n18) );
  ND4P U23 ( .A(n833), .B(n832), .C(n831), .D(n830), .Z(n834) );
  AO2 U24 ( .A(n281), .B(n782), .C(n781), .D(n222), .Z(n789) );
  B4I U25 ( .A(r2[30]), .Z(n1044) );
  IVI U26 ( .A(n24), .Z(n19) );
  IVDAP U27 ( .A(r1[8]), .Y(n24), .Z(n25) );
  AO3 U28 ( .A(n961), .B(n101), .C(n960), .D(n959), .Z(n962) );
  IVI U29 ( .A(n275), .Z(n20) );
  IVI U30 ( .A(n441), .Z(n21) );
  IVI U31 ( .A(n489), .Z(n22) );
  B3I U32 ( .A(r2[19]), .Z1(n40), .Z2(n41) );
  B2I U33 ( .A(r2[9]), .Z2(n23) );
  AN2I U34 ( .A(n587), .B(n377), .Z(n26) );
  AO3 U35 ( .A(n270), .B(n176), .C(n776), .D(n775), .Z(n777) );
  AO2 U36 ( .A(n74), .B(n601), .C(n203), .D(n54), .Z(n568) );
  IVI U37 ( .A(n60), .Z(n907) );
  AO2 U38 ( .A(n843), .B(n16), .C(n281), .D(n973), .Z(n833) );
  AO2 U39 ( .A(n852), .B(n843), .C(n190), .D(n338), .Z(n768) );
  IVDAP U40 ( .A(n368), .Y(n27), .Z(n28) );
  B3I U41 ( .A(n496), .Z1(n29), .Z2(n30) );
  IVDAP U42 ( .A(n371), .Y(n31), .Z(n32) );
  IVDAP U43 ( .A(r1[3]), .Y(n33), .Z(n34) );
  B2IP U44 ( .A(n312), .Z2(n35) );
  ND3P U45 ( .A(control[1]), .B(n401), .C(n421), .Z(n36) );
  IVDAP U46 ( .A(r1[6]), .Y(n37), .Z(n38) );
  AN2I U47 ( .A(n381), .B(n421), .Z(n39) );
  IVDAP U48 ( .A(r1[28]), .Y(n42), .Z(n43) );
  B3I U49 ( .A(r1[27]), .Z1(n44), .Z2(n45) );
  OR2I U50 ( .A(r2[25]), .B(r2[23]), .Z(n46) );
  B3I U51 ( .A(r2[22]), .Z1(n47), .Z2(n127) );
  B2IP U52 ( .A(r2[2]), .Z2(n48) );
  B3I U53 ( .A(n329), .Z1(n330), .Z2(n331) );
  IVDAP U54 ( .A(r1[16]), .Y(n49), .Z(n50) );
  IVDAP U55 ( .A(r1[20]), .Y(n51), .Z(n52) );
  IVDAP U56 ( .A(n876), .Y(n6), .Z(n53) );
  IVDA U57 ( .A(r1[4]), .Y(n54), .Z(n55) );
  AN2I U58 ( .A(r1[31]), .B(n102), .Z(n56) );
  AN4P U59 ( .A(n775), .B(n819), .C(n859), .D(n738), .Z(n57) );
  AN4P U60 ( .A(n861), .B(n895), .C(n931), .D(n817), .Z(n58) );
  B4IP U61 ( .A(r1[1]), .Z(n523) );
  AN2I U62 ( .A(r1[0]), .B(n278), .Z(n59) );
  IVDAP U63 ( .A(n285), .Y(n291), .Z(n292) );
  AO2P U64 ( .A(n334), .B(n953), .C(n994), .D(n934), .Z(n935) );
  ND2I U65 ( .A(n61), .B(n62), .Z(n60) );
  ND2I U66 ( .A(n16), .B(n272), .Z(n61) );
  ND2I U67 ( .A(n26), .B(n1020), .Z(n62) );
  AN2I U68 ( .A(n373), .B(n48), .Z(n63) );
  B4I U69 ( .A(n63), .Z(n661) );
  ND2I U70 ( .A(n261), .B(n924), .Z(n64) );
  IVI U71 ( .A(n306), .Z(n65) );
  IVI U72 ( .A(n65), .Z(n66) );
  IVDA U73 ( .A(r2[26]), .Z(n67) );
  AO7 U74 ( .A(n936), .B(n378), .C(n935), .Z(n937) );
  IVI U75 ( .A(n289), .Z(n180) );
  IVI U76 ( .A(n292), .Z(n68) );
  AO2P U77 ( .A(n171), .B(n33), .C(n119), .D(n37), .Z(n567) );
  AN2I U78 ( .A(n152), .B(n938), .Z(n69) );
  AN2I U79 ( .A(n300), .B(n937), .Z(n70) );
  NR2I U80 ( .A(n69), .B(n70), .Z(n941) );
  AN2I U81 ( .A(n169), .B(n695), .Z(n71) );
  NR2I U82 ( .A(n71), .B(n228), .Z(n696) );
  IVI U83 ( .A(n289), .Z(n72) );
  ND2I U84 ( .A(n20), .B(n317), .Z(n73) );
  IVI U85 ( .A(n177), .Z(n74) );
  B3I U86 ( .A(n289), .Z1(n278), .Z2(n287) );
  ND2I U87 ( .A(n64), .B(n404), .Z(n75) );
  B4I U88 ( .A(n370), .Z(n343) );
  B4IP U89 ( .A(r1[2]), .Z(n542) );
  MUX21LP U90 ( .A(n267), .B(n34), .S(n124), .Z(n466) );
  AN2I U91 ( .A(n173), .B(n478), .Z(n76) );
  AN2I U92 ( .A(n292), .B(n33), .Z(n77) );
  NR2I U93 ( .A(n76), .B(n77), .Z(n479) );
  AO2P U94 ( .A(n169), .B(n542), .C(n278), .D(n601), .Z(n543) );
  AN2I U95 ( .A(n168), .B(n1050), .Z(n78) );
  AN2I U96 ( .A(n290), .B(n42), .Z(n79) );
  NR2I U97 ( .A(n78), .B(n79), .Z(n408) );
  AO2 U98 ( .A(n1016), .B(n760), .C(n759), .D(n222), .Z(n767) );
  MUX21L U99 ( .A(n1058), .B(n1050), .S(n124), .Z(n457) );
  IVI U100 ( .A(r1[0]), .Z(n478) );
  AO2 U101 ( .A(r2[27]), .B(n975), .C(n306), .D(n974), .Z(n980) );
  AO2 U102 ( .A(n52), .B(n845), .C(n844), .D(n212), .Z(n854) );
  AO2 U103 ( .A(n251), .B(n580), .C(n341), .D(n579), .Z(n591) );
  AO4 U104 ( .A(n216), .B(n823), .C(n495), .D(n1062), .Z(n505) );
  AN4P U105 ( .A(n860), .B(n818), .C(n774), .D(n892), .Z(n80) );
  MUX21H U106 ( .A(n334), .B(n862), .S(n344), .Z(n81) );
  AN4P U107 ( .A(n932), .B(n894), .C(n858), .D(n965), .Z(n82) );
  B4I U108 ( .A(n191), .Z(n103) );
  AN2I U109 ( .A(n545), .B(n375), .Z(n83) );
  AN2I U110 ( .A(n597), .B(n377), .Z(n84) );
  AN2I U111 ( .A(n620), .B(n378), .Z(n85) );
  AN4P U112 ( .A(n917), .B(n916), .C(n915), .D(n64), .Z(n86) );
  AN4P U113 ( .A(n756), .B(n719), .C(n678), .D(n794), .Z(n87) );
  AN2I U114 ( .A(n636), .B(n378), .Z(n88) );
  AN4P U115 ( .A(n840), .B(n839), .C(n838), .D(n837), .Z(n89) );
  AN2I U116 ( .A(n700), .B(n699), .Z(n90) );
  B2I U117 ( .A(n708), .Z2(n91) );
  AN3 U118 ( .A(n422), .B(n421), .C(control[2]), .Z(n93) );
  AO3 U119 ( .A(n259), .B(n206), .C(n659), .D(n658), .Z(n737) );
  ND4 U120 ( .A(n697), .B(n659), .C(n622), .D(n739), .Z(n440) );
  IVI U121 ( .A(n95), .Z(n94) );
  IVI U122 ( .A(n301), .Z(n95) );
  IVI U123 ( .A(n95), .Z(n96) );
  IVI U124 ( .A(n288), .Z(n97) );
  ND4 U125 ( .A(n591), .B(n590), .C(n589), .D(n588), .Z(result[7]) );
  IVDAP U126 ( .A(n316), .Y(n124), .Z(n123) );
  NR2I U127 ( .A(n141), .B(n142), .Z(n98) );
  IVI U128 ( .A(r1[4]), .Z(n99) );
  IVI U129 ( .A(r1[4]), .Z(n256) );
  ND4P U130 ( .A(n453), .B(n452), .C(n451), .D(n450), .Z(result[1]) );
  ND4P U131 ( .A(n530), .B(n529), .C(n528), .D(n527), .Z(result[4]) );
  ND4P U132 ( .A(n628), .B(n627), .C(n626), .D(n625), .Z(result[9]) );
  AO2P U133 ( .A(N201), .B(n39), .C(N40), .D(n35), .Z(n625) );
  AO6 U134 ( .A(n273), .B(n234), .C(n997), .Z(n998) );
  B4I U135 ( .A(n680), .Z(n259) );
  ND4P U136 ( .A(n574), .B(n573), .C(n572), .D(n571), .Z(result[6]) );
  AO2P U137 ( .A(n147), .B(n556), .C(n342), .D(n555), .Z(n574) );
  ND4P U138 ( .A(n705), .B(n704), .C(n703), .D(n702), .Z(result[13]) );
  AO2P U139 ( .A(N205), .B(n39), .C(N44), .D(n35), .Z(n702) );
  ND4P U140 ( .A(n728), .B(n727), .C(n726), .D(n725), .Z(result[14]) );
  AO2P U141 ( .A(N206), .B(n39), .C(N45), .D(n35), .Z(n725) );
  IVI U142 ( .A(n1006), .Z(n100) );
  IVI U143 ( .A(n100), .Z(n101) );
  ND4P U144 ( .A(n549), .B(n548), .C(n547), .D(n546), .Z(result[5]) );
  AO2P U145 ( .A(n224), .B(n536), .C(n340), .D(n535), .Z(n549) );
  ND4P U146 ( .A(n917), .B(n951), .C(n559), .D(n53), .Z(n709) );
  ND4P U147 ( .A(n477), .B(n476), .C(n475), .D(n474), .Z(result[2]) );
  IVI U148 ( .A(n68), .Z(n102) );
  ND4P U149 ( .A(n752), .B(n751), .C(n750), .D(n749), .Z(result[15]) );
  ND2I U150 ( .A(n104), .B(n105), .Z(n997) );
  OR2P U151 ( .A(n996), .B(n42), .Z(n104) );
  OR2I U152 ( .A(n1032), .B(n183), .Z(n105) );
  IVI U153 ( .A(n657), .Z(n106) );
  IVI U154 ( .A(n208), .Z(n107) );
  AO2 U155 ( .A(n169), .B(n99), .C(n180), .D(n208), .Z(n108) );
  IVI U156 ( .A(n176), .Z(n109) );
  IVI U157 ( .A(n168), .Z(n176) );
  ND2I U158 ( .A(n328), .B(n37), .Z(n110) );
  ND2I U159 ( .A(n202), .B(n601), .Z(n111) );
  AN2I U160 ( .A(n110), .B(n111), .Z(n586) );
  AN2I U161 ( .A(n48), .B(n198), .Z(n112) );
  AN2I U162 ( .A(n373), .B(n744), .Z(n113) );
  NR2I U163 ( .A(n112), .B(n113), .Z(n660) );
  B5I U164 ( .A(n167), .Z(n174) );
  B3IP U165 ( .A(n329), .Z1(n332), .Z2(n333) );
  IVI U166 ( .A(n1042), .Z(n114) );
  IVI U167 ( .A(n114), .Z(n115) );
  IVI U168 ( .A(n1044), .Z(n116) );
  ND2I U169 ( .A(n120), .B(n953), .Z(n117) );
  ND2I U170 ( .A(n952), .B(n994), .Z(n118) );
  AN2I U171 ( .A(n117), .B(n118), .Z(n954) );
  B5IP U172 ( .A(n971), .Z(n994) );
  AO7 U173 ( .A(n955), .B(n378), .C(n954), .Z(n956) );
  AN4P U174 ( .A(n878), .B(n877), .C(n876), .D(n875), .Z(n120) );
  OR2I U175 ( .A(r2[10]), .B(r2[9]), .Z(n122) );
  IVDAP U176 ( .A(n286), .Y(n119), .Z(n288) );
  IVI U177 ( .A(n286), .Z(n125) );
  IVAP U178 ( .A(n370), .Z(n344) );
  IVI U179 ( .A(n981), .Z(n126) );
  ND2I U180 ( .A(n89), .B(n953), .Z(n128) );
  ND2I U181 ( .A(n994), .B(n86), .Z(n129) );
  AN2I U182 ( .A(n128), .B(n129), .Z(n918) );
  B4IP U183 ( .A(n970), .Z(n953) );
  B4IP U184 ( .A(r1[25]), .Z(n942) );
  ND2I U185 ( .A(n167), .B(n24), .Z(n130) );
  ND2I U186 ( .A(n179), .B(n657), .Z(n131) );
  AN2I U187 ( .A(n130), .B(n131), .Z(n658) );
  AO3P U188 ( .A(n259), .B(n207), .C(n659), .D(n658), .Z(n132) );
  ND2I U189 ( .A(n74), .B(n489), .Z(n133) );
  ND2I U190 ( .A(n63), .B(n744), .Z(n134) );
  ND2I U191 ( .A(n994), .B(n898), .Z(n135) );
  AN2I U192 ( .A(n134), .B(n135), .Z(n745) );
  NR3P U193 ( .A(n393), .B(r2[24]), .C(n46), .Z(n397) );
  AN2I U194 ( .A(n169), .B(n1058), .Z(n136) );
  NR2I U195 ( .A(n136), .B(n482), .Z(n483) );
  ND2I U196 ( .A(n648), .B(n32), .Z(n137) );
  ND2I U197 ( .A(n137), .B(n492), .Z(n823) );
  B5IP U198 ( .A(n265), .Z(n266) );
  IVI U199 ( .A(n387), .Z(n138) );
  EON1P U200 ( .A(n246), .B(n230), .C(n81), .D(n281), .Z(n872) );
  IVI U201 ( .A(n1016), .Z(n283) );
  ND2I U202 ( .A(n949), .B(n558), .Z(n139) );
  ND2I U203 ( .A(n98), .B(n140), .Z(n708) );
  IVI U204 ( .A(n139), .Z(n140) );
  NR2I U205 ( .A(r1[28]), .B(n207), .Z(n141) );
  NR2I U206 ( .A(r1[27]), .B(n177), .Z(n142) );
  IVI U207 ( .A(n290), .Z(n143) );
  B4I U208 ( .A(r1[24]), .Z(n924) );
  EO1P U209 ( .A(n48), .B(n805), .C(n376), .D(n319), .Z(n642) );
  IVI U210 ( .A(r2[10]), .Z(n144) );
  ND2I U211 ( .A(N159), .B(n93), .Z(n423) );
  AN2I U212 ( .A(N47), .B(n35), .Z(n145) );
  NR2I U213 ( .A(n145), .B(n769), .Z(n770) );
  AO2P U214 ( .A(n29), .B(n517), .C(n342), .D(n516), .Z(n530) );
  AO7P U215 ( .A(n4), .B(n1068), .C(n310), .Z(n416) );
  MUX21LP U216 ( .A(n689), .B(n221), .S(n373), .Z(n539) );
  MUX21LP U217 ( .A(n732), .B(n1070), .S(n373), .Z(n900) );
  IVDAP U218 ( .A(r2[0]), .Y(n264), .Z(n349) );
  IVI U219 ( .A(n1006), .Z(n209) );
  MUX21LP U220 ( .A(n577), .B(n57), .S(n48), .Z(n653) );
  MUX21LP U221 ( .A(n553), .B(n551), .S(n48), .Z(n632) );
  MUX21LP U222 ( .A(n533), .B(n531), .S(n48), .Z(n615) );
  MUX21LP U223 ( .A(n514), .B(n87), .S(n48), .Z(n593) );
  MUX21LP U224 ( .A(n80), .B(n82), .S(n48), .Z(n612) );
  AO4P U225 ( .A(n804), .B(n803), .C(n335), .D(n2), .Z(n810) );
  IVI U226 ( .A(r2[6]), .Z(n146) );
  B4IP U227 ( .A(n146), .Z(n147) );
  AO2P U228 ( .A(N207), .B(n39), .C(N46), .D(n35), .Z(n749) );
  OR2I U229 ( .A(n1009), .B(n103), .Z(n641) );
  AO3 U230 ( .A(n19), .B(n206), .C(n641), .D(n640), .Z(n148) );
  IVI U231 ( .A(n670), .Z(n149) );
  IVI U232 ( .A(n149), .Z(n150) );
  IVI U233 ( .A(r2[25]), .Z(n151) );
  B4IP U234 ( .A(n151), .Z(n152) );
  ND2I U235 ( .A(n328), .B(n499), .Z(n153) );
  AO2P U236 ( .A(n311), .B(n805), .C(n953), .D(n714), .Z(n722) );
  IVI U237 ( .A(n629), .Z(n154) );
  AO7P U238 ( .A(r1[31]), .B(n143), .C(n1053), .Z(n1057) );
  IVI U239 ( .A(n184), .Z(n155) );
  IVI U240 ( .A(n184), .Z(n156) );
  IVI U241 ( .A(n184), .Z(n185) );
  ND2I U242 ( .A(n180), .B(n801), .Z(n157) );
  IVI U243 ( .A(n805), .Z(n158) );
  IVI U244 ( .A(n158), .Z(n159) );
  EON1P U245 ( .A(n414), .B(n1062), .C(n412), .D(n29), .Z(n417) );
  AO3P U246 ( .A(n43), .B(n332), .C(n1055), .D(n483), .Z(n484) );
  IVI U247 ( .A(n291), .Z(n160) );
  IVI U248 ( .A(n215), .Z(n161) );
  AO3 U249 ( .A(n672), .B(n971), .C(n661), .D(n520), .Z(n162) );
  NR2I U250 ( .A(n406), .B(n405), .Z(n163) );
  IVI U251 ( .A(n242), .Z(n164) );
  IVI U252 ( .A(n164), .Z(n165) );
  IVI U253 ( .A(n803), .Z(n166) );
  MUX21LP U254 ( .A(n583), .B(n56), .S(n48), .Z(n648) );
  IVI U255 ( .A(n186), .Z(n167) );
  IVI U256 ( .A(n1007), .Z(n168) );
  IVI U257 ( .A(n1007), .Z(n169) );
  IVI U258 ( .A(n1007), .Z(n170) );
  IVI U259 ( .A(n1007), .Z(n171) );
  IVI U260 ( .A(n186), .Z(n172) );
  IVI U261 ( .A(n1007), .Z(n173) );
  IVI U262 ( .A(n167), .Z(n175) );
  ND2I U263 ( .A(n349), .B(n265), .Z(n177) );
  AN4P U264 ( .A(n839), .B(n153), .C(n9), .D(n875), .Z(n178) );
  IVI U265 ( .A(n286), .Z(n179) );
  IVI U266 ( .A(n319), .Z(n181) );
  B3IP U267 ( .A(n285), .Z1(n289), .Z2(n290) );
  IVI U268 ( .A(n394), .Z(n182) );
  IVI U269 ( .A(n668), .Z(n183) );
  B3IP U270 ( .A(r2[1]), .Z1(n265), .Z2(n350) );
  B2I U271 ( .A(n494), .Z1(n231), .Z2(n232) );
  IVI U272 ( .A(r2[16]), .Z(n184) );
  ND2I U273 ( .A(n350), .B(n349), .Z(n186) );
  ND2I U274 ( .A(n163), .B(n950), .Z(n187) );
  IVI U275 ( .A(n215), .Z(n197) );
  IVI U276 ( .A(r2[20]), .Z(n188) );
  B4IP U277 ( .A(n188), .Z(n189) );
  IVI U278 ( .A(n412), .Z(n190) );
  EO1P U279 ( .A(N200), .B(n39), .C(n321), .D(n302), .Z(n609) );
  IVI U280 ( .A(r1[9]), .Z(n191) );
  IVI U281 ( .A(n1076), .Z(n192) );
  IVI U282 ( .A(r2[21]), .Z(n193) );
  B4IP U283 ( .A(n193), .Z(n194) );
  IVI U284 ( .A(r2[29]), .Z(n195) );
  IVI U285 ( .A(n382), .Z(n196) );
  AO2P U286 ( .A(n266), .B(n478), .C(n197), .D(n523), .Z(n454) );
  ND2I U287 ( .A(n586), .B(n108), .Z(n198) );
  IVI U288 ( .A(n1008), .Z(n199) );
  AO3P U289 ( .A(n982), .B(n302), .C(n980), .D(n979), .Z(n983) );
  AO2P U290 ( .A(n45), .B(n978), .C(n977), .D(n234), .Z(n979) );
  ND4P U291 ( .A(n511), .B(n510), .C(n509), .D(n508), .Z(result[3]) );
  IVI U292 ( .A(n1010), .Z(n200) );
  IVI U293 ( .A(n1010), .Z(n201) );
  IVI U294 ( .A(n1010), .Z(n202) );
  IVI U295 ( .A(n1010), .Z(n203) );
  IVI U296 ( .A(n271), .Z(n204) );
  IVI U297 ( .A(n271), .Z(n205) );
  IVI U298 ( .A(n271), .Z(n206) );
  IVI U299 ( .A(n271), .Z(n207) );
  AO3P U300 ( .A(n925), .B(n924), .C(n923), .D(n922), .Z(n926) );
  IVI U301 ( .A(r1[7]), .Z(n208) );
  IVI U302 ( .A(r2[13]), .Z(n210) );
  B4IP U303 ( .A(n210), .Z(n211) );
  IVI U304 ( .A(n899), .Z(n212) );
  AO2P U305 ( .A(n326), .B(n99), .C(n201), .D(n33), .Z(n544) );
  IVI U306 ( .A(r2[17]), .Z(n213) );
  IVI U307 ( .A(n213), .Z(n214) );
  IVI U308 ( .A(n348), .Z(n215) );
  IVI U309 ( .A(n227), .Z(n216) );
  AO2P U310 ( .A(n939), .B(n234), .C(n85), .D(n338), .Z(n940) );
  IVI U311 ( .A(n394), .Z(n217) );
  B5I U312 ( .A(n144), .Z(n218) );
  IVI U313 ( .A(r2[31]), .Z(n219) );
  IVI U314 ( .A(n1076), .Z(n220) );
  IVI U315 ( .A(n1018), .Z(n221) );
  OR2P U316 ( .A(n248), .B(n249), .Z(n889) );
  IVI U317 ( .A(n806), .Z(n222) );
  AO1P U318 ( .A(N52), .B(n35), .C(n872), .D(n871), .Z(n873) );
  AO3P U319 ( .A(n18), .B(n870), .C(n869), .D(n868), .Z(n871) );
  IVI U320 ( .A(r2[5]), .Z(n223) );
  B4IP U321 ( .A(n223), .Z(n224) );
  AO2 U322 ( .A(n161), .B(n1058), .C(n266), .D(n1050), .Z(n432) );
  MUX21LP U323 ( .A(n467), .B(n314), .S(n266), .Z(n468) );
  IVI U324 ( .A(n394), .Z(n225) );
  IVI U325 ( .A(n99), .Z(n226) );
  IVI U326 ( .A(n496), .Z(n227) );
  AO2P U327 ( .A(n881), .B(n901), .C(n10), .D(n1020), .Z(n886) );
  MUX21LP U328 ( .A(n150), .B(n183), .S(n344), .Z(n597) );
  B4IP U329 ( .A(r1[30]), .Z(n1058) );
  AN2I U330 ( .A(n290), .B(n441), .Z(n228) );
  IVI U331 ( .A(n286), .Z(n229) );
  IVI U332 ( .A(n779), .Z(n230) );
  ND4P U333 ( .A(n40), .B(n847), .C(n392), .D(n47), .Z(n393) );
  ND2I U334 ( .A(n480), .B(n479), .Z(n233) );
  IVI U335 ( .A(n284), .Z(n234) );
  IVI U336 ( .A(n783), .Z(n1020) );
  ND2I U337 ( .A(n235), .B(n236), .Z(n274) );
  ND2I U338 ( .A(n953), .B(n753), .Z(n235) );
  ND2I U339 ( .A(n994), .B(n758), .Z(n236) );
  IVI U340 ( .A(n228), .Z(n237) );
  ND2I U341 ( .A(N56), .B(n312), .Z(n238) );
  IVI U342 ( .A(n944), .Z(n239) );
  AN2I U343 ( .A(n238), .B(n239), .Z(n945) );
  IVI U344 ( .A(n287), .Z(n240) );
  AO3P U345 ( .A(n943), .B(n942), .C(n941), .D(n940), .Z(n944) );
  B5I U346 ( .A(n657), .Z(n241) );
  AN4P U347 ( .A(n797), .B(n796), .C(n795), .D(n794), .Z(n242) );
  OR2I U348 ( .A(n848), .B(n847), .Z(n243) );
  OR2I U349 ( .A(n245), .B(n846), .Z(n244) );
  ND2I U350 ( .A(n243), .B(n244), .Z(n851) );
  AO1P U351 ( .A(n852), .B(n222), .C(n851), .D(n850), .Z(n853) );
  AO3P U352 ( .A(n902), .B(n971), .C(n661), .D(n660), .Z(n662) );
  AO2P U353 ( .A(r2[24]), .B(n921), .C(n94), .D(n920), .Z(n923) );
  AO4P U354 ( .A(n1036), .B(n1060), .C(n1068), .D(n1035), .Z(n1040) );
  MUX21LP U355 ( .A(n159), .B(n181), .S(n344), .Z(n569) );
  IVI U356 ( .A(n339), .Z(n245) );
  EO1P U357 ( .A(n84), .B(n338), .C(n607), .D(n284), .Z(n922) );
  IVI U358 ( .A(n212), .Z(n246) );
  ND4P U359 ( .A(n426), .B(n425), .C(n424), .D(n423), .Z(result[0]) );
  AO1P U360 ( .A(n606), .B(n1016), .C(n420), .D(n419), .Z(n424) );
  AO2P U361 ( .A(n306), .B(n1073), .C(r1[31]), .D(n1072), .Z(n1074) );
  OR2I U362 ( .A(n606), .B(n377), .Z(n247) );
  ND2I U363 ( .A(n247), .B(n605), .Z(n607) );
  OR2I U364 ( .A(n823), .B(n337), .Z(n324) );
  AO2P U365 ( .A(n864), .B(n901), .C(n83), .D(n234), .Z(n869) );
  IVI U366 ( .A(r2[3]), .Z(n374) );
  NR3P U367 ( .A(n386), .B(r2[11]), .C(n122), .Z(n399) );
  NR2I U368 ( .A(n1036), .B(n282), .Z(n248) );
  NR2I U369 ( .A(n246), .B(n879), .Z(n249) );
  IVI U370 ( .A(r2[7]), .Z(n250) );
  B4IP U371 ( .A(n250), .Z(n251) );
  MUX21LP U372 ( .A(n120), .B(n242), .S(n344), .Z(n1036) );
  AO7P U373 ( .A(n919), .B(n31), .C(n918), .Z(n920) );
  AO2P U374 ( .A(n63), .B(n320), .C(n994), .D(n879), .Z(n721) );
  ND4P U375 ( .A(n951), .B(n950), .C(n949), .D(n948), .Z(n1035) );
  NR2I U376 ( .A(n1059), .B(n282), .Z(n252) );
  NR2I U377 ( .A(n8), .B(n898), .Z(n253) );
  OR2P U378 ( .A(n252), .B(n253), .Z(n910) );
  MUX21LP U379 ( .A(n897), .B(n896), .S(n344), .Z(n1059) );
  AO3 U380 ( .A(n990), .B(n283), .C(n854), .D(n853), .Z(n855) );
  AN2I U381 ( .A(N59), .B(n35), .Z(n254) );
  NR2I U382 ( .A(n254), .B(n1002), .Z(n1003) );
  ND4P U383 ( .A(n933), .B(n932), .C(n931), .D(n930), .Z(n1013) );
  MUX21LP U384 ( .A(n862), .B(n779), .S(n344), .Z(n936) );
  AO7 U385 ( .A(n606), .B(n377), .C(n605), .Z(n321) );
  MUX21LP U386 ( .A(n841), .B(n844), .S(n344), .Z(n919) );
  AN2I U387 ( .A(N51), .B(n35), .Z(n255) );
  NR2I U388 ( .A(n255), .B(n855), .Z(n856) );
  AO2P U389 ( .A(n311), .B(n187), .C(n953), .D(n519), .Z(n411) );
  IVI U390 ( .A(n256), .Z(n257) );
  AO2P U391 ( .A(n328), .B(n1008), .C(n201), .D(n1058), .Z(n409) );
  AO2P U392 ( .A(n311), .B(n824), .C(n953), .D(n737), .Z(n746) );
  IVI U393 ( .A(n695), .Z(n258) );
  IVI U394 ( .A(n439), .Z(n260) );
  AO3P U395 ( .A(r1[8]), .B(n204), .C(n641), .D(n640), .Z(n714) );
  IVI U396 ( .A(n286), .Z(n261) );
  AN2I U397 ( .A(n953), .B(n604), .Z(n262) );
  AN2I U398 ( .A(n994), .B(n753), .Z(n263) );
  NR2I U399 ( .A(n262), .B(n263), .Z(n605) );
  ND4P U400 ( .A(n839), .B(n153), .C(n754), .D(n875), .Z(n512) );
  AO3P U401 ( .A(n1069), .B(n1068), .C(n1067), .D(n1066), .Z(n1075) );
  AO2P U402 ( .A(n333), .B(n542), .C(n203), .D(n523), .Z(n480) );
  ND4P U403 ( .A(n895), .B(n894), .C(n893), .D(n892), .Z(n969) );
  AO2P U404 ( .A(n173), .B(n54), .C(n72), .D(n208), .Z(n585) );
  IVI U405 ( .A(n542), .Z(n267) );
  ND2I U406 ( .A(n63), .B(n995), .Z(n268) );
  ND2I U407 ( .A(n994), .B(n512), .Z(n269) );
  AN2I U408 ( .A(n268), .B(n269), .Z(n410) );
  IVI U409 ( .A(n462), .Z(n270) );
  MUX21LP U410 ( .A(n198), .B(n233), .S(n344), .Z(n587) );
  AN2I U411 ( .A(n350), .B(n264), .Z(n271) );
  AO6P U412 ( .A(n229), .B(n695), .C(n639), .Z(n640) );
  AO3P U413 ( .A(n267), .B(n291), .C(n174), .D(n454), .Z(n807) );
  ND2I U414 ( .A(n350), .B(n349), .Z(n1007) );
  AO2P U415 ( .A(n958), .B(n234), .C(n88), .D(n338), .Z(n959) );
  AO3P U416 ( .A(n1077), .B(n1076), .C(n1075), .D(n1074), .Z(n1078) );
  IVI U417 ( .A(n806), .Z(n272) );
  IVI U418 ( .A(n806), .Z(n901) );
  AO3P U419 ( .A(n1001), .B(n283), .C(n999), .D(n998), .Z(n1002) );
  AO3P U420 ( .A(n199), .B(n288), .C(n175), .D(n432), .Z(n687) );
  AO3P U421 ( .A(n881), .B(n971), .C(n661), .D(n642), .Z(n643) );
  AO6P U422 ( .A(n526), .B(n32), .C(n274), .Z(n273) );
  AO3P U423 ( .A(n38), .B(n176), .C(n622), .D(n621), .Z(n694) );
  ND2I U424 ( .A(n1042), .B(n30), .Z(n275) );
  IVI U425 ( .A(n801), .Z(n276) );
  IVI U426 ( .A(n275), .Z(n277) );
  AO6P U427 ( .A(N58), .B(n35), .C(n983), .Z(n984) );
  MUX21LP U428 ( .A(n708), .B(n1033), .S(n344), .Z(n636) );
  MUX21LP U429 ( .A(n154), .B(n91), .S(n344), .Z(n712) );
  OR2I U430 ( .A(n808), .B(n320), .Z(n279) );
  OR2I U431 ( .A(n806), .B(n159), .Z(n280) );
  ND2I U432 ( .A(n279), .B(n280), .Z(n809) );
  NR3P U433 ( .A(n284), .B(n526), .C(n32), .Z(n850) );
  AO3P U434 ( .A(n336), .B(n887), .C(n886), .D(n885), .Z(n888) );
  IVI U435 ( .A(n1000), .Z(n281) );
  IVI U436 ( .A(n1016), .Z(n282) );
  AO1P U437 ( .A(N53), .B(n35), .C(n889), .D(n888), .Z(n890) );
  AO2P U438 ( .A(n67), .B(n957), .C(n301), .D(n956), .Z(n960) );
  ND2I U439 ( .A(n313), .B(n317), .Z(n284) );
  MUX21LP U440 ( .A(n759), .B(n59), .S(n344), .Z(n526) );
  B3IP U441 ( .A(n1054), .Z1(n285), .Z2(n286) );
  AO3P U442 ( .A(n955), .B(n283), .C(n812), .D(n811), .Z(n813) );
  B5I U443 ( .A(n439), .Z(n293) );
  AN2I U444 ( .A(n171), .B(n601), .Z(n294) );
  NR2I U445 ( .A(n294), .B(n600), .Z(n602) );
  AO1P U446 ( .A(n418), .B(n593), .C(n417), .D(n416), .Z(n419) );
  AO6P U447 ( .A(N57), .B(n35), .C(n962), .Z(n963) );
  ND2I U448 ( .A(n318), .B(n277), .Z(n295) );
  AN3P U449 ( .A(control[0]), .B(control[2]), .C(n422), .Z(n318) );
  AO6P U450 ( .A(n29), .B(n1065), .C(n1064), .Z(n1066) );
  AO6P U451 ( .A(N55), .B(n312), .C(n926), .Z(n927) );
  AN2I U452 ( .A(n318), .B(n277), .Z(n296) );
  IVI U453 ( .A(r2[12]), .Z(n297) );
  B4IP U454 ( .A(n297), .Z(n298) );
  IVI U455 ( .A(n388), .Z(n299) );
  ND4P U456 ( .A(n790), .B(n789), .C(n788), .D(n787), .Z(n791) );
  AO2P U457 ( .A(n864), .B(n843), .C(n773), .D(n341), .Z(n790) );
  ND2I U458 ( .A(n989), .B(n31), .Z(n1000) );
  AO3P U459 ( .A(n672), .B(n971), .C(n661), .D(n520), .Z(n846) );
  B2I U460 ( .A(r2[0]), .Z1(n316), .Z2(n348) );
  IVI U461 ( .A(n981), .Z(n300) );
  IVI U462 ( .A(n73), .Z(n301) );
  IVI U463 ( .A(n300), .Z(n302) );
  IVI U464 ( .A(n73), .Z(n989) );
  IVI U465 ( .A(n296), .Z(n337) );
  ND2I U466 ( .A(N62), .B(n35), .Z(n303) );
  IVI U467 ( .A(n1078), .Z(n304) );
  AN2I U468 ( .A(n303), .B(n304), .Z(n1079) );
  AO1P U469 ( .A(N54), .B(n35), .C(n910), .D(n909), .Z(n911) );
  AO3P U470 ( .A(n908), .B(n336), .C(n907), .D(n906), .Z(n909) );
  AO6P U471 ( .A(N48), .B(n312), .C(n791), .Z(n792) );
  AO2P U472 ( .A(n373), .B(n995), .C(n48), .D(n670), .Z(n520) );
  ND3P U473 ( .A(n195), .B(n1044), .C(n219), .Z(n395) );
  ND4P U474 ( .A(n385), .B(n384), .C(n383), .D(n382), .Z(n386) );
  ND4P U475 ( .A(n916), .B(n133), .C(n837), .D(n948), .Z(n519) );
  AO2P U476 ( .A(n307), .B(n992), .C(r2[28]), .D(n991), .Z(n999) );
  NR4P U477 ( .A(n395), .B(r2[28]), .C(r2[27]), .D(r2[26]), .Z(n396) );
  ND4P U478 ( .A(n768), .B(n767), .C(n766), .D(n765), .Z(n769) );
  ND4P U479 ( .A(n390), .B(n389), .C(n388), .D(n387), .Z(n391) );
  AO6P U480 ( .A(n170), .B(n680), .C(n679), .Z(n681) );
  AO3P U481 ( .A(n241), .B(n332), .C(n682), .D(n681), .Z(n758) );
  AO4P U482 ( .A(n1063), .B(n1062), .C(n1061), .D(n1060), .Z(n1064) );
  AN2I U483 ( .A(n338), .B(n373), .Z(n305) );
  AN2I U484 ( .A(n339), .B(n31), .Z(n306) );
  AN2I U485 ( .A(n300), .B(n373), .Z(n307) );
  AN2I U486 ( .A(n301), .B(n994), .Z(n308) );
  MUX21L U487 ( .A(n57), .B(n58), .S(n344), .Z(n733) );
  AN2I U488 ( .A(n667), .B(n994), .Z(n309) );
  B4I U489 ( .A(n354), .Z(n364) );
  IVI U490 ( .A(n368), .Z(n365) );
  IVI U491 ( .A(n368), .Z(n367) );
  IVI U492 ( .A(n368), .Z(n366) );
  AO2 U493 ( .A(n953), .B(n582), .C(n994), .D(n575), .Z(n492) );
  AO2 U494 ( .A(n333), .B(n33), .C(n201), .D(n542), .Z(n525) );
  MUX21L U495 ( .A(n619), .B(n221), .S(n344), .Z(n620) );
  AN2I U496 ( .A(n318), .B(n115), .Z(n310) );
  AN2I U497 ( .A(n373), .B(n370), .Z(n311) );
  AN3 U498 ( .A(n421), .B(n401), .C(n422), .Z(n312) );
  IVI U499 ( .A(n319), .Z(n320) );
  AO2 U500 ( .A(n327), .B(n24), .C(n201), .D(n208), .Z(n621) );
  AN2I U501 ( .A(n29), .B(n1042), .Z(n313) );
  AO3 U502 ( .A(r1[13]), .B(n174), .C(n756), .D(n755), .Z(n757) );
  MUX21H U503 ( .A(n257), .B(n34), .S(n123), .Z(n315) );
  AN3 U504 ( .A(control[0]), .B(control[1]), .C(n401), .Z(n317) );
  IVI U505 ( .A(n807), .Z(n319) );
  AN2I U506 ( .A(N49), .B(n312), .Z(n322) );
  NR2I U507 ( .A(n322), .B(n813), .Z(n814) );
  AN2I U508 ( .A(N50), .B(n312), .Z(n323) );
  NR2I U509 ( .A(n323), .B(n834), .Z(n835) );
  ND2I U510 ( .A(n825), .B(n272), .Z(n325) );
  AN2I U511 ( .A(n324), .B(n325), .Z(n832) );
  AO3P U512 ( .A(n293), .B(n330), .C(n697), .D(n696), .Z(n863) );
  IVI U513 ( .A(n177), .Z(n326) );
  IVI U514 ( .A(n177), .Z(n327) );
  IVI U515 ( .A(n1009), .Z(n328) );
  IVI U516 ( .A(n1009), .Z(n329) );
  AN4P U517 ( .A(n861), .B(n860), .C(n859), .D(n858), .Z(n334) );
  IVI U518 ( .A(n296), .Z(n335) );
  IVI U519 ( .A(n296), .Z(n336) );
  IVI U520 ( .A(n295), .Z(n338) );
  IVI U521 ( .A(n295), .Z(n339) );
  IVI U522 ( .A(n336), .Z(n340) );
  IVI U523 ( .A(n337), .Z(n341) );
  IVI U524 ( .A(n337), .Z(n342) );
  NR4P U525 ( .A(n391), .B(r2[18]), .C(r2[17]), .D(n185), .Z(n398) );
  ND2I U526 ( .A(n350), .B(n264), .Z(n1010) );
  ND2I U527 ( .A(n494), .B(n264), .Z(n1054) );
  AO3P U528 ( .A(n107), .B(n332), .C(n603), .D(n602), .Z(n753) );
  B4IP U529 ( .A(n374), .Z(n373) );
  B2IP U530 ( .A(n1029), .Z1(n92), .Z2(n345) );
  B2IP U531 ( .A(n92), .Z2(n346) );
  B2IP U532 ( .A(n92), .Z2(n347) );
  IVI U533 ( .A(n363), .Z(n351) );
  IVI U534 ( .A(n363), .Z(n352) );
  IVI U535 ( .A(n363), .Z(n353) );
  IVI U536 ( .A(n360), .Z(n354) );
  IVI U537 ( .A(n362), .Z(n355) );
  IVI U538 ( .A(n362), .Z(n356) );
  IVI U539 ( .A(n362), .Z(n357) );
  IVI U540 ( .A(n360), .Z(n358) );
  IVI U541 ( .A(n360), .Z(n359) );
  IVI U542 ( .A(n1030), .Z(n360) );
  IVI U543 ( .A(n1030), .Z(n361) );
  IVI U544 ( .A(n1030), .Z(n362) );
  IVI U545 ( .A(n1030), .Z(n363) );
  IVI U546 ( .A(n36), .Z(n368) );
  IVI U547 ( .A(n36), .Z(n369) );
  IVI U548 ( .A(r2[2]), .Z(n370) );
  IVI U549 ( .A(n372), .Z(n371) );
  IVI U550 ( .A(r2[3]), .Z(n372) );
  IVI U551 ( .A(n371), .Z(n375) );
  IVI U552 ( .A(n371), .Z(n376) );
  IVI U553 ( .A(n371), .Z(n377) );
  IVI U554 ( .A(n371), .Z(n378) );
  IVI U555 ( .A(control[0]), .Z(n421) );
  IVI U556 ( .A(control[2]), .Z(n401) );
  IVI U557 ( .A(control[1]), .Z(n422) );
  ND2I U558 ( .A(control[2]), .B(control[1]), .Z(n379) );
  IVI U559 ( .A(n379), .Z(n381) );
  ND2I U560 ( .A(control[0]), .B(n381), .Z(n1030) );
  AO7 U561 ( .A(r1[0]), .B(n355), .C(n365), .Z(n380) );
  AO2 U562 ( .A(N31), .B(n35), .C(n161), .D(n380), .Z(n426) );
  ND2I U563 ( .A(N192), .B(n39), .Z(n425) );
  IVI U564 ( .A(r2[1]), .Z(n494) );
  ND2I U565 ( .A(n59), .B(n370), .Z(n761) );
  IVI U566 ( .A(n761), .Z(n606) );
  IVI U567 ( .A(r2[5]), .Z(n385) );
  IVI U568 ( .A(r2[6]), .Z(n384) );
  IVI U569 ( .A(r2[7]), .Z(n383) );
  IVI U570 ( .A(r2[8]), .Z(n382) );
  IVI U571 ( .A(r2[12]), .Z(n390) );
  IVI U572 ( .A(r2[13]), .Z(n389) );
  IVI U573 ( .A(r2[14]), .Z(n388) );
  IVI U574 ( .A(r2[15]), .Z(n387) );
  IVI U575 ( .A(r2[20]), .Z(n847) );
  IVI U576 ( .A(r2[21]), .Z(n392) );
  IVI U577 ( .A(r2[29]), .Z(n394) );
  IVI U578 ( .A(r2[31]), .Z(n1076) );
  ND4 U579 ( .A(n399), .B(n398), .C(n397), .D(n396), .Z(n400) );
  IVI U580 ( .A(n400), .Z(n1042) );
  IVI U581 ( .A(r2[4]), .Z(n496) );
  ND2I U582 ( .A(n20), .B(n317), .Z(n981) );
  IVI U583 ( .A(n1000), .Z(n1016) );
  ND3 U584 ( .A(control[0]), .B(n401), .C(n422), .Z(n1029) );
  MUX21L U585 ( .A(n364), .B(n346), .S(n124), .Z(n402) );
  AO6 U586 ( .A(n402), .B(n365), .C(n478), .Z(n420) );
  ND2I U587 ( .A(n373), .B(n30), .Z(n1060) );
  IVI U588 ( .A(n1060), .Z(n418) );
  IVI U589 ( .A(r1[10]), .Z(n695) );
  ND2I U590 ( .A(n201), .B(n695), .Z(n682) );
  ND2I U591 ( .A(n349), .B(n265), .Z(n1009) );
  IVI U592 ( .A(r1[9]), .Z(n680) );
  ND2I U593 ( .A(n229), .B(n24), .Z(n599) );
  IVI U594 ( .A(r1[11]), .Z(n657) );
  ND2I U595 ( .A(n172), .B(n657), .Z(n716) );
  ND4 U596 ( .A(n682), .B(n641), .C(n599), .D(n716), .Z(n403) );
  IVI U597 ( .A(n403), .Z(n514) );
  IVI U598 ( .A(r1[14]), .Z(n462) );
  ND2I U599 ( .A(n200), .B(n462), .Z(n756) );
  IVI U600 ( .A(r1[13]), .Z(n441) );
  ND2I U601 ( .A(n333), .B(n441), .Z(n719) );
  IVI U602 ( .A(r1[12]), .Z(n439) );
  ND2I U603 ( .A(n179), .B(n439), .Z(n678) );
  IVI U604 ( .A(r1[15]), .Z(n500) );
  ND2I U605 ( .A(n170), .B(n500), .Z(n794) );
  NR2I U606 ( .A(r1[26]), .B(n205), .Z(n406) );
  ND2I U607 ( .A(n125), .B(n924), .Z(n914) );
  ND2I U608 ( .A(n172), .B(n44), .Z(n404) );
  ND2I U609 ( .A(n914), .B(n404), .Z(n405) );
  NR2I U610 ( .A(n406), .B(n75), .Z(n407) );
  ND2I U611 ( .A(n326), .B(n942), .Z(n950) );
  ND2I U612 ( .A(n407), .B(n950), .Z(n670) );
  ND2I U613 ( .A(n48), .B(n31), .Z(n970) );
  IVI U614 ( .A(r1[22]), .Z(n490) );
  ND2I U615 ( .A(n202), .B(n490), .Z(n916) );
  IVI U616 ( .A(r1[21]), .Z(n489) );
  ND2I U617 ( .A(n328), .B(n489), .Z(n877) );
  ND2I U618 ( .A(n179), .B(n51), .Z(n837) );
  IVI U619 ( .A(r1[23]), .Z(n487) );
  ND2I U620 ( .A(n168), .B(n487), .Z(n948) );
  IVI U621 ( .A(r1[29]), .Z(n1008) );
  IVI U622 ( .A(r1[31]), .Z(n1050) );
  ND2I U623 ( .A(n409), .B(n408), .Z(n995) );
  ND2I U624 ( .A(n370), .B(n375), .Z(n971) );
  IVI U625 ( .A(r1[18]), .Z(n801) );
  ND2I U626 ( .A(n271), .B(n801), .Z(n839) );
  IVI U627 ( .A(r1[17]), .Z(n499) );
  ND2I U628 ( .A(n74), .B(n499), .Z(n796) );
  ND2I U629 ( .A(n261), .B(n49), .Z(n754) );
  IVI U630 ( .A(r1[19]), .Z(n491) );
  ND2I U631 ( .A(n172), .B(n491), .Z(n875) );
  ND2I U632 ( .A(n411), .B(n410), .Z(n412) );
  AO4 U633 ( .A(r1[0]), .B(n288), .C(r1[1]), .D(n177), .Z(n413) );
  AO6 U634 ( .A(n266), .B(n466), .C(n413), .Z(n414) );
  ND2I U635 ( .A(n994), .B(n30), .Z(n1062) );
  ND2I U636 ( .A(n203), .B(n37), .Z(n603) );
  ND2I U637 ( .A(n172), .B(n208), .Z(n638) );
  AO3 U638 ( .A(n231), .B(n314), .C(n603), .D(n638), .Z(n415) );
  IVI U639 ( .A(n415), .Z(n513) );
  ND2I U640 ( .A(n953), .B(n216), .Z(n1068) );
  AO7 U641 ( .A(r1[1]), .B(n355), .C(n365), .Z(n428) );
  MUX21L U642 ( .A(n523), .B(n478), .S(n124), .Z(n427) );
  ND2I U643 ( .A(n427), .B(n232), .Z(n698) );
  IVI U644 ( .A(n698), .Z(n785) );
  AO2 U645 ( .A(n266), .B(n428), .C(n308), .D(n785), .Z(n453) );
  NR2I U646 ( .A(r1[27]), .B(n207), .Z(n430) );
  ND2I U647 ( .A(n171), .B(n42), .Z(n1053) );
  ND2I U648 ( .A(n160), .B(n942), .Z(n930) );
  ND2I U649 ( .A(n1053), .B(n930), .Z(n429) );
  NR2I U650 ( .A(n430), .B(n429), .Z(n431) );
  IVI U651 ( .A(r1[26]), .Z(n1006) );
  ND2I U652 ( .A(n326), .B(n1006), .Z(n967) );
  ND2I U653 ( .A(n431), .B(n967), .Z(n619) );
  ND2I U654 ( .A(n311), .B(n619), .Z(n434) );
  ND2I U655 ( .A(n63), .B(n687), .Z(n433) );
  AN2I U656 ( .A(n434), .B(n433), .Z(n436) );
  ND2I U657 ( .A(n203), .B(n491), .Z(n860) );
  ND2I U658 ( .A(n74), .B(n801), .Z(n818) );
  ND2I U659 ( .A(n292), .B(n499), .Z(n774) );
  ND2I U660 ( .A(n171), .B(n51), .Z(n892) );
  ND2I U661 ( .A(n202), .B(n487), .Z(n932) );
  ND2I U662 ( .A(n327), .B(n490), .Z(n894) );
  ND2I U663 ( .A(n229), .B(n489), .Z(n858) );
  ND2I U664 ( .A(n169), .B(n924), .Z(n965) );
  ND2I U665 ( .A(n612), .B(n378), .Z(n435) );
  ND2I U666 ( .A(n436), .B(n435), .Z(n772) );
  AO4 U667 ( .A(n291), .B(n523), .C(n330), .D(n542), .Z(n437) );
  AO6 U668 ( .A(n266), .B(n315), .C(n437), .Z(n438) );
  AO4 U669 ( .A(n216), .B(n772), .C(n438), .D(n1062), .Z(n447) );
  ND2I U670 ( .A(n202), .B(n657), .Z(n697) );
  ND2I U671 ( .A(n328), .B(n695), .Z(n659) );
  ND2I U672 ( .A(n160), .B(n680), .Z(n622) );
  ND2I U673 ( .A(n173), .B(n439), .Z(n739) );
  IVI U674 ( .A(n440), .Z(n533) );
  ND2I U675 ( .A(n200), .B(n500), .Z(n776) );
  ND2I U676 ( .A(n74), .B(n462), .Z(n742) );
  ND2I U677 ( .A(n167), .B(n49), .Z(n816) );
  ND4 U678 ( .A(n776), .B(n742), .C(n237), .D(n816), .Z(n442) );
  IVI U679 ( .A(n442), .Z(n531) );
  AO2 U680 ( .A(n38), .B(n326), .C(n107), .D(n200), .Z(n444) );
  AO2 U681 ( .A(n19), .B(n173), .C(r1[5]), .D(n180), .Z(n443) );
  ND2I U682 ( .A(n444), .B(n443), .Z(n532) );
  IVI U683 ( .A(n532), .Z(n445) );
  AO4 U684 ( .A(n615), .B(n1060), .C(n445), .D(n1068), .Z(n446) );
  AO7 U685 ( .A(n447), .B(n446), .C(n310), .Z(n452) );
  MUX21L U686 ( .A(n364), .B(n347), .S(n231), .Z(n448) );
  ND2I U687 ( .A(n448), .B(n365), .Z(n449) );
  AO2 U688 ( .A(r1[1]), .B(n449), .C(N193), .D(n39), .Z(n451) );
  ND2I U689 ( .A(N32), .B(n35), .Z(n450) );
  AO7 U690 ( .A(n267), .B(n355), .C(n365), .Z(n456) );
  IVI U691 ( .A(n181), .Z(n455) );
  AO2 U692 ( .A(n48), .B(n456), .C(n308), .D(n455), .Z(n477) );
  ND2I U693 ( .A(n173), .B(n1008), .Z(n558) );
  ND2I U694 ( .A(n292), .B(n1006), .Z(n949) );
  ND2I U695 ( .A(n326), .B(n487), .Z(n917) );
  ND2I U696 ( .A(n200), .B(n924), .Z(n951) );
  ND2I U697 ( .A(n169), .B(n942), .Z(n559) );
  ND2I U698 ( .A(n125), .B(n490), .Z(n876) );
  AO2 U699 ( .A(n311), .B(n708), .C(n953), .D(n709), .Z(n459) );
  ND2I U700 ( .A(n457), .B(n232), .Z(n1033) );
  ND2I U701 ( .A(n331), .B(n491), .Z(n840) );
  ND2I U702 ( .A(n202), .B(n51), .Z(n878) );
  ND2I U703 ( .A(n171), .B(n489), .Z(n915) );
  ND2I U704 ( .A(n261), .B(n801), .Z(n795) );
  AO2 U705 ( .A(n63), .B(n1033), .C(n994), .D(n550), .Z(n458) );
  ND2I U706 ( .A(n459), .B(n458), .Z(n802) );
  AO2 U707 ( .A(n241), .B(n326), .C(n293), .D(n203), .Z(n461) );
  AO2 U708 ( .A(r1[13]), .B(n109), .C(n258), .D(n102), .Z(n460) );
  ND2I U709 ( .A(n461), .B(n460), .Z(n553) );
  ND2I U710 ( .A(n333), .B(n500), .Z(n755) );
  ND2I U711 ( .A(n200), .B(n49), .Z(n797) );
  ND2I U712 ( .A(n171), .B(n499), .Z(n838) );
  ND2I U713 ( .A(n72), .B(n462), .Z(n715) );
  ND4 U714 ( .A(n755), .B(n797), .C(n838), .D(n715), .Z(n463) );
  IVI U715 ( .A(n463), .Z(n551) );
  AO4 U716 ( .A(n216), .B(n802), .C(n1060), .D(n632), .Z(n471) );
  AO2 U717 ( .A(n107), .B(n327), .C(n19), .D(n200), .Z(n465) );
  AO2 U718 ( .A(n259), .B(n109), .C(n38), .D(n240), .Z(n464) );
  ND2I U719 ( .A(n465), .B(n464), .Z(n552) );
  IVI U720 ( .A(n552), .Z(n469) );
  IVI U721 ( .A(n466), .Z(n467) );
  AO4 U722 ( .A(n469), .B(n1068), .C(n468), .D(n1062), .Z(n470) );
  AO7 U723 ( .A(n471), .B(n470), .C(n310), .Z(n476) );
  MUX21L U724 ( .A(n364), .B(n346), .S(n48), .Z(n472) );
  ND2I U725 ( .A(n472), .B(n365), .Z(n473) );
  AO2 U726 ( .A(n267), .B(n473), .C(N194), .D(n39), .Z(n475) );
  ND2I U727 ( .A(N33), .B(n35), .Z(n474) );
  AO7 U728 ( .A(n34), .B(n355), .C(n365), .Z(n481) );
  ND2I U729 ( .A(n480), .B(n479), .Z(n744) );
  IVI U730 ( .A(n233), .Z(n828) );
  AO2 U731 ( .A(n373), .B(n481), .C(n308), .D(n828), .Z(n511) );
  ND2I U732 ( .A(n202), .B(n1008), .Z(n1055) );
  ND2I U733 ( .A(n261), .B(n44), .Z(n966) );
  IVI U734 ( .A(n966), .Z(n482) );
  IVI U735 ( .A(n484), .Z(n583) );
  IVI U736 ( .A(n648), .Z(n974) );
  NR2I U737 ( .A(n209), .B(n175), .Z(n486) );
  ND2I U738 ( .A(n271), .B(n942), .Z(n968) );
  ND2I U739 ( .A(n326), .B(n924), .Z(n933) );
  ND2I U740 ( .A(n968), .B(n933), .Z(n485) );
  NR2I U741 ( .A(n486), .B(n485), .Z(n488) );
  ND2I U742 ( .A(n229), .B(n487), .Z(n893) );
  ND2I U743 ( .A(n488), .B(n893), .Z(n582) );
  ND2I U744 ( .A(n327), .B(n51), .Z(n861) );
  ND2I U745 ( .A(n201), .B(n489), .Z(n895) );
  ND2I U746 ( .A(n170), .B(n490), .Z(n931) );
  ND2I U747 ( .A(n179), .B(n491), .Z(n817) );
  ND4 U748 ( .A(n861), .B(n895), .C(n931), .D(n817), .Z(n575) );
  IVI U749 ( .A(r1[5]), .Z(n601) );
  AO4 U750 ( .A(n174), .B(n37), .C(n204), .D(n601), .Z(n493) );
  AO6 U751 ( .A(n315), .B(n232), .C(n493), .Z(n495) );
  AO2 U752 ( .A(n293), .B(n331), .C(r1[13]), .D(n203), .Z(n498) );
  AO2 U753 ( .A(n270), .B(n109), .C(n241), .D(n102), .Z(n497) );
  ND2I U754 ( .A(n498), .B(n497), .Z(n577) );
  ND2I U755 ( .A(n327), .B(n49), .Z(n775) );
  ND2I U756 ( .A(n203), .B(n499), .Z(n819) );
  ND2I U757 ( .A(n170), .B(n801), .Z(n859) );
  ND2I U758 ( .A(n229), .B(n500), .Z(n738) );
  AO2 U759 ( .A(n19), .B(n327), .C(n259), .D(n202), .Z(n502) );
  AO2 U760 ( .A(n258), .B(n109), .C(n107), .D(n97), .Z(n501) );
  ND2I U761 ( .A(n502), .B(n501), .Z(n576) );
  IVI U762 ( .A(n576), .Z(n503) );
  AO4 U763 ( .A(n1060), .B(n653), .C(n503), .D(n1068), .Z(n504) );
  AO7 U764 ( .A(n505), .B(n504), .C(n310), .Z(n510) );
  MUX21L U765 ( .A(n364), .B(n347), .S(n373), .Z(n506) );
  ND2I U766 ( .A(n506), .B(n365), .Z(n507) );
  AO2 U767 ( .A(n34), .B(n507), .C(N195), .D(n39), .Z(n509) );
  ND2I U768 ( .A(N34), .B(n35), .Z(n508) );
  AO7 U769 ( .A(n55), .B(n355), .C(n365), .Z(n517) );
  MUX21L U770 ( .A(n87), .B(n178), .S(n344), .Z(n674) );
  AO2 U771 ( .A(n514), .B(n953), .C(n513), .D(n994), .Z(n515) );
  AO7 U772 ( .A(n674), .B(n31), .C(n515), .Z(n516) );
  MUX21L U773 ( .A(n362), .B(n346), .S(n29), .Z(n518) );
  ND2I U774 ( .A(n518), .B(n366), .Z(n522) );
  ND2I U775 ( .A(n313), .B(n318), .Z(n729) );
  IVI U776 ( .A(n729), .Z(n667) );
  IVI U777 ( .A(n519), .Z(n672) );
  IVI U778 ( .A(n162), .Z(n521) );
  AO2 U779 ( .A(n55), .B(n522), .C(n667), .D(n521), .Z(n529) );
  AO2 U780 ( .A(n173), .B(n523), .C(n119), .D(n99), .Z(n524) );
  ND2I U781 ( .A(n525), .B(n524), .Z(n604) );
  IVI U782 ( .A(n604), .Z(n759) );
  IVI U783 ( .A(n526), .Z(n849) );
  AO2 U784 ( .A(n281), .B(n849), .C(N196), .D(n39), .Z(n528) );
  ND2I U785 ( .A(N35), .B(n35), .Z(n527) );
  AO7 U786 ( .A(r1[5]), .B(n355), .C(n366), .Z(n536) );
  MUX21L U787 ( .A(n531), .B(n80), .S(n344), .Z(n690) );
  AO2 U788 ( .A(n533), .B(n953), .C(n994), .D(n532), .Z(n534) );
  AO7 U789 ( .A(n690), .B(n31), .C(n534), .Z(n535) );
  MUX21L U790 ( .A(n362), .B(n347), .S(n224), .Z(n537) );
  ND2I U791 ( .A(n537), .B(n366), .Z(n541) );
  IVI U792 ( .A(n619), .Z(n538) );
  MUX21L U793 ( .A(n82), .B(n538), .S(n344), .Z(n689) );
  ND2I U794 ( .A(n539), .B(n661), .Z(n870) );
  IVI U795 ( .A(n870), .Z(n540) );
  AO2 U796 ( .A(r1[5]), .B(n541), .C(n667), .D(n540), .Z(n548) );
  ND2I U797 ( .A(n544), .B(n543), .Z(n780) );
  MUX21L U798 ( .A(n780), .B(n698), .S(n344), .Z(n545) );
  AO2 U799 ( .A(n83), .B(n300), .C(N197), .D(n39), .Z(n547) );
  ND2I U800 ( .A(N36), .B(n35), .Z(n546) );
  AO7 U801 ( .A(n38), .B(n356), .C(n366), .Z(n556) );
  IVI U802 ( .A(n550), .Z(n630) );
  MUX21L U803 ( .A(n551), .B(n630), .S(n344), .Z(n710) );
  AO2 U804 ( .A(n953), .B(n553), .C(n994), .D(n552), .Z(n554) );
  AO7 U805 ( .A(n710), .B(n375), .C(n554), .Z(n555) );
  MUX21L U806 ( .A(n362), .B(n346), .S(n147), .Z(n557) );
  ND2I U807 ( .A(n557), .B(n366), .Z(n566) );
  ND4 U808 ( .A(n953), .B(n949), .C(n558), .D(n5), .Z(n563) );
  IVI U809 ( .A(n559), .Z(n560) );
  NR2I U810 ( .A(n560), .B(n971), .Z(n561) );
  ND4 U811 ( .A(n561), .B(n951), .C(n917), .D(n7), .Z(n562) );
  AO3 U812 ( .A(n376), .B(n1033), .C(n563), .D(n562), .Z(n564) );
  ND2I U813 ( .A(n564), .B(n661), .Z(n887) );
  IVI U814 ( .A(n887), .Z(n565) );
  AO2 U815 ( .A(n38), .B(n566), .C(n667), .D(n565), .Z(n573) );
  ND2I U816 ( .A(n568), .B(n567), .Z(n805) );
  ND2I U817 ( .A(n569), .B(n376), .Z(n570) );
  IVI U818 ( .A(n570), .Z(n880) );
  AO2 U819 ( .A(n880), .B(n301), .C(N198), .D(n39), .Z(n572) );
  ND2I U820 ( .A(N37), .B(n35), .Z(n571) );
  AO7 U821 ( .A(n107), .B(n356), .C(n366), .Z(n580) );
  AO2 U822 ( .A(n953), .B(n577), .C(n994), .D(n576), .Z(n578) );
  AO7 U823 ( .A(n733), .B(n376), .C(n578), .Z(n579) );
  MUX21L U824 ( .A(n361), .B(n347), .S(n251), .Z(n581) );
  ND2I U825 ( .A(n581), .B(n366), .Z(n584) );
  IVI U826 ( .A(n582), .Z(n651) );
  MUX21L U827 ( .A(n651), .B(n583), .S(n344), .Z(n732) );
  ND2I U828 ( .A(n56), .B(n370), .Z(n1070) );
  AO2 U829 ( .A(n107), .B(n584), .C(n667), .D(n900), .Z(n590) );
  ND2I U830 ( .A(n586), .B(n585), .Z(n824) );
  AO2 U831 ( .A(n26), .B(n300), .C(N199), .D(n39), .Z(n589) );
  ND2I U832 ( .A(N38), .B(n35), .Z(n588) );
  AO7 U833 ( .A(n19), .B(n356), .C(n366), .Z(n595) );
  AO2 U834 ( .A(n178), .B(n311), .C(n672), .D(n63), .Z(n592) );
  AO7 U835 ( .A(n373), .B(n593), .C(n592), .Z(n594) );
  AO2 U836 ( .A(n196), .B(n595), .C(n342), .D(n594), .Z(n611) );
  MUX21L U837 ( .A(n361), .B(n346), .S(n196), .Z(n596) );
  ND2I U838 ( .A(n596), .B(n366), .Z(n598) );
  AO2 U839 ( .A(n25), .B(n598), .C(n667), .D(n84), .Z(n610) );
  IVI U840 ( .A(n599), .Z(n600) );
  ND2I U841 ( .A(N39), .B(n35), .Z(n608) );
  AO7 U842 ( .A(n259), .B(n357), .C(n367), .Z(n614) );
  IVI U843 ( .A(n612), .Z(n613) );
  AO2 U844 ( .A(n23), .B(n614), .C(n305), .D(n613), .Z(n628) );
  IVI U845 ( .A(n615), .Z(n618) );
  MUX21L U846 ( .A(n362), .B(n347), .S(n23), .Z(n616) );
  ND2I U847 ( .A(n616), .B(n367), .Z(n617) );
  AO2 U848 ( .A(n66), .B(n618), .C(n259), .D(n617), .Z(n627) );
  IVI U849 ( .A(n694), .Z(n864) );
  AO2 U850 ( .A(n48), .B(n780), .C(n373), .D(n698), .Z(n623) );
  AO3 U851 ( .A(n864), .B(n971), .C(n661), .D(n623), .Z(n624) );
  IVI U852 ( .A(n624), .Z(n939) );
  AO2 U853 ( .A(n667), .B(n85), .C(n939), .D(n300), .Z(n626) );
  AO7 U854 ( .A(n258), .B(n357), .C(n367), .Z(n634) );
  IVI U855 ( .A(n709), .Z(n629) );
  AO2 U856 ( .A(n630), .B(n311), .C(n629), .D(n63), .Z(n631) );
  AO7 U857 ( .A(n373), .B(n632), .C(n631), .Z(n633) );
  AO2 U858 ( .A(n218), .B(n634), .C(n341), .D(n633), .Z(n647) );
  MUX21L U859 ( .A(n362), .B(n346), .S(n218), .Z(n635) );
  ND2I U860 ( .A(n635), .B(n367), .Z(n637) );
  AO2 U861 ( .A(n258), .B(n637), .C(n667), .D(n88), .Z(n646) );
  IVI U862 ( .A(n638), .Z(n639) );
  IVI U863 ( .A(n148), .Z(n881) );
  IVI U864 ( .A(n643), .Z(n958) );
  AO2 U865 ( .A(n958), .B(n96), .C(N202), .D(n39), .Z(n645) );
  ND2I U866 ( .A(N41), .B(n35), .Z(n644) );
  ND4 U867 ( .A(n647), .B(n646), .C(n645), .D(n644), .Z(result[10]) );
  NR2I U868 ( .A(n648), .B(n729), .Z(n650) );
  AO7 U869 ( .A(n241), .B(n357), .C(n367), .Z(n649) );
  AO2 U870 ( .A(n650), .B(n378), .C(r2[11]), .D(n649), .Z(n666) );
  AO2 U871 ( .A(n58), .B(n311), .C(n651), .D(n63), .Z(n652) );
  AO7 U872 ( .A(n373), .B(n653), .C(n652), .Z(n656) );
  MUX21L U873 ( .A(n363), .B(n347), .S(r2[11]), .Z(n654) );
  ND2I U874 ( .A(n654), .B(n367), .Z(n655) );
  AO2 U875 ( .A(n341), .B(n656), .C(n241), .D(n655), .Z(n665) );
  IVI U876 ( .A(n132), .Z(n902) );
  IVI U877 ( .A(n662), .Z(n977) );
  AO2 U878 ( .A(n977), .B(n300), .C(N203), .D(n39), .Z(n664) );
  ND2I U879 ( .A(N42), .B(n35), .Z(n663) );
  ND4 U880 ( .A(n666), .B(n665), .C(n664), .D(n663), .Z(result[11]) );
  AO7 U881 ( .A(n293), .B(n355), .C(n367), .Z(n669) );
  IVI U882 ( .A(n995), .Z(n668) );
  AO2 U883 ( .A(n298), .B(n669), .C(n309), .D(n668), .Z(n686) );
  IVI U884 ( .A(n187), .Z(n671) );
  AO2 U885 ( .A(n672), .B(n311), .C(n671), .D(n63), .Z(n673) );
  AO7 U886 ( .A(n373), .B(n674), .C(n673), .Z(n677) );
  MUX21L U887 ( .A(n363), .B(n346), .S(n298), .Z(n675) );
  ND2I U888 ( .A(n675), .B(n367), .Z(n676) );
  AO2 U889 ( .A(n340), .B(n677), .C(n293), .D(n676), .Z(n685) );
  IVI U890 ( .A(n678), .Z(n679) );
  AO2 U891 ( .A(n273), .B(n96), .C(N204), .D(n39), .Z(n684) );
  ND2I U892 ( .A(N43), .B(n35), .Z(n683) );
  ND4 U893 ( .A(n686), .B(n685), .C(n684), .D(n683), .Z(result[12]) );
  AO7 U894 ( .A(r1[13]), .B(n355), .C(n367), .Z(n688) );
  IVI U895 ( .A(n687), .Z(n1018) );
  AO2 U896 ( .A(n211), .B(n688), .C(n309), .D(n1018), .Z(n705) );
  IVI U897 ( .A(n689), .Z(n692) );
  IVI U898 ( .A(n690), .Z(n691) );
  AO2 U899 ( .A(n305), .B(n692), .C(n66), .D(n691), .Z(n704) );
  MUX21L U900 ( .A(n364), .B(n347), .S(n211), .Z(n693) );
  ND2I U901 ( .A(n693), .B(n366), .Z(n701) );
  AO2 U902 ( .A(n311), .B(n780), .C(n953), .D(n694), .Z(n700) );
  AO2 U903 ( .A(n63), .B(n698), .C(n994), .D(n863), .Z(n699) );
  AO2 U904 ( .A(n21), .B(n701), .C(n90), .D(n300), .Z(n703) );
  AO7 U905 ( .A(n270), .B(n355), .C(n367), .Z(n707) );
  IVI U906 ( .A(n1033), .Z(n706) );
  AO2 U907 ( .A(r2[14]), .B(n707), .C(n309), .D(n706), .Z(n728) );
  IVI U908 ( .A(n710), .Z(n711) );
  AO2 U909 ( .A(n305), .B(n712), .C(n306), .D(n711), .Z(n727) );
  MUX21L U910 ( .A(n364), .B(n346), .S(r2[14]), .Z(n713) );
  ND2I U911 ( .A(n713), .B(n367), .Z(n724) );
  NR2I U912 ( .A(n293), .B(n206), .Z(n718) );
  ND2I U913 ( .A(n716), .B(n715), .Z(n717) );
  NR2I U914 ( .A(n718), .B(n717), .Z(n720) );
  ND2I U915 ( .A(n720), .B(n719), .Z(n879) );
  ND2I U916 ( .A(n722), .B(n721), .Z(n723) );
  IVI U917 ( .A(n723), .Z(n1041) );
  AO2 U918 ( .A(n270), .B(n724), .C(n301), .D(n1041), .Z(n726) );
  NR2I U919 ( .A(n1070), .B(n729), .Z(n731) );
  AO7 U920 ( .A(r1[15]), .B(n355), .C(n366), .Z(n730) );
  AO2 U921 ( .A(n731), .B(n378), .C(n138), .D(n730), .Z(n752) );
  IVI U922 ( .A(n732), .Z(n735) );
  IVI U923 ( .A(n733), .Z(n734) );
  AO2 U924 ( .A(n305), .B(n735), .C(n306), .D(n734), .Z(n751) );
  MUX21L U925 ( .A(n364), .B(n347), .S(n138), .Z(n736) );
  ND2I U926 ( .A(n736), .B(n366), .Z(n748) );
  NR2I U927 ( .A(r1[13]), .B(n204), .Z(n741) );
  ND2I U928 ( .A(n739), .B(n738), .Z(n740) );
  NR2I U929 ( .A(n741), .B(n740), .Z(n743) );
  ND2I U930 ( .A(n743), .B(n742), .Z(n898) );
  ND2I U931 ( .A(n746), .B(n745), .Z(n1065) );
  IVI U932 ( .A(n1065), .Z(n747) );
  AO2 U933 ( .A(r1[15]), .B(n748), .C(n747), .D(n300), .Z(n750) );
  ND2I U934 ( .A(N208), .B(n39), .Z(n771) );
  IVI U935 ( .A(n753), .Z(n852) );
  ND2I U936 ( .A(n989), .B(n311), .Z(n899) );
  IVI U937 ( .A(n899), .Z(n843) );
  NR2I U938 ( .A(n121), .B(n757), .Z(n841) );
  IVI U939 ( .A(n758), .Z(n844) );
  IVI U940 ( .A(n919), .Z(n760) );
  ND2I U941 ( .A(n126), .B(n63), .Z(n806) );
  ND2I U942 ( .A(n313), .B(n317), .Z(n783) );
  NR2I U943 ( .A(n783), .B(n761), .Z(n763) );
  AO7 U944 ( .A(n50), .B(n357), .C(n367), .Z(n762) );
  AO2 U945 ( .A(n763), .B(n31), .C(n155), .D(n762), .Z(n766) );
  MUX21L U946 ( .A(n354), .B(n345), .S(n156), .Z(n764) );
  AO7 U947 ( .A(n28), .B(n764), .C(n50), .Z(n765) );
  ND2I U948 ( .A(n771), .B(n770), .Z(result[16]) );
  ND2I U949 ( .A(N209), .B(n39), .Z(n793) );
  IVI U950 ( .A(n772), .Z(n773) );
  IVI U951 ( .A(n774), .Z(n778) );
  NR2I U952 ( .A(n778), .B(n777), .Z(n862) );
  IVI U953 ( .A(n863), .Z(n779) );
  IVI U954 ( .A(n936), .Z(n782) );
  IVI U955 ( .A(n780), .Z(n781) );
  ND2I U956 ( .A(n1020), .B(n994), .Z(n808) );
  IVI U957 ( .A(n808), .Z(n827) );
  AO7 U958 ( .A(r1[17]), .B(n351), .C(n365), .Z(n784) );
  AO2 U959 ( .A(n785), .B(n827), .C(n214), .D(n784), .Z(n788) );
  MUX21L U960 ( .A(n353), .B(n345), .S(n214), .Z(n786) );
  AO7 U961 ( .A(n28), .B(n786), .C(r1[17]), .Z(n787) );
  ND2I U962 ( .A(n793), .B(n792), .Z(result[17]) );
  ND2I U963 ( .A(N210), .B(n39), .Z(n815) );
  IVI U964 ( .A(n879), .Z(n798) );
  MUX21L U965 ( .A(n165), .B(n798), .S(n344), .Z(n955) );
  MUX21L U966 ( .A(n364), .B(n346), .S(n166), .Z(n799) );
  ND2I U967 ( .A(n799), .B(n366), .Z(n800) );
  AO2 U968 ( .A(n276), .B(n800), .C(n881), .D(n843), .Z(n812) );
  AO6 U969 ( .A(n362), .B(n801), .C(n368), .Z(n804) );
  IVI U970 ( .A(r2[18]), .Z(n803) );
  NR2I U971 ( .A(n810), .B(n809), .Z(n811) );
  ND2I U972 ( .A(n815), .B(n814), .Z(result[18]) );
  ND2I U973 ( .A(N211), .B(n39), .Z(n836) );
  ND4 U974 ( .A(n819), .B(n818), .C(n817), .D(n816), .Z(n820) );
  IVI U975 ( .A(n820), .Z(n896) );
  IVI U976 ( .A(n898), .Z(n821) );
  MUX21L U977 ( .A(n896), .B(n821), .S(n344), .Z(n822) );
  IVI U978 ( .A(n822), .Z(n973) );
  IVI U979 ( .A(n198), .Z(n825) );
  AO7 U980 ( .A(r1[19]), .B(n353), .C(n366), .Z(n826) );
  AO2 U981 ( .A(n828), .B(n827), .C(n41), .D(n826), .Z(n831) );
  MUX21L U982 ( .A(n353), .B(n345), .S(r2[19]), .Z(n829) );
  AO7 U983 ( .A(n28), .B(n829), .C(r1[19]), .Z(n830) );
  ND2I U984 ( .A(n836), .B(n835), .Z(result[19]) );
  ND2I U985 ( .A(N212), .B(n39), .Z(n857) );
  MUX21L U986 ( .A(n89), .B(n841), .S(n344), .Z(n990) );
  MUX21L U987 ( .A(n364), .B(n347), .S(n189), .Z(n842) );
  ND2I U988 ( .A(n842), .B(n27), .Z(n845) );
  AO6 U989 ( .A(n361), .B(n51), .C(n369), .Z(n848) );
  ND2I U990 ( .A(n857), .B(n856), .Z(result[20]) );
  ND2I U991 ( .A(N213), .B(n39), .Z(n874) );
  AO7 U992 ( .A(n22), .B(n359), .C(n27), .Z(n867) );
  MUX21L U993 ( .A(n364), .B(n346), .S(n194), .Z(n865) );
  ND2I U994 ( .A(n865), .B(n27), .Z(n866) );
  AO2 U995 ( .A(n194), .B(n867), .C(n22), .D(n866), .Z(n868) );
  ND2I U996 ( .A(n874), .B(n873), .Z(result[21]) );
  ND2I U997 ( .A(N214), .B(n39), .Z(n891) );
  AO7 U998 ( .A(r1[22]), .B(n358), .C(n27), .Z(n884) );
  MUX21L U999 ( .A(n364), .B(n347), .S(n127), .Z(n882) );
  ND2I U1000 ( .A(n882), .B(n27), .Z(n883) );
  AO2 U1001 ( .A(n127), .B(n884), .C(r1[22]), .D(n883), .Z(n885) );
  ND2I U1002 ( .A(n891), .B(n890), .Z(result[22]) );
  ND2I U1003 ( .A(N215), .B(n39), .Z(n912) );
  IVI U1004 ( .A(n969), .Z(n897) );
  IVI U1005 ( .A(n900), .Z(n908) );
  AO7 U1006 ( .A(r1[23]), .B(n358), .C(n27), .Z(n905) );
  MUX21L U1007 ( .A(n364), .B(n346), .S(r2[23]), .Z(n903) );
  ND2I U1008 ( .A(n903), .B(n27), .Z(n904) );
  AO2 U1009 ( .A(r2[23]), .B(n905), .C(r1[23]), .D(n904), .Z(n906) );
  ND2I U1010 ( .A(n912), .B(n911), .Z(result[23]) );
  ND2I U1011 ( .A(N216), .B(n39), .Z(n928) );
  MUX21L U1012 ( .A(n353), .B(n345), .S(r2[24]), .Z(n913) );
  NR2I U1013 ( .A(n28), .B(n913), .Z(n925) );
  AO7 U1014 ( .A(r1[24]), .B(n358), .C(n27), .Z(n921) );
  ND2I U1015 ( .A(n928), .B(n927), .Z(result[24]) );
  ND2I U1016 ( .A(N217), .B(n39), .Z(n946) );
  MUX21L U1017 ( .A(n353), .B(n345), .S(n152), .Z(n929) );
  NR2I U1018 ( .A(n369), .B(n929), .Z(n943) );
  AO7 U1019 ( .A(r1[25]), .B(n359), .C(n27), .Z(n938) );
  IVI U1020 ( .A(n1013), .Z(n934) );
  ND2I U1021 ( .A(n946), .B(n945), .Z(result[25]) );
  ND2I U1022 ( .A(N218), .B(n39), .Z(n964) );
  MUX21L U1023 ( .A(n352), .B(n345), .S(r2[26]), .Z(n947) );
  NR2I U1024 ( .A(n369), .B(n947), .Z(n961) );
  AO7 U1025 ( .A(n209), .B(n359), .C(n367), .Z(n957) );
  IVI U1026 ( .A(n1035), .Z(n952) );
  ND2I U1027 ( .A(n964), .B(n963), .Z(result[26]) );
  ND2I U1028 ( .A(N219), .B(n39), .Z(n985) );
  ND4 U1029 ( .A(n968), .B(n967), .C(n966), .D(n965), .Z(n1051) );
  AO4 U1030 ( .A(n971), .B(n1051), .C(n970), .D(n969), .Z(n972) );
  AO6 U1031 ( .A(n373), .B(n973), .C(n972), .Z(n982) );
  AO7 U1032 ( .A(r1[27]), .B(n359), .C(n365), .Z(n975) );
  MUX21L U1033 ( .A(n364), .B(n347), .S(r2[27]), .Z(n976) );
  ND2I U1034 ( .A(n976), .B(n366), .Z(n978) );
  ND2I U1035 ( .A(n985), .B(n984), .Z(result[27]) );
  ND2I U1036 ( .A(N220), .B(n39), .Z(n1004) );
  AO2 U1037 ( .A(n45), .B(n327), .C(n209), .D(n201), .Z(n987) );
  AO2 U1038 ( .A(r1[25]), .B(n109), .C(n43), .D(n240), .Z(n986) );
  ND2I U1039 ( .A(n987), .B(n986), .Z(n988) );
  MUX21L U1040 ( .A(n988), .B(n86), .S(n344), .Z(n1001) );
  IVI U1041 ( .A(n990), .Z(n992) );
  AO7 U1042 ( .A(n43), .B(n356), .C(n366), .Z(n991) );
  MUX21L U1043 ( .A(n352), .B(n345), .S(r2[28]), .Z(n993) );
  NR2I U1044 ( .A(n369), .B(n993), .Z(n996) );
  ND2I U1045 ( .A(n296), .B(n994), .Z(n1032) );
  ND2I U1046 ( .A(n1004), .B(n1003), .Z(result[28]) );
  AO7 U1047 ( .A(n199), .B(n354), .C(n367), .Z(n1005) );
  ND2I U1048 ( .A(n182), .B(n1005), .Z(n1028) );
  ND2I U1049 ( .A(n307), .B(n81), .Z(n1027) );
  AO4 U1050 ( .A(n291), .B(n1008), .C(n175), .D(n101), .Z(n1012) );
  AO4 U1051 ( .A(n206), .B(n44), .C(n330), .D(n42), .Z(n1011) );
  NR2I U1052 ( .A(n1012), .B(n1011), .Z(n1014) );
  MUX21L U1053 ( .A(n1014), .B(n1013), .S(n48), .Z(n1015) );
  ND2I U1054 ( .A(n281), .B(n1015), .Z(n1026) );
  MUX21L U1055 ( .A(n351), .B(n345), .S(n182), .Z(n1017) );
  AO7 U1056 ( .A(n28), .B(n1017), .C(n199), .Z(n1025) );
  IVI U1057 ( .A(n1032), .Z(n1019) );
  ND2I U1058 ( .A(n1019), .B(n1018), .Z(n1024) );
  ND2I U1059 ( .A(n234), .B(n90), .Z(n1023) );
  ND2I U1060 ( .A(N60), .B(n35), .Z(n1022) );
  ND2I U1061 ( .A(N221), .B(n39), .Z(n1021) );
  ND8 U1062 ( .A(n1028), .B(n1027), .C(n1026), .D(n1025), .E(n1024), .F(n1023), 
        .G(n1022), .H(n1021), .Z(result[29]) );
  ND2I U1063 ( .A(N222), .B(n39), .Z(n1049) );
  MUX21L U1064 ( .A(n351), .B(n345), .S(r2[30]), .Z(n1031) );
  NR2I U1065 ( .A(n28), .B(n1031), .Z(n1034) );
  AO4 U1066 ( .A(n1034), .B(n1058), .C(n1033), .D(n1032), .Z(n1047) );
  AO6 U1067 ( .A(n362), .B(n1058), .C(n28), .Z(n1045) );
  AO2 U1068 ( .A(r1[29]), .B(n326), .C(n43), .D(n201), .Z(n1038) );
  AO2 U1069 ( .A(r1[27]), .B(n173), .C(r1[30]), .D(n97), .Z(n1037) );
  AO6 U1070 ( .A(n1038), .B(n1037), .C(n1062), .Z(n1039) );
  AO1P U1071 ( .A(n1041), .B(n29), .C(n1040), .D(n1039), .Z(n1043) );
  ND2I U1072 ( .A(n317), .B(n115), .Z(n1052) );
  AO4 U1073 ( .A(n1045), .B(n1044), .C(n1043), .D(n1052), .Z(n1046) );
  AO1P U1074 ( .A(N61), .B(n35), .C(n1047), .D(n1046), .Z(n1048) );
  ND2I U1075 ( .A(n1049), .B(n1048), .Z(result[30]) );
  ND2I U1076 ( .A(N223), .B(n39), .Z(n1080) );
  AO6 U1077 ( .A(n362), .B(n1050), .C(n28), .Z(n1077) );
  IVI U1078 ( .A(n1051), .Z(n1069) );
  IVI U1079 ( .A(n1052), .Z(n1067) );
  IVI U1080 ( .A(n1055), .Z(n1056) );
  AO1P U1081 ( .A(n333), .B(n1058), .C(n1057), .D(n1056), .Z(n1063) );
  IVI U1082 ( .A(n1059), .Z(n1061) );
  IVI U1083 ( .A(n1070), .Z(n1073) );
  MUX21L U1084 ( .A(n364), .B(n346), .S(n220), .Z(n1071) );
  ND2I U1085 ( .A(n1071), .B(n366), .Z(n1072) );
  ND2I U1086 ( .A(n1080), .B(n1079), .Z(result[31]) );
endmodule


module forward_stall ( gpr_wr_addr, m_gpr_wr_addr, mw_opcode, xm_opcode, xm_rt, 
        dx_gpr_rd_addr1, dx_rt, dx_isSLL_SRL, dx_opcode, fd_opcode, fd_funct, 
        fd_rs, fd_rt, gpr_rd_addr1, d_fwd_rs, d_fwd_rt, d_stall, 
        x_fwd_alu_src1, x_fwd_alu_src2, Port20 );
  input [4:0] gpr_wr_addr;
  input [4:0] m_gpr_wr_addr;
  input [5:0] mw_opcode;
  input [5:0] xm_opcode;
  input [4:0] xm_rt;
  input [4:0] dx_gpr_rd_addr1;
  input [4:0] dx_rt;
  input [5:0] dx_opcode;
  input [5:0] fd_opcode;
  input [5:0] fd_funct;
  input [4:0] fd_rs;
  input [4:0] fd_rt;
  input [4:0] gpr_rd_addr1;
  output [1:0] d_fwd_rs;
  output [1:0] d_fwd_rt;
  output [1:0] x_fwd_alu_src1;
  output [1:0] x_fwd_alu_src2;
  input dx_isSLL_SRL, Port20;
  output d_stall;
  wire   mw_opcode_3, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143;
  assign d_stall = 1'b0;
  assign mw_opcode_3 = mw_opcode[3];

  B2I U2 ( .A(fd_rt[4]), .Z1(n1), .Z2(n2) );
  IVDA U3 ( .A(fd_rt[3]), .Y(n3), .Z(n4) );
  IVDA U4 ( .A(fd_rt[2]), .Y(n5), .Z(n6) );
  IVI U5 ( .A(n27), .Z(n7) );
  ND2I U6 ( .A(n40), .B(n66), .Z(n8) );
  IVI U7 ( .A(m_gpr_wr_addr[3]), .Z(n9) );
  IVI U8 ( .A(fd_rs[0]), .Z(n12) );
  AN2I U9 ( .A(n85), .B(n113), .Z(n10) );
  AN2I U10 ( .A(n102), .B(n113), .Z(n11) );
  ENI U11 ( .A(n122), .B(n12), .Z(n129) );
  ND3P U12 ( .A(n94), .B(n95), .C(n11), .Z(n97) );
  IVI U13 ( .A(m_gpr_wr_addr[0]), .Z(n13) );
  ND2I U14 ( .A(n14), .B(n34), .Z(n15) );
  ND2I U15 ( .A(n15), .B(n33), .Z(d_fwd_rt[1]) );
  IVI U16 ( .A(n121), .Z(n14) );
  OR2I U17 ( .A(n8), .B(n53), .Z(n16) );
  OR2I U18 ( .A(n89), .B(n88), .Z(n17) );
  ND2I U19 ( .A(n16), .B(n17), .Z(x_fwd_alu_src2[1]) );
  ND2I U20 ( .A(n18), .B(n19), .Z(n22) );
  EOI U21 ( .A(dx_gpr_rd_addr1[3]), .B(n9), .Z(n18) );
  EOI U22 ( .A(dx_gpr_rd_addr1[1]), .B(n61), .Z(n19) );
  NR2I U23 ( .A(n21), .B(n54), .Z(n20) );
  ENI U24 ( .A(gpr_wr_addr[3]), .B(n79), .Z(n21) );
  ND2I U25 ( .A(n24), .B(n25), .Z(n23) );
  ENI U26 ( .A(gpr_wr_addr[2]), .B(dx_gpr_rd_addr1[2]), .Z(n24) );
  ENI U27 ( .A(n7), .B(dx_gpr_rd_addr1[1]), .Z(n25) );
  AN2I U28 ( .A(n20), .B(n87), .Z(n26) );
  AN2I U29 ( .A(n88), .B(n26), .Z(x_fwd_alu_src2[0]) );
  IVI U30 ( .A(gpr_wr_addr[1]), .Z(n27) );
  IVI U31 ( .A(n27), .Z(n28) );
  IVI U32 ( .A(gpr_wr_addr[2]), .Z(n29) );
  IVI U33 ( .A(n29), .Z(n30) );
  ND2I U34 ( .A(n140), .B(n139), .Z(n31) );
  IVI U35 ( .A(n122), .Z(n32) );
  NR2I U36 ( .A(n51), .B(n22), .Z(n98) );
  ND2I U37 ( .A(n118), .B(n117), .Z(n33) );
  IVI U38 ( .A(n120), .Z(n34) );
  NR3P U39 ( .A(n96), .B(n97), .C(n23), .Z(n101) );
  ND2I U40 ( .A(n36), .B(n125), .Z(n35) );
  EOI U41 ( .A(fd_rs[1]), .B(n61), .Z(n36) );
  OR2I U42 ( .A(n143), .B(n142), .Z(n37) );
  ND2I U43 ( .A(n37), .B(n31), .Z(d_fwd_rs[1]) );
  B3IP U44 ( .A(m_gpr_wr_addr[1]), .Z1(n61), .Z2(n60) );
  IVI U45 ( .A(n119), .Z(d_fwd_rt[0]) );
  IVI U46 ( .A(gpr_wr_addr[3]), .Z(n38) );
  IVI U47 ( .A(n38), .Z(n39) );
  ND4P U48 ( .A(n100), .B(n125), .C(n99), .D(n98), .Z(n104) );
  AN2I U49 ( .A(n67), .B(n68), .Z(n40) );
  AN4 U50 ( .A(n41), .B(n42), .C(n43), .D(n44), .Z(n117) );
  ENI U51 ( .A(n6), .B(n30), .Z(n41) );
  ENI U52 ( .A(gpr_wr_addr[0]), .B(n64), .Z(n42) );
  ENI U53 ( .A(n4), .B(n39), .Z(n43) );
  ENI U54 ( .A(n62), .B(n28), .Z(n44) );
  AN2I U55 ( .A(n120), .B(n52), .Z(n118) );
  AN4 U56 ( .A(n45), .B(n46), .C(n47), .D(n48), .Z(n139) );
  ENI U57 ( .A(fd_rs[2]), .B(n30), .Z(n45) );
  ENI U58 ( .A(fd_rs[0]), .B(gpr_wr_addr[0]), .Z(n46) );
  ENI U59 ( .A(fd_rs[3]), .B(n39), .Z(n47) );
  ENI U60 ( .A(fd_rs[1]), .B(n28), .Z(n48) );
  NR2I U61 ( .A(n56), .B(n35), .Z(n126) );
  ND2I U62 ( .A(n102), .B(n49), .Z(n50) );
  ND2I U63 ( .A(n50), .B(n103), .Z(x_fwd_alu_src1[1]) );
  IVI U64 ( .A(n104), .Z(n49) );
  ENI U65 ( .A(n124), .B(dx_gpr_rd_addr1[4]), .Z(n51) );
  ENI U66 ( .A(n93), .B(n78), .Z(n86) );
  NR3P U67 ( .A(n116), .B(n121), .C(n138), .Z(n52) );
  NR3P U68 ( .A(n110), .B(n109), .C(n108), .Z(n111) );
  IVI U69 ( .A(n20), .Z(n53) );
  ND2I U70 ( .A(n86), .B(n10), .Z(n54) );
  AN3 U71 ( .A(n58), .B(n57), .C(n113), .Z(n55) );
  AN2I U72 ( .A(n142), .B(n55), .Z(n140) );
  IVI U73 ( .A(n143), .Z(n57) );
  NR3P U74 ( .A(xm_opcode[5]), .B(n74), .C(n73), .Z(n76) );
  ENI U75 ( .A(n124), .B(fd_rs[4]), .Z(n56) );
  ENI U76 ( .A(fd_rs[4]), .B(gpr_wr_addr[4]), .Z(n58) );
  ENI U77 ( .A(dx_gpr_rd_addr1[3]), .B(gpr_wr_addr[3]), .Z(n95) );
  NR4 U78 ( .A(fd_opcode[4]), .B(fd_opcode[5]), .C(fd_opcode[1]), .D(
        fd_opcode[3]), .Z(n59) );
  NR3 U79 ( .A(dx_gpr_rd_addr1[2]), .B(dx_gpr_rd_addr1[1]), .C(
        dx_gpr_rd_addr1[0]), .Z(n92) );
  ND4P U80 ( .A(n129), .B(n128), .C(n127), .D(n126), .Z(n142) );
  AO3P U81 ( .A(dx_opcode[4]), .B(n84), .C(n83), .D(n82), .Z(n89) );
  IVI U82 ( .A(n63), .Z(n62) );
  IVI U83 ( .A(fd_rt[1]), .Z(n63) );
  IVI U84 ( .A(n65), .Z(n64) );
  IVI U85 ( .A(fd_rt[0]), .Z(n65) );
  ENI U86 ( .A(gpr_wr_addr[2]), .B(dx_rt[2]), .Z(n67) );
  ENI U87 ( .A(gpr_wr_addr[0]), .B(dx_rt[0]), .Z(n66) );
  ENI U88 ( .A(gpr_wr_addr[1]), .B(dx_rt[1]), .Z(n68) );
  ND2I U89 ( .A(n40), .B(n66), .Z(n90) );
  IVI U90 ( .A(n90), .Z(n87) );
  ENI U91 ( .A(m_gpr_wr_addr[2]), .B(dx_rt[2]), .Z(n70) );
  ENI U92 ( .A(m_gpr_wr_addr[4]), .B(dx_rt[4]), .Z(n69) );
  ND2I U93 ( .A(n70), .B(n69), .Z(n74) );
  ENI U94 ( .A(m_gpr_wr_addr[3]), .B(dx_rt[3]), .Z(n72) );
  ENI U95 ( .A(n60), .B(dx_rt[1]), .Z(n71) );
  ND2I U96 ( .A(n72), .B(n71), .Z(n73) );
  ENI U97 ( .A(dx_rt[0]), .B(n32), .Z(n75) );
  ND2I U98 ( .A(n76), .B(n75), .Z(n88) );
  IVI U99 ( .A(dx_rt[4]), .Z(n78) );
  IVI U100 ( .A(dx_rt[3]), .Z(n79) );
  IVI U101 ( .A(dx_opcode[3]), .Z(n77) );
  ND2I U102 ( .A(dx_opcode[5]), .B(n77), .Z(n84) );
  NR2I U103 ( .A(dx_rt[1]), .B(dx_rt[0]), .Z(n81) );
  IVI U104 ( .A(dx_rt[2]), .Z(n80) );
  ND4 U105 ( .A(n81), .B(n80), .C(n79), .D(n78), .Z(n83) );
  IVI U106 ( .A(dx_isSLL_SRL), .Z(n82) );
  IVI U107 ( .A(n89), .Z(n85) );
  ND2I U108 ( .A(mw_opcode_3), .B(mw_opcode[5]), .Z(n113) );
  NR2I U109 ( .A(dx_gpr_rd_addr1[3]), .B(dx_gpr_rd_addr1[4]), .Z(n91) );
  ND2I U110 ( .A(n92), .B(n91), .Z(n102) );
  IVI U111 ( .A(gpr_wr_addr[4]), .Z(n93) );
  EOI U112 ( .A(n93), .B(dx_gpr_rd_addr1[4]), .Z(n94) );
  EOI U113 ( .A(dx_gpr_rd_addr1[0]), .B(gpr_wr_addr[0]), .Z(n96) );
  IVI U114 ( .A(m_gpr_wr_addr[2]), .Z(n123) );
  EOI U115 ( .A(n123), .B(dx_gpr_rd_addr1[2]), .Z(n100) );
  IVI U116 ( .A(xm_opcode[5]), .Z(n125) );
  IVI U117 ( .A(m_gpr_wr_addr[0]), .Z(n122) );
  EOI U118 ( .A(dx_gpr_rd_addr1[0]), .B(n122), .Z(n99) );
  IVI U119 ( .A(m_gpr_wr_addr[4]), .Z(n124) );
  ND2I U120 ( .A(n101), .B(n104), .Z(n103) );
  IVI U121 ( .A(n103), .Z(x_fwd_alu_src1[0]) );
  ENI U122 ( .A(n123), .B(n6), .Z(n105) );
  NR2I U123 ( .A(xm_opcode[5]), .B(n105), .Z(n112) );
  ENI U124 ( .A(n13), .B(n64), .Z(n110) );
  ENI U125 ( .A(n124), .B(n2), .Z(n109) );
  ENI U126 ( .A(m_gpr_wr_addr[3]), .B(n4), .Z(n107) );
  ENI U127 ( .A(n62), .B(n60), .Z(n106) );
  ND2I U128 ( .A(n107), .B(n106), .Z(n108) );
  ND2I U129 ( .A(n112), .B(n111), .Z(n120) );
  EOI U130 ( .A(gpr_wr_addr[4]), .B(n2), .Z(n116) );
  IVI U131 ( .A(n113), .Z(n138) );
  NR2I U132 ( .A(n62), .B(n64), .Z(n114) );
  ND4 U133 ( .A(n114), .B(n5), .C(n3), .D(n1), .Z(n115) );
  ND3 U134 ( .A(fd_opcode[2]), .B(n59), .C(n115), .Z(n121) );
  ND2I U135 ( .A(n118), .B(n117), .Z(n119) );
  EOI U136 ( .A(fd_rs[2]), .B(n123), .Z(n128) );
  EOI U137 ( .A(fd_rs[3]), .B(n9), .Z(n127) );
  IVI U138 ( .A(fd_funct[3]), .Z(n130) );
  OR4 U139 ( .A(fd_funct[0]), .B(n130), .C(fd_funct[2]), .D(fd_funct[1]), .Z(
        n131) );
  NR4 U140 ( .A(n131), .B(fd_opcode[0]), .C(fd_funct[5]), .D(fd_funct[4]), .Z(
        n137) );
  NR2I U141 ( .A(fd_rs[1]), .B(fd_rs[0]), .Z(n135) );
  IVI U142 ( .A(fd_rs[2]), .Z(n134) );
  IVI U143 ( .A(fd_rs[3]), .Z(n133) );
  IVI U144 ( .A(fd_rs[4]), .Z(n132) );
  ND4 U145 ( .A(n135), .B(n134), .C(n133), .D(n132), .Z(n136) );
  AO3 U146 ( .A(fd_opcode[2]), .B(n137), .C(n59), .D(n136), .Z(n143) );
  ND2I U147 ( .A(n140), .B(n139), .Z(n141) );
  IVI U148 ( .A(n141), .Z(d_fwd_rs[0]) );
endmodule


module processor ( clock, reset, PC, Inst, MemRead, MemWrite, Addr, Din, Dout
 );
  output [31:0] PC;
  input [31:0] Inst;
  output [31:0] Addr;
  output [31:0] Din;
  input [31:0] Dout;
  input clock, reset;
  output MemRead, MemWrite;
  wire   d_PCSrc1, d_PCSrc2, d_PCSrc3, dx_Inst_5, dx_Inst_4, dx_Inst_3,
         dx_Inst_2, dx_Inst_1, dx_Inst_0, mw_Inst_5, mw_Inst_4, mw_Inst_3,
         mw_Inst_2, mw_Inst_1, mw_Inst_0, xm_Inst_5, xm_Inst_4, xm_Inst_3,
         xm_Inst_2, xm_Inst_1, xm_Inst_0, w_RegWrite, w_RegDest, w_MemtoReg,
         w_isJAL, m_isJAL, m_RegDest, x_ALUSrc, x_isSLL_SRL, d_isSLL_SRL, n4,
         n6, n30, n31, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139;
  wire   [31:0] Inst_stall_b_j;
  wire   [31:0] fd_Inst_stall;
  wire   [31:0] d_pc_plus_8;
  wire   [31:0] gpr_rd_data2;
  wire   [31:11] dx_Inst;
  wire   [31:0] dx_pc_plus_8;
  wire   [31:0] x_ALU_Result;
  wire   [31:0] dx_Inst_15_0_signext;
  wire   [31:0] dx_shamt;
  wire   [31:0] dx_gpr_rd_data1;
  wire   [4:0] dx_gpr_rd_addr1;
  wire   [31:11] mw_Inst;
  wire   [31:0] mw_pc_plus_8;
  wire   [31:0] mw_Dout;
  wire   [31:0] mw_ALU_Result;
  wire   [31:0] xm_pc_plus_8;
  wire   [31:11] xm_Inst;
  wire   [31:0] dx_gpr_rd_data2;
  wire   [31:0] d_Inst_15_0_signext;
  wire   [31:0] gpr_rd_data1;
  wire   [4:0] gpr_rd_addr1;
  wire   [31:0] d_br_signext_sl2;
  wire   [31:0] mem_alu_data_out;
  wire   [1:0] d_fwd_rs;
  wire   [31:0] fwd_data_DECODE_src1;
  wire   [31:0] fwd_gpr_rd_data1;
  wire   [1:0] d_fwd_rt;
  wire   [31:0] fwd_data_DECODE_src2;
  wire   [31:0] fwd_gpr_rd_data2;
  wire   [2:0] x_ALU_Control;
  wire   [4:0] gpr_wr_addr0;
  wire   [4:0] gpr_wr_addr;
  wire   [4:0] m_gpr_wr_addr0;
  wire   [4:0] m_gpr_wr_addr;
  wire   [31:0] gpr_wr_data;
  wire   [31:0] x_gpr_rd_data2_I;
  wire   [31:0] x_gpr_rd_data2_I_shamt;
  wire   [1:0] x_fwd_alu_src1;
  wire   [31:0] fwd_data_ALU_src1;
  wire   [1:0] x_fwd_alu_src2;
  wire   [31:0] fwd_data_ALU_src2;
  wire   [31:0] ALU_datain1;
  wire   [31:0] ALU_datain2;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  FD2 \mw_Dout_reg[31]  ( .D(Dout[31]), .CP(clock), .CD(n139), .Q(mw_Dout[31])
         );
  FD2 \mw_Dout_reg[30]  ( .D(Dout[30]), .CP(clock), .CD(n139), .Q(mw_Dout[30])
         );
  FD2 \mw_Dout_reg[29]  ( .D(Dout[29]), .CP(clock), .CD(n139), .Q(mw_Dout[29])
         );
  FD2 \mw_Dout_reg[28]  ( .D(Dout[28]), .CP(clock), .CD(n139), .Q(mw_Dout[28])
         );
  FD2 \mw_Dout_reg[27]  ( .D(Dout[27]), .CP(clock), .CD(n139), .Q(mw_Dout[27])
         );
  FD2 \mw_Dout_reg[26]  ( .D(Dout[26]), .CP(clock), .CD(n139), .Q(mw_Dout[26])
         );
  FD2 \mw_Dout_reg[25]  ( .D(Dout[25]), .CP(clock), .CD(n139), .Q(mw_Dout[25])
         );
  FD2 \mw_Dout_reg[24]  ( .D(Dout[24]), .CP(clock), .CD(n139), .Q(mw_Dout[24])
         );
  FD2 \mw_Dout_reg[23]  ( .D(Dout[23]), .CP(clock), .CD(n139), .Q(mw_Dout[23])
         );
  FD2 \mw_Dout_reg[22]  ( .D(Dout[22]), .CP(clock), .CD(n139), .Q(mw_Dout[22])
         );
  FD2 \mw_Dout_reg[21]  ( .D(Dout[21]), .CP(clock), .CD(n139), .Q(mw_Dout[21])
         );
  FD2 \mw_Dout_reg[20]  ( .D(Dout[20]), .CP(clock), .CD(n139), .Q(mw_Dout[20])
         );
  FD2 \mw_Dout_reg[19]  ( .D(Dout[19]), .CP(clock), .CD(n139), .Q(mw_Dout[19])
         );
  FD2 \mw_Dout_reg[18]  ( .D(Dout[18]), .CP(clock), .CD(n139), .Q(mw_Dout[18])
         );
  FD2 \mw_Dout_reg[17]  ( .D(Dout[17]), .CP(clock), .CD(n139), .Q(mw_Dout[17])
         );
  FD2 \mw_Dout_reg[16]  ( .D(Dout[16]), .CP(clock), .CD(n139), .Q(mw_Dout[16])
         );
  FD2 \mw_Dout_reg[15]  ( .D(Dout[15]), .CP(clock), .CD(n139), .Q(mw_Dout[15])
         );
  FD2 \mw_Dout_reg[14]  ( .D(Dout[14]), .CP(clock), .CD(n139), .Q(mw_Dout[14])
         );
  FD2 \mw_Dout_reg[13]  ( .D(Dout[13]), .CP(clock), .CD(n139), .Q(mw_Dout[13])
         );
  FD2 \mw_Dout_reg[12]  ( .D(Dout[12]), .CP(clock), .CD(n139), .Q(mw_Dout[12])
         );
  FD2 \mw_Dout_reg[11]  ( .D(Dout[11]), .CP(clock), .CD(n139), .Q(mw_Dout[11])
         );
  FD2 \mw_Dout_reg[10]  ( .D(Dout[10]), .CP(clock), .CD(n139), .Q(mw_Dout[10])
         );
  FD2 \mw_Dout_reg[9]  ( .D(Dout[9]), .CP(clock), .CD(n139), .Q(mw_Dout[9]) );
  FD2 \mw_Dout_reg[8]  ( .D(Dout[8]), .CP(clock), .CD(n139), .Q(mw_Dout[8]) );
  FD2 \mw_Dout_reg[7]  ( .D(Dout[7]), .CP(clock), .CD(n139), .Q(mw_Dout[7]) );
  FD2 \mw_Dout_reg[6]  ( .D(Dout[6]), .CP(clock), .CD(n139), .Q(mw_Dout[6]) );
  FD2 \mw_Dout_reg[5]  ( .D(Dout[5]), .CP(clock), .CD(n139), .Q(mw_Dout[5]) );
  FD2 \mw_Dout_reg[4]  ( .D(Dout[4]), .CP(clock), .CD(n139), .Q(mw_Dout[4]) );
  FD2 \mw_Dout_reg[3]  ( .D(Dout[3]), .CP(clock), .CD(n139), .Q(mw_Dout[3]) );
  FD2 \mw_Dout_reg[2]  ( .D(Dout[2]), .CP(clock), .CD(n139), .Q(mw_Dout[2]) );
  FD2 \mw_Dout_reg[1]  ( .D(Dout[1]), .CP(clock), .CD(n139), .Q(mw_Dout[1]) );
  FD2 \mw_Dout_reg[0]  ( .D(Dout[0]), .CP(clock), .CD(n139), .Q(mw_Dout[0]) );
  FD2 \mw_pc_plus_8_reg[0]  ( .D(xm_pc_plus_8[0]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[0]) );
  FD2 \xm_gpr_rd_data2_reg[0]  ( .D(dx_gpr_rd_data2[0]), .CP(clock), .CD(n139), 
        .Q(Din[0]) );
  FD2 \dx_gpr_rd_data2_reg[1]  ( .D(gpr_rd_data2[1]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[1]) );
  FD2 \xm_gpr_rd_data2_reg[1]  ( .D(dx_gpr_rd_data2[1]), .CP(clock), .CD(n139), 
        .Q(Din[1]) );
  FD2 \dx_gpr_rd_data2_reg[2]  ( .D(gpr_rd_data2[2]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[2]) );
  FD2 \xm_gpr_rd_data2_reg[2]  ( .D(dx_gpr_rd_data2[2]), .CP(clock), .CD(n139), 
        .Q(Din[2]) );
  FD2 \dx_gpr_rd_data2_reg[3]  ( .D(gpr_rd_data2[3]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[3]) );
  FD2 \xm_gpr_rd_data2_reg[3]  ( .D(dx_gpr_rd_data2[3]), .CP(clock), .CD(n139), 
        .Q(Din[3]) );
  FD2 \dx_gpr_rd_data2_reg[4]  ( .D(gpr_rd_data2[4]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[4]) );
  FD2 \xm_gpr_rd_data2_reg[4]  ( .D(dx_gpr_rd_data2[4]), .CP(clock), .CD(n139), 
        .Q(Din[4]) );
  FD2 \dx_gpr_rd_data2_reg[5]  ( .D(gpr_rd_data2[5]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[5]) );
  FD2 \dx_gpr_rd_data2_reg[6]  ( .D(gpr_rd_data2[6]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[6]) );
  FD2 \dx_gpr_rd_data2_reg[7]  ( .D(gpr_rd_data2[7]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[7]) );
  FD2 \dx_gpr_rd_data2_reg[8]  ( .D(gpr_rd_data2[8]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[8]) );
  FD2 \dx_gpr_rd_data2_reg[10]  ( .D(gpr_rd_data2[10]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[10]) );
  FD2 \dx_gpr_rd_data2_reg[11]  ( .D(gpr_rd_data2[11]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[11]) );
  FD2 \dx_gpr_rd_data2_reg[12]  ( .D(gpr_rd_data2[12]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[12]) );
  FD2 \dx_gpr_rd_data2_reg[13]  ( .D(gpr_rd_data2[13]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[13]) );
  FD2 \dx_gpr_rd_data2_reg[15]  ( .D(gpr_rd_data2[15]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[15]) );
  FD2 \dx_gpr_rd_data2_reg[16]  ( .D(gpr_rd_data2[16]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[16]) );
  FD2 \dx_gpr_rd_data2_reg[17]  ( .D(gpr_rd_data2[17]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[17]) );
  FD2 \dx_gpr_rd_data2_reg[18]  ( .D(gpr_rd_data2[18]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[18]) );
  FD2 \dx_gpr_rd_data2_reg[19]  ( .D(gpr_rd_data2[19]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[19]) );
  FD2 \dx_gpr_rd_data2_reg[20]  ( .D(gpr_rd_data2[20]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[20]) );
  FD2 \dx_gpr_rd_data2_reg[21]  ( .D(gpr_rd_data2[21]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[21]) );
  FD2 \dx_gpr_rd_data2_reg[22]  ( .D(gpr_rd_data2[22]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[22]) );
  FD2 \dx_gpr_rd_data2_reg[24]  ( .D(gpr_rd_data2[24]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[24]) );
  FD2 \dx_gpr_rd_data2_reg[25]  ( .D(gpr_rd_data2[25]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[25]) );
  FD2 \dx_gpr_rd_data2_reg[26]  ( .D(gpr_rd_data2[26]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[26]) );
  FD2 \dx_gpr_rd_data2_reg[27]  ( .D(gpr_rd_data2[27]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[27]) );
  FD2 \dx_gpr_rd_data2_reg[28]  ( .D(gpr_rd_data2[28]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[28]) );
  FD2 \dx_gpr_rd_data2_reg[30]  ( .D(gpr_rd_data2[30]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[30]) );
  FD2 \dx_gpr_rd_data2_reg[31]  ( .D(gpr_rd_data2[31]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[31]) );
  FD2 \dx_gpr_rd_data1_reg[4]  ( .D(gpr_rd_data1[4]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[4]) );
  FD2 \fd_Inst_reg[9]  ( .D(Inst_stall_b_j[9]), .CP(clock), .CD(n139), .Q(n125) );
  FD2 \dx_shamt_reg[3]  ( .D(n125), .CP(clock), .CD(n139), .Q(dx_shamt[3]) );
  FD2 \fd_Inst_reg[8]  ( .D(Inst_stall_b_j[8]), .CP(clock), .CD(n139), .Q(n126) );
  FD2 \dx_shamt_reg[2]  ( .D(n126), .CP(clock), .CD(n139), .Q(dx_shamt[2]) );
  FD2 \fd_Inst_reg[7]  ( .D(Inst_stall_b_j[7]), .CP(clock), .CD(n139), .Q(n127) );
  FD2 \dx_shamt_reg[1]  ( .D(n127), .CP(clock), .CD(n139), .Q(dx_shamt[1]) );
  FD2 \fd_Inst_reg[6]  ( .D(Inst_stall_b_j[6]), .CP(clock), .CD(n139), .Q(n128) );
  FD2 \dx_shamt_reg[0]  ( .D(n128), .CP(clock), .CD(n139), .Q(dx_shamt[0]) );
  FD2 \fd_Inst_reg[5]  ( .D(Inst_stall_b_j[5]), .CP(clock), .CD(n139), .Q(n112), .QN(n96) );
  FD2 \dx_Inst_reg[5]  ( .D(n97), .CP(clock), .CD(n139), .Q(dx_Inst_5) );
  FD2 \xm_Inst_reg[5]  ( .D(dx_Inst_5), .CP(clock), .CD(n139), .Q(xm_Inst_5)
         );
  FD2 \mw_Inst_reg[5]  ( .D(xm_Inst_5), .CP(clock), .CD(n139), .Q(mw_Inst_5)
         );
  FD2 \fd_Inst_reg[4]  ( .D(Inst_stall_b_j[4]), .CP(clock), .CD(n139), .Q(n93)
         );
  FD2 \xm_Inst_reg[4]  ( .D(dx_Inst_4), .CP(clock), .CD(n139), .Q(xm_Inst_4)
         );
  FD2 \mw_Inst_reg[4]  ( .D(xm_Inst_4), .CP(clock), .CD(n139), .Q(mw_Inst_4)
         );
  FD2 \fd_Inst_reg[3]  ( .D(Inst_stall_b_j[3]), .CP(clock), .CD(n139), .Q(n91), 
        .QN(n30) );
  FD2 \dx_Inst_reg[3]  ( .D(fd_Inst_stall[3]), .CP(clock), .CD(n139), .Q(
        dx_Inst_3) );
  FD2 \xm_Inst_reg[3]  ( .D(dx_Inst_3), .CP(clock), .CD(n139), .Q(xm_Inst_3)
         );
  FD2 \mw_Inst_reg[3]  ( .D(xm_Inst_3), .CP(clock), .CD(n139), .Q(mw_Inst_3)
         );
  FD2 \dx_Inst_reg[31]  ( .D(n74), .CP(clock), .CD(n139), .Q(dx_Inst[31]) );
  FD2 \xm_Inst_reg[31]  ( .D(dx_Inst[31]), .CP(clock), .CD(n139), .Q(
        xm_Inst[31]), .QN(n104) );
  FD2 \mw_Inst_reg[31]  ( .D(n105), .CP(clock), .CD(n139), .Q(mw_Inst[31]), 
        .QN(n76) );
  FD2 \fd_Inst_reg[30]  ( .D(Inst_stall_b_j[30]), .CP(clock), .CD(n139), .Q(
        fd_Inst_stall[30]) );
  FD2 \dx_Inst_reg[30]  ( .D(fd_Inst_stall[30]), .CP(clock), .CD(n139), .Q(
        dx_Inst[30]) );
  FD2 \xm_Inst_reg[30]  ( .D(dx_Inst[30]), .CP(clock), .CD(n139), .Q(
        xm_Inst[30]), .QN(n98) );
  FD2 \mw_Inst_reg[30]  ( .D(n99), .CP(clock), .CD(n139), .Q(mw_Inst[30]) );
  FD2 \fd_Inst_reg[2]  ( .D(Inst_stall_b_j[2]), .CP(clock), .CD(n139), .Q(n88), 
        .QN(n31) );
  FD2 \xm_Inst_reg[2]  ( .D(dx_Inst_2), .CP(clock), .CD(n139), .Q(xm_Inst_2)
         );
  FD2 \mw_Inst_reg[2]  ( .D(xm_Inst_2), .CP(clock), .CD(n139), .Q(mw_Inst_2)
         );
  FD2 \fd_Inst_reg[29]  ( .D(Inst_stall_b_j[29]), .CP(clock), .CD(n139), .Q(
        n83), .QN(n4) );
  FD2 \dx_Inst_reg[29]  ( .D(fd_Inst_stall[29]), .CP(clock), .CD(n139), .Q(
        dx_Inst[29]) );
  FD2 \xm_Inst_reg[29]  ( .D(dx_Inst[29]), .CP(clock), .CD(n139), .Q(
        xm_Inst[29]), .QN(n100) );
  FD2 \mw_Inst_reg[29]  ( .D(n101), .CP(clock), .CD(n139), .Q(mw_Inst[29]), 
        .QN(n106) );
  FD2 \fd_Inst_reg[28]  ( .D(Inst_stall_b_j[28]), .CP(clock), .CD(n139), .Q(
        fd_Inst_stall[28]) );
  FD2 \dx_Inst_reg[28]  ( .D(fd_Inst_stall[28]), .CP(clock), .CD(n139), .Q(
        dx_Inst[28]) );
  FD2 \xm_Inst_reg[28]  ( .D(dx_Inst[28]), .CP(clock), .CD(n139), .Q(
        xm_Inst[28]), .QN(n102) );
  FD2 \mw_Inst_reg[28]  ( .D(n103), .CP(clock), .CD(n139), .Q(mw_Inst[28]) );
  FD2 \fd_Inst_reg[27]  ( .D(Inst_stall_b_j[27]), .CP(clock), .CD(n139), .Q(
        n75), .QN(n6) );
  FD2 \dx_Inst_reg[27]  ( .D(fd_Inst_stall[27]), .CP(clock), .CD(n139), .Q(
        dx_Inst[27]) );
  FD2 \xm_Inst_reg[27]  ( .D(dx_Inst[27]), .CP(clock), .CD(n139), .Q(
        xm_Inst[27]), .QN(n86) );
  FD2 \mw_Inst_reg[27]  ( .D(n87), .CP(clock), .CD(n139), .Q(mw_Inst[27]) );
  FD2 \fd_Inst_reg[26]  ( .D(Inst_stall_b_j[26]), .CP(clock), .CD(n139), .Q(
        n80), .QN(n71) );
  FD2 \dx_Inst_reg[26]  ( .D(n72), .CP(clock), .CD(n139), .Q(dx_Inst[26]) );
  FD2 \xm_Inst_reg[26]  ( .D(dx_Inst[26]), .CP(clock), .CD(n139), .Q(
        xm_Inst[26]), .QN(n84) );
  FD2 \mw_Inst_reg[26]  ( .D(n85), .CP(clock), .CD(n139), .Q(mw_Inst[26]) );
  FD2 \fd_Inst_reg[25]  ( .D(Inst_stall_b_j[25]), .CP(clock), .CD(n139), .Q(
        n129) );
  FD2 \dx_Inst_reg[25]  ( .D(n129), .CP(clock), .CD(n139), .Q(dx_Inst[25]) );
  FD2 \mw_Inst_reg[25]  ( .D(xm_Inst[25]), .CP(clock), .CD(n139), .Q(
        mw_Inst[25]) );
  FD2 \fd_Inst_reg[24]  ( .D(Inst_stall_b_j[24]), .CP(clock), .CD(n139), .Q(
        n130) );
  FD2 \dx_Inst_reg[24]  ( .D(n130), .CP(clock), .CD(n139), .Q(dx_Inst[24]) );
  FD2 \mw_Inst_reg[24]  ( .D(xm_Inst[24]), .CP(clock), .CD(n139), .Q(
        mw_Inst[24]) );
  FD2 \fd_Inst_reg[23]  ( .D(Inst_stall_b_j[23]), .CP(clock), .CD(n139), .Q(
        n131) );
  FD2 \dx_Inst_reg[23]  ( .D(n131), .CP(clock), .CD(n139), .Q(dx_Inst[23]) );
  FD2 \mw_Inst_reg[23]  ( .D(xm_Inst[23]), .CP(clock), .CD(n139), .Q(
        mw_Inst[23]) );
  FD2 \fd_Inst_reg[22]  ( .D(Inst_stall_b_j[22]), .CP(clock), .CD(n139), .Q(
        n132) );
  FD2 \dx_Inst_reg[22]  ( .D(n132), .CP(clock), .CD(n139), .Q(dx_Inst[22]) );
  FD2 \mw_Inst_reg[22]  ( .D(xm_Inst[22]), .CP(clock), .CD(n139), .Q(
        mw_Inst[22]) );
  FD2 \fd_Inst_reg[21]  ( .D(Inst_stall_b_j[21]), .CP(clock), .CD(n139), .Q(
        n133) );
  FD2 \dx_Inst_reg[21]  ( .D(n133), .CP(clock), .CD(n139), .Q(dx_Inst[21]) );
  FD2 \mw_Inst_reg[21]  ( .D(xm_Inst[21]), .CP(clock), .CD(n139), .Q(
        mw_Inst[21]) );
  FD2 \fd_Inst_reg[20]  ( .D(Inst_stall_b_j[20]), .CP(clock), .CD(n139), .Q(
        n134) );
  FD2 \dx_Inst_reg[20]  ( .D(n134), .CP(clock), .CD(n139), .Q(dx_Inst[20]) );
  FD2 \xm_Inst_reg[20]  ( .D(dx_Inst[20]), .CP(clock), .CD(n139), .Q(
        xm_Inst[20]) );
  FD2 \mw_Inst_reg[20]  ( .D(xm_Inst[20]), .CP(clock), .CD(n139), .Q(
        mw_Inst[20]) );
  FD2 \fd_Inst_reg[1]  ( .D(Inst_stall_b_j[1]), .CP(clock), .CD(n139), .Q(
        fd_Inst_stall[1]) );
  FD2 \dx_Inst_reg[1]  ( .D(fd_Inst_stall[1]), .CP(clock), .CD(n139), .Q(
        dx_Inst_1) );
  FD2 \xm_Inst_reg[1]  ( .D(dx_Inst_1), .CP(clock), .CD(n139), .Q(xm_Inst_1)
         );
  FD2 \mw_Inst_reg[1]  ( .D(xm_Inst_1), .CP(clock), .CD(n139), .Q(mw_Inst_1)
         );
  FD2 \fd_Inst_reg[19]  ( .D(Inst_stall_b_j[19]), .CP(clock), .CD(n139), .Q(
        n135) );
  FD2 \dx_Inst_reg[19]  ( .D(n135), .CP(clock), .CD(n139), .Q(dx_Inst[19]) );
  FD2 \xm_Inst_reg[19]  ( .D(dx_Inst[19]), .CP(clock), .CD(n139), .Q(
        xm_Inst[19]) );
  FD2 \mw_Inst_reg[19]  ( .D(xm_Inst[19]), .CP(clock), .CD(n139), .Q(
        mw_Inst[19]) );
  FD2 \fd_Inst_reg[18]  ( .D(Inst_stall_b_j[18]), .CP(clock), .CD(n139), .Q(
        n136) );
  FD2 \dx_Inst_reg[18]  ( .D(n136), .CP(clock), .CD(n139), .Q(dx_Inst[18]) );
  FD2 \xm_Inst_reg[18]  ( .D(dx_Inst[18]), .CP(clock), .CD(n139), .Q(
        xm_Inst[18]) );
  FD2 \mw_Inst_reg[18]  ( .D(xm_Inst[18]), .CP(clock), .CD(n139), .Q(
        mw_Inst[18]) );
  FD2 \fd_Inst_reg[17]  ( .D(Inst_stall_b_j[17]), .CP(clock), .CD(n139), .Q(
        n137) );
  FD2 \dx_Inst_reg[17]  ( .D(n137), .CP(clock), .CD(n139), .Q(dx_Inst[17]) );
  FD2 \xm_Inst_reg[17]  ( .D(dx_Inst[17]), .CP(clock), .CD(n139), .Q(
        xm_Inst[17]) );
  FD2 \mw_Inst_reg[17]  ( .D(xm_Inst[17]), .CP(clock), .CD(n139), .Q(
        mw_Inst[17]) );
  FD2 \fd_Inst_reg[16]  ( .D(Inst_stall_b_j[16]), .CP(clock), .CD(n139), .Q(
        n138) );
  FD2 \dx_Inst_reg[16]  ( .D(n138), .CP(clock), .CD(n139), .Q(dx_Inst[16]) );
  FD2 \xm_Inst_reg[16]  ( .D(dx_Inst[16]), .CP(clock), .CD(n139), .Q(
        xm_Inst[16]) );
  FD2 \mw_Inst_reg[16]  ( .D(xm_Inst[16]), .CP(clock), .CD(n139), .Q(
        mw_Inst[16]) );
  FD2 \dx_gpr_rd_addr1_reg[0]  ( .D(gpr_rd_addr1[0]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_addr1[0]) );
  FD2 \dx_gpr_rd_addr1_reg[1]  ( .D(gpr_rd_addr1[1]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_addr1[1]) );
  FD2 \fd_Inst_reg[15]  ( .D(Inst_stall_b_j[15]), .CP(clock), .CD(n139), .Q(
        n119) );
  FD2 \dx_Inst_reg[15]  ( .D(n119), .CP(clock), .CD(n139), .Q(dx_Inst[15]) );
  FD2 \xm_Inst_reg[15]  ( .D(dx_Inst[15]), .CP(clock), .CD(n139), .Q(
        xm_Inst[15]) );
  FD2 \mw_Inst_reg[15]  ( .D(xm_Inst[15]), .CP(clock), .CD(n139), .Q(
        mw_Inst[15]) );
  FD2 \fd_Inst_reg[14]  ( .D(Inst_stall_b_j[14]), .CP(clock), .CD(n139), .Q(
        n120) );
  FD2 \dx_Inst_reg[14]  ( .D(n120), .CP(clock), .CD(n139), .Q(dx_Inst[14]) );
  FD2 \xm_Inst_reg[14]  ( .D(dx_Inst[14]), .CP(clock), .CD(n139), .Q(
        xm_Inst[14]) );
  FD2 \mw_Inst_reg[14]  ( .D(xm_Inst[14]), .CP(clock), .CD(n139), .Q(
        mw_Inst[14]) );
  FD2 \fd_Inst_reg[13]  ( .D(Inst_stall_b_j[13]), .CP(clock), .CD(n139), .Q(
        n121) );
  FD2 \dx_Inst_reg[13]  ( .D(n121), .CP(clock), .CD(n139), .Q(dx_Inst[13]) );
  FD2 \xm_Inst_reg[13]  ( .D(dx_Inst[13]), .CP(clock), .CD(n139), .Q(
        xm_Inst[13]) );
  FD2 \mw_Inst_reg[13]  ( .D(xm_Inst[13]), .CP(clock), .CD(n139), .Q(
        mw_Inst[13]) );
  FD2 \fd_Inst_reg[12]  ( .D(Inst_stall_b_j[12]), .CP(clock), .CD(n139), .Q(
        n122) );
  FD2 \dx_Inst_reg[12]  ( .D(n122), .CP(clock), .CD(n139), .Q(dx_Inst[12]) );
  FD2 \xm_Inst_reg[12]  ( .D(dx_Inst[12]), .CP(clock), .CD(n139), .Q(
        xm_Inst[12]) );
  FD2 \mw_Inst_reg[12]  ( .D(xm_Inst[12]), .CP(clock), .CD(n139), .Q(
        mw_Inst[12]) );
  FD2 \fd_Inst_reg[11]  ( .D(Inst_stall_b_j[11]), .CP(clock), .CD(n139), .Q(
        n123) );
  FD2 \dx_Inst_reg[11]  ( .D(n123), .CP(clock), .CD(n139), .Q(dx_Inst[11]) );
  FD2 \xm_Inst_reg[11]  ( .D(dx_Inst[11]), .CP(clock), .CD(n139), .Q(
        xm_Inst[11]) );
  FD2 \mw_Inst_reg[11]  ( .D(xm_Inst[11]), .CP(clock), .CD(n139), .Q(
        mw_Inst[11]) );
  FD2 \fd_Inst_reg[10]  ( .D(Inst_stall_b_j[10]), .CP(clock), .CD(n139), .Q(
        n124) );
  FD2 \dx_shamt_reg[4]  ( .D(n124), .CP(clock), .CD(n139), .Q(dx_shamt[4]) );
  FD2 \fd_Inst_reg[0]  ( .D(Inst_stall_b_j[0]), .CP(clock), .CD(n139), .Q(n92), 
        .QN(n60) );
  FD2 \dx_Inst_reg[0]  ( .D(fd_Inst_stall[0]), .CP(clock), .CD(n139), .Q(
        dx_Inst_0) );
  FD2 \xm_Inst_reg[0]  ( .D(dx_Inst_0), .CP(clock), .CD(n139), .Q(xm_Inst_0)
         );
  FD2 \mw_Inst_reg[0]  ( .D(xm_Inst_0), .CP(clock), .CD(n139), .Q(mw_Inst_0)
         );
  FD2 \dx_Inst_15_0_signext_reg[0]  ( .D(d_Inst_15_0_signext[0]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[0]) );
  FD2 \dx_Inst_15_0_signext_reg[1]  ( .D(d_Inst_15_0_signext[1]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[1]) );
  FD2 \dx_Inst_15_0_signext_reg[2]  ( .D(d_Inst_15_0_signext[2]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[2]) );
  FD2 \dx_Inst_15_0_signext_reg[3]  ( .D(d_Inst_15_0_signext[3]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[3]) );
  FD2 \dx_Inst_15_0_signext_reg[4]  ( .D(d_Inst_15_0_signext[4]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[4]) );
  FD2 \dx_Inst_15_0_signext_reg[5]  ( .D(d_Inst_15_0_signext[5]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[5]) );
  FD2 \dx_Inst_15_0_signext_reg[6]  ( .D(d_Inst_15_0_signext[6]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[6]) );
  FD2 \dx_Inst_15_0_signext_reg[7]  ( .D(d_Inst_15_0_signext[7]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[7]) );
  FD2 \dx_Inst_15_0_signext_reg[8]  ( .D(d_Inst_15_0_signext[8]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[8]) );
  FD2 \dx_Inst_15_0_signext_reg[9]  ( .D(d_Inst_15_0_signext[9]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[9]) );
  FD2 \dx_Inst_15_0_signext_reg[10]  ( .D(d_Inst_15_0_signext[10]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[10]) );
  FD2 \dx_Inst_15_0_signext_reg[11]  ( .D(d_Inst_15_0_signext[11]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[11]) );
  FD2 \dx_Inst_15_0_signext_reg[12]  ( .D(d_Inst_15_0_signext[12]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[12]) );
  FD2 \dx_Inst_15_0_signext_reg[13]  ( .D(d_Inst_15_0_signext[13]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[13]) );
  FD2 \dx_Inst_15_0_signext_reg[14]  ( .D(d_Inst_15_0_signext[14]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[14]) );
  FD2 \dx_Inst_15_0_signext_reg[15]  ( .D(d_Inst_15_0_signext[15]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[15]) );
  FD2 \dx_Inst_15_0_signext_reg[16]  ( .D(d_Inst_15_0_signext[16]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[16]) );
  FD2 \dx_Inst_15_0_signext_reg[17]  ( .D(d_Inst_15_0_signext[17]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[17]) );
  FD2 \dx_Inst_15_0_signext_reg[18]  ( .D(d_Inst_15_0_signext[18]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[18]) );
  FD2 \dx_Inst_15_0_signext_reg[19]  ( .D(d_Inst_15_0_signext[19]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[19]) );
  FD2 \dx_Inst_15_0_signext_reg[20]  ( .D(d_Inst_15_0_signext[20]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[20]) );
  FD2 \dx_Inst_15_0_signext_reg[21]  ( .D(d_Inst_15_0_signext[21]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[21]) );
  FD2 \dx_Inst_15_0_signext_reg[22]  ( .D(d_Inst_15_0_signext[22]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[22]) );
  FD2 \dx_Inst_15_0_signext_reg[23]  ( .D(d_Inst_15_0_signext[23]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[23]) );
  FD2 \dx_Inst_15_0_signext_reg[24]  ( .D(d_Inst_15_0_signext[24]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[24]) );
  FD2 \dx_Inst_15_0_signext_reg[25]  ( .D(d_Inst_15_0_signext[25]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[25]) );
  FD2 \dx_Inst_15_0_signext_reg[26]  ( .D(d_Inst_15_0_signext[26]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[26]) );
  FD2 \dx_Inst_15_0_signext_reg[27]  ( .D(d_Inst_15_0_signext[27]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[27]) );
  FD2 \dx_Inst_15_0_signext_reg[28]  ( .D(d_Inst_15_0_signext[28]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[28]) );
  FD2 \dx_Inst_15_0_signext_reg[29]  ( .D(d_Inst_15_0_signext[29]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[29]) );
  FD2 \dx_Inst_15_0_signext_reg[30]  ( .D(d_Inst_15_0_signext[30]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[30]) );
  FD2 \dx_Inst_15_0_signext_reg[31]  ( .D(d_Inst_15_0_signext[31]), .CP(clock), 
        .CD(n139), .Q(dx_Inst_15_0_signext[31]) );
  FD2 \xm_ALU_Result_reg[0]  ( .D(x_ALU_Result[0]), .CP(clock), .CD(n139), .Q(
        Addr[0]) );
  FD2 \mw_ALU_Result_reg[0]  ( .D(Addr[0]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[0]) );
  FD2 \xm_ALU_Result_reg[1]  ( .D(x_ALU_Result[1]), .CP(clock), .CD(n139), .Q(
        Addr[1]) );
  FD2 \mw_ALU_Result_reg[1]  ( .D(Addr[1]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[1]) );
  FD2 \xm_ALU_Result_reg[2]  ( .D(x_ALU_Result[2]), .CP(clock), .CD(n139), .Q(
        Addr[2]) );
  FD2 \mw_ALU_Result_reg[2]  ( .D(Addr[2]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[2]) );
  FD2 \xm_ALU_Result_reg[3]  ( .D(x_ALU_Result[3]), .CP(clock), .CD(n139), .Q(
        Addr[3]) );
  FD2 \mw_ALU_Result_reg[3]  ( .D(Addr[3]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[3]) );
  FD2 \xm_ALU_Result_reg[4]  ( .D(x_ALU_Result[4]), .CP(clock), .CD(n139), .Q(
        Addr[4]) );
  FD2 \mw_ALU_Result_reg[4]  ( .D(Addr[4]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[4]) );
  FD2 \xm_ALU_Result_reg[5]  ( .D(x_ALU_Result[5]), .CP(clock), .CD(n139), .Q(
        Addr[5]) );
  FD2 \mw_ALU_Result_reg[5]  ( .D(Addr[5]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[5]) );
  FD2 \xm_ALU_Result_reg[6]  ( .D(x_ALU_Result[6]), .CP(clock), .CD(n139), .Q(
        Addr[6]) );
  FD2 \mw_ALU_Result_reg[6]  ( .D(Addr[6]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[6]) );
  FD2 \xm_ALU_Result_reg[7]  ( .D(x_ALU_Result[7]), .CP(clock), .CD(n139), .Q(
        Addr[7]) );
  FD2 \mw_ALU_Result_reg[7]  ( .D(Addr[7]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[7]) );
  FD2 \xm_ALU_Result_reg[8]  ( .D(x_ALU_Result[8]), .CP(clock), .CD(n139), .Q(
        Addr[8]) );
  FD2 \mw_ALU_Result_reg[8]  ( .D(Addr[8]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[8]) );
  FD2 \xm_ALU_Result_reg[9]  ( .D(x_ALU_Result[9]), .CP(clock), .CD(n139), .Q(
        Addr[9]) );
  FD2 \mw_ALU_Result_reg[9]  ( .D(Addr[9]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[9]) );
  FD2 \xm_ALU_Result_reg[10]  ( .D(x_ALU_Result[10]), .CP(clock), .CD(n139), 
        .Q(Addr[10]) );
  FD2 \mw_ALU_Result_reg[10]  ( .D(Addr[10]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[10]) );
  FD2 \xm_ALU_Result_reg[11]  ( .D(x_ALU_Result[11]), .CP(clock), .CD(n139), 
        .Q(Addr[11]) );
  FD2 \mw_ALU_Result_reg[11]  ( .D(Addr[11]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[11]) );
  FD2 \xm_ALU_Result_reg[12]  ( .D(x_ALU_Result[12]), .CP(clock), .CD(n139), 
        .Q(Addr[12]) );
  FD2 \mw_ALU_Result_reg[12]  ( .D(Addr[12]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[12]) );
  FD2 \xm_ALU_Result_reg[13]  ( .D(x_ALU_Result[13]), .CP(clock), .CD(n139), 
        .Q(Addr[13]) );
  FD2 \mw_ALU_Result_reg[13]  ( .D(Addr[13]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[13]) );
  FD2 \xm_ALU_Result_reg[14]  ( .D(x_ALU_Result[14]), .CP(clock), .CD(n139), 
        .Q(Addr[14]) );
  FD2 \mw_ALU_Result_reg[14]  ( .D(Addr[14]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[14]) );
  FD2 \xm_ALU_Result_reg[15]  ( .D(x_ALU_Result[15]), .CP(clock), .CD(n139), 
        .Q(Addr[15]) );
  FD2 \mw_ALU_Result_reg[15]  ( .D(Addr[15]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[15]) );
  FD2 \xm_ALU_Result_reg[16]  ( .D(x_ALU_Result[16]), .CP(clock), .CD(n139), 
        .Q(Addr[16]) );
  FD2 \mw_ALU_Result_reg[16]  ( .D(Addr[16]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[16]) );
  FD2 \xm_ALU_Result_reg[17]  ( .D(x_ALU_Result[17]), .CP(clock), .CD(n139), 
        .Q(Addr[17]) );
  FD2 \mw_ALU_Result_reg[17]  ( .D(Addr[17]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[17]) );
  FD2 \xm_ALU_Result_reg[18]  ( .D(x_ALU_Result[18]), .CP(clock), .CD(n139), 
        .Q(Addr[18]) );
  FD2 \mw_ALU_Result_reg[18]  ( .D(Addr[18]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[18]) );
  FD2 \xm_ALU_Result_reg[19]  ( .D(x_ALU_Result[19]), .CP(clock), .CD(n139), 
        .Q(Addr[19]) );
  FD2 \mw_ALU_Result_reg[19]  ( .D(Addr[19]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[19]) );
  FD2 \xm_ALU_Result_reg[20]  ( .D(x_ALU_Result[20]), .CP(clock), .CD(n139), 
        .Q(Addr[20]) );
  FD2 \mw_ALU_Result_reg[20]  ( .D(Addr[20]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[20]) );
  FD2 \xm_ALU_Result_reg[21]  ( .D(x_ALU_Result[21]), .CP(clock), .CD(n139), 
        .Q(Addr[21]) );
  FD2 \mw_ALU_Result_reg[21]  ( .D(Addr[21]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[21]) );
  FD2 \xm_ALU_Result_reg[22]  ( .D(x_ALU_Result[22]), .CP(clock), .CD(n139), 
        .Q(Addr[22]) );
  FD2 \mw_ALU_Result_reg[22]  ( .D(Addr[22]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[22]) );
  FD2 \xm_ALU_Result_reg[23]  ( .D(x_ALU_Result[23]), .CP(clock), .CD(n139), 
        .Q(Addr[23]) );
  FD2 \mw_ALU_Result_reg[23]  ( .D(Addr[23]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[23]) );
  FD2 \xm_ALU_Result_reg[24]  ( .D(x_ALU_Result[24]), .CP(clock), .CD(n139), 
        .Q(Addr[24]) );
  FD2 \mw_ALU_Result_reg[24]  ( .D(Addr[24]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[24]) );
  FD2 \xm_ALU_Result_reg[25]  ( .D(x_ALU_Result[25]), .CP(clock), .CD(n139), 
        .Q(Addr[25]) );
  FD2 \mw_ALU_Result_reg[25]  ( .D(Addr[25]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[25]) );
  FD2 \xm_ALU_Result_reg[26]  ( .D(x_ALU_Result[26]), .CP(clock), .CD(n139), 
        .Q(Addr[26]) );
  FD2 \mw_ALU_Result_reg[26]  ( .D(Addr[26]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[26]) );
  FD2 \xm_ALU_Result_reg[27]  ( .D(x_ALU_Result[27]), .CP(clock), .CD(n139), 
        .Q(Addr[27]) );
  FD2 \mw_ALU_Result_reg[27]  ( .D(Addr[27]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[27]) );
  FD2 \xm_ALU_Result_reg[28]  ( .D(x_ALU_Result[28]), .CP(clock), .CD(n139), 
        .Q(Addr[28]) );
  FD2 \mw_ALU_Result_reg[28]  ( .D(Addr[28]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[28]) );
  FD2 \xm_ALU_Result_reg[29]  ( .D(x_ALU_Result[29]), .CP(clock), .CD(n139), 
        .Q(Addr[29]) );
  FD2 \mw_ALU_Result_reg[29]  ( .D(Addr[29]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[29]) );
  FD2 \xm_ALU_Result_reg[30]  ( .D(x_ALU_Result[30]), .CP(clock), .CD(n139), 
        .Q(Addr[30]) );
  FD2 \mw_ALU_Result_reg[30]  ( .D(Addr[30]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[30]) );
  FD2 \xm_ALU_Result_reg[31]  ( .D(x_ALU_Result[31]), .CP(clock), .CD(n139), 
        .Q(Addr[31]) );
  FD2 \mw_ALU_Result_reg[31]  ( .D(Addr[31]), .CP(clock), .CD(n139), .Q(
        mw_ALU_Result[31]) );
  FD2 \dx_pc_plus_8_reg[0]  ( .D(d_pc_plus_8[0]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[0]) );
  FD2 \dx_pc_plus_8_reg[1]  ( .D(d_pc_plus_8[1]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[1]) );
  FD2 \mw_pc_plus_8_reg[1]  ( .D(xm_pc_plus_8[1]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[1]) );
  FD2 \dx_pc_plus_8_reg[2]  ( .D(d_pc_plus_8[2]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[2]) );
  FD2 \mw_pc_plus_8_reg[2]  ( .D(xm_pc_plus_8[2]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[2]) );
  FD2 \dx_pc_plus_8_reg[3]  ( .D(d_pc_plus_8[3]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[3]) );
  FD2 \mw_pc_plus_8_reg[3]  ( .D(xm_pc_plus_8[3]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[3]) );
  FD2 \dx_pc_plus_8_reg[4]  ( .D(d_pc_plus_8[4]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[4]) );
  FD2 \mw_pc_plus_8_reg[4]  ( .D(xm_pc_plus_8[4]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[4]) );
  FD2 \dx_pc_plus_8_reg[5]  ( .D(d_pc_plus_8[5]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[5]) );
  FD2 \mw_pc_plus_8_reg[5]  ( .D(xm_pc_plus_8[5]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[5]) );
  FD2 \dx_pc_plus_8_reg[6]  ( .D(d_pc_plus_8[6]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[6]) );
  FD2 \mw_pc_plus_8_reg[6]  ( .D(xm_pc_plus_8[6]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[6]) );
  FD2 \dx_pc_plus_8_reg[7]  ( .D(d_pc_plus_8[7]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[7]) );
  FD2 \mw_pc_plus_8_reg[7]  ( .D(xm_pc_plus_8[7]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[7]) );
  FD2 \dx_pc_plus_8_reg[8]  ( .D(d_pc_plus_8[8]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[8]) );
  FD2 \mw_pc_plus_8_reg[8]  ( .D(xm_pc_plus_8[8]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[8]) );
  FD2 \dx_pc_plus_8_reg[9]  ( .D(d_pc_plus_8[9]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[9]) );
  FD2 \mw_pc_plus_8_reg[9]  ( .D(xm_pc_plus_8[9]), .CP(clock), .CD(n139), .Q(
        mw_pc_plus_8[9]) );
  FD2 \dx_pc_plus_8_reg[10]  ( .D(d_pc_plus_8[10]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[10]) );
  FD2 \mw_pc_plus_8_reg[10]  ( .D(xm_pc_plus_8[10]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[10]) );
  FD2 \dx_pc_plus_8_reg[11]  ( .D(d_pc_plus_8[11]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[11]) );
  FD2 \mw_pc_plus_8_reg[11]  ( .D(xm_pc_plus_8[11]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[11]) );
  FD2 \dx_pc_plus_8_reg[12]  ( .D(d_pc_plus_8[12]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[12]) );
  FD2 \mw_pc_plus_8_reg[12]  ( .D(xm_pc_plus_8[12]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[12]) );
  FD2 \dx_pc_plus_8_reg[13]  ( .D(d_pc_plus_8[13]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[13]) );
  FD2 \mw_pc_plus_8_reg[13]  ( .D(xm_pc_plus_8[13]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[13]) );
  FD2 \dx_pc_plus_8_reg[14]  ( .D(d_pc_plus_8[14]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[14]) );
  FD2 \mw_pc_plus_8_reg[14]  ( .D(xm_pc_plus_8[14]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[14]) );
  FD2 \dx_pc_plus_8_reg[15]  ( .D(d_pc_plus_8[15]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[15]) );
  FD2 \mw_pc_plus_8_reg[15]  ( .D(xm_pc_plus_8[15]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[15]) );
  FD2 \dx_pc_plus_8_reg[16]  ( .D(d_pc_plus_8[16]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[16]) );
  FD2 \mw_pc_plus_8_reg[16]  ( .D(xm_pc_plus_8[16]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[16]) );
  FD2 \dx_pc_plus_8_reg[17]  ( .D(d_pc_plus_8[17]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[17]) );
  FD2 \mw_pc_plus_8_reg[17]  ( .D(xm_pc_plus_8[17]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[17]) );
  FD2 \dx_pc_plus_8_reg[18]  ( .D(d_pc_plus_8[18]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[18]) );
  FD2 \mw_pc_plus_8_reg[18]  ( .D(xm_pc_plus_8[18]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[18]) );
  FD2 \dx_pc_plus_8_reg[19]  ( .D(d_pc_plus_8[19]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[19]) );
  FD2 \mw_pc_plus_8_reg[19]  ( .D(xm_pc_plus_8[19]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[19]) );
  FD2 \dx_pc_plus_8_reg[20]  ( .D(d_pc_plus_8[20]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[20]) );
  FD2 \mw_pc_plus_8_reg[20]  ( .D(xm_pc_plus_8[20]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[20]) );
  FD2 \dx_pc_plus_8_reg[21]  ( .D(d_pc_plus_8[21]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[21]) );
  FD2 \mw_pc_plus_8_reg[21]  ( .D(xm_pc_plus_8[21]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[21]) );
  FD2 \dx_pc_plus_8_reg[22]  ( .D(d_pc_plus_8[22]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[22]) );
  FD2 \mw_pc_plus_8_reg[22]  ( .D(xm_pc_plus_8[22]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[22]) );
  FD2 \dx_pc_plus_8_reg[23]  ( .D(d_pc_plus_8[23]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[23]) );
  FD2 \mw_pc_plus_8_reg[23]  ( .D(xm_pc_plus_8[23]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[23]) );
  FD2 \dx_pc_plus_8_reg[24]  ( .D(d_pc_plus_8[24]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[24]) );
  FD2 \mw_pc_plus_8_reg[24]  ( .D(xm_pc_plus_8[24]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[24]) );
  FD2 \dx_pc_plus_8_reg[25]  ( .D(d_pc_plus_8[25]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[25]) );
  FD2 \mw_pc_plus_8_reg[25]  ( .D(xm_pc_plus_8[25]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[25]) );
  FD2 \dx_pc_plus_8_reg[26]  ( .D(d_pc_plus_8[26]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[26]) );
  FD2 \mw_pc_plus_8_reg[26]  ( .D(xm_pc_plus_8[26]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[26]) );
  FD2 \dx_pc_plus_8_reg[27]  ( .D(d_pc_plus_8[27]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[27]) );
  FD2 \mw_pc_plus_8_reg[27]  ( .D(xm_pc_plus_8[27]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[27]) );
  FD2 \dx_pc_plus_8_reg[28]  ( .D(d_pc_plus_8[28]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[28]) );
  FD2 \mw_pc_plus_8_reg[28]  ( .D(xm_pc_plus_8[28]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[28]) );
  FD2 \dx_pc_plus_8_reg[29]  ( .D(d_pc_plus_8[29]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[29]) );
  FD2 \mw_pc_plus_8_reg[29]  ( .D(xm_pc_plus_8[29]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[29]) );
  FD2 \dx_pc_plus_8_reg[30]  ( .D(d_pc_plus_8[30]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[30]) );
  FD2 \mw_pc_plus_8_reg[30]  ( .D(xm_pc_plus_8[30]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[30]) );
  FD2 \dx_pc_plus_8_reg[31]  ( .D(d_pc_plus_8[31]), .CP(clock), .CD(n139), .Q(
        dx_pc_plus_8[31]) );
  FD2 \mw_pc_plus_8_reg[31]  ( .D(xm_pc_plus_8[31]), .CP(clock), .CD(n139), 
        .Q(mw_pc_plus_8[31]) );
  signext signext_u0 ( .ip({n119, n120, n121, n122, n123, n124, n125, n126, 
        n127, n128, n97, n57, fd_Inst_stall[3], n90, fd_Inst_stall[1:0]}), 
        .op(d_Inst_15_0_signext) );
  lshift lshift_u0 ( .ip(d_Inst_15_0_signext), .op({d_br_signext_sl2[31:2], 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  mux_2x1_DATA_WIDTH32_0 mux_2x1_FWD_D1 ( .ip1(mem_alu_data_out), .ip0(Addr), 
        .sel(d_fwd_rs[0]), .out(fwd_data_DECODE_src1) );
  mux_2x1_DATA_WIDTH32_11 mux_2x1_FWD_D2 ( .ip1(fwd_data_DECODE_src1), .ip0(
        gpr_rd_data1), .sel(d_fwd_rs[1]), .out(fwd_gpr_rd_data1) );
  mux_2x1_DATA_WIDTH32_10 mux_2x1_FWD_D3 ( .ip1(mem_alu_data_out), .ip0(Addr), 
        .sel(d_fwd_rt[0]), .out(fwd_data_DECODE_src2) );
  mux_2x1_DATA_WIDTH32_9 mux_2x1_FWD_D4 ( .ip1(fwd_data_DECODE_src2), .ip0(
        gpr_rd_data2), .sel(d_fwd_rt[1]), .out(fwd_gpr_rd_data2) );
  pc pc_u0 ( .clk(clock), .rst(reset), .fd_br_signext_sl2({
        d_br_signext_sl2[31:2], 1'b0, 1'b0}), .fd_Inst_25_0({n129, n130, n131, 
        n132, n133, n134, n135, n136, n137, n138, n119, n120, n121, n122, n123, 
        n124, n125, n126, n127, n128, n97, n57, fd_Inst_stall[3], n90, 
        fd_Inst_stall[1:0]}), .fwd_gpr_rd_data1(fwd_gpr_rd_data1), .d_stall(
        1'b0), .jump(d_PCSrc1), .branch(d_PCSrc2), .jump_reg(d_PCSrc3), .pc(PC), .d_pc_plus_8(d_pc_plus_8) );
  control_unit control_unit_u0 ( .mw_opcode(mw_Inst[31:26]), .mw_funct({
        mw_Inst_5, mw_Inst_4, mw_Inst_3, mw_Inst_2, mw_Inst_1, mw_Inst_0}), 
        .mw_rs(mw_Inst[25:21]), .mw_rt(mw_Inst[20:16]), .mw_rd(mw_Inst[15:11]), 
        .xm_opcode(xm_Inst[31:26]), .dx_opcode(dx_Inst[31:26]), .dx_funct({
        dx_Inst_5, dx_Inst_4, dx_Inst_3, dx_Inst_2, dx_Inst_1, dx_Inst_0}), 
        .fd_opcode({n111, fd_Inst_stall[30], n83, fd_Inst_stall[28], n75, n80}), .fd_funct({n112, n93, n91, n88, fd_Inst_stall[1], n92}), .fwd_gpr_rd_data1(
        fwd_gpr_rd_data1), .fwd_gpr_rd_data2(fwd_gpr_rd_data2), .w_RegWrite(
        w_RegWrite), .w_RegDest(w_RegDest), .w_MemtoReg(w_MemtoReg), .w_isJAL(
        w_isJAL), .m_MemRead(MemRead), .m_MemWrite(MemWrite), .m_isJAL(m_isJAL), .m_RegDest(m_RegDest), .x_ALUSrc(x_ALUSrc), .x_isSLL_SRL(x_isSLL_SRL), 
        .x_ALU_Control(x_ALU_Control), .d_PCSrc1(d_PCSrc1), .d_PCSrc2(d_PCSrc2), .d_PCSrc3(d_PCSrc3), .d_isSLL_SRL(d_isSLL_SRL) );
  mux_2x1_DATA_WIDTH5_0 mux_2x1_u0 ( .ip1(mw_Inst[15:11]), .ip0(mw_Inst[20:16]), .sel(w_RegDest), .out(gpr_wr_addr0) );
  mux_2x1_DATA_WIDTH5_4 mux_2x1_u1 ( .ip1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .ip0(gpr_wr_addr0), .sel(w_isJAL), .out(gpr_wr_addr) );
  mux_2x1_DATA_WIDTH5_3 mux_2x1_u2 ( .ip1(xm_Inst[15:11]), .ip0(xm_Inst[20:16]), .sel(m_RegDest), .out(m_gpr_wr_addr0) );
  mux_2x1_DATA_WIDTH5_2 mux_2x1_u3 ( .ip1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .ip0(m_gpr_wr_addr0), .sel(m_isJAL), .out(m_gpr_wr_addr) );
  mux_2x1_DATA_WIDTH32_8 mux_2x1_u4 ( .ip1(mw_Dout), .ip0(mw_ALU_Result), 
        .sel(w_MemtoReg), .out(mem_alu_data_out) );
  mux_2x1_DATA_WIDTH32_7 mux_2x1_u5 ( .ip1(mw_pc_plus_8), .ip0(
        mem_alu_data_out), .sel(w_isJAL), .out(gpr_wr_data) );
  mux_2x1_DATA_WIDTH5_1 mux_2x1_u6 ( .ip1({n134, n135, n136, n137, n138}), 
        .ip0({n129, n130, n131, n132, n133}), .sel(n110), .out(gpr_rd_addr1)
         );
  gpr gpr_u0 ( .clk(clock), .RegWrite(w_RegWrite), .rd_addr1(gpr_rd_addr1), 
        .rd_addr2({n134, n135, n136, n137, n138}), .wr_addr({n58, n59, n82, 
        n79, n95}), .wr_data(gpr_wr_data), .rd_data1(gpr_rd_data1), .rd_data2(
        gpr_rd_data2) );
  mux_2x1_DATA_WIDTH32_6 mux_2x1_u7 ( .ip1(dx_Inst_15_0_signext), .ip0(
        dx_gpr_rd_data2), .sel(x_ALUSrc), .out(x_gpr_rd_data2_I) );
  mux_2x1_DATA_WIDTH32_5 mux_2x1_u8 ( .ip1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, dx_shamt[4:0]}), 
        .ip0(x_gpr_rd_data2_I), .sel(x_isSLL_SRL), .out(x_gpr_rd_data2_I_shamt) );
  mux_2x1_DATA_WIDTH32_4 mux_2x1_u9 ( .ip1(mem_alu_data_out), .ip0(Addr), 
        .sel(x_fwd_alu_src1[0]), .out(fwd_data_ALU_src1) );
  mux_2x1_DATA_WIDTH32_3 mux_2x1_u10 ( .ip1(mem_alu_data_out), .ip0(Addr), 
        .sel(x_fwd_alu_src2[0]), .out(fwd_data_ALU_src2) );
  mux_2x1_DATA_WIDTH32_2 mux_2x1_u11 ( .ip1(fwd_data_ALU_src1), .ip0(
        dx_gpr_rd_data1), .sel(x_fwd_alu_src1[1]), .out(ALU_datain1) );
  mux_2x1_DATA_WIDTH32_1 mux_2x1_u12 ( .ip1(fwd_data_ALU_src2), .ip0(
        x_gpr_rd_data2_I_shamt), .sel(x_fwd_alu_src2[1]), .out(ALU_datain2) );
  alu alu_u0 ( .r1(ALU_datain1), .r2(ALU_datain2), .control(x_ALU_Control), 
        .result(x_ALU_Result) );
  forward_stall forward_stall_u0 ( .gpr_wr_addr(gpr_wr_addr), .m_gpr_wr_addr(
        m_gpr_wr_addr), .mw_opcode({n77, mw_Inst[30], n107, mw_Inst[28:26]}), 
        .xm_opcode({n105, n99, n101, n103, n87, n85}), .xm_rt(xm_Inst[20:16]), 
        .dx_gpr_rd_addr1(dx_gpr_rd_addr1), .dx_rt(dx_Inst[20:16]), 
        .dx_isSLL_SRL(n110), .dx_opcode(dx_Inst[31:26]), .fd_opcode({n74, 
        fd_Inst_stall[30:27], n72}), .fd_funct({n97, n57, n91, 
        fd_Inst_stall[2:1], n92}), .fd_rs({n129, n130, n131, n132, n133}), 
        .fd_rt({n134, n135, n136, n137, n138}), .gpr_rd_addr1(gpr_rd_addr1), 
        .d_fwd_rs(d_fwd_rs), .d_fwd_rt(d_fwd_rt), .x_fwd_alu_src1(
        x_fwd_alu_src1), .x_fwd_alu_src2(x_fwd_alu_src2), .Port20(1'b0) );
  FD2 \xm_pc_plus_8_reg[31]  ( .D(dx_pc_plus_8[31]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[31]) );
  FD2 \xm_pc_plus_8_reg[30]  ( .D(dx_pc_plus_8[30]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[30]) );
  FD2 \xm_pc_plus_8_reg[29]  ( .D(dx_pc_plus_8[29]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[29]) );
  FD2 \xm_pc_plus_8_reg[28]  ( .D(dx_pc_plus_8[28]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[28]) );
  FD2 \xm_pc_plus_8_reg[27]  ( .D(dx_pc_plus_8[27]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[27]) );
  FD2 \xm_pc_plus_8_reg[26]  ( .D(dx_pc_plus_8[26]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[26]) );
  FD2 \xm_pc_plus_8_reg[25]  ( .D(dx_pc_plus_8[25]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[25]) );
  FD2 \xm_pc_plus_8_reg[24]  ( .D(dx_pc_plus_8[24]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[24]) );
  FD2 \xm_pc_plus_8_reg[23]  ( .D(dx_pc_plus_8[23]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[23]) );
  FD2 \xm_pc_plus_8_reg[22]  ( .D(dx_pc_plus_8[22]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[22]) );
  FD2 \xm_pc_plus_8_reg[21]  ( .D(dx_pc_plus_8[21]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[21]) );
  FD2 \xm_pc_plus_8_reg[20]  ( .D(dx_pc_plus_8[20]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[20]) );
  FD2 \xm_pc_plus_8_reg[19]  ( .D(dx_pc_plus_8[19]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[19]) );
  FD2 \xm_pc_plus_8_reg[18]  ( .D(dx_pc_plus_8[18]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[18]) );
  FD2 \xm_pc_plus_8_reg[17]  ( .D(dx_pc_plus_8[17]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[17]) );
  FD2 \xm_pc_plus_8_reg[16]  ( .D(dx_pc_plus_8[16]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[16]) );
  FD2 \xm_pc_plus_8_reg[15]  ( .D(dx_pc_plus_8[15]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[15]) );
  FD2 \xm_pc_plus_8_reg[14]  ( .D(dx_pc_plus_8[14]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[14]) );
  FD2 \xm_pc_plus_8_reg[13]  ( .D(dx_pc_plus_8[13]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[13]) );
  FD2 \xm_pc_plus_8_reg[12]  ( .D(dx_pc_plus_8[12]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[12]) );
  FD2 \xm_pc_plus_8_reg[11]  ( .D(dx_pc_plus_8[11]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[11]) );
  FD2 \xm_pc_plus_8_reg[10]  ( .D(dx_pc_plus_8[10]), .CP(clock), .CD(n139), 
        .Q(xm_pc_plus_8[10]) );
  FD2 \xm_pc_plus_8_reg[9]  ( .D(dx_pc_plus_8[9]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[9]) );
  FD2 \xm_pc_plus_8_reg[8]  ( .D(dx_pc_plus_8[8]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[8]) );
  FD2 \xm_pc_plus_8_reg[7]  ( .D(dx_pc_plus_8[7]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[7]) );
  FD2 \xm_pc_plus_8_reg[6]  ( .D(dx_pc_plus_8[6]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[6]) );
  FD2 \xm_pc_plus_8_reg[5]  ( .D(dx_pc_plus_8[5]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[5]) );
  FD2 \xm_pc_plus_8_reg[4]  ( .D(dx_pc_plus_8[4]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[4]) );
  FD2 \xm_pc_plus_8_reg[3]  ( .D(dx_pc_plus_8[3]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[3]) );
  FD2 \xm_pc_plus_8_reg[2]  ( .D(dx_pc_plus_8[2]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[2]) );
  FD2 \xm_pc_plus_8_reg[1]  ( .D(dx_pc_plus_8[1]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[1]) );
  FD2 \xm_pc_plus_8_reg[0]  ( .D(dx_pc_plus_8[0]), .CP(clock), .CD(n139), .Q(
        xm_pc_plus_8[0]) );
  FD2 \xm_Inst_reg[25]  ( .D(dx_Inst[25]), .CP(clock), .CD(n139), .Q(
        xm_Inst[25]) );
  FD2 \xm_Inst_reg[24]  ( .D(dx_Inst[24]), .CP(clock), .CD(n139), .Q(
        xm_Inst[24]) );
  FD2 \xm_Inst_reg[23]  ( .D(dx_Inst[23]), .CP(clock), .CD(n139), .Q(
        xm_Inst[23]) );
  FD2 \xm_Inst_reg[22]  ( .D(dx_Inst[22]), .CP(clock), .CD(n139), .Q(
        xm_Inst[22]) );
  FD2 \xm_Inst_reg[21]  ( .D(dx_Inst[21]), .CP(clock), .CD(n139), .Q(
        xm_Inst[21]) );
  FD2 \xm_gpr_rd_data2_reg[31]  ( .D(dx_gpr_rd_data2[31]), .CP(clock), .CD(
        n139), .Q(Din[31]) );
  FD2 \xm_gpr_rd_data2_reg[30]  ( .D(dx_gpr_rd_data2[30]), .CP(clock), .CD(
        n139), .Q(Din[30]) );
  FD2 \xm_gpr_rd_data2_reg[29]  ( .D(dx_gpr_rd_data2[29]), .CP(clock), .CD(
        n139), .Q(Din[29]) );
  FD2 \xm_gpr_rd_data2_reg[28]  ( .D(dx_gpr_rd_data2[28]), .CP(clock), .CD(
        n139), .Q(Din[28]) );
  FD2 \xm_gpr_rd_data2_reg[27]  ( .D(dx_gpr_rd_data2[27]), .CP(clock), .CD(
        n139), .Q(Din[27]) );
  FD2 \xm_gpr_rd_data2_reg[26]  ( .D(dx_gpr_rd_data2[26]), .CP(clock), .CD(
        n139), .Q(Din[26]) );
  FD2 \xm_gpr_rd_data2_reg[25]  ( .D(dx_gpr_rd_data2[25]), .CP(clock), .CD(
        n139), .Q(Din[25]) );
  FD2 \xm_gpr_rd_data2_reg[24]  ( .D(dx_gpr_rd_data2[24]), .CP(clock), .CD(
        n139), .Q(Din[24]) );
  FD2 \xm_gpr_rd_data2_reg[23]  ( .D(dx_gpr_rd_data2[23]), .CP(clock), .CD(
        n139), .Q(Din[23]) );
  FD2 \xm_gpr_rd_data2_reg[22]  ( .D(dx_gpr_rd_data2[22]), .CP(clock), .CD(
        n139), .Q(Din[22]) );
  FD2 \xm_gpr_rd_data2_reg[21]  ( .D(dx_gpr_rd_data2[21]), .CP(clock), .CD(
        n139), .Q(Din[21]) );
  FD2 \xm_gpr_rd_data2_reg[20]  ( .D(dx_gpr_rd_data2[20]), .CP(clock), .CD(
        n139), .Q(Din[20]) );
  FD2 \xm_gpr_rd_data2_reg[19]  ( .D(dx_gpr_rd_data2[19]), .CP(clock), .CD(
        n139), .Q(Din[19]) );
  FD2 \xm_gpr_rd_data2_reg[18]  ( .D(dx_gpr_rd_data2[18]), .CP(clock), .CD(
        n139), .Q(Din[18]) );
  FD2 \xm_gpr_rd_data2_reg[17]  ( .D(dx_gpr_rd_data2[17]), .CP(clock), .CD(
        n139), .Q(Din[17]) );
  FD2 \xm_gpr_rd_data2_reg[16]  ( .D(dx_gpr_rd_data2[16]), .CP(clock), .CD(
        n139), .Q(Din[16]) );
  FD2 \xm_gpr_rd_data2_reg[15]  ( .D(dx_gpr_rd_data2[15]), .CP(clock), .CD(
        n139), .Q(Din[15]) );
  FD2 \xm_gpr_rd_data2_reg[14]  ( .D(dx_gpr_rd_data2[14]), .CP(clock), .CD(
        n139), .Q(Din[14]) );
  FD2 \xm_gpr_rd_data2_reg[13]  ( .D(dx_gpr_rd_data2[13]), .CP(clock), .CD(
        n139), .Q(Din[13]) );
  FD2 \xm_gpr_rd_data2_reg[12]  ( .D(dx_gpr_rd_data2[12]), .CP(clock), .CD(
        n139), .Q(Din[12]) );
  FD2 \xm_gpr_rd_data2_reg[11]  ( .D(dx_gpr_rd_data2[11]), .CP(clock), .CD(
        n139), .Q(Din[11]) );
  FD2 \xm_gpr_rd_data2_reg[10]  ( .D(dx_gpr_rd_data2[10]), .CP(clock), .CD(
        n139), .Q(Din[10]) );
  FD2 \xm_gpr_rd_data2_reg[9]  ( .D(dx_gpr_rd_data2[9]), .CP(clock), .CD(n139), 
        .Q(Din[9]) );
  FD2 \xm_gpr_rd_data2_reg[8]  ( .D(dx_gpr_rd_data2[8]), .CP(clock), .CD(n139), 
        .Q(Din[8]) );
  FD2 \xm_gpr_rd_data2_reg[7]  ( .D(dx_gpr_rd_data2[7]), .CP(clock), .CD(n139), 
        .Q(Din[7]) );
  FD2 \xm_gpr_rd_data2_reg[6]  ( .D(dx_gpr_rd_data2[6]), .CP(clock), .CD(n139), 
        .Q(Din[6]) );
  FD2 \xm_gpr_rd_data2_reg[5]  ( .D(dx_gpr_rd_data2[5]), .CP(clock), .CD(n139), 
        .Q(Din[5]) );
  FD2 \dx_gpr_rd_data1_reg[6]  ( .D(gpr_rd_data1[6]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[6]) );
  FD2 \dx_gpr_rd_data1_reg[9]  ( .D(gpr_rd_data1[9]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[9]) );
  FD2 \dx_gpr_rd_data1_reg[14]  ( .D(gpr_rd_data1[14]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[14]) );
  FD2 \dx_gpr_rd_data1_reg[11]  ( .D(gpr_rd_data1[11]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[11]) );
  FD2 \dx_gpr_rd_data1_reg[19]  ( .D(gpr_rd_data1[19]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[19]) );
  FD2 \dx_gpr_rd_data1_reg[13]  ( .D(gpr_rd_data1[13]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[13]) );
  FD2 \dx_gpr_rd_data1_reg[27]  ( .D(gpr_rd_data1[27]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[27]) );
  FD2 \dx_gpr_rd_data1_reg[30]  ( .D(gpr_rd_data1[30]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[30]) );
  FD2 \dx_gpr_rd_data1_reg[31]  ( .D(gpr_rd_data1[31]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[31]) );
  FD2 \dx_gpr_rd_data1_reg[15]  ( .D(gpr_rd_data1[15]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[15]) );
  FD2 \dx_gpr_rd_data1_reg[7]  ( .D(gpr_rd_data1[7]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[7]) );
  FD2 \dx_gpr_rd_data1_reg[5]  ( .D(gpr_rd_data1[5]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[5]) );
  FD2 \dx_gpr_rd_data1_reg[3]  ( .D(gpr_rd_data1[3]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[3]) );
  FD2 \dx_gpr_rd_data1_reg[8]  ( .D(gpr_rd_data1[8]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[8]) );
  FD2 \dx_gpr_rd_data1_reg[10]  ( .D(gpr_rd_data1[10]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[10]) );
  FD2 \dx_gpr_rd_data1_reg[20]  ( .D(gpr_rd_data1[20]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[20]) );
  FD2 \dx_gpr_rd_data1_reg[12]  ( .D(gpr_rd_data1[12]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[12]) );
  FD2 \dx_gpr_rd_data1_reg[26]  ( .D(gpr_rd_data1[26]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[26]) );
  FD2 \dx_gpr_rd_data1_reg[22]  ( .D(gpr_rd_data1[22]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[22]) );
  FD2 \dx_gpr_rd_data1_reg[29]  ( .D(gpr_rd_data1[29]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[29]) );
  FD2 \dx_gpr_rd_data1_reg[1]  ( .D(gpr_rd_data1[1]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[1]) );
  FD2 \dx_gpr_rd_data1_reg[28]  ( .D(gpr_rd_data1[28]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[28]) );
  FD2 \dx_gpr_rd_data1_reg[25]  ( .D(gpr_rd_data1[25]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[25]) );
  FD2 \dx_gpr_rd_data1_reg[24]  ( .D(gpr_rd_data1[24]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[24]) );
  FD2 \dx_gpr_rd_data1_reg[23]  ( .D(gpr_rd_data1[23]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[23]) );
  FD2 \dx_gpr_rd_data1_reg[21]  ( .D(gpr_rd_data1[21]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[21]) );
  FD2 \dx_gpr_rd_data1_reg[18]  ( .D(gpr_rd_data1[18]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[18]) );
  FD2 \dx_gpr_rd_data1_reg[17]  ( .D(gpr_rd_data1[17]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[17]) );
  FD2 \dx_gpr_rd_data1_reg[16]  ( .D(gpr_rd_data1[16]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[16]) );
  FD2 \dx_gpr_rd_data1_reg[0]  ( .D(gpr_rd_data1[0]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[0]) );
  FD2 \dx_gpr_rd_data1_reg[2]  ( .D(gpr_rd_data1[2]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data1[2]) );
  FD2 \dx_gpr_rd_data2_reg[14]  ( .D(gpr_rd_data2[14]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[14]) );
  FD2 \dx_gpr_rd_data2_reg[23]  ( .D(gpr_rd_data2[23]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[23]) );
  FD2 \dx_gpr_rd_data2_reg[29]  ( .D(gpr_rd_data2[29]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[29]) );
  FD2 \dx_gpr_rd_data2_reg[9]  ( .D(gpr_rd_data2[9]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[9]) );
  FD2 \dx_gpr_rd_data2_reg[0]  ( .D(gpr_rd_data2[0]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_data2[0]) );
  FD2 \dx_gpr_rd_addr1_reg[4]  ( .D(gpr_rd_addr1[4]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_addr1[4]) );
  FD2 \dx_gpr_rd_addr1_reg[3]  ( .D(gpr_rd_addr1[3]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_addr1[3]) );
  FD2 \dx_gpr_rd_addr1_reg[2]  ( .D(gpr_rd_addr1[2]), .CP(clock), .CD(n139), 
        .Q(dx_gpr_rd_addr1[2]) );
  FD2 \dx_Inst_reg[4]  ( .D(n93), .CP(clock), .CD(n139), .Q(dx_Inst_4) );
  FD2 \dx_Inst_reg[2]  ( .D(n90), .CP(clock), .CD(n139), .Q(dx_Inst_2) );
  FD2 \fd_Inst_reg[31]  ( .D(Inst_stall_b_j[31]), .CP(clock), .CD(n139), .Q(
        n111), .QN(n73) );
  B5I U99 ( .A(n38), .Z(Inst_stall_b_j[9]) );
  IVI U100 ( .A(n39), .Z(Inst_stall_b_j[7]) );
  IVI U101 ( .A(n40), .Z(Inst_stall_b_j[5]) );
  IVI U102 ( .A(n41), .Z(Inst_stall_b_j[30]) );
  IVI U103 ( .A(n42), .Z(Inst_stall_b_j[29]) );
  IVI U104 ( .A(n43), .Z(Inst_stall_b_j[27]) );
  IVI U105 ( .A(n44), .Z(Inst_stall_b_j[26]) );
  B5I U106 ( .A(n45), .Z(Inst_stall_b_j[20]) );
  IVI U107 ( .A(n46), .Z(Inst_stall_b_j[1]) );
  IVI U108 ( .A(n47), .Z(Inst_stall_b_j[19]) );
  IVI U109 ( .A(n48), .Z(Inst_stall_b_j[18]) );
  IVI U110 ( .A(n49), .Z(Inst_stall_b_j[17]) );
  IVI U111 ( .A(n50), .Z(Inst_stall_b_j[16]) );
  IVI U112 ( .A(n51), .Z(Inst_stall_b_j[15]) );
  IVI U113 ( .A(n52), .Z(Inst_stall_b_j[14]) );
  IVI U114 ( .A(n53), .Z(Inst_stall_b_j[13]) );
  IVI U115 ( .A(n54), .Z(Inst_stall_b_j[11]) );
  IVI U116 ( .A(n55), .Z(Inst_stall_b_j[10]) );
  IVI U117 ( .A(n56), .Z(Inst_stall_b_j[0]) );
  ND2I U118 ( .A(Inst[9]), .B(n69), .Z(n38) );
  ND2I U119 ( .A(Inst[7]), .B(n113), .Z(n39) );
  ND2I U120 ( .A(Inst[5]), .B(n69), .Z(n40) );
  ND2I U121 ( .A(Inst[30]), .B(n70), .Z(n41) );
  ND2I U122 ( .A(Inst[29]), .B(n69), .Z(n42) );
  ND2I U123 ( .A(Inst[27]), .B(n113), .Z(n43) );
  ND2I U124 ( .A(Inst[26]), .B(n70), .Z(n44) );
  ND2I U125 ( .A(Inst[20]), .B(n115), .Z(n45) );
  ND2I U126 ( .A(Inst[1]), .B(n114), .Z(n46) );
  ND2I U127 ( .A(Inst[19]), .B(n114), .Z(n47) );
  ND2I U128 ( .A(Inst[18]), .B(n115), .Z(n48) );
  ND2I U129 ( .A(Inst[17]), .B(n114), .Z(n49) );
  ND2I U130 ( .A(Inst[16]), .B(n115), .Z(n50) );
  ND2I U131 ( .A(Inst[15]), .B(n113), .Z(n51) );
  ND2I U132 ( .A(Inst[14]), .B(n70), .Z(n52) );
  ND2I U133 ( .A(Inst[13]), .B(n69), .Z(n53) );
  ND2I U134 ( .A(Inst[11]), .B(n113), .Z(n54) );
  ND2I U135 ( .A(Inst[10]), .B(n70), .Z(n55) );
  ND2I U136 ( .A(Inst[0]), .B(n66), .Z(n56) );
  IVI U137 ( .A(n81), .Z(n82) );
  IVDAP U138 ( .A(n93), .Z(n57) );
  B2I U139 ( .A(gpr_wr_addr[4]), .Z2(n58) );
  B2I U140 ( .A(gpr_wr_addr[3]), .Z2(n59) );
  IVI U141 ( .A(n61), .Z(Inst_stall_b_j[6]) );
  IVI U142 ( .A(n62), .Z(Inst_stall_b_j[3]) );
  IVI U143 ( .A(n63), .Z(Inst_stall_b_j[2]) );
  IVI U144 ( .A(n64), .Z(Inst_stall_b_j[22]) );
  IVI U145 ( .A(n65), .Z(Inst_stall_b_j[21]) );
  ND2I U146 ( .A(Inst[6]), .B(n66), .Z(n61) );
  ND2I U147 ( .A(Inst[3]), .B(n114), .Z(n62) );
  ND2I U148 ( .A(Inst[2]), .B(n115), .Z(n63) );
  ND2I U149 ( .A(Inst[22]), .B(n66), .Z(n64) );
  ND2I U150 ( .A(Inst[21]), .B(n66), .Z(n65) );
  IVI U151 ( .A(n67), .Z(n66) );
  ND3P U152 ( .A(n118), .B(n117), .C(n116), .Z(n67) );
  ND3P U153 ( .A(n118), .B(n117), .C(n116), .Z(n68) );
  IVI U154 ( .A(n67), .Z(n114) );
  AN3P U155 ( .A(n118), .B(n117), .C(n116), .Z(n108) );
  IVI U156 ( .A(n68), .Z(n69) );
  IVI U157 ( .A(n68), .Z(n70) );
  IVI U158 ( .A(n71), .Z(n72) );
  IVI U159 ( .A(n73), .Z(n74) );
  IVI U160 ( .A(n60), .Z(fd_Inst_stall[0]) );
  IVI U161 ( .A(n76), .Z(n77) );
  IVI U162 ( .A(gpr_wr_addr[1]), .Z(n78) );
  B5I U163 ( .A(n78), .Z(n79) );
  IVI U164 ( .A(gpr_wr_addr[2]), .Z(n81) );
  IVI U165 ( .A(n84), .Z(n85) );
  IVI U166 ( .A(n86), .Z(n87) );
  IVI U167 ( .A(n88), .Z(n89) );
  IVI U168 ( .A(n31), .Z(n90) );
  IVI U169 ( .A(n89), .Z(fd_Inst_stall[2]) );
  IVI U170 ( .A(n30), .Z(fd_Inst_stall[3]) );
  IVI U171 ( .A(gpr_wr_addr[0]), .Z(n94) );
  B5I U172 ( .A(n94), .Z(n95) );
  IVI U173 ( .A(n96), .Z(n97) );
  IVI U174 ( .A(n98), .Z(n99) );
  IVI U175 ( .A(n100), .Z(n101) );
  IVI U176 ( .A(n102), .Z(n103) );
  IVI U177 ( .A(n104), .Z(n105) );
  IVI U178 ( .A(n106), .Z(n107) );
  IVI U179 ( .A(d_isSLL_SRL), .Z(n109) );
  IVI U180 ( .A(n109), .Z(n110) );
  IVI U181 ( .A(n68), .Z(n113) );
  IVI U182 ( .A(n67), .Z(n115) );
  IVI U183 ( .A(d_PCSrc3), .Z(n118) );
  IVI U184 ( .A(d_PCSrc2), .Z(n117) );
  IVI U185 ( .A(d_PCSrc1), .Z(n116) );
  IVI U186 ( .A(reset), .Z(n139) );
  AN2I U187 ( .A(Inst[23]), .B(n108), .Z(Inst_stall_b_j[23]) );
  AN2I U188 ( .A(Inst[24]), .B(n108), .Z(Inst_stall_b_j[24]) );
  AN2I U189 ( .A(Inst[25]), .B(n108), .Z(Inst_stall_b_j[25]) );
  AN2I U190 ( .A(Inst[4]), .B(n108), .Z(Inst_stall_b_j[4]) );
  IVI U191 ( .A(n6), .Z(fd_Inst_stall[27]) );
  AN2I U192 ( .A(Inst[28]), .B(n108), .Z(Inst_stall_b_j[28]) );
  IVI U193 ( .A(n4), .Z(fd_Inst_stall[29]) );
  AN2I U194 ( .A(Inst[31]), .B(n108), .Z(Inst_stall_b_j[31]) );
  AN2I U195 ( .A(Inst[8]), .B(n108), .Z(Inst_stall_b_j[8]) );
  AN2I U196 ( .A(Inst[12]), .B(n108), .Z(Inst_stall_b_j[12]) );
endmodule

