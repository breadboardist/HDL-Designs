
module sfilt_DW01_add_2 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n83, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n133, n134, n135, n136, n137, n138, n139,
         n140, n142, n145, n146, n147, n148, n149, n150, n151, n153, n154,
         n155, n156, n157, n158, n159, n160, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n179, n180,
         n181, n182, n183, n184, n185, n186, n188, n191, n192, n193, n194,
         n195, n196, n197, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n235,
         n236, n237, n238, n239, n240, n243, n244, n245, n246, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n267, n268, n269, n270, n271, n272, n273, n274,
         n276, n279, n280, n281, n282, n283, n284, n285, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n323, n324, n325, n326, n327, n328, n331,
         n332, n333, n334, n335, n336, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n351, n352, n353, n354, n355, n356, n357,
         n360, n361, n362, n363, n364, n365, n366, n369, n370, n373, n374,
         n375, n376, n379, n380, n381, n382, n383, n384, n385, n386, n389,
         n390, n391, n392, n394, n397, n398, n399, n401, n402, n403, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n425, n426, n427, n428, n429,
         n430, n431, n432, n434, n437, n438, n439, n440, n441, n442, n443,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n481, n482, n483, n484,
         n485, n486, n489, n490, n491, n492, n493, n494, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n509, n510, n511, n512,
         n513, n514, n515, n518, n519, n520, n521, n522, n523, n524, n527,
         n528, n531, n532, n533, n534, n537, n538, n539, n540, n541, n542,
         n543, n544, n547, n548, n549, n550, n552, n555, n556, n557, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n574, n575, n576, n577, n578, n579, n580, n583, n584,
         n585, n586, n588, n589, n590, n591, n592, n593, n594, n595, n598,
         n599, n600, n601, n602, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n915, n916, n917;

  COND1X1 U123 ( .A(n163), .B(n206), .C(n164), .Z(n5) );
  COND1X1 U347 ( .A(n339), .B(n374), .C(n340), .Z(n334) );
  COND1X1 U553 ( .A(n497), .B(n532), .C(n498), .Z(n492) );
  COND1X1 U723 ( .A(n619), .B(n639), .C(n620), .Z(n618) );
  CANR1XL U784 ( .A(n492), .B(n407), .C(n408), .Z(n406) );
  CNIVX4 U785 ( .A(n2), .Z(n917) );
  CNR2XL U786 ( .A(n486), .B(n481), .Z(n475) );
  CNR2XL U787 ( .A(n222), .B(n213), .Z(n211) );
  CNR2XL U788 ( .A(n544), .B(n539), .Z(n537) );
  CNR2XL U789 ( .A(B[24]), .B(A[24]), .Z(n486) );
  CND2XL U790 ( .A(B[2]), .B(A[2]), .Z(n646) );
  CND2X1 U791 ( .A(B[36]), .B(A[36]), .Z(n369) );
  CNR2XL U792 ( .A(n615), .B(n612), .Z(n610) );
  CNR2XL U793 ( .A(n560), .B(n555), .Z(n549) );
  CNR2XL U794 ( .A(B[40]), .B(A[40]), .Z(n328) );
  CNR2XL U795 ( .A(B[16]), .B(A[16]), .Z(n560) );
  CNR2XL U796 ( .A(B[28]), .B(A[28]), .Z(n446) );
  CNR2X1 U797 ( .A(n592), .B(n566), .Z(n564) );
  CNR2X1 U798 ( .A(n589), .B(n584), .Z(n580) );
  COND1XL U799 ( .A(n251), .B(n294), .C(n252), .Z(n250) );
  CANR1XL U800 ( .A(n140), .B(n119), .C(n120), .Z(n118) );
  CANR1XL U801 ( .A(n648), .B(n640), .C(n641), .Z(n639) );
  COND1XL U802 ( .A(n561), .B(n555), .C(n556), .Z(n550) );
  COND1XL U803 ( .A(n447), .B(n437), .C(n438), .Z(n432) );
  CNR2X1 U804 ( .A(B[44]), .B(A[44]), .Z(n288) );
  CNR2XL U805 ( .A(n4), .B(n159), .Z(n157) );
  CNR2XL U806 ( .A(n4), .B(n89), .Z(n87) );
  CNR2XL U807 ( .A(n4), .B(n113), .Z(n111) );
  CND2XL U808 ( .A(n6), .B(n91), .Z(n89) );
  CND2XL U809 ( .A(n6), .B(n115), .Z(n113) );
  CNR2XL U810 ( .A(n335), .B(n260), .Z(n258) );
  CNR2XL U811 ( .A(n493), .B(n418), .Z(n416) );
  CANR1X1 U812 ( .A(n618), .B(n564), .C(n565), .Z(n563) );
  COND1X1 U813 ( .A(n405), .B(n563), .C(n406), .Z(n2) );
  CND2XL U814 ( .A(n375), .B(n357), .Z(n355) );
  CND2XL U815 ( .A(n533), .B(n515), .Z(n513) );
  CND2XL U816 ( .A(n6), .B(n128), .Z(n126) );
  CND2XL U817 ( .A(n6), .B(n139), .Z(n137) );
  CND2XL U818 ( .A(n6), .B(n660), .Z(n150) );
  CND2XL U819 ( .A(n229), .B(n666), .Z(n218) );
  CND2XL U820 ( .A(n174), .B(n207), .Z(n172) );
  CND2XL U821 ( .A(n207), .B(n185), .Z(n183) );
  CND2XL U822 ( .A(n453), .B(n431), .Z(n429) );
  CANR1X1 U823 ( .A(n230), .B(n211), .C(n212), .Z(n206) );
  CANR1X1 U824 ( .A(n392), .B(n379), .C(n380), .Z(n374) );
  CANR1X1 U825 ( .A(n550), .B(n537), .C(n538), .Z(n532) );
  CNR2XL U826 ( .A(n645), .B(n642), .Z(n640) );
  CANR1X1 U827 ( .A(n611), .B(n598), .C(n599), .Z(n593) );
  CANR1X1 U828 ( .A(n476), .B(n457), .C(n458), .Z(n452) );
  CNR2XL U829 ( .A(n328), .B(n323), .Z(n317) );
  CNR2XL U830 ( .A(n154), .B(n145), .Z(n139) );
  CNR2XL U831 ( .A(n288), .B(n279), .Z(n273) );
  CNR2XL U832 ( .A(n106), .B(n97), .Z(n95) );
  CNR2XL U833 ( .A(n626), .B(n623), .Z(n621) );
  CND2XL U834 ( .A(n629), .B(n621), .Z(n619) );
  CNR2XL U835 ( .A(n402), .B(n397), .Z(n391) );
  CNR2XL U836 ( .A(n605), .B(n600), .Z(n598) );
  CNR2XL U837 ( .A(n468), .B(n459), .Z(n457) );
  CNR2XL U838 ( .A(n575), .B(n570), .Z(n568) );
  CNR2XL U839 ( .A(n386), .B(n381), .Z(n379) );
  CNR2XL U840 ( .A(n310), .B(n301), .Z(n299) );
  CNR2XL U841 ( .A(n422), .B(n413), .Z(n411) );
  CNR2XL U842 ( .A(n348), .B(n343), .Z(n341) );
  CNR2XL U843 ( .A(n264), .B(n255), .Z(n253) );
  CNR2XL U844 ( .A(n130), .B(n121), .Z(n119) );
  CNR2XL U845 ( .A(n636), .B(n631), .Z(n629) );
  CNR2IXL U846 ( .B(n139), .A(n130), .Z(n128) );
  CNR2XL U847 ( .A(n355), .B(n348), .Z(n346) );
  CNR2XL U848 ( .A(n513), .B(n506), .Z(n504) );
  CNR2XL U849 ( .A(B[8]), .B(A[8]), .Z(n615) );
  CNR2XL U850 ( .A(B[4]), .B(A[4]), .Z(n636) );
  CNR2XL U851 ( .A(B[32]), .B(A[32]), .Z(n402) );
  CNR2XL U852 ( .A(B[56]), .B(A[56]), .Z(n154) );
  CND2XL U853 ( .A(B[18]), .B(A[18]), .Z(n547) );
  CND2XL U854 ( .A(B[22]), .B(A[22]), .Z(n509) );
  CND2XL U855 ( .A(B[6]), .B(A[6]), .Z(n627) );
  CND2XL U856 ( .A(B[30]), .B(A[30]), .Z(n425) );
  CND2XL U857 ( .A(B[34]), .B(A[34]), .Z(n389) );
  CND2XL U858 ( .A(B[58]), .B(A[58]), .Z(n133) );
  CND2XL U859 ( .A(B[46]), .B(A[46]), .Z(n267) );
  CND2XL U860 ( .A(B[38]), .B(A[38]), .Z(n351) );
  CND2XL U861 ( .A(B[1]), .B(A[1]), .Z(n650) );
  CEOXL U862 ( .A(n22), .B(n244), .Z(SUM[48]) );
  CEOXL U863 ( .A(n23), .B(n257), .Z(SUM[47]) );
  CEOXL U864 ( .A(n24), .B(n268), .Z(SUM[46]) );
  CEOXL U865 ( .A(n25), .B(n281), .Z(SUM[45]) );
  CEOXL U866 ( .A(n26), .B(n290), .Z(SUM[44]) );
  CEOXL U867 ( .A(n27), .B(n303), .Z(SUM[43]) );
  CEOXL U868 ( .A(n28), .B(n312), .Z(SUM[42]) );
  CEOXL U869 ( .A(n29), .B(n325), .Z(SUM[41]) );
  CEOXL U870 ( .A(n30), .B(n332), .Z(SUM[40]) );
  CEOXL U871 ( .A(n31), .B(n345), .Z(SUM[39]) );
  CEOXL U872 ( .A(n32), .B(n352), .Z(SUM[38]) );
  CEOXL U873 ( .A(n33), .B(n363), .Z(SUM[37]) );
  CEOXL U874 ( .A(n34), .B(n370), .Z(SUM[36]) );
  CEOXL U875 ( .A(n35), .B(n383), .Z(SUM[35]) );
  CEOXL U876 ( .A(n36), .B(n390), .Z(SUM[34]) );
  CEOXL U877 ( .A(n37), .B(n399), .Z(SUM[33]) );
  CEOXL U878 ( .A(n7), .B(n73), .Z(SUM[63]) );
  CEOXL U879 ( .A(n8), .B(n86), .Z(SUM[62]) );
  CEOXL U880 ( .A(n9), .B(n99), .Z(SUM[61]) );
  CEOXL U881 ( .A(n10), .B(n110), .Z(SUM[60]) );
  CEOXL U882 ( .A(n11), .B(n123), .Z(SUM[59]) );
  CEOXL U883 ( .A(n12), .B(n134), .Z(SUM[58]) );
  CEOXL U884 ( .A(n13), .B(n147), .Z(SUM[57]) );
  CEOXL U885 ( .A(n14), .B(n156), .Z(SUM[56]) );
  CEOXL U886 ( .A(n15), .B(n169), .Z(SUM[55]) );
  CEOXL U887 ( .A(n16), .B(n180), .Z(SUM[54]) );
  CEOXL U888 ( .A(n17), .B(n193), .Z(SUM[53]) );
  CEOXL U889 ( .A(n18), .B(n202), .Z(SUM[52]) );
  CEOXL U890 ( .A(n19), .B(n215), .Z(SUM[51]) );
  CEOXL U891 ( .A(n20), .B(n224), .Z(SUM[50]) );
  CEOXL U892 ( .A(n21), .B(n237), .Z(SUM[49]) );
  CEOXL U893 ( .A(n39), .B(n415), .Z(SUM[31]) );
  CEOXL U894 ( .A(n40), .B(n426), .Z(SUM[30]) );
  CEOXL U895 ( .A(n41), .B(n439), .Z(SUM[29]) );
  CEOXL U896 ( .A(n42), .B(n448), .Z(SUM[28]) );
  CEOXL U897 ( .A(n43), .B(n461), .Z(SUM[27]) );
  CEOXL U898 ( .A(n44), .B(n470), .Z(SUM[26]) );
  CEOXL U899 ( .A(n45), .B(n483), .Z(SUM[25]) );
  CEOXL U900 ( .A(n46), .B(n490), .Z(SUM[24]) );
  CEOXL U901 ( .A(n47), .B(n503), .Z(SUM[23]) );
  CEOXL U902 ( .A(n48), .B(n510), .Z(SUM[22]) );
  CEOXL U903 ( .A(n49), .B(n521), .Z(SUM[21]) );
  CEOXL U904 ( .A(n50), .B(n528), .Z(SUM[20]) );
  CEOXL U905 ( .A(n51), .B(n541), .Z(SUM[19]) );
  CEOXL U906 ( .A(n52), .B(n548), .Z(SUM[18]) );
  CEOXL U907 ( .A(n53), .B(n557), .Z(SUM[17]) );
  CEOXL U908 ( .A(n55), .B(n572), .Z(SUM[15]) );
  CEOXL U909 ( .A(n57), .B(n586), .Z(SUM[13]) );
  CEOXL U910 ( .A(n59), .B(n602), .Z(SUM[11]) );
  CEOXL U911 ( .A(n64), .B(n628), .Z(SUM[6]) );
  CND2IXL U912 ( .B(n651), .A(n652), .Z(n70) );
  CND2X1 U913 ( .A(n333), .B(n249), .Z(n4) );
  CNR2XL U914 ( .A(n4), .B(n76), .Z(n74) );
  CNR2X1 U915 ( .A(n205), .B(n163), .Z(n6) );
  CNR2X1 U916 ( .A(n373), .B(n339), .Z(n333) );
  CNR2X1 U917 ( .A(n293), .B(n251), .Z(n249) );
  CIVX2 U918 ( .A(n563), .Z(n562) );
  CNR2X1 U919 ( .A(n531), .B(n497), .Z(n491) );
  CNR2X1 U920 ( .A(n117), .B(n93), .Z(n91) );
  CNR2X1 U921 ( .A(n451), .B(n409), .Z(n407) );
  CNR2XL U922 ( .A(n4), .B(n102), .Z(n100) );
  CNR2XL U923 ( .A(n4), .B(n126), .Z(n124) );
  CNR2XL U924 ( .A(n4), .B(n137), .Z(n135) );
  CNR2XL U925 ( .A(n4), .B(n150), .Z(n148) );
  CNR2XL U926 ( .A(n4), .B(n172), .Z(n170) );
  CNR2XL U927 ( .A(n4), .B(n183), .Z(n181) );
  CNR2XL U928 ( .A(n4), .B(n196), .Z(n194) );
  CNR2XL U929 ( .A(n4), .B(n205), .Z(n203) );
  CNR2XL U930 ( .A(n4), .B(n218), .Z(n216) );
  CNR2XL U931 ( .A(n4), .B(n227), .Z(n225) );
  CNR2XL U932 ( .A(n335), .B(n271), .Z(n269) );
  CNR2XL U933 ( .A(n335), .B(n284), .Z(n282) );
  CNR2XL U934 ( .A(n335), .B(n293), .Z(n291) );
  CNR2XL U935 ( .A(n335), .B(n306), .Z(n304) );
  CNR2XL U936 ( .A(n335), .B(n315), .Z(n313) );
  CNR2XL U937 ( .A(n493), .B(n429), .Z(n427) );
  CNR2XL U938 ( .A(n493), .B(n442), .Z(n440) );
  CNR2XL U939 ( .A(n493), .B(n451), .Z(n449) );
  CNR2XL U940 ( .A(n493), .B(n464), .Z(n462) );
  CNR2XL U941 ( .A(n493), .B(n473), .Z(n471) );
  CND2XL U942 ( .A(n6), .B(n78), .Z(n76) );
  CANR1XL U943 ( .A(n629), .B(n638), .C(n630), .Z(n628) );
  COND1XL U944 ( .A(n578), .B(n617), .C(n579), .Z(n577) );
  CND2X1 U945 ( .A(n594), .B(n580), .Z(n578) );
  CANR1XL U946 ( .A(n580), .B(n595), .C(n583), .Z(n579) );
  COND1XL U947 ( .A(n592), .B(n617), .C(n593), .Z(n591) );
  COND1XL U948 ( .A(n608), .B(n617), .C(n609), .Z(n607) );
  COND1XL U949 ( .A(n566), .B(n593), .C(n567), .Z(n565) );
  CND2X1 U950 ( .A(n580), .B(n568), .Z(n566) );
  CANR1XL U951 ( .A(n357), .B(n376), .C(n360), .Z(n356) );
  CANR1XL U952 ( .A(n515), .B(n534), .C(n518), .Z(n514) );
  CND2XL U953 ( .A(n491), .B(n407), .Z(n405) );
  CNR2X1 U954 ( .A(n117), .B(n80), .Z(n78) );
  CND2X1 U955 ( .A(n139), .B(n119), .Z(n117) );
  COND1XL U956 ( .A(n89), .B(n3), .C(n90), .Z(n88) );
  CANR1XL U957 ( .A(n91), .B(n5), .C(n92), .Z(n90) );
  COND1XL U958 ( .A(n93), .B(n118), .C(n94), .Z(n92) );
  COND1XL U959 ( .A(n113), .B(n3), .C(n114), .Z(n112) );
  CANR1XL U960 ( .A(n115), .B(n5), .C(n116), .Z(n114) );
  COND1XL U961 ( .A(n137), .B(n3), .C(n138), .Z(n136) );
  CANR1XL U962 ( .A(n139), .B(n5), .C(n140), .Z(n138) );
  COND1XL U963 ( .A(n159), .B(n3), .C(n160), .Z(n158) );
  COND1XL U964 ( .A(n183), .B(n3), .C(n184), .Z(n182) );
  CANR1XL U965 ( .A(n185), .B(n208), .C(n186), .Z(n184) );
  COND1XL U966 ( .A(n205), .B(n3), .C(n206), .Z(n204) );
  COND1XL U967 ( .A(n227), .B(n3), .C(n228), .Z(n226) );
  COND1XL U968 ( .A(n271), .B(n336), .C(n272), .Z(n270) );
  CANR1XL U969 ( .A(n273), .B(n296), .C(n274), .Z(n272) );
  COND1XL U970 ( .A(n293), .B(n336), .C(n294), .Z(n292) );
  COND1XL U971 ( .A(n315), .B(n336), .C(n316), .Z(n314) );
  COND1XL U972 ( .A(n429), .B(n494), .C(n430), .Z(n428) );
  CANR1XL U973 ( .A(n431), .B(n454), .C(n432), .Z(n430) );
  COND1XL U974 ( .A(n451), .B(n494), .C(n452), .Z(n450) );
  COND1XL U975 ( .A(n473), .B(n494), .C(n474), .Z(n472) );
  CND2X1 U976 ( .A(n229), .B(n211), .Z(n205) );
  CND2X1 U977 ( .A(n475), .B(n457), .Z(n451) );
  CND2X1 U978 ( .A(n317), .B(n299), .Z(n293) );
  CND2X1 U979 ( .A(n549), .B(n537), .Z(n531) );
  CND2X1 U980 ( .A(n391), .B(n379), .Z(n373) );
  CND2X1 U981 ( .A(n610), .B(n598), .Z(n592) );
  CND2X1 U982 ( .A(n515), .B(n499), .Z(n497) );
  CND2X1 U983 ( .A(n185), .B(n165), .Z(n163) );
  CND2X1 U984 ( .A(n357), .B(n341), .Z(n339) );
  CND2X1 U985 ( .A(n273), .B(n253), .Z(n251) );
  CND2X1 U986 ( .A(n431), .B(n411), .Z(n409) );
  CND2X1 U987 ( .A(n317), .B(n674), .Z(n306) );
  CND2X1 U988 ( .A(n475), .B(n690), .Z(n464) );
  CND2XL U989 ( .A(n6), .B(n104), .Z(n102) );
  CND2X1 U990 ( .A(n207), .B(n664), .Z(n196) );
  CND2X1 U991 ( .A(n295), .B(n273), .Z(n271) );
  CND2X1 U992 ( .A(n295), .B(n672), .Z(n284) );
  CND2X1 U993 ( .A(n453), .B(n688), .Z(n442) );
  CND2X1 U994 ( .A(n262), .B(n295), .Z(n260) );
  CND2X1 U995 ( .A(n420), .B(n453), .Z(n418) );
  CANR1XL U996 ( .A(n274), .B(n253), .C(n254), .Z(n252) );
  COND1XL U997 ( .A(n267), .B(n255), .C(n256), .Z(n254) );
  CANR1XL U998 ( .A(n186), .B(n165), .C(n166), .Z(n164) );
  COND1XL U999 ( .A(n179), .B(n167), .C(n168), .Z(n166) );
  COND1XL U1000 ( .A(n133), .B(n121), .C(n122), .Z(n120) );
  CANR1XL U1001 ( .A(n360), .B(n341), .C(n342), .Z(n340) );
  COND1XL U1002 ( .A(n351), .B(n343), .C(n344), .Z(n342) );
  COND1XL U1003 ( .A(n606), .B(n600), .C(n601), .Z(n599) );
  CANR1XL U1004 ( .A(n318), .B(n299), .C(n300), .Z(n294) );
  COND1XL U1005 ( .A(n311), .B(n301), .C(n302), .Z(n300) );
  COND1XL U1006 ( .A(n469), .B(n459), .C(n460), .Z(n458) );
  COND1XL U1007 ( .A(n223), .B(n213), .C(n214), .Z(n212) );
  COND1XL U1008 ( .A(n547), .B(n539), .C(n540), .Z(n538) );
  COND1XL U1009 ( .A(n389), .B(n381), .C(n382), .Z(n380) );
  CANR1XL U1010 ( .A(n518), .B(n499), .C(n500), .Z(n498) );
  COND1XL U1011 ( .A(n509), .B(n501), .C(n502), .Z(n500) );
  COND1XL U1012 ( .A(n289), .B(n279), .C(n280), .Z(n274) );
  COND1XL U1013 ( .A(n403), .B(n397), .C(n398), .Z(n392) );
  COND1XL U1014 ( .A(n201), .B(n191), .C(n192), .Z(n186) );
  COND1XL U1015 ( .A(n155), .B(n145), .C(n146), .Z(n140) );
  COND1XL U1016 ( .A(n331), .B(n323), .C(n324), .Z(n318) );
  COND1XL U1017 ( .A(n489), .B(n481), .C(n482), .Z(n476) );
  COND1XL U1018 ( .A(n243), .B(n235), .C(n236), .Z(n230) );
  COND1XL U1019 ( .A(n646), .B(n642), .C(n643), .Z(n641) );
  CNR2X1 U1020 ( .A(n200), .B(n191), .Z(n185) );
  CNR2X1 U1021 ( .A(n446), .B(n437), .Z(n431) );
  CANR1XL U1022 ( .A(n630), .B(n621), .C(n622), .Z(n620) );
  COND1XL U1023 ( .A(n652), .B(n649), .C(n650), .Z(n648) );
  COND1XL U1024 ( .A(n616), .B(n612), .C(n613), .Z(n611) );
  COND1XL U1025 ( .A(n109), .B(n97), .C(n98), .Z(n96) );
  CNR2X1 U1026 ( .A(n240), .B(n235), .Z(n229) );
  CNR2X1 U1027 ( .A(n524), .B(n519), .Z(n515) );
  CNR2X1 U1028 ( .A(n366), .B(n361), .Z(n357) );
  COND1XL U1029 ( .A(n527), .B(n519), .C(n520), .Z(n518) );
  COND1XL U1030 ( .A(n637), .B(n631), .C(n632), .Z(n630) );
  COND1XL U1031 ( .A(n369), .B(n361), .C(n362), .Z(n360) );
  COND1XL U1032 ( .A(n590), .B(n584), .C(n585), .Z(n583) );
  CANR1XL U1033 ( .A(n583), .B(n568), .C(n569), .Z(n567) );
  COND1XL U1034 ( .A(n576), .B(n570), .C(n571), .Z(n569) );
  CNR2X1 U1035 ( .A(n117), .B(n106), .Z(n104) );
  CNR2X1 U1036 ( .A(n506), .B(n501), .Z(n499) );
  CNR2X1 U1037 ( .A(n176), .B(n167), .Z(n165) );
  COND1XL U1038 ( .A(n409), .B(n452), .C(n410), .Z(n408) );
  CANR1XL U1039 ( .A(n432), .B(n411), .C(n412), .Z(n410) );
  COND1XL U1040 ( .A(n425), .B(n413), .C(n414), .Z(n412) );
  COND1XL U1041 ( .A(n627), .B(n623), .C(n624), .Z(n622) );
  COND1XL U1042 ( .A(n76), .B(n3), .C(n77), .Z(n75) );
  CANR1XL U1043 ( .A(n78), .B(n5), .C(n79), .Z(n77) );
  COND1XL U1044 ( .A(n80), .B(n118), .C(n81), .Z(n79) );
  CANR1XL U1045 ( .A(n915), .B(n96), .C(n83), .Z(n81) );
  COND1XL U1046 ( .A(n102), .B(n3), .C(n103), .Z(n101) );
  CANR1XL U1047 ( .A(n104), .B(n5), .C(n105), .Z(n103) );
  COND1XL U1048 ( .A(n106), .B(n118), .C(n109), .Z(n105) );
  COND1XL U1049 ( .A(n126), .B(n3), .C(n127), .Z(n125) );
  CANR1XL U1050 ( .A(n128), .B(n5), .C(n129), .Z(n127) );
  COND1XL U1051 ( .A(n130), .B(n142), .C(n133), .Z(n129) );
  COND1XL U1052 ( .A(n150), .B(n3), .C(n151), .Z(n149) );
  CANR1XL U1053 ( .A(n660), .B(n5), .C(n153), .Z(n151) );
  COND1XL U1054 ( .A(n172), .B(n3), .C(n173), .Z(n171) );
  CANR1XL U1055 ( .A(n208), .B(n174), .C(n175), .Z(n173) );
  COND1XL U1056 ( .A(n176), .B(n188), .C(n179), .Z(n175) );
  COND1XL U1057 ( .A(n196), .B(n3), .C(n197), .Z(n195) );
  CANR1XL U1058 ( .A(n664), .B(n208), .C(n199), .Z(n197) );
  COND1XL U1059 ( .A(n218), .B(n3), .C(n219), .Z(n217) );
  CANR1XL U1060 ( .A(n666), .B(n230), .C(n221), .Z(n219) );
  COND1XL U1061 ( .A(n240), .B(n3), .C(n243), .Z(n239) );
  COND1XL U1062 ( .A(n366), .B(n374), .C(n369), .Z(n365) );
  COND1XL U1063 ( .A(n386), .B(n394), .C(n389), .Z(n385) );
  COND1XL U1064 ( .A(n524), .B(n532), .C(n527), .Z(n523) );
  COND1XL U1065 ( .A(n544), .B(n552), .C(n547), .Z(n543) );
  COND1XL U1066 ( .A(n260), .B(n336), .C(n261), .Z(n259) );
  CANR1XL U1067 ( .A(n296), .B(n262), .C(n263), .Z(n261) );
  COND1XL U1068 ( .A(n264), .B(n276), .C(n267), .Z(n263) );
  COND1XL U1069 ( .A(n284), .B(n336), .C(n285), .Z(n283) );
  CANR1XL U1070 ( .A(n672), .B(n296), .C(n287), .Z(n285) );
  COND1XL U1071 ( .A(n306), .B(n336), .C(n307), .Z(n305) );
  CANR1XL U1072 ( .A(n674), .B(n318), .C(n309), .Z(n307) );
  COND1XL U1073 ( .A(n328), .B(n336), .C(n331), .Z(n327) );
  COND1XL U1074 ( .A(n418), .B(n494), .C(n419), .Z(n417) );
  CANR1XL U1075 ( .A(n454), .B(n420), .C(n421), .Z(n419) );
  COND1XL U1076 ( .A(n422), .B(n434), .C(n425), .Z(n421) );
  COND1XL U1077 ( .A(n442), .B(n494), .C(n443), .Z(n441) );
  CANR1XL U1078 ( .A(n688), .B(n454), .C(n445), .Z(n443) );
  COND1XL U1079 ( .A(n464), .B(n494), .C(n465), .Z(n463) );
  CANR1XL U1080 ( .A(n690), .B(n476), .C(n467), .Z(n465) );
  COND1XL U1081 ( .A(n486), .B(n494), .C(n489), .Z(n485) );
  COND1XL U1082 ( .A(n348), .B(n356), .C(n351), .Z(n347) );
  COND1XL U1083 ( .A(n506), .B(n514), .C(n509), .Z(n505) );
  CNR2IXL U1084 ( .B(n185), .A(n176), .Z(n174) );
  CNR2IXL U1085 ( .B(n273), .A(n264), .Z(n262) );
  CNR2IXL U1086 ( .B(n431), .A(n422), .Z(n420) );
  CNR2XL U1087 ( .A(n373), .B(n366), .Z(n364) );
  CNR2XL U1088 ( .A(n531), .B(n524), .Z(n522) );
  CNR2XL U1089 ( .A(n4), .B(n240), .Z(n238) );
  CNR2XL U1090 ( .A(n335), .B(n328), .Z(n326) );
  CNR2XL U1091 ( .A(n493), .B(n486), .Z(n484) );
  CNR2IXL U1092 ( .B(n391), .A(n386), .Z(n384) );
  CNR2IXL U1093 ( .B(n549), .A(n544), .Z(n542) );
  CND2X1 U1094 ( .A(n95), .B(n915), .Z(n80) );
  CNR2X1 U1095 ( .A(B[48]), .B(A[48]), .Z(n240) );
  CNR2X1 U1096 ( .A(B[20]), .B(A[20]), .Z(n524) );
  CNR2X1 U1097 ( .A(B[34]), .B(A[34]), .Z(n386) );
  CNR2X1 U1098 ( .A(B[18]), .B(A[18]), .Z(n544) );
  CNR2X1 U1099 ( .A(B[22]), .B(A[22]), .Z(n506) );
  CNR2X1 U1100 ( .A(B[46]), .B(A[46]), .Z(n264) );
  CNR2X1 U1101 ( .A(B[38]), .B(A[38]), .Z(n348) );
  CNR2X1 U1102 ( .A(B[36]), .B(A[36]), .Z(n366) );
  CNR2X1 U1103 ( .A(B[54]), .B(A[54]), .Z(n176) );
  CNR2X1 U1104 ( .A(B[30]), .B(A[30]), .Z(n422) );
  CNR2X1 U1105 ( .A(B[58]), .B(A[58]), .Z(n130) );
  CNR2X1 U1106 ( .A(B[60]), .B(A[60]), .Z(n106) );
  CNR2X1 U1107 ( .A(B[47]), .B(A[47]), .Z(n255) );
  CNR2X1 U1108 ( .A(B[23]), .B(A[23]), .Z(n501) );
  CNR2X1 U1109 ( .A(B[41]), .B(A[41]), .Z(n323) );
  CNR2X1 U1110 ( .A(B[45]), .B(A[45]), .Z(n279) );
  CNR2X1 U1111 ( .A(B[25]), .B(A[25]), .Z(n481) );
  CNR2X1 U1112 ( .A(B[49]), .B(A[49]), .Z(n235) );
  CNR2X1 U1113 ( .A(B[17]), .B(A[17]), .Z(n555) );
  CNR2X1 U1114 ( .A(B[35]), .B(A[35]), .Z(n381) );
  CNR2X1 U1115 ( .A(B[11]), .B(A[11]), .Z(n600) );
  CNR2X1 U1116 ( .A(B[21]), .B(A[21]), .Z(n519) );
  CNR2X1 U1117 ( .A(B[19]), .B(A[19]), .Z(n539) );
  CNR2X1 U1118 ( .A(B[53]), .B(A[53]), .Z(n191) );
  CNR2X1 U1119 ( .A(B[43]), .B(A[43]), .Z(n301) );
  CNR2X1 U1120 ( .A(B[39]), .B(A[39]), .Z(n343) );
  CNR2X1 U1121 ( .A(B[29]), .B(A[29]), .Z(n437) );
  CNR2X1 U1122 ( .A(B[33]), .B(A[33]), .Z(n397) );
  CNR2X1 U1123 ( .A(B[15]), .B(A[15]), .Z(n570) );
  CNR2X1 U1124 ( .A(B[27]), .B(A[27]), .Z(n459) );
  CNR2X1 U1125 ( .A(B[37]), .B(A[37]), .Z(n361) );
  CNR2X1 U1126 ( .A(B[13]), .B(A[13]), .Z(n584) );
  CNR2X1 U1127 ( .A(B[51]), .B(A[51]), .Z(n213) );
  CNR2X1 U1128 ( .A(B[9]), .B(A[9]), .Z(n612) );
  CNR2X1 U1129 ( .A(B[31]), .B(A[31]), .Z(n413) );
  CNR2X1 U1130 ( .A(B[7]), .B(A[7]), .Z(n623) );
  CNR2X1 U1131 ( .A(B[55]), .B(A[55]), .Z(n167) );
  CNR2X1 U1132 ( .A(B[5]), .B(A[5]), .Z(n631) );
  CNR2X1 U1133 ( .A(B[57]), .B(A[57]), .Z(n145) );
  CNR2X1 U1134 ( .A(B[3]), .B(A[3]), .Z(n642) );
  CNR2X1 U1135 ( .A(B[59]), .B(A[59]), .Z(n121) );
  CNR2X1 U1136 ( .A(B[61]), .B(A[61]), .Z(n97) );
  CNR2X1 U1137 ( .A(B[6]), .B(A[6]), .Z(n626) );
  CNR2X1 U1138 ( .A(B[2]), .B(A[2]), .Z(n645) );
  CNR2X1 U1139 ( .A(B[52]), .B(A[52]), .Z(n200) );
  CNR2X1 U1140 ( .A(B[42]), .B(A[42]), .Z(n310) );
  CNR2X1 U1141 ( .A(B[50]), .B(A[50]), .Z(n222) );
  CNR2X1 U1142 ( .A(B[26]), .B(A[26]), .Z(n468) );
  CNR2X1 U1143 ( .A(B[10]), .B(A[10]), .Z(n605) );
  CNR2X1 U1144 ( .A(B[12]), .B(A[12]), .Z(n589) );
  CNR2X1 U1145 ( .A(B[14]), .B(A[14]), .Z(n575) );
  CND2X1 U1146 ( .A(B[0]), .B(A[0]), .Z(n652) );
  CNR2X1 U1147 ( .A(B[1]), .B(A[1]), .Z(n649) );
  COR2X1 U1148 ( .A(B[62]), .B(A[62]), .Z(n915) );
  CNR2XL U1149 ( .A(B[0]), .B(A[0]), .Z(n651) );
  COR2X1 U1150 ( .A(B[63]), .B(A[63]), .Z(n916) );
  CND2X1 U1151 ( .A(B[16]), .B(A[16]), .Z(n561) );
  CND2X1 U1152 ( .A(B[10]), .B(A[10]), .Z(n606) );
  CND2X1 U1153 ( .A(B[32]), .B(A[32]), .Z(n403) );
  CND2X1 U1154 ( .A(B[44]), .B(A[44]), .Z(n289) );
  CND2X1 U1155 ( .A(B[42]), .B(A[42]), .Z(n311) );
  CND2X1 U1156 ( .A(B[4]), .B(A[4]), .Z(n637) );
  CND2X1 U1157 ( .A(B[26]), .B(A[26]), .Z(n469) );
  CND2X1 U1158 ( .A(B[28]), .B(A[28]), .Z(n447) );
  CND2X1 U1159 ( .A(B[14]), .B(A[14]), .Z(n576) );
  CND2X1 U1160 ( .A(B[12]), .B(A[12]), .Z(n590) );
  CND2X1 U1161 ( .A(B[50]), .B(A[50]), .Z(n223) );
  CND2X1 U1162 ( .A(B[52]), .B(A[52]), .Z(n201) );
  CND2X1 U1163 ( .A(B[56]), .B(A[56]), .Z(n155) );
  CND2X1 U1164 ( .A(B[40]), .B(A[40]), .Z(n331) );
  CND2X1 U1165 ( .A(B[8]), .B(A[8]), .Z(n616) );
  CND2X1 U1166 ( .A(B[24]), .B(A[24]), .Z(n489) );
  CND2X1 U1167 ( .A(B[48]), .B(A[48]), .Z(n243) );
  CND2XL U1168 ( .A(B[20]), .B(A[20]), .Z(n527) );
  CND2XL U1169 ( .A(B[54]), .B(A[54]), .Z(n179) );
  CND2X1 U1170 ( .A(B[60]), .B(A[60]), .Z(n109) );
  CND2X1 U1171 ( .A(B[62]), .B(A[62]), .Z(n85) );
  CND2XL U1172 ( .A(B[47]), .B(A[47]), .Z(n256) );
  CND2XL U1173 ( .A(B[23]), .B(A[23]), .Z(n502) );
  CND2XL U1174 ( .A(B[11]), .B(A[11]), .Z(n601) );
  CND2XL U1175 ( .A(B[33]), .B(A[33]), .Z(n398) );
  CND2XL U1176 ( .A(B[45]), .B(A[45]), .Z(n280) );
  CND2XL U1177 ( .A(B[41]), .B(A[41]), .Z(n324) );
  CND2XL U1178 ( .A(B[17]), .B(A[17]), .Z(n556) );
  CND2XL U1179 ( .A(B[9]), .B(A[9]), .Z(n613) );
  CND2XL U1180 ( .A(B[35]), .B(A[35]), .Z(n382) );
  CND2XL U1181 ( .A(B[39]), .B(A[39]), .Z(n344) );
  CND2XL U1182 ( .A(B[43]), .B(A[43]), .Z(n302) );
  CND2XL U1183 ( .A(B[3]), .B(A[3]), .Z(n643) );
  CND2XL U1184 ( .A(B[25]), .B(A[25]), .Z(n482) );
  CND2XL U1185 ( .A(B[19]), .B(A[19]), .Z(n540) );
  CND2XL U1186 ( .A(B[27]), .B(A[27]), .Z(n460) );
  CND2XL U1187 ( .A(B[15]), .B(A[15]), .Z(n571) );
  CND2XL U1188 ( .A(B[7]), .B(A[7]), .Z(n624) );
  CND2XL U1189 ( .A(B[31]), .B(A[31]), .Z(n414) );
  CND2XL U1190 ( .A(B[13]), .B(A[13]), .Z(n585) );
  CND2XL U1191 ( .A(B[29]), .B(A[29]), .Z(n438) );
  CND2XL U1192 ( .A(B[5]), .B(A[5]), .Z(n632) );
  CND2XL U1193 ( .A(B[37]), .B(A[37]), .Z(n362) );
  CND2XL U1194 ( .A(B[21]), .B(A[21]), .Z(n520) );
  CND2XL U1195 ( .A(B[49]), .B(A[49]), .Z(n236) );
  CND2XL U1196 ( .A(B[51]), .B(A[51]), .Z(n214) );
  CND2XL U1197 ( .A(B[55]), .B(A[55]), .Z(n168) );
  CND2XL U1198 ( .A(B[57]), .B(A[57]), .Z(n146) );
  CND2XL U1199 ( .A(B[53]), .B(A[53]), .Z(n192) );
  CND2XL U1200 ( .A(B[59]), .B(A[59]), .Z(n122) );
  CND2XL U1201 ( .A(B[61]), .B(A[61]), .Z(n98) );
  CND2X1 U1202 ( .A(B[63]), .B(A[63]), .Z(n72) );
  CND2X1 U1203 ( .A(n916), .B(n72), .Z(n7) );
  CANR1XL U1204 ( .A(n74), .B(n917), .C(n75), .Z(n73) );
  CND2XL U1205 ( .A(n915), .B(n85), .Z(n8) );
  CANR1XL U1206 ( .A(n87), .B(n917), .C(n88), .Z(n86) );
  CND2XL U1207 ( .A(n655), .B(n98), .Z(n9) );
  CANR1XL U1208 ( .A(n100), .B(n917), .C(n101), .Z(n99) );
  CND2XL U1209 ( .A(n656), .B(n109), .Z(n10) );
  CANR1XL U1210 ( .A(n111), .B(n917), .C(n112), .Z(n110) );
  CND2XL U1211 ( .A(n657), .B(n122), .Z(n11) );
  CANR1XL U1212 ( .A(n124), .B(n917), .C(n125), .Z(n123) );
  CND2XL U1213 ( .A(n658), .B(n133), .Z(n12) );
  CANR1XL U1214 ( .A(n135), .B(n917), .C(n136), .Z(n134) );
  CND2XL U1215 ( .A(n659), .B(n146), .Z(n13) );
  CANR1XL U1216 ( .A(n148), .B(n917), .C(n149), .Z(n147) );
  CND2XL U1217 ( .A(n660), .B(n155), .Z(n14) );
  CANR1XL U1218 ( .A(n157), .B(n917), .C(n158), .Z(n156) );
  CND2XL U1219 ( .A(n661), .B(n168), .Z(n15) );
  CANR1XL U1220 ( .A(n170), .B(n917), .C(n171), .Z(n169) );
  CND2XL U1221 ( .A(n662), .B(n179), .Z(n16) );
  CANR1XL U1222 ( .A(n181), .B(n917), .C(n182), .Z(n180) );
  CND2XL U1223 ( .A(n663), .B(n192), .Z(n17) );
  CANR1XL U1224 ( .A(n194), .B(n917), .C(n195), .Z(n193) );
  CND2XL U1225 ( .A(n664), .B(n201), .Z(n18) );
  CANR1XL U1226 ( .A(n203), .B(n917), .C(n204), .Z(n202) );
  CND2XL U1227 ( .A(n665), .B(n214), .Z(n19) );
  CANR1XL U1228 ( .A(n216), .B(n917), .C(n217), .Z(n215) );
  CND2XL U1229 ( .A(n666), .B(n223), .Z(n20) );
  CANR1XL U1230 ( .A(n225), .B(n917), .C(n226), .Z(n224) );
  CND2XL U1231 ( .A(n667), .B(n236), .Z(n21) );
  CANR1XL U1232 ( .A(n238), .B(n917), .C(n239), .Z(n237) );
  CND2XL U1233 ( .A(n668), .B(n243), .Z(n22) );
  CANR1XL U1234 ( .A(n245), .B(n917), .C(n246), .Z(n244) );
  CND2XL U1235 ( .A(n669), .B(n256), .Z(n23) );
  CANR1XL U1236 ( .A(n258), .B(n917), .C(n259), .Z(n257) );
  CND2XL U1237 ( .A(n670), .B(n267), .Z(n24) );
  CANR1XL U1238 ( .A(n269), .B(n917), .C(n270), .Z(n268) );
  CND2XL U1239 ( .A(n671), .B(n280), .Z(n25) );
  CANR1XL U1240 ( .A(n282), .B(n917), .C(n283), .Z(n281) );
  CND2XL U1241 ( .A(n672), .B(n289), .Z(n26) );
  CANR1XL U1242 ( .A(n291), .B(n917), .C(n292), .Z(n290) );
  CND2XL U1243 ( .A(n673), .B(n302), .Z(n27) );
  CANR1XL U1244 ( .A(n304), .B(n917), .C(n305), .Z(n303) );
  CND2XL U1245 ( .A(n674), .B(n311), .Z(n28) );
  CANR1XL U1246 ( .A(n313), .B(n917), .C(n314), .Z(n312) );
  CND2XL U1247 ( .A(n675), .B(n324), .Z(n29) );
  CANR1XL U1248 ( .A(n326), .B(n917), .C(n327), .Z(n325) );
  CND2XL U1249 ( .A(n676), .B(n331), .Z(n30) );
  CANR1XL U1250 ( .A(n333), .B(n917), .C(n334), .Z(n332) );
  CND2XL U1251 ( .A(n677), .B(n344), .Z(n31) );
  CANR1XL U1252 ( .A(n346), .B(n917), .C(n347), .Z(n345) );
  CND2XL U1253 ( .A(n678), .B(n351), .Z(n32) );
  CANR1XL U1254 ( .A(n353), .B(n917), .C(n354), .Z(n352) );
  CND2XL U1255 ( .A(n679), .B(n362), .Z(n33) );
  CANR1XL U1256 ( .A(n364), .B(n917), .C(n365), .Z(n363) );
  CND2XL U1257 ( .A(n680), .B(n369), .Z(n34) );
  CANR1XL U1258 ( .A(n375), .B(n917), .C(n376), .Z(n370) );
  CND2XL U1259 ( .A(n681), .B(n382), .Z(n35) );
  CANR1XL U1260 ( .A(n384), .B(n917), .C(n385), .Z(n383) );
  CND2XL U1261 ( .A(n682), .B(n389), .Z(n36) );
  CANR1XL U1262 ( .A(n391), .B(n917), .C(n392), .Z(n390) );
  CND2XL U1263 ( .A(n683), .B(n398), .Z(n37) );
  CANR1XL U1264 ( .A(n684), .B(n917), .C(n401), .Z(n399) );
  CEOXL U1265 ( .A(n62), .B(n617), .Z(SUM[8]) );
  CND2XL U1266 ( .A(n708), .B(n616), .Z(n62) );
  CND2XL U1267 ( .A(n710), .B(n627), .Z(n64) );
  CEOX1 U1268 ( .A(n65), .B(n633), .Z(SUM[5]) );
  CND2XL U1269 ( .A(n711), .B(n632), .Z(n65) );
  CANR1XL U1270 ( .A(n712), .B(n638), .C(n635), .Z(n633) );
  CENX1 U1271 ( .A(n644), .B(n67), .Z(SUM[3]) );
  CND2XL U1272 ( .A(n713), .B(n643), .Z(n67) );
  COND1XL U1273 ( .A(n645), .B(n647), .C(n646), .Z(n644) );
  CND2XL U1274 ( .A(n701), .B(n571), .Z(n55) );
  CANR1XL U1275 ( .A(n702), .B(n577), .C(n574), .Z(n572) );
  CND2XL U1276 ( .A(n703), .B(n585), .Z(n57) );
  CANR1XL U1277 ( .A(n704), .B(n591), .C(n588), .Z(n586) );
  CND2XL U1278 ( .A(n705), .B(n601), .Z(n59) );
  CANR1XL U1279 ( .A(n706), .B(n607), .C(n604), .Z(n602) );
  CENX1 U1280 ( .A(n917), .B(n38), .Z(SUM[32]) );
  CND2XL U1281 ( .A(n684), .B(n403), .Z(n38) );
  CND2XL U1282 ( .A(n685), .B(n414), .Z(n39) );
  CANR1XL U1283 ( .A(n416), .B(n562), .C(n417), .Z(n415) );
  CND2XL U1284 ( .A(n686), .B(n425), .Z(n40) );
  CANR1XL U1285 ( .A(n427), .B(n562), .C(n428), .Z(n426) );
  CND2XL U1286 ( .A(n687), .B(n438), .Z(n41) );
  CANR1XL U1287 ( .A(n440), .B(n562), .C(n441), .Z(n439) );
  CND2XL U1288 ( .A(n688), .B(n447), .Z(n42) );
  CANR1XL U1289 ( .A(n449), .B(n562), .C(n450), .Z(n448) );
  CND2XL U1290 ( .A(n689), .B(n460), .Z(n43) );
  CANR1XL U1291 ( .A(n462), .B(n562), .C(n463), .Z(n461) );
  CND2XL U1292 ( .A(n690), .B(n469), .Z(n44) );
  CANR1XL U1293 ( .A(n471), .B(n562), .C(n472), .Z(n470) );
  CND2XL U1294 ( .A(n691), .B(n482), .Z(n45) );
  CANR1XL U1295 ( .A(n484), .B(n562), .C(n485), .Z(n483) );
  CND2XL U1296 ( .A(n692), .B(n489), .Z(n46) );
  CANR1XL U1297 ( .A(n491), .B(n562), .C(n492), .Z(n490) );
  CND2XL U1298 ( .A(n693), .B(n502), .Z(n47) );
  CANR1XL U1299 ( .A(n504), .B(n562), .C(n505), .Z(n503) );
  CND2XL U1300 ( .A(n694), .B(n509), .Z(n48) );
  CANR1XL U1301 ( .A(n511), .B(n562), .C(n512), .Z(n510) );
  CND2XL U1302 ( .A(n695), .B(n520), .Z(n49) );
  CANR1XL U1303 ( .A(n522), .B(n562), .C(n523), .Z(n521) );
  CND2XL U1304 ( .A(n696), .B(n527), .Z(n50) );
  CANR1XL U1305 ( .A(n533), .B(n562), .C(n534), .Z(n528) );
  CND2XL U1306 ( .A(n697), .B(n540), .Z(n51) );
  CANR1XL U1307 ( .A(n542), .B(n562), .C(n543), .Z(n541) );
  CND2XL U1308 ( .A(n698), .B(n547), .Z(n52) );
  CANR1XL U1309 ( .A(n549), .B(n562), .C(n550), .Z(n548) );
  CND2XL U1310 ( .A(n699), .B(n556), .Z(n53) );
  CANR1XL U1311 ( .A(n700), .B(n562), .C(n559), .Z(n557) );
  CENX1 U1312 ( .A(n562), .B(n54), .Z(SUM[16]) );
  CND2XL U1313 ( .A(n700), .B(n561), .Z(n54) );
  CENX1 U1314 ( .A(n577), .B(n56), .Z(SUM[14]) );
  CND2XL U1315 ( .A(n702), .B(n576), .Z(n56) );
  CENX1 U1316 ( .A(n591), .B(n58), .Z(SUM[12]) );
  CND2XL U1317 ( .A(n704), .B(n590), .Z(n58) );
  CENX1 U1318 ( .A(n607), .B(n60), .Z(SUM[10]) );
  CND2XL U1319 ( .A(n706), .B(n606), .Z(n60) );
  CENX1 U1320 ( .A(n625), .B(n63), .Z(SUM[7]) );
  CND2XL U1321 ( .A(n709), .B(n624), .Z(n63) );
  COND1XL U1322 ( .A(n626), .B(n628), .C(n627), .Z(n625) );
  CENX1 U1323 ( .A(n614), .B(n61), .Z(SUM[9]) );
  CND2XL U1324 ( .A(n707), .B(n613), .Z(n61) );
  COND1XL U1325 ( .A(n615), .B(n617), .C(n616), .Z(n614) );
  CENX1 U1326 ( .A(n638), .B(n66), .Z(SUM[4]) );
  CND2XL U1327 ( .A(n712), .B(n637), .Z(n66) );
  CEOX1 U1328 ( .A(n68), .B(n647), .Z(SUM[2]) );
  CND2XL U1329 ( .A(n714), .B(n646), .Z(n68) );
  CEOXL U1330 ( .A(n652), .B(n69), .Z(SUM[1]) );
  CND2XL U1331 ( .A(n715), .B(n650), .Z(n69) );
  CANR1X2 U1332 ( .A(n334), .B(n249), .C(n250), .Z(n3) );
  CIVX2 U1333 ( .A(n96), .Z(n94) );
  CIVX2 U1334 ( .A(n95), .Z(n93) );
  CIVX2 U1335 ( .A(n85), .Z(n83) );
  CIVX2 U1336 ( .A(n649), .Z(n715) );
  CIVX2 U1337 ( .A(n645), .Z(n714) );
  CIVX2 U1338 ( .A(n642), .Z(n713) );
  CIVX2 U1339 ( .A(n631), .Z(n711) );
  CIVX2 U1340 ( .A(n626), .Z(n710) );
  CIVX2 U1341 ( .A(n623), .Z(n709) );
  CIVX2 U1342 ( .A(n615), .Z(n708) );
  CIVX2 U1343 ( .A(n612), .Z(n707) );
  CIVX2 U1344 ( .A(n600), .Z(n705) );
  CIVX2 U1345 ( .A(n584), .Z(n703) );
  CIVX2 U1346 ( .A(n570), .Z(n701) );
  CIVX2 U1347 ( .A(n555), .Z(n699) );
  CIVX2 U1348 ( .A(n544), .Z(n698) );
  CIVX2 U1349 ( .A(n539), .Z(n697) );
  CIVX2 U1350 ( .A(n524), .Z(n696) );
  CIVX2 U1351 ( .A(n519), .Z(n695) );
  CIVX2 U1352 ( .A(n506), .Z(n694) );
  CIVX2 U1353 ( .A(n501), .Z(n693) );
  CIVX2 U1354 ( .A(n486), .Z(n692) );
  CIVX2 U1355 ( .A(n481), .Z(n691) );
  CIVX2 U1356 ( .A(n459), .Z(n689) );
  CIVX2 U1357 ( .A(n437), .Z(n687) );
  CIVX2 U1358 ( .A(n422), .Z(n686) );
  CIVX2 U1359 ( .A(n413), .Z(n685) );
  CIVX2 U1360 ( .A(n397), .Z(n683) );
  CIVX2 U1361 ( .A(n386), .Z(n682) );
  CIVX2 U1362 ( .A(n381), .Z(n681) );
  CIVX2 U1363 ( .A(n366), .Z(n680) );
  CIVX2 U1364 ( .A(n361), .Z(n679) );
  CIVX2 U1365 ( .A(n348), .Z(n678) );
  CIVX2 U1366 ( .A(n343), .Z(n677) );
  CIVX2 U1367 ( .A(n328), .Z(n676) );
  CIVX2 U1368 ( .A(n323), .Z(n675) );
  CIVX2 U1369 ( .A(n301), .Z(n673) );
  CIVX2 U1370 ( .A(n279), .Z(n671) );
  CIVX2 U1371 ( .A(n264), .Z(n670) );
  CIVX2 U1372 ( .A(n255), .Z(n669) );
  CIVX2 U1373 ( .A(n240), .Z(n668) );
  CIVX2 U1374 ( .A(n235), .Z(n667) );
  CIVX2 U1375 ( .A(n213), .Z(n665) );
  CIVX2 U1376 ( .A(n191), .Z(n663) );
  CIVX2 U1377 ( .A(n176), .Z(n662) );
  CIVX2 U1378 ( .A(n167), .Z(n661) );
  CIVX2 U1379 ( .A(n145), .Z(n659) );
  CIVX2 U1380 ( .A(n130), .Z(n658) );
  CIVX2 U1381 ( .A(n121), .Z(n657) );
  CIVX2 U1382 ( .A(n106), .Z(n656) );
  CIVX2 U1383 ( .A(n97), .Z(n655) );
  CIVX2 U1384 ( .A(n648), .Z(n647) );
  CIVX2 U1385 ( .A(n639), .Z(n638) );
  CIVX2 U1386 ( .A(n637), .Z(n635) );
  CIVX2 U1387 ( .A(n636), .Z(n712) );
  CIVX2 U1388 ( .A(n618), .Z(n617) );
  CIVX2 U1389 ( .A(n611), .Z(n609) );
  CIVX2 U1390 ( .A(n610), .Z(n608) );
  CIVX2 U1391 ( .A(n606), .Z(n604) );
  CIVX2 U1392 ( .A(n605), .Z(n706) );
  CIVX2 U1393 ( .A(n593), .Z(n595) );
  CIVX2 U1394 ( .A(n592), .Z(n594) );
  CIVX2 U1395 ( .A(n590), .Z(n588) );
  CIVX2 U1396 ( .A(n589), .Z(n704) );
  CIVX2 U1397 ( .A(n576), .Z(n574) );
  CIVX2 U1398 ( .A(n575), .Z(n702) );
  CIVX2 U1399 ( .A(n561), .Z(n559) );
  CIVX2 U1400 ( .A(n560), .Z(n700) );
  CIVX2 U1401 ( .A(n550), .Z(n552) );
  CIVX2 U1402 ( .A(n532), .Z(n534) );
  CIVX2 U1403 ( .A(n531), .Z(n533) );
  CIVX2 U1404 ( .A(n514), .Z(n512) );
  CIVX2 U1405 ( .A(n513), .Z(n511) );
  CIVX2 U1406 ( .A(n492), .Z(n494) );
  CIVX2 U1407 ( .A(n491), .Z(n493) );
  CIVX2 U1408 ( .A(n476), .Z(n474) );
  CIVX2 U1409 ( .A(n475), .Z(n473) );
  CIVX2 U1410 ( .A(n469), .Z(n467) );
  CIVX2 U1411 ( .A(n468), .Z(n690) );
  CIVX2 U1412 ( .A(n452), .Z(n454) );
  CIVX2 U1413 ( .A(n451), .Z(n453) );
  CIVX2 U1414 ( .A(n447), .Z(n445) );
  CIVX2 U1415 ( .A(n446), .Z(n688) );
  CIVX2 U1416 ( .A(n432), .Z(n434) );
  CIVX2 U1417 ( .A(n403), .Z(n401) );
  CIVX2 U1418 ( .A(n402), .Z(n684) );
  CIVX2 U1419 ( .A(n392), .Z(n394) );
  CIVX2 U1420 ( .A(n374), .Z(n376) );
  CIVX2 U1421 ( .A(n373), .Z(n375) );
  CIVX2 U1422 ( .A(n356), .Z(n354) );
  CIVX2 U1423 ( .A(n355), .Z(n353) );
  CIVX2 U1424 ( .A(n334), .Z(n336) );
  CIVX2 U1425 ( .A(n333), .Z(n335) );
  CIVX2 U1426 ( .A(n318), .Z(n316) );
  CIVX2 U1427 ( .A(n317), .Z(n315) );
  CIVX2 U1428 ( .A(n311), .Z(n309) );
  CIVX2 U1429 ( .A(n310), .Z(n674) );
  CIVX2 U1430 ( .A(n294), .Z(n296) );
  CIVX2 U1431 ( .A(n293), .Z(n295) );
  CIVX2 U1432 ( .A(n289), .Z(n287) );
  CIVX2 U1433 ( .A(n288), .Z(n672) );
  CIVX2 U1434 ( .A(n274), .Z(n276) );
  CIVX2 U1435 ( .A(n3), .Z(n246) );
  CIVX2 U1436 ( .A(n4), .Z(n245) );
  CIVX2 U1437 ( .A(n230), .Z(n228) );
  CIVX2 U1438 ( .A(n229), .Z(n227) );
  CIVX2 U1439 ( .A(n223), .Z(n221) );
  CIVX2 U1440 ( .A(n222), .Z(n666) );
  CIVX2 U1441 ( .A(n206), .Z(n208) );
  CIVX2 U1442 ( .A(n205), .Z(n207) );
  CIVX2 U1443 ( .A(n201), .Z(n199) );
  CIVX2 U1444 ( .A(n200), .Z(n664) );
  CIVX2 U1445 ( .A(n186), .Z(n188) );
  CIVX2 U1446 ( .A(n5), .Z(n160) );
  CIVX2 U1447 ( .A(n6), .Z(n159) );
  CIVX2 U1448 ( .A(n155), .Z(n153) );
  CIVX2 U1449 ( .A(n154), .Z(n660) );
  CIVX2 U1450 ( .A(n140), .Z(n142) );
  CIVX2 U1451 ( .A(n118), .Z(n116) );
  CIVX2 U1452 ( .A(n117), .Z(n115) );
  CIVX2 U1453 ( .A(n70), .Z(SUM[0]) );
endmodule


module sfilt_DW01_add_3 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31, n32,
         n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n68, n69, n70, n71, n72, n73, n74, n75, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n216, n217, n218, n219, n220, n221, n222,
         n223, n225, n226, n227, n228, n229, n230, n231, n232, n233, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n260, n261, n262, n263, n264, n265, n266, n267, n269, n270,
         n271;
  assign n13 = A[56];
  assign n17 = A[55];
  assign n24 = A[54];
  assign n28 = A[53];
  assign n33 = A[52];
  assign n37 = A[51];
  assign n43 = A[50];
  assign n47 = A[49];
  assign n52 = A[48];
  assign n56 = A[47];
  assign n64 = A[46];
  assign n68 = A[45];
  assign n73 = A[44];
  assign n77 = A[43];
  assign n83 = A[42];
  assign n87 = A[41];
  assign n92 = A[40];
  assign n96 = A[39];
  assign n104 = A[38];
  assign n108 = A[37];
  assign n113 = A[36];
  assign n117 = A[35];
  assign n123 = A[34];
  assign n127 = A[33];
  assign n132 = A[32];
  assign n135 = A[31];
  assign n143 = A[30];
  assign n146 = A[29];
  assign n150 = A[28];
  assign n153 = A[27];
  assign n160 = A[26];
  assign n163 = A[25];
  assign n167 = A[24];
  assign n170 = A[23];
  assign n177 = A[22];
  assign n180 = A[21];
  assign n184 = A[20];
  assign n187 = A[19];
  assign n194 = A[18];
  assign n197 = A[17];
  assign n201 = A[16];
  assign n205 = A[15];
  assign n212 = A[14];
  assign n216 = A[13];
  assign n221 = A[12];
  assign n225 = A[11];
  assign n231 = A[10];
  assign n235 = A[9];
  assign n240 = A[8];
  assign n243 = A[7];
  assign n249 = A[6];
  assign n252 = A[5];
  assign n256 = A[4];
  assign n260 = A[3];
  assign n265 = A[2];
  assign n269 = A[1];

  CHA1X1 U2 ( .A(A[62]), .B(n4), .CO(n3), .S(SUM[62]) );
  CHA1X1 U3 ( .A(A[61]), .B(n5), .CO(n4), .S(SUM[61]) );
  CHA1X1 U4 ( .A(A[60]), .B(n6), .CO(n5), .S(SUM[60]) );
  CHA1X1 U5 ( .A(A[59]), .B(n7), .CO(n6), .S(SUM[59]) );
  CHA1X1 U6 ( .A(A[58]), .B(n8), .CO(n7), .S(SUM[58]) );
  CHA1X1 U7 ( .A(A[57]), .B(n9), .CO(n8), .S(SUM[57]) );
  CIVXL U334 ( .A(n138), .Z(n137) );
  CIVX1 U335 ( .A(n208), .Z(n207) );
  CIVXL U336 ( .A(n246), .Z(n245) );
  CIVX1 U337 ( .A(n263), .Z(n262) );
  CNR2XL U338 ( .A(n1), .B(n270), .Z(n267) );
  CEOXL U339 ( .A(n1), .B(n270), .Z(SUM[1]) );
  CNR2XL U340 ( .A(A[0]), .B(B[0]), .Z(n271) );
  CNR2X1 U341 ( .A(n155), .B(n149), .Z(n148) );
  CNR2X1 U342 ( .A(n172), .B(n166), .Z(n165) );
  CNR2X1 U343 ( .A(n189), .B(n183), .Z(n182) );
  CNR2X1 U344 ( .A(n19), .B(n18), .Z(n15) );
  CNR2X1 U345 ( .A(n30), .B(n29), .Z(n26) );
  CNR2X1 U346 ( .A(n40), .B(n38), .Z(n35) );
  CNR2X1 U347 ( .A(n49), .B(n48), .Z(n45) );
  CNR2X1 U348 ( .A(n70), .B(n69), .Z(n66) );
  CNR2X1 U349 ( .A(n80), .B(n78), .Z(n75) );
  CNR2X1 U350 ( .A(n89), .B(n88), .Z(n85) );
  CNR2X1 U351 ( .A(n110), .B(n109), .Z(n106) );
  CNR2X1 U352 ( .A(n129), .B(n128), .Z(n125) );
  CNR2X1 U353 ( .A(n172), .B(n157), .Z(n156) );
  CNR2X1 U354 ( .A(n207), .B(n174), .Z(n173) );
  CNR2X1 U355 ( .A(n207), .B(n191), .Z(n190) );
  CND2X1 U356 ( .A(n58), .B(n20), .Z(n19) );
  CND2X1 U357 ( .A(n39), .B(n31), .Z(n30) );
  CND2X1 U358 ( .A(n58), .B(n50), .Z(n49) );
  CND2X1 U359 ( .A(n79), .B(n71), .Z(n70) );
  CND2X1 U360 ( .A(n98), .B(n90), .Z(n89) );
  CND2X1 U361 ( .A(n119), .B(n111), .Z(n110) );
  CND2X1 U362 ( .A(n137), .B(n130), .Z(n129) );
  CND2X1 U363 ( .A(n139), .B(n208), .Z(n138) );
  CNR2X1 U364 ( .A(n174), .B(n140), .Z(n139) );
  CND2X1 U365 ( .A(n158), .B(n141), .Z(n140) );
  CNR2X1 U366 ( .A(n149), .B(n142), .Z(n141) );
  CND2X1 U367 ( .A(n58), .B(n41), .Z(n40) );
  CND2X1 U368 ( .A(n137), .B(n60), .Z(n59) );
  CND2X1 U369 ( .A(n98), .B(n81), .Z(n80) );
  CND2X1 U370 ( .A(n137), .B(n100), .Z(n99) );
  CND2X1 U371 ( .A(n137), .B(n121), .Z(n120) );
  CNR2X1 U372 ( .A(n207), .B(n200), .Z(n199) );
  CNR2X1 U373 ( .A(n262), .B(n255), .Z(n254) );
  CNR2X1 U374 ( .A(n59), .B(n57), .Z(n54) );
  CNR2X1 U375 ( .A(n99), .B(n97), .Z(n94) );
  CNR2X1 U376 ( .A(n120), .B(n118), .Z(n115) );
  CNR2X1 U377 ( .A(n207), .B(n206), .Z(n203) );
  CNR2X1 U378 ( .A(n218), .B(n217), .Z(n214) );
  CNR2X1 U379 ( .A(n228), .B(n226), .Z(n223) );
  CNR2X1 U380 ( .A(n237), .B(n236), .Z(n233) );
  CNR2X1 U381 ( .A(n262), .B(n261), .Z(n258) );
  CND2X1 U382 ( .A(n227), .B(n219), .Z(n218) );
  CND2X1 U383 ( .A(n245), .B(n238), .Z(n237) );
  CND2X1 U384 ( .A(n245), .B(n229), .Z(n228) );
  CENX1 U385 ( .A(n15), .B(n14), .Z(SUM[56]) );
  CEOX1 U386 ( .A(n18), .B(n19), .Z(SUM[55]) );
  CENX1 U387 ( .A(n26), .B(n25), .Z(SUM[54]) );
  CEOX1 U388 ( .A(n29), .B(n30), .Z(SUM[53]) );
  CENX1 U389 ( .A(n35), .B(n34), .Z(SUM[52]) );
  CENX1 U390 ( .A(n39), .B(n38), .Z(SUM[51]) );
  CENX1 U391 ( .A(n45), .B(n44), .Z(SUM[50]) );
  CEOX1 U392 ( .A(n48), .B(n49), .Z(SUM[49]) );
  CENX1 U393 ( .A(n58), .B(n57), .Z(SUM[47]) );
  CENX1 U394 ( .A(n66), .B(n65), .Z(SUM[46]) );
  CEOX1 U395 ( .A(n69), .B(n70), .Z(SUM[45]) );
  CENX1 U396 ( .A(n75), .B(n74), .Z(SUM[44]) );
  CENX1 U397 ( .A(n79), .B(n78), .Z(SUM[43]) );
  CENX1 U398 ( .A(n85), .B(n84), .Z(SUM[42]) );
  CEOX1 U399 ( .A(n88), .B(n89), .Z(SUM[41]) );
  CENX1 U400 ( .A(n106), .B(n105), .Z(SUM[38]) );
  CEOX1 U401 ( .A(n109), .B(n110), .Z(SUM[37]) );
  CENX1 U402 ( .A(n125), .B(n124), .Z(SUM[34]) );
  CEOX1 U403 ( .A(n144), .B(n145), .Z(SUM[30]) );
  CENX1 U404 ( .A(n148), .B(n147), .Z(SUM[29]) );
  CEOX1 U405 ( .A(n151), .B(n152), .Z(SUM[28]) );
  CEOX1 U406 ( .A(n154), .B(n155), .Z(SUM[27]) );
  CEOX1 U407 ( .A(n161), .B(n162), .Z(SUM[26]) );
  CENX1 U408 ( .A(n165), .B(n164), .Z(SUM[25]) );
  CEOX1 U409 ( .A(n178), .B(n179), .Z(SUM[22]) );
  CENX1 U410 ( .A(n182), .B(n181), .Z(SUM[21]) );
  CND2X1 U411 ( .A(A[0]), .B(B[0]), .Z(n1) );
  CNR2X1 U412 ( .A(n239), .B(n230), .Z(n229) );
  CND2X1 U413 ( .A(n235), .B(n231), .Z(n230) );
  CNR2X1 U414 ( .A(n131), .B(n122), .Z(n121) );
  CND2X1 U415 ( .A(n127), .B(n123), .Z(n122) );
  CNR2X1 U416 ( .A(n91), .B(n82), .Z(n81) );
  CND2X1 U417 ( .A(n87), .B(n83), .Z(n82) );
  CNR2X1 U418 ( .A(n51), .B(n42), .Z(n41) );
  CND2X1 U419 ( .A(n47), .B(n43), .Z(n42) );
  CNR2X1 U420 ( .A(n101), .B(n61), .Z(n60) );
  CND2X1 U421 ( .A(n81), .B(n62), .Z(n61) );
  CNR2X1 U422 ( .A(n72), .B(n63), .Z(n62) );
  CND2X1 U423 ( .A(n68), .B(n64), .Z(n63) );
  CNR2X1 U424 ( .A(n264), .B(n1), .Z(n263) );
  CND2X1 U425 ( .A(n269), .B(n265), .Z(n264) );
  CNR2X1 U426 ( .A(n209), .B(n246), .Z(n208) );
  CND2X1 U427 ( .A(n229), .B(n210), .Z(n209) );
  CNR2X1 U428 ( .A(n220), .B(n211), .Z(n210) );
  CND2X1 U429 ( .A(n216), .B(n212), .Z(n211) );
  CNR2X1 U430 ( .A(n166), .B(n159), .Z(n158) );
  CND2X1 U431 ( .A(n163), .B(n160), .Z(n159) );
  CNR2X1 U432 ( .A(n10), .B(n138), .Z(n9) );
  CND2X1 U433 ( .A(n60), .B(n11), .Z(n10) );
  CNR2X1 U434 ( .A(n21), .B(n12), .Z(n11) );
  CND2X1 U435 ( .A(n260), .B(n256), .Z(n255) );
  CND2X1 U436 ( .A(n205), .B(n201), .Z(n200) );
  CND2X1 U437 ( .A(n187), .B(n184), .Z(n183) );
  CND2X1 U438 ( .A(n170), .B(n167), .Z(n166) );
  CND2X1 U439 ( .A(n153), .B(n150), .Z(n149) );
  CND2X1 U440 ( .A(n192), .B(n175), .Z(n174) );
  CNR2X1 U441 ( .A(n183), .B(n176), .Z(n175) );
  CND2X1 U442 ( .A(n180), .B(n177), .Z(n176) );
  CND2X1 U443 ( .A(n247), .B(n263), .Z(n246) );
  CNR2X1 U444 ( .A(n255), .B(n248), .Z(n247) );
  CND2X1 U445 ( .A(n252), .B(n249), .Z(n248) );
  CND2X1 U446 ( .A(n243), .B(n240), .Z(n239) );
  CND2X1 U447 ( .A(n225), .B(n221), .Z(n220) );
  CND2X1 U448 ( .A(n135), .B(n132), .Z(n131) );
  CND2X1 U449 ( .A(n117), .B(n113), .Z(n112) );
  CND2X1 U450 ( .A(n96), .B(n92), .Z(n91) );
  CND2X1 U451 ( .A(n77), .B(n73), .Z(n72) );
  CND2X1 U452 ( .A(n56), .B(n52), .Z(n51) );
  CND2X1 U453 ( .A(n37), .B(n33), .Z(n32) );
  CND2X1 U454 ( .A(n121), .B(n102), .Z(n101) );
  CNR2X1 U455 ( .A(n112), .B(n103), .Z(n102) );
  CND2X1 U456 ( .A(n108), .B(n104), .Z(n103) );
  CND2X1 U457 ( .A(n41), .B(n22), .Z(n21) );
  CNR2X1 U458 ( .A(n32), .B(n23), .Z(n22) );
  CND2X1 U459 ( .A(n28), .B(n24), .Z(n23) );
  CND2X1 U460 ( .A(n148), .B(n146), .Z(n145) );
  CND2X1 U461 ( .A(n156), .B(n153), .Z(n152) );
  CND2X1 U462 ( .A(n165), .B(n163), .Z(n162) );
  CND2X1 U463 ( .A(n182), .B(n180), .Z(n179) );
  CEOX1 U464 ( .A(A[63]), .B(n3), .Z(SUM[63]) );
  CND2X1 U465 ( .A(n146), .B(n143), .Z(n142) );
  CNR2X1 U466 ( .A(n200), .B(n193), .Z(n192) );
  CND2X1 U467 ( .A(n197), .B(n194), .Z(n193) );
  CND2X1 U468 ( .A(n17), .B(n13), .Z(n12) );
  CENX1 U469 ( .A(n54), .B(n53), .Z(SUM[48]) );
  CENX1 U470 ( .A(n94), .B(n93), .Z(SUM[40]) );
  CENX1 U471 ( .A(n98), .B(n97), .Z(SUM[39]) );
  CENX1 U472 ( .A(n115), .B(n114), .Z(SUM[36]) );
  CENX1 U473 ( .A(n119), .B(n118), .Z(SUM[35]) );
  CEOX1 U474 ( .A(n128), .B(n129), .Z(SUM[33]) );
  CEOX1 U475 ( .A(n133), .B(n134), .Z(SUM[32]) );
  CENX1 U476 ( .A(n137), .B(n136), .Z(SUM[31]) );
  CEOX1 U477 ( .A(n168), .B(n169), .Z(SUM[24]) );
  CEOX1 U478 ( .A(n171), .B(n172), .Z(SUM[23]) );
  CEOX1 U479 ( .A(n185), .B(n186), .Z(SUM[20]) );
  CEOX1 U480 ( .A(n188), .B(n189), .Z(SUM[19]) );
  CEOX1 U481 ( .A(n195), .B(n196), .Z(SUM[18]) );
  CENX1 U482 ( .A(n199), .B(n198), .Z(SUM[17]) );
  CENX1 U483 ( .A(n203), .B(n202), .Z(SUM[16]) );
  CEOX1 U484 ( .A(n206), .B(n207), .Z(SUM[15]) );
  CENX1 U485 ( .A(n214), .B(n213), .Z(SUM[14]) );
  CEOX1 U486 ( .A(n217), .B(n218), .Z(SUM[13]) );
  CENX1 U487 ( .A(n223), .B(n222), .Z(SUM[12]) );
  CENX1 U488 ( .A(n227), .B(n226), .Z(SUM[11]) );
  CENX1 U489 ( .A(n233), .B(n232), .Z(SUM[10]) );
  CEOX1 U490 ( .A(n236), .B(n237), .Z(SUM[9]) );
  CEOX1 U491 ( .A(n241), .B(n242), .Z(SUM[8]) );
  CENX1 U492 ( .A(n245), .B(n244), .Z(SUM[7]) );
  CEOX1 U493 ( .A(n250), .B(n251), .Z(SUM[6]) );
  CENX1 U494 ( .A(n258), .B(n257), .Z(SUM[4]) );
  CENX1 U495 ( .A(n267), .B(n266), .Z(SUM[2]) );
  CENX1 U496 ( .A(n254), .B(n253), .Z(SUM[5]) );
  CND2X1 U497 ( .A(n137), .B(n135), .Z(n134) );
  CND2X1 U498 ( .A(n173), .B(n170), .Z(n169) );
  CND2X1 U499 ( .A(n190), .B(n187), .Z(n186) );
  CND2X1 U500 ( .A(n199), .B(n197), .Z(n196) );
  CND2X1 U501 ( .A(n245), .B(n243), .Z(n242) );
  CND2X1 U502 ( .A(n254), .B(n252), .Z(n251) );
  CEOX1 U503 ( .A(n261), .B(n262), .Z(SUM[3]) );
  CND2IX1 U504 ( .B(n271), .A(n1), .Z(n2) );
  CIVX2 U505 ( .A(n99), .Z(n98) );
  CIVX2 U506 ( .A(n96), .Z(n97) );
  CIVX2 U507 ( .A(n92), .Z(n93) );
  CIVX2 U508 ( .A(n91), .Z(n90) );
  CIVX2 U509 ( .A(n87), .Z(n88) );
  CIVX2 U510 ( .A(n83), .Z(n84) );
  CIVX2 U511 ( .A(n80), .Z(n79) );
  CIVX2 U512 ( .A(n77), .Z(n78) );
  CIVX2 U513 ( .A(n73), .Z(n74) );
  CIVX2 U514 ( .A(n72), .Z(n71) );
  CIVX2 U515 ( .A(n68), .Z(n69) );
  CIVX2 U516 ( .A(n64), .Z(n65) );
  CIVX2 U517 ( .A(n59), .Z(n58) );
  CIVX2 U518 ( .A(n56), .Z(n57) );
  CIVX2 U519 ( .A(n52), .Z(n53) );
  CIVX2 U520 ( .A(n51), .Z(n50) );
  CIVX2 U521 ( .A(n47), .Z(n48) );
  CIVX2 U522 ( .A(n43), .Z(n44) );
  CIVX2 U523 ( .A(n40), .Z(n39) );
  CIVX2 U524 ( .A(n37), .Z(n38) );
  CIVX2 U525 ( .A(n33), .Z(n34) );
  CIVX2 U526 ( .A(n32), .Z(n31) );
  CIVX2 U527 ( .A(n28), .Z(n29) );
  CIVX2 U528 ( .A(n269), .Z(n270) );
  CIVX2 U529 ( .A(n265), .Z(n266) );
  CIVX2 U530 ( .A(n260), .Z(n261) );
  CIVX2 U531 ( .A(n256), .Z(n257) );
  CIVX2 U532 ( .A(n252), .Z(n253) );
  CIVX2 U533 ( .A(n249), .Z(n250) );
  CIVX2 U534 ( .A(n24), .Z(n25) );
  CIVX2 U535 ( .A(n243), .Z(n244) );
  CIVX2 U536 ( .A(n240), .Z(n241) );
  CIVX2 U537 ( .A(n239), .Z(n238) );
  CIVX2 U538 ( .A(n235), .Z(n236) );
  CIVX2 U539 ( .A(n231), .Z(n232) );
  CIVX2 U540 ( .A(n228), .Z(n227) );
  CIVX2 U541 ( .A(n225), .Z(n226) );
  CIVX2 U542 ( .A(n221), .Z(n222) );
  CIVX2 U543 ( .A(n220), .Z(n219) );
  CIVX2 U544 ( .A(n216), .Z(n217) );
  CIVX2 U545 ( .A(n212), .Z(n213) );
  CIVX2 U546 ( .A(n205), .Z(n206) );
  CIVX2 U547 ( .A(n201), .Z(n202) );
  CIVX2 U548 ( .A(n21), .Z(n20) );
  CIVX2 U549 ( .A(n197), .Z(n198) );
  CIVX2 U550 ( .A(n194), .Z(n195) );
  CIVX2 U551 ( .A(n192), .Z(n191) );
  CIVX2 U552 ( .A(n190), .Z(n189) );
  CIVX2 U553 ( .A(n187), .Z(n188) );
  CIVX2 U554 ( .A(n184), .Z(n185) );
  CIVX2 U555 ( .A(n180), .Z(n181) );
  CIVX2 U556 ( .A(n177), .Z(n178) );
  CIVX2 U557 ( .A(n173), .Z(n172) );
  CIVX2 U558 ( .A(n170), .Z(n171) );
  CIVX2 U559 ( .A(n167), .Z(n168) );
  CIVX2 U560 ( .A(n163), .Z(n164) );
  CIVX2 U561 ( .A(n160), .Z(n161) );
  CIVX2 U562 ( .A(n17), .Z(n18) );
  CIVX2 U563 ( .A(n158), .Z(n157) );
  CIVX2 U564 ( .A(n156), .Z(n155) );
  CIVX2 U565 ( .A(n153), .Z(n154) );
  CIVX2 U566 ( .A(n150), .Z(n151) );
  CIVX2 U567 ( .A(n146), .Z(n147) );
  CIVX2 U568 ( .A(n143), .Z(n144) );
  CIVX2 U569 ( .A(n13), .Z(n14) );
  CIVX2 U570 ( .A(n135), .Z(n136) );
  CIVX2 U571 ( .A(n132), .Z(n133) );
  CIVX2 U572 ( .A(n131), .Z(n130) );
  CIVX2 U573 ( .A(n127), .Z(n128) );
  CIVX2 U574 ( .A(n123), .Z(n124) );
  CIVX2 U575 ( .A(n120), .Z(n119) );
  CIVX2 U576 ( .A(n117), .Z(n118) );
  CIVX2 U577 ( .A(n113), .Z(n114) );
  CIVX2 U578 ( .A(n112), .Z(n111) );
  CIVX2 U579 ( .A(n108), .Z(n109) );
  CIVX2 U580 ( .A(n104), .Z(n105) );
  CIVX2 U581 ( .A(n101), .Z(n100) );
  CIVX2 U582 ( .A(n2), .Z(SUM[0]) );
endmodule


module sfilt_DW_mult_tc_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n9, n12, n18, n21, n24, n27, n30, n33, n36, n39, n42, n48,
         n51, n54, n57, n63, n66, n75, n81, n84, n87, n90, n93, n99, n102,
         n105, n108, n111, n117, n120, n126, n129, n132, n135, n136, n144,
         n145, n149, n150, n152, n153, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n173, n174, n175, n176, n178, n179, n184, n185, n187, n188, n190,
         n191, n192, n193, n194, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n213, n214, n216, n218,
         n219, n220, n221, n222, n223, n224, n225, n241, n246, n247, n248,
         n249, n254, n255, n256, n257, n258, n259, n260, n261, n262, n274,
         n279, n280, n281, n282, n283, n286, n287, n289, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n301, n302, n303, n304, n306,
         n308, n309, n310, n314, n315, n316, n317, n318, n319, n320, n323,
         n324, n327, n328, n329, n330, n331, n332, n333, n334, n340, n342,
         n343, n344, n345, n349, n351, n352, n353, n354, n355, n356, n360,
         n361, n362, n363, n364, n365, n366, n369, n370, n371, n372, n373,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n392, n393, n394, n395, n396, n397, n399, n402, n403,
         n404, n405, n406, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n424, n426, n427, n428, n432, n434, n435,
         n438, n439, n440, n441, n444, n445, n448, n449, n450, n451, n452,
         n456, n458, n459, n460, n461, n462, n463, n467, n468, n469, n470,
         n471, n472, n474, n478, n480, n486, n487, n488, n489, n490, n495,
         n496, n497, n498, n501, n506, n507, n508, n510, n511, n513, n516,
         n517, n520, n522, n524, n525, n526, n528, n529, n530, n531, n532,
         n534, n535, n540, n541, n542, n543, n544, n546, n548, n550, n551,
         n552, n553, n554, n555, n559, n560, n561, n564, n567, n568, n569,
         n571, n572, n573, n574, n576, n578, n583, n584, n585, n586, n590,
         n591, n592, n593, n594, n596, n597, n603, n604, n605, n606, n613,
         n618, n619, n620, n621, n622, n623, n624, n626, n627, n628, n629,
         n631, n634, n635, n636, n642, n643, n644, n649, n650, n651, n652,
         n654, n656, n657, n658, n659, n660, n661, n662, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n681, n683, n684, n686, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n704,
         n706, n707, n708, n709, n710, n712, n714, n718, n720, n721, n722,
         n723, n724, n726, n728, n729, n730, n731, n735, n738, n739, n740,
         n741, n744, n745, n746, n747, n748, n749, n751, n753, n754, n756,
         n757, n758, n760, n762, n763, n764, n766, n767, n768, n770, n772,
         n773, n774, n776, n778, n779, n780, n781, n784, n785, n786, n791,
         n793, n794, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1108, n1110, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1136, n1137, n1138, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1164,
         n1165, n1166, n1170, n1171, n1172, n1173, n1176, n1177, n1178, n1179,
         n1180, n1181, n1184, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1199, n1201, n1204, n1206, n1207,
         n1208, n1209, n1214, n1215, n1216, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2812, n2813, n2814,
         n2816, n2818, n2819, n2820, n2821, n2822, n2823, n2825, n2826, n2827,
         net15963, net15979, net15975, net15985, net15993, net16005, net16001,
         net15999, net16019, net16015, net16027, net16023, net16389, net16391,
         net16393, net16399, net16403, net16407, net16539, net16549, net16554,
         net16580, net16593, net16606, net16605, net16617, net16623, net16621,
         net16633, net16639, net16638, net16637, net16645, net16649, net16671,
         net16670, net16676, net16684, net16683, net18090, net18096, net18255,
         net18264, net18274, net18280, net18282, net18408, net18407, net18430,
         net18429, net18455, net18453, net18486, net18485, net18492, net18510,
         net18509, net18520, net18538, net18537, net18546, net18545, net18568,
         net18570, net18572, net18573, net18607, net18613, net18612, net18617,
         net18700, net18703, net18736, net18734, net18745, net18744, net18772,
         net18783, net18811, net18809, net18827, net18832, net18830, net18839,
         net18844, net18843, net18867, net18869, net18868, net18887, net18902,
         net18906, net18944, net18953, net18952, net18951, net18983, net18982,
         net19011, net19026, net19025, net19035, net19034, net19148, net19162,
         net19184, net19200, net19203, net19209, net19208, net19253, net19288,
         net19290, net19319, net19358, net19362, net19382, net19384, net19385,
         net19415, net19414, net19422, net19442, net19448, net19447, net19446,
         net19491, net19522, net19521, net19520, net19526, net19538, net19536,
         net19560, net19619, net19618, net19617, net19689, net19695, net19702,
         net19754, net19753, net19757, net19794, net19793, net19845, net19877,
         net19890, net19927, net19953, net19965, net19977, net19987, net19996,
         net20002, net20005, net20022, net20025, net18491, net16682, net16021,
         net16017, n2543, n2017, net19939, net18901, n521, n514, n646, n637,
         n632, n630, n616, n614, n608, n601, n595, n582, n579, n577, n575,
         n556, n549, n547, net21345, net21418, net21540, net21539, net21556,
         net21555, net21565, net21564, net21572, net21576, net21583, net21601,
         net21614, net22007, net22025, net22026, net19048, net18516, net16675,
         net15989, n2373, n2372, n1111, net18254, n795, n229, n227, n151,
         net22015, net21559, net21373, net21367, net19259, net19232, net19207,
         n2815, n114, n512, n1133, net18270, n253, n244, n242, n236, n233,
         n232, n231, n230, net19762, net19760, n78, net18276, net16579,
         net16578, net16577, net21569, net15959, n2311, n2310, n1971, n1853,
         n1796, n1211, n1210, n1205, net18964, net18962, n2156, n1766, n1213,
         n1212, n1200, n1198, n1185, n1175, n1174, n1167, net19249, net19248,
         net16513, net16512, net16511, n485, n484, n1106, n2187, n1203, n1202,
         net19780, net15965, n2155, n1940, n1765, n1183, n1182, n1169, n1168,
         n1163, n1162, n1139, n1135, n1134, net19300, net19299, net18635,
         net18411, net18380, n505, n499, n491, n482, n1132, net18753, net18752,
         net18751, net18750, net18278, n1109, n1107, n736, n266, n265, n264,
         n154, net19938, net19456, net18412, n515, n494, n483, n481, n479,
         n359, n277, n275, n273, n272, n269, n268, n267, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n57 = a[13];
  assign n66 = a[15];
  assign n75 = a[17];
  assign n84 = a[19];
  assign n93 = a[21];
  assign n102 = a[23];
  assign n111 = a[25];
  assign n120 = a[27];
  assign n129 = a[29];
  assign n136 = a[31];
  assign n145 = b[0];
  assign n2780 = b[31];
  assign n2781 = b[30];
  assign n2782 = b[29];
  assign n2783 = b[28];
  assign n2784 = b[27];
  assign n2785 = b[26];
  assign n2786 = b[25];
  assign n2787 = b[24];
  assign n2788 = b[23];
  assign n2789 = b[22];
  assign n2790 = b[21];
  assign n2791 = b[20];
  assign n2792 = b[19];
  assign n2793 = b[18];
  assign n2794 = b[17];
  assign n2795 = b[16];
  assign n2796 = b[15];
  assign n2797 = b[14];
  assign n2798 = b[13];
  assign n2799 = b[12];
  assign n2800 = b[11];
  assign n2801 = b[10];
  assign n2802 = b[9];
  assign n2803 = b[8];
  assign n2804 = b[7];
  assign n2805 = b[6];
  assign n2806 = b[5];
  assign n2807 = b[4];
  assign n2808 = b[3];
  assign n2809 = b[2];
  assign n2810 = b[1];

  CND2X2 U187 ( .A(n735), .B(net18255), .Z(n241) );
  COND1X1 U208 ( .A(n257), .B(net18429), .C(n258), .Z(n256) );
  CND2X2 U229 ( .A(n283), .B(net18264), .Z(n274) );
  COND1X1 U238 ( .A(n281), .B(net18429), .C(n282), .Z(n280) );
  CNR2X2 U243 ( .A(n333), .B(n287), .Z(n283) );
  COND1X1 U244 ( .A(n287), .B(n334), .C(n3941), .Z(n286) );
  CNR2X2 U247 ( .A(n291), .B(n324), .Z(n289) );
  CND2X2 U249 ( .A(n293), .B(n740), .Z(n291) );
  CANR1X1 U250 ( .A(n314), .B(n293), .C(n294), .Z(n292) );
  CNR2X2 U251 ( .A(n302), .B(n295), .Z(n293) );
  COND1X1 U252 ( .A(n295), .B(n303), .C(n296), .Z(n294) );
  CNR2X2 U255 ( .A(n813), .B(n818), .Z(n295) );
  CNR2X2 U265 ( .A(n826), .B(n819), .Z(n302) );
  CND2X2 U266 ( .A(n826), .B(n819), .Z(n303) );
  COND1X1 U268 ( .A(n3121), .B(net18429), .C(n306), .Z(n304) );
  COND1X1 U284 ( .A(n318), .B(net18430), .C(n319), .Z(n317) );
  CNR2X2 U295 ( .A(n835), .B(n844), .Z(n324) );
  COND1X1 U298 ( .A(n329), .B(net18429), .C(n330), .Z(n328) );
  COND1X1 U328 ( .A(n353), .B(net18430), .C(net18839), .Z(n352) );
  CNR2X2 U339 ( .A(n365), .B(n389), .Z(n363) );
  CND2X2 U341 ( .A(n745), .B(n744), .Z(n365) );
  CNR2X2 U347 ( .A(n878), .B(n867), .Z(n369) );
  COND1X1 U350 ( .A(n372), .B(net18430), .C(n373), .Z(n371) );
  CNR2X2 U375 ( .A(n893), .B(n906), .Z(n389) );
  COND1X1 U378 ( .A(n394), .B(net18430), .C(n395), .Z(n393) );
  CNR2X2 U385 ( .A(n402), .B(n409), .Z(n396) );
  CND2X2 U400 ( .A(n923), .B(n938), .Z(n410) );
  COND1X1 U402 ( .A(n412), .B(net18430), .C(n413), .Z(n411) );
  CNR2X2 U417 ( .A(n939), .B(n956), .Z(n424) );
  COND1X1 U420 ( .A(n427), .B(n149), .C(n428), .Z(n426) );
  COND1X1 U432 ( .A(n440), .B(net18429), .C(net19526), .Z(n435) );
  CNR2X2 U447 ( .A(n975), .B(n994), .Z(n448) );
  COND1X1 U450 ( .A(n451), .B(net18429), .C(n452), .Z(n450) );
  CNR2X2 U473 ( .A(n3803), .B(n1036), .Z(n468) );
  COND1X1 U476 ( .A(n3144), .B(net18429), .C(n3809), .Z(n470) );
  CNR2X2 U555 ( .A(n1187), .B(n1214), .Z(n529) );
  CNR2X2 U565 ( .A(n3911), .B(n543), .Z(n534) );
  CNR2X2 U608 ( .A(n1333), .B(n1360), .Z(n567) );
  COND1X1 U725 ( .A(n668), .B(n651), .C(n652), .Z(n650) );
  CFA1X1 U858 ( .A(n800), .B(n1771), .CI(n1741), .CO(n796), .S(n797) );
  CFA1X1 U859 ( .A(n1772), .B(n804), .CI(n801), .CO(n798), .S(n799) );
  CFA1X1 U861 ( .A(n1803), .B(n805), .CI(n808), .CO(n802), .S(n803) );
  CFA1X1 U862 ( .A(n810), .B(n1773), .CI(n1742), .CO(n804), .S(n805) );
  CFA1X1 U863 ( .A(n816), .B(n814), .CI(n809), .CO(n806), .S(n807) );
  CFA1X1 U864 ( .A(n1743), .B(n811), .CI(n1804), .CO(n808), .S(n809) );
  CFA1X1 U866 ( .A(n817), .B(n815), .CI(n820), .CO(n812), .S(n813) );
  CFA1X1 U867 ( .A(n1744), .B(n822), .CI(n1834), .CO(n814), .S(n815) );
  CFA1X1 U868 ( .A(n824), .B(n1805), .CI(n1774), .CO(n816), .S(n817) );
  CFA1X1 U869 ( .A(n823), .B(n821), .CI(n828), .CO(n818), .S(n819) );
  CFA1X1 U870 ( .A(n825), .B(n830), .CI(n832), .CO(n820), .S(n821) );
  CFA1X1 U873 ( .A(n838), .B(n829), .CI(n836), .CO(n826), .S(n827) );
  CFA1X1 U874 ( .A(n840), .B(n831), .CI(n833), .CO(n828), .S(n829) );
  CFA1X1 U875 ( .A(n1746), .B(n1864), .CI(n1776), .CO(n830), .S(n831) );
  CFA1X1 U876 ( .A(n842), .B(n1836), .CI(n1806), .CO(n832), .S(n833) );
  CFA1X1 U877 ( .A(n839), .B(n837), .CI(n846), .CO(n834), .S(n835) );
  CFA1X1 U878 ( .A(n850), .B(n848), .CI(n841), .CO(n836), .S(n837) );
  CFA1X1 U879 ( .A(n1837), .B(n852), .CI(n843), .CO(n838), .S(n839) );
  CFA1X1 U880 ( .A(n1777), .B(n1865), .CI(n1747), .CO(n840), .S(n841) );
  CFA1X1 U882 ( .A(n849), .B(n847), .CI(n856), .CO(n844), .S(n845) );
  CFA1X1 U883 ( .A(n851), .B(n858), .CI(n853), .CO(n846), .S(n847) );
  CFA1X1 U884 ( .A(n1895), .B(n860), .CI(n862), .CO(n848), .S(n849) );
  CFA1X1 U887 ( .A(n859), .B(n857), .CI(n868), .CO(n854), .S(n855) );
  CFA1X1 U888 ( .A(n861), .B(n870), .CI(n872), .CO(n856), .S(n857) );
  CFA1X1 U889 ( .A(n876), .B(n863), .CI(n874), .CO(n858), .S(n859) );
  CFA1X1 U890 ( .A(n1867), .B(n865), .CI(n1779), .CO(n860), .S(n861) );
  CFA1X1 U893 ( .A(n871), .B(n869), .CI(n880), .CO(n866), .S(n867) );
  CFA1X1 U894 ( .A(n884), .B(n882), .CI(n873), .CO(n868), .S(n869) );
  CFA1X1 U895 ( .A(n886), .B(n877), .CI(n875), .CO(n870), .S(n871) );
  CFA1X1 U896 ( .A(n1780), .B(n888), .CI(n1927), .CO(n872), .S(n873) );
  CFA1X1 U897 ( .A(n1839), .B(n1868), .CI(n1750), .CO(n874), .S(n875) );
  CFA1X1 U900 ( .A(n898), .B(n896), .CI(n885), .CO(n880), .S(n881) );
  CFA1X1 U901 ( .A(n900), .B(n889), .CI(n887), .CO(n882), .S(n883) );
  CFA1X1 U902 ( .A(n891), .B(n902), .CI(n904), .CO(n884), .S(n885) );
  CFA1X1 U904 ( .A(n1810), .B(n1928), .CI(n1781), .CO(n888), .S(n889) );
  CFA1X1 U908 ( .A(n905), .B(n914), .CI(n901), .CO(n896), .S(n897) );
  CFA1X1 U909 ( .A(n918), .B(n903), .CI(n916), .CO(n898), .S(n899) );
  CFA1X1 U910 ( .A(n920), .B(n1958), .CI(n1899), .CO(n900), .S(n901) );
  CFA1X1 U911 ( .A(n1870), .B(n1840), .CI(n1782), .CO(n902), .S(n903) );
  CFA1X1 U912 ( .A(n1752), .B(n1929), .CI(n1811), .CO(n904), .S(n905) );
  CFA1X1 U913 ( .A(n911), .B(n909), .CI(n924), .CO(n906), .S(n907) );
  CFA1X1 U914 ( .A(n928), .B(n926), .CI(n913), .CO(n908), .S(n909) );
  CFA1X1 U915 ( .A(n919), .B(n915), .CI(n930), .CO(n910), .S(n911) );
  CFA1X1 U916 ( .A(n934), .B(n917), .CI(n932), .CO(n912), .S(n913) );
  CFA1X1 U919 ( .A(n1812), .B(n1959), .CI(n1753), .CO(n918), .S(n919) );
  CFA1X1 U921 ( .A(n927), .B(n925), .CI(n940), .CO(n922), .S(n923) );
  CFA1X1 U922 ( .A(n944), .B(n942), .CI(n929), .CO(n924), .S(n925) );
  CFA1X1 U923 ( .A(n937), .B(n931), .CI(n946), .CO(n926), .S(n927) );
  CFA1X1 U924 ( .A(n948), .B(n935), .CI(n933), .CO(n928), .S(n929) );
  CFA1X1 U925 ( .A(n1990), .B(n950), .CI(n952), .CO(n930), .S(n931) );
  CFA1X1 U926 ( .A(n1841), .B(n3120), .CI(n1901), .CO(n932), .S(n933) );
  CFA1X1 U927 ( .A(n1872), .B(n1813), .CI(n1784), .CO(n934), .S(n935) );
  CFA1X1 U928 ( .A(n1754), .B(n1960), .CI(n954), .CO(n936), .S(n937) );
  CFA1X1 U929 ( .A(n943), .B(n941), .CI(n958), .CO(n938), .S(n939) );
  CFA1X1 U930 ( .A(n945), .B(n960), .CI(n962), .CO(n940), .S(n941) );
  CFA1X1 U931 ( .A(n966), .B(n947), .CI(n964), .CO(n942), .S(n943) );
  CFA1X1 U932 ( .A(n951), .B(n949), .CI(n953), .CO(n944), .S(n945) );
  CFA1X1 U933 ( .A(n972), .B(n970), .CI(n968), .CO(n946), .S(n947) );
  CFA1X1 U934 ( .A(n1961), .B(n955), .CI(n1932), .CO(n948), .S(n949) );
  CFA1X1 U935 ( .A(n1785), .B(n1902), .CI(n1814), .CO(n950), .S(n951) );
  CFA1X1 U938 ( .A(n961), .B(n959), .CI(n976), .CO(n956), .S(n957) );
  CFA1X1 U941 ( .A(n971), .B(n984), .CI(n973), .CO(n962), .S(n963) );
  CFA1X1 U943 ( .A(n1962), .B(n990), .CI(n2022), .CO(n966), .S(n967) );
  CFA1X1 U944 ( .A(n1933), .B(n1873), .CI(n1843), .CO(n968), .S(n969) );
  CFA1X1 U945 ( .A(n1903), .B(n1786), .CI(n1815), .CO(n970), .S(n971) );
  CFA1X1 U946 ( .A(n992), .B(n1992), .CI(n1756), .CO(n972), .S(n973) );
  CFA1X1 U948 ( .A(n1000), .B(n998), .CI(n981), .CO(n976), .S(n977) );
  CFA1X1 U950 ( .A(n989), .B(n1004), .CI(n991), .CO(n980), .S(n981) );
  CFA1X1 U951 ( .A(n1008), .B(n987), .CI(n1006), .CO(n982), .S(n983) );
  CFA1X1 U952 ( .A(n993), .B(n1010), .CI(n1012), .CO(n984), .S(n985) );
  CFA1X1 U953 ( .A(n1934), .B(n1904), .CI(n1963), .CO(n986), .S(n987) );
  CFA1X1 U954 ( .A(n1816), .B(n3045), .CI(n1993), .CO(n988), .S(n989) );
  CFA1X1 U957 ( .A(n999), .B(n997), .CI(n1016), .CO(n994), .S(n995) );
  CFA1X1 U959 ( .A(n1022), .B(n1003), .CI(n1005), .CO(n998), .S(n999) );
  CFA1X1 U960 ( .A(n1007), .B(n1024), .CI(n1026), .CO(n1000), .S(n1001) );
  CFA1X1 U962 ( .A(n1032), .B(n1030), .CI(n1028), .CO(n1004), .S(n1005) );
  CFA1X1 U963 ( .A(n1994), .B(n2055), .CI(n1964), .CO(n1006), .S(n1007) );
  CFA1X1 U964 ( .A(n1817), .B(n1935), .CI(n1874), .CO(n1008), .S(n1009) );
  CFA1X1 U966 ( .A(n1034), .B(n2024), .CI(n1758), .CO(n1012), .S(n1013) );
  CFA1X1 U967 ( .A(n1019), .B(n1017), .CI(n1038), .CO(n1014), .S(n1015) );
  CFA1X1 U969 ( .A(n1044), .B(n1023), .CI(n1025), .CO(n1018), .S(n1019) );
  CFA1X1 U971 ( .A(n1033), .B(n1031), .CI(n1029), .CO(n1022), .S(n1023) );
  CFA1X1 U972 ( .A(n1054), .B(n1052), .CI(n1050), .CO(n1024), .S(n1025) );
  CFA1X1 U973 ( .A(n1965), .B(n1056), .CI(n1035), .CO(n1026), .S(n1027) );
  CFA1X1 U974 ( .A(n1936), .B(n1995), .CI(n1818), .CO(n1028), .S(n1029) );
  CFA1X1 U975 ( .A(n1846), .B(n1789), .CI(n2025), .CO(n1030), .S(n1031) );
  CFA1X1 U978 ( .A(n1041), .B(n1039), .CI(n1060), .CO(n1036), .S(n1037) );
  CFA1X1 U980 ( .A(n1047), .B(n1045), .CI(n1066), .CO(n1040), .S(n1041) );
  CFA1X1 U981 ( .A(n1070), .B(n1068), .CI(n1049), .CO(n1042), .S(n1043) );
  CFA1X1 U985 ( .A(n2026), .B(n1996), .CI(n1876), .CO(n1050), .S(n1051) );
  CFA1X1 U986 ( .A(n1906), .B(n1966), .CI(n1847), .CO(n1052), .S(n1053) );
  CFA1X1 U987 ( .A(n1937), .B(n1790), .CI(n1819), .CO(n1054), .S(n1055) );
  CFA1X1 U988 ( .A(n1760), .B(n2057), .CI(n3038), .CO(n1056), .S(n1057) );
  CFA1X1 U992 ( .A(n1094), .B(n1071), .CI(n1092), .CO(n1064), .S(n1065) );
  CFA1X1 U993 ( .A(n1079), .B(n1096), .CI(n1073), .CO(n1066), .S(n1067) );
  CFA1X1 U995 ( .A(n1104), .B(n1100), .CI(n1098), .CO(n1070), .S(n1071) );
  CFA1X1 U998 ( .A(n2027), .B(n2058), .CI(n1877), .CO(n1076), .S(n1077) );
  CFA1X1 U1002 ( .A(n1112), .B(n1110), .CI(n1089), .CO(n1084), .S(n1085) );
  CFA1X1 U1003 ( .A(n1093), .B(n1091), .CI(n1114), .CO(n1086), .S(n1087) );
  CFA1X1 U1007 ( .A(n1122), .B(n1124), .CI(n1126), .CO(n1094), .S(n1095) );
  CFA1X1 U1010 ( .A(n1938), .B(n1878), .CI(n1849), .CO(n1100), .S(n1101) );
  CFA1X1 U1011 ( .A(n1908), .B(n1821), .CI(n1792), .CO(n1102), .S(n1103) );
  CFA1X1 U1012 ( .A(n1762), .B(n2090), .CI(n2059), .CO(n1104), .S(n1105) );
  CFA1X1 U1016 ( .A(n1144), .B(n1142), .CI(n1119), .CO(n1112), .S(n1113) );
  CFA1X1 U1018 ( .A(n1127), .B(n1123), .CI(n1129), .CO(n1116), .S(n1117) );
  CFA1X1 U1021 ( .A(n2029), .B(n1999), .CI(n2060), .CO(n1122), .S(n1123) );
  CFA1X1 U1022 ( .A(n1969), .B(n2091), .CI(n1850), .CO(n1124), .S(n1125) );
  CFA1X1 U1023 ( .A(n1879), .B(n1822), .CI(n1763), .CO(n1126), .S(n1127) );
  CFA1X1 U1024 ( .A(n1909), .B(n1793), .CI(n2122), .CO(n1128), .S(n1129) );
  CFA1X1 U1031 ( .A(n1155), .B(n1149), .CI(n1157), .CO(n1142), .S(n1143) );
  CFA1X1 U1034 ( .A(n2061), .B(n2154), .CI(n2030), .CO(n1148), .S(n1149) );
  CFA1X1 U1035 ( .A(n1880), .B(n1910), .CI(n2000), .CO(n1150), .S(n1151) );
  CFA1X1 U1036 ( .A(n1970), .B(n1184), .CI(n1851), .CO(n1152), .S(n1153) );
  CFA1X1 U1037 ( .A(n1823), .B(n1939), .CI(n1794), .CO(n1154), .S(n1155) );
  CFA1X1 U1038 ( .A(n1764), .B(n2123), .CI(n2092), .CO(n1156), .S(n1157) );
  CFA1X1 U1048 ( .A(n2124), .B(n2031), .CI(n2062), .CO(n1176), .S(n1177) );
  CFA1X1 U1049 ( .A(n1881), .B(n2001), .CI(n1852), .CO(n1178), .S(n1179) );
  CFA1X1 U1050 ( .A(n1911), .B(n1824), .CI(n1795), .CO(n1180), .S(n1181) );
  CFA1X1 U1053 ( .A(n3490), .B(n1216), .CI(n3914), .CO(n1186), .S(n1187) );
  CFA1X1 U1054 ( .A(n1193), .B(n1218), .CI(n1220), .CO(n1188), .S(n1189) );
  CFA1X1 U1056 ( .A(n1201), .B(n1224), .CI(n1199), .CO(n1192), .S(n1193) );
  CFA1X1 U1063 ( .A(n1825), .B(n2063), .CI(n2032), .CO(n1206), .S(n1207) );
  CFA1X1 U1064 ( .A(n2002), .B(n1912), .CI(n1882), .CO(n1208), .S(n1209) );
  CFA1X1 U1067 ( .A(n3048), .B(n3469), .CI(n1246), .CO(n1214), .S(n1215) );
  CFA1X1 U1071 ( .A(n1258), .B(n1231), .CI(n1256), .CO(n1222), .S(n1223) );
  CFA1X1 U1075 ( .A(n1272), .B(n1264), .CI(n1266), .CO(n1230), .S(n1231) );
  CFA1X1 U1076 ( .A(n2033), .B(n1243), .CI(n2064), .CO(n1232), .S(n1233) );
  CFA1X1 U1082 ( .A(n1249), .B(n1247), .CI(n1276), .CO(n1244), .S(n1245) );
  CFA1X1 U1084 ( .A(n1255), .B(n1280), .CI(n1282), .CO(n1248), .S(n1249) );
  CFA1X1 U1087 ( .A(n1267), .B(n1290), .CI(n1263), .CO(n1254), .S(n1255) );
  CFA1X1 U1089 ( .A(n1292), .B(n1298), .CI(n1300), .CO(n1258), .S(n1259) );
  CFA1X1 U1090 ( .A(n1273), .B(n1296), .CI(n1294), .CO(n1260), .S(n1261) );
  CFA1X1 U1092 ( .A(n2127), .B(n2158), .CI(n2065), .CO(n1264), .S(n1265) );
  CFA1X1 U1095 ( .A(n1768), .B(n2189), .CI(n1973), .CO(n1270), .S(n1271) );
  COR2X1 U1097 ( .A(n1798), .B(n2034), .Z(n1272) );
  CFA1X1 U1098 ( .A(n1279), .B(n3900), .CI(n1306), .CO(n1274), .S(n1275) );
  CFA1X1 U1099 ( .A(n1283), .B(n1308), .CI(n1281), .CO(n1276), .S(n1277) );
  CFA1X1 U1104 ( .A(n1301), .B(n1299), .CI(n1293), .CO(n1286), .S(n1287) );
  CFA1X1 U1105 ( .A(n1322), .B(n1324), .CI(n1326), .CO(n1288), .S(n1289) );
  CFA1X1 U1106 ( .A(n1303), .B(n1328), .CI(n1330), .CO(n1290), .S(n1291) );
  CFA1X1 U1107 ( .A(n1885), .B(n1944), .CI(n2035), .CO(n1292), .S(n1293) );
  CFA1X1 U1109 ( .A(n2128), .B(n2097), .CI(n1915), .CO(n1296), .S(n1297) );
  CFA1X1 U1110 ( .A(n2190), .B(n2159), .CI(n1974), .CO(n1298), .S(n1299) );
  CFA1X1 U1111 ( .A(n2221), .B(n1799), .CI(n2004), .CO(n1300), .S(n1301) );
  CHA1X1 U1112 ( .A(n1724), .B(n1769), .CO(n1302), .S(n1303) );
  CFA1X1 U1117 ( .A(n1346), .B(n1321), .CI(n1344), .CO(n1312), .S(n1313) );
  CFA1X1 U1120 ( .A(n1352), .B(n1354), .CI(n1356), .CO(n1318), .S(n1319) );
  CFA1X1 U1121 ( .A(n2129), .B(n1350), .CI(n3955), .CO(n1320), .S(n1321) );
  CFA1X1 U1122 ( .A(n2067), .B(n2160), .CI(n2098), .CO(n1322), .S(n1323) );
  CFA1X1 U1123 ( .A(n1916), .B(n1975), .CI(n1945), .CO(n1324), .S(n1325) );
  CFA1X1 U1126 ( .A(n1770), .B(n2036), .CI(n1829), .CO(n1330), .S(n1331) );
  CFA1X1 U1128 ( .A(n1341), .B(n1364), .CI(n1339), .CO(n1334), .S(n1335) );
  CFA1X1 U1131 ( .A(n1374), .B(n1372), .CI(n1349), .CO(n1340), .S(n1341) );
  CFA1X1 U1132 ( .A(n1355), .B(n1357), .CI(n1353), .CO(n1342), .S(n1343) );
  CFA1X1 U1134 ( .A(n1384), .B(n1380), .CI(n1382), .CO(n1346), .S(n1347) );
  CFA1X1 U1135 ( .A(n2006), .B(n1359), .CI(n2068), .CO(n1348), .S(n1349) );
  CFA1X1 U1136 ( .A(n2099), .B(n1976), .CI(n1917), .CO(n1350), .S(n1351) );
  CFA1X1 U1137 ( .A(n1830), .B(n1887), .CI(n1858), .CO(n1352), .S(n1353) );
  CFA1X1 U1138 ( .A(n2130), .B(n1946), .CI(n2161), .CO(n1354), .S(n1355) );
  CFA1X1 U1139 ( .A(n2037), .B(n2223), .CI(n2192), .CO(n1356), .S(n1357) );
  CFA1X1 U1141 ( .A(n1365), .B(n1363), .CI(n1388), .CO(n1360), .S(n1361) );
  CFA1X1 U1142 ( .A(n1392), .B(n1390), .CI(n1367), .CO(n1362), .S(n1363) );
  CFA1X1 U1143 ( .A(n1371), .B(n1369), .CI(n1394), .CO(n1364), .S(n1365) );
  CFA1X1 U1145 ( .A(n1400), .B(n1398), .CI(n1379), .CO(n1368), .S(n1369) );
  CFA1X1 U1147 ( .A(n1406), .B(n1385), .CI(n1408), .CO(n1372), .S(n1373) );
  CFA1X1 U1148 ( .A(n1410), .B(n1404), .CI(n1402), .CO(n1374), .S(n1375) );
  CFA1X1 U1149 ( .A(n2100), .B(n2038), .CI(n1977), .CO(n1376), .S(n1377) );
  CFA1X1 U1150 ( .A(n2131), .B(n1947), .CI(n1918), .CO(n1378), .S(n1379) );
  CFA1X1 U1151 ( .A(n2162), .B(n1888), .CI(n1831), .CO(n1380), .S(n1381) );
  CFA1X1 U1152 ( .A(n2007), .B(n2224), .CI(n2193), .CO(n1382), .S(n1383) );
  CFA1X1 U1153 ( .A(n1802), .B(n2069), .CI(n1859), .CO(n1384), .S(n1385) );
  CFA1X1 U1155 ( .A(n1395), .B(n1416), .CI(n1393), .CO(n1388), .S(n1389) );
  CFA1X1 U1156 ( .A(n1420), .B(n1418), .CI(n1397), .CO(n1390), .S(n1391) );
  CFA1X1 U1157 ( .A(n1401), .B(n1399), .CI(n1422), .CO(n1392), .S(n1393) );
  CFA1X1 U1163 ( .A(n2163), .B(n1948), .CI(n1919), .CO(n1404), .S(n1405) );
  CFA1X1 U1164 ( .A(n2008), .B(n2194), .CI(n1889), .CO(n1406), .S(n1407) );
  CFA1X1 U1165 ( .A(n1860), .B(n2039), .CI(n2225), .CO(n1408), .S(n1409) );
  CFA1X1 U1169 ( .A(n1425), .B(n1421), .CI(n1423), .CO(n1416), .S(n1417) );
  CFA1X1 U1171 ( .A(n1431), .B(n1427), .CI(n1433), .CO(n1420), .S(n1421) );
  CFA1X1 U1172 ( .A(n1454), .B(n1429), .CI(n1435), .CO(n1422), .S(n1423) );
  CFA1X1 U1173 ( .A(n1456), .B(n1452), .CI(n1450), .CO(n1424), .S(n1425) );
  CFA1X1 U1174 ( .A(n3794), .B(n1458), .CI(n2102), .CO(n1426), .S(n1427) );
  CFA1X1 U1178 ( .A(n1833), .B(n1890), .CI(n2071), .CO(n1434), .S(n1435) );
  CFA1X1 U1181 ( .A(n1468), .B(n1445), .CI(n1447), .CO(n1440), .S(n1441) );
  CFA1X1 U1182 ( .A(n1472), .B(n1449), .CI(n1470), .CO(n1442), .S(n1443) );
  CFA1X1 U1185 ( .A(n1459), .B(n1478), .CI(n1480), .CO(n1448), .S(n1449) );
  CFA1X1 U1186 ( .A(n2041), .B(n2134), .CI(n2103), .CO(n1450), .S(n1451) );
  CFA1X1 U1187 ( .A(n2010), .B(n2165), .CI(n1950), .CO(n1452), .S(n1453) );
  CFA1X1 U1188 ( .A(n1891), .B(n1921), .CI(n1980), .CO(n1454), .S(n1455) );
  CFA1X1 U1189 ( .A(n2072), .B(n2227), .CI(n2196), .CO(n1456), .S(n1457) );
  CFA1X1 U1191 ( .A(n1465), .B(n1463), .CI(n1484), .CO(n1460), .S(n1461) );
  CFA1X1 U1195 ( .A(n1475), .B(n1477), .CI(n1479), .CO(n1468), .S(n1469) );
  CFA1X1 U1196 ( .A(n1498), .B(n1481), .CI(n1496), .CO(n1470), .S(n1471) );
  CFA1X1 U1197 ( .A(n2104), .B(n1500), .CI(n1502), .CO(n1472), .S(n1473) );
  CFA1X1 U1198 ( .A(n2135), .B(n2011), .CI(n1981), .CO(n1474), .S(n1475) );
  CFA1X1 U1199 ( .A(n2197), .B(n2166), .CI(n1951), .CO(n1476), .S(n1477) );
  CFA1X1 U1200 ( .A(n1892), .B(n2042), .CI(n2228), .CO(n1478), .S(n1479) );
  CFA1X1 U1201 ( .A(n1863), .B(n2073), .CI(n1922), .CO(n1480), .S(n1481) );
  CFA1X1 U1202 ( .A(n1487), .B(n1485), .CI(n1506), .CO(n1482), .S(n1483) );
  CFA1X1 U1206 ( .A(n1520), .B(n1499), .CI(n1497), .CO(n1490), .S(n1491) );
  CFA1X1 U1207 ( .A(n1518), .B(n1522), .CI(n1516), .CO(n1492), .S(n1493) );
  CFA1X1 U1208 ( .A(n2105), .B(n1503), .CI(n2043), .CO(n1494), .S(n1495) );
  CFA1X1 U1209 ( .A(n2136), .B(n1982), .CI(n1952), .CO(n1496), .S(n1497) );
  CFA1X1 U1210 ( .A(n2012), .B(n2167), .CI(n2198), .CO(n1498), .S(n1499) );
  CFA1X1 U1211 ( .A(n2074), .B(n2229), .CI(n1923), .CO(n1500), .S(n1501) );
  CFA1X1 U1214 ( .A(n1513), .B(n1528), .CI(n1511), .CO(n1506), .S(n1507) );
  CFA1X1 U1215 ( .A(n1515), .B(n1530), .CI(n1532), .CO(n1508), .S(n1509) );
  CFA1X1 U1216 ( .A(n1519), .B(n1534), .CI(n1521), .CO(n1510), .S(n1511) );
  CFA1X1 U1217 ( .A(n1536), .B(n1517), .CI(n1523), .CO(n1512), .S(n1513) );
  CFA1X1 U1218 ( .A(n1542), .B(n1538), .CI(n1540), .CO(n1514), .S(n1515) );
  CFA1X1 U1220 ( .A(n1983), .B(n2013), .CI(n2199), .CO(n1518), .S(n1519) );
  CFA1X1 U1221 ( .A(n2044), .B(n2230), .CI(n1924), .CO(n1520), .S(n1521) );
  CFA1X1 U1222 ( .A(n1894), .B(n1953), .CI(n2106), .CO(n1522), .S(n1523) );
  CFA1X1 U1223 ( .A(n1529), .B(n1527), .CI(n1546), .CO(n1524), .S(n1525) );
  CFA1X1 U1224 ( .A(n1533), .B(n1548), .CI(n1531), .CO(n1526), .S(n1527) );
  CFA1X1 U1225 ( .A(n1552), .B(n1550), .CI(n1535), .CO(n1528), .S(n1529) );
  CFA1X1 U1226 ( .A(n1541), .B(n1554), .CI(n1539), .CO(n1530), .S(n1531) );
  CFA1X1 U1227 ( .A(n1558), .B(n1537), .CI(n1556), .CO(n1532), .S(n1533) );
  CFA1X1 U1228 ( .A(n2045), .B(n1560), .CI(n1543), .CO(n1534), .S(n1535) );
  CFA1X1 U1229 ( .A(n2107), .B(n1984), .CI(n1954), .CO(n1536), .S(n1537) );
  CFA1X1 U1230 ( .A(n2138), .B(n2014), .CI(n2169), .CO(n1538), .S(n1539) );
  CFA1X1 U1231 ( .A(n2231), .B(n2200), .CI(n2076), .CO(n1540), .S(n1541) );
  CHA1X1 U1232 ( .A(n1729), .B(n1925), .CO(n1542), .S(n1543) );
  CFA1X1 U1233 ( .A(n1549), .B(n3209), .CI(n1564), .CO(n1544), .S(n1545) );
  CFA1X1 U1235 ( .A(n1555), .B(n1568), .CI(n1570), .CO(n1548), .S(n1549) );
  CFA1X1 U1236 ( .A(n1561), .B(n1557), .CI(n1559), .CO(n1550), .S(n1551) );
  CFA1X1 U1237 ( .A(n1576), .B(n1574), .CI(n1572), .CO(n1552), .S(n1553) );
  CFA1X1 U1239 ( .A(n2201), .B(n3151), .CI(n2015), .CO(n1556), .S(n1557) );
  CFA1X1 U1240 ( .A(n2077), .B(n2232), .CI(n1955), .CO(n1558), .S(n1559) );
  CFA1X1 U1241 ( .A(n1926), .B(n2108), .CI(n1985), .CO(n1560), .S(n1561) );
  CFA1X1 U1242 ( .A(n1567), .B(n1565), .CI(n1582), .CO(n1562), .S(n1563) );
  CFA1X1 U1244 ( .A(n1577), .B(n1586), .CI(n1588), .CO(n1566), .S(n1567) );
  CFA1X1 U1246 ( .A(n1592), .B(n1579), .CI(n1594), .CO(n1570), .S(n1571) );
  CFA1X1 U1247 ( .A(n2171), .B(n2140), .CI(n2047), .CO(n1572), .S(n1573) );
  CFA1X1 U1248 ( .A(n2078), .B(n2016), .CI(n2202), .CO(n1574), .S(n1575) );
  CFA1X1 U1249 ( .A(n2109), .B(n2233), .CI(n1986), .CO(n1576), .S(n1577) );
  CFA1X1 U1251 ( .A(n1585), .B(n1583), .CI(n1598), .CO(n1580), .S(n1581) );
  CFA1X1 U1253 ( .A(n1593), .B(n1602), .CI(n1604), .CO(n1584), .S(n1585) );
  CFA1X1 U1255 ( .A(n3125), .B(n1608), .CI(n1610), .CO(n1588), .S(n1589) );
  CFA1X1 U1256 ( .A(n2079), .B(n2203), .CI(n2048), .CO(n1590), .S(n1591) );
  CFA1X1 U1257 ( .A(n2110), .B(n2234), .CI(n1987), .CO(n1592), .S(n1593) );
  CFA1X1 U1259 ( .A(n1601), .B(n1599), .CI(n1614), .CO(n1596), .S(n1597) );
  CFA1X1 U1260 ( .A(n1605), .B(n1616), .CI(n1603), .CO(n1598), .S(n1599) );
  CFA1X1 U1261 ( .A(n1607), .B(n1618), .CI(n1609), .CO(n1600), .S(n1601) );
  CFA1X1 U1262 ( .A(n1624), .B(n1622), .CI(n1620), .CO(n1602), .S(n1603) );
  CFA1X1 U1264 ( .A(n2049), .B(n2080), .CI(n2018), .CO(n1606), .S(n1607) );
  CFA1X1 U1265 ( .A(n2111), .B(n2235), .CI(n2204), .CO(n1608), .S(n1609) );
  CHA1X1 U1266 ( .A(n1731), .B(n1988), .CO(n1610), .S(n1611) );
  CFA1X1 U1267 ( .A(n1617), .B(n1615), .CI(n1628), .CO(n1612), .S(n1613) );
  CFA1X1 U1268 ( .A(n1632), .B(n1630), .CI(n1619), .CO(n1614), .S(n1615) );
  CFA1X1 U1269 ( .A(n1625), .B(n1621), .CI(n1623), .CO(n1616), .S(n1617) );
  CFA1X1 U1272 ( .A(n2236), .B(n2112), .CI(n2019), .CO(n1622), .S(n1623) );
  CFA1X1 U1274 ( .A(n1631), .B(n1629), .CI(n1642), .CO(n1626), .S(n1627) );
  CFA1X1 U1275 ( .A(n1646), .B(n1644), .CI(n1633), .CO(n1628), .S(n1629) );
  CFA1X1 U1276 ( .A(n1648), .B(n1637), .CI(n1635), .CO(n1630), .S(n1631) );
  CFA1X1 U1277 ( .A(n2175), .B(n1650), .CI(n1639), .CO(n1632), .S(n1633) );
  CHA1X1 U1280 ( .A(n2051), .B(n2020), .CO(n1638), .S(n1639) );
  CFA1X1 U1281 ( .A(n1645), .B(n1643), .CI(n1654), .CO(n1640), .S(n1641) );
  CFA1X1 U1282 ( .A(n1649), .B(n1656), .CI(n1647), .CO(n1642), .S(n1643) );
  CFA1X1 U1283 ( .A(n1660), .B(n1651), .CI(n1658), .CO(n1644), .S(n1645) );
  CFA1X1 U1284 ( .A(n2207), .B(n1662), .CI(n2114), .CO(n1646), .S(n1647) );
  CFA1X1 U1285 ( .A(n3473), .B(n2238), .CI(n3070), .CO(n1648), .S(n1649) );
  CFA1X1 U1286 ( .A(n2021), .B(n3488), .CI(n2083), .CO(n1650), .S(n1651) );
  CFA1X1 U1287 ( .A(n1657), .B(n1655), .CI(n1666), .CO(n1652), .S(n1653) );
  CFA1X1 U1288 ( .A(n1659), .B(n1668), .CI(n1661), .CO(n1654), .S(n1655) );
  CFA1X1 U1289 ( .A(n1663), .B(n1670), .CI(n1672), .CO(n1656), .S(n1657) );
  CFA1X1 U1291 ( .A(n2146), .B(n2239), .CI(n2208), .CO(n1660), .S(n1661) );
  CHA1X1 U1292 ( .A(n2084), .B(n2053), .CO(n1662), .S(n1663) );
  CFA1X1 U1293 ( .A(n1676), .B(n1667), .CI(n1669), .CO(n1664), .S(n1665) );
  CFA1X1 U1294 ( .A(n1673), .B(n1678), .CI(n1671), .CO(n1666), .S(n1667) );
  CFA1X1 U1295 ( .A(n2209), .B(n1680), .CI(n1682), .CO(n1668), .S(n1669) );
  CFA1X1 U1296 ( .A(n2147), .B(n2240), .CI(n2085), .CO(n1670), .S(n1671) );
  CFA1X1 U1297 ( .A(n2054), .B(n2178), .CI(n2116), .CO(n1672), .S(n1673) );
  CFA1X1 U1298 ( .A(n1679), .B(n1677), .CI(n1686), .CO(n1674), .S(n1675) );
  CFA1X1 U1299 ( .A(n1690), .B(n1681), .CI(n1688), .CO(n1676), .S(n1677) );
  CFA1X1 U1300 ( .A(n2148), .B(n1683), .CI(n1734), .CO(n1678), .S(n1679) );
  CFA1X1 U1301 ( .A(n2179), .B(n2241), .CI(n2210), .CO(n1680), .S(n1681) );
  CFA1X1 U1303 ( .A(n1689), .B(n1687), .CI(n1694), .CO(n1684), .S(n1685) );
  CFA1X1 U1304 ( .A(n1698), .B(n1691), .CI(n1696), .CO(n1686), .S(n1687) );
  CFA1X1 U1305 ( .A(n2180), .B(n2242), .CI(n2118), .CO(n1688), .S(n1689) );
  CFA1X1 U1306 ( .A(n2087), .B(n2211), .CI(n2149), .CO(n1690), .S(n1691) );
  CFA1X1 U1307 ( .A(n1697), .B(n1695), .CI(n1702), .CO(n1692), .S(n1693) );
  CFA1X1 U1308 ( .A(n2212), .B(n1704), .CI(n1699), .CO(n1694), .S(n1695) );
  CFA1X1 U1309 ( .A(n2181), .B(n2243), .CI(n3337), .CO(n1696), .S(n1697) );
  CHA1X1 U1310 ( .A(n2150), .B(n2119), .CO(n1698), .S(n1699) );
  CFA1X1 U1311 ( .A(n1708), .B(n1703), .CI(n1705), .CO(n1700), .S(n1701) );
  CFA1X1 U1312 ( .A(n2182), .B(n1710), .CI(n2244), .CO(n1702), .S(n1703) );
  CFA1X1 U1313 ( .A(n2120), .B(n2213), .CI(n2151), .CO(n1704), .S(n1705) );
  CFA1X1 U1314 ( .A(n1711), .B(n1709), .CI(n1714), .CO(n1706), .S(n1707) );
  CFA1X1 U1315 ( .A(n2214), .B(n2245), .CI(n2183), .CO(n1708), .S(n1709) );
  CHA1X1 U1316 ( .A(n1736), .B(n2152), .CO(n1710), .S(n1711) );
  CFA1X1 U1317 ( .A(n2246), .B(n1715), .CI(n1718), .CO(n1712), .S(n1713) );
  CFA1X1 U1318 ( .A(n2215), .B(n2153), .CI(n2184), .CO(n1714), .S(n1715) );
  CFA1X1 U1319 ( .A(n2216), .B(n1719), .CI(n2247), .CO(n1716), .S(n1717) );
  CHA1X1 U1320 ( .A(n1737), .B(n2185), .CO(n1718), .S(n1719) );
  CFA1X1 U1321 ( .A(n2186), .B(n2248), .CI(n2217), .CO(n1720), .S(n1721) );
  CHA1X1 U1322 ( .A(n1738), .B(n2249), .CO(n1722), .S(n1723) );
  COND2X1 U1323 ( .A(n144), .B(n3921), .C(net16617), .D(n2284), .Z(n1724) );
  COND2X1 U1332 ( .A(net18570), .B(n2260), .C(net16617), .D(n2259), .Z(n1746)
         );
  COND2X1 U1333 ( .A(n3705), .B(n2261), .C(net16617), .D(n2260), .Z(n1747) );
  COND2X1 U1335 ( .A(net18570), .B(n2263), .C(net16617), .D(n2262), .Z(n1749)
         );
  COND2X1 U1339 ( .A(n3705), .B(n2267), .C(net16617), .D(n2266), .Z(n1753) );
  COND2X1 U1340 ( .A(n3705), .B(n2268), .C(net16617), .D(n2267), .Z(n1754) );
  COND2X1 U1341 ( .A(n144), .B(n2269), .C(net16617), .D(n2268), .Z(n1755) );
  COND2X1 U1342 ( .A(net18570), .B(n2270), .C(net16617), .D(n2269), .Z(n1756)
         );
  COND2X1 U1343 ( .A(n3705), .B(n2271), .C(net16617), .D(n2270), .Z(n1757) );
  COND2X1 U1344 ( .A(net18570), .B(n2272), .C(net16617), .D(n2271), .Z(n1758)
         );
  COND2X1 U1346 ( .A(n3705), .B(n2274), .C(net16617), .D(n2273), .Z(n1760) );
  COND2X1 U1348 ( .A(net18570), .B(n2276), .C(net16617), .D(n2275), .Z(n1762)
         );
  COND2X1 U1349 ( .A(net18570), .B(n2277), .C(net16617), .D(n2276), .Z(n1763)
         );
  COND2X1 U1350 ( .A(net18570), .B(n2278), .C(net16617), .D(n2277), .Z(n1764)
         );
  COND2X1 U1354 ( .A(net18570), .B(n2282), .C(net16617), .D(n2281), .Z(n1768)
         );
  COND2X1 U1355 ( .A(n144), .B(n2283), .C(net16617), .D(n2282), .Z(n1769) );
  CND2IX1 U1389 ( .B(n3998), .A(n3920), .Z(n2284) );
  CAOR1X1 U1391 ( .A(net18772), .B(n3915), .C(n2285), .Z(n1771) );
  COND2X1 U1393 ( .A(n2286), .B(net18772), .C(n2287), .D(n3915), .Z(n1773) );
  COND2X1 U1395 ( .A(n3915), .B(n2289), .C(net18772), .D(n2288), .Z(n1774) );
  COND2X1 U1396 ( .A(n3915), .B(n2290), .C(net18772), .D(n2289), .Z(n1775) );
  COND2X1 U1399 ( .A(n3915), .B(n2293), .C(net18772), .D(n2292), .Z(n1778) );
  COND2X1 U1400 ( .A(n3915), .B(n2294), .C(net18772), .D(n2293), .Z(n1779) );
  COND2X1 U1402 ( .A(net18573), .B(n2296), .C(net18772), .D(n2295), .Z(n1781)
         );
  COND2X1 U1403 ( .A(net18573), .B(n2297), .C(net18772), .D(n2296), .Z(n1782)
         );
  COND2X1 U1404 ( .A(n3915), .B(n2298), .C(net18772), .D(n2297), .Z(n1783) );
  COND2X1 U1405 ( .A(net18573), .B(n2299), .C(net18772), .D(n2298), .Z(n1784)
         );
  COND2X1 U1406 ( .A(n3915), .B(n2300), .C(net18772), .D(n2299), .Z(n1785) );
  COND2X1 U1407 ( .A(n3915), .B(n2301), .C(net18772), .D(n2300), .Z(n1786) );
  COND2X1 U1409 ( .A(net18573), .B(n2303), .C(net18772), .D(n2302), .Z(n1788)
         );
  COND2X1 U1411 ( .A(n3915), .B(n2305), .C(net18772), .D(n2304), .Z(n1790) );
  COND2X1 U1414 ( .A(n2308), .B(net18573), .C(net18772), .D(n2307), .Z(n1793)
         );
  COND2X1 U1415 ( .A(n135), .B(n2309), .C(net18772), .D(n2308), .Z(n1794) );
  COND2X1 U1416 ( .A(n3710), .B(net18573), .C(net18772), .D(n2309), .Z(n1795)
         );
  COND2X1 U1418 ( .A(n135), .B(n2312), .C(net18772), .D(n3507), .Z(n1797) );
  COND2X1 U1419 ( .A(net18573), .B(n2313), .C(net18772), .D(n2312), .Z(n1798)
         );
  COND2X1 U1420 ( .A(n3915), .B(n2314), .C(net18772), .D(n2313), .Z(n1799) );
  COND2X1 U1421 ( .A(n3915), .B(n2315), .C(net18772), .D(n2314), .Z(n1800) );
  CND2IX1 U1456 ( .B(n3998), .A(net15963), .Z(n2317) );
  COND2X1 U1459 ( .A(n2319), .B(n3682), .C(net16623), .D(n2318), .Z(n1804) );
  COND2X1 U1460 ( .A(n2319), .B(net16623), .C(n2320), .D(n3682), .Z(n1805) );
  COND2X1 U1461 ( .A(n3682), .B(n2321), .C(net16623), .D(n2320), .Z(n824) );
  COND2X1 U1462 ( .A(n3682), .B(n2322), .C(net16623), .D(n2321), .Z(n1806) );
  COND2X1 U1463 ( .A(n3682), .B(n2323), .C(net16623), .D(n2322), .Z(n842) );
  COND2X1 U1464 ( .A(n3682), .B(n2324), .C(net16623), .D(n2323), .Z(n1807) );
  COND2X1 U1465 ( .A(n3682), .B(n2325), .C(net16623), .D(n2324), .Z(n1808) );
  COND2X1 U1467 ( .A(n3682), .B(n2327), .C(net16623), .D(n2326), .Z(n1810) );
  COND2X1 U1468 ( .A(n3682), .B(n2328), .C(net16623), .D(n2327), .Z(n1811) );
  COND2X1 U1469 ( .A(n3682), .B(n2329), .C(net16623), .D(n2328), .Z(n1812) );
  COND2X1 U1471 ( .A(n3682), .B(n2331), .C(net16623), .D(n2330), .Z(n1814) );
  COND2X1 U1472 ( .A(n3682), .B(n2332), .C(net16623), .D(n2331), .Z(n1815) );
  COND2X1 U1473 ( .A(n3682), .B(n2333), .C(net16623), .D(n2332), .Z(n1816) );
  COND2X1 U1474 ( .A(n126), .B(n2334), .C(net16621), .D(n2333), .Z(n1817) );
  COND2X1 U1476 ( .A(n3682), .B(n2336), .C(net16623), .D(n2335), .Z(n1819) );
  COND2X1 U1477 ( .A(n3682), .B(n2337), .C(net16623), .D(n2336), .Z(n1820) );
  COND2X1 U1478 ( .A(n3682), .B(n2338), .C(net16623), .D(n2337), .Z(n1821) );
  COND2X1 U1479 ( .A(n3682), .B(n2339), .C(net16623), .D(n2338), .Z(n1822) );
  COND2X1 U1480 ( .A(n3682), .B(n2340), .C(net16623), .D(n2339), .Z(n1823) );
  COND2X1 U1481 ( .A(n3682), .B(n2341), .C(net16623), .D(n2340), .Z(n1824) );
  COND2X1 U1482 ( .A(n3682), .B(n3485), .C(net16623), .D(n2341), .Z(n1825) );
  COND2X1 U1483 ( .A(n3682), .B(n2343), .C(net16623), .D(n2342), .Z(n1826) );
  COND2X1 U1487 ( .A(n3682), .B(n2347), .C(net16623), .D(n2346), .Z(n1830) );
  COND2X1 U1488 ( .A(n3682), .B(n2348), .C(net16623), .D(n2347), .Z(n1831) );
  COND2X1 U1489 ( .A(n3682), .B(n2349), .C(net16623), .D(n2348), .Z(n1832) );
  COND2X1 U1531 ( .A(n3172), .B(n2357), .C(n2356), .D(net16605), .Z(n1839) );
  COND2X1 U1532 ( .A(n3173), .B(n2358), .C(net16606), .D(n2357), .Z(n890) );
  COND2X1 U1534 ( .A(n3172), .B(n2360), .C(net16605), .D(n2359), .Z(n920) );
  COND2X1 U1535 ( .A(n3172), .B(n2361), .C(net16606), .D(n2360), .Z(n1841) );
  COND2X1 U1537 ( .A(n117), .B(n2363), .C(net16605), .D(n2362), .Z(n1843) );
  COND2X1 U1538 ( .A(n3172), .B(n2364), .C(net16605), .D(n2363), .Z(n1844) );
  COND2X1 U1540 ( .A(n3173), .B(n2366), .C(n2365), .D(net16606), .Z(n1846) );
  COND2X1 U1541 ( .A(n3172), .B(n2367), .C(net16605), .D(n2366), .Z(n1847) );
  COND2X1 U1542 ( .A(n3173), .B(n2368), .C(n2367), .D(net16605), .Z(n1848) );
  COND2X1 U1543 ( .A(n3173), .B(n2369), .C(n2368), .D(net16605), .Z(n1849) );
  COND2X1 U1544 ( .A(n3172), .B(n2370), .C(n2369), .D(net16606), .Z(n1850) );
  COND2X1 U1545 ( .A(n3172), .B(n2371), .C(net16605), .D(n2370), .Z(n1851) );
  COND2X1 U1550 ( .A(n3173), .B(n2376), .C(n2375), .D(net16605), .Z(n1856) );
  COND2X1 U1551 ( .A(n3172), .B(n2377), .C(net16605), .D(n2376), .Z(n1857) );
  COND2X1 U1552 ( .A(n3173), .B(n2378), .C(net16605), .D(n2377), .Z(n1858) );
  COND2X1 U1554 ( .A(n117), .B(n2380), .C(net16605), .D(n2379), .Z(n1860) );
  COND2X1 U1555 ( .A(net18572), .B(n3050), .C(net21572), .D(n2380), .Z(n1861)
         );
  CAOR1X1 U1592 ( .A(n3479), .B(n3747), .C(n2384), .Z(n1864) );
  COND2X1 U1593 ( .A(n2385), .B(n108), .C(n3479), .D(n2384), .Z(n1865) );
  COND2X1 U1594 ( .A(n2385), .B(n3472), .C(n2386), .D(n108), .Z(n1866) );
  COND2X1 U1595 ( .A(n3747), .B(n2387), .C(n3472), .D(n2386), .Z(n1867) );
  COND2X1 U1596 ( .A(n108), .B(n2388), .C(n3472), .D(n2387), .Z(n1868) );
  COND2X1 U1597 ( .A(n3747), .B(n2389), .C(n3957), .D(n2388), .Z(n1869) );
  COND2X1 U1598 ( .A(n3747), .B(n2390), .C(n3957), .D(n2389), .Z(n1870) );
  COND2X1 U1599 ( .A(n108), .B(n2391), .C(n3472), .D(n2390), .Z(n1871) );
  COND2X1 U1600 ( .A(n3747), .B(n2392), .C(n3957), .D(n2391), .Z(n1872) );
  COND2X1 U1602 ( .A(n2394), .B(n3747), .C(n3957), .D(n2393), .Z(n1873) );
  COND2X1 U1604 ( .A(n108), .B(n2396), .C(n3957), .D(n2395), .Z(n1874) );
  COND2X1 U1607 ( .A(n108), .B(n2399), .C(n3957), .D(n2398), .Z(n1877) );
  COND2X1 U1609 ( .A(n3747), .B(n2401), .C(n3957), .D(n2400), .Z(n1879) );
  COND2X1 U1610 ( .A(n108), .B(n2402), .C(n3957), .D(n2401), .Z(n1880) );
  COND2X1 U1611 ( .A(n108), .B(n2403), .C(n3957), .D(n2402), .Z(n1881) );
  COND2X1 U1612 ( .A(n108), .B(n2404), .C(n3957), .D(n2403), .Z(n1882) );
  COND2X1 U1613 ( .A(n3747), .B(n2405), .C(n3957), .D(n2404), .Z(n1883) );
  COND2X1 U1617 ( .A(n108), .B(n2409), .C(n3957), .D(n2408), .Z(n1887) );
  COND2X1 U1618 ( .A(n3747), .B(n2410), .C(n3957), .D(n2409), .Z(n1888) );
  COND2X1 U1619 ( .A(n108), .B(n2411), .C(n3957), .D(n2410), .Z(n1889) );
  COND2X1 U1621 ( .A(n2413), .B(n3747), .C(n3957), .D(n2412), .Z(n1891) );
  COND2X1 U1622 ( .A(n3747), .B(n2414), .C(n3957), .D(n2413), .Z(n1892) );
  CND2IX1 U1657 ( .B(n3998), .A(net18520), .Z(n2416) );
  COND2X1 U1658 ( .A(n3332), .B(net19200), .C(n3333), .D(n2449), .Z(n1729) );
  COND2X1 U1662 ( .A(n3331), .B(n2420), .C(n3023), .D(n2419), .Z(n1898) );
  COND2X1 U1663 ( .A(n3331), .B(n2421), .C(n3335), .D(n2420), .Z(n1899) );
  COND2X1 U1665 ( .A(n3332), .B(n2423), .C(n3333), .D(n2422), .Z(n1901) );
  COND2X1 U1666 ( .A(n3332), .B(n2424), .C(n3334), .D(n2423), .Z(n1902) );
  COND2X1 U1667 ( .A(n3336), .B(n2425), .C(n3335), .D(n2424), .Z(n1903) );
  COND2X1 U1668 ( .A(n3332), .B(n2426), .C(n3334), .D(n2425), .Z(n1904) );
  COND2X1 U1669 ( .A(n99), .B(n2427), .C(n3333), .D(n2426), .Z(n1905) );
  COND2X1 U1671 ( .A(n3331), .B(n2429), .C(n3023), .D(n2428), .Z(n1906) );
  COND2X1 U1672 ( .A(n3331), .B(n2430), .C(n3334), .D(n2429), .Z(n1907) );
  COND2X1 U1673 ( .A(n3332), .B(n2431), .C(n3023), .D(n2430), .Z(n1908) );
  COND2X1 U1674 ( .A(n3336), .B(n2432), .C(n3023), .D(n2431), .Z(n1909) );
  COND2X1 U1675 ( .A(n3331), .B(n2433), .C(n3334), .D(n2432), .Z(n1910) );
  COND2X1 U1676 ( .A(n3336), .B(n2434), .C(n3023), .D(n2433), .Z(n1911) );
  COND2X1 U1677 ( .A(n3331), .B(n2435), .C(n3334), .D(n3486), .Z(n1912) );
  COND2X1 U1678 ( .A(n99), .B(n2436), .C(n3023), .D(n2435), .Z(n1913) );
  COND2X1 U1679 ( .A(n3332), .B(n2437), .C(n3335), .D(n2436), .Z(n1914) );
  COND2X1 U1680 ( .A(n99), .B(n2438), .C(n3023), .D(n2437), .Z(n1915) );
  COND2X1 U1681 ( .A(n3331), .B(n2439), .C(n3023), .D(n2438), .Z(n1916) );
  COND2X1 U1683 ( .A(n3331), .B(n2441), .C(n3023), .D(n2440), .Z(n1918) );
  COND2X1 U1684 ( .A(n99), .B(n2442), .C(n3023), .D(n2441), .Z(n1919) );
  COND2X1 U1686 ( .A(n3332), .B(n3802), .C(n3023), .D(n2443), .Z(n1921) );
  COND2X1 U1687 ( .A(n3332), .B(n2445), .C(n3023), .D(n2444), .Z(n1922) );
  COND2X1 U1688 ( .A(n3336), .B(n2446), .C(n3023), .D(n2445), .Z(n1923) );
  COND2X1 U1689 ( .A(n3331), .B(n2447), .C(n3333), .D(n2446), .Z(n1924) );
  COND2X1 U1690 ( .A(n2448), .B(n99), .C(n3333), .D(n2447), .Z(n1925) );
  COND2X1 U1732 ( .A(n3913), .B(n2456), .C(n87), .D(n2455), .Z(n1933) );
  COND2X1 U1733 ( .A(net22025), .B(n2457), .C(net19996), .D(n2456), .Z(n1934)
         );
  COND2X1 U1734 ( .A(net22025), .B(n3160), .C(net19996), .D(n2457), .Z(n1935)
         );
  COND2X1 U1736 ( .A(n3913), .B(n2460), .C(net19996), .D(n2459), .Z(n1937) );
  COND2X1 U1738 ( .A(net22025), .B(n2462), .C(net19996), .D(n2461), .Z(n1938)
         );
  COND2X1 U1739 ( .A(n90), .B(n2463), .C(net19996), .D(n2462), .Z(n1130) );
  COND2X1 U1742 ( .A(n90), .B(n2466), .C(net19422), .D(n2465), .Z(n1941) );
  COND2X1 U1744 ( .A(n90), .B(n2468), .C(net19422), .D(n2467), .Z(n1943) );
  COND2X1 U1746 ( .A(n90), .B(n2470), .C(net19996), .D(n2469), .Z(n1945) );
  COND2X1 U1747 ( .A(n90), .B(n2471), .C(net19422), .D(n2470), .Z(n1946) );
  COND2X1 U1749 ( .A(net22025), .B(n2473), .C(net19996), .D(n2472), .Z(n1948)
         );
  COND2X1 U1750 ( .A(net22025), .B(n2474), .C(net19422), .D(n2473), .Z(n1949)
         );
  COND2X1 U1751 ( .A(n90), .B(n2475), .C(net19422), .D(n2474), .Z(n1950) );
  COND2X1 U1752 ( .A(net22025), .B(n2476), .C(net19996), .D(n2475), .Z(n1951)
         );
  COND2X1 U1753 ( .A(net22025), .B(n2477), .C(net19996), .D(n2476), .Z(n1952)
         );
  COND2X1 U1754 ( .A(net22025), .B(n2478), .C(net19996), .D(n2477), .Z(n1953)
         );
  COND2X1 U1756 ( .A(net22025), .B(n2480), .C(net19996), .D(n2479), .Z(n1955)
         );
  CENX2 U1776 ( .A(n3988), .B(net16671), .Z(n2467) );
  COND2X1 U1792 ( .A(n3188), .B(n3493), .C(n3285), .D(n2515), .Z(n1731) );
  COND2X1 U1795 ( .A(n2484), .B(net18902), .C(n2485), .D(n3080), .Z(n1960) );
  COND2X1 U1796 ( .A(n3189), .B(n2486), .C(n3285), .D(n2485), .Z(n1961) );
  COND2X1 U1798 ( .A(n3189), .B(n2488), .C(n3484), .D(n2487), .Z(n1963) );
  COND2X1 U1799 ( .A(n3080), .B(n2489), .C(n3285), .D(n2488), .Z(n1964) );
  COND2X1 U1801 ( .A(n3189), .B(n2491), .C(n3285), .D(n2490), .Z(n1966) );
  COND2X1 U1803 ( .A(n3080), .B(n2493), .C(n3285), .D(n2492), .Z(n1968) );
  COND2X1 U1804 ( .A(n3080), .B(n2494), .C(n3285), .D(n2493), .Z(n1969) );
  COND2X1 U1805 ( .A(n3080), .B(n2495), .C(net21576), .D(n2494), .Z(n1970) );
  COND2X1 U1811 ( .A(n3189), .B(n2501), .C(n3285), .D(n2500), .Z(n1975) );
  COND2X1 U1812 ( .A(n3080), .B(n2502), .C(n3484), .D(n2501), .Z(n1976) );
  COND2X1 U1813 ( .A(n3080), .B(n2503), .C(net18902), .D(n2502), .Z(n1977) );
  COND2X1 U1814 ( .A(n3189), .B(n2504), .C(n3484), .D(n2503), .Z(n1978) );
  COND2X1 U1815 ( .A(n2505), .B(n81), .C(n3345), .D(n2504), .Z(n1979) );
  COND2X1 U1816 ( .A(n81), .B(n2506), .C(n3345), .D(n2505), .Z(n1980) );
  COND2X1 U1817 ( .A(n81), .B(n2507), .C(n3484), .D(n2506), .Z(n1981) );
  COND2X1 U1819 ( .A(n3189), .B(n2509), .C(net18902), .D(n2508), .Z(n1983) );
  COND2X1 U1820 ( .A(n3080), .B(n2510), .C(n3285), .D(n2509), .Z(n1984) );
  COND2X1 U1822 ( .A(n3189), .B(n2512), .C(n3285), .D(n2511), .Z(n1986) );
  COND2X1 U1823 ( .A(n2513), .B(n3188), .C(net18902), .D(n2512), .Z(n1987) );
  COND2X1 U1824 ( .A(n2514), .B(n3080), .C(n3285), .D(n2513), .Z(n1988) );
  COND2X1 U1865 ( .A(n2521), .B(net18612), .C(net16684), .D(n2520), .Z(n1995)
         );
  COND2X1 U1867 ( .A(n3340), .B(n2523), .C(net16683), .D(n2522), .Z(n1997) );
  COND2X1 U1868 ( .A(n2524), .B(net18612), .C(net16684), .D(n2523), .Z(n1998)
         );
  COND2X1 U1869 ( .A(n3026), .B(net18612), .C(net16684), .D(n2524), .Z(n1999)
         );
  COND2X1 U1870 ( .A(n2526), .B(net18612), .C(net16684), .D(n2525), .Z(n2000)
         );
  COND2X1 U1871 ( .A(net18612), .B(n2527), .C(net16684), .D(n2526), .Z(n2001)
         );
  COND2X1 U1872 ( .A(n3158), .B(n3044), .C(net16684), .D(n2527), .Z(n2002) );
  COND2X1 U1875 ( .A(n2531), .B(n3340), .C(net16683), .D(n3864), .Z(n2004) );
  COND2X1 U1879 ( .A(n2535), .B(n3044), .C(net16684), .D(n2534), .Z(n2008) );
  COND2X1 U1880 ( .A(n3340), .B(n2536), .C(net16683), .D(n2535), .Z(n2009) );
  COND2X1 U1881 ( .A(n2537), .B(net18613), .C(net16683), .D(n2536), .Z(n2010)
         );
  COND2X1 U1883 ( .A(n3044), .B(n2539), .C(net16684), .D(n2538), .Z(n2012) );
  COND2X1 U1884 ( .A(n2540), .B(n3044), .C(net16684), .D(n2539), .Z(n2013) );
  COND2X1 U1885 ( .A(n3044), .B(n2541), .C(net16684), .D(n2540), .Z(n2014) );
  COND2X1 U1890 ( .A(n3340), .B(n2546), .C(net16683), .D(n2545), .Z(n2019) );
  COND2X1 U1929 ( .A(n2550), .B(n3355), .C(n2551), .D(n63), .Z(n2024) );
  COND2X1 U1930 ( .A(n2552), .B(n3058), .C(n3355), .D(n2551), .Z(n2025) );
  COND2X1 U1931 ( .A(n63), .B(n2553), .C(n2552), .D(n3355), .Z(n2026) );
  COND2X1 U1932 ( .A(n63), .B(n2554), .C(n3355), .D(n2553), .Z(n2027) );
  COND2X1 U1934 ( .A(n3058), .B(n2556), .C(n3355), .D(n2555), .Z(n2029) );
  COND2X1 U1935 ( .A(n63), .B(n2557), .C(n3355), .D(n2556), .Z(n2030) );
  COND2X1 U1936 ( .A(n63), .B(n2558), .C(n3037), .D(n2557), .Z(n2031) );
  COND2X1 U1937 ( .A(n2559), .B(n3059), .C(n3355), .D(n2558), .Z(n2032) );
  COND2X1 U1938 ( .A(n2560), .B(n3916), .C(n2559), .D(n3918), .Z(n2033) );
  COND2X1 U1942 ( .A(n63), .B(n2564), .C(n3355), .D(n2563), .Z(n2037) );
  COND2X1 U1943 ( .A(n3059), .B(n2565), .C(n3037), .D(n2564), .Z(n2038) );
  COND2X1 U1945 ( .A(n3059), .B(n2567), .C(n3355), .D(n2566), .Z(n2040) );
  COND2X1 U1946 ( .A(n63), .B(n2568), .C(n3355), .D(n2567), .Z(n2041) );
  COND2X1 U1947 ( .A(n3058), .B(n2569), .C(n3571), .D(n2568), .Z(n2042) );
  COND2X1 U1949 ( .A(n3059), .B(n2571), .C(n3055), .D(n2570), .Z(n2044) );
  COND2X1 U1952 ( .A(n63), .B(n2574), .C(n3355), .D(n2573), .Z(n2047) );
  COND2X1 U1996 ( .A(n2583), .B(n3267), .C(n2584), .D(n3352), .Z(n2057) );
  COND2X1 U1998 ( .A(n3353), .B(n2586), .C(n51), .D(n3165), .Z(n2059) );
  COND2X1 U1999 ( .A(n3353), .B(n3036), .C(n3267), .D(n2586), .Z(n2060) );
  COND2X1 U2000 ( .A(n3352), .B(n2588), .C(n51), .D(n2587), .Z(n2061) );
  COND2X1 U2001 ( .A(n54), .B(n2589), .C(n3267), .D(n2588), .Z(n2062) );
  COND2X1 U2003 ( .A(n54), .B(n2591), .C(n3733), .D(n2590), .Z(n2064) );
  COND2X1 U2004 ( .A(n54), .B(n2592), .C(n3267), .D(n2591), .Z(n2065) );
  COND2X1 U2005 ( .A(n3912), .B(n2593), .C(n3267), .D(n2592), .Z(n2066) );
  COND2X1 U2006 ( .A(n54), .B(n2594), .C(n51), .D(n2593), .Z(n2067) );
  COND2X1 U2009 ( .A(n54), .B(n2597), .C(n51), .D(n2596), .Z(n2070) );
  COND2X1 U2011 ( .A(n2599), .B(n54), .C(n3267), .D(n3032), .Z(n2072) );
  COND2X1 U2012 ( .A(n3352), .B(n2600), .C(n51), .D(n2599), .Z(n2073) );
  COND2X1 U2013 ( .A(n54), .B(n2601), .C(n3267), .D(n2600), .Z(n2074) );
  COND2X1 U2015 ( .A(n2603), .B(n3912), .C(n3267), .D(n2602), .Z(n2076) );
  COND2X1 U2016 ( .A(n2604), .B(n3352), .C(n51), .D(n2603), .Z(n2077) );
  COND2X1 U2017 ( .A(n3353), .B(n3342), .C(n3267), .D(n2604), .Z(n2078) );
  COND2X1 U2018 ( .A(n3912), .B(n2606), .C(n3267), .D(n2605), .Z(n2079) );
  COND2X1 U2021 ( .A(n3353), .B(n2609), .C(n3267), .D(n2608), .Z(n2082) );
  COND2X1 U2022 ( .A(n3352), .B(n2610), .C(n51), .D(n2609), .Z(n2083) );
  COND2X1 U2024 ( .A(n3352), .B(n2612), .C(n3267), .D(n2611), .Z(n2085) );
  COND2X1 U2062 ( .A(n2616), .B(n3904), .C(n3832), .D(n2615), .Z(n2089) );
  COND2X1 U2063 ( .A(n2616), .B(n3833), .C(n2617), .D(n3904), .Z(n2090) );
  COND2X1 U2067 ( .A(n3903), .B(n2621), .C(n3832), .D(n2620), .Z(n2094) );
  COND2X1 U2068 ( .A(n3904), .B(n2622), .C(n3959), .D(n2621), .Z(n2095) );
  COND2X1 U2069 ( .A(n3904), .B(n2623), .C(n3832), .D(n2622), .Z(n2096) );
  COND2X1 U2070 ( .A(n3904), .B(n2624), .C(n3832), .D(n2623), .Z(n2097) );
  COND2X1 U2071 ( .A(n3904), .B(n2625), .C(n3833), .D(n2624), .Z(n2098) );
  COND2X1 U2072 ( .A(n3904), .B(n2626), .C(n42), .D(n2625), .Z(n2099) );
  COND2X1 U2073 ( .A(n3904), .B(n2627), .C(n3832), .D(n2626), .Z(n2100) );
  COND2X1 U2076 ( .A(n3903), .B(n2630), .C(n3833), .D(n2629), .Z(n2103) );
  COND2X1 U2079 ( .A(n3904), .B(n2633), .C(n3832), .D(n2632), .Z(n2106) );
  COND2X1 U2080 ( .A(n3904), .B(n2634), .C(n3832), .D(n2633), .Z(n2107) );
  COND2X1 U2081 ( .A(n3904), .B(n2635), .C(n3833), .D(n2634), .Z(n2108) );
  COND2X1 U2082 ( .A(n3904), .B(n2636), .C(n3832), .D(n2635), .Z(n2109) );
  COND2X1 U2083 ( .A(n3903), .B(n2637), .C(n2636), .D(n3833), .Z(n2110) );
  COND2X1 U2084 ( .A(n3904), .B(n2638), .C(n3832), .D(n2637), .Z(n2111) );
  COND2X1 U2085 ( .A(n3904), .B(n3035), .C(n3833), .D(n2638), .Z(n2112) );
  COND2X1 U2086 ( .A(n3903), .B(n2640), .C(n3832), .D(n2639), .Z(n2113) );
  COND2X1 U2088 ( .A(n3904), .B(n2642), .C(n3832), .D(n2641), .Z(n2115) );
  COND2X1 U2129 ( .A(n2649), .B(n36), .C(n3425), .D(n2648), .Z(n2122) );
  COND2X1 U2131 ( .A(n3163), .B(n2651), .C(n3424), .D(n2650), .Z(n2124) );
  COND2X1 U2135 ( .A(n36), .B(n2655), .C(n3425), .D(n2654), .Z(n2128) );
  COND2X1 U2137 ( .A(n3163), .B(n2657), .C(n3655), .D(n2656), .Z(n2130) );
  COND2X1 U2138 ( .A(n3163), .B(n2658), .C(n3424), .D(n2657), .Z(n2131) );
  COND2X1 U2142 ( .A(n36), .B(n2662), .C(n3424), .D(n2661), .Z(n2135) );
  COND2X1 U2143 ( .A(n3163), .B(n2663), .C(n3425), .D(n2662), .Z(n2136) );
  COND2X1 U2144 ( .A(n3163), .B(n2664), .C(n3425), .D(n2663), .Z(n2137) );
  COND2X1 U2145 ( .A(n3163), .B(n2665), .C(n3425), .D(n2664), .Z(n2138) );
  COND2X1 U2146 ( .A(n3163), .B(n2666), .C(n3425), .D(n2665), .Z(n2139) );
  COND2X1 U2147 ( .A(n3163), .B(n2667), .C(n3425), .D(n2666), .Z(n2140) );
  COND2X1 U2149 ( .A(n3163), .B(n2669), .C(n3655), .D(n2668), .Z(n2142) );
  COND2X1 U2153 ( .A(n3163), .B(n2673), .C(n3425), .D(n2672), .Z(n2146) );
  COND2X1 U2154 ( .A(n3163), .B(n2674), .C(n3424), .D(n2673), .Z(n2147) );
  COND2X1 U2155 ( .A(n3163), .B(n2675), .C(n3424), .D(n2674), .Z(n2148) );
  COND2X1 U2156 ( .A(n3163), .B(n2676), .C(n3655), .D(n2675), .Z(n2149) );
  COND2X1 U2157 ( .A(n3163), .B(n2677), .C(n3424), .D(n2676), .Z(n2150) );
  CAOR1X1 U2195 ( .A(net18545), .B(n27), .C(n2681), .Z(n2154) );
  COND2X1 U2198 ( .A(n27), .B(n2684), .C(net18545), .D(n2683), .Z(n2157) );
  COND2X1 U2200 ( .A(n27), .B(n2686), .C(net18545), .D(n2685), .Z(n2159) );
  COND2X1 U2201 ( .A(n27), .B(n2687), .C(net18546), .D(n2686), .Z(n2160) );
  COND2X1 U2202 ( .A(n27), .B(n2688), .C(net18546), .D(n2687), .Z(n2161) );
  COND2X1 U2203 ( .A(n27), .B(n2689), .C(net18546), .D(n2688), .Z(n2162) );
  COND2X1 U2204 ( .A(n27), .B(n2690), .C(net18546), .D(n2689), .Z(n2163) );
  COND2X1 U2215 ( .A(n27), .B(n2701), .C(net18545), .D(n2700), .Z(n2174) );
  COND2X1 U2216 ( .A(net19977), .B(n2702), .C(net18545), .D(n2701), .Z(n2175)
         );
  COND2X1 U2220 ( .A(n27), .B(n2706), .C(net18545), .D(n2705), .Z(n2179) );
  COND2X1 U2221 ( .A(net20002), .B(n2707), .C(net18545), .D(n2706), .Z(n2180)
         );
  COND2X1 U2222 ( .A(n27), .B(n2708), .C(net18545), .D(n2707), .Z(n2181) );
  COND2X1 U2223 ( .A(net19794), .B(n2709), .C(net18545), .D(n2708), .Z(n2182)
         );
  COND2X1 U2225 ( .A(net20022), .B(n2711), .C(net18545), .D(n2710), .Z(n2184)
         );
  COND2X1 U2263 ( .A(n2715), .B(n3743), .C(net16638), .D(n2714), .Z(n2188) );
  COND2X1 U2265 ( .A(n3743), .B(n2717), .C(net16638), .D(n2716), .Z(n2190) );
  COND2X1 U2266 ( .A(n3743), .B(n2718), .C(net16639), .D(n2717), .Z(n2191) );
  COND2X1 U2267 ( .A(n18), .B(n2719), .C(net16638), .D(n2718), .Z(n2192) );
  COND2X1 U2268 ( .A(n3743), .B(n2720), .C(net16639), .D(n2719), .Z(n2193) );
  COND2X1 U2269 ( .A(n18), .B(n2721), .C(net16639), .D(n2720), .Z(n2194) );
  COND2X1 U2271 ( .A(n3743), .B(n2723), .C(net16638), .D(n2722), .Z(n2196) );
  COND2X1 U2272 ( .A(n3743), .B(n2724), .C(net16638), .D(n2723), .Z(n2197) );
  COND2X1 U2273 ( .A(n18), .B(n2725), .C(net16638), .D(n2724), .Z(n2198) );
  COND2X1 U2274 ( .A(n3743), .B(n2726), .C(net16639), .D(n2725), .Z(n2199) );
  COND2X1 U2275 ( .A(n18), .B(n2727), .C(n2726), .D(net16638), .Z(n2200) );
  COND2X1 U2276 ( .A(n2728), .B(n18), .C(net16638), .D(n2727), .Z(n2201) );
  COND2X1 U2277 ( .A(n3743), .B(n2729), .C(net16639), .D(n2728), .Z(n2202) );
  COND2X1 U2278 ( .A(n18), .B(n2730), .C(net16639), .D(n2729), .Z(n2203) );
  COND2X1 U2279 ( .A(n18), .B(n2731), .C(net16638), .D(n2730), .Z(n2204) );
  COND2X1 U2280 ( .A(n18), .B(n2732), .C(net16639), .D(n2731), .Z(n2205) );
  COND2X1 U2281 ( .A(n2733), .B(n3743), .C(net16638), .D(n3043), .Z(n2206) );
  COND2X1 U2282 ( .A(n18), .B(n2734), .C(net16638), .D(n2733), .Z(n2207) );
  COND2X1 U2283 ( .A(n18), .B(n2735), .C(net16638), .D(n2734), .Z(n2208) );
  COND2X1 U2284 ( .A(n18), .B(n2736), .C(net16638), .D(n2735), .Z(n2209) );
  COND2X1 U2285 ( .A(n18), .B(n2737), .C(net16639), .D(n2736), .Z(n2210) );
  COND2X1 U2287 ( .A(net18700), .B(n2739), .C(net16638), .D(n2738), .Z(n2212)
         );
  COND2X1 U2288 ( .A(n18), .B(n2740), .C(net16638), .D(n2739), .Z(n2213) );
  COND2X1 U2291 ( .A(n18), .B(n2743), .C(net16639), .D(n2742), .Z(n2216) );
  COND2X1 U2292 ( .A(n18), .B(n2744), .C(net16638), .D(n2743), .Z(n2217) );
  COND2X1 U2293 ( .A(n2745), .B(net18700), .C(net16639), .D(n2744), .Z(n2218)
         );
  CAOR1X1 U2329 ( .A(n6), .B(n9), .C(n2747), .Z(n2220) );
  COND2X1 U2331 ( .A(n2748), .B(n6), .C(n2749), .D(n9), .Z(n2222) );
  COND2X1 U2332 ( .A(n9), .B(n2750), .C(n6), .D(n2749), .Z(n2223) );
  COND2X1 U2333 ( .A(n9), .B(n2751), .C(n6), .D(n2750), .Z(n2224) );
  COND2X1 U2334 ( .A(n9), .B(n2752), .C(n6), .D(n2751), .Z(n2225) );
  COND2X1 U2335 ( .A(n3022), .B(n3905), .C(n6), .D(n2752), .Z(n2226) );
  COND2X1 U2336 ( .A(n2754), .B(n9), .C(n6), .D(n2753), .Z(n2227) );
  COND2X1 U2337 ( .A(n9), .B(n2755), .C(n6), .D(n2754), .Z(n2228) );
  COND2X1 U2340 ( .A(n9), .B(n2758), .C(n6), .D(n2757), .Z(n2231) );
  COND2X1 U2341 ( .A(n9), .B(n2759), .C(n6), .D(n2758), .Z(n2232) );
  COND2X1 U2343 ( .A(n3905), .B(n2761), .C(n6), .D(n2760), .Z(n2234) );
  COND2X1 U2344 ( .A(n9), .B(n2762), .C(n6), .D(n2761), .Z(n2235) );
  COND2X1 U2345 ( .A(n3905), .B(n2763), .C(n6), .D(n2762), .Z(n2236) );
  COND2X1 U2349 ( .A(n9), .B(n2767), .C(n6), .D(n2766), .Z(n2240) );
  COND2X1 U2355 ( .A(n3906), .B(n2773), .C(n6), .D(n2772), .Z(n2246) );
  COND2X1 U2356 ( .A(n3906), .B(n2774), .C(n6), .D(n2773), .Z(n2247) );
  COND2X1 U2360 ( .A(n2778), .B(n3906), .C(n6), .D(n2777), .Z(n2251) );
  COND2X1 U1887 ( .A(n3044), .B(n2543), .C(net16684), .D(n2542), .Z(n2016) );
  COND2X1 U1889 ( .A(n2545), .B(n3044), .C(n3360), .D(net16684), .Z(n2018) );
  CFA1X1 U1258 ( .A(n1957), .B(n2141), .CI(n2017), .CO(n1594), .S(n1595) );
  COND2X1 U1888 ( .A(n3340), .B(n3360), .C(net16683), .D(n2543), .Z(n2017) );
  COND2X1 U1546 ( .A(n3051), .B(n3168), .C(net21572), .D(n2371), .Z(n1852) );
  CANR1X1 U188 ( .A(net18255), .B(n253), .C(n244), .Z(n242) );
  CNR2X2 U181 ( .A(n274), .B(n3127), .Z(n233) );
  COND1X1 U176 ( .A(n231), .B(net18430), .C(n232), .Z(n230) );
  COND2X1 U1808 ( .A(n2498), .B(n81), .C(net18902), .D(n2497), .Z(n1972) );
  COND2X1 U1547 ( .A(net18572), .B(n2373), .C(net21572), .D(n2372), .Z(n1853)
         );
  COND2X1 U1417 ( .A(n135), .B(n2311), .C(net18772), .D(n2310), .Z(n1796) );
  CFA1X1 U1046 ( .A(n1206), .B(n1204), .CI(n1210), .CO(n1172), .S(n1173) );
  CFA1X1 U1065 ( .A(n1853), .B(n1796), .CI(n1971), .CO(n1210), .S(n1211) );
  COND2X1 U2197 ( .A(n2682), .B(net18545), .C(n2683), .D(n27), .Z(n2156) );
  COND2X1 U1352 ( .A(n144), .B(n2280), .C(net16617), .D(n2279), .Z(n1766) );
  CFA1X1 U1047 ( .A(n2093), .B(n1212), .CI(n1185), .CO(n1174), .S(n1175) );
  CAOR1X1 U2262 ( .A(net16639), .B(n18), .C(n2714), .Z(n2187) );
  CFA1X1 U1061 ( .A(n2187), .B(n1238), .CI(n1240), .CO(n1202), .S(n1203) );
  COND2X1 U1351 ( .A(net18570), .B(n2279), .C(net16617), .D(n2278), .Z(n1765)
         );
  COND2X1 U2196 ( .A(n2682), .B(n27), .C(net18546), .D(n2681), .Z(n2155) );
  CFA1X1 U1033 ( .A(n1178), .B(n1180), .CI(n1182), .CO(n1146), .S(n1147) );
  CFA1X1 U1051 ( .A(n1765), .B(n1940), .CI(n2155), .CO(n1182), .S(n1183) );
  CFA1X1 U1041 ( .A(n1194), .B(n1167), .CI(n1169), .CO(n1162), .S(n1163) );
  CFA1X1 U1027 ( .A(n1139), .B(n1162), .CI(n1164), .CO(n1134), .S(n1135) );
  CND2X2 U333 ( .A(n359), .B(n438), .Z(n353) );
  COND1X1 U182 ( .A(n3127), .B(n275), .C(net18270), .Z(n236) );
  CND2X2 U213 ( .A(n272), .B(n736), .Z(n261) );
  CANR1X1 U214 ( .A(n736), .B(n273), .C(n264), .Z(n262) );
  COND1X1 U222 ( .A(n268), .B(net18430), .C(n269), .Z(n267) );
  CND2X1 U2507 ( .A(n1417), .B(n3543), .Z(n3544) );
  CENXL U2508 ( .A(n3994), .B(n3999), .Z(n3022) );
  CIVX3 U2509 ( .A(net19148), .Z(n3023) );
  CIVX2 U2510 ( .A(net19148), .Z(net16633) );
  CIVX2 U2511 ( .A(n3319), .Z(n3321) );
  CND2X1 U2512 ( .A(net21373), .B(n3262), .Z(net21367) );
  COND2X2 U2513 ( .A(n36), .B(n2654), .C(n3655), .D(n2653), .Z(n2127) );
  CENX1 U2514 ( .A(n2792), .B(net18486), .Z(n2429) );
  CAN2X1 U2515 ( .A(n1563), .B(n1580), .Z(n3124) );
  CNR2X1 U2516 ( .A(n3579), .B(n1562), .Z(n3596) );
  CENX2 U2517 ( .A(n3024), .B(n881), .Z(n3375) );
  CIVX20 U2518 ( .A(n883), .Z(n3024) );
  CIVXL U2519 ( .A(n3214), .Z(n3025) );
  CIVX2 U2520 ( .A(n39), .Z(n3157) );
  CENXL U2521 ( .A(n2789), .B(net18510), .Z(n3026) );
  CNIVXL U2522 ( .A(n1084), .Z(n3027) );
  CIVXL U2523 ( .A(n1227), .Z(n3028) );
  CIVX1 U2524 ( .A(n3028), .Z(n3029) );
  CENX2 U2525 ( .A(n3191), .B(net18491), .Z(net18887) );
  CIVDX4 U2526 ( .A(a[16]), .Z0(n3191) );
  CENX2 U2527 ( .A(n3989), .B(net18520), .Z(n2400) );
  CENXL U2528 ( .A(net16389), .B(n3961), .Z(n3030) );
  COND1XL U2529 ( .A(n628), .B(n622), .C(n623), .Z(n3031) );
  CENXL U2530 ( .A(n3989), .B(n3806), .Z(n3032) );
  CIVXL U2531 ( .A(n1338), .Z(n3033) );
  CIVX2 U2532 ( .A(n3033), .Z(n3034) );
  CEOX1 U2533 ( .A(n1337), .B(n1362), .Z(n3379) );
  CENXL U2534 ( .A(n2804), .B(n4011), .Z(n3035) );
  CENXL U2535 ( .A(n3995), .B(n3961), .Z(n3036) );
  CENX1 U2536 ( .A(n3997), .B(net16676), .Z(n2382) );
  CND2X2 U2537 ( .A(n3250), .B(n3251), .Z(n2346) );
  COND2X2 U2538 ( .A(n3913), .B(n2479), .C(net19422), .D(n2478), .Z(n1954) );
  CND2XL U2539 ( .A(net19446), .B(n3421), .Z(n3423) );
  COND2XL U2540 ( .A(n108), .B(n2400), .C(n3957), .D(n2399), .Z(n1878) );
  COND2XL U2541 ( .A(n3747), .B(net19695), .C(n3957), .D(n2416), .Z(n1728) );
  CIVX1 U2542 ( .A(n3957), .Z(n3478) );
  COND2X1 U2543 ( .A(n2415), .B(n3747), .C(n3957), .D(n2414), .Z(n1893) );
  CENX1 U2544 ( .A(n3993), .B(net18510), .Z(n2523) );
  CIVXL U2545 ( .A(n3935), .Z(n3037) );
  CND2XL U2546 ( .A(n1383), .B(n1381), .Z(n3547) );
  COND2X1 U2547 ( .A(n90), .B(n2461), .C(n87), .D(n2460), .Z(n3038) );
  COND2XL U2548 ( .A(n90), .B(n2461), .C(n87), .D(n2460), .Z(n1080) );
  CEOXL U2549 ( .A(n3201), .B(n4017), .Z(n2496) );
  CIVX1 U2550 ( .A(n954), .Z(n955) );
  CIVXL U2551 ( .A(n1978), .Z(n3039) );
  CIVX1 U2552 ( .A(n3039), .Z(n3040) );
  CENX1 U2553 ( .A(n3992), .B(n4015), .Z(n2590) );
  CENXL U2554 ( .A(net16393), .B(net16676), .Z(n3041) );
  CENX2 U2555 ( .A(n3990), .B(net18520), .Z(n2399) );
  CIVXL U2556 ( .A(n3166), .Z(n3042) );
  CND2XL U2557 ( .A(n1320), .B(n1297), .Z(n3497) );
  CEOX1 U2558 ( .A(n3183), .B(n1260), .Z(n1225) );
  CND2XL U2559 ( .A(n1260), .B(n1237), .Z(n3184) );
  CND2XL U2560 ( .A(n1260), .B(n1241), .Z(n3185) );
  CND2XL U2561 ( .A(n3126), .B(n1261), .Z(n3301) );
  CIVXL U2562 ( .A(n668), .Z(n667) );
  CENXL U2563 ( .A(n667), .B(n197), .Z(product[15]) );
  CENXL U2564 ( .A(n3987), .B(n4004), .Z(n3043) );
  CIVX4 U2565 ( .A(net19442), .Z(net18772) );
  CIVX2 U2566 ( .A(net18096), .Z(net16638) );
  CND2X4 U2567 ( .A(n3371), .B(net16682), .Z(n3044) );
  CND2X2 U2568 ( .A(n3371), .B(net16682), .Z(net18612) );
  CEO3XL U2569 ( .A(n1590), .B(n1573), .C(n1575), .Z(n1569) );
  CIVX3 U2570 ( .A(n3327), .Z(n3334) );
  CNIVX1 U2571 ( .A(n1787), .Z(n3045) );
  COND2X1 U2572 ( .A(n108), .B(n2397), .C(n3957), .D(n2396), .Z(n3343) );
  COND2XL U2573 ( .A(n27), .B(n2701), .C(net18545), .D(n2700), .Z(n3046) );
  CENX1 U2574 ( .A(n3986), .B(n3348), .Z(n2700) );
  CIVXL U2575 ( .A(n3167), .Z(n3047) );
  CENX2 U2576 ( .A(net19780), .B(n1145), .Z(n1139) );
  CND2X2 U2577 ( .A(n3190), .B(a[16]), .Z(n3193) );
  CIVX3 U2578 ( .A(n4017), .Z(n3190) );
  CNIVX1 U2579 ( .A(n1219), .Z(n3048) );
  CENX1 U2580 ( .A(n3795), .B(n3489), .Z(n1219) );
  CENXL U2581 ( .A(n3201), .B(n3493), .Z(n3049) );
  CIVX1 U2582 ( .A(n2793), .Z(n3201) );
  CENXL U2583 ( .A(n3572), .B(n3182), .Z(n3050) );
  CENX1 U2584 ( .A(n3572), .B(n3182), .Z(n2381) );
  CIVX2 U2585 ( .A(net15975), .Z(n3182) );
  CEOXL U2586 ( .A(net16391), .B(net16675), .Z(n3051) );
  COND2XL U2587 ( .A(n2517), .B(n3044), .C(net16684), .D(n2516), .Z(n3052) );
  COND2XL U2588 ( .A(n2517), .B(n3044), .C(net16684), .D(n2516), .Z(n1991) );
  COND2XL U2589 ( .A(n90), .B(n2468), .C(net19422), .D(n2467), .Z(n3053) );
  CENXL U2590 ( .A(n2789), .B(net18510), .Z(n2525) );
  CENXL U2591 ( .A(n2783), .B(net16023), .Z(n2552) );
  CENXL U2592 ( .A(n2806), .B(net16549), .Z(n2575) );
  CENXL U2593 ( .A(n3986), .B(net16549), .Z(n2568) );
  CENXL U2594 ( .A(n3989), .B(net16027), .Z(n2565) );
  CIVX1 U2595 ( .A(n864), .Z(n865) );
  CFA1X1 U2596 ( .A(n1866), .B(n864), .CI(n1807), .CO(n852), .S(n853) );
  COND2X1 U2597 ( .A(n3173), .B(n2356), .C(net16606), .D(n2355), .Z(n864) );
  CIVX1 U2598 ( .A(n3355), .Z(n3054) );
  CIVX1 U2599 ( .A(n3054), .Z(n3055) );
  COND2X2 U2600 ( .A(n3352), .B(n3165), .C(n3432), .D(n2584), .Z(n2058) );
  CENX2 U2601 ( .A(n2794), .B(net16645), .Z(n3864) );
  CENXL U2602 ( .A(n3921), .B(a[30]), .Z(n3056) );
  CENX1 U2603 ( .A(n3921), .B(a[30]), .Z(n3057) );
  CIVDX4 U2604 ( .A(n136), .Z0(n3921), .Z1(n3920) );
  CENX1 U2605 ( .A(n3921), .B(a[30]), .Z(n2812) );
  COND2X1 U2606 ( .A(n3336), .B(n2428), .C(n3023), .D(n2427), .Z(n1034) );
  CNR2X1 U2607 ( .A(n3908), .B(n1244), .Z(n540) );
  CND2X2 U2608 ( .A(n3918), .B(n2821), .Z(n3058) );
  CND2X2 U2609 ( .A(n3918), .B(n2821), .Z(n3059) );
  CND2X1 U2610 ( .A(n3918), .B(n2821), .Z(n3916) );
  CIVXL U2611 ( .A(n505), .Z(n3060) );
  CIVXL U2612 ( .A(n3060), .Z(n3061) );
  CENXL U2613 ( .A(n3989), .B(n3806), .Z(n2598) );
  CND2XL U2614 ( .A(n3447), .B(n3406), .Z(n3408) );
  CIVX2 U2615 ( .A(n4015), .Z(n3735) );
  CNIVXL U2616 ( .A(n1198), .Z(n3266) );
  CENX1 U2617 ( .A(net16403), .B(n4021), .Z(n2345) );
  COAN1X1 U2618 ( .A(n613), .B(n3653), .C(net19203), .Z(n3062) );
  CNIVX1 U2619 ( .A(n2206), .Z(n3063) );
  CENX1 U2620 ( .A(n3064), .B(n1636), .Z(n1619) );
  CENX1 U2621 ( .A(n1638), .B(n1634), .Z(n3064) );
  COND1XL U2622 ( .A(n287), .B(n334), .C(n3941), .Z(n3065) );
  COND1XL U2623 ( .A(n224), .B(net19414), .C(n225), .Z(n3066) );
  COAN1X1 U2624 ( .A(n327), .B(n291), .C(n292), .Z(n3941) );
  CANR1X1 U2625 ( .A(net18254), .B(n236), .C(n227), .Z(n225) );
  CENXL U2626 ( .A(n560), .B(n3067), .Z(product[30]) );
  CAN2XL U2627 ( .A(n764), .B(n3801), .Z(n3067) );
  CENXL U2628 ( .A(n569), .B(n3068), .Z(product[29]) );
  CAN2XL U2629 ( .A(n568), .B(n3781), .Z(n3068) );
  CIVX1 U2630 ( .A(n514), .Z(n516) );
  CIVXL U2631 ( .A(net19456), .Z(n3069) );
  CND2X1 U2632 ( .A(n3202), .B(n1040), .Z(n3205) );
  CND2XL U2633 ( .A(n1040), .B(n1042), .Z(n3751) );
  CNR2X1 U2634 ( .A(n671), .B(n674), .Z(n669) );
  COND1X1 U2635 ( .A(n674), .B(n676), .C(n675), .Z(n673) );
  CIVXL U2636 ( .A(n674), .Z(n781) );
  CNR2X2 U2637 ( .A(n1653), .B(n1664), .Z(n674) );
  CNIVX1 U2638 ( .A(n1223), .Z(n3795) );
  CNR2X2 U2639 ( .A(n460), .B(n444), .Z(n438) );
  CIVXL U2640 ( .A(n460), .Z(n462) );
  CNIVX2 U2641 ( .A(n2052), .Z(n3070) );
  CENX1 U2642 ( .A(n1307), .B(n3071), .Z(n1305) );
  CENX1 U2643 ( .A(n1309), .B(n1334), .Z(n3071) );
  CEO3X1 U2644 ( .A(n1019), .B(n1038), .C(n3084), .Z(n3803) );
  CND3X2 U2645 ( .A(n3583), .B(n3584), .C(n3585), .Z(n1038) );
  CAN2X2 U2646 ( .A(n3215), .B(n3216), .Z(n3153) );
  CIVX2 U2647 ( .A(a[24]), .Z(n3072) );
  CIVX4 U2648 ( .A(n3072), .Z(n3073) );
  CND2X2 U2649 ( .A(net18887), .B(n3346), .Z(n81) );
  CIVX3 U2650 ( .A(a[16]), .Z(n3074) );
  CIVX4 U2651 ( .A(n3074), .Z(n3075) );
  COND2X1 U2652 ( .A(n3353), .B(n2590), .C(n3267), .D(n2589), .Z(n2063) );
  CNIVXL U2653 ( .A(n2081), .Z(n3076) );
  CENXL U2654 ( .A(n3994), .B(n4011), .Z(n2621) );
  CENXL U2655 ( .A(n2804), .B(n4011), .Z(n2639) );
  CIVXL U2656 ( .A(n129), .Z(n3077) );
  CIVX3 U2657 ( .A(n4022), .Z(n3475) );
  CIVX4 U2658 ( .A(n4022), .Z(n4020) );
  CENX2 U2659 ( .A(a[28]), .B(n4022), .Z(net19442) );
  COND2XL U2660 ( .A(n3353), .B(n2608), .C(n3267), .D(n2607), .Z(n2081) );
  COND2XL U2661 ( .A(n3353), .B(n2611), .C(n51), .D(n2610), .Z(n2084) );
  CIVXL U2662 ( .A(n1467), .Z(n3078) );
  CIVXL U2663 ( .A(n3078), .Z(n3079) );
  CND2X2 U2664 ( .A(net18887), .B(n3346), .Z(n3080) );
  CND2X1 U2665 ( .A(n3422), .B(n3423), .Z(n3360) );
  CAN2XL U2666 ( .A(n1261), .B(n3296), .Z(n3081) );
  CAN2X2 U2667 ( .A(n1288), .B(n3295), .Z(n3082) );
  CENX1 U2668 ( .A(net16403), .B(n3166), .Z(n2543) );
  CNIVXL U2669 ( .A(n1301), .Z(n3083) );
  CND2X2 U2670 ( .A(n3128), .B(n3268), .Z(n3209) );
  CND2X2 U2671 ( .A(n1581), .B(n1596), .Z(n644) );
  CND2X2 U2672 ( .A(n1222), .B(n1197), .Z(n3892) );
  CNIVX1 U2673 ( .A(n1017), .Z(n3084) );
  COR2X1 U2674 ( .A(n3234), .B(n1014), .Z(n3419) );
  COND1X2 U2675 ( .A(n444), .B(n3161), .C(n445), .Z(net21583) );
  CEO3X1 U2676 ( .A(n1087), .B(n1108), .C(net19382), .Z(net18635) );
  COND1X2 U2677 ( .A(n573), .B(n567), .C(n568), .Z(n3162) );
  CANR1X2 U2678 ( .A(n3854), .B(n3162), .C(n550), .Z(n548) );
  CND2X2 U2679 ( .A(n1413), .B(n1436), .Z(n592) );
  CIVXL U2680 ( .A(n3214), .Z(n3085) );
  CIVX1 U2681 ( .A(n2009), .Z(n3214) );
  CND3X1 U2682 ( .A(n3649), .B(n3650), .C(n3651), .Z(n1144) );
  COND2X2 U2683 ( .A(n27), .B(n2685), .C(net18545), .D(n2684), .Z(n2158) );
  CEOX2 U2684 ( .A(n1183), .B(n1181), .Z(n3086) );
  CEOX2 U2685 ( .A(n3086), .B(n1202), .Z(n1169) );
  CND2X1 U2686 ( .A(n1202), .B(n1181), .Z(n3087) );
  CND2X1 U2687 ( .A(n1202), .B(n1183), .Z(n3088) );
  CND2XL U2688 ( .A(n1181), .B(n1183), .Z(n3089) );
  CND3X2 U2689 ( .A(n3087), .B(n3088), .C(n3089), .Z(n1168) );
  CIVX3 U2690 ( .A(n3326), .Z(n3333) );
  COND2X1 U2691 ( .A(n3705), .B(n2281), .C(net16617), .D(n2280), .Z(n1767) );
  CEOX2 U2692 ( .A(n3691), .B(n3383), .Z(n1399) );
  COND2XL U2693 ( .A(n3915), .B(n2306), .C(net18772), .D(n2305), .Z(n1791) );
  CENXL U2694 ( .A(net16399), .B(net18538), .Z(n3710) );
  CENXL U2695 ( .A(n3987), .B(net18538), .Z(n2303) );
  CENX1 U2696 ( .A(n3990), .B(net18538), .Z(n2300) );
  CENXL U2697 ( .A(n3995), .B(n3999), .Z(n2752) );
  CENXL U2698 ( .A(n3993), .B(n3999), .Z(n2754) );
  CENXL U2699 ( .A(n3994), .B(n3999), .Z(n2753) );
  CENXL U2700 ( .A(n3992), .B(n3999), .Z(n2755) );
  CENX2 U2701 ( .A(n3987), .B(net16671), .Z(n2468) );
  CND2X2 U2702 ( .A(n3816), .B(n3817), .Z(n3090) );
  CND2X2 U2703 ( .A(n3816), .B(n3817), .Z(n2821) );
  CEO3X1 U2704 ( .A(n1219), .B(n1246), .C(n3469), .Z(n3908) );
  CND2XL U2705 ( .A(net16407), .B(net18492), .Z(n3093) );
  CND2X1 U2706 ( .A(n3091), .B(n3092), .Z(n3094) );
  CND2X1 U2707 ( .A(n3093), .B(n3094), .Z(n2545) );
  CIVXL U2708 ( .A(net16407), .Z(n3091) );
  CIVXL U2709 ( .A(net18492), .Z(n3092) );
  CEOX2 U2710 ( .A(n979), .B(n996), .Z(n3095) );
  CEOX2 U2711 ( .A(n3095), .B(n977), .Z(n975) );
  CND2XL U2712 ( .A(n977), .B(n996), .Z(n3096) );
  CND2X1 U2713 ( .A(n977), .B(n979), .Z(n3097) );
  CND2XL U2714 ( .A(n996), .B(n979), .Z(n3098) );
  CND3X1 U2715 ( .A(n3096), .B(n3097), .C(n3098), .Z(n974) );
  CND3X2 U2716 ( .A(n3114), .B(n3115), .C(n3116), .Z(n996) );
  CND2X1 U2717 ( .A(n1329), .B(n1331), .Z(n3454) );
  CEN3X1 U2718 ( .A(n1046), .B(n1048), .C(n1027), .Z(n3099) );
  CEOX1 U2719 ( .A(n1074), .B(n1072), .Z(n3100) );
  CEOX1 U2720 ( .A(n3100), .B(n1051), .Z(n1047) );
  CND2X1 U2721 ( .A(n1051), .B(n1072), .Z(n3101) );
  CND2X1 U2722 ( .A(n1051), .B(n1074), .Z(n3102) );
  CND2X1 U2723 ( .A(n1072), .B(n1074), .Z(n3103) );
  CND3X2 U2724 ( .A(n3101), .B(n3102), .C(n3103), .Z(n1046) );
  CNR2X1 U2725 ( .A(n3864), .B(net18613), .Z(n3307) );
  CND2XL U2726 ( .A(n1140), .B(n3323), .Z(n3106) );
  CND2X1 U2727 ( .A(n3104), .B(n3105), .Z(n3107) );
  CND2X1 U2728 ( .A(n3106), .B(n3107), .Z(n1111) );
  CIVXL U2729 ( .A(n1140), .Z(n3104) );
  CIVX1 U2730 ( .A(n3323), .Z(n3105) );
  CND2X1 U2731 ( .A(n1109), .B(n1111), .Z(net16512) );
  CIVX2 U2732 ( .A(n3699), .Z(n1243) );
  CENXL U2733 ( .A(n2782), .B(net16023), .Z(n2551) );
  CENXL U2734 ( .A(n3992), .B(net16023), .Z(n2557) );
  CENXL U2735 ( .A(n2784), .B(net16023), .Z(n2553) );
  CENXL U2736 ( .A(n2792), .B(net16023), .Z(n2561) );
  CND2X2 U2737 ( .A(n2815), .B(n114), .Z(net18572) );
  CIVX3 U2738 ( .A(net21569), .Z(net15959) );
  CENX2 U2739 ( .A(n3108), .B(n1587), .Z(n1583) );
  CENX2 U2740 ( .A(n1589), .B(n1600), .Z(n3108) );
  CENX1 U2741 ( .A(n2794), .B(n4018), .Z(n2497) );
  CNR2X2 U2742 ( .A(n1641), .B(n1652), .Z(n671) );
  COND2X1 U2743 ( .A(n3915), .B(n2304), .C(net18772), .D(n2303), .Z(n1789) );
  CENX1 U2744 ( .A(net18510), .B(n2792), .Z(n2528) );
  CIVX1 U2745 ( .A(n369), .Z(n744) );
  CENXL U2746 ( .A(n3995), .B(n4017), .Z(n2488) );
  CND2X1 U2747 ( .A(n4015), .B(n3736), .Z(n3111) );
  CND2X2 U2748 ( .A(n3109), .B(n3110), .Z(n3112) );
  CND2X2 U2749 ( .A(n3112), .B(n3111), .Z(n2822) );
  CIVX2 U2750 ( .A(n4015), .Z(n3109) );
  CIVX1 U2751 ( .A(n3736), .Z(n3110) );
  CIVX2 U2752 ( .A(a[10]), .Z(n3736) );
  CIVXL U2753 ( .A(n1979), .Z(n3213) );
  CND2XL U2754 ( .A(n3214), .B(n1979), .Z(n3215) );
  CND2XL U2755 ( .A(n3350), .B(n1767), .Z(n3725) );
  CEOX2 U2756 ( .A(n3217), .B(n1869), .Z(n887) );
  CND2XL U2757 ( .A(n1869), .B(n1898), .Z(n3218) );
  CEOX2 U2758 ( .A(n1020), .B(n1001), .Z(n3113) );
  CEOX2 U2759 ( .A(n3113), .B(n1018), .Z(n997) );
  CND2XL U2760 ( .A(n1018), .B(n1001), .Z(n3114) );
  CND2XL U2761 ( .A(n1018), .B(n1020), .Z(n3115) );
  CND2XL U2762 ( .A(n1001), .B(n1020), .Z(n3116) );
  COR2X2 U2763 ( .A(n126), .B(n2335), .Z(n3117) );
  COR2X1 U2764 ( .A(net16623), .B(n2334), .Z(n3118) );
  CND2X2 U2765 ( .A(n3117), .B(n3118), .Z(n1818) );
  CND3X1 U2766 ( .A(n3555), .B(n3556), .C(n3557), .Z(n1020) );
  COND2XL U2767 ( .A(net18573), .B(n2291), .C(net18772), .D(n2290), .Z(n1776)
         );
  COND2XL U2768 ( .A(net18573), .B(n2302), .C(net18772), .D(n2301), .Z(n1787)
         );
  CANR1X2 U2769 ( .A(net18282), .B(n608), .C(n601), .Z(n595) );
  CND2XL U2770 ( .A(n3230), .B(n3042), .Z(n3232) );
  CND2XL U2771 ( .A(net18491), .B(net21418), .Z(n3414) );
  CIVX3 U2772 ( .A(net18491), .Z(net18492) );
  CANR1X2 U2773 ( .A(n363), .B(n397), .C(n364), .Z(n362) );
  COND2X2 U2774 ( .A(n3705), .B(n2265), .C(net16617), .D(n2264), .Z(n1751) );
  CIVX1 U2775 ( .A(net19760), .Z(net19762) );
  CENX1 U2776 ( .A(n3344), .B(net19762), .Z(n2535) );
  CIVX1 U2777 ( .A(n3744), .Z(n3645) );
  CAOR1XL U2778 ( .A(net16684), .B(n3044), .C(n2516), .Z(n1990) );
  COR2X1 U2779 ( .A(net21601), .B(n2510), .Z(n3625) );
  CNIVX4 U2780 ( .A(net15959), .Z(net18538) );
  CENXL U2781 ( .A(net16391), .B(net18538), .Z(n2306) );
  CENXL U2782 ( .A(net16399), .B(net18538), .Z(n2310) );
  CANR1X1 U2783 ( .A(n739), .B(n308), .C(n301), .Z(n299) );
  CENX4 U2784 ( .A(n3075), .B(n3167), .Z(n3285) );
  CAN2X2 U2785 ( .A(net18411), .B(net18412), .Z(net22007) );
  CNIVX4 U2786 ( .A(n2799), .Z(n3986) );
  CNIVX4 U2787 ( .A(n2798), .Z(n3987) );
  CNIVX1 U2788 ( .A(n1426), .Z(n3804) );
  COND1X1 U2789 ( .A(n392), .B(n365), .C(n366), .Z(n364) );
  COAN1XL U2790 ( .A(n369), .B(n379), .C(n370), .Z(n366) );
  CEOX1 U2791 ( .A(n1407), .B(n1405), .Z(n3562) );
  CND2X1 U2792 ( .A(n233), .B(net18254), .Z(n224) );
  CENX1 U2793 ( .A(n2808), .B(net16671), .Z(n2478) );
  CND2X1 U2794 ( .A(n3573), .B(n3574), .Z(n2414) );
  CIVX2 U2795 ( .A(n84), .Z(net16580) );
  CIVX2 U2796 ( .A(n3736), .Z(n3487) );
  COND2X1 U2797 ( .A(n27), .B(n2696), .C(net18546), .D(n2695), .Z(n2169) );
  CHA1X1 U2798 ( .A(n1727), .B(n1862), .CO(n1458), .S(n1459) );
  CIVX2 U2799 ( .A(net15999), .Z(net19319) );
  CND2X1 U2800 ( .A(n3447), .B(net21345), .Z(n3449) );
  CENX1 U2801 ( .A(net16389), .B(net16671), .Z(n2470) );
  CENX1 U2802 ( .A(n3995), .B(n3956), .Z(n2686) );
  CND2X1 U2803 ( .A(n1208), .B(n1177), .Z(n3640) );
  CND2X1 U2804 ( .A(n1208), .B(n1179), .Z(n3639) );
  CND2X1 U2805 ( .A(n1179), .B(n1177), .Z(n3641) );
  CNIVX4 U2806 ( .A(n2787), .Z(n3993) );
  CNIVX4 U2807 ( .A(n2785), .Z(n3995) );
  CNIVX4 U2808 ( .A(n2795), .Z(n3990) );
  CENX1 U2809 ( .A(n3991), .B(net18520), .Z(n2394) );
  CNIVX4 U2810 ( .A(n2805), .Z(net16399) );
  CNR2IX1 U2811 ( .B(n3998), .A(n3484), .Z(n1989) );
  CIVX1 U2812 ( .A(n3986), .Z(n3344) );
  COND2X1 U2813 ( .A(n90), .B(n2469), .C(n2468), .D(net19996), .Z(n1944) );
  CND2X1 U2814 ( .A(n1230), .B(n1207), .Z(n3440) );
  CND2X1 U2815 ( .A(n1230), .B(n1209), .Z(n3441) );
  CND2X1 U2816 ( .A(n1153), .B(n1151), .Z(n3651) );
  CND2X1 U2817 ( .A(n1176), .B(n1153), .Z(n3649) );
  COND2X1 U2818 ( .A(n2583), .B(n3912), .C(n51), .D(n2582), .Z(n2056) );
  COND2X1 U2819 ( .A(net18573), .B(n2307), .C(net18772), .D(n2306), .Z(n1792)
         );
  CND2X1 U2820 ( .A(n3679), .B(n3680), .Z(n3749) );
  CFA1X1 U2821 ( .A(n1490), .B(n1469), .CI(n1471), .CO(n1464), .S(n1465) );
  CNIVX1 U2822 ( .A(n1226), .Z(net19702) );
  CEOX1 U2823 ( .A(n3660), .B(n1075), .Z(n1069) );
  CEOX1 U2824 ( .A(n1102), .B(n1077), .Z(n3660) );
  CIVX4 U2825 ( .A(net18090), .Z(net16623) );
  CEOX1 U2826 ( .A(n3415), .B(n895), .Z(n893) );
  CNR2X1 U2827 ( .A(n3159), .B(n922), .Z(n3384) );
  CND2X1 U2828 ( .A(n1545), .B(n1562), .Z(n634) );
  CND2X1 U2829 ( .A(n3134), .B(n1386), .Z(n573) );
  CND2X1 U2830 ( .A(n3908), .B(n1244), .Z(n541) );
  CNR2X1 U2831 ( .A(n353), .B(n261), .Z(n259) );
  CANR1XL U2832 ( .A(n740), .B(n323), .C(n314), .Z(n310) );
  CND2X1 U2833 ( .A(n893), .B(n906), .Z(n392) );
  CND2X1 U2834 ( .A(n939), .B(n956), .Z(n3712) );
  CANR1XL U2835 ( .A(n779), .B(n667), .C(n664), .Z(n662) );
  CIVXL U2836 ( .A(n660), .Z(n778) );
  CANR1XL U2837 ( .A(n554), .B(n574), .C(n555), .Z(n553) );
  CAN2X2 U2838 ( .A(n3177), .B(n3178), .Z(n3119) );
  CNIVX1 U2839 ( .A(n1931), .Z(n3120) );
  COR2XL U2840 ( .A(n353), .B(n309), .Z(n3121) );
  CIVXL U2841 ( .A(net18703), .Z(net18700) );
  CENX4 U2842 ( .A(a[30]), .B(net15965), .Z(n3122) );
  CAN2X1 U2843 ( .A(n3301), .B(n3300), .Z(n3123) );
  CNIVX1 U2844 ( .A(n2172), .Z(n3125) );
  CAN2X1 U2845 ( .A(n1286), .B(n1288), .Z(n3126) );
  COR2X1 U2846 ( .A(n265), .B(n241), .Z(n3127) );
  CAN2X1 U2847 ( .A(n3273), .B(n3274), .Z(n3128) );
  CAN2XL U2848 ( .A(n1566), .B(n1553), .Z(n3129) );
  CAN2XL U2849 ( .A(n1286), .B(n3295), .Z(n3130) );
  CIVX1 U2850 ( .A(a[8]), .Z(n3235) );
  CIVX2 U2851 ( .A(n424), .Z(n749) );
  CIVX2 U2852 ( .A(a[22]), .Z(net18453) );
  CIVX1 U2853 ( .A(n708), .Z(n3925) );
  CNIVX4 U2854 ( .A(n2809), .Z(net16407) );
  CIVX2 U2855 ( .A(net16407), .Z(n3258) );
  CENXL U2856 ( .A(n629), .B(n191), .Z(product[21]) );
  CANR1X1 U2857 ( .A(n773), .B(n629), .C(n626), .Z(n624) );
  CIVXL U2858 ( .A(n3653), .Z(n629) );
  CENXL U2859 ( .A(n3131), .B(n619), .Z(product[23]) );
  CAN2XL U2860 ( .A(net19288), .B(n618), .Z(n3131) );
  COND1X1 U2861 ( .A(n585), .B(n3062), .C(n586), .Z(n584) );
  COR2X1 U2862 ( .A(net16684), .B(n2546), .Z(n3180) );
  CENX1 U2863 ( .A(n3984), .B(n3166), .Z(n2546) );
  CENXL U2864 ( .A(n3132), .B(n662), .Z(product[16]) );
  CAN2XL U2865 ( .A(n778), .B(n661), .Z(n3132) );
  CIVX1 U2866 ( .A(n683), .Z(n681) );
  CND2X1 U2867 ( .A(n780), .B(n672), .Z(n198) );
  CND2X1 U2868 ( .A(n1641), .B(n1652), .Z(n672) );
  CIVXL U2869 ( .A(n30), .Z(n3133) );
  CEO3XL U2870 ( .A(n1365), .B(n1363), .C(n1388), .Z(n3134) );
  CENXL U2871 ( .A(n657), .B(n3135), .Z(product[17]) );
  CAN2XL U2872 ( .A(n3944), .B(n656), .Z(n3135) );
  CENXL U2873 ( .A(n3136), .B(n3069), .Z(product[32]) );
  CAN2XL U2874 ( .A(n762), .B(n3865), .Z(n3136) );
  CIVX1 U2875 ( .A(n3697), .Z(n3357) );
  CIVX1 U2876 ( .A(n3697), .Z(n4006) );
  CIVX3 U2877 ( .A(n21), .Z(n3697) );
  CENXL U2878 ( .A(n3137), .B(n593), .Z(product[26]) );
  CND2XL U2879 ( .A(n768), .B(n592), .Z(n3137) );
  CIVX2 U2880 ( .A(n4002), .Z(n4001) );
  CENX1 U2881 ( .A(n3138), .B(n1443), .Z(n1439) );
  CENX1 U2882 ( .A(n1466), .B(n1464), .Z(n3138) );
  CENXL U2883 ( .A(n3139), .B(n553), .Z(product[31]) );
  CAN2XL U2884 ( .A(n552), .B(n763), .Z(n3139) );
  COND2XL U2885 ( .A(n63), .B(n2577), .C(n3037), .D(n2576), .Z(n3140) );
  COND2XL U2886 ( .A(n63), .B(n2577), .C(n3355), .D(n2576), .Z(n2050) );
  CEO3XL U2887 ( .A(n927), .B(n940), .C(n925), .Z(n3141) );
  CNIVXL U2888 ( .A(n396), .Z(n3142) );
  COAN1XL U2889 ( .A(n213), .B(net18430), .C(n214), .Z(product[63]) );
  CIVXL U2890 ( .A(n754), .Z(n3144) );
  CEOX2 U2891 ( .A(n3811), .B(n3395), .Z(n1267) );
  CNIVXL U2892 ( .A(n1827), .Z(n3145) );
  CND3XL U2893 ( .A(n3962), .B(n3963), .C(n3964), .Z(n3146) );
  CND3XL U2894 ( .A(n3962), .B(n3963), .C(n3964), .Z(n3147) );
  CANR1XL U2895 ( .A(n419), .B(n387), .C(n388), .Z(n386) );
  COND1XL U2896 ( .A(n693), .B(n697), .C(n694), .Z(n3148) );
  COND1X1 U2897 ( .A(n693), .B(n697), .C(n694), .Z(n692) );
  CIVX2 U2898 ( .A(n3305), .Z(n3294) );
  CIVXL U2899 ( .A(n3592), .Z(n3149) );
  CIVXL U2900 ( .A(n2046), .Z(n3150) );
  CIVX1 U2901 ( .A(n3150), .Z(n3151) );
  CENX1 U2902 ( .A(net19702), .B(net18867), .Z(n1195) );
  CND3X2 U2903 ( .A(n3636), .B(n3637), .C(n3638), .Z(n1160) );
  CIVX1 U2904 ( .A(net16633), .Z(n3326) );
  CIVXL U2905 ( .A(n3656), .Z(n3152) );
  CEO3X1 U2906 ( .A(n1943), .B(n1855), .C(n3145), .Z(n1269) );
  COND2X1 U2907 ( .A(n2481), .B(net22025), .C(net19996), .D(n2480), .Z(n1956)
         );
  CENX2 U2908 ( .A(n1138), .B(n1113), .Z(n3194) );
  CENX1 U2909 ( .A(n3153), .B(n2164), .Z(n1429) );
  CND3X2 U2910 ( .A(n3536), .B(n3537), .C(n3538), .Z(n1568) );
  CND2X1 U2911 ( .A(n1590), .B(n1573), .Z(n3536) );
  CND2X1 U2912 ( .A(n1419), .B(n1440), .Z(n3785) );
  CENX2 U2913 ( .A(n2784), .B(n3956), .Z(n2685) );
  CENX1 U2914 ( .A(n1262), .B(n3154), .Z(n1227) );
  CENX1 U2915 ( .A(n1233), .B(n1239), .Z(n3154) );
  CEOX1 U2916 ( .A(n3675), .B(n965), .Z(n961) );
  CEOXL U2917 ( .A(n967), .B(n982), .Z(n3675) );
  CIVX1 U2918 ( .A(n409), .Z(n748) );
  CNR2IX1 U2919 ( .B(n396), .A(n389), .Z(n387) );
  CND2X4 U2920 ( .A(n3264), .B(n3265), .Z(n114) );
  CENX1 U2921 ( .A(n3987), .B(n3348), .Z(n2699) );
  COND2X1 U2922 ( .A(n36), .B(n2652), .C(n3655), .D(n2651), .Z(n2125) );
  CENXL U2923 ( .A(n2784), .B(n4009), .Z(n2652) );
  CENX1 U2924 ( .A(n2789), .B(net16001), .Z(n2459) );
  COND1X2 U2925 ( .A(n700), .B(n702), .C(n701), .Z(n699) );
  CEN3X1 U2926 ( .A(n1191), .B(n1216), .C(n1189), .Z(n3552) );
  COND2XL U2927 ( .A(n126), .B(n2326), .C(net16623), .D(n2325), .Z(n1809) );
  CIVXL U2928 ( .A(n664), .Z(n3155) );
  CENX1 U2929 ( .A(n2793), .B(n4024), .Z(n2265) );
  CANR1X2 U2930 ( .A(n669), .B(n677), .C(n670), .Z(n668) );
  CND2X1 U2931 ( .A(n1165), .B(n1192), .Z(n3637) );
  CENX1 U2932 ( .A(n3987), .B(n4020), .Z(n2336) );
  COR2XL U2933 ( .A(n1082), .B(n3311), .Z(n3156) );
  CENXL U2934 ( .A(n3995), .B(n4021), .Z(n2323) );
  CIVX4 U2935 ( .A(n3347), .Z(n3348) );
  CANR1X1 U2936 ( .A(n621), .B(net19288), .C(n616), .Z(n614) );
  CND2X2 U2937 ( .A(net19208), .B(net19209), .Z(n2816) );
  CIVX2 U2938 ( .A(n39), .Z(n4014) );
  CEN3X2 U2939 ( .A(n1293), .B(n3083), .C(n1299), .Z(n3187) );
  COND2X1 U2940 ( .A(n90), .B(n2467), .C(net19996), .D(n2466), .Z(n1942) );
  CENXL U2941 ( .A(net16393), .B(n4018), .Z(n2505) );
  CENXL U2942 ( .A(n2792), .B(n3166), .Z(n3158) );
  CENX1 U2943 ( .A(n3989), .B(net18486), .Z(n2433) );
  CND2X1 U2944 ( .A(n1443), .B(n1466), .Z(n3256) );
  COND2XL U2945 ( .A(n3905), .B(n2771), .C(n6), .D(n2770), .Z(n2244) );
  COND2XL U2946 ( .A(n3905), .B(n2772), .C(n6), .D(n2771), .Z(n2245) );
  COND2XL U2947 ( .A(n3905), .B(n2777), .C(n6), .D(n2776), .Z(n2250) );
  COND2XL U2948 ( .A(n3905), .B(n2769), .C(n6), .D(n2768), .Z(n2242) );
  COND2XL U2949 ( .A(n3905), .B(n2776), .C(n6), .D(n2775), .Z(n2249) );
  COND2XL U2950 ( .A(n3905), .B(n2766), .C(n6), .D(n2765), .Z(n2239) );
  COND2XL U2951 ( .A(n3905), .B(n2770), .C(n6), .D(n2769), .Z(n2243) );
  COND2XL U2952 ( .A(n3905), .B(n2775), .C(n6), .D(n2774), .Z(n2248) );
  COND2XL U2953 ( .A(n3905), .B(n2768), .C(n6), .D(n2767), .Z(n2241) );
  COND2XL U2954 ( .A(n3905), .B(n2765), .C(n6), .D(n2764), .Z(n2238) );
  COND2XL U2955 ( .A(n3905), .B(n2760), .C(n6), .D(n2759), .Z(n2233) );
  COND2XL U2956 ( .A(n3905), .B(n2756), .C(n6), .D(n2755), .Z(n2229) );
  CEO3XL U2957 ( .A(n911), .B(n924), .C(n909), .Z(n3159) );
  CENX1 U2958 ( .A(net16399), .B(n3475), .Z(n2343) );
  CND2X1 U2959 ( .A(n1448), .B(n1444), .Z(n3838) );
  CNIVX2 U2960 ( .A(n2458), .Z(n3160) );
  CANR1X1 U2961 ( .A(n753), .B(n474), .C(n467), .Z(n3161) );
  CANR1X1 U2962 ( .A(n753), .B(n474), .C(n467), .Z(n461) );
  COND2XL U2963 ( .A(n3904), .B(n2645), .C(n3833), .D(n2644), .Z(n2118) );
  COND2X2 U2964 ( .A(n99), .B(n2440), .C(n3333), .D(n2439), .Z(n1917) );
  COND2X1 U2965 ( .A(n63), .B(n2575), .C(n3355), .D(n2574), .Z(n2048) );
  CIVX1 U2966 ( .A(n353), .Z(n355) );
  CNR2XL U2967 ( .A(n353), .B(n224), .Z(n222) );
  CIVXL U2968 ( .A(n992), .Z(n993) );
  CENX1 U2969 ( .A(n3990), .B(net16645), .Z(n2531) );
  CNIVX1 U2970 ( .A(n1430), .Z(n3383) );
  CND2IX4 U2971 ( .B(n3934), .A(n33), .Z(n3163) );
  CND2IX2 U2972 ( .B(n3934), .A(n33), .Z(n36) );
  CIVX1 U2973 ( .A(n2585), .Z(n3164) );
  CIVX2 U2974 ( .A(n3164), .Z(n3165) );
  CND2X2 U2975 ( .A(n2823), .B(n42), .Z(n3903) );
  CIVX3 U2976 ( .A(net18491), .Z(n3166) );
  CIVX3 U2977 ( .A(net18491), .Z(n3167) );
  CND2XL U2978 ( .A(n1972), .B(n1883), .Z(n3404) );
  CND2X2 U2979 ( .A(n114), .B(net21559), .Z(n3168) );
  CND2X1 U2980 ( .A(n114), .B(net21559), .Z(n117) );
  CND2X2 U2981 ( .A(net22015), .B(net21367), .Z(net21559) );
  CENX2 U2982 ( .A(n1061), .B(net19385), .Z(n3311) );
  CIVXL U2983 ( .A(n2191), .Z(n3169) );
  CIVXL U2984 ( .A(n3169), .Z(n3170) );
  CENX2 U2985 ( .A(a[26]), .B(net19232), .Z(n3171) );
  CENX2 U2986 ( .A(a[26]), .B(net19232), .Z(net18090) );
  CND2X2 U2987 ( .A(n2815), .B(n114), .Z(n3172) );
  CND2X2 U2988 ( .A(n2815), .B(n114), .Z(n3173) );
  CENX1 U2989 ( .A(n1473), .B(n3174), .Z(n1467) );
  CENX1 U2990 ( .A(n1494), .B(n1492), .Z(n3174) );
  CND2XL U2991 ( .A(n93), .B(a[20]), .Z(n3177) );
  CND2X1 U2992 ( .A(n3175), .B(n3176), .Z(n3178) );
  CIVXL U2993 ( .A(n93), .Z(n3175) );
  CIVX1 U2994 ( .A(a[20]), .Z(n3176) );
  CIVX2 U2995 ( .A(net16539), .Z(net19011) );
  CEOXL U2996 ( .A(n2806), .B(n4019), .Z(n2509) );
  CIVX4 U2997 ( .A(n3654), .Z(n3424) );
  CND2XL U2998 ( .A(n1147), .B(n1145), .Z(n3652) );
  CIVX2 U2999 ( .A(n3902), .Z(n3657) );
  CNIVX4 U3000 ( .A(n1248), .Z(n3483) );
  COND2X1 U3001 ( .A(n27), .B(n2703), .C(net18546), .D(n2702), .Z(n2176) );
  COR2XL U3002 ( .A(n2547), .B(net18613), .Z(n3179) );
  CND2X1 U3003 ( .A(n3179), .B(n3180), .Z(n2020) );
  CND3X1 U3004 ( .A(n3501), .B(n3502), .C(n3503), .Z(n1488) );
  CND2IXL U3005 ( .B(n3465), .A(n3181), .Z(n3897) );
  CEOXL U3006 ( .A(n2793), .B(net16645), .Z(n3181) );
  CENX4 U3007 ( .A(n3549), .B(n4008), .Z(n3832) );
  CENXL U3008 ( .A(net16389), .B(net19259), .Z(n2404) );
  CIVX3 U3009 ( .A(n4002), .Z(n4000) );
  CIVX3 U3010 ( .A(n4002), .Z(n3999) );
  CND2X1 U3011 ( .A(n1195), .B(n1197), .Z(n3891) );
  CENXL U3012 ( .A(n3987), .B(n4004), .Z(n2732) );
  CENX1 U3013 ( .A(n3996), .B(n4004), .Z(n2714) );
  CEOX2 U3014 ( .A(n1241), .B(n1237), .Z(n3183) );
  CND2XL U3015 ( .A(n1237), .B(n1241), .Z(n3186) );
  CND3X1 U3016 ( .A(n3184), .B(n3185), .C(n3186), .Z(n1224) );
  CEO3X2 U3017 ( .A(n2126), .B(net21556), .C(n1826), .Z(n1237) );
  CEO3X1 U3018 ( .A(n1201), .B(n3397), .C(n1224), .Z(n3799) );
  CENX2 U3019 ( .A(n3706), .B(n3187), .Z(n1281) );
  CIVX2 U3020 ( .A(net16539), .Z(net16549) );
  CIVX2 U3021 ( .A(net16539), .Z(net16027) );
  CND2X2 U3022 ( .A(n2819), .B(n78), .Z(n3188) );
  CND2X2 U3023 ( .A(n2819), .B(n78), .Z(n3189) );
  CND2X1 U3024 ( .A(n4017), .B(n3191), .Z(n3192) );
  CND2X2 U3025 ( .A(n3192), .B(n3193), .Z(n2819) );
  CENX2 U3026 ( .A(n3194), .B(n1136), .Z(n1109) );
  CEO3X2 U3027 ( .A(n1606), .B(n1591), .C(n1595), .Z(n1587) );
  CND2X1 U3028 ( .A(n1606), .B(n1591), .Z(n3195) );
  CND2X1 U3029 ( .A(n1606), .B(n1595), .Z(n3196) );
  CND2X1 U3030 ( .A(n1591), .B(n1595), .Z(n3197) );
  CND3X2 U3031 ( .A(n3195), .B(n3196), .C(n3197), .Z(n1586) );
  CND2XL U3032 ( .A(n1589), .B(n1600), .Z(n3198) );
  CND2XL U3033 ( .A(n1589), .B(n1587), .Z(n3199) );
  CND2XL U3034 ( .A(n1600), .B(n1587), .Z(n3200) );
  CND3X1 U3035 ( .A(n3198), .B(n3199), .C(n3200), .Z(n1582) );
  CENXL U3036 ( .A(net16389), .B(n4009), .Z(n2668) );
  CND2X2 U3037 ( .A(n3943), .B(n749), .Z(n416) );
  CEOX2 U3038 ( .A(n3450), .B(n1327), .Z(n1317) );
  CND2IX1 U3039 ( .B(net19034), .A(net19035), .Z(n3807) );
  CENX1 U3040 ( .A(n3990), .B(n4020), .Z(n2333) );
  CND3X1 U3041 ( .A(net18843), .B(net18844), .C(n3866), .Z(n1058) );
  CND2X1 U3042 ( .A(n3749), .B(n3203), .Z(n3204) );
  CND2X2 U3043 ( .A(n3204), .B(n3205), .Z(n1017) );
  CIVX2 U3044 ( .A(n3749), .Z(n3202) );
  CIVXL U3045 ( .A(n1040), .Z(n3203) );
  CEOX2 U3046 ( .A(n1432), .B(n1428), .Z(n3691) );
  CFA1X1 U3047 ( .A(n2040), .B(n2226), .CI(n1861), .CO(n1432), .S(n1433) );
  CNIVXL U3048 ( .A(n417), .Z(n3206) );
  CANR1X2 U3049 ( .A(n432), .B(n749), .C(n3711), .Z(n417) );
  CIVXL U3050 ( .A(n485), .Z(n3207) );
  CIVXL U3051 ( .A(n3207), .Z(n3208) );
  CND3X2 U3052 ( .A(n3965), .B(n3967), .C(n3966), .Z(n1256) );
  CIVX1 U3053 ( .A(n3348), .Z(n3857) );
  CNIVX1 U3054 ( .A(n30), .Z(n3700) );
  CIVX3 U3055 ( .A(net19927), .Z(net19422) );
  CIVX2 U3056 ( .A(net21569), .Z(net18408) );
  CIVX1 U3057 ( .A(n1009), .Z(n3592) );
  CND2XL U3058 ( .A(net19619), .B(n3607), .Z(n3397) );
  CND2X2 U3059 ( .A(n2820), .B(n3465), .Z(net18613) );
  CND2X2 U3060 ( .A(n3737), .B(n3738), .Z(n3210) );
  CND3XL U3061 ( .A(n3613), .B(n3612), .C(n3614), .Z(n3211) );
  CIVXL U3062 ( .A(n4016), .Z(n3212) );
  CND2X1 U3063 ( .A(n3737), .B(n3738), .Z(n3860) );
  COND2XL U3064 ( .A(n3189), .B(n2487), .C(n3285), .D(n2486), .Z(n1962) );
  CAOR1XL U3065 ( .A(n3285), .B(n3188), .C(n2483), .Z(n1958) );
  CENX1 U3066 ( .A(n1101), .B(n1118), .Z(n3744) );
  CND3X1 U3067 ( .A(n3608), .B(n3609), .C(n3610), .Z(n1118) );
  CNIVX1 U3068 ( .A(net18887), .Z(net21576) );
  CIVXL U3069 ( .A(n4014), .Z(n3559) );
  CIVX2 U3070 ( .A(n4014), .Z(n4011) );
  CIVX3 U3071 ( .A(n3681), .Z(n3733) );
  CEOX2 U3072 ( .A(n3375), .B(n894), .Z(n879) );
  CND2XL U3073 ( .A(n1251), .B(n1278), .Z(n3823) );
  CIVX4 U3074 ( .A(n3171), .Z(net16621) );
  CND2X1 U3075 ( .A(n3213), .B(n2009), .Z(n3216) );
  CEOX2 U3076 ( .A(n1751), .B(n1898), .Z(n3217) );
  CND2XL U3077 ( .A(n1869), .B(n1751), .Z(n3219) );
  CND2XL U3078 ( .A(n1898), .B(n1751), .Z(n3220) );
  CND3XL U3079 ( .A(n3218), .B(n3219), .C(n3220), .Z(n886) );
  CENX1 U3080 ( .A(n3989), .B(n3348), .Z(n2697) );
  CEO3X1 U3081 ( .A(n1322), .B(n1324), .C(n1326), .Z(n3221) );
  CENX1 U3082 ( .A(n3222), .B(n969), .Z(n965) );
  CENX1 U3083 ( .A(n986), .B(n988), .Z(n3222) );
  CND2X1 U3084 ( .A(n3221), .B(n3224), .Z(n3225) );
  CND2X2 U3085 ( .A(n3223), .B(n1314), .Z(n3226) );
  CND2X2 U3086 ( .A(n3225), .B(n3226), .Z(n3706) );
  CIVX2 U3087 ( .A(n1289), .Z(n3223) );
  CIVX2 U3088 ( .A(n1314), .Z(n3224) );
  CEO3X2 U3089 ( .A(n1342), .B(n1319), .C(n1317), .Z(n1311) );
  CND2X1 U3090 ( .A(n1342), .B(n1317), .Z(n3227) );
  CND2XL U3091 ( .A(n1342), .B(n1319), .Z(n3228) );
  CND2X1 U3092 ( .A(n1317), .B(n1319), .Z(n3229) );
  CND3X2 U3093 ( .A(n3227), .B(n3228), .C(n3229), .Z(n1310) );
  CIVX2 U3094 ( .A(n1109), .Z(net18751) );
  CND2XL U3095 ( .A(n2791), .B(net18510), .Z(n3231) );
  CND2X1 U3096 ( .A(n3231), .B(n3232), .Z(n2527) );
  CIVXL U3097 ( .A(n2791), .Z(n3230) );
  CENXL U3098 ( .A(n2784), .B(net18486), .Z(n2421) );
  CENXL U3099 ( .A(n2789), .B(net18486), .Z(n2426) );
  CENX1 U3100 ( .A(n3987), .B(net18486), .Z(n2435) );
  CENXL U3101 ( .A(n1491), .B(n1508), .Z(n3233) );
  CEO3XL U3102 ( .A(n999), .B(n997), .C(n1016), .Z(n3234) );
  CND3X2 U3103 ( .A(n3848), .B(n3849), .C(n3850), .Z(n1396) );
  CENX1 U3104 ( .A(n2783), .B(n4004), .Z(n2717) );
  CND2X1 U3105 ( .A(a[8]), .B(n3700), .Z(n3237) );
  CND2X2 U3106 ( .A(n3235), .B(n3236), .Z(n3238) );
  CND2X4 U3107 ( .A(n3237), .B(n3238), .Z(n42) );
  CIVX2 U3108 ( .A(n3700), .Z(n3236) );
  CND2X4 U3109 ( .A(n2823), .B(n42), .Z(n3904) );
  CEOX2 U3110 ( .A(n1055), .B(n1053), .Z(n3239) );
  CEOX2 U3111 ( .A(n1057), .B(n3239), .Z(n1045) );
  CND2X1 U3112 ( .A(n1057), .B(n1053), .Z(n3240) );
  CND2XL U3113 ( .A(n1057), .B(n1055), .Z(n3241) );
  CND2XL U3114 ( .A(n1053), .B(n1055), .Z(n3242) );
  CND3X1 U3115 ( .A(n3240), .B(n3241), .C(n3242), .Z(n1044) );
  CEO3X2 U3116 ( .A(n1242), .B(n2156), .C(n1766), .Z(n1213) );
  CND2XL U3117 ( .A(n1242), .B(n1766), .Z(n3243) );
  CND2XL U3118 ( .A(n1242), .B(n2156), .Z(n3244) );
  CND2XL U3119 ( .A(n1766), .B(n2156), .Z(n3245) );
  CND3X1 U3120 ( .A(n3243), .B(n3244), .C(n3245), .Z(n1212) );
  CENXL U3121 ( .A(n2793), .B(net16645), .Z(n3246) );
  CENXL U3122 ( .A(n2793), .B(net16645), .Z(n3247) );
  CENX1 U3123 ( .A(n2808), .B(n4024), .Z(n2280) );
  CANR1X1 U3124 ( .A(n3854), .B(n3162), .C(n550), .Z(net19491) );
  CND2XL U3125 ( .A(n4021), .B(n2808), .Z(n3250) );
  CND2X1 U3126 ( .A(n3248), .B(n3249), .Z(n3251) );
  CIVXL U3127 ( .A(n2808), .Z(n3248) );
  CIVXL U3128 ( .A(n4021), .Z(n3249) );
  CAOR1XL U3129 ( .A(net16623), .B(n3682), .C(n2318), .Z(n1803) );
  CEOX1 U3130 ( .A(n2808), .B(net16675), .Z(n2379) );
  CEO3X2 U3131 ( .A(n1842), .B(n3052), .C(n1755), .Z(n953) );
  CND2XL U3132 ( .A(n1842), .B(n1755), .Z(n3252) );
  CND2XL U3133 ( .A(n1991), .B(n1842), .Z(n3253) );
  CND2XL U3134 ( .A(n1755), .B(n1991), .Z(n3254) );
  CND3X1 U3135 ( .A(n3252), .B(n3253), .C(n3254), .Z(n952) );
  COND2XL U3136 ( .A(net18572), .B(n2362), .C(n2361), .D(net21572), .Z(n1842)
         );
  CND2XL U3137 ( .A(n1464), .B(n1443), .Z(n3255) );
  CND2XL U3138 ( .A(n1464), .B(n1466), .Z(n3257) );
  CND3X1 U3139 ( .A(n3255), .B(n3256), .C(n3257), .Z(n1438) );
  CND2XL U3140 ( .A(net16407), .B(net18516), .Z(n3260) );
  CND2X1 U3141 ( .A(n3258), .B(n3259), .Z(n3261) );
  CND2X1 U3142 ( .A(n3260), .B(n3261), .Z(n2413) );
  CIVXL U3143 ( .A(net18516), .Z(n3259) );
  CND3X1 U3144 ( .A(n3515), .B(n3516), .C(n3517), .Z(n1466) );
  CENX1 U3145 ( .A(n3994), .B(n4008), .Z(n2654) );
  CENXL U3146 ( .A(n584), .B(n185), .Z(product[27]) );
  CND2X2 U3147 ( .A(n2820), .B(n3465), .Z(n3340) );
  CND3X2 U3148 ( .A(n3567), .B(n3568), .C(n3569), .Z(n1604) );
  CND2X1 U3149 ( .A(n1611), .B(n2142), .Z(n3567) );
  CND2X1 U3150 ( .A(a[24]), .B(net19259), .Z(n3264) );
  CND2X2 U3151 ( .A(n3262), .B(n3263), .Z(n3265) );
  CIVX2 U3152 ( .A(a[24]), .Z(n3262) );
  CIVX2 U3153 ( .A(net19259), .Z(n3263) );
  CND2X2 U3154 ( .A(n3719), .B(n3720), .Z(n3420) );
  CND2X1 U3155 ( .A(n1611), .B(n2173), .Z(n3568) );
  CIVX3 U3156 ( .A(n3681), .Z(n3267) );
  CND2X2 U3157 ( .A(n3269), .B(n3270), .Z(n1546) );
  CIVX1 U3158 ( .A(n1553), .Z(n3271) );
  CIVXL U3159 ( .A(n1566), .Z(n3272) );
  CND2XL U3160 ( .A(n3272), .B(n3283), .Z(n3274) );
  CND2X1 U3161 ( .A(n3272), .B(n3276), .Z(n3275) );
  CND2X1 U3162 ( .A(n1551), .B(n3129), .Z(n3277) );
  CND2XL U3163 ( .A(n1553), .B(n1551), .Z(n3278) );
  CND2XL U3164 ( .A(n1566), .B(n1551), .Z(n3279) );
  CND2XL U3165 ( .A(n1566), .B(n1553), .Z(n3269) );
  CND2XL U3166 ( .A(n1551), .B(n3271), .Z(n3280) );
  CIVX1 U3167 ( .A(n3280), .Z(n3276) );
  CND2X1 U3168 ( .A(n3275), .B(n3277), .Z(n3281) );
  CIVX2 U3169 ( .A(n3281), .Z(n3268) );
  CND2X1 U3170 ( .A(n3278), .B(n3279), .Z(n3282) );
  CIVX2 U3171 ( .A(n3282), .Z(n3270) );
  CNR2XL U3172 ( .A(n3271), .B(n1551), .Z(n3283) );
  CAN2XL U3173 ( .A(n1566), .B(n3271), .Z(n3284) );
  CND2IX1 U3174 ( .B(n1551), .A(n3284), .Z(n3273) );
  CND2XL U3175 ( .A(n1391), .B(n1414), .Z(n3979) );
  CND3X2 U3176 ( .A(n3621), .B(n3622), .C(n3623), .Z(n1462) );
  CND2X1 U3177 ( .A(n3079), .B(n1486), .Z(n3623) );
  CND2X1 U3178 ( .A(n3572), .B(net19695), .Z(n3574) );
  CND2XL U3179 ( .A(n1043), .B(n1062), .Z(n3585) );
  CND2X1 U3180 ( .A(n1064), .B(n1062), .Z(n3584) );
  CIVX2 U3181 ( .A(n3328), .Z(n3325) );
  CIVX1 U3182 ( .A(n3984), .Z(n3572) );
  CENX2 U3183 ( .A(n3075), .B(n3166), .Z(net18902) );
  CENX1 U3184 ( .A(n3606), .B(n3286), .Z(n1033) );
  CENX1 U3185 ( .A(n2056), .B(n3343), .Z(n3286) );
  CND2XL U3186 ( .A(n482), .B(n498), .Z(n3287) );
  CND2IX1 U3187 ( .B(a[16]), .A(net19446), .Z(n3361) );
  CND2X2 U3188 ( .A(n3288), .B(n3289), .Z(n1876) );
  CIVX1 U3189 ( .A(n2397), .Z(n3290) );
  CIVX1 U3190 ( .A(n3957), .Z(n3291) );
  CND2X1 U3191 ( .A(n3290), .B(n3291), .Z(n3288) );
  CND2X1 U3192 ( .A(n2816), .B(n3292), .Z(n3289) );
  CNR2IX2 U3193 ( .B(n3958), .A(n2398), .Z(n3292) );
  CENX2 U3194 ( .A(n2794), .B(net18520), .Z(n2398) );
  CNR2XL U3195 ( .A(n1627), .B(n1640), .Z(n665) );
  CIVX2 U3196 ( .A(n468), .Z(n753) );
  CIVX2 U3197 ( .A(n469), .Z(n467) );
  CND2X4 U3198 ( .A(n3420), .B(n87), .Z(n90) );
  CND2X4 U3199 ( .A(n2818), .B(n87), .Z(net22025) );
  CND2X2 U3200 ( .A(n1190), .B(n1192), .Z(n3638) );
  CIVX2 U3201 ( .A(net19384), .Z(net19617) );
  CIVXL U3202 ( .A(n573), .Z(n571) );
  CNR2IX1 U3203 ( .B(n561), .A(n3899), .Z(n554) );
  CENX1 U3204 ( .A(n1064), .B(n1043), .Z(n3362) );
  COND1X1 U3205 ( .A(n675), .B(n671), .C(n672), .Z(n670) );
  CIVXL U3206 ( .A(n671), .Z(n780) );
  COND2X1 U3207 ( .A(n3030), .B(n3353), .C(n51), .D(n2601), .Z(n2075) );
  CND2IX2 U3208 ( .B(n3191), .A(net18510), .Z(net19447) );
  CENX1 U3209 ( .A(n2791), .B(n3999), .Z(n2758) );
  CIVXL U3210 ( .A(n677), .Z(n676) );
  CENX2 U3211 ( .A(n2791), .B(net18485), .Z(n2428) );
  CENX1 U3212 ( .A(net16403), .B(net18408), .Z(n2312) );
  CND2X2 U3213 ( .A(n3293), .B(n3123), .Z(n1253) );
  CIVX1 U3214 ( .A(n1261), .Z(n3295) );
  CIVX1 U3215 ( .A(n1288), .Z(n3296) );
  CIVXL U3216 ( .A(n1286), .Z(n3297) );
  CND2X1 U3217 ( .A(n3296), .B(n3130), .Z(n3298) );
  CND2X1 U3218 ( .A(n3297), .B(n3082), .Z(n3299) );
  CND2X1 U3219 ( .A(n3297), .B(n3081), .Z(n3300) );
  CND2XL U3220 ( .A(n1288), .B(n1261), .Z(n3302) );
  CND2X1 U3221 ( .A(n1286), .B(n1261), .Z(n3303) );
  CND2X1 U3222 ( .A(n3298), .B(n3299), .Z(n3304) );
  CIVX2 U3223 ( .A(n3304), .Z(n3293) );
  CND2X1 U3224 ( .A(n3302), .B(n3303), .Z(n3305) );
  CND2IX2 U3225 ( .B(n3126), .A(n3294), .Z(n1252) );
  CIVX1 U3226 ( .A(n3308), .Z(n481) );
  CEOX2 U3227 ( .A(n3989), .B(n3635), .Z(n2730) );
  CND3X1 U3228 ( .A(n3764), .B(n3765), .C(n3766), .Z(n1504) );
  COND1XL U3229 ( .A(n3384), .B(n410), .C(n403), .Z(n3306) );
  COND1X1 U3230 ( .A(n410), .B(n3384), .C(n403), .Z(n397) );
  CIVXL U3231 ( .A(n410), .Z(n408) );
  CIVXL U3232 ( .A(n594), .Z(n596) );
  CND2IX1 U3233 ( .B(n3307), .A(n3897), .Z(n2003) );
  CENX1 U3234 ( .A(n3988), .B(n3476), .Z(n2335) );
  CNIVX4 U3235 ( .A(n2797), .Z(n3988) );
  CND2XL U3236 ( .A(net18411), .B(net18412), .Z(n3308) );
  CIVX2 U3237 ( .A(n483), .Z(net18412) );
  CENXL U3238 ( .A(n267), .B(n154), .Z(product[58]) );
  CANR1X1 U3239 ( .A(n272), .B(n356), .C(n273), .Z(n269) );
  CIVX1 U3240 ( .A(n275), .Z(n273) );
  CIVX2 U3241 ( .A(n3310), .Z(n356) );
  CANR1X1 U3242 ( .A(n359), .B(n439), .C(n360), .Z(n3310) );
  CIVX2 U3243 ( .A(n274), .Z(n272) );
  CND2XL U3244 ( .A(n355), .B(n272), .Z(n268) );
  CANR1X2 U3245 ( .A(net19938), .B(net19456), .C(n479), .Z(net18430) );
  COND1X1 U3246 ( .A(n480), .B(n515), .C(n481), .Z(n479) );
  COND1X1 U3247 ( .A(n494), .B(n484), .C(n485), .Z(n483) );
  CND2XL U3248 ( .A(net18635), .B(n1106), .Z(n494) );
  CANR1X1 U3249 ( .A(n520), .B(n535), .C(n3309), .Z(n515) );
  COND1X1 U3250 ( .A(n530), .B(n522), .C(net19253), .Z(n3309) );
  COND1X1 U3251 ( .A(n547), .B(n575), .C(n548), .Z(net19456) );
  CNR2X1 U3252 ( .A(n514), .B(n480), .Z(net19938) );
  CANR1X2 U3253 ( .A(net18264), .B(n286), .C(n277), .Z(n275) );
  CIVX2 U3254 ( .A(n279), .Z(n277) );
  CNR2X2 U3255 ( .A(n361), .B(n416), .Z(n359) );
  CANR1X1 U3256 ( .A(n359), .B(n439), .C(n360), .Z(net19414) );
  CANR1X1 U3257 ( .A(n359), .B(net21583), .C(net19415), .Z(n354) );
  CND2XL U3258 ( .A(n736), .B(n266), .Z(n154) );
  CIVX2 U3259 ( .A(n265), .Z(n736) );
  CND2X1 U3260 ( .A(n806), .B(n803), .Z(n266) );
  CIVX1 U3261 ( .A(n266), .Z(n264) );
  COAN1XL U3262 ( .A(n266), .B(n241), .C(n242), .Z(net18270) );
  CNR2X1 U3263 ( .A(n806), .B(n803), .Z(n265) );
  CND2X2 U3264 ( .A(net18752), .B(net18753), .Z(n1107) );
  CND2X1 U3265 ( .A(n1107), .B(net19299), .Z(n505) );
  CNR2X1 U3266 ( .A(n1107), .B(n1132), .Z(net18380) );
  CNR2X1 U3267 ( .A(net19300), .B(n1107), .Z(net18745) );
  CND2X2 U3268 ( .A(net18750), .B(net18751), .Z(net18753) );
  CIVX1 U3269 ( .A(net18278), .Z(net18750) );
  CND2X1 U3270 ( .A(net18278), .B(n1109), .Z(net18752) );
  CND2XL U3271 ( .A(n1109), .B(net19249), .Z(net16511) );
  CENX1 U3272 ( .A(n1111), .B(n1134), .Z(net18278) );
  CND2X1 U3273 ( .A(n1136), .B(n1138), .Z(net19521) );
  CND2X1 U3274 ( .A(n1136), .B(n1113), .Z(net19520) );
  CND2XL U3275 ( .A(n1113), .B(n1138), .Z(net19522) );
  CND2XL U3276 ( .A(net19249), .B(n1111), .Z(net16513) );
  CIVXL U3277 ( .A(n1134), .Z(net19248) );
  CND2X1 U3278 ( .A(n482), .B(n499), .Z(net18411) );
  CNR2X1 U3279 ( .A(n484), .B(n491), .Z(n482) );
  CND2X1 U3280 ( .A(n482), .B(n498), .Z(n480) );
  CNR2X1 U3281 ( .A(net18635), .B(n1106), .Z(n491) );
  COND1X1 U3282 ( .A(n512), .B(net18380), .C(n505), .Z(n499) );
  CIVXL U3283 ( .A(n499), .Z(n501) );
  CND3XL U3284 ( .A(net16578), .B(net16579), .C(net16577), .Z(n1132) );
  CND2XL U3285 ( .A(net18635), .B(n1106), .Z(net18783) );
  CNR2XL U3286 ( .A(n1083), .B(n1106), .Z(net18617) );
  CIVXL U3287 ( .A(n512), .Z(n510) );
  CND3XL U3288 ( .A(net16577), .B(net16578), .C(net16579), .Z(net19300) );
  CND3XL U3289 ( .A(net16577), .B(net16579), .C(net16578), .Z(net19299) );
  CENX1 U3290 ( .A(net18276), .B(n1135), .Z(n1133) );
  CND2XL U3291 ( .A(n1135), .B(n1137), .Z(net16578) );
  CND2XL U3292 ( .A(n1135), .B(n1160), .Z(net16577) );
  CENX1 U3293 ( .A(n1147), .B(n1168), .Z(net19780) );
  CEO3X2 U3294 ( .A(n1163), .B(n1188), .C(n1161), .Z(net18607) );
  CIVX1 U3295 ( .A(n1163), .Z(net19034) );
  CND2XL U3296 ( .A(n1188), .B(n1163), .Z(net19026) );
  CND2XL U3297 ( .A(n1161), .B(n1163), .Z(net19025) );
  CND2XL U3298 ( .A(n1168), .B(n1145), .Z(net19538) );
  CND2XL U3299 ( .A(n1147), .B(n1168), .Z(net19536) );
  CNIVX4 U3300 ( .A(net16593), .Z(net18546) );
  COND2X1 U3301 ( .A(n2465), .B(net22025), .C(net19422), .D(n2464), .Z(n1940)
         );
  CIVX8 U3302 ( .A(n3122), .Z(net16617) );
  CIVX2 U3303 ( .A(n129), .Z(net15965) );
  CIVXL U3304 ( .A(net15965), .Z(net22026) );
  CENX1 U3305 ( .A(n1228), .B(n1203), .Z(net18867) );
  CND2X1 U3306 ( .A(n1226), .B(n1203), .Z(net18830) );
  CND2X1 U3307 ( .A(n1228), .B(n1203), .Z(net18832) );
  CIVX2 U3308 ( .A(net18096), .Z(net16639) );
  CNR2X2 U3309 ( .A(n3311), .B(n1082), .Z(n484) );
  CND2X1 U3310 ( .A(n3311), .B(n3211), .Z(n485) );
  CND2X1 U3311 ( .A(n3156), .B(n3208), .Z(n173) );
  CND3X1 U3312 ( .A(net16511), .B(net16512), .C(net16513), .Z(n1106) );
  CIVXL U3313 ( .A(net19248), .Z(net19249) );
  CND2X1 U3314 ( .A(n1061), .B(n1063), .Z(net18844) );
  CND2XL U3315 ( .A(n3027), .B(n1061), .Z(net18843) );
  CEO3X1 U3316 ( .A(n1200), .B(n1198), .C(n1175), .Z(n1167) );
  CND3X1 U3317 ( .A(n3313), .B(n3314), .C(n3315), .Z(n1200) );
  CIVXL U3318 ( .A(n1200), .Z(net19753) );
  CND2X1 U3319 ( .A(n1232), .B(n1234), .Z(n3315) );
  CND2X1 U3320 ( .A(n1236), .B(n1234), .Z(n3314) );
  CND2XL U3321 ( .A(n1232), .B(n1236), .Z(n3313) );
  CND3X2 U3322 ( .A(net18962), .B(n3312), .C(net18964), .Z(n1198) );
  CND2XL U3323 ( .A(n3266), .B(net19754), .Z(net18951) );
  CND2XL U3324 ( .A(n3266), .B(n1175), .Z(net18953) );
  CND2X1 U3325 ( .A(n1211), .B(n1205), .Z(net18964) );
  CND2X1 U3326 ( .A(n1213), .B(n1205), .Z(n3312) );
  CND2X1 U3327 ( .A(n1211), .B(n1213), .Z(net18962) );
  CND2X1 U3328 ( .A(n1174), .B(n1172), .Z(net18983) );
  CND2XL U3329 ( .A(n1174), .B(n1170), .Z(net18982) );
  CEO3X2 U3330 ( .A(n1174), .B(n1170), .C(n1172), .Z(n1141) );
  CND2XL U3331 ( .A(net19754), .B(n1175), .Z(net18952) );
  CIVXL U3332 ( .A(n1184), .Z(n1185) );
  CENX1 U3333 ( .A(n1213), .B(n1211), .Z(net19384) );
  COND2X1 U3334 ( .A(n3188), .B(n2497), .C(n3316), .D(n2496), .Z(n1971) );
  CND2X1 U3335 ( .A(net19447), .B(net19448), .Z(n3316) );
  CNIVX2 U3336 ( .A(net15959), .Z(net18537) );
  CND2IX1 U3337 ( .B(net15959), .A(a[28]), .Z(net18811) );
  CIVX2 U3338 ( .A(n129), .Z(net21569) );
  CIVX1 U3339 ( .A(n3077), .Z(net15963) );
  CIVX1 U3340 ( .A(net21569), .Z(net18407) );
  CENXL U3341 ( .A(n2806), .B(net18408), .Z(n2311) );
  CEO3X2 U3342 ( .A(n2094), .B(n1941), .C(n2125), .Z(n1205) );
  CIVXL U3343 ( .A(n1205), .Z(net19618) );
  CND2X1 U3344 ( .A(net19384), .B(n1205), .Z(net19619) );
  COND2X1 U3345 ( .A(n3049), .B(n3189), .C(net21576), .D(n2495), .Z(n1184) );
  CND2X1 U3346 ( .A(net19447), .B(net19448), .Z(net21601) );
  CND2XL U3347 ( .A(n1160), .B(n1137), .Z(net16579) );
  CENX1 U3348 ( .A(n1137), .B(n1160), .Z(net18276) );
  CND2X2 U3349 ( .A(n3317), .B(n3318), .Z(n78) );
  CND2X1 U3350 ( .A(n3191), .B(net19762), .Z(n3318) );
  COR2XL U3351 ( .A(net18613), .B(n3047), .Z(net19162) );
  CIVXL U3352 ( .A(net16021), .Z(net19760) );
  CND2X1 U3353 ( .A(a[16]), .B(net19760), .Z(n3317) );
  CIVX2 U3354 ( .A(n66), .Z(net16021) );
  CENXL U3355 ( .A(n230), .B(n151), .Z(product[61]) );
  CANR1X1 U3356 ( .A(n233), .B(n356), .C(n236), .Z(n232) );
  CND2XL U3357 ( .A(n355), .B(n233), .Z(n231) );
  CIVX2 U3358 ( .A(n246), .Z(n244) );
  CIVX2 U3359 ( .A(n255), .Z(n253) );
  CANR1XL U3360 ( .A(n735), .B(n260), .C(n253), .Z(n249) );
  CND2X1 U3361 ( .A(n1158), .B(n1133), .Z(n512) );
  CNR2X1 U3362 ( .A(n1158), .B(n1133), .Z(n511) );
  CND2X2 U3363 ( .A(net21367), .B(n3322), .Z(n2815) );
  CND2X2 U3364 ( .A(net16675), .B(n3073), .Z(n3322) );
  CND2X1 U3365 ( .A(n3321), .B(a[24]), .Z(net22015) );
  CIVX4 U3366 ( .A(n3320), .Z(n3319) );
  CIVX8 U3367 ( .A(n3319), .Z(net16675) );
  CIVX2 U3368 ( .A(n111), .Z(n3320) );
  CIVX1 U3369 ( .A(net19207), .Z(net19259) );
  CIVXL U3370 ( .A(n102), .Z(net19207) );
  CND2IXL U3371 ( .B(net18453), .A(net19207), .Z(net19208) );
  CIVXL U3372 ( .A(net19232), .Z(net21373) );
  CIVX4 U3373 ( .A(n111), .Z(net19232) );
  CIVX3 U3374 ( .A(net19232), .Z(net15975) );
  CIVX1 U3375 ( .A(net19232), .Z(net15979) );
  CIVX2 U3376 ( .A(n102), .Z(net15989) );
  CND2XL U3377 ( .A(n102), .B(net18453), .Z(net19209) );
  CND2X1 U3378 ( .A(net18254), .B(n229), .Z(n151) );
  COR2X1 U3379 ( .A(n796), .B(n795), .Z(net18254) );
  CIVX2 U3380 ( .A(n794), .Z(n795) );
  CND2X1 U3381 ( .A(n796), .B(n795), .Z(n229) );
  CIVX2 U3382 ( .A(n229), .Z(n227) );
  CENXL U3383 ( .A(n1117), .B(n1115), .Z(n3323) );
  CNR2X2 U3384 ( .A(net19953), .B(n529), .Z(n520) );
  CENX1 U3385 ( .A(net16393), .B(net16676), .Z(n2373) );
  COND2X1 U3386 ( .A(n117), .B(n2374), .C(net16606), .D(n3041), .Z(n1854) );
  CIVX8 U3387 ( .A(net16675), .Z(net16676) );
  CEOX1 U3388 ( .A(net16391), .B(n3321), .Z(n2372) );
  CENXL U3389 ( .A(n3258), .B(net16675), .Z(n2380) );
  CNIVX4 U3390 ( .A(n2802), .Z(net16393) );
  CENX2 U3391 ( .A(n3073), .B(net18516), .Z(net21572) );
  CNIVX4 U3392 ( .A(net19048), .Z(net18516) );
  CENX2 U3393 ( .A(n3073), .B(net18516), .Z(net16606) );
  CIVX2 U3394 ( .A(net15989), .Z(net19048) );
  CNIVX4 U3395 ( .A(net19048), .Z(net19890) );
  CNIVX4 U3396 ( .A(net19048), .Z(net18944) );
  CIVX2 U3397 ( .A(net15989), .Z(net15985) );
  CNIVX4 U3398 ( .A(n2801), .Z(net16391) );
  CAOR1XL U3399 ( .A(n3055), .B(n3058), .C(n2549), .Z(n2022) );
  CND2X2 U3400 ( .A(n2818), .B(n87), .Z(n3913) );
  CND2X2 U3401 ( .A(n2826), .B(net16637), .Z(n3743) );
  COND1X1 U3402 ( .A(n547), .B(n575), .C(net19491), .Z(n3324) );
  CEO3X2 U3403 ( .A(n1453), .B(n1455), .C(n1457), .Z(n1445) );
  CIVX2 U3404 ( .A(net18096), .Z(net16637) );
  CND2X1 U3405 ( .A(n1325), .B(n1323), .Z(n3770) );
  COND1X1 U3406 ( .A(n540), .B(n544), .C(n541), .Z(n535) );
  COND2X1 U3407 ( .A(n3044), .B(n2533), .C(net16684), .D(n2532), .Z(n2006) );
  CIVX2 U3408 ( .A(n93), .Z(net21614) );
  CND2X2 U3409 ( .A(net16633), .B(n3119), .Z(n3336) );
  CIVX4 U3410 ( .A(n3325), .Z(net16649) );
  CND2XL U3411 ( .A(n93), .B(a[22]), .Z(net18455) );
  CND2X2 U3412 ( .A(net16633), .B(n3119), .Z(n99) );
  CENXL U3413 ( .A(net16005), .B(a[20]), .Z(n3330) );
  CENX2 U3414 ( .A(a[20]), .B(net16005), .Z(net19148) );
  CND2X2 U3415 ( .A(net19560), .B(n3119), .Z(n3331) );
  CND2X2 U3416 ( .A(net19560), .B(n3119), .Z(n3332) );
  CIVX2 U3417 ( .A(net16633), .Z(n3327) );
  CIVX1 U3418 ( .A(net21614), .Z(n3328) );
  CIVX2 U3419 ( .A(n3329), .Z(n3335) );
  CIVX2 U3420 ( .A(net16633), .Z(n3329) );
  CND2X1 U3421 ( .A(n1448), .B(n3825), .Z(n3826) );
  CND2X2 U3422 ( .A(n3826), .B(n3827), .Z(n3837) );
  CNIVX2 U3423 ( .A(n1735), .Z(n3337) );
  CENX1 U3424 ( .A(n2806), .B(net16671), .Z(n2476) );
  CENXL U3425 ( .A(n1489), .B(n3233), .Z(n3338) );
  CENX1 U3426 ( .A(n1489), .B(n3433), .Z(n1485) );
  CENX1 U3427 ( .A(n1491), .B(n1508), .Z(n3433) );
  CND3XL U3428 ( .A(n3831), .B(n3830), .C(n3829), .Z(n3339) );
  CENX1 U3429 ( .A(n3553), .B(n1171), .Z(n1165) );
  COR2XL U3430 ( .A(n1244), .B(n1215), .Z(n3341) );
  CIVXL U3431 ( .A(n530), .Z(n528) );
  CND3XL U3432 ( .A(n3786), .B(n3787), .C(n3788), .Z(n1412) );
  CIVX4 U3433 ( .A(n4005), .Z(n3982) );
  CENXL U3434 ( .A(n3985), .B(n3961), .Z(n3342) );
  CIVX2 U3435 ( .A(n4005), .Z(n4003) );
  CND2X1 U3436 ( .A(net19447), .B(net19448), .Z(n3345) );
  COND2X1 U3437 ( .A(n108), .B(n2412), .C(n3957), .D(n2411), .Z(n1890) );
  CEOX2 U3438 ( .A(n4017), .B(a[16]), .Z(n3346) );
  CIVX2 U3439 ( .A(n4007), .Z(n3347) );
  COND1X1 U3440 ( .A(n444), .B(n461), .C(n445), .Z(n439) );
  CANR1XL U3441 ( .A(n520), .B(n535), .C(n521), .Z(n3349) );
  COND2XL U3442 ( .A(n90), .B(n2467), .C(net19996), .D(n2466), .Z(n3350) );
  COND2XL U3443 ( .A(n90), .B(n2467), .C(net19996), .D(n2466), .Z(n3351) );
  CEO3X2 U3444 ( .A(n2005), .B(n2222), .C(n1800), .Z(n1329) );
  CND2XL U3445 ( .A(n1800), .B(n2222), .Z(n3877) );
  CIVX2 U3446 ( .A(net19890), .Z(net19695) );
  COND2XL U3447 ( .A(n3905), .B(n2757), .C(n6), .D(n2756), .Z(n2230) );
  CENX1 U3448 ( .A(n3985), .B(net19890), .Z(n2407) );
  COND2X1 U3449 ( .A(n3340), .B(n2534), .C(net16683), .D(n2533), .Z(n2007) );
  COND2XL U3450 ( .A(n2418), .B(n3334), .C(n2419), .D(n3331), .Z(n1897) );
  CNR2XL U3451 ( .A(n3336), .B(n2443), .Z(n3695) );
  CEOXL U3452 ( .A(n921), .B(n1900), .Z(n3385) );
  CFA1XL U3453 ( .A(n890), .B(n1897), .CI(n1809), .CO(n876), .S(n877) );
  CIVX1 U3454 ( .A(n3477), .Z(n1035) );
  CND2X1 U3455 ( .A(n3448), .B(n3449), .Z(n2378) );
  CIVXL U3456 ( .A(n1972), .Z(net21564) );
  CIVX1 U3457 ( .A(net21564), .Z(net21565) );
  CND2X2 U3458 ( .A(n3210), .B(n51), .Z(n3352) );
  CND2X2 U3459 ( .A(n3860), .B(n51), .Z(n3353) );
  CND2X2 U3460 ( .A(n3210), .B(n51), .Z(n3912) );
  COND2XL U3461 ( .A(n3705), .B(n2281), .C(net16617), .D(n2280), .Z(n3354) );
  CIVX2 U3462 ( .A(a[18]), .Z(n3718) );
  CENX1 U3463 ( .A(n1569), .B(n3427), .Z(n1565) );
  CND2XL U3464 ( .A(n1571), .B(n1569), .Z(n3540) );
  CIVXL U3465 ( .A(n1854), .Z(net21555) );
  CIVX1 U3466 ( .A(net21555), .Z(net21556) );
  CIVX4 U3467 ( .A(n3935), .Z(n3355) );
  CIVX4 U3468 ( .A(n3935), .Z(n3918) );
  CND2XL U3469 ( .A(a[4]), .B(n3697), .Z(n3358) );
  CND2X1 U3470 ( .A(n3356), .B(n4007), .Z(n3359) );
  CND2X2 U3471 ( .A(n3358), .B(n3359), .Z(n2825) );
  CIVXL U3472 ( .A(a[4]), .Z(n3356) );
  CND2XL U3473 ( .A(n1439), .B(n1441), .Z(n3975) );
  CND2IX1 U3474 ( .B(net16015), .A(a[14]), .Z(net18736) );
  CND3X2 U3475 ( .A(net19520), .B(net19521), .C(net19522), .Z(n1108) );
  CIVXL U3476 ( .A(n2094), .Z(net21539) );
  CIVXL U3477 ( .A(net21539), .Z(net21540) );
  CIVX2 U3478 ( .A(n3330), .Z(net19560) );
  CENX1 U3479 ( .A(n1062), .B(n3362), .Z(n1039) );
  CEO3X2 U3480 ( .A(n2096), .B(n1302), .C(n2220), .Z(n1263) );
  CND2XL U3481 ( .A(n2096), .B(n1302), .Z(n3363) );
  CND2X1 U3482 ( .A(n2096), .B(n2220), .Z(n3364) );
  CND2XL U3483 ( .A(n1302), .B(n2220), .Z(n3365) );
  CND3X1 U3484 ( .A(n3363), .B(n3364), .C(n3365), .Z(n1262) );
  CND2XL U3485 ( .A(n1233), .B(n1239), .Z(n3366) );
  CND2XL U3486 ( .A(n1233), .B(n1262), .Z(n3367) );
  CND2XL U3487 ( .A(n1239), .B(n1262), .Z(n3368) );
  CND3X1 U3488 ( .A(n3366), .B(n3367), .C(n3368), .Z(n1226) );
  CIVXL U3489 ( .A(n456), .Z(n3369) );
  CIVXL U3490 ( .A(n3099), .Z(n3370) );
  CIVX2 U3491 ( .A(n4005), .Z(n4004) );
  CND2X2 U3492 ( .A(n3896), .B(net18736), .Z(n3371) );
  CND2X2 U3493 ( .A(n3896), .B(net18736), .Z(n2820) );
  CEO3X2 U3494 ( .A(n912), .B(n910), .C(n899), .Z(n895) );
  CND2XL U3495 ( .A(n912), .B(n910), .Z(n3372) );
  CND2X1 U3496 ( .A(n912), .B(n899), .Z(n3373) );
  CND2XL U3497 ( .A(n910), .B(n899), .Z(n3374) );
  CND3X1 U3498 ( .A(n3372), .B(n3373), .C(n3374), .Z(n894) );
  CND2XL U3499 ( .A(n883), .B(n881), .Z(n3376) );
  CND2XL U3500 ( .A(n883), .B(n894), .Z(n3377) );
  CND2XL U3501 ( .A(n881), .B(n894), .Z(n3378) );
  CND3X1 U3502 ( .A(n3376), .B(n3377), .C(n3378), .Z(n878) );
  CNIVX3 U3503 ( .A(n48), .Z(n3961) );
  CEOX2 U3504 ( .A(n3379), .B(n1335), .Z(n1333) );
  CND2XL U3505 ( .A(n1335), .B(n1362), .Z(n3380) );
  CND2X1 U3506 ( .A(n1335), .B(n1337), .Z(n3381) );
  CND2XL U3507 ( .A(n1362), .B(n1337), .Z(n3382) );
  CND3X1 U3508 ( .A(n3380), .B(n3381), .C(n3382), .Z(n1332) );
  CEOX1 U3509 ( .A(n3777), .B(n1366), .Z(n1337) );
  CNR2X2 U3510 ( .A(n1305), .B(n1332), .Z(n3873) );
  COND2XL U3511 ( .A(n2286), .B(net18573), .C(net18772), .D(n2285), .Z(n1772)
         );
  COND2XL U3512 ( .A(net18573), .B(n2288), .C(net18772), .D(n2287), .Z(n810)
         );
  COND2XL U3513 ( .A(net18573), .B(n2292), .C(net18772), .D(n2291), .Z(n1777)
         );
  COND2XL U3514 ( .A(net18573), .B(n2295), .C(net18772), .D(n2294), .Z(n1780)
         );
  CENX1 U3515 ( .A(n1571), .B(n1584), .Z(n3427) );
  CENXL U3516 ( .A(n2782), .B(n4008), .Z(n2650) );
  CND2IXL U3517 ( .B(n1042), .A(n1021), .Z(n3680) );
  CND2X1 U3518 ( .A(n1065), .B(n1088), .Z(n3511) );
  CIVX1 U3519 ( .A(n448), .Z(n751) );
  CND2X2 U3520 ( .A(n3936), .B(n3937), .Z(n33) );
  CND2X1 U3521 ( .A(n1165), .B(n1190), .Z(n3636) );
  CNR2X1 U3522 ( .A(n578), .B(n594), .Z(n576) );
  CIVX2 U3523 ( .A(n591), .Z(n768) );
  CND2XL U3524 ( .A(n1173), .B(n1171), .Z(n3643) );
  CENX1 U3525 ( .A(n1173), .B(n1196), .Z(n3553) );
  CND2X1 U3526 ( .A(n1271), .B(n1269), .Z(n3967) );
  CND2X1 U3527 ( .A(n1271), .B(n1265), .Z(n3965) );
  COND2X1 U3528 ( .A(n2722), .B(n18), .C(net16638), .D(n2721), .Z(n2195) );
  CIVX3 U3529 ( .A(n12), .Z(n4005) );
  CENX1 U3530 ( .A(net16391), .B(net16671), .Z(n2471) );
  CND2X1 U3531 ( .A(n3146), .B(n1270), .Z(n3431) );
  CNR2XL U3532 ( .A(n1387), .B(n1412), .Z(n582) );
  CNR2X1 U3533 ( .A(n907), .B(n922), .Z(n402) );
  CEOX1 U3534 ( .A(n3385), .B(n936), .Z(n915) );
  CND2XL U3535 ( .A(n936), .B(n1900), .Z(n3386) );
  CND2XL U3536 ( .A(n936), .B(n921), .Z(n3387) );
  CND2XL U3537 ( .A(n1900), .B(n921), .Z(n3388) );
  CND3X1 U3538 ( .A(n3386), .B(n3387), .C(n3388), .Z(n914) );
  CIVXL U3539 ( .A(n920), .Z(n921) );
  CIVX2 U3540 ( .A(n1438), .Z(n3543) );
  CNR2XL U3541 ( .A(n514), .B(n3287), .Z(n3389) );
  CENX2 U3542 ( .A(n3483), .B(n3805), .Z(n3469) );
  CND2X1 U3543 ( .A(n969), .B(n988), .Z(n3390) );
  CND2X1 U3544 ( .A(n969), .B(n986), .Z(n3391) );
  CND2XL U3545 ( .A(n988), .B(n986), .Z(n3392) );
  CND3X1 U3546 ( .A(n3390), .B(n3391), .C(n3392), .Z(n964) );
  CND2X1 U3547 ( .A(n1488), .B(n1486), .Z(n3622) );
  CENX1 U3548 ( .A(n3551), .B(n1486), .Z(n1463) );
  CANR1X1 U3549 ( .A(n3550), .B(n384), .C(n377), .Z(n373) );
  CENX1 U3550 ( .A(n3994), .B(net18510), .Z(n2522) );
  COND1XL U3551 ( .A(n668), .B(n651), .C(n652), .Z(n3393) );
  CENX1 U3552 ( .A(n4005), .B(a[2]), .Z(n2826) );
  CND2IX2 U3553 ( .B(a[16]), .A(net19446), .Z(net19448) );
  CIVX1 U3554 ( .A(net19793), .Z(net20022) );
  CIVXL U3555 ( .A(n2003), .Z(n3394) );
  CIVX1 U3556 ( .A(n3394), .Z(n3395) );
  CEO3X2 U3557 ( .A(n1220), .B(n3799), .C(n3746), .Z(n3914) );
  CIVXL U3558 ( .A(n665), .Z(n779) );
  CNR2X1 U3559 ( .A(n514), .B(n3287), .Z(n478) );
  CND2XL U3560 ( .A(n1638), .B(n1636), .Z(n3760) );
  COND1XL U3561 ( .A(n540), .B(n544), .C(n541), .Z(n3396) );
  CND2X1 U3562 ( .A(n1245), .B(n1274), .Z(n544) );
  CIVX2 U3563 ( .A(n48), .Z(n3398) );
  CIVX2 U3564 ( .A(n48), .Z(n4016) );
  CND3X2 U3565 ( .A(n3783), .B(n3784), .C(n3785), .Z(n1414) );
  CND2X1 U3566 ( .A(n1442), .B(n1440), .Z(n3784) );
  CIVX2 U3567 ( .A(n378), .Z(n745) );
  CANR1X1 U3568 ( .A(n699), .B(n691), .C(n692), .Z(n690) );
  COND2XL U3569 ( .A(n18), .B(n2741), .C(net16639), .D(n2740), .Z(n2214) );
  CENXL U3570 ( .A(net16399), .B(n4004), .Z(n2739) );
  CENXL U3571 ( .A(n2806), .B(n4004), .Z(n2740) );
  CENXL U3572 ( .A(net16389), .B(n4004), .Z(n2734) );
  CENXL U3573 ( .A(net16391), .B(n4004), .Z(n2735) );
  CENXL U3574 ( .A(n3984), .B(n4004), .Z(n2744) );
  CENXL U3575 ( .A(net16393), .B(n4004), .Z(n2736) );
  CENXL U3576 ( .A(net16407), .B(n4004), .Z(n2743) );
  CENXL U3577 ( .A(n3985), .B(n4004), .Z(n2737) );
  CENXL U3578 ( .A(n3986), .B(n4004), .Z(n2733) );
  CENXL U3579 ( .A(n3988), .B(n4003), .Z(n2731) );
  CENXL U3580 ( .A(n3990), .B(n4004), .Z(n2729) );
  CENXL U3581 ( .A(n2808), .B(n4004), .Z(n2742) );
  CIVX1 U3582 ( .A(n4003), .Z(n3635) );
  CEO3X1 U3583 ( .A(n2113), .B(n3063), .C(n2082), .Z(n1635) );
  CND2XL U3584 ( .A(n2206), .B(n2082), .Z(n3399) );
  CND2XL U3585 ( .A(n2206), .B(n2113), .Z(n3400) );
  CND2XL U3586 ( .A(n2082), .B(n2113), .Z(n3401) );
  CND3X1 U3587 ( .A(n3399), .B(n3400), .C(n3401), .Z(n1634) );
  CENX2 U3588 ( .A(net16399), .B(net16671), .Z(n2475) );
  CIVDX3 U3589 ( .A(n4019), .Z0(n4018), .Z1(n3493) );
  CEO3X2 U3590 ( .A(n1883), .B(net21565), .C(n2095), .Z(n1235) );
  CND2XL U3591 ( .A(n2095), .B(n1972), .Z(n3402) );
  CND2XL U3592 ( .A(n1883), .B(n2095), .Z(n3403) );
  CND3X1 U3593 ( .A(n3402), .B(n3403), .C(n3404), .Z(n1234) );
  CEOX2 U3594 ( .A(n1236), .B(n1232), .Z(n3405) );
  CEOX2 U3595 ( .A(n3405), .B(n1234), .Z(n1201) );
  CND2XL U3596 ( .A(net16403), .B(n3212), .Z(n3407) );
  CND2X1 U3597 ( .A(n3407), .B(n3408), .Z(n2609) );
  CIVXL U3598 ( .A(n3961), .Z(n3406) );
  CEOX1 U3599 ( .A(n2101), .B(n1411), .Z(n3409) );
  CEOX1 U3600 ( .A(n3409), .B(n1434), .Z(n1401) );
  CND2XL U3601 ( .A(n1434), .B(n1411), .Z(n3410) );
  CND2X1 U3602 ( .A(n1434), .B(n2101), .Z(n3411) );
  CND2XL U3603 ( .A(n1411), .B(n2101), .Z(n3412) );
  CND3X1 U3604 ( .A(n3410), .B(n3411), .C(n3412), .Z(n1400) );
  CENX2 U3605 ( .A(n2793), .B(net18520), .Z(n2397) );
  CFA1XL U3606 ( .A(n2177), .B(n2115), .CI(n1733), .CO(n1658), .S(n1659) );
  CND2XL U3607 ( .A(net16389), .B(n3167), .Z(n3413) );
  CND2X1 U3608 ( .A(n3413), .B(n3414), .Z(n2536) );
  CIVXL U3609 ( .A(net16389), .Z(net21418) );
  CNIVX4 U3610 ( .A(n2800), .Z(net16389) );
  CIVX2 U3611 ( .A(n4010), .Z(n3930) );
  CEOX2 U3612 ( .A(n897), .B(n908), .Z(n3415) );
  CND2XL U3613 ( .A(n895), .B(n908), .Z(n3416) );
  CND2X1 U3614 ( .A(n895), .B(n897), .Z(n3417) );
  CND2XL U3615 ( .A(n908), .B(n897), .Z(n3418) );
  CND3XL U3616 ( .A(n3416), .B(n3417), .C(n3418), .Z(n892) );
  CIVX1 U3617 ( .A(n389), .Z(n746) );
  CND2XL U3618 ( .A(n3167), .B(n2808), .Z(n3422) );
  CIVXL U3619 ( .A(n2808), .Z(n3421) );
  CIVX4 U3620 ( .A(n3654), .Z(n3425) );
  CIVX4 U3621 ( .A(n3654), .Z(n3655) );
  CENX2 U3622 ( .A(n3426), .B(n1284), .Z(n1251) );
  CENX2 U3623 ( .A(n1259), .B(n1257), .Z(n3426) );
  CEOX2 U3624 ( .A(n1270), .B(n1268), .Z(n3428) );
  CEOX2 U3625 ( .A(n3428), .B(n1235), .Z(n1229) );
  CND2X1 U3626 ( .A(n1235), .B(n3147), .Z(n3429) );
  CND2X1 U3627 ( .A(n1235), .B(n1270), .Z(n3430) );
  CND3X2 U3628 ( .A(n3429), .B(n3430), .C(n3431), .Z(n1228) );
  CNIVX1 U3629 ( .A(n3733), .Z(n3432) );
  CNR2X1 U3630 ( .A(n440), .B(n385), .Z(n383) );
  CIVXL U3631 ( .A(n739), .Z(n3434) );
  CND2IXL U3632 ( .B(n353), .A(n3435), .Z(n298) );
  CNR2X1 U3633 ( .A(n309), .B(n3434), .Z(n3435) );
  CND2X2 U3634 ( .A(n3436), .B(n3437), .Z(n3438) );
  CND2X2 U3635 ( .A(n3892), .B(n3438), .Z(n3792) );
  CIVX1 U3636 ( .A(n1197), .Z(n3436) );
  CIVX2 U3637 ( .A(n1222), .Z(n3437) );
  CEOX2 U3638 ( .A(n1209), .B(n1207), .Z(n3439) );
  CEOX2 U3639 ( .A(n3439), .B(n1230), .Z(n1197) );
  CND2XL U3640 ( .A(n1207), .B(n1209), .Z(n3442) );
  CND3X2 U3641 ( .A(n3440), .B(n3441), .C(n3442), .Z(n1196) );
  CND2X1 U3642 ( .A(n3714), .B(n3444), .Z(n3445) );
  CND2X1 U3643 ( .A(n3443), .B(n1345), .Z(n3446) );
  CND2X1 U3644 ( .A(n3445), .B(n3446), .Z(n1339) );
  CIVX2 U3645 ( .A(n3714), .Z(n3443) );
  CIVXL U3646 ( .A(n1345), .Z(n3444) );
  CND2XL U3647 ( .A(net16403), .B(net16676), .Z(n3448) );
  CIVXL U3648 ( .A(net16403), .Z(n3447) );
  CIVX1 U3649 ( .A(net16676), .Z(net21345) );
  CEO3X1 U3650 ( .A(n1378), .B(n1376), .C(n1351), .Z(n1345) );
  CND2X1 U3651 ( .A(n1370), .B(n1347), .Z(n3717) );
  COND2X1 U3652 ( .A(n135), .B(net19987), .C(net18772), .D(n2317), .Z(n1725)
         );
  CND2X2 U3653 ( .A(n2813), .B(n132), .Z(n135) );
  CEO3X2 U3654 ( .A(n2191), .B(n1857), .C(n1886), .Z(n1327) );
  CEOX2 U3655 ( .A(n1329), .B(n1331), .Z(n3450) );
  CND2XL U3656 ( .A(n3170), .B(n1857), .Z(n3451) );
  CND2XL U3657 ( .A(n3170), .B(n1886), .Z(n3452) );
  CND2XL U3658 ( .A(n1857), .B(n1886), .Z(n3453) );
  CND3X1 U3659 ( .A(n3451), .B(n3452), .C(n3453), .Z(n1326) );
  CND2XL U3660 ( .A(n1329), .B(n1327), .Z(n3455) );
  CND2XL U3661 ( .A(n1331), .B(n1327), .Z(n3456) );
  CND3X1 U3662 ( .A(n3456), .B(n3455), .C(n3454), .Z(n1316) );
  COR2XL U3663 ( .A(n108), .B(n2408), .Z(n3457) );
  COR2XL U3664 ( .A(n3957), .B(n2407), .Z(n3458) );
  CND2X1 U3665 ( .A(n3457), .B(n3458), .Z(n1886) );
  CENXL U3666 ( .A(n2804), .B(net18520), .Z(n2408) );
  CNR2X1 U3667 ( .A(n1186), .B(net18607), .Z(net19953) );
  COND2X1 U3668 ( .A(n3747), .B(n2407), .C(n3957), .D(n2406), .Z(n1885) );
  COND2X1 U3669 ( .A(n2316), .B(n135), .C(n132), .D(n2315), .Z(n1801) );
  CND2XL U3670 ( .A(n2126), .B(n1826), .Z(n3459) );
  CND2X1 U3671 ( .A(n2126), .B(n1854), .Z(n3460) );
  CND2X1 U3672 ( .A(n1826), .B(n1854), .Z(n3461) );
  CND3X1 U3673 ( .A(n3459), .B(n3460), .C(n3461), .Z(n1236) );
  COND2X1 U3674 ( .A(n3163), .B(n2653), .C(n3424), .D(n2652), .Z(n2126) );
  CIVX2 U3675 ( .A(a[14]), .Z(net18734) );
  CIVX2 U3676 ( .A(n57), .Z(net16539) );
  CIVX8 U3677 ( .A(n3463), .Z(net16684) );
  CIVX4 U3678 ( .A(n3462), .Z(n3463) );
  CNIVX4 U3679 ( .A(n57), .Z(n3464) );
  CENX2 U3680 ( .A(a[14]), .B(n3464), .Z(n3462) );
  CENX2 U3681 ( .A(a[14]), .B(n3464), .Z(n3465) );
  CENX2 U3682 ( .A(a[14]), .B(n3464), .Z(net16683) );
  CENX2 U3683 ( .A(a[14]), .B(n3464), .Z(net16682) );
  CANR1X1 U3684 ( .A(n3389), .B(n3324), .C(net20025), .Z(n149) );
  CANR1X2 U3685 ( .A(net19939), .B(n3324), .C(net18901), .Z(net18429) );
  CND2X2 U3686 ( .A(n561), .B(n549), .Z(n547) );
  COND1X1 U3687 ( .A(n547), .B(n575), .C(n548), .Z(n546) );
  CNR2X2 U3688 ( .A(net16554), .B(n556), .Z(n549) );
  CNR2X1 U3689 ( .A(n1305), .B(n1332), .Z(n556) );
  CANR1X2 U3690 ( .A(n576), .B(n3466), .C(n577), .Z(n575) );
  CIVXL U3691 ( .A(n575), .Z(n574) );
  COND1X2 U3692 ( .A(n578), .B(n595), .C(n579), .Z(n577) );
  COAN1X1 U3693 ( .A(n582), .B(n592), .C(n583), .Z(n579) );
  CIVX2 U3694 ( .A(n603), .Z(n601) );
  CANR1XL U3695 ( .A(n608), .B(net18282), .C(n601), .Z(net18827) );
  CIVX1 U3696 ( .A(n606), .Z(n608) );
  COND1X1 U3697 ( .A(n613), .B(n630), .C(n614), .Z(n3466) );
  CIVX2 U3698 ( .A(n618), .Z(n616) );
  CANR1XL U3699 ( .A(net18280), .B(n3031), .C(n616), .Z(net19203) );
  CANR1X1 U3700 ( .A(n631), .B(n650), .C(n632), .Z(n630) );
  COND1X1 U3701 ( .A(n3596), .B(n637), .C(n634), .Z(n632) );
  CANR1X1 U3702 ( .A(n646), .B(net18274), .C(n3124), .Z(n637) );
  CANR1XL U3703 ( .A(n646), .B(net18274), .C(n3124), .Z(net19965) );
  CIVXL U3704 ( .A(n3124), .Z(net19362) );
  CIVX2 U3705 ( .A(n644), .Z(n646) );
  COND1X1 U3706 ( .A(n480), .B(n3467), .C(net22007), .Z(net18901) );
  CNR2X1 U3707 ( .A(n514), .B(n3287), .Z(net19939) );
  CANR1X1 U3708 ( .A(n3396), .B(n520), .C(n521), .Z(n3467) );
  CIVXL U3709 ( .A(n3349), .Z(n517) );
  COND1X1 U3710 ( .A(n530), .B(n522), .C(net19253), .Z(n521) );
  CND2X2 U3711 ( .A(n534), .B(n520), .Z(n514) );
  CANR1XL U3712 ( .A(n498), .B(n517), .C(net18744), .Z(n497) );
  CND2XL U3713 ( .A(n516), .B(n498), .Z(n496) );
  CNR2IXL U3714 ( .B(n498), .A(net18617), .Z(n489) );
  CANR1X1 U3715 ( .A(n520), .B(n535), .C(n3468), .Z(net18906) );
  COND1X1 U3716 ( .A(n530), .B(n522), .C(net19253), .Z(n3468) );
  CIVX4 U3717 ( .A(net16017), .Z(net18491) );
  CIVX2 U3718 ( .A(net16021), .Z(net16017) );
  CIVX1 U3719 ( .A(net16021), .Z(net16015) );
  CIVXL U3720 ( .A(net16021), .Z(net16019) );
  CNIVX4 U3721 ( .A(n2807), .Z(net16403) );
  COND1XL U3722 ( .A(n480), .B(net18906), .C(net22007), .Z(net20025) );
  COND2X2 U3723 ( .A(n2379), .B(n3168), .C(net16605), .D(n2378), .Z(n1859) );
  CIVX1 U3724 ( .A(n27), .Z(net19793) );
  COND2XL U3725 ( .A(n2352), .B(n3173), .C(net16606), .D(n2351), .Z(n1835) );
  COND2XL U3726 ( .A(n3172), .B(n2354), .C(net16606), .D(n2353), .Z(n1837) );
  COND2XL U3727 ( .A(n117), .B(n2365), .C(n2364), .D(net16605), .Z(n1845) );
  CFA1XL U3728 ( .A(n1778), .B(n1838), .CI(n1748), .CO(n850), .S(n851) );
  CIVX1 U3729 ( .A(n890), .Z(n891) );
  CFA1XL U3730 ( .A(n1745), .B(n1835), .CI(n1775), .CO(n822), .S(n823) );
  CIVXL U3731 ( .A(n415), .Z(n413) );
  COND2XL U3732 ( .A(n2670), .B(n36), .C(n3424), .D(n2669), .Z(n3470) );
  COND2XL U3733 ( .A(n3163), .B(n2670), .C(n3655), .D(n2669), .Z(n2143) );
  CENX1 U3734 ( .A(n3471), .B(n1797), .Z(n1239) );
  CENX1 U3735 ( .A(n2157), .B(n1913), .Z(n3471) );
  CND2XL U3736 ( .A(n1634), .B(n1636), .Z(n3761) );
  CIVX2 U3737 ( .A(n3478), .Z(n3472) );
  CIVXL U3738 ( .A(net16676), .Z(net20005) );
  CIVXL U3739 ( .A(net19793), .Z(net20002) );
  CIVX4 U3740 ( .A(net19927), .Z(net19996) );
  CNIVX2 U3741 ( .A(n2145), .Z(n3473) );
  CND3X1 U3742 ( .A(n3495), .B(n3496), .C(n3497), .Z(n1284) );
  CENXL U3743 ( .A(n3474), .B(n2168), .Z(n1517) );
  CENXL U3744 ( .A(n2137), .B(n2075), .Z(n3474) );
  CIVXL U3745 ( .A(net18537), .Z(net19987) );
  CIVX2 U3746 ( .A(n4022), .Z(n3476) );
  COND2XL U3747 ( .A(n3336), .B(n2428), .C(n3023), .D(n2427), .Z(n3477) );
  COND2XL U3748 ( .A(n126), .B(n2330), .C(net16623), .D(n2329), .Z(n1813) );
  CIVXL U3749 ( .A(n628), .Z(n626) );
  CIVX1 U3750 ( .A(n627), .Z(n773) );
  CND2XL U3751 ( .A(n634), .B(n774), .Z(n192) );
  CENX1 U3752 ( .A(net16391), .B(net19890), .Z(n2405) );
  CIVXL U3753 ( .A(net19793), .Z(net19977) );
  CIVX4 U3754 ( .A(n3983), .Z(n87) );
  CENXL U3755 ( .A(n2789), .B(n4007), .Z(n2690) );
  CENXL U3756 ( .A(n3992), .B(n4007), .Z(n2689) );
  CIVX1 U3757 ( .A(n3478), .Z(n3479) );
  CND2XL U3758 ( .A(n1495), .B(n1514), .Z(n3503) );
  CENX1 U3759 ( .A(n2808), .B(net16549), .Z(n2577) );
  CNR2X2 U3760 ( .A(n1413), .B(n1436), .Z(n591) );
  CND2XL U3761 ( .A(net18282), .B(n603), .Z(n187) );
  CND2X1 U3762 ( .A(n770), .B(net18282), .Z(n594) );
  COND1XL U3763 ( .A(n3596), .B(net19965), .C(n634), .Z(n3480) );
  CND2X1 U3764 ( .A(net18274), .B(n776), .Z(n636) );
  CIVXL U3765 ( .A(n776), .Z(n3481) );
  CNIVXL U3766 ( .A(n33), .Z(n3482) );
  CIVX1 U3767 ( .A(n438), .Z(n440) );
  CND2X2 U3768 ( .A(net19447), .B(n3361), .Z(n3484) );
  CENXL U3769 ( .A(n2804), .B(n4020), .Z(n3485) );
  CENX1 U3770 ( .A(n3990), .B(n4001), .Z(n2762) );
  CENX1 U3771 ( .A(n3989), .B(n4001), .Z(n2763) );
  CENXL U3772 ( .A(n3988), .B(net15979), .Z(n2368) );
  CENXL U3773 ( .A(n3989), .B(net15979), .Z(n2367) );
  CENXL U3774 ( .A(n2793), .B(net15975), .Z(n2364) );
  CENXL U3775 ( .A(n2794), .B(net15975), .Z(n2365) );
  CENXL U3776 ( .A(n3990), .B(net15975), .Z(n2366) );
  CENXL U3777 ( .A(n3987), .B(net15975), .Z(n2369) );
  CND2IXL U3778 ( .B(n3998), .A(net15975), .Z(n2383) );
  CENXL U3779 ( .A(n2791), .B(net15975), .Z(n2362) );
  CENXL U3780 ( .A(n3988), .B(net18485), .Z(n3486) );
  CIVX4 U3781 ( .A(net19200), .Z(net18485) );
  COND2XL U3782 ( .A(n126), .B(n2344), .C(net16623), .D(n2343), .Z(n1827) );
  CANR1X1 U3783 ( .A(n3942), .B(n356), .C(n349), .Z(n345) );
  CNIVX1 U3784 ( .A(n2176), .Z(n3488) );
  COND2X2 U3785 ( .A(n3913), .B(n2459), .C(net19996), .D(n3160), .Z(n1936) );
  CENX1 U3786 ( .A(n1225), .B(n1252), .Z(n3489) );
  CNIVX2 U3787 ( .A(n1191), .Z(n3490) );
  CENXL U3788 ( .A(n3792), .B(n1195), .Z(n1191) );
  COND2XL U3789 ( .A(n27), .B(n2684), .C(net18545), .D(n2683), .Z(n3491) );
  COND2XL U3790 ( .A(net18570), .B(n2257), .C(net16617), .D(n2256), .Z(n1743)
         );
  CENX1 U3791 ( .A(n3492), .B(n3728), .Z(n1241) );
  CENXL U3792 ( .A(n2188), .B(n3351), .Z(n3492) );
  CENX2 U3793 ( .A(a[18]), .B(n4019), .Z(net19927) );
  CENX2 U3794 ( .A(a[18]), .B(n4019), .Z(n3983) );
  CENXL U3795 ( .A(n2806), .B(n4012), .Z(n2641) );
  CENXL U3796 ( .A(n3984), .B(n4012), .Z(n2645) );
  CENXL U3797 ( .A(net16393), .B(n4012), .Z(n2637) );
  CENXL U3798 ( .A(net16399), .B(n4012), .Z(n2640) );
  CENXL U3799 ( .A(net16407), .B(n4012), .Z(n2644) );
  CENXL U3800 ( .A(net16389), .B(n4012), .Z(n2635) );
  CENXL U3801 ( .A(n3986), .B(n4012), .Z(n2634) );
  CENXL U3802 ( .A(n3993), .B(n4011), .Z(n2622) );
  CENXL U3803 ( .A(n2781), .B(n4011), .Z(n2616) );
  CENXL U3804 ( .A(n3995), .B(n4011), .Z(n2620) );
  CENXL U3805 ( .A(n3992), .B(n4011), .Z(n2623) );
  CENXL U3806 ( .A(n2783), .B(n4011), .Z(n2618) );
  CENXL U3807 ( .A(n2784), .B(n4011), .Z(n2619) );
  CENXL U3808 ( .A(n2789), .B(n4011), .Z(n2624) );
  CENXL U3809 ( .A(n2782), .B(n4011), .Z(n2617) );
  CENXL U3810 ( .A(n2792), .B(n4011), .Z(n2627) );
  CENXL U3811 ( .A(n2791), .B(n4011), .Z(n2626) );
  CEOX2 U3812 ( .A(n3989), .B(n3493), .Z(n2499) );
  COND2XL U3813 ( .A(net18570), .B(n2255), .C(net16617), .D(n2254), .Z(n800)
         );
  COND2XL U3814 ( .A(n2253), .B(n3705), .C(net16617), .D(n2252), .Z(n794) );
  CAOR1XL U3815 ( .A(n3023), .B(n3332), .C(n2417), .Z(n1895) );
  COND2XL U3816 ( .A(n2418), .B(n3332), .C(n3023), .D(n2417), .Z(n1896) );
  COND2XL U3817 ( .A(n3332), .B(n2422), .C(n3334), .D(n2421), .Z(n1900) );
  CND2XL U3818 ( .A(n1797), .B(n1913), .Z(n3668) );
  CFA1XL U3819 ( .A(n1808), .B(n1896), .CI(n1749), .CO(n862), .S(n863) );
  CENXL U3820 ( .A(n3494), .B(n3076), .Z(n1621) );
  CENXL U3821 ( .A(n3046), .B(n2205), .Z(n3494) );
  CND2XL U3822 ( .A(n1011), .B(n3149), .Z(n3685) );
  CENX1 U3823 ( .A(net16403), .B(net16649), .Z(n2444) );
  CEOX1 U3824 ( .A(n3729), .B(n1128), .Z(n1097) );
  CND2XL U3825 ( .A(n3053), .B(n1827), .Z(n3963) );
  CEO3X1 U3826 ( .A(n1295), .B(n1320), .C(n1297), .Z(n1285) );
  CND2XL U3827 ( .A(n1295), .B(n1320), .Z(n3495) );
  CND2XL U3828 ( .A(n1295), .B(n1297), .Z(n3496) );
  CND2XL U3829 ( .A(n1259), .B(n1257), .Z(n3498) );
  CND2XL U3830 ( .A(n1259), .B(n1284), .Z(n3499) );
  CND2XL U3831 ( .A(n1257), .B(n1284), .Z(n3500) );
  CND3X2 U3832 ( .A(n3498), .B(n3499), .C(n3500), .Z(n1250) );
  CENX1 U3833 ( .A(n3993), .B(n3933), .Z(n2688) );
  COND2X1 U3834 ( .A(n2613), .B(n3353), .C(n51), .D(n2612), .Z(n2086) );
  CND2X1 U3835 ( .A(n4007), .B(n3698), .Z(n3936) );
  CEO3X2 U3836 ( .A(n1501), .B(n1495), .C(n1514), .Z(n1489) );
  CND2X1 U3837 ( .A(n1501), .B(n1495), .Z(n3501) );
  CND2X1 U3838 ( .A(n1501), .B(n1514), .Z(n3502) );
  CND2XL U3839 ( .A(n1491), .B(n1508), .Z(n3504) );
  CND2X1 U3840 ( .A(n1491), .B(n1489), .Z(n3505) );
  CND2XL U3841 ( .A(n1508), .B(n1489), .Z(n3506) );
  CND3X1 U3842 ( .A(n3504), .B(n3505), .C(n3506), .Z(n1484) );
  CHA1XL U3843 ( .A(n1893), .B(n1728), .CO(n1502), .S(n1503) );
  CND3X1 U3844 ( .A(n3724), .B(n3725), .C(n3726), .Z(n1240) );
  CENXL U3845 ( .A(n2806), .B(net18408), .Z(n3507) );
  CEOX2 U3846 ( .A(n1088), .B(n1065), .Z(n3508) );
  CEOX2 U3847 ( .A(n3508), .B(n1086), .Z(n1061) );
  CND2X1 U3848 ( .A(n1086), .B(n1065), .Z(n3509) );
  CND2X1 U3849 ( .A(n1086), .B(n1088), .Z(n3510) );
  CND3X2 U3850 ( .A(n3509), .B(n3510), .C(n3511), .Z(n1060) );
  CND3X1 U3851 ( .A(n3615), .B(n3616), .C(n3617), .Z(n1088) );
  CIVXL U3852 ( .A(net19319), .Z(net19877) );
  CIVXL U3853 ( .A(n543), .Z(n762) );
  COND2X1 U3854 ( .A(n3905), .B(n2764), .C(n6), .D(n2763), .Z(n2237) );
  CND2X1 U3855 ( .A(n1476), .B(n1451), .Z(n3834) );
  CND2X1 U3856 ( .A(n1451), .B(n1474), .Z(n3836) );
  CANR1X1 U3857 ( .A(n283), .B(n356), .C(n3065), .Z(n282) );
  CANR1X1 U3858 ( .A(n320), .B(n356), .C(n323), .Z(n319) );
  CANR1X1 U3859 ( .A(n331), .B(n356), .C(n332), .Z(n330) );
  CENX1 U3860 ( .A(n2782), .B(n3961), .Z(n2584) );
  CND2XL U3861 ( .A(n2168), .B(n2075), .Z(n3512) );
  CND2XL U3862 ( .A(n2168), .B(n2137), .Z(n3513) );
  CND2XL U3863 ( .A(n2075), .B(n2137), .Z(n3514) );
  CND3X1 U3864 ( .A(n3512), .B(n3513), .C(n3514), .Z(n1516) );
  CND2XL U3865 ( .A(n1473), .B(n1492), .Z(n3515) );
  CND2X1 U3866 ( .A(n1473), .B(n1494), .Z(n3516) );
  CND2XL U3867 ( .A(n1492), .B(n1494), .Z(n3517) );
  COND2XL U3868 ( .A(n27), .B(n2695), .C(net18546), .D(n2694), .Z(n2168) );
  CENX1 U3869 ( .A(n1488), .B(n1467), .Z(n3551) );
  CENXL U3870 ( .A(n3996), .B(net18538), .Z(n2285) );
  CENXL U3871 ( .A(n3994), .B(net18538), .Z(n2291) );
  CENXL U3872 ( .A(n3995), .B(net18538), .Z(n2290) );
  CENXL U3873 ( .A(n2793), .B(net18538), .Z(n2298) );
  CEOX2 U3874 ( .A(n1375), .B(n1396), .Z(n3518) );
  CEOX2 U3875 ( .A(n3518), .B(n1373), .Z(n1367) );
  CND2X1 U3876 ( .A(n1373), .B(n1396), .Z(n3519) );
  CND2X1 U3877 ( .A(n1373), .B(n1375), .Z(n3520) );
  CND2X1 U3878 ( .A(n1396), .B(n1375), .Z(n3521) );
  CND3X2 U3879 ( .A(n3519), .B(n3520), .C(n3521), .Z(n1366) );
  COND1X1 U3880 ( .A(n361), .B(n417), .C(n362), .Z(n360) );
  CIVXL U3881 ( .A(n529), .Z(n760) );
  CIVXL U3882 ( .A(n308), .Z(n306) );
  CND2XL U3883 ( .A(n1424), .B(n1407), .Z(n3564) );
  CND2XL U3884 ( .A(n1424), .B(n1405), .Z(n3563) );
  CEOX1 U3885 ( .A(n3562), .B(n1424), .Z(n1395) );
  CEO3X2 U3886 ( .A(n1998), .B(n1968), .C(n1130), .Z(n1099) );
  CEOX2 U3887 ( .A(n1103), .B(n1105), .Z(n3522) );
  CEOX2 U3888 ( .A(n3522), .B(n1099), .Z(n1093) );
  CND2XL U3889 ( .A(n1998), .B(n1968), .Z(n3523) );
  CND2XL U3890 ( .A(n1998), .B(n1130), .Z(n3524) );
  CND2XL U3891 ( .A(n1968), .B(n1130), .Z(n3525) );
  CND3X1 U3892 ( .A(n3523), .B(n3524), .C(n3525), .Z(n1098) );
  CND2XL U3893 ( .A(n1103), .B(n1105), .Z(n3526) );
  CND2XL U3894 ( .A(n1103), .B(n1099), .Z(n3527) );
  CND2XL U3895 ( .A(n1105), .B(n1099), .Z(n3528) );
  CND3X1 U3896 ( .A(n3526), .B(n3527), .C(n3528), .Z(n1092) );
  CIVXL U3897 ( .A(net16580), .Z(net19845) );
  CENXL U3898 ( .A(n2793), .B(net16027), .Z(n2562) );
  CEO3X2 U3899 ( .A(n985), .B(n983), .C(n1002), .Z(n979) );
  CND2X1 U3900 ( .A(n985), .B(n983), .Z(n3529) );
  CND2XL U3901 ( .A(n985), .B(n1002), .Z(n3530) );
  CND2X1 U3902 ( .A(n983), .B(n1002), .Z(n3531) );
  CND3X2 U3903 ( .A(n3529), .B(n3530), .C(n3531), .Z(n978) );
  CEOX2 U3904 ( .A(n980), .B(n963), .Z(n3532) );
  CEOX2 U3905 ( .A(n978), .B(n3532), .Z(n959) );
  CND2XL U3906 ( .A(n963), .B(n980), .Z(n3533) );
  CND2XL U3907 ( .A(n980), .B(n978), .Z(n3534) );
  CND2XL U3908 ( .A(n963), .B(n978), .Z(n3535) );
  CND3X1 U3909 ( .A(n3533), .B(n3534), .C(n3535), .Z(n958) );
  CND3X2 U3910 ( .A(n3834), .B(n3835), .C(n3836), .Z(n1446) );
  CND2X1 U3911 ( .A(n1590), .B(n1575), .Z(n3537) );
  CND2X1 U3912 ( .A(n1573), .B(n1575), .Z(n3538) );
  CND2XL U3913 ( .A(n1571), .B(n1584), .Z(n3539) );
  CND2XL U3914 ( .A(n1584), .B(n1569), .Z(n3541) );
  CND3X1 U3915 ( .A(n3539), .B(n3540), .C(n3541), .Z(n1564) );
  CND3X2 U3916 ( .A(n3692), .B(n3693), .C(n3694), .Z(n1398) );
  CND2X1 U3917 ( .A(n1438), .B(n3542), .Z(n3545) );
  CND2X2 U3918 ( .A(n3545), .B(n3544), .Z(n3782) );
  CIVXL U3919 ( .A(n1417), .Z(n3542) );
  CND2X1 U3920 ( .A(n658), .B(n3944), .Z(n651) );
  CIVXL U3921 ( .A(net19793), .Z(net19794) );
  CEO3X2 U3922 ( .A(n1383), .B(n1381), .C(n1377), .Z(n1371) );
  CND2XL U3923 ( .A(n1383), .B(n1377), .Z(n3546) );
  CND2X1 U3924 ( .A(n1377), .B(n1381), .Z(n3548) );
  CND3X2 U3925 ( .A(n3546), .B(n3547), .C(n3548), .Z(n1370) );
  CNIVX4 U3926 ( .A(a[8]), .Z(n3549) );
  COND2X1 U3927 ( .A(n3904), .B(n2629), .C(n3959), .D(n2628), .Z(n2102) );
  CENX1 U3928 ( .A(n3549), .B(n4008), .Z(n3959) );
  CDLY1XL U3929 ( .A(n745), .Z(n3550) );
  CENX1 U3930 ( .A(net16399), .B(net16649), .Z(n2442) );
  CND2IX2 U3931 ( .B(n3552), .A(n1214), .Z(n530) );
  CND2XL U3932 ( .A(n867), .B(n878), .Z(n370) );
  CIVXL U3933 ( .A(n379), .Z(n377) );
  CENX1 U3934 ( .A(n3984), .B(n3476), .Z(n2348) );
  CND2XL U3935 ( .A(n462), .B(n3419), .Z(n451) );
  CENXL U3936 ( .A(n2794), .B(net16027), .Z(n2563) );
  CIVXL U3937 ( .A(n532), .Z(net19757) );
  CIVXL U3938 ( .A(net19753), .Z(net19754) );
  COND2X1 U3939 ( .A(n2550), .B(n3058), .C(n3055), .D(n2549), .Z(n2023) );
  CFA1X1 U3940 ( .A(n1844), .B(n2023), .CI(n1757), .CO(n990), .S(n991) );
  CENX1 U3941 ( .A(n2806), .B(net16649), .Z(n2443) );
  CEO3XL U3942 ( .A(n1487), .B(n1506), .C(n3338), .Z(n3554) );
  CIVX1 U3943 ( .A(n605), .Z(n770) );
  CEOX1 U3944 ( .A(n1509), .B(n1526), .Z(n3763) );
  CND2XL U3945 ( .A(n1526), .B(n1509), .Z(n3766) );
  CIVXL U3946 ( .A(n3384), .Z(n747) );
  CND2X1 U3947 ( .A(n1221), .B(n1250), .Z(n3886) );
  CEO3X1 U3948 ( .A(n1046), .B(n1048), .C(n1027), .Z(n1021) );
  CND2XL U3949 ( .A(n1046), .B(n1027), .Z(n3555) );
  CND2XL U3950 ( .A(n1046), .B(n1048), .Z(n3556) );
  CND2X1 U3951 ( .A(n1027), .B(n1048), .Z(n3557) );
  CENXL U3952 ( .A(n2781), .B(n4017), .Z(n2484) );
  CENXL U3953 ( .A(n2783), .B(n4017), .Z(n2486) );
  CENXL U3954 ( .A(n3994), .B(n4017), .Z(n2489) );
  CENXL U3955 ( .A(n2782), .B(n4017), .Z(n2485) );
  CENXL U3956 ( .A(n3992), .B(n4017), .Z(n2491) );
  CENXL U3957 ( .A(n3991), .B(n4017), .Z(n2493) );
  CENXL U3958 ( .A(n2789), .B(n4017), .Z(n2492) );
  CENXL U3959 ( .A(n2784), .B(n4017), .Z(n2487) );
  CENXL U3960 ( .A(n2791), .B(n4017), .Z(n2494) );
  CENXL U3961 ( .A(n3993), .B(n4017), .Z(n2490) );
  CENXL U3962 ( .A(n2792), .B(n4017), .Z(n2495) );
  CENXL U3963 ( .A(n2804), .B(n4017), .Z(n2507) );
  CENXL U3964 ( .A(n187), .B(n604), .Z(product[25]) );
  CND2XL U3965 ( .A(n3159), .B(n922), .Z(n3558) );
  CND2XL U3966 ( .A(n4014), .B(a[8]), .Z(n3560) );
  CND2X1 U3967 ( .A(n3559), .B(n3235), .Z(n3561) );
  CND2X2 U3968 ( .A(n3560), .B(n3561), .Z(n2823) );
  CND2X1 U3969 ( .A(n1305), .B(n1332), .Z(n559) );
  CND2XL U3970 ( .A(n1405), .B(n1407), .Z(n3565) );
  CND3X1 U3971 ( .A(n3563), .B(n3564), .C(n3565), .Z(n1394) );
  CEOX1 U3972 ( .A(n2173), .B(n2142), .Z(n3566) );
  CEOX1 U3973 ( .A(n3566), .B(n1611), .Z(n1605) );
  CND2XL U3974 ( .A(n2142), .B(n2173), .Z(n3569) );
  CIVXL U3975 ( .A(n3918), .Z(n3570) );
  CIVXL U3976 ( .A(n3570), .Z(n3571) );
  CENX1 U3977 ( .A(n3995), .B(n3930), .Z(n2653) );
  CND3X2 U3978 ( .A(n3740), .B(n3739), .C(n3741), .Z(n1220) );
  CND2X1 U3979 ( .A(n1254), .B(n1227), .Z(n3739) );
  CIVXL U3980 ( .A(n458), .Z(n456) );
  COND2X1 U3981 ( .A(n3353), .B(n2607), .C(n51), .D(n2606), .Z(n2080) );
  CENX2 U3982 ( .A(a[0]), .B(n4002), .Z(n2827) );
  CND2X2 U3983 ( .A(n396), .B(n363), .Z(n361) );
  CNR2X2 U3984 ( .A(net16554), .B(n3873), .Z(n3854) );
  CENX2 U3985 ( .A(n3917), .B(n3972), .Z(n1359) );
  CENX1 U3986 ( .A(n3986), .B(net18944), .Z(n2403) );
  CND2XL U3987 ( .A(n3984), .B(net18944), .Z(n3573) );
  CNIVX4 U3988 ( .A(n2810), .Z(n3984) );
  CND2X2 U3989 ( .A(n1015), .B(n1036), .Z(n469) );
  CND2X1 U3990 ( .A(n1009), .B(n3593), .Z(n3594) );
  CANR1X1 U3991 ( .A(n478), .B(n546), .C(n3855), .Z(n3922) );
  CIVX1 U3992 ( .A(n418), .Z(net19689) );
  CIVXL U3993 ( .A(n416), .Z(n418) );
  CIVX1 U3994 ( .A(n1188), .Z(net19035) );
  CND2X1 U3995 ( .A(n1347), .B(n3576), .Z(n3577) );
  CND2X2 U3996 ( .A(n3575), .B(n1370), .Z(n3578) );
  CND2X2 U3997 ( .A(n3577), .B(n3578), .Z(n3714) );
  CIVX1 U3998 ( .A(n1347), .Z(n3575) );
  CIVX1 U3999 ( .A(n1370), .Z(n3576) );
  COND2X1 U4000 ( .A(net22025), .B(n2455), .C(net19996), .D(n2454), .Z(n1932)
         );
  CEO3XL U4001 ( .A(n1549), .B(n1564), .C(n3209), .Z(n3579) );
  CND2X2 U4002 ( .A(n3056), .B(net16617), .Z(n144) );
  CND2X1 U4003 ( .A(n1253), .B(n1278), .Z(n3822) );
  CENX1 U4004 ( .A(n3991), .B(net16023), .Z(n2559) );
  CEO3X2 U4005 ( .A(n1069), .B(n1067), .C(n1090), .Z(n1063) );
  CND2X1 U4006 ( .A(n1069), .B(n1067), .Z(n3580) );
  CND2XL U4007 ( .A(n1069), .B(n1090), .Z(n3581) );
  CND2X1 U4008 ( .A(n1067), .B(n1090), .Z(n3582) );
  CND3X2 U4009 ( .A(n3580), .B(n3581), .C(n3582), .Z(n1062) );
  CND2XL U4010 ( .A(n1064), .B(n1043), .Z(n3583) );
  CEO3X2 U4011 ( .A(n1081), .B(n1848), .C(n1967), .Z(n1073) );
  CND2XL U4012 ( .A(n1081), .B(n1967), .Z(n3586) );
  CND2XL U4013 ( .A(n1081), .B(n1848), .Z(n3587) );
  CND2XL U4014 ( .A(n1967), .B(n1848), .Z(n3588) );
  CND3X1 U4015 ( .A(n3586), .B(n3587), .C(n3588), .Z(n1072) );
  COND2XL U4016 ( .A(n3189), .B(n2492), .C(net18902), .D(n2491), .Z(n1967) );
  CIVX1 U4017 ( .A(n1080), .Z(n1081) );
  CND2XL U4018 ( .A(n2081), .B(n2205), .Z(n3589) );
  CND2XL U4019 ( .A(n2174), .B(n2081), .Z(n3590) );
  CND2XL U4020 ( .A(n2205), .B(n2174), .Z(n3591) );
  CND3X1 U4021 ( .A(n3589), .B(n3591), .C(n3590), .Z(n1620) );
  CND2X1 U4022 ( .A(n3592), .B(n1013), .Z(n3595) );
  CND2X2 U4023 ( .A(n3594), .B(n3595), .Z(n3683) );
  CIVX1 U4024 ( .A(n1013), .Z(n3593) );
  CND2XL U4025 ( .A(n2188), .B(n1942), .Z(n3726) );
  CND2XL U4026 ( .A(n1378), .B(n1351), .Z(n3597) );
  CND2XL U4027 ( .A(n1378), .B(n1376), .Z(n3598) );
  CND2XL U4028 ( .A(n1351), .B(n1376), .Z(n3599) );
  CND3X1 U4029 ( .A(n3597), .B(n3598), .C(n3599), .Z(n1344) );
  COR2XL U4030 ( .A(n3913), .B(n2472), .Z(n3600) );
  COR2XL U4031 ( .A(net19422), .B(n2471), .Z(n3601) );
  CND2X1 U4032 ( .A(n3600), .B(n3601), .Z(n1947) );
  CENX1 U4033 ( .A(net16393), .B(net19890), .Z(n2406) );
  CENX1 U4034 ( .A(n2782), .B(n3357), .Z(n2683) );
  COND2X1 U4035 ( .A(net18613), .B(n3247), .C(net16683), .D(n2528), .Z(n3699)
         );
  CND2XL U4036 ( .A(n3343), .B(n1759), .Z(n3602) );
  CND2XL U4037 ( .A(n1759), .B(n2056), .Z(n3603) );
  CND2XL U4038 ( .A(n2056), .B(n3343), .Z(n3604) );
  CND3X1 U4039 ( .A(n3602), .B(n3603), .C(n3604), .Z(n1032) );
  CIVXL U4040 ( .A(n1759), .Z(n3605) );
  CIVX2 U4041 ( .A(n3605), .Z(n3606) );
  COND2XL U4042 ( .A(n3705), .B(n2273), .C(net16617), .D(n2272), .Z(n1759) );
  CND2X2 U4043 ( .A(net19617), .B(net19618), .Z(n3607) );
  CND2X2 U4044 ( .A(net19619), .B(n3607), .Z(n1199) );
  CNIVX4 U4045 ( .A(net16019), .Z(net16645) );
  CFA1X1 U4046 ( .A(n1930), .B(n1871), .CI(n1783), .CO(n916), .S(n917) );
  COND2X1 U4047 ( .A(net22025), .B(n2453), .C(net19996), .D(n2452), .Z(n1930)
         );
  CHA1XL U4048 ( .A(n2086), .B(n2117), .CO(n1682), .S(n1683) );
  CEO3X2 U4049 ( .A(n1150), .B(n1148), .C(n1152), .Z(n1119) );
  CND2XL U4050 ( .A(n1150), .B(n1152), .Z(n3608) );
  CND2X1 U4051 ( .A(n1150), .B(n1148), .Z(n3609) );
  CND2X1 U4052 ( .A(n1152), .B(n1148), .Z(n3610) );
  COND2X1 U4053 ( .A(n126), .B(n2346), .C(net16621), .D(n2345), .Z(n1829) );
  CEOXL U4054 ( .A(n1087), .B(n1108), .Z(n3611) );
  CEOXL U4055 ( .A(n3611), .B(n1085), .Z(n1083) );
  CND2XL U4056 ( .A(n1085), .B(n1108), .Z(n3612) );
  CND2XL U4057 ( .A(n1085), .B(n1087), .Z(n3613) );
  CND2XL U4058 ( .A(n1108), .B(n1087), .Z(n3614) );
  CND3X1 U4059 ( .A(n3612), .B(n3613), .C(n3614), .Z(n1082) );
  CEO3X2 U4060 ( .A(n1116), .B(n1097), .C(n1095), .Z(n1089) );
  CND2XL U4061 ( .A(n1116), .B(n1095), .Z(n3615) );
  CND2XL U4062 ( .A(n1116), .B(n1097), .Z(n3616) );
  CND2X1 U4063 ( .A(n1095), .B(n1097), .Z(n3617) );
  CENXL U4064 ( .A(n3996), .B(net16649), .Z(n2417) );
  CENXL U4065 ( .A(n3984), .B(net16649), .Z(n2447) );
  CENX1 U4066 ( .A(net16393), .B(net16649), .Z(n2439) );
  CENX1 U4067 ( .A(n3985), .B(net16649), .Z(n2440) );
  CEO3X2 U4068 ( .A(n1512), .B(n1493), .C(n1510), .Z(n1487) );
  CND2X1 U4069 ( .A(n1512), .B(n1510), .Z(n3618) );
  CND2X1 U4070 ( .A(n1512), .B(n1493), .Z(n3619) );
  CND2X1 U4071 ( .A(n1510), .B(n1493), .Z(n3620) );
  CND3X2 U4072 ( .A(n3618), .B(n3619), .C(n3620), .Z(n1486) );
  CND2XL U4073 ( .A(n1467), .B(n1488), .Z(n3621) );
  COR2X1 U4074 ( .A(n3188), .B(n2511), .Z(n3624) );
  CND2X2 U4075 ( .A(n3624), .B(n3625), .Z(n1985) );
  CIVX1 U4076 ( .A(a[28]), .Z(net18809) );
  CND2X1 U4077 ( .A(n1287), .B(n1314), .Z(n3707) );
  CND2X1 U4078 ( .A(n1287), .B(n3221), .Z(n3708) );
  CENXL U4079 ( .A(n3992), .B(n4003), .Z(n2722) );
  CIVX4 U4080 ( .A(net19200), .Z(net18486) );
  CIVXL U4081 ( .A(n3162), .Z(n564) );
  CEO3X2 U4082 ( .A(n2089), .B(n1907), .C(n3634), .Z(n1079) );
  CND2XL U4083 ( .A(n1907), .B(n2089), .Z(n3626) );
  CND2XL U4084 ( .A(n1907), .B(n1791), .Z(n3627) );
  CND2X1 U4085 ( .A(n2089), .B(n1791), .Z(n3628) );
  CND3X1 U4086 ( .A(n3626), .B(n3627), .C(n3628), .Z(n1078) );
  CEOX2 U4087 ( .A(n2088), .B(n1076), .Z(n3629) );
  CEOX2 U4088 ( .A(n1078), .B(n3629), .Z(n1049) );
  CND2XL U4089 ( .A(n2088), .B(n1076), .Z(n3630) );
  CND2X1 U4090 ( .A(n2088), .B(n1078), .Z(n3631) );
  CND2XL U4091 ( .A(n1076), .B(n1078), .Z(n3632) );
  CND3X1 U4092 ( .A(n3630), .B(n3631), .C(n3632), .Z(n1048) );
  CIVXL U4093 ( .A(n1791), .Z(n3633) );
  CIVX1 U4094 ( .A(n3633), .Z(n3634) );
  CENXL U4095 ( .A(n2806), .B(n3961), .Z(n2608) );
  CENXL U4096 ( .A(n3988), .B(n3961), .Z(n2599) );
  CENXL U4097 ( .A(n2793), .B(n3961), .Z(n3901) );
  CENXL U4098 ( .A(net16399), .B(n3961), .Z(n2607) );
  CENXL U4099 ( .A(n3996), .B(n3961), .Z(n2582) );
  CENXL U4100 ( .A(n2808), .B(n3961), .Z(n2610) );
  CENXL U4101 ( .A(net16407), .B(n3961), .Z(n2611) );
  CENXL U4102 ( .A(n3987), .B(n3212), .Z(n2600) );
  CENXL U4103 ( .A(n3990), .B(n4015), .Z(n2597) );
  CENXL U4104 ( .A(n3994), .B(n4015), .Z(n2588) );
  CND2IXL U4105 ( .B(n3998), .A(n3806), .Z(n2614) );
  CND2XL U4106 ( .A(n2827), .B(n6), .Z(n3906) );
  CND2X4 U4107 ( .A(n2827), .B(n6), .Z(n9) );
  CND2X2 U4108 ( .A(net16637), .B(n2826), .Z(n18) );
  CEO3X1 U4109 ( .A(n1192), .B(n1165), .C(n1190), .Z(n1161) );
  CEO3X2 U4110 ( .A(n1208), .B(n1179), .C(n1177), .Z(n1171) );
  CND3X2 U4111 ( .A(n3639), .B(n3640), .C(n3641), .Z(n1170) );
  CND2XL U4112 ( .A(n1173), .B(n1196), .Z(n3642) );
  CND2XL U4113 ( .A(n1196), .B(n1171), .Z(n3644) );
  CND3X1 U4114 ( .A(n3642), .B(n3643), .C(n3644), .Z(n1164) );
  CENX1 U4115 ( .A(n2793), .B(net16671), .Z(n2463) );
  CND2X1 U4116 ( .A(n3744), .B(n1120), .Z(n3647) );
  CND2X2 U4117 ( .A(n3645), .B(n3646), .Z(n3648) );
  CND2X2 U4118 ( .A(n3647), .B(n3648), .Z(n1091) );
  CIVXL U4119 ( .A(n1120), .Z(n3646) );
  CND2IXL U4120 ( .B(a[6]), .A(n3697), .Z(n3937) );
  CEO3X2 U4121 ( .A(n1176), .B(n1153), .C(n1151), .Z(n1145) );
  CND2X1 U4122 ( .A(n1176), .B(n1151), .Z(n3650) );
  CND3X1 U4123 ( .A(net19536), .B(n3652), .C(net19538), .Z(n1138) );
  CIVXL U4124 ( .A(net21583), .Z(net19526) );
  COND2X1 U4125 ( .A(n3168), .B(net20005), .C(n2383), .D(net21572), .Z(n1727)
         );
  COND2XL U4126 ( .A(n3058), .B(n2579), .C(n3355), .D(n2578), .Z(n2052) );
  COND2XL U4127 ( .A(n63), .B(n2566), .C(n3355), .D(n2565), .Z(n2039) );
  COND2X1 U4128 ( .A(n2562), .B(n3059), .C(n3355), .D(n2561), .Z(n2035) );
  CENXL U4129 ( .A(n2781), .B(net18485), .Z(n2418) );
  CENXL U4130 ( .A(n3995), .B(net18485), .Z(n2422) );
  CENXL U4131 ( .A(n3993), .B(net18485), .Z(n2424) );
  CENXL U4132 ( .A(n3994), .B(net18485), .Z(n2423) );
  CENXL U4133 ( .A(n3988), .B(net18485), .Z(n2434) );
  CENX1 U4134 ( .A(n3986), .B(net18485), .Z(n2436) );
  CENXL U4135 ( .A(a[6]), .B(n30), .Z(n3934) );
  COND2X2 U4136 ( .A(n3747), .B(n2393), .C(n3957), .D(n2392), .Z(n954) );
  CANR1XL U4137 ( .A(n631), .B(n3393), .C(n3480), .Z(n3653) );
  CIVX8 U4138 ( .A(n3960), .Z(n3654) );
  CND2X1 U4139 ( .A(n3152), .B(n3902), .Z(n3658) );
  CND2X2 U4140 ( .A(n3656), .B(n3657), .Z(n3659) );
  CND2X2 U4141 ( .A(n3658), .B(n3659), .Z(n1257) );
  CIVXL U4142 ( .A(n1269), .Z(n3656) );
  CENXL U4143 ( .A(n2781), .B(net18510), .Z(n2517) );
  CENXL U4144 ( .A(n2783), .B(n3167), .Z(n2519) );
  CENXL U4145 ( .A(n3995), .B(net18510), .Z(n2521) );
  CENXL U4146 ( .A(n3992), .B(net18510), .Z(n2524) );
  CENXL U4147 ( .A(n3991), .B(net18510), .Z(n2526) );
  CENXL U4148 ( .A(n2804), .B(net18510), .Z(n2540) );
  CEO3X2 U4149 ( .A(n1997), .B(n1820), .C(n1761), .Z(n1075) );
  CND2X1 U4150 ( .A(n1997), .B(n1820), .Z(n3661) );
  CND2XL U4151 ( .A(n1997), .B(n1761), .Z(n3662) );
  CND2XL U4152 ( .A(n1820), .B(n1761), .Z(n3663) );
  CND3X1 U4153 ( .A(n3661), .B(n3662), .C(n3663), .Z(n1074) );
  CND2XL U4154 ( .A(n1102), .B(n1077), .Z(n3664) );
  CND2XL U4155 ( .A(n1102), .B(n1075), .Z(n3665) );
  CND2XL U4156 ( .A(n1077), .B(n1075), .Z(n3666) );
  CND3X1 U4157 ( .A(n3664), .B(n3665), .C(n3666), .Z(n1068) );
  COND2XL U4158 ( .A(n144), .B(n2275), .C(net16617), .D(n2274), .Z(n1761) );
  CENXL U4159 ( .A(n3996), .B(n4006), .Z(n2681) );
  CENXL U4160 ( .A(n3667), .B(n524), .Z(product[35]) );
  CND2XL U4161 ( .A(net19253), .B(n3980), .Z(n3667) );
  CND2XL U4162 ( .A(n1797), .B(n3491), .Z(n3669) );
  CND2XL U4163 ( .A(n1913), .B(n3491), .Z(n3670) );
  CND3X1 U4164 ( .A(n3668), .B(n3669), .C(n3670), .Z(n1238) );
  COND2X1 U4165 ( .A(n3173), .B(n2359), .C(net16606), .D(n2358), .Z(n1840) );
  COND1X1 U4166 ( .A(n261), .B(n354), .C(n262), .Z(n260) );
  CNR2X2 U4167 ( .A(n1215), .B(n1244), .Z(n3911) );
  CND2X2 U4168 ( .A(net18537), .B(net18809), .Z(n3883) );
  CEOX1 U4169 ( .A(n2066), .B(n1828), .Z(n3671) );
  CEOX1 U4170 ( .A(n3671), .B(n1856), .Z(n1295) );
  CND2XL U4171 ( .A(n1856), .B(n1828), .Z(n3672) );
  CND2XL U4172 ( .A(n1856), .B(n2066), .Z(n3673) );
  CND2XL U4173 ( .A(n1828), .B(n2066), .Z(n3674) );
  CND3X1 U4174 ( .A(n3672), .B(n3673), .C(n3674), .Z(n1294) );
  COND2X1 U4175 ( .A(n3682), .B(n2345), .C(net16623), .D(n2344), .Z(n1828) );
  CND2X1 U4176 ( .A(n965), .B(n982), .Z(n3676) );
  CND2X1 U4177 ( .A(n965), .B(n967), .Z(n3677) );
  CND2X1 U4178 ( .A(n982), .B(n967), .Z(n3678) );
  CND3X2 U4179 ( .A(n3676), .B(n3677), .C(n3678), .Z(n960) );
  CND2X1 U4180 ( .A(n1042), .B(n3099), .Z(n3679) );
  CND3X1 U4181 ( .A(n3893), .B(n3745), .C(n3895), .Z(n3746) );
  CENX2 U4182 ( .A(a[10]), .B(n3157), .Z(n3681) );
  CENX2 U4183 ( .A(a[10]), .B(n4014), .Z(n3981) );
  CND2X4 U4184 ( .A(n2814), .B(net16621), .Z(n3682) );
  CND2X2 U4185 ( .A(n2814), .B(net16621), .Z(n126) );
  CIVX2 U4186 ( .A(net18492), .Z(net19446) );
  CND2X2 U4187 ( .A(n1159), .B(n1186), .Z(net19253) );
  CIVX4 U4188 ( .A(n4022), .Z(n4021) );
  CND2XL U4189 ( .A(n1941), .B(net21540), .Z(n3845) );
  CND2IXL U4190 ( .B(n3998), .A(net16671), .Z(n2482) );
  CENXL U4191 ( .A(n3996), .B(net16001), .Z(n2450) );
  CENX1 U4192 ( .A(n2794), .B(net16671), .Z(n2464) );
  CENXL U4193 ( .A(n3985), .B(net19877), .Z(n2473) );
  CENXL U4194 ( .A(net16393), .B(net16671), .Z(n2472) );
  CENX2 U4195 ( .A(n3989), .B(net16671), .Z(n2466) );
  CEOX2 U4196 ( .A(n1011), .B(n3683), .Z(n1003) );
  CND2XL U4197 ( .A(n1011), .B(n1013), .Z(n3684) );
  CND2XL U4198 ( .A(n1013), .B(n1009), .Z(n3686) );
  CND3X1 U4199 ( .A(n3684), .B(n3685), .C(n3686), .Z(n1002) );
  CIVXL U4200 ( .A(n4011), .Z(n3687) );
  CENXL U4201 ( .A(n3985), .B(net18408), .Z(n2308) );
  CENXL U4202 ( .A(net16389), .B(net18408), .Z(n2305) );
  CENXL U4203 ( .A(n3988), .B(net18408), .Z(n2302) );
  CENXL U4204 ( .A(n3991), .B(net18408), .Z(n2295) );
  COND1XL U4205 ( .A(n361), .B(n417), .C(n362), .Z(net19415) );
  CANR1XL U4206 ( .A(n3142), .B(n415), .C(n3306), .Z(n395) );
  CANR1XL U4207 ( .A(n748), .B(n415), .C(n408), .Z(n406) );
  CENX1 U4208 ( .A(net16403), .B(net19890), .Z(n2411) );
  CEO3X2 U4209 ( .A(n2195), .B(n1949), .C(n1920), .Z(n1431) );
  CND2XL U4210 ( .A(n2195), .B(n1949), .Z(n3688) );
  CND2XL U4211 ( .A(n2195), .B(n1920), .Z(n3689) );
  CND2XL U4212 ( .A(n1949), .B(n1920), .Z(n3690) );
  CND3X1 U4213 ( .A(n3688), .B(n3689), .C(n3690), .Z(n1430) );
  CND2X1 U4214 ( .A(n1432), .B(n1428), .Z(n3692) );
  CND2X1 U4215 ( .A(n1432), .B(n1430), .Z(n3693) );
  CND2X1 U4216 ( .A(n1428), .B(n1430), .Z(n3694) );
  CNR2XL U4217 ( .A(n3333), .B(n2442), .Z(n3696) );
  COR2X1 U4218 ( .A(n3695), .B(n3696), .Z(n1920) );
  CIVXL U4219 ( .A(n3596), .Z(n774) );
  CENXL U4220 ( .A(n635), .B(n192), .Z(product[20]) );
  CIVXL U4221 ( .A(n572), .Z(n766) );
  CENX2 U4222 ( .A(a[26]), .B(n4022), .Z(n2814) );
  CIVX4 U4223 ( .A(n4010), .Z(n4008) );
  CIVX2 U4224 ( .A(n3712), .Z(n3711) );
  CNIVX4 U4225 ( .A(a[6]), .Z(n3698) );
  CENX2 U4226 ( .A(n1063), .B(n1084), .Z(net19385) );
  CENX1 U4227 ( .A(n2808), .B(net19890), .Z(n2412) );
  COND2X1 U4228 ( .A(net18613), .B(n3246), .C(net16683), .D(n2528), .Z(n1242)
         );
  CEO3XL U4229 ( .A(n1112), .B(n3339), .C(n1089), .Z(net19382) );
  CEOXL U4230 ( .A(n2121), .B(n2028), .Z(n3729) );
  COND2X1 U4231 ( .A(n3747), .B(n2395), .C(n3957), .D(n2394), .Z(n992) );
  CENX2 U4232 ( .A(n3701), .B(n1278), .Z(n1247) );
  CENX2 U4233 ( .A(n1253), .B(n1251), .Z(n3701) );
  CEO3X1 U4234 ( .A(n2139), .B(n2170), .C(n1578), .Z(n1555) );
  CND2XL U4235 ( .A(n2139), .B(n1578), .Z(n3702) );
  CND2XL U4236 ( .A(n2139), .B(n2170), .Z(n3703) );
  CND2XL U4237 ( .A(n1578), .B(n2170), .Z(n3704) );
  CND3X1 U4238 ( .A(n3702), .B(n3703), .C(n3704), .Z(n1554) );
  COND2XL U4239 ( .A(n27), .B(n2697), .C(n2696), .D(net18545), .Z(n2170) );
  CHA1XL U4240 ( .A(n1730), .B(n1956), .CO(n1578), .S(n1579) );
  CND2X4 U4241 ( .A(n3057), .B(net16617), .Z(n3705) );
  CND2X1 U4242 ( .A(n1314), .B(n3221), .Z(n3709) );
  CND3X2 U4243 ( .A(n3707), .B(n3708), .C(n3709), .Z(n1280) );
  CIVX8 U4244 ( .A(net16670), .Z(net16671) );
  CND2XL U4245 ( .A(n414), .B(n3142), .Z(n394) );
  CND2XL U4246 ( .A(n414), .B(n748), .Z(n405) );
  CNR2X2 U4247 ( .A(n440), .B(net19689), .Z(n414) );
  CIVXL U4248 ( .A(n510), .Z(net19358) );
  CND2X2 U4249 ( .A(n957), .B(n974), .Z(n434) );
  CENXL U4250 ( .A(n3987), .B(n4001), .Z(n2765) );
  CENXL U4251 ( .A(n2794), .B(n4001), .Z(n2761) );
  CENXL U4252 ( .A(n3988), .B(n4001), .Z(n2764) );
  CENXL U4253 ( .A(n2793), .B(n4001), .Z(n2760) );
  CND3X2 U4254 ( .A(net18830), .B(n3874), .C(net18832), .Z(n1194) );
  COND2X1 U4255 ( .A(n27), .B(n2705), .C(net18546), .D(n2704), .Z(n2178) );
  COAN1X1 U4256 ( .A(n458), .B(n448), .C(n449), .Z(n445) );
  CND2XL U4257 ( .A(n3354), .B(n2188), .Z(n3724) );
  COND2X1 U4258 ( .A(n27), .B(n2694), .C(net18546), .D(n2693), .Z(n2167) );
  CNR2X1 U4259 ( .A(n1361), .B(n1386), .Z(n572) );
  CENX1 U4260 ( .A(n3713), .B(net19184), .Z(n1159) );
  CND2X1 U4261 ( .A(n3808), .B(n3807), .Z(n3713) );
  CND2X1 U4262 ( .A(n1345), .B(n1370), .Z(n3715) );
  CND2X1 U4263 ( .A(n1345), .B(n1347), .Z(n3716) );
  CND3X2 U4264 ( .A(n3715), .B(n3716), .C(n3717), .Z(n1338) );
  CND2X1 U4265 ( .A(net15999), .B(n3718), .Z(n3719) );
  CND2X2 U4266 ( .A(net19319), .B(a[18]), .Z(n3720) );
  CND2X2 U4267 ( .A(n3719), .B(n3720), .Z(n2818) );
  CEOX2 U4268 ( .A(n3879), .B(n3034), .Z(n1309) );
  CEOX1 U4269 ( .A(n3767), .B(n1348), .Z(n1315) );
  CNIVX4 U4270 ( .A(n2780), .Z(n3996) );
  CENX1 U4271 ( .A(n3996), .B(n4000), .Z(n2747) );
  CENXL U4272 ( .A(n3994), .B(net19845), .Z(n2456) );
  CND2XL U4273 ( .A(n3085), .B(n2164), .Z(n3721) );
  CND2XL U4274 ( .A(n1979), .B(n2164), .Z(n3722) );
  CND2XL U4275 ( .A(n1979), .B(n3025), .Z(n3723) );
  CND3X1 U4276 ( .A(n3721), .B(n3722), .C(n3723), .Z(n1428) );
  COND2X1 U4277 ( .A(n27), .B(n2691), .C(net18545), .D(n2690), .Z(n2164) );
  CND3X1 U4278 ( .A(n3753), .B(n3754), .C(n3755), .Z(n1282) );
  CIVXL U4279 ( .A(n546), .Z(net19290) );
  COND2X1 U4280 ( .A(n3080), .B(n2508), .C(n3285), .D(n2507), .Z(n1982) );
  COR2X1 U4281 ( .A(n1504), .B(n1483), .Z(net19288) );
  CND2X1 U4282 ( .A(n1461), .B(n1482), .Z(n606) );
  CNR2X1 U4283 ( .A(n1461), .B(n1482), .Z(n605) );
  CNR2X1 U4284 ( .A(n636), .B(n3596), .Z(n631) );
  CIVXL U4285 ( .A(n1767), .Z(n3727) );
  CIVX1 U4286 ( .A(n3727), .Z(n3728) );
  CAOR1XL U4287 ( .A(n3832), .B(n3904), .C(n2615), .Z(n2088) );
  COND2XL U4288 ( .A(n3904), .B(n2641), .C(n2640), .D(n3833), .Z(n2114) );
  COND2XL U4289 ( .A(n3904), .B(n2628), .C(n3832), .D(n2627), .Z(n2101) );
  COND2XL U4290 ( .A(n3904), .B(n2632), .C(n3833), .D(n2631), .Z(n2105) );
  CND2XL U4291 ( .A(n1128), .B(n2028), .Z(n3730) );
  CND2XL U4292 ( .A(n1128), .B(n2121), .Z(n3731) );
  CND2XL U4293 ( .A(n2028), .B(n2121), .Z(n3732) );
  CND3X1 U4294 ( .A(n3730), .B(n3731), .C(n3732), .Z(n1096) );
  CNR2X2 U4295 ( .A(n3909), .B(n1304), .Z(n551) );
  CEOX1 U4296 ( .A(n1315), .B(n1340), .Z(n3879) );
  CIVXL U4297 ( .A(n3306), .Z(n399) );
  CND3X2 U4298 ( .A(n3890), .B(n3891), .C(n3892), .Z(n1190) );
  CENXL U4299 ( .A(n2792), .B(n3999), .Z(n2759) );
  CENXL U4300 ( .A(n2784), .B(n3999), .Z(n2751) );
  CENXL U4301 ( .A(n2789), .B(n3999), .Z(n2756) );
  CENXL U4302 ( .A(n3991), .B(n3999), .Z(n2757) );
  CENXL U4303 ( .A(n2783), .B(n3999), .Z(n2750) );
  CENXL U4304 ( .A(n2782), .B(n3999), .Z(n2749) );
  CENXL U4305 ( .A(n2794), .B(n3930), .Z(n2662) );
  CENXL U4306 ( .A(n3986), .B(n3930), .Z(n2667) );
  CENXL U4307 ( .A(n2806), .B(n3930), .Z(n2674) );
  CENXL U4308 ( .A(n3990), .B(n3930), .Z(n2663) );
  CENXL U4309 ( .A(n3984), .B(n3930), .Z(n2678) );
  CENXL U4310 ( .A(n3985), .B(n3930), .Z(n2671) );
  CENXL U4311 ( .A(n2793), .B(n3930), .Z(n2661) );
  COND2XL U4312 ( .A(n36), .B(n2672), .C(n3425), .D(n2671), .Z(n2145) );
  CIVX4 U4313 ( .A(n3981), .Z(n51) );
  CNR2XL U4314 ( .A(n1387), .B(n1412), .Z(n3734) );
  CENX2 U4315 ( .A(n1250), .B(n1221), .Z(n3805) );
  CNR2IX1 U4316 ( .B(n3998), .A(net16623), .Z(n1833) );
  COND2XL U4317 ( .A(n36), .B(n2678), .C(n3655), .D(n2677), .Z(n2151) );
  CND2X1 U4318 ( .A(n4015), .B(n3736), .Z(n3737) );
  CND2X2 U4319 ( .A(n3735), .B(n3487), .Z(n3738) );
  CEOX1 U4320 ( .A(n1343), .B(n1368), .Z(n3777) );
  CEO3X2 U4321 ( .A(n1283), .B(n1281), .C(n1308), .Z(n3900) );
  CIVX2 U4322 ( .A(net16580), .Z(net16001) );
  CEO3X2 U4323 ( .A(n1254), .B(n1229), .C(n3029), .Z(n1221) );
  CND2XL U4324 ( .A(n1254), .B(n1229), .Z(n3740) );
  CND2X1 U4325 ( .A(n1227), .B(n1229), .Z(n3741) );
  COND2X1 U4326 ( .A(n2563), .B(n3916), .C(n3355), .D(n2562), .Z(n2036) );
  COND2X1 U4327 ( .A(n2649), .B(n3424), .C(n2650), .D(n3163), .Z(n2123) );
  COND2XL U4328 ( .A(n2679), .B(n3163), .C(n3425), .D(n2678), .Z(n2152) );
  CND2XL U4329 ( .A(net21540), .B(n2125), .Z(n3847) );
  CND2XL U4330 ( .A(n1387), .B(n1412), .Z(n583) );
  CENXL U4331 ( .A(n2804), .B(net16023), .Z(n3742) );
  CND2XL U4332 ( .A(n1223), .B(n1225), .Z(n3745) );
  COND2X2 U4333 ( .A(n27), .B(n2698), .C(n2697), .D(net18545), .Z(n2171) );
  CENX1 U4334 ( .A(net16399), .B(net16549), .Z(n2574) );
  CNR2X1 U4335 ( .A(n693), .B(n696), .Z(n691) );
  CIVXL U4336 ( .A(n693), .Z(n784) );
  CND2X4 U4337 ( .A(n2816), .B(n3958), .Z(n3747) );
  COND2X2 U4338 ( .A(n2748), .B(n9), .C(n6), .D(n2747), .Z(n2221) );
  CIVXL U4339 ( .A(n474), .Z(n3748) );
  CNIVX4 U4340 ( .A(net21614), .Z(net19200) );
  COND2XL U4341 ( .A(n3080), .B(n2490), .C(n3285), .D(n2489), .Z(n1965) );
  COND2XL U4342 ( .A(n2484), .B(n3080), .C(n3285), .D(n2483), .Z(n1959) );
  COND2X1 U4343 ( .A(n81), .B(n2500), .C(n2499), .D(net18902), .Z(n1974) );
  CENXL U4344 ( .A(n2791), .B(n3476), .Z(n2329) );
  CENXL U4345 ( .A(n2781), .B(n4020), .Z(n2319) );
  CENXL U4346 ( .A(n3991), .B(n3475), .Z(n2328) );
  CENXL U4347 ( .A(n2789), .B(n3476), .Z(n2327) );
  CENXL U4348 ( .A(n3994), .B(n3476), .Z(n2324) );
  CENXL U4349 ( .A(n2784), .B(n4020), .Z(n2322) );
  CENXL U4350 ( .A(n2792), .B(n3476), .Z(n2330) );
  CENXL U4351 ( .A(n3992), .B(n3475), .Z(n2326) );
  CENXL U4352 ( .A(n2804), .B(n3475), .Z(n2342) );
  CENXL U4353 ( .A(n2794), .B(n3476), .Z(n2332) );
  CENXL U4354 ( .A(n3989), .B(n4021), .Z(n2334) );
  CENXL U4355 ( .A(n2793), .B(n4020), .Z(n2331) );
  CND3X2 U4356 ( .A(n3768), .B(n3769), .C(n3770), .Z(n1314) );
  CIVX4 U4357 ( .A(n120), .Z(n4022) );
  CIVX2 U4358 ( .A(n84), .Z(net16005) );
  CND2X4 U4359 ( .A(n2822), .B(n3733), .Z(n54) );
  CENX1 U4360 ( .A(n3798), .B(n1121), .Z(n1115) );
  CENX1 U4361 ( .A(n1125), .B(n1146), .Z(n3798) );
  COND2X1 U4362 ( .A(n2451), .B(net22025), .C(net19996), .D(n2450), .Z(n1928)
         );
  CIVXL U4363 ( .A(n1161), .Z(net19184) );
  CND2XL U4364 ( .A(n1040), .B(n3370), .Z(n3750) );
  CND2XL U4365 ( .A(n1021), .B(n1042), .Z(n3752) );
  CND3X1 U4366 ( .A(n3750), .B(n3751), .C(n3752), .Z(n1016) );
  CNR2IX1 U4367 ( .B(n3998), .A(n3267), .Z(n2087) );
  CIVX4 U4368 ( .A(net15999), .Z(net16670) );
  CENX1 U4369 ( .A(net16403), .B(net16671), .Z(n2477) );
  COND2X1 U4370 ( .A(n3705), .B(n2264), .C(net16617), .D(n2263), .Z(n1750) );
  CANR1X2 U4371 ( .A(n349), .B(n3946), .C(n340), .Z(n334) );
  CIVX1 U4372 ( .A(n351), .Z(n349) );
  CND2IXL U4373 ( .B(n3998), .A(n4004), .Z(n2746) );
  CENXL U4374 ( .A(n2794), .B(n4004), .Z(n2728) );
  CENXL U4375 ( .A(n2793), .B(n4003), .Z(n2727) );
  COND2X1 U4376 ( .A(n3340), .B(n2532), .C(net16683), .D(n2531), .Z(n2005) );
  COND2X1 U4377 ( .A(n54), .B(n2598), .C(n3733), .D(n2597), .Z(n2071) );
  CNR2IX1 U4378 ( .B(n3998), .A(net16606), .Z(n1863) );
  CENXL U4379 ( .A(n2781), .B(net22026), .Z(n2286) );
  CENXL U4380 ( .A(n3993), .B(net22026), .Z(n2292) );
  CENXL U4381 ( .A(n3992), .B(net22026), .Z(n2293) );
  CENXL U4382 ( .A(n2791), .B(net18407), .Z(n2296) );
  CENXL U4383 ( .A(n3986), .B(net18407), .Z(n2304) );
  CENXL U4384 ( .A(n2794), .B(net18407), .Z(n2299) );
  CENXL U4385 ( .A(n2804), .B(net18407), .Z(n2309) );
  CNR2X2 U4386 ( .A(n1713), .B(n1716), .Z(n708) );
  COND1X1 U4387 ( .A(n666), .B(n660), .C(n661), .Z(n659) );
  CIVXL U4388 ( .A(n666), .Z(n664) );
  CNR2X2 U4389 ( .A(n511), .B(net18745), .Z(n498) );
  CEO3X2 U4390 ( .A(n1316), .B(n1318), .C(n1291), .Z(n1283) );
  CND2XL U4391 ( .A(n1316), .B(n1291), .Z(n3753) );
  CND2XL U4392 ( .A(n1316), .B(n1318), .Z(n3754) );
  CND2X1 U4393 ( .A(n1291), .B(n1318), .Z(n3755) );
  CEO3X1 U4394 ( .A(n2237), .B(n2144), .C(n1732), .Z(n1637) );
  CND2XL U4395 ( .A(n2237), .B(n2144), .Z(n3756) );
  CND2XL U4396 ( .A(n2237), .B(n1732), .Z(n3757) );
  CND2XL U4397 ( .A(n2144), .B(n1732), .Z(n3758) );
  CND3X1 U4398 ( .A(n3756), .B(n3757), .C(n3758), .Z(n1636) );
  CND2XL U4399 ( .A(n1638), .B(n1634), .Z(n3759) );
  CND3X1 U4400 ( .A(n3759), .B(n3760), .C(n3761), .Z(n1618) );
  COR2XL U4401 ( .A(n2548), .B(net16683), .Z(n3762) );
  CND2X1 U4402 ( .A(net19162), .B(n3762), .Z(n1732) );
  CND2IXL U4403 ( .B(n3998), .A(n3167), .Z(n2548) );
  CEOX2 U4404 ( .A(n3763), .B(n1507), .Z(n1505) );
  CND2XL U4405 ( .A(n1507), .B(n1526), .Z(n3764) );
  CND2XL U4406 ( .A(n1507), .B(n1509), .Z(n3765) );
  CND3X2 U4407 ( .A(n3842), .B(n3843), .C(n3844), .Z(n1136) );
  CND2X1 U4408 ( .A(n1143), .B(n1141), .Z(n3842) );
  CND2X4 U4409 ( .A(n2813), .B(n132), .Z(n3915) );
  CEOX2 U4410 ( .A(n1323), .B(n1325), .Z(n3767) );
  CND2X1 U4411 ( .A(n1348), .B(n1325), .Z(n3768) );
  CND2X1 U4412 ( .A(n1348), .B(n1323), .Z(n3769) );
  CIVX4 U4413 ( .A(net16539), .Z(net16023) );
  CEO3X2 U4414 ( .A(n1313), .B(n1336), .C(n1311), .Z(n1307) );
  CND2XL U4415 ( .A(n1313), .B(n1336), .Z(n3771) );
  CND2X1 U4416 ( .A(n1313), .B(n1311), .Z(n3772) );
  CND2X1 U4417 ( .A(n1336), .B(n1311), .Z(n3773) );
  CND3X2 U4418 ( .A(n3771), .B(n3772), .C(n3773), .Z(n1306) );
  CND2XL U4419 ( .A(n1309), .B(n1334), .Z(n3774) );
  CND2X1 U4420 ( .A(n1309), .B(n1307), .Z(n3775) );
  CND2X1 U4421 ( .A(n1334), .B(n1307), .Z(n3776) );
  CND3X2 U4422 ( .A(n3774), .B(n3775), .C(n3776), .Z(n1304) );
  CND2X1 U4423 ( .A(n1366), .B(n1368), .Z(n3778) );
  CND2X1 U4424 ( .A(n1366), .B(n1343), .Z(n3779) );
  CND2XL U4425 ( .A(n1368), .B(n1343), .Z(n3780) );
  CND3X2 U4426 ( .A(n3778), .B(n3779), .C(n3780), .Z(n1336) );
  COR2XL U4427 ( .A(n1360), .B(n1333), .Z(n3781) );
  CEO3X2 U4428 ( .A(n1442), .B(n1419), .C(n1440), .Z(n1415) );
  CEOX2 U4429 ( .A(n1415), .B(n3782), .Z(n1413) );
  CND2X1 U4430 ( .A(n1442), .B(n1419), .Z(n3783) );
  CND2XL U4431 ( .A(n1438), .B(n1417), .Z(n3786) );
  CND2XL U4432 ( .A(n1417), .B(n1415), .Z(n3787) );
  CND2XL U4433 ( .A(n1438), .B(n1415), .Z(n3788) );
  CND2XL U4434 ( .A(n1453), .B(n1457), .Z(n3789) );
  CND2X1 U4435 ( .A(n1453), .B(n1455), .Z(n3790) );
  CND2X1 U4436 ( .A(n1457), .B(n1455), .Z(n3791) );
  CND3X2 U4437 ( .A(n3789), .B(n3790), .C(n3791), .Z(n1444) );
  CIVX2 U4438 ( .A(n472), .Z(n474) );
  CENXL U4439 ( .A(n2793), .B(n3357), .Z(n2694) );
  CENXL U4440 ( .A(n3988), .B(n4006), .Z(n2698) );
  CENXL U4441 ( .A(n2794), .B(n3357), .Z(n2695) );
  CIVX1 U4442 ( .A(n2133), .Z(n3793) );
  CIVX2 U4443 ( .A(n3793), .Z(n3794) );
  CND2XL U4444 ( .A(n784), .B(n694), .Z(n202) );
  CND2XL U4445 ( .A(net18274), .B(net19362), .Z(n193) );
  COND2X1 U4446 ( .A(n3059), .B(n2561), .C(n3037), .D(n2560), .Z(n2034) );
  CNIVX4 U4447 ( .A(n2786), .Z(n3994) );
  COND2X1 U4448 ( .A(n2520), .B(n3044), .C(net16684), .D(n2519), .Z(n1994) );
  CAOR1XL U4449 ( .A(n3432), .B(n3352), .C(n2582), .Z(n2055) );
  CENXL U4450 ( .A(n2784), .B(net18510), .Z(n2520) );
  CIVXL U4451 ( .A(n2143), .Z(n3796) );
  CIVX1 U4452 ( .A(n3796), .Z(n3797) );
  CNR2IX1 U4453 ( .B(n3998), .A(n3957), .Z(n1894) );
  CENX1 U4454 ( .A(n1265), .B(n1271), .Z(n3902) );
  CENXL U4455 ( .A(n3996), .B(n4020), .Z(n2318) );
  CENXL U4456 ( .A(net16389), .B(n3475), .Z(n2338) );
  CENXL U4457 ( .A(net16391), .B(n4020), .Z(n2339) );
  CENXL U4458 ( .A(n3986), .B(n3475), .Z(n2337) );
  CENXL U4459 ( .A(net16393), .B(n4020), .Z(n2340) );
  CENXL U4460 ( .A(n3985), .B(n3475), .Z(n2341) );
  CENXL U4461 ( .A(net16407), .B(n3476), .Z(n2347) );
  CENXL U4462 ( .A(n2806), .B(n3475), .Z(n2344) );
  CENX4 U4463 ( .A(a[28]), .B(n4021), .Z(n132) );
  CND3X1 U4464 ( .A(n3875), .B(n3876), .C(n3877), .Z(n1328) );
  CIVXL U4465 ( .A(n559), .Z(n3800) );
  CIVXL U4466 ( .A(n3800), .Z(n3801) );
  CND2X1 U4467 ( .A(n620), .B(net18280), .Z(n613) );
  COND2XL U4468 ( .A(n63), .B(n2572), .C(n3037), .D(n2571), .Z(n2045) );
  CENXL U4469 ( .A(net16403), .B(net16649), .Z(n3802) );
  CNIVX16 U4470 ( .A(net15985), .Z(net18520) );
  CENXL U4471 ( .A(n3996), .B(n4018), .Z(n2483) );
  CND2IXL U4472 ( .B(n3998), .A(n4018), .Z(n2515) );
  CENXL U4473 ( .A(n3998), .B(n4018), .Z(n2514) );
  CENXL U4474 ( .A(net16407), .B(n4018), .Z(n2512) );
  CENXL U4475 ( .A(net16399), .B(n4018), .Z(n2508) );
  CENXL U4476 ( .A(net16391), .B(n4018), .Z(n2504) );
  CENXL U4477 ( .A(n3984), .B(n4018), .Z(n2513) );
  CENXL U4478 ( .A(n3987), .B(n4018), .Z(n2501) );
  CENXL U4479 ( .A(n3988), .B(n4018), .Z(n2500) );
  CENXL U4480 ( .A(n3986), .B(n4018), .Z(n2502) );
  CENXL U4481 ( .A(n3990), .B(n4018), .Z(n2498) );
  CENXL U4482 ( .A(n3985), .B(n4018), .Z(n2506) );
  CENXL U4483 ( .A(n2808), .B(n4018), .Z(n2511) );
  CENXL U4484 ( .A(net16389), .B(n4018), .Z(n2503) );
  CENXL U4485 ( .A(n2781), .B(net16001), .Z(n2451) );
  CENXL U4486 ( .A(n2784), .B(net16001), .Z(n2454) );
  CENXL U4487 ( .A(n2792), .B(net16001), .Z(n2462) );
  CENXL U4488 ( .A(n3992), .B(net15999), .Z(n2458) );
  CENXL U4489 ( .A(n2783), .B(net16001), .Z(n2453) );
  CENXL U4490 ( .A(n3993), .B(net16001), .Z(n2457) );
  CENXL U4491 ( .A(n3995), .B(net16001), .Z(n2455) );
  CENXL U4492 ( .A(n2791), .B(net16001), .Z(n2461) );
  CENXL U4493 ( .A(n2782), .B(net16001), .Z(n2452) );
  CENXL U4494 ( .A(n2804), .B(net16001), .Z(n2474) );
  CND2XL U4495 ( .A(n1121), .B(n1146), .Z(n3887) );
  COND1XL U4496 ( .A(n605), .B(n3062), .C(net18869), .Z(n604) );
  CEO3X2 U4497 ( .A(n1989), .B(n3797), .C(n3140), .Z(n1625) );
  CND2XL U4498 ( .A(n1989), .B(n3470), .Z(n3863) );
  COND2X1 U4499 ( .A(n3904), .B(n2619), .C(n42), .D(n2618), .Z(n2092) );
  CNIVX4 U4500 ( .A(n105), .Z(n3958) );
  COND2X1 U4501 ( .A(n2451), .B(net19996), .C(n2452), .D(net22025), .Z(n1929)
         );
  CAOR1XL U4502 ( .A(net19996), .B(net22025), .C(n2450), .Z(n1927) );
  COND2XL U4503 ( .A(net22025), .B(n2454), .C(net19422), .D(n2453), .Z(n1931)
         );
  CND3X1 U4504 ( .A(n3840), .B(n3839), .C(n3838), .Z(n1418) );
  CND2XL U4505 ( .A(n1448), .B(n1446), .Z(n3839) );
  CND2X1 U4506 ( .A(n1226), .B(n1228), .Z(n3874) );
  CIVXL U4507 ( .A(n3398), .Z(n3806) );
  CND2X4 U4508 ( .A(n3883), .B(net18811), .Z(n2813) );
  CND2XL U4509 ( .A(n1188), .B(net19034), .Z(n3808) );
  CIVXL U4510 ( .A(n474), .Z(n3809) );
  CND2XL U4511 ( .A(n1188), .B(n1161), .Z(n3810) );
  CND3X1 U4512 ( .A(n3810), .B(net19025), .C(net19026), .Z(n1158) );
  CEOX1 U4513 ( .A(n1914), .B(n1884), .Z(n3811) );
  CND2XL U4514 ( .A(n2003), .B(n1884), .Z(n3812) );
  CND2XL U4515 ( .A(n2003), .B(n1914), .Z(n3813) );
  CND2XL U4516 ( .A(n1884), .B(n1914), .Z(n3814) );
  CND3X1 U4517 ( .A(n3812), .B(n3813), .C(n3814), .Z(n1266) );
  COND2X1 U4518 ( .A(n3168), .B(n2382), .C(net21572), .D(n2381), .Z(n1862) );
  CND2X1 U4519 ( .A(a[12]), .B(net16539), .Z(n3816) );
  CND2X2 U4520 ( .A(n3815), .B(net19011), .Z(n3817) );
  CIVXL U4521 ( .A(a[12]), .Z(n3815) );
  CENX1 U4522 ( .A(n3986), .B(net16676), .Z(n2370) );
  CND2X1 U4523 ( .A(n3858), .B(n3859), .Z(n2682) );
  CENXL U4524 ( .A(n2804), .B(n4008), .Z(n2672) );
  CENXL U4525 ( .A(n3988), .B(n4008), .Z(n2665) );
  CENXL U4526 ( .A(n2789), .B(n4008), .Z(n2657) );
  CENXL U4527 ( .A(n3989), .B(n4008), .Z(n2664) );
  CENXL U4528 ( .A(n3992), .B(n4008), .Z(n2656) );
  CENXL U4529 ( .A(n3993), .B(n4008), .Z(n2655) );
  CENXL U4530 ( .A(n3987), .B(n4008), .Z(n2666) );
  CENXL U4531 ( .A(n3991), .B(n4008), .Z(n2658) );
  CENXL U4532 ( .A(net16393), .B(n4008), .Z(n2670) );
  CENXL U4533 ( .A(n2792), .B(n4008), .Z(n2660) );
  CNR2X2 U4534 ( .A(n3141), .B(n938), .Z(n409) );
  COND2X1 U4535 ( .A(n2517), .B(n3465), .C(n2518), .D(net18612), .Z(n1992) );
  CENXL U4536 ( .A(n2782), .B(net18510), .Z(n2518) );
  CEO3X2 U4537 ( .A(n1285), .B(n1310), .C(n1312), .Z(n1279) );
  CND2X1 U4538 ( .A(n1285), .B(n1310), .Z(n3818) );
  CND2X1 U4539 ( .A(n1285), .B(n1312), .Z(n3819) );
  CND2X1 U4540 ( .A(n1310), .B(n1312), .Z(n3820) );
  CND3X2 U4541 ( .A(n3818), .B(n3819), .C(n3820), .Z(n1278) );
  CND2XL U4542 ( .A(n1253), .B(n1251), .Z(n3821) );
  CND3X2 U4543 ( .A(n3823), .B(n3822), .C(n3821), .Z(n1246) );
  CIVX4 U4544 ( .A(n3398), .Z(n4015) );
  CIVX1 U4545 ( .A(n1444), .Z(n3825) );
  CND2XL U4546 ( .A(n1444), .B(n1446), .Z(n3840) );
  COND2XL U4547 ( .A(net20022), .B(n2699), .C(net18546), .D(n2698), .Z(n2172)
         );
  COND2XL U4548 ( .A(n27), .B(n2710), .C(net18546), .D(n2709), .Z(n2183) );
  COND2XL U4549 ( .A(n27), .B(n2700), .C(net18546), .D(n2699), .Z(n2173) );
  COND2XL U4550 ( .A(n2712), .B(n27), .C(net18546), .D(n2711), .Z(n2185) );
  COND2XL U4551 ( .A(n27), .B(n2704), .C(net18546), .D(n2703), .Z(n2177) );
  CNR2IX1 U4552 ( .B(n3998), .A(n3334), .Z(n1926) );
  CND2X1 U4553 ( .A(n3824), .B(n1444), .Z(n3827) );
  CIVXL U4554 ( .A(n1448), .Z(n3824) );
  CND2XL U4555 ( .A(n1170), .B(n1172), .Z(n3828) );
  CND3X1 U4556 ( .A(net18982), .B(n3828), .C(net18983), .Z(n1140) );
  CND2XL U4557 ( .A(n1115), .B(n1117), .Z(n3829) );
  CND2XL U4558 ( .A(n1117), .B(n1140), .Z(n3830) );
  CND2XL U4559 ( .A(n1115), .B(n1140), .Z(n3831) );
  CND3X1 U4560 ( .A(n3831), .B(n3830), .C(n3829), .Z(n1110) );
  CNR2IX1 U4561 ( .B(n3998), .A(net16617), .Z(n1770) );
  CENX2 U4562 ( .A(n3549), .B(n4008), .Z(n3833) );
  CNIVX4 U4563 ( .A(n2788), .Z(n3992) );
  CANR1X1 U4564 ( .A(n686), .B(n3948), .C(n681), .Z(n679) );
  CNIVX1 U4565 ( .A(n4007), .Z(n3933) );
  CEO3X1 U4566 ( .A(n1476), .B(n1451), .C(n1474), .Z(n1447) );
  CND2X1 U4567 ( .A(n1476), .B(n1474), .Z(n3835) );
  CEOX2 U4568 ( .A(n3837), .B(n1446), .Z(n1419) );
  CND3X1 U4569 ( .A(net18951), .B(net18952), .C(net18953), .Z(n1166) );
  CEOX2 U4570 ( .A(n1143), .B(n1141), .Z(n3841) );
  CEOX2 U4571 ( .A(n3841), .B(n1166), .Z(n1137) );
  CND2X1 U4572 ( .A(n1143), .B(n1166), .Z(n3843) );
  CND2X1 U4573 ( .A(n1141), .B(n1166), .Z(n3844) );
  CND2XL U4574 ( .A(n1941), .B(n2125), .Z(n3846) );
  CND3X1 U4575 ( .A(n3845), .B(n3846), .C(n3847), .Z(n1204) );
  COND2X1 U4576 ( .A(n2576), .B(n63), .C(n3355), .D(n2575), .Z(n2049) );
  CENXL U4577 ( .A(n3991), .B(n4011), .Z(n2625) );
  CAN2X2 U4578 ( .A(n3917), .B(n3973), .Z(n3955) );
  COND2X1 U4579 ( .A(n3163), .B(n2671), .C(n3482), .D(n2670), .Z(n2144) );
  CIVX1 U4580 ( .A(n511), .Z(n758) );
  COND2X1 U4581 ( .A(n3044), .B(n2522), .C(net16684), .D(n2521), .Z(n1996) );
  CIVX1 U4582 ( .A(n3157), .Z(n4013) );
  CIVX3 U4583 ( .A(n3157), .Z(n4012) );
  CNIVX4 U4584 ( .A(n2803), .Z(n3985) );
  COND2XL U4585 ( .A(n3058), .B(n2555), .C(n3037), .D(n2554), .Z(n2028) );
  COND2XL U4586 ( .A(n63), .B(n2570), .C(n3355), .D(n2569), .Z(n2043) );
  COND2XL U4587 ( .A(n63), .B(n3742), .C(n3355), .D(n2572), .Z(n2046) );
  CIVX3 U4588 ( .A(n3), .Z(n4002) );
  CND2X4 U4589 ( .A(n2827), .B(n6), .Z(n3905) );
  CND2IXL U4590 ( .B(n3998), .A(n3348), .Z(n2713) );
  COND2X1 U4591 ( .A(n27), .B(n2692), .C(net18546), .D(n2691), .Z(n2165) );
  COND2X1 U4592 ( .A(n2693), .B(n27), .C(net18545), .D(n2692), .Z(n2166) );
  CENXL U4593 ( .A(n3990), .B(n3357), .Z(n2696) );
  COND2X1 U4594 ( .A(n3044), .B(n2538), .C(net16684), .D(n2537), .Z(n2011) );
  CIVX1 U4595 ( .A(net21583), .Z(n441) );
  CNR2X2 U4596 ( .A(n572), .B(n567), .Z(n561) );
  CEO3X2 U4597 ( .A(n1403), .B(n3804), .C(n1409), .Z(n1397) );
  CND2X1 U4598 ( .A(n1403), .B(n1409), .Z(n3848) );
  CND2XL U4599 ( .A(n1403), .B(n1426), .Z(n3849) );
  CND2X1 U4600 ( .A(n1409), .B(n1426), .Z(n3850) );
  CEO3X1 U4601 ( .A(n2132), .B(n3040), .C(n2070), .Z(n1403) );
  CND2XL U4602 ( .A(n2132), .B(n2070), .Z(n3851) );
  CND2XL U4603 ( .A(n2132), .B(n1978), .Z(n3852) );
  CND2X1 U4604 ( .A(n2070), .B(n1978), .Z(n3853) );
  CND3X1 U4605 ( .A(n3851), .B(n3852), .C(n3853), .Z(n1402) );
  COND2X1 U4606 ( .A(n3163), .B(n2659), .C(n3424), .D(n2658), .Z(n2132) );
  COND2X1 U4607 ( .A(n3044), .B(n2519), .C(net16684), .D(n2518), .Z(n1993) );
  CND2X4 U4608 ( .A(n2813), .B(n132), .Z(net18573) );
  CENXL U4609 ( .A(n3991), .B(n4015), .Z(n2592) );
  CENX1 U4610 ( .A(n2791), .B(n3956), .Z(n2692) );
  COND2X1 U4611 ( .A(net18570), .B(n2266), .C(net16617), .D(n2265), .Z(n1752)
         );
  COND1X1 U4612 ( .A(n480), .B(net18906), .C(net22007), .Z(n3855) );
  CND2XL U4613 ( .A(n2781), .B(n3956), .Z(n3858) );
  CND2X1 U4614 ( .A(n3856), .B(n3857), .Z(n3859) );
  CIVXL U4615 ( .A(n2781), .Z(n3856) );
  CND2XL U4616 ( .A(n2050), .B(n1989), .Z(n3861) );
  CND2XL U4617 ( .A(n2050), .B(n3470), .Z(n3862) );
  CND3X1 U4618 ( .A(n3861), .B(n3862), .C(n3863), .Z(n1624) );
  CND2X2 U4619 ( .A(net18509), .B(net18734), .Z(n3896) );
  CND2XL U4620 ( .A(n1245), .B(n1274), .Z(n3865) );
  COND2XL U4621 ( .A(n3904), .B(n2631), .C(n3833), .D(n2630), .Z(n2104) );
  CIVX2 U4622 ( .A(n30), .Z(n4010) );
  COND2XL U4623 ( .A(n2660), .B(n36), .C(n3425), .D(n2659), .Z(n2133) );
  CAOR1XL U4624 ( .A(n3424), .B(n3163), .C(n2648), .Z(n2121) );
  COND2X1 U4625 ( .A(n3163), .B(n2661), .C(n3424), .D(n2660), .Z(n2134) );
  CND2X2 U4626 ( .A(net18455), .B(n3923), .Z(n105) );
  CND2X1 U4627 ( .A(n1613), .B(n1626), .Z(n661) );
  CIVXL U4628 ( .A(n606), .Z(net18868) );
  CIVXL U4629 ( .A(net18868), .Z(net18869) );
  CENXL U4630 ( .A(n574), .B(n184), .Z(product[28]) );
  CANR1XL U4631 ( .A(n766), .B(n574), .C(n571), .Z(n569) );
  CND2XL U4632 ( .A(n3027), .B(n1063), .Z(n3866) );
  CEO3X2 U4633 ( .A(n1131), .B(n1154), .C(n1156), .Z(n1121) );
  CND2XL U4634 ( .A(n1131), .B(n1154), .Z(n3867) );
  CND2X1 U4635 ( .A(n1131), .B(n1156), .Z(n3868) );
  CND2XL U4636 ( .A(n1154), .B(n1156), .Z(n3869) );
  CND3X1 U4637 ( .A(n3867), .B(n3868), .C(n3869), .Z(n1120) );
  CND2XL U4638 ( .A(n1101), .B(n1118), .Z(n3870) );
  CND2X1 U4639 ( .A(n1101), .B(n1120), .Z(n3871) );
  CND2XL U4640 ( .A(n1118), .B(n1120), .Z(n3872) );
  CND3X1 U4641 ( .A(n3872), .B(n3871), .C(n3870), .Z(n1090) );
  CIVXL U4642 ( .A(n356), .Z(net18839) );
  COND2X1 U4643 ( .A(n3044), .B(n2542), .C(net16683), .D(n2541), .Z(n2015) );
  CND2X1 U4644 ( .A(n3878), .B(n1800), .Z(n3875) );
  CND2XL U4645 ( .A(n3878), .B(n2222), .Z(n3876) );
  COND2XL U4646 ( .A(n3044), .B(n2532), .C(net16684), .D(n2531), .Z(n3878) );
  CND2X1 U4647 ( .A(n1338), .B(n1340), .Z(n3880) );
  CND2X1 U4648 ( .A(n1338), .B(n1315), .Z(n3881) );
  CND2X1 U4649 ( .A(n1340), .B(n1315), .Z(n3882) );
  CND3X2 U4650 ( .A(n3880), .B(n3881), .C(n3882), .Z(n1308) );
  CND2X1 U4651 ( .A(n1221), .B(n1248), .Z(n3884) );
  CND2X1 U4652 ( .A(n1248), .B(n1250), .Z(n3885) );
  CND3X2 U4653 ( .A(n3884), .B(n3885), .C(n3886), .Z(n1216) );
  CENX1 U4654 ( .A(n2806), .B(net16676), .Z(n2377) );
  CENX1 U4655 ( .A(net16399), .B(net16676), .Z(n2376) );
  CND2X1 U4656 ( .A(n1121), .B(n1125), .Z(n3888) );
  CND2XL U4657 ( .A(n1146), .B(n1125), .Z(n3889) );
  CND3X1 U4658 ( .A(n3887), .B(n3888), .C(n3889), .Z(n1114) );
  CNIVX2 U4659 ( .A(n1725), .Z(n3917) );
  COND2X1 U4660 ( .A(n3163), .B(n2668), .C(n3655), .D(n2667), .Z(n2141) );
  COND1X1 U4661 ( .A(n405), .B(n149), .C(n406), .Z(n404) );
  COND1XL U4662 ( .A(n460), .B(n3922), .C(n3919), .Z(n459) );
  CENXL U4663 ( .A(n3985), .B(n3167), .Z(n2539) );
  CENXL U4664 ( .A(net16393), .B(n3166), .Z(n2538) );
  CENXL U4665 ( .A(n3996), .B(n3167), .Z(n2516) );
  CENXL U4666 ( .A(net16399), .B(n3167), .Z(n2541) );
  CENXL U4667 ( .A(n2806), .B(n3166), .Z(n2542) );
  CENXL U4668 ( .A(net16391), .B(net18492), .Z(n2537) );
  CND2X1 U4669 ( .A(n1195), .B(n1222), .Z(n3890) );
  CIVXL U4670 ( .A(n501), .Z(net18744) );
  CND2X1 U4671 ( .A(n1223), .B(n1252), .Z(n3893) );
  CND2X1 U4672 ( .A(n1223), .B(n1225), .Z(n3894) );
  CND2X1 U4673 ( .A(n1252), .B(n1225), .Z(n3895) );
  CND3X2 U4674 ( .A(n3893), .B(n3895), .C(n3894), .Z(n1218) );
  CNIVX2 U4675 ( .A(net16015), .Z(net18509) );
  CENX2 U4676 ( .A(a[12]), .B(n4016), .Z(n3935) );
  CENXL U4677 ( .A(n3898), .B(n149), .Z(product[40]) );
  CAN2XL U4678 ( .A(n754), .B(n3748), .Z(n3898) );
  CENXL U4679 ( .A(n2791), .B(n4003), .Z(n2725) );
  CENXL U4680 ( .A(n3991), .B(n4003), .Z(n2724) );
  CENXL U4681 ( .A(n2792), .B(n4003), .Z(n2726) );
  CENXL U4682 ( .A(n3993), .B(n4003), .Z(n2721) );
  CENXL U4683 ( .A(n3994), .B(n4003), .Z(n2720) );
  CENXL U4684 ( .A(n2782), .B(n4003), .Z(n2716) );
  CENXL U4685 ( .A(n2789), .B(n4003), .Z(n2723) );
  CENXL U4686 ( .A(n3995), .B(n4003), .Z(n2719) );
  CENXL U4687 ( .A(n2784), .B(n4003), .Z(n2718) );
  CENXL U4688 ( .A(n2781), .B(n4003), .Z(n2715) );
  CIVXL U4689 ( .A(n764), .Z(n3899) );
  CIVXL U4690 ( .A(n3873), .Z(n764) );
  CENXL U4691 ( .A(n3996), .B(net18520), .Z(n2384) );
  CENXL U4692 ( .A(n2806), .B(net19890), .Z(n2410) );
  CENXL U4693 ( .A(net16399), .B(net18944), .Z(n2409) );
  CIVXL U4694 ( .A(n18), .Z(net18703) );
  CIVXL U4695 ( .A(n592), .Z(n590) );
  COND1XL U4696 ( .A(n298), .B(n3922), .C(n299), .Z(n297) );
  COND2X1 U4697 ( .A(n126), .B(n3910), .C(net16623), .D(n2350), .Z(n1726) );
  CHA1X1 U4698 ( .A(n1726), .B(n1832), .CO(n1410), .S(n1411) );
  CENXL U4699 ( .A(n2793), .B(n3806), .Z(n2595) );
  CENXL U4700 ( .A(n426), .B(n167), .Z(product[45]) );
  CIVXL U4701 ( .A(n223), .Z(n221) );
  COND1XL U4702 ( .A(n381), .B(n3922), .C(n382), .Z(n380) );
  CENXL U4703 ( .A(n459), .B(n170), .Z(product[42]) );
  CENXL U4704 ( .A(n380), .B(n163), .Z(product[49]) );
  COND2X1 U4705 ( .A(n90), .B(n2464), .C(net19996), .D(n2463), .Z(n1939) );
  COND1XL U4706 ( .A(n220), .B(n3922), .C(n221), .Z(n219) );
  COND1XL U4707 ( .A(n344), .B(n3922), .C(n345), .Z(n343) );
  CENXL U4708 ( .A(n404), .B(n165), .Z(product[47]) );
  CENXL U4709 ( .A(n3986), .B(n3961), .Z(n2601) );
  CENXL U4710 ( .A(n3985), .B(n3961), .Z(n2605) );
  CENXL U4711 ( .A(net16393), .B(n3961), .Z(n2604) );
  CENXL U4712 ( .A(net16389), .B(n3961), .Z(n2602) );
  CENXL U4713 ( .A(net16391), .B(n3961), .Z(n2603) );
  CENXL U4714 ( .A(n3984), .B(n3961), .Z(n2612) );
  CFA1X1 U4715 ( .A(n1905), .B(n1845), .CI(n1788), .CO(n1010), .S(n1011) );
  CIVX1 U4716 ( .A(n1130), .Z(n1131) );
  CEO3X1 U4717 ( .A(n1279), .B(n1306), .C(n1277), .Z(n3909) );
  CENXL U4718 ( .A(n3984), .B(net16671), .Z(n2480) );
  COND1X1 U4719 ( .A(n628), .B(n622), .C(n623), .Z(n621) );
  CNR2X2 U4720 ( .A(n1505), .B(n1524), .Z(n622) );
  CNIVX4 U4721 ( .A(n2790), .Z(n3991) );
  COND1XL U4722 ( .A(n224), .B(net19414), .C(n225), .Z(n223) );
  CIVXL U4723 ( .A(n260), .Z(n258) );
  COND2XL U4724 ( .A(n3912), .B(n2595), .C(n3267), .D(n2594), .Z(n2068) );
  CENXL U4725 ( .A(n343), .B(n160), .Z(product[52]) );
  CAOR1XL U4726 ( .A(net16617), .B(net18570), .C(n2252), .Z(n1740) );
  COND2XL U4727 ( .A(n2253), .B(net16617), .C(n2254), .D(n3705), .Z(n1741) );
  COND2XL U4728 ( .A(n3705), .B(n2256), .C(net16617), .D(n2255), .Z(n1742) );
  COND2XL U4729 ( .A(n3705), .B(n2258), .C(net16617), .D(n2257), .Z(n1744) );
  COND2XL U4730 ( .A(n3705), .B(n2262), .C(net16617), .D(n2261), .Z(n1748) );
  COND2XL U4731 ( .A(net18570), .B(n2259), .C(net16617), .D(n2258), .Z(n1745)
         );
  CIVXL U4732 ( .A(net16554), .Z(n763) );
  CNR2X2 U4733 ( .A(n1275), .B(n1304), .Z(net16554) );
  CIVX1 U4734 ( .A(n384), .Z(n382) );
  COND1X1 U4735 ( .A(n385), .B(n441), .C(n386), .Z(n384) );
  CIVXL U4736 ( .A(net18827), .Z(n597) );
  CENXL U4737 ( .A(n3997), .B(n4004), .Z(n2745) );
  CENXL U4738 ( .A(n3997), .B(n4008), .Z(n2679) );
  CENXL U4739 ( .A(n3997), .B(net16645), .Z(n2547) );
  CENXL U4740 ( .A(n3997), .B(net16671), .Z(n2481) );
  CENXL U4741 ( .A(n3997), .B(net18944), .Z(n2415) );
  CENXL U4742 ( .A(n3997), .B(net16649), .Z(n2448) );
  CENXL U4743 ( .A(n3997), .B(n4020), .Z(n2349) );
  CENXL U4744 ( .A(n3997), .B(net18407), .Z(n2316) );
  CENXL U4745 ( .A(n2794), .B(n3961), .Z(n3907) );
  CENXL U4746 ( .A(n2794), .B(n3806), .Z(n2596) );
  CIVXL U4747 ( .A(n534), .Z(n532) );
  CENXL U4748 ( .A(n176), .B(n513), .Z(product[36]) );
  CND2X2 U4749 ( .A(n754), .B(n753), .Z(n460) );
  COND1X1 U4750 ( .A(n309), .B(net19414), .C(n310), .Z(n308) );
  CIVXL U4751 ( .A(n4020), .Z(n3910) );
  CENXL U4752 ( .A(n3996), .B(net16549), .Z(n2549) );
  CENXL U4753 ( .A(net16407), .B(net16549), .Z(n2578) );
  CENXL U4754 ( .A(n3985), .B(net16549), .Z(n2572) );
  CENXL U4755 ( .A(net16389), .B(net16549), .Z(n2569) );
  CENXL U4756 ( .A(net16403), .B(net16549), .Z(n2576) );
  CENXL U4757 ( .A(n3990), .B(net16027), .Z(n2564) );
  CENXL U4758 ( .A(n3988), .B(net16027), .Z(n2566) );
  CENXL U4759 ( .A(net16391), .B(net16027), .Z(n2570) );
  CENXL U4760 ( .A(net16393), .B(net16027), .Z(n2571) );
  CNR2IX1 U4761 ( .B(n3998), .A(net18772), .Z(n1802) );
  CENXL U4762 ( .A(n3996), .B(n4023), .Z(n2252) );
  CENXL U4763 ( .A(n2804), .B(n4023), .Z(n2276) );
  CENXL U4764 ( .A(net16391), .B(n4023), .Z(n2273) );
  CENXL U4765 ( .A(n3985), .B(n4023), .Z(n2275) );
  CENXL U4766 ( .A(n3986), .B(n4023), .Z(n2271) );
  CENXL U4767 ( .A(net16389), .B(n4023), .Z(n2272) );
  CENXL U4768 ( .A(n3997), .B(n4023), .Z(n2283) );
  CENXL U4769 ( .A(net16393), .B(n4023), .Z(n2274) );
  CENXL U4770 ( .A(n3984), .B(n4023), .Z(n2282) );
  CENXL U4771 ( .A(net16407), .B(n4023), .Z(n2281) );
  CENXL U4772 ( .A(net16399), .B(n4023), .Z(n2277) );
  CENXL U4773 ( .A(n2806), .B(n4023), .Z(n2278) );
  CIVX4 U4774 ( .A(n3921), .Z(n4023) );
  COND2X1 U4775 ( .A(n18), .B(n2738), .C(net16639), .D(n2737), .Z(n2211) );
  CENXL U4776 ( .A(n2804), .B(n4003), .Z(n2738) );
  CENXL U4777 ( .A(n178), .B(n531), .Z(product[34]) );
  CND2XL U4778 ( .A(net18783), .B(n756), .Z(n174) );
  CENXL U4779 ( .A(n179), .B(n542), .Z(product[33]) );
  CENX1 U4780 ( .A(net16389), .B(net16676), .Z(n2371) );
  CND2XL U4781 ( .A(n757), .B(n3061), .Z(n175) );
  COND2X1 U4782 ( .A(n108), .B(n2406), .C(n3957), .D(n2405), .Z(n1884) );
  CIVX4 U4783 ( .A(n3921), .Z(n4024) );
  COND2XL U4784 ( .A(n3904), .B(n2618), .C(n3832), .D(n2617), .Z(n2091) );
  COND2XL U4785 ( .A(n2620), .B(n3904), .C(n3833), .D(n2619), .Z(n2093) );
  CENXL U4786 ( .A(n2808), .B(n4012), .Z(n2643) );
  CENXL U4787 ( .A(n3985), .B(n4012), .Z(n2638) );
  CENXL U4788 ( .A(net16391), .B(n4012), .Z(n2636) );
  CENXL U4789 ( .A(n3996), .B(n4012), .Z(n2615) );
  CENXL U4790 ( .A(n3996), .B(net16676), .Z(n2351) );
  CENXL U4791 ( .A(n3985), .B(net16676), .Z(n2374) );
  CENXL U4792 ( .A(n2808), .B(n3348), .Z(n2709) );
  CENXL U4793 ( .A(n3998), .B(n3348), .Z(n2712) );
  CENXL U4794 ( .A(net16399), .B(n3348), .Z(n2706) );
  CENXL U4795 ( .A(net16407), .B(n3348), .Z(n2710) );
  CENXL U4796 ( .A(n3984), .B(n3348), .Z(n2711) );
  CENXL U4797 ( .A(n2806), .B(n3348), .Z(n2707) );
  CENXL U4798 ( .A(n3985), .B(n3357), .Z(n2704) );
  CENXL U4799 ( .A(net16393), .B(n4006), .Z(n2703) );
  CENXL U4800 ( .A(net16389), .B(n4006), .Z(n2701) );
  CENXL U4801 ( .A(net16391), .B(n4007), .Z(n2702) );
  CNR2X1 U4802 ( .A(n1274), .B(n1245), .Z(n543) );
  CIVXL U4803 ( .A(n417), .Z(n419) );
  CENXL U4804 ( .A(n450), .B(n169), .Z(product[43]) );
  CENXL U4805 ( .A(n435), .B(n168), .Z(product[44]) );
  CENXL U4806 ( .A(n328), .B(n159), .Z(product[53]) );
  CENXL U4807 ( .A(n470), .B(n171), .Z(product[41]) );
  CENXL U4808 ( .A(n297), .B(n156), .Z(product[56]) );
  CIVX4 U4809 ( .A(net16580), .Z(net15999) );
  CENXL U4810 ( .A(n3991), .B(net19845), .Z(n2460) );
  CNIVX4 U4811 ( .A(n4007), .Z(n3956) );
  COND2X1 U4812 ( .A(n54), .B(n3907), .C(n3267), .D(n3901), .Z(n2069) );
  COND2X1 U4813 ( .A(n2715), .B(net16639), .C(n3743), .D(n2716), .Z(n2189) );
  CND2X4 U4814 ( .A(net16617), .B(n2812), .Z(net18570) );
  CENXL U4815 ( .A(net16403), .B(n3348), .Z(n2708) );
  CENXL U4816 ( .A(net16403), .B(n3930), .Z(n2675) );
  CENXL U4817 ( .A(net16403), .B(n4004), .Z(n2741) );
  CENXL U4818 ( .A(net16403), .B(n4012), .Z(n2642) );
  CENXL U4819 ( .A(net16403), .B(n4018), .Z(n2510) );
  CENXL U4820 ( .A(net16403), .B(n4023), .Z(n2279) );
  CENXL U4821 ( .A(n173), .B(n486), .Z(product[39]) );
  CENXL U4822 ( .A(n174), .B(n495), .Z(product[38]) );
  CENXL U4823 ( .A(n175), .B(n506), .Z(product[37]) );
  CENX2 U4824 ( .A(a[4]), .B(n3982), .Z(n24) );
  CIVXL U4825 ( .A(n517), .Z(net18568) );
  CIVXL U4826 ( .A(net18617), .Z(n756) );
  CAOR1XL U4827 ( .A(net16606), .B(n3172), .C(n2351), .Z(n1834) );
  COND2XL U4828 ( .A(n3173), .B(n2355), .C(net16606), .D(n2354), .Z(n1838) );
  COND2XL U4829 ( .A(n2352), .B(net16605), .C(n2353), .D(n3173), .Z(n1836) );
  CENXL U4830 ( .A(n411), .B(n166), .Z(product[46]) );
  CENXL U4831 ( .A(n393), .B(n164), .Z(product[48]) );
  CENXL U4832 ( .A(n371), .B(n162), .Z(product[50]) );
  CENXL U4833 ( .A(n352), .B(n161), .Z(product[51]) );
  CENXL U4834 ( .A(n317), .B(n158), .Z(product[54]) );
  CIVX2 U4835 ( .A(n1801), .Z(n3972) );
  CENX4 U4836 ( .A(n3073), .B(net18944), .Z(net16605) );
  CNR2X1 U4837 ( .A(n1581), .B(n1596), .Z(n643) );
  CENXL U4838 ( .A(n2804), .B(n3956), .Z(n2705) );
  CENXL U4839 ( .A(n2792), .B(n3956), .Z(n2693) );
  CANR1X2 U4840 ( .A(n3949), .B(n707), .C(n704), .Z(n702) );
  CND2X2 U4841 ( .A(n3926), .B(n709), .Z(n707) );
  CNIVX4 U4842 ( .A(net16593), .Z(net18545) );
  CENX2 U4843 ( .A(a[4]), .B(n3982), .Z(net16593) );
  CENX2 U4844 ( .A(n2783), .B(n3956), .Z(n2684) );
  CENXL U4845 ( .A(n2783), .B(net15975), .Z(n2354) );
  CENXL U4846 ( .A(n2781), .B(net15975), .Z(n2352) );
  CENXL U4847 ( .A(n2784), .B(net15975), .Z(n2355) );
  CENXL U4848 ( .A(n3995), .B(net15979), .Z(n2356) );
  CENXL U4849 ( .A(n3994), .B(net15979), .Z(n2357) );
  CENXL U4850 ( .A(n3993), .B(net15975), .Z(n2358) );
  CENXL U4851 ( .A(n2789), .B(net15975), .Z(n2360) );
  CENXL U4852 ( .A(n3992), .B(net15975), .Z(n2359) );
  CENXL U4853 ( .A(n3991), .B(net15975), .Z(n2361) );
  CENXL U4854 ( .A(n2804), .B(net15979), .Z(n2375) );
  CENXL U4855 ( .A(n2792), .B(net15979), .Z(n2363) );
  CENXL U4856 ( .A(n3989), .B(n4013), .Z(n2631) );
  CENXL U4857 ( .A(n2793), .B(n4013), .Z(n2628) );
  CND2IXL U4858 ( .B(n3998), .A(n4013), .Z(n2647) );
  CENXL U4859 ( .A(n3988), .B(n4013), .Z(n2632) );
  CENXL U4860 ( .A(n3987), .B(n4013), .Z(n2633) );
  CENXL U4861 ( .A(n2794), .B(n4013), .Z(n2629) );
  CENXL U4862 ( .A(n3990), .B(n4013), .Z(n2630) );
  CNR2X2 U4863 ( .A(n1613), .B(n1626), .Z(n660) );
  CENXL U4864 ( .A(n2806), .B(n4000), .Z(n2773) );
  CENXL U4865 ( .A(n3997), .B(n4000), .Z(n2778) );
  CENXL U4866 ( .A(n2804), .B(n4000), .Z(n2771) );
  CENXL U4867 ( .A(net16391), .B(n4000), .Z(n2768) );
  CENXL U4868 ( .A(net16399), .B(n4000), .Z(n2772) );
  CENXL U4869 ( .A(n3984), .B(n4000), .Z(n2777) );
  CENXL U4870 ( .A(net16389), .B(n4000), .Z(n2767) );
  CENXL U4871 ( .A(net16393), .B(n4000), .Z(n2769) );
  CENXL U4872 ( .A(n3985), .B(n4000), .Z(n2770) );
  CENXL U4873 ( .A(n3986), .B(n4000), .Z(n2766) );
  CENXL U4874 ( .A(net16407), .B(n4000), .Z(n2776) );
  CENXL U4875 ( .A(n2808), .B(n4000), .Z(n2775) );
  CENXL U4876 ( .A(net16403), .B(n4000), .Z(n2774) );
  CENXL U4877 ( .A(n3998), .B(net16023), .Z(n2580) );
  CENXL U4878 ( .A(n3995), .B(net16023), .Z(n2554) );
  CENXL U4879 ( .A(n2781), .B(net16023), .Z(n2550) );
  CENXL U4880 ( .A(n3994), .B(net16023), .Z(n2555) );
  CENXL U4881 ( .A(n3993), .B(net16023), .Z(n2556) );
  CENXL U4882 ( .A(n3984), .B(net16023), .Z(n2579) );
  CENXL U4883 ( .A(n2804), .B(net16023), .Z(n2573) );
  CENXL U4884 ( .A(n2791), .B(net16023), .Z(n2560) );
  CENXL U4885 ( .A(n2789), .B(net16023), .Z(n2558) );
  CIVXL U4886 ( .A(n3393), .Z(n649) );
  CENXL U4887 ( .A(n2781), .B(n4015), .Z(n2583) );
  CENXL U4888 ( .A(n2804), .B(n4015), .Z(n2606) );
  CENXL U4889 ( .A(n2783), .B(n4015), .Z(n2585) );
  CENXL U4890 ( .A(n2784), .B(n4015), .Z(n2586) );
  CENXL U4891 ( .A(n3995), .B(n3961), .Z(n2587) );
  CENXL U4892 ( .A(n2792), .B(n4015), .Z(n2594) );
  CENXL U4893 ( .A(n3993), .B(n3212), .Z(n2589) );
  CENXL U4894 ( .A(n2789), .B(n4015), .Z(n2591) );
  CENXL U4895 ( .A(n2791), .B(n4015), .Z(n2593) );
  CNIVX4 U4896 ( .A(net16015), .Z(net18510) );
  CANR1X2 U4897 ( .A(n3945), .B(n3950), .C(n712), .Z(n710) );
  CIVX4 U4898 ( .A(n75), .Z(n4019) );
  CIVXL U4899 ( .A(n463), .Z(n3919) );
  CIVXL U4900 ( .A(n461), .Z(n463) );
  COND1X1 U4901 ( .A(net19689), .B(n441), .C(n3206), .Z(n415) );
  CIVX4 U4902 ( .A(a[0]), .Z(n6) );
  CNIVX4 U4903 ( .A(n105), .Z(n3957) );
  CIVX1 U4904 ( .A(n4010), .Z(n3929) );
  CND2X1 U4905 ( .A(net18453), .B(net21614), .Z(n3923) );
  COND1X1 U4906 ( .A(n678), .B(n690), .C(n679), .Z(n677) );
  CENX1 U4907 ( .A(n205), .B(n707), .Z(product[7]) );
  CND2X1 U4908 ( .A(n3924), .B(n3925), .Z(n3926) );
  CIVX2 U4909 ( .A(n710), .Z(n3924) );
  COR2XL U4910 ( .A(n18), .B(n2742), .Z(n3927) );
  COR2XL U4911 ( .A(net16638), .B(n2741), .Z(n3928) );
  CND2X1 U4912 ( .A(n3927), .B(n3928), .Z(n2215) );
  CNR2XL U4913 ( .A(n3903), .B(n2643), .Z(n3931) );
  CNR2XL U4914 ( .A(n3959), .B(n2642), .Z(n3932) );
  COR2X1 U4915 ( .A(n3932), .B(n3931), .Z(n2116) );
  COR2X1 U4916 ( .A(n2250), .B(n2219), .Z(n3952) );
  CND2XL U4917 ( .A(n799), .B(n802), .Z(n255) );
  CNIVX2 U4918 ( .A(n145), .Z(n3998) );
  CENXL U4919 ( .A(n3997), .B(n3212), .Z(n2613) );
  CENXL U4920 ( .A(n3997), .B(n4012), .Z(n2646) );
  CND2X2 U4921 ( .A(n767), .B(n768), .Z(n578) );
  CND2X2 U4922 ( .A(n751), .B(n3419), .Z(n444) );
  CENXL U4923 ( .A(n208), .B(n721), .Z(product[4]) );
  COND2XL U4924 ( .A(n2580), .B(n3059), .C(n3355), .D(n2579), .Z(n2053) );
  COND2X1 U4925 ( .A(n3188), .B(n2499), .C(net21601), .D(n2498), .Z(n1973) );
  CNIVX1 U4926 ( .A(n145), .Z(n3997) );
  CND2XL U4927 ( .A(n355), .B(n331), .Z(n329) );
  CANR1X1 U4928 ( .A(n3944), .B(n659), .C(n654), .Z(n652) );
  CND2X1 U4929 ( .A(n879), .B(n892), .Z(n379) );
  CND2X1 U4930 ( .A(n3942), .B(n3946), .Z(n333) );
  CND2XL U4931 ( .A(n786), .B(n701), .Z(n204) );
  CND2X1 U4932 ( .A(n827), .B(n834), .Z(n316) );
  CENX1 U4933 ( .A(n3994), .B(n3933), .Z(n2687) );
  CIVX8 U4934 ( .A(n4019), .Z(n4017) );
  CND2XL U4935 ( .A(n516), .B(n758), .Z(n507) );
  CND2XL U4936 ( .A(n3419), .B(n3369), .Z(n170) );
  CND2XL U4937 ( .A(n392), .B(n746), .Z(n164) );
  CND2XL U4938 ( .A(n3943), .B(n434), .Z(n168) );
  CND2XL U4939 ( .A(n3942), .B(n351), .Z(n161) );
  CND2XL U4940 ( .A(n747), .B(n3558), .Z(n165) );
  CND2XL U4941 ( .A(n383), .B(n3550), .Z(n372) );
  CIVXL U4942 ( .A(n383), .Z(n381) );
  CEOXL U4943 ( .A(n190), .B(n624), .Z(product[22]) );
  CND2XL U4944 ( .A(n772), .B(n623), .Z(n190) );
  CND2XL U4945 ( .A(n779), .B(n3155), .Z(n197) );
  CND2XL U4946 ( .A(n3948), .B(n3947), .Z(n678) );
  CND2XL U4947 ( .A(n738), .B(n296), .Z(n156) );
  CND2XL U4948 ( .A(n355), .B(n320), .Z(n318) );
  CND2XL U4949 ( .A(n355), .B(n3942), .Z(n344) );
  CND2XL U4950 ( .A(n3946), .B(n342), .Z(n160) );
  CND2XL U4951 ( .A(n741), .B(n327), .Z(n159) );
  CND2XL U4952 ( .A(n355), .B(n283), .Z(n281) );
  CND2XL U4953 ( .A(net18264), .B(n279), .Z(n155) );
  CEOXL U4954 ( .A(n200), .B(n684), .Z(product[12]) );
  CND2XL U4955 ( .A(n3948), .B(n683), .Z(n200) );
  CND2XL U4956 ( .A(n781), .B(n675), .Z(n199) );
  CND2XL U4957 ( .A(n785), .B(n697), .Z(n203) );
  CEOXL U4958 ( .A(n702), .B(n204), .Z(product[8]) );
  CND2XL U4959 ( .A(n3947), .B(n688), .Z(n201) );
  CANR1X1 U4960 ( .A(n729), .B(n3952), .C(n726), .Z(n724) );
  CIVXL U4961 ( .A(n222), .Z(n220) );
  CIVXL U4962 ( .A(n259), .Z(n257) );
  CENXL U4963 ( .A(n247), .B(n152), .Z(product[60]) );
  CND2XL U4964 ( .A(net18255), .B(n246), .Z(n152) );
  CND2XL U4965 ( .A(n1701), .B(n1706), .Z(n701) );
  CND2XL U4966 ( .A(n1685), .B(n1692), .Z(n694) );
  CND2XL U4967 ( .A(n3949), .B(n706), .Z(n205) );
  CND2XL U4968 ( .A(n3952), .B(n728), .Z(n210) );
  CND2XL U4969 ( .A(n3951), .B(n720), .Z(n208) );
  CND2XL U4970 ( .A(n3950), .B(n714), .Z(n207) );
  CND2XL U4971 ( .A(n1713), .B(n1716), .Z(n709) );
  CND2XL U4972 ( .A(n1723), .B(n2218), .Z(n723) );
  COND2XL U4973 ( .A(n2646), .B(n3904), .C(n3832), .D(n2645), .Z(n2119) );
  CNR2IX1 U4974 ( .B(n3998), .A(net18545), .Z(n2186) );
  COND2XL U4975 ( .A(n3058), .B(n2578), .C(n3918), .D(n2577), .Z(n2051) );
  CNR2IXL U4976 ( .B(n3998), .A(n3918), .Z(n2054) );
  COND2XL U4977 ( .A(n3163), .B(n2656), .C(n3424), .D(n2655), .Z(n2129) );
  COND2XL U4978 ( .A(n3903), .B(n2644), .C(n2643), .D(n3833), .Z(n2117) );
  CENXL U4979 ( .A(n2782), .B(net15975), .Z(n2353) );
  CIVX8 U4980 ( .A(n3697), .Z(n4007) );
  CANR1XL U4981 ( .A(n699), .B(n691), .C(n3148), .Z(n3938) );
  CND2XL U4982 ( .A(net19757), .B(n760), .Z(n525) );
  CND2XL U4983 ( .A(n489), .B(n516), .Z(n487) );
  CANR1XL U4984 ( .A(n758), .B(n517), .C(n510), .Z(n508) );
  CANR1XL U4985 ( .A(n489), .B(n517), .C(n490), .Z(n488) );
  COND1XL U4986 ( .A(n501), .B(net18617), .C(net18783), .Z(n490) );
  CANR1XL U4987 ( .A(n3419), .B(n463), .C(n456), .Z(n452) );
  CND2XL U4988 ( .A(n751), .B(n449), .Z(n169) );
  COND1XL U4989 ( .A(n507), .B(net19290), .C(n508), .Z(n506) );
  COND1XL U4990 ( .A(net19290), .B(n496), .C(n497), .Z(n495) );
  COND1XL U4991 ( .A(n487), .B(n3069), .C(n488), .Z(n486) );
  CND2XL U4992 ( .A(n3341), .B(n541), .Z(n179) );
  COND1XL U4993 ( .A(n543), .B(net19290), .C(n3865), .Z(n542) );
  CND2XL U4994 ( .A(n760), .B(n530), .Z(n178) );
  COND1XL U4995 ( .A(n532), .B(net19290), .C(n3970), .Z(n531) );
  CND2XL U4996 ( .A(n758), .B(net19358), .Z(n176) );
  COND1XL U4997 ( .A(n514), .B(net19290), .C(net18568), .Z(n513) );
  CND2XL U4998 ( .A(n766), .B(n573), .Z(n184) );
  CND2XL U4999 ( .A(n583), .B(n767), .Z(n185) );
  CND2XL U5000 ( .A(n596), .B(n768), .Z(n585) );
  CANR1XL U5001 ( .A(n561), .B(n574), .C(n3162), .Z(n560) );
  CANR1XL U5002 ( .A(n620), .B(n629), .C(n3031), .Z(n619) );
  CND2XL U5003 ( .A(n753), .B(n469), .Z(n171) );
  CND2X1 U5004 ( .A(n387), .B(n418), .Z(n385) );
  CANR1XL U5005 ( .A(n768), .B(n597), .C(n590), .Z(n586) );
  CEOXL U5006 ( .A(n3062), .B(n188), .Z(product[24]) );
  CND2XL U5007 ( .A(n770), .B(net18869), .Z(n188) );
  COND1XL U5008 ( .A(n389), .B(n399), .C(n392), .Z(n388) );
  CANR1XL U5009 ( .A(n3943), .B(net21583), .C(n432), .Z(n428) );
  CND2XL U5010 ( .A(n749), .B(n3712), .Z(n167) );
  CND2XL U5011 ( .A(n438), .B(n3943), .Z(n427) );
  CND2XL U5012 ( .A(n748), .B(n410), .Z(n166) );
  COND1XL U5013 ( .A(n525), .B(n3069), .C(n526), .Z(n524) );
  COND1X1 U5014 ( .A(n551), .B(n559), .C(n552), .Z(n550) );
  CNR2X1 U5015 ( .A(n627), .B(n622), .Z(n620) );
  CNR2X1 U5016 ( .A(n665), .B(n660), .Z(n658) );
  CNR2X1 U5017 ( .A(n1037), .B(n1058), .Z(n471) );
  COR2X1 U5018 ( .A(n1460), .B(n1437), .Z(net18282) );
  CND2XL U5019 ( .A(n744), .B(n370), .Z(n162) );
  CND2XL U5020 ( .A(n3550), .B(n379), .Z(n163) );
  COR2X1 U5021 ( .A(n3554), .B(n1504), .Z(net18280) );
  CND2X1 U5022 ( .A(n1037), .B(n1058), .Z(n472) );
  CND2X1 U5023 ( .A(n3909), .B(n1304), .Z(n552) );
  CND2X1 U5024 ( .A(n995), .B(n1014), .Z(n458) );
  CND2X1 U5025 ( .A(n975), .B(n994), .Z(n449) );
  CND2X1 U5026 ( .A(n1437), .B(n1460), .Z(n603) );
  CND2X1 U5027 ( .A(n3554), .B(n1504), .Z(n618) );
  CND2X1 U5028 ( .A(n1333), .B(n1360), .Z(n568) );
  CND2XL U5029 ( .A(n773), .B(n628), .Z(n191) );
  CENX1 U5030 ( .A(n642), .B(n193), .Z(product[19]) );
  COND1XL U5031 ( .A(n3481), .B(n649), .C(n644), .Z(n642) );
  COND1XL U5032 ( .A(n636), .B(n649), .C(net19965), .Z(n635) );
  CANR1XL U5033 ( .A(n658), .B(n667), .C(n659), .Z(n657) );
  CEOXL U5034 ( .A(n194), .B(n649), .Z(product[18]) );
  CND2XL U5035 ( .A(n776), .B(n644), .Z(n194) );
  CENX1 U5036 ( .A(n1389), .B(n3939), .Z(n1387) );
  CENX1 U5037 ( .A(n1414), .B(n1391), .Z(n3939) );
  CENX1 U5038 ( .A(n3940), .B(n1439), .Z(n1437) );
  CENX1 U5039 ( .A(n1441), .B(n1462), .Z(n3940) );
  CND2XL U5040 ( .A(n739), .B(n303), .Z(n157) );
  CND2XL U5041 ( .A(n740), .B(n316), .Z(n158) );
  CNR2X1 U5042 ( .A(n1525), .B(n1544), .Z(n627) );
  COR2X1 U5043 ( .A(n1580), .B(n1563), .Z(net18274) );
  COR2X1 U5044 ( .A(n855), .B(n866), .Z(n3942) );
  COR2X1 U5045 ( .A(n974), .B(n957), .Z(n3943) );
  CNR2X1 U5046 ( .A(n879), .B(n892), .Z(n378) );
  COR2X1 U5047 ( .A(n1597), .B(n1612), .Z(n3944) );
  CND2X1 U5048 ( .A(n1525), .B(n1544), .Z(n628) );
  CND2X1 U5049 ( .A(n1627), .B(n1640), .Z(n666) );
  CND2X1 U5050 ( .A(n855), .B(n866), .Z(n351) );
  CND2X1 U5051 ( .A(n1597), .B(n1612), .Z(n656) );
  CND2X1 U5052 ( .A(n907), .B(n922), .Z(n403) );
  CND2X1 U5053 ( .A(n1505), .B(n1524), .Z(n623) );
  CNR2XL U5054 ( .A(n333), .B(n324), .Z(n320) );
  COND1XL U5055 ( .A(n324), .B(n334), .C(n327), .Z(n323) );
  CENX1 U5056 ( .A(n673), .B(n198), .Z(product[14]) );
  CENX1 U5057 ( .A(n689), .B(n201), .Z(product[11]) );
  CENX1 U5058 ( .A(n202), .B(n695), .Z(product[10]) );
  COND1XL U5059 ( .A(n696), .B(n698), .C(n697), .Z(n695) );
  CANR1XL U5060 ( .A(n3947), .B(n689), .C(n686), .Z(n684) );
  CEOXL U5061 ( .A(n199), .B(n676), .Z(product[13]) );
  CEOXL U5062 ( .A(n698), .B(n203), .Z(product[9]) );
  CND2XL U5063 ( .A(n320), .B(n740), .Z(n309) );
  COND1XL U5064 ( .A(n724), .B(n722), .C(n723), .Z(n721) );
  CNR2X1 U5065 ( .A(n1693), .B(n1700), .Z(n696) );
  CNR2X1 U5066 ( .A(n1685), .B(n1692), .Z(n693) );
  CND2X1 U5067 ( .A(n3953), .B(n218), .Z(n150) );
  CND2XL U5068 ( .A(n735), .B(n255), .Z(n153) );
  COND1XL U5069 ( .A(n248), .B(n3922), .C(n249), .Z(n247) );
  CND2XL U5070 ( .A(n259), .B(n735), .Z(n248) );
  CAOR1X1 U5071 ( .A(n721), .B(n3951), .C(n718), .Z(n3945) );
  CNR2X1 U5072 ( .A(n827), .B(n834), .Z(n315) );
  CNR2X1 U5073 ( .A(n1701), .B(n1706), .Z(n700) );
  COR2X1 U5074 ( .A(n845), .B(n854), .Z(n3946) );
  COR2X1 U5075 ( .A(n1675), .B(n1684), .Z(n3947) );
  COR2X1 U5076 ( .A(n1674), .B(n1665), .Z(n3948) );
  CND2X1 U5077 ( .A(n1653), .B(n1664), .Z(n675) );
  CND2X1 U5078 ( .A(n1693), .B(n1700), .Z(n697) );
  CND2X1 U5079 ( .A(n845), .B(n854), .Z(n342) );
  CND2X1 U5080 ( .A(n1675), .B(n1684), .Z(n688) );
  CND2X1 U5081 ( .A(n1665), .B(n1674), .Z(n683) );
  CND2XL U5082 ( .A(n222), .B(n3953), .Z(n213) );
  CANR1XL U5083 ( .A(n3953), .B(n3066), .C(n216), .Z(n214) );
  CENX1 U5084 ( .A(n207), .B(n3945), .Z(product[5]) );
  CEOXL U5085 ( .A(n724), .B(n209), .Z(product[3]) );
  CND2X1 U5086 ( .A(n791), .B(n723), .Z(n209) );
  CEOXL U5087 ( .A(n710), .B(n206), .Z(product[6]) );
  CND2X1 U5088 ( .A(n3925), .B(n709), .Z(n206) );
  COR2X1 U5089 ( .A(n807), .B(n812), .Z(net18264) );
  CND2X1 U5090 ( .A(n835), .B(n844), .Z(n327) );
  CND2X1 U5091 ( .A(n807), .B(n812), .Z(n279) );
  CND2X1 U5092 ( .A(n813), .B(n818), .Z(n296) );
  CENX1 U5093 ( .A(n210), .B(n729), .Z(product[2]) );
  CNR2X1 U5094 ( .A(n1723), .B(n2218), .Z(n722) );
  COR2X1 U5095 ( .A(n1707), .B(n1712), .Z(n3949) );
  COR2X1 U5096 ( .A(n1717), .B(n1720), .Z(n3950) );
  CENX1 U5097 ( .A(n1798), .B(n2034), .Z(n1273) );
  CND2X1 U5098 ( .A(n1721), .B(n1722), .Z(n720) );
  CND2X1 U5099 ( .A(n1717), .B(n1720), .Z(n714) );
  CND2X1 U5100 ( .A(n2250), .B(n2219), .Z(n728) );
  CND2X1 U5101 ( .A(n1707), .B(n1712), .Z(n706) );
  COR2X1 U5102 ( .A(n1721), .B(n1722), .Z(n3951) );
  CNR2X1 U5103 ( .A(n799), .B(n802), .Z(n254) );
  COR2X1 U5104 ( .A(n798), .B(n797), .Z(net18255) );
  COR2X1 U5105 ( .A(n1740), .B(n794), .Z(n3953) );
  CND2X1 U5106 ( .A(n798), .B(n797), .Z(n246) );
  CND2X1 U5107 ( .A(n1740), .B(n794), .Z(n218) );
  CAN2XL U5108 ( .A(n793), .B(n731), .Z(product[1]) );
  CENX1 U5109 ( .A(n2782), .B(net18486), .Z(n2419) );
  CENX1 U5110 ( .A(n2808), .B(net15963), .Z(n2313) );
  CENX1 U5111 ( .A(n2783), .B(n4009), .Z(n2651) );
  CENX1 U5112 ( .A(net16407), .B(net18407), .Z(n2314) );
  CENX1 U5113 ( .A(n3990), .B(net18485), .Z(n2432) );
  CENX1 U5114 ( .A(n2794), .B(net18486), .Z(n2431) );
  CENX1 U5115 ( .A(net16393), .B(net18407), .Z(n2307) );
  CENX1 U5116 ( .A(n3992), .B(net18485), .Z(n2425) );
  CENX1 U5117 ( .A(n2793), .B(net15993), .Z(n2430) );
  CENX1 U5118 ( .A(n3991), .B(net15993), .Z(n2427) );
  CENX1 U5119 ( .A(n2804), .B(net18486), .Z(n2441) );
  CENX1 U5120 ( .A(n2808), .B(net16649), .Z(n2445) );
  CENX1 U5121 ( .A(n3987), .B(net16027), .Z(n2567) );
  CENX1 U5122 ( .A(n2808), .B(n4009), .Z(n2676) );
  CENX1 U5123 ( .A(net16399), .B(n3929), .Z(n2673) );
  CENX1 U5124 ( .A(net16407), .B(n3929), .Z(n2677) );
  CENX1 U5125 ( .A(n2781), .B(n3999), .Z(n2748) );
  CENX1 U5126 ( .A(n2781), .B(n4009), .Z(n2649) );
  CENX1 U5127 ( .A(n3996), .B(n3929), .Z(n2648) );
  CENX1 U5128 ( .A(n3984), .B(net15963), .Z(n2315) );
  CNR2IXL U5129 ( .B(n3998), .A(net16639), .Z(n2219) );
  CENX1 U5130 ( .A(net16389), .B(net16649), .Z(n2437) );
  CENX1 U5131 ( .A(net16391), .B(net16649), .Z(n2438) );
  CENX1 U5132 ( .A(n3987), .B(net18520), .Z(n2402) );
  CENX1 U5133 ( .A(n3989), .B(net16645), .Z(n2532) );
  CENX1 U5134 ( .A(n3990), .B(net16671), .Z(n2465) );
  CENX1 U5135 ( .A(n3988), .B(net16645), .Z(n2533) );
  CENX1 U5136 ( .A(n2791), .B(net18520), .Z(n2395) );
  CENX1 U5137 ( .A(n3989), .B(net15963), .Z(n2301) );
  CENX1 U5138 ( .A(n3988), .B(net18520), .Z(n2401) );
  CENX1 U5139 ( .A(n3992), .B(net18520), .Z(n2392) );
  CENX1 U5140 ( .A(n2789), .B(net18520), .Z(n2393) );
  CENX1 U5141 ( .A(n3987), .B(net16645), .Z(n2534) );
  CENX1 U5142 ( .A(n2792), .B(net18520), .Z(n2396) );
  CENX1 U5143 ( .A(net16407), .B(net18486), .Z(n2446) );
  CENX1 U5144 ( .A(n3991), .B(n3956), .Z(n2691) );
  CENX1 U5145 ( .A(n3989), .B(n4024), .Z(n2268) );
  CENX1 U5146 ( .A(n3987), .B(n4024), .Z(n2270) );
  CENX1 U5147 ( .A(n3988), .B(n4024), .Z(n2269) );
  CENX1 U5148 ( .A(n3990), .B(n4024), .Z(n2267) );
  CENX1 U5149 ( .A(n2792), .B(n4024), .Z(n2264) );
  CNR2IX1 U5150 ( .B(n3998), .A(net19996), .Z(n1957) );
  CNR2IXL U5151 ( .B(n3998), .A(n3833), .Z(n2120) );
  CNR2IXL U5152 ( .B(n3998), .A(n3425), .Z(n2153) );
  CNR2IXL U5153 ( .B(n3998), .A(net16682), .Z(n2021) );
  CENX1 U5154 ( .A(n2782), .B(n3475), .Z(n2320) );
  CENX1 U5155 ( .A(n2782), .B(net18408), .Z(n2287) );
  CENX1 U5156 ( .A(n2783), .B(n3476), .Z(n2321) );
  CENX1 U5157 ( .A(n2789), .B(net18408), .Z(n2294) );
  CENX1 U5158 ( .A(n2784), .B(net18408), .Z(n2289) );
  CENX1 U5159 ( .A(n3993), .B(n3475), .Z(n2325) );
  CENX1 U5160 ( .A(n2783), .B(net15963), .Z(n2288) );
  CENX1 U5161 ( .A(n2792), .B(net15963), .Z(n2297) );
  CENX1 U5162 ( .A(n2783), .B(net18486), .Z(n2420) );
  CENX1 U5163 ( .A(n2782), .B(net18520), .Z(n2386) );
  CENX1 U5164 ( .A(n2782), .B(n3920), .Z(n2254) );
  CENX1 U5165 ( .A(n2783), .B(net18520), .Z(n2387) );
  CENX1 U5166 ( .A(n3994), .B(net18520), .Z(n2390) );
  CENX1 U5167 ( .A(n3993), .B(net18520), .Z(n2391) );
  CENX1 U5168 ( .A(n3995), .B(net18520), .Z(n2389) );
  CENX1 U5169 ( .A(n2784), .B(net18520), .Z(n2388) );
  CENX1 U5170 ( .A(n2794), .B(n4024), .Z(n2266) );
  CENX1 U5171 ( .A(n2791), .B(n4024), .Z(n2263) );
  CENX1 U5172 ( .A(n3991), .B(n4024), .Z(n2262) );
  CENX1 U5173 ( .A(n3993), .B(n4024), .Z(n2259) );
  CENX1 U5174 ( .A(n2789), .B(n4024), .Z(n2261) );
  CENX1 U5175 ( .A(n3992), .B(n4024), .Z(n2260) );
  CENX1 U5176 ( .A(n3994), .B(n4024), .Z(n2258) );
  CENX1 U5177 ( .A(n3995), .B(n3920), .Z(n2257) );
  CENX1 U5178 ( .A(n2784), .B(n3920), .Z(n2256) );
  CENX1 U5179 ( .A(n2783), .B(n3920), .Z(n2255) );
  CENX1 U5180 ( .A(n2781), .B(net18520), .Z(n2385) );
  CENX1 U5181 ( .A(n2781), .B(n3920), .Z(n2253) );
  CNR2IX1 U5182 ( .B(n3998), .A(n6), .Z(product[0]) );
  CNIVX8 U5183 ( .A(n2796), .Z(n3989) );
  CEOX2 U5184 ( .A(n3), .B(a[2]), .Z(net18096) );
  CENXL U5185 ( .A(n304), .B(n157), .Z(product[55]) );
  CENXL U5186 ( .A(n150), .B(n219), .Z(product[62]) );
  CND2IXL U5187 ( .B(n3998), .A(net18485), .Z(n2449) );
  COND2XL U5188 ( .A(n3904), .B(n3687), .C(n3959), .D(n2647), .Z(n1735) );
  CIVXL U5189 ( .A(n3175), .Z(net15993) );
  CENX1 U5190 ( .A(net16407), .B(net16671), .Z(n2479) );
  CENX1 U5191 ( .A(n3986), .B(net16671), .Z(n2469) );
  CENX4 U5192 ( .A(n3698), .B(n4007), .Z(n3960) );
  CENXL U5193 ( .A(n256), .B(n153), .Z(product[59]) );
  CENXL U5194 ( .A(n280), .B(n155), .Z(product[57]) );
  CND2IXL U5195 ( .B(n3998), .A(net16027), .Z(n2581) );
  CND2IXL U5196 ( .B(n3998), .A(n4020), .Z(n2350) );
  CIVX1 U5197 ( .A(n3133), .Z(n4009) );
  CENX1 U5198 ( .A(net16391), .B(n3929), .Z(n2669) );
  CND2IXL U5199 ( .B(n3998), .A(n3930), .Z(n2680) );
  CENX1 U5200 ( .A(n2791), .B(n3929), .Z(n2659) );
  CND2XL U5201 ( .A(n3053), .B(n1855), .Z(n3962) );
  CND2XL U5202 ( .A(n1855), .B(n1827), .Z(n3964) );
  CND3X1 U5203 ( .A(n3962), .B(n3963), .C(n3964), .Z(n1268) );
  CND2X1 U5204 ( .A(n1265), .B(n1269), .Z(n3966) );
  CNR2XL U5205 ( .A(n117), .B(n2375), .Z(n3968) );
  CNR2XL U5206 ( .A(net16605), .B(n2374), .Z(n3969) );
  COR2X1 U5207 ( .A(n3968), .B(n3969), .Z(n1855) );
  COND1XL U5208 ( .A(n3873), .B(n564), .C(n3801), .Z(n555) );
  COND2XL U5209 ( .A(n27), .B(n3857), .C(net18545), .D(n2713), .Z(n1737) );
  COAN1XL U5210 ( .A(n3865), .B(n3911), .C(n541), .Z(n3970) );
  CIVXL U5211 ( .A(n3970), .Z(n3971) );
  CANR1XL U5212 ( .A(n760), .B(n3971), .C(n528), .Z(n526) );
  CIVX1 U5213 ( .A(n3972), .Z(n3973) );
  CND2XL U5214 ( .A(n1439), .B(n1462), .Z(n3974) );
  CND2XL U5215 ( .A(n1462), .B(n1441), .Z(n3976) );
  CND3X1 U5216 ( .A(n3974), .B(n3975), .C(n3976), .Z(n1436) );
  CND2XL U5217 ( .A(n1389), .B(n1391), .Z(n3977) );
  CND2XL U5218 ( .A(n1389), .B(n1414), .Z(n3978) );
  CND3XL U5219 ( .A(n3977), .B(n3978), .C(n3979), .Z(n1386) );
  COND2XL U5220 ( .A(n3905), .B(n4002), .C(n6), .D(n2779), .Z(n1739) );
  CND2IXL U5221 ( .B(n3998), .A(n4001), .Z(n2779) );
  CND2X1 U5222 ( .A(n2251), .B(n1739), .Z(n731) );
  CNR2XL U5223 ( .A(n2251), .B(n1739), .Z(n730) );
  COR2XL U5224 ( .A(n1186), .B(net18607), .Z(n3980) );
  CIVX1 U5225 ( .A(n3734), .Z(n767) );
  CNR2X2 U5226 ( .A(n1186), .B(net18607), .Z(n522) );
  COND2XL U5227 ( .A(n63), .B(net16539), .C(n3355), .D(n2581), .Z(n1733) );
  COND2XL U5228 ( .A(n3352), .B(n3735), .C(n51), .D(n2614), .Z(n1734) );
  COND2XL U5229 ( .A(n18), .B(n3635), .C(n2746), .D(net16639), .Z(n1738) );
  COND2XL U5230 ( .A(net22025), .B(net19319), .C(net19996), .D(n2482), .Z(
        n1730) );
  COND2XL U5231 ( .A(n3163), .B(n3133), .C(n3424), .D(n2680), .Z(n1736) );
  COND1XL U5232 ( .A(n594), .B(n3062), .C(net18827), .Z(n593) );
  CIVXL U5233 ( .A(net18745), .Z(n757) );
  CND2X4 U5234 ( .A(n2825), .B(n24), .Z(n27) );
  CND2X4 U5235 ( .A(n3918), .B(n3090), .Z(n63) );
  CND2X4 U5236 ( .A(n2816), .B(n3958), .Z(n108) );
  CIVX2 U5237 ( .A(n842), .Z(n843) );
  CIVX2 U5238 ( .A(n824), .Z(n825) );
  CIVX2 U5239 ( .A(n810), .Z(n811) );
  CIVX2 U5240 ( .A(n800), .Z(n801) );
  CIVX2 U5241 ( .A(n730), .Z(n793) );
  CIVX2 U5242 ( .A(n722), .Z(n791) );
  CIVX2 U5243 ( .A(n700), .Z(n786) );
  CIVX2 U5244 ( .A(n696), .Z(n785) );
  CIVX2 U5245 ( .A(n622), .Z(n772) );
  CIVX2 U5246 ( .A(n324), .Z(n741) );
  CIVX2 U5247 ( .A(n295), .Z(n738) );
  CIVX2 U5248 ( .A(n731), .Z(n729) );
  CIVX2 U5249 ( .A(n728), .Z(n726) );
  CIVX2 U5250 ( .A(n720), .Z(n718) );
  CIVX2 U5251 ( .A(n714), .Z(n712) );
  CIVX2 U5252 ( .A(n706), .Z(n704) );
  CIVX2 U5253 ( .A(n699), .Z(n698) );
  CIVX2 U5254 ( .A(n3938), .Z(n689) );
  CIVX2 U5255 ( .A(n688), .Z(n686) );
  CIVX2 U5256 ( .A(n656), .Z(n654) );
  CIVX2 U5257 ( .A(n643), .Z(n776) );
  CIVX2 U5258 ( .A(n471), .Z(n754) );
  CIVX2 U5259 ( .A(n434), .Z(n432) );
  CIVX2 U5260 ( .A(n414), .Z(n412) );
  CIVX2 U5261 ( .A(n342), .Z(n340) );
  CIVX2 U5262 ( .A(n334), .Z(n332) );
  CIVX2 U5263 ( .A(n333), .Z(n331) );
  CIVX2 U5264 ( .A(n316), .Z(n314) );
  CIVX2 U5265 ( .A(n315), .Z(n740) );
  CIVX2 U5266 ( .A(n303), .Z(n301) );
  CIVX2 U5267 ( .A(n302), .Z(n739) );
  CIVX2 U5268 ( .A(n289), .Z(n287) );
  CIVX2 U5269 ( .A(n254), .Z(n735) );
  CIVX2 U5270 ( .A(n218), .Z(n216) );
endmodule


module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push0, en0_p0, en1_p0, push0_p0, push0_p2, push0_p1, en0_p1, en1_p1,
         en2_p1, en2_p2, en0_p2_d1, en1_p2_d1, en1_p2, en0_p2, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N398, N399, N400, N401, N402, N403, N404, N405, roundit,
         _pushout_d, N418, N419, N420, N421, N422, N423, N424, N425, N426,
         N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437,
         N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, n12,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276;
  wire   [1:0] cmd0;
  wire   [1:0] cmd0_p0;
  wire   [1:0] cmd0_p2;
  wire   [1:0] cmd0_p1;
  wire   [63:0] out0_p0;
  wire   [63:0] out0_p2;
  wire   [63:0] out0_p1;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] acc_cmd1;
  wire   [63:0] acc;
  wire   [63:0] out1_p2;
  wire   [63:0] out1_p0;
  wire   [63:0] out1_p1;
  wire   [63:0] acc_cmd2;
  wire   [63:0] out2_p2;
  wire   [6:0] h0_p1;
  wire   [6:0] h0_p0;

  CAOR2X1 U369 ( .A(h0_p0[0]), .B(en2_p1), .C(n1323), .D(n1949), .Z(n612) );
  CAOR2X1 U372 ( .A(h0_p0[1]), .B(en2_p1), .C(n1330), .D(n1949), .Z(n615) );
  CAOR2X1 U375 ( .A(h0_p0[2]), .B(en2_p1), .C(n1239), .D(n1949), .Z(n618) );
  CAOR2X1 U378 ( .A(h0_p0[3]), .B(en2_p1), .C(n1336), .D(n1949), .Z(n621) );
  CAOR2X1 U381 ( .A(h0_p0[4]), .B(en2_p1), .C(n1244), .D(n1949), .Z(n624) );
  CAOR2X1 U384 ( .A(h0_p0[5]), .B(en2_p1), .C(n1250), .D(n1949), .Z(n627) );
  CAOR2X1 U387 ( .A(h0_p0[6]), .B(en2_p1), .C(n1251), .D(n1949), .Z(n630) );
  CFD2QX2 \q0_reg[30]  ( .D(n688), .CP(clk), .CD(n1271), .Q(q0[30]) );
  CFD2QX2 \q0_reg[25]  ( .D(n683), .CP(clk), .CD(n1283), .Q(q0[25]) );
  CFD2QX2 \q0_reg[20]  ( .D(n1116), .CP(clk), .CD(n1283), .Q(q0[20]) );
  CFD2QX2 \q0_reg[4]  ( .D(n1113), .CP(clk), .CD(n1285), .Q(q0[4]) );
  CFD2QX2 \q0_reg[2]  ( .D(n1112), .CP(clk), .CD(n1285), .Q(q0[2]) );
  CFD2QX2 \q0_reg[0]  ( .D(n1111), .CP(clk), .CD(n1285), .Q(q0[0]) );
  sfilt_DW01_add_2 add_148 ( .A(out1_p1), .B(acc_cmd1), .CI(1'b0), .SUM({N271, 
        N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, 
        N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, 
        N210, N209, N208}) );
  sfilt_DW01_add_3 add_251 ( .A(out2_p2), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, roundit}), 
        .CI(1'b0), .SUM({N481, N480, N479, N478, N477, N476, N475, N474, N473, 
        N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, 
        N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, 
        N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, 
        N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, 
        N424, N423, N422, N421, N420, N419, N418}) );
  sfilt_DW_mult_tc_1 r304 ( .a({q0[31:15], n1236, q0[13:0]}), .b(h0), 
        .product({N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, 
        N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, 
        N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, 
        N23, N22, N21, N20, N19, N18, N17, N16, N15, N14}) );
  CFD2QX1 \q0_reg[27]  ( .D(n685), .CP(clk), .CD(n1271), .Q(q0[27]) );
  CFD2QX1 \q0_reg[15]  ( .D(n673), .CP(clk), .CD(n1284), .Q(q0[15]) );
  CFD2QX1 \q0_reg[13]  ( .D(n671), .CP(clk), .CD(n1284), .Q(q0[13]) );
  CFD2QX1 \q0_reg[3]  ( .D(n661), .CP(clk), .CD(n1285), .Q(q0[3]) );
  CFD2QX1 \q0_reg[19]  ( .D(n677), .CP(clk), .CD(n1284), .Q(q0[19]) );
  CFD2QX1 \q0_reg[7]  ( .D(n665), .CP(clk), .CD(n1284), .Q(q0[7]) );
  CFD2QX1 \q0_reg[29]  ( .D(n687), .CP(clk), .CD(n1271), .Q(q0[29]) );
  CFD2QXL \out0_p0_reg[42]  ( .D(N56), .CP(clk), .CD(n1308), .Q(out0_p0[42])
         );
  CFD2QXL \out1_p0_reg[42]  ( .D(N56), .CP(clk), .CD(n1272), .Q(out1_p0[42])
         );
  CFD2QXL \out0_p0_reg[43]  ( .D(N57), .CP(clk), .CD(n1308), .Q(out0_p0[43])
         );
  CFD2QXL \out1_p0_reg[43]  ( .D(N57), .CP(clk), .CD(n1272), .Q(out1_p0[43])
         );
  CFD2QXL \out0_p0_reg[44]  ( .D(N58), .CP(clk), .CD(n1307), .Q(out0_p0[44])
         );
  CFD2QXL \out1_p0_reg[44]  ( .D(N58), .CP(clk), .CD(n1272), .Q(out1_p0[44])
         );
  CFD2QXL \out0_p0_reg[45]  ( .D(N59), .CP(clk), .CD(n1307), .Q(out0_p0[45])
         );
  CFD2QXL \out1_p0_reg[45]  ( .D(N59), .CP(clk), .CD(n1272), .Q(out1_p0[45])
         );
  CFD2QXL \out0_p0_reg[46]  ( .D(N60), .CP(clk), .CD(n1307), .Q(out0_p0[46])
         );
  CFD2QXL \out1_p0_reg[46]  ( .D(N60), .CP(clk), .CD(n1271), .Q(out1_p0[46])
         );
  CFD2QXL \out0_p0_reg[47]  ( .D(N61), .CP(clk), .CD(n1306), .Q(out0_p0[47])
         );
  CFD2QXL \out1_p0_reg[47]  ( .D(N61), .CP(clk), .CD(n1271), .Q(out1_p0[47])
         );
  CFD2QXL \out0_p0_reg[48]  ( .D(N62), .CP(clk), .CD(n1306), .Q(out0_p0[48])
         );
  CFD2QXL \out1_p0_reg[48]  ( .D(N62), .CP(clk), .CD(n1271), .Q(out1_p0[48])
         );
  CFD2QXL \out0_p0_reg[49]  ( .D(N63), .CP(clk), .CD(n1305), .Q(out0_p0[49])
         );
  CFD2QXL \out1_p0_reg[49]  ( .D(N63), .CP(clk), .CD(n1292), .Q(out1_p0[49])
         );
  CFD2QXL \out0_p0_reg[50]  ( .D(N64), .CP(clk), .CD(n1305), .Q(out0_p0[50])
         );
  CFD2QXL \out1_p0_reg[50]  ( .D(N64), .CP(clk), .CD(n1292), .Q(out1_p0[50])
         );
  CFD2QXL \out0_p0_reg[51]  ( .D(N65), .CP(clk), .CD(n1311), .Q(out0_p0[51])
         );
  CFD2QXL \out1_p0_reg[51]  ( .D(N65), .CP(clk), .CD(n1292), .Q(out1_p0[51])
         );
  CFD2QXL \out0_p0_reg[52]  ( .D(N66), .CP(clk), .CD(n1283), .Q(out0_p0[52])
         );
  CFD2QXL \out1_p0_reg[52]  ( .D(N66), .CP(clk), .CD(n1292), .Q(out1_p0[52])
         );
  CFD2QXL \out0_p0_reg[53]  ( .D(N67), .CP(clk), .CD(n1282), .Q(out0_p0[53])
         );
  CFD2QXL \out1_p0_reg[53]  ( .D(N67), .CP(clk), .CD(n1292), .Q(out1_p0[53])
         );
  CFD2QXL \out0_p0_reg[54]  ( .D(N68), .CP(clk), .CD(n1282), .Q(out0_p0[54])
         );
  CFD2QXL \out1_p0_reg[54]  ( .D(N68), .CP(clk), .CD(n1291), .Q(out1_p0[54])
         );
  CFD2QXL \out0_p0_reg[55]  ( .D(N69), .CP(clk), .CD(n1282), .Q(out0_p0[55])
         );
  CFD2QXL \out1_p0_reg[55]  ( .D(N69), .CP(clk), .CD(n1291), .Q(out1_p0[55])
         );
  CFD2QXL \out0_p0_reg[56]  ( .D(N70), .CP(clk), .CD(n1281), .Q(out0_p0[56])
         );
  CFD2QXL \out1_p0_reg[56]  ( .D(N70), .CP(clk), .CD(n1291), .Q(out1_p0[56])
         );
  CFD2QXL \out0_p0_reg[57]  ( .D(N71), .CP(clk), .CD(n1281), .Q(out0_p0[57])
         );
  CFD2QXL \out1_p0_reg[57]  ( .D(N71), .CP(clk), .CD(n1291), .Q(out1_p0[57])
         );
  CFD2QXL \out0_p0_reg[58]  ( .D(N72), .CP(clk), .CD(n1280), .Q(out0_p0[58])
         );
  CFD2QXL \out1_p0_reg[58]  ( .D(N72), .CP(clk), .CD(n1291), .Q(out1_p0[58])
         );
  CFD2QXL \out0_p0_reg[59]  ( .D(N73), .CP(clk), .CD(n1280), .Q(out0_p0[59])
         );
  CFD2QXL \out1_p0_reg[59]  ( .D(N73), .CP(clk), .CD(n1291), .Q(out1_p0[59])
         );
  CFD2QXL \out0_p0_reg[60]  ( .D(N74), .CP(clk), .CD(n1280), .Q(out0_p0[60])
         );
  CFD2QXL \out1_p0_reg[60]  ( .D(N74), .CP(clk), .CD(n1290), .Q(out1_p0[60])
         );
  CFD2QXL \out0_p0_reg[61]  ( .D(N75), .CP(clk), .CD(n1279), .Q(out0_p0[61])
         );
  CFD2QXL \out1_p0_reg[61]  ( .D(N75), .CP(clk), .CD(n1290), .Q(out1_p0[61])
         );
  CFD2QXL \out0_p0_reg[62]  ( .D(N76), .CP(clk), .CD(n1279), .Q(out0_p0[62])
         );
  CFD2QXL \out1_p0_reg[62]  ( .D(N76), .CP(clk), .CD(n1290), .Q(out1_p0[62])
         );
  CFD2QX1 \q0_reg[14]  ( .D(n672), .CP(clk), .CD(n1284), .Q(q0[14]) );
  CFD2QXL \out1_p0_reg[41]  ( .D(N55), .CP(clk), .CD(n1272), .Q(out1_p0[41])
         );
  CFD2QXL \out1_p1_reg[41]  ( .D(n1075), .CP(clk), .CD(n1272), .Q(out1_p1[41])
         );
  CFD2QXL \out0_p1_reg[63]  ( .D(n1060), .CP(clk), .CD(n1288), .Q(out0_p1[63])
         );
  CFD2QXL \out0_p1_reg[62]  ( .D(n1058), .CP(clk), .CD(n1279), .Q(out0_p1[62])
         );
  CFD2QXL \out0_p1_reg[61]  ( .D(n1056), .CP(clk), .CD(n1279), .Q(out0_p1[61])
         );
  CFD2QXL \out0_p1_reg[60]  ( .D(n1054), .CP(clk), .CD(n1280), .Q(out0_p1[60])
         );
  CFD2QXL \out0_p1_reg[59]  ( .D(n1052), .CP(clk), .CD(n1280), .Q(out0_p1[59])
         );
  CFD2QXL \out0_p1_reg[58]  ( .D(n1050), .CP(clk), .CD(n1281), .Q(out0_p1[58])
         );
  CFD2QXL \out0_p1_reg[57]  ( .D(n1048), .CP(clk), .CD(n1281), .Q(out0_p1[57])
         );
  CFD2QXL \out0_p1_reg[56]  ( .D(n1046), .CP(clk), .CD(n1281), .Q(out0_p1[56])
         );
  CFD2QXL \out0_p1_reg[55]  ( .D(n1044), .CP(clk), .CD(n1282), .Q(out0_p1[55])
         );
  CFD2QXL \out0_p1_reg[54]  ( .D(n1042), .CP(clk), .CD(n1282), .Q(out0_p1[54])
         );
  CFD2QXL \out0_p1_reg[53]  ( .D(n1040), .CP(clk), .CD(n1282), .Q(out0_p1[53])
         );
  CFD2QXL \out0_p1_reg[52]  ( .D(n1038), .CP(clk), .CD(n1283), .Q(out0_p1[52])
         );
  CFD2QXL \out0_p1_reg[51]  ( .D(n1036), .CP(clk), .CD(n1305), .Q(out0_p1[51])
         );
  CFD2QXL \out0_p1_reg[50]  ( .D(n1034), .CP(clk), .CD(n1305), .Q(out0_p1[50])
         );
  CFD2QXL \out0_p1_reg[49]  ( .D(n1032), .CP(clk), .CD(n1305), .Q(out0_p1[49])
         );
  CFD2QXL \out0_p1_reg[48]  ( .D(n1030), .CP(clk), .CD(n1306), .Q(out0_p1[48])
         );
  CFD2QXL \out0_p1_reg[47]  ( .D(n1028), .CP(clk), .CD(n1306), .Q(out0_p1[47])
         );
  CFD2QXL \out0_p1_reg[46]  ( .D(n1026), .CP(clk), .CD(n1307), .Q(out0_p1[46])
         );
  CFD2QXL \out0_p1_reg[45]  ( .D(n1024), .CP(clk), .CD(n1307), .Q(out0_p1[45])
         );
  CFD2QXL \out0_p1_reg[44]  ( .D(n1022), .CP(clk), .CD(n1307), .Q(out0_p1[44])
         );
  CFD2QXL \out0_p1_reg[43]  ( .D(n1020), .CP(clk), .CD(n1308), .Q(out0_p1[43])
         );
  CFD2QXL \out0_p1_reg[42]  ( .D(n1018), .CP(clk), .CD(n1308), .Q(out0_p1[42])
         );
  CFD2QXL \out0_p1_reg[41]  ( .D(n1016), .CP(clk), .CD(n1309), .Q(out0_p1[41])
         );
  CFD2QXL \out0_p1_reg[40]  ( .D(n1014), .CP(clk), .CD(n1309), .Q(out0_p1[40])
         );
  CFD2QXL \out0_p1_reg[39]  ( .D(n1012), .CP(clk), .CD(n1309), .Q(out0_p1[39])
         );
  CFD2QXL \out0_p1_reg[38]  ( .D(n1010), .CP(clk), .CD(n1310), .Q(out0_p1[38])
         );
  CFD2QXL \out0_p1_reg[37]  ( .D(n1008), .CP(clk), .CD(n1310), .Q(out0_p1[37])
         );
  CFD2QXL \out0_p1_reg[36]  ( .D(n1006), .CP(clk), .CD(n1310), .Q(out0_p1[36])
         );
  CFD2QXL \out0_p1_reg[35]  ( .D(n1004), .CP(clk), .CD(n1311), .Q(out0_p1[35])
         );
  CFD2QXL \out0_p1_reg[34]  ( .D(n1002), .CP(clk), .CD(n1311), .Q(out0_p1[34])
         );
  CFD2QXL \out0_p1_reg[33]  ( .D(n1000), .CP(clk), .CD(n1312), .Q(out0_p1[33])
         );
  CFD2QXL \out0_p1_reg[32]  ( .D(n998), .CP(clk), .CD(n1312), .Q(out0_p1[32])
         );
  CFD2QXL \out0_p1_reg[31]  ( .D(n996), .CP(clk), .CD(n1313), .Q(out0_p1[31])
         );
  CFD2QXL \out0_p1_reg[30]  ( .D(n994), .CP(clk), .CD(n1313), .Q(out0_p1[30])
         );
  CFD2QXL \out0_p1_reg[29]  ( .D(n992), .CP(clk), .CD(n1312), .Q(out0_p1[29])
         );
  CFD2QXL \out0_p1_reg[28]  ( .D(n990), .CP(clk), .CD(n1314), .Q(out0_p1[28])
         );
  CFD2QXL \out0_p1_reg[27]  ( .D(n988), .CP(clk), .CD(n1314), .Q(out0_p1[27])
         );
  CFD2QXL \out0_p1_reg[26]  ( .D(n986), .CP(clk), .CD(n1314), .Q(out0_p1[26])
         );
  CFD2QXL \out0_p1_reg[25]  ( .D(n984), .CP(clk), .CD(n1315), .Q(out0_p1[25])
         );
  CFD2QXL \out0_p1_reg[24]  ( .D(n982), .CP(clk), .CD(n1315), .Q(out0_p1[24])
         );
  CFD2QXL \out0_p1_reg[23]  ( .D(n980), .CP(clk), .CD(n1316), .Q(out0_p1[23])
         );
  CFD2QXL \out0_p1_reg[22]  ( .D(n978), .CP(clk), .CD(n1316), .Q(out0_p1[22])
         );
  CFD2QXL \out0_p1_reg[21]  ( .D(n976), .CP(clk), .CD(n1316), .Q(out0_p1[21])
         );
  CFD2QXL \out0_p1_reg[20]  ( .D(n974), .CP(clk), .CD(n1317), .Q(out0_p1[20])
         );
  CFD2QXL \out0_p1_reg[19]  ( .D(n972), .CP(clk), .CD(n1292), .Q(out0_p1[19])
         );
  CFD2QXL \out0_p1_reg[18]  ( .D(n970), .CP(clk), .CD(n1293), .Q(out0_p1[18])
         );
  CFD2QXL \out0_p1_reg[17]  ( .D(n968), .CP(clk), .CD(n1293), .Q(out0_p1[17])
         );
  CFD2QXL \out0_p1_reg[16]  ( .D(n966), .CP(clk), .CD(n1293), .Q(out0_p1[16])
         );
  CFD2QXL \out0_p1_reg[15]  ( .D(n964), .CP(clk), .CD(n1294), .Q(out0_p1[15])
         );
  CFD2QXL \out0_p1_reg[14]  ( .D(n962), .CP(clk), .CD(n1294), .Q(out0_p1[14])
         );
  CFD2QXL \out0_p1_reg[13]  ( .D(n960), .CP(clk), .CD(n1295), .Q(out0_p1[13])
         );
  CFD2QXL \out0_p1_reg[12]  ( .D(n958), .CP(clk), .CD(n1295), .Q(out0_p1[12])
         );
  CFD2QXL \out0_p1_reg[11]  ( .D(n956), .CP(clk), .CD(n1295), .Q(out0_p1[11])
         );
  CFD2QXL \out0_p1_reg[10]  ( .D(n954), .CP(clk), .CD(n1296), .Q(out0_p1[10])
         );
  CFD2QXL \out0_p1_reg[9]  ( .D(n952), .CP(clk), .CD(n1296), .Q(out0_p1[9]) );
  CFD2QXL \out0_p1_reg[8]  ( .D(n950), .CP(clk), .CD(n1297), .Q(out0_p1[8]) );
  CFD2QXL \out0_p1_reg[7]  ( .D(n948), .CP(clk), .CD(n1297), .Q(out0_p1[7]) );
  CFD2QXL \out0_p1_reg[6]  ( .D(n946), .CP(clk), .CD(n1297), .Q(out0_p1[6]) );
  CFD2QXL \out0_p1_reg[5]  ( .D(n944), .CP(clk), .CD(n1298), .Q(out0_p1[5]) );
  CFD2QXL \out0_p1_reg[4]  ( .D(n942), .CP(clk), .CD(n1298), .Q(out0_p1[4]) );
  CFD2QXL \out0_p1_reg[3]  ( .D(n940), .CP(clk), .CD(n1305), .Q(out0_p1[3]) );
  CFD2QXL \out0_p1_reg[2]  ( .D(n938), .CP(clk), .CD(n1299), .Q(out0_p1[2]) );
  CFD2QXL \out0_p1_reg[1]  ( .D(n936), .CP(clk), .CD(n1299), .Q(out0_p1[1]) );
  CFD2QXL \out0_p1_reg[0]  ( .D(n934), .CP(clk), .CD(n1300), .Q(out0_p1[0]) );
  CFD2QXL \dout_reg[31]  ( .D(n786), .CP(clk), .CD(n1305), .Q(z[31]) );
  CFD2QXL \dout_reg[30]  ( .D(n785), .CP(clk), .CD(n1304), .Q(z[30]) );
  CFD2QXL \dout_reg[29]  ( .D(n784), .CP(clk), .CD(n1304), .Q(z[29]) );
  CFD2QXL \dout_reg[28]  ( .D(n783), .CP(clk), .CD(n1304), .Q(z[28]) );
  CFD2QXL \dout_reg[27]  ( .D(n782), .CP(clk), .CD(n1304), .Q(z[27]) );
  CFD2QXL \dout_reg[26]  ( .D(n781), .CP(clk), .CD(n1304), .Q(z[26]) );
  CFD2QXL \dout_reg[25]  ( .D(n780), .CP(clk), .CD(n1304), .Q(z[25]) );
  CFD2QXL \dout_reg[24]  ( .D(n779), .CP(clk), .CD(n1304), .Q(z[24]) );
  CFD2QXL \dout_reg[23]  ( .D(n778), .CP(clk), .CD(n1304), .Q(z[23]) );
  CFD2QXL \dout_reg[22]  ( .D(n777), .CP(clk), .CD(n1304), .Q(z[22]) );
  CFD2QXL \dout_reg[21]  ( .D(n776), .CP(clk), .CD(n1304), .Q(z[21]) );
  CFD2QXL \dout_reg[20]  ( .D(n775), .CP(clk), .CD(n1304), .Q(z[20]) );
  CFD2QXL \dout_reg[19]  ( .D(n774), .CP(clk), .CD(n1304), .Q(z[19]) );
  CFD2QXL \dout_reg[18]  ( .D(n773), .CP(clk), .CD(n1304), .Q(z[18]) );
  CFD2QXL \dout_reg[17]  ( .D(n772), .CP(clk), .CD(n1303), .Q(z[17]) );
  CFD2QXL \dout_reg[16]  ( .D(n771), .CP(clk), .CD(n1303), .Q(z[16]) );
  CFD2QXL \dout_reg[15]  ( .D(n770), .CP(clk), .CD(n1303), .Q(z[15]) );
  CFD2QXL \dout_reg[14]  ( .D(n769), .CP(clk), .CD(n1303), .Q(z[14]) );
  CFD2QXL \dout_reg[13]  ( .D(n768), .CP(clk), .CD(n1303), .Q(z[13]) );
  CFD2QXL \dout_reg[12]  ( .D(n767), .CP(clk), .CD(n1303), .Q(z[12]) );
  CFD2QXL \dout_reg[11]  ( .D(n766), .CP(clk), .CD(n1303), .Q(z[11]) );
  CFD2QXL \dout_reg[10]  ( .D(n765), .CP(clk), .CD(n1303), .Q(z[10]) );
  CFD2QXL \dout_reg[9]  ( .D(n764), .CP(clk), .CD(n1303), .Q(z[9]) );
  CFD2QXL \dout_reg[8]  ( .D(n763), .CP(clk), .CD(n1303), .Q(z[8]) );
  CFD2QXL \dout_reg[7]  ( .D(n762), .CP(clk), .CD(n1303), .Q(z[7]) );
  CFD2QXL \dout_reg[6]  ( .D(n761), .CP(clk), .CD(n1303), .Q(z[6]) );
  CFD2QXL \dout_reg[5]  ( .D(n760), .CP(clk), .CD(n1303), .Q(z[5]) );
  CFD2QXL \dout_reg[4]  ( .D(n759), .CP(clk), .CD(n1302), .Q(z[4]) );
  CFD2QXL \dout_reg[3]  ( .D(n758), .CP(clk), .CD(n1302), .Q(z[3]) );
  CFD2QXL \dout_reg[2]  ( .D(n757), .CP(clk), .CD(n1302), .Q(z[2]) );
  CFD2QXL \dout_reg[1]  ( .D(n756), .CP(clk), .CD(n1302), .Q(z[1]) );
  CFD2QXL \dout_reg[0]  ( .D(n755), .CP(clk), .CD(n1302), .Q(z[0]) );
  CFD2QXL \h0_p0_reg[6]  ( .D(n932), .CP(clk), .CD(n1302), .Q(h0_p0[6]) );
  CFD2QXL \h0_p0_reg[5]  ( .D(n930), .CP(clk), .CD(n1302), .Q(h0_p0[5]) );
  CFD2QXL \h0_p0_reg[4]  ( .D(n929), .CP(clk), .CD(n1302), .Q(h0_p0[4]) );
  CFD2QXL \h0_p0_reg[3]  ( .D(n928), .CP(clk), .CD(n1302), .Q(h0_p0[3]) );
  CFD2QXL \h0_p0_reg[2]  ( .D(n926), .CP(clk), .CD(n1302), .Q(h0_p0[2]) );
  CFD2QXL \h0_p0_reg[1]  ( .D(n924), .CP(clk), .CD(n1302), .Q(h0_p0[1]) );
  CFD2QXL \h0_p0_reg[0]  ( .D(n923), .CP(clk), .CD(n1302), .Q(h0_p0[0]) );
  CFD2QXL \h0_p1_reg[6]  ( .D(n630), .CP(clk), .CD(n1301), .Q(h0_p1[6]) );
  CFD2QXL \h0_p1_reg[5]  ( .D(n627), .CP(clk), .CD(n1300), .Q(h0_p1[5]) );
  CFD2QXL \out1_p1_reg[63]  ( .D(n921), .CP(clk), .CD(n1290), .Q(out1_p1[63])
         );
  CFD2QXL \out1_p1_reg[62]  ( .D(n919), .CP(clk), .CD(n1290), .Q(out1_p1[62])
         );
  CFD2QXL \out1_p1_reg[61]  ( .D(n917), .CP(clk), .CD(n1290), .Q(out1_p1[61])
         );
  CFD2QXL \out1_p1_reg[60]  ( .D(n915), .CP(clk), .CD(n1291), .Q(out1_p1[60])
         );
  CFD2QXL \out1_p1_reg[54]  ( .D(n913), .CP(clk), .CD(n1291), .Q(out1_p1[54])
         );
  CFD2QXL \out0_p2_reg[63]  ( .D(n690), .CP(clk), .CD(n1288), .Q(out0_p2[63])
         );
  CFD2QXL \cmd0_p2_reg[0]  ( .D(n911), .CP(clk), .CD(n1301), .Q(cmd0_p2[0]) );
  CFD2QXL \cmd0_p2_reg[1]  ( .D(n909), .CP(clk), .CD(n1301), .Q(cmd0_p2[1]) );
  CFD2QXL \h0_p1_reg[3]  ( .D(n621), .CP(clk), .CD(n1300), .Q(h0_p1[3]) );
  CFD2QXL push0_reg ( .D(n1344), .CP(clk), .CD(n1301), .Q(push0) );
  CFD2QXL en0_p2_reg ( .D(n907), .CP(clk), .CD(n1288), .Q(en0_p2) );
  CFD2QXL \h0_p1_reg[2]  ( .D(n618), .CP(clk), .CD(n1300), .Q(h0_p1[2]) );
  CFD2QXL en2_p1_reg ( .D(n787), .CP(clk), .CD(n1301), .Q(en2_p1) );
  CFD2QXL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n1301), .Q(cmd0[0]) );
  CFD2QXL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n1302), .Q(cmd0[1]) );
  CFD2QXL \h0_p1_reg[4]  ( .D(n624), .CP(clk), .CD(n1300), .Q(h0_p1[4]) );
  CFD2QXL \h0_p1_reg[1]  ( .D(n615), .CP(clk), .CD(n1300), .Q(h0_p1[1]) );
  CFD2QXL \acc_reg[63]  ( .D(n546), .CP(clk), .CD(n1300), .Q(acc[63]) );
  CFD2QXL \acc_reg[32]  ( .D(n480), .CP(clk), .CD(n1312), .Q(acc[32]) );
  CFD2QXL \acc_reg[33]  ( .D(n478), .CP(clk), .CD(n1312), .Q(acc[33]) );
  CFD2QXL \acc_reg[34]  ( .D(n476), .CP(clk), .CD(n1312), .Q(acc[34]) );
  CFD2QXL \acc_reg[35]  ( .D(n474), .CP(clk), .CD(n1311), .Q(acc[35]) );
  CFD2QXL \acc_reg[36]  ( .D(n472), .CP(clk), .CD(n1311), .Q(acc[36]) );
  CFD2QXL \acc_reg[37]  ( .D(n470), .CP(clk), .CD(n1310), .Q(acc[37]) );
  CFD2QXL \acc_reg[38]  ( .D(n468), .CP(clk), .CD(n1310), .Q(acc[38]) );
  CFD2QXL \acc_reg[39]  ( .D(n466), .CP(clk), .CD(n1310), .Q(acc[39]) );
  CFD2QXL \acc_reg[40]  ( .D(n464), .CP(clk), .CD(n1309), .Q(acc[40]) );
  CFD2QXL \acc_reg[41]  ( .D(n462), .CP(clk), .CD(n1309), .Q(acc[41]) );
  CFD2QXL \acc_reg[42]  ( .D(n460), .CP(clk), .CD(n1308), .Q(acc[42]) );
  CFD2QXL \acc_reg[43]  ( .D(n458), .CP(clk), .CD(n1308), .Q(acc[43]) );
  CFD2QXL \acc_reg[44]  ( .D(n456), .CP(clk), .CD(n1308), .Q(acc[44]) );
  CFD2QXL \acc_reg[45]  ( .D(n454), .CP(clk), .CD(n1307), .Q(acc[45]) );
  CFD2QXL \acc_reg[46]  ( .D(n452), .CP(clk), .CD(n1307), .Q(acc[46]) );
  CFD2QXL \acc_reg[47]  ( .D(n450), .CP(clk), .CD(n1306), .Q(acc[47]) );
  CFD2QXL \acc_reg[48]  ( .D(n448), .CP(clk), .CD(n1306), .Q(acc[48]) );
  CFD2QXL \acc_reg[49]  ( .D(n446), .CP(clk), .CD(n1306), .Q(acc[49]) );
  CFD2QXL \acc_reg[50]  ( .D(n444), .CP(clk), .CD(n1305), .Q(acc[50]) );
  CFD2QXL \acc_reg[51]  ( .D(n442), .CP(clk), .CD(n1305), .Q(acc[51]) );
  CFD2QXL \acc_reg[52]  ( .D(n440), .CP(clk), .CD(n1283), .Q(acc[52]) );
  CFD2QXL \acc_reg[53]  ( .D(n438), .CP(clk), .CD(n1283), .Q(acc[53]) );
  CFD2QXL \acc_reg[54]  ( .D(n436), .CP(clk), .CD(n1282), .Q(acc[54]) );
  CFD2QXL \acc_reg[55]  ( .D(n434), .CP(clk), .CD(n1282), .Q(acc[55]) );
  CFD2QXL \acc_reg[56]  ( .D(n432), .CP(clk), .CD(n1282), .Q(acc[56]) );
  CFD2QXL \acc_reg[57]  ( .D(n430), .CP(clk), .CD(n1281), .Q(acc[57]) );
  CFD2QXL \acc_reg[58]  ( .D(n428), .CP(clk), .CD(n1281), .Q(acc[58]) );
  CFD2QXL \acc_reg[59]  ( .D(n426), .CP(clk), .CD(n1280), .Q(acc[59]) );
  CFD2QXL \acc_reg[60]  ( .D(n424), .CP(clk), .CD(n1280), .Q(acc[60]) );
  CFD2QXL \acc_reg[61]  ( .D(n422), .CP(clk), .CD(n1280), .Q(acc[61]) );
  CFD2QXL \acc_reg[62]  ( .D(n420), .CP(clk), .CD(n1279), .Q(acc[62]) );
  CFD2QXL \h0_p1_reg[0]  ( .D(n612), .CP(clk), .CD(n1300), .Q(h0_p1[0]) );
  CFD1QXL roundit_reg ( .D(n611), .CP(clk), .Q(roundit) );
  CFD2QXL \out1_p1_reg[59]  ( .D(n905), .CP(clk), .CD(n1291), .Q(out1_p1[59])
         );
  CFD2QXL \out1_p1_reg[58]  ( .D(n903), .CP(clk), .CD(n1291), .Q(out1_p1[58])
         );
  CFD2QXL \out1_p1_reg[57]  ( .D(n901), .CP(clk), .CD(n1291), .Q(out1_p1[57])
         );
  CFD2QXL \out1_p1_reg[56]  ( .D(n899), .CP(clk), .CD(n1291), .Q(out1_p1[56])
         );
  CFD2QXL \out1_p1_reg[55]  ( .D(n897), .CP(clk), .CD(n1291), .Q(out1_p1[55])
         );
  CFD2QXL \out1_p1_reg[53]  ( .D(n895), .CP(clk), .CD(n1292), .Q(out1_p1[53])
         );
  CFD2QXL \out1_p1_reg[52]  ( .D(n893), .CP(clk), .CD(n1292), .Q(out1_p1[52])
         );
  CFD2QXL \out1_p1_reg[51]  ( .D(n891), .CP(clk), .CD(n1292), .Q(out1_p1[51])
         );
  CFD2QXL \out1_p1_reg[50]  ( .D(n889), .CP(clk), .CD(n1292), .Q(out1_p1[50])
         );
  CFD2QXL \out1_p1_reg[49]  ( .D(n887), .CP(clk), .CD(n1277), .Q(out1_p1[49])
         );
  CFD2QXL \out1_p1_reg[48]  ( .D(n885), .CP(clk), .CD(n1271), .Q(out1_p1[48])
         );
  CFD2QXL \out1_p1_reg[47]  ( .D(n883), .CP(clk), .CD(n1271), .Q(out1_p1[47])
         );
  CFD2QXL \out1_p1_reg[46]  ( .D(n881), .CP(clk), .CD(n1271), .Q(out1_p1[46])
         );
  CFD2QXL \out1_p1_reg[45]  ( .D(n879), .CP(clk), .CD(n1271), .Q(out1_p1[45])
         );
  CFD2QXL \out1_p1_reg[44]  ( .D(n877), .CP(clk), .CD(n1272), .Q(out1_p1[44])
         );
  CFD2QXL \out1_p1_reg[43]  ( .D(n875), .CP(clk), .CD(n1272), .Q(out1_p1[43])
         );
  CFD2QXL \out1_p1_reg[42]  ( .D(n873), .CP(clk), .CD(n1272), .Q(out1_p1[42])
         );
  CFD2QXL \out1_p1_reg[40]  ( .D(n871), .CP(clk), .CD(n1272), .Q(out1_p1[40])
         );
  CFD2QXL \out1_p1_reg[39]  ( .D(n869), .CP(clk), .CD(n1272), .Q(out1_p1[39])
         );
  CFD2QXL \out1_p1_reg[38]  ( .D(n867), .CP(clk), .CD(n1273), .Q(out1_p1[38])
         );
  CFD2QXL \out1_p1_reg[37]  ( .D(n865), .CP(clk), .CD(n1273), .Q(out1_p1[37])
         );
  CFD2QXL \out1_p1_reg[36]  ( .D(n863), .CP(clk), .CD(n1273), .Q(out1_p1[36])
         );
  CFD2QXL \out1_p1_reg[35]  ( .D(n861), .CP(clk), .CD(n1273), .Q(out1_p1[35])
         );
  CFD2QXL \out1_p1_reg[34]  ( .D(n859), .CP(clk), .CD(n1273), .Q(out1_p1[34])
         );
  CFD2QXL \out1_p1_reg[33]  ( .D(n857), .CP(clk), .CD(n1273), .Q(out1_p1[33])
         );
  CFD2QXL \out1_p1_reg[32]  ( .D(n855), .CP(clk), .CD(n1274), .Q(out1_p1[32])
         );
  CFD2QXL \out1_p1_reg[31]  ( .D(n853), .CP(clk), .CD(n1274), .Q(out1_p1[31])
         );
  CFD2QXL \out1_p1_reg[30]  ( .D(n851), .CP(clk), .CD(n1274), .Q(out1_p1[30])
         );
  CFD2QXL \out1_p1_reg[29]  ( .D(n849), .CP(clk), .CD(n1274), .Q(out1_p1[29])
         );
  CFD2QXL \out1_p1_reg[28]  ( .D(n847), .CP(clk), .CD(n1274), .Q(out1_p1[28])
         );
  CFD2QXL \out1_p1_reg[27]  ( .D(n845), .CP(clk), .CD(n1274), .Q(out1_p1[27])
         );
  CFD2QXL \out1_p1_reg[26]  ( .D(n843), .CP(clk), .CD(n1274), .Q(out1_p1[26])
         );
  CFD2QXL \out1_p1_reg[25]  ( .D(n841), .CP(clk), .CD(n1275), .Q(out1_p1[25])
         );
  CFD2QXL \out1_p1_reg[24]  ( .D(n839), .CP(clk), .CD(n1275), .Q(out1_p1[24])
         );
  CFD2QXL \out1_p1_reg[23]  ( .D(n837), .CP(clk), .CD(n1275), .Q(out1_p1[23])
         );
  CFD2QXL \out1_p1_reg[22]  ( .D(n835), .CP(clk), .CD(n1275), .Q(out1_p1[22])
         );
  CFD2QXL \out1_p1_reg[21]  ( .D(n833), .CP(clk), .CD(n1275), .Q(out1_p1[21])
         );
  CFD2QXL \out1_p1_reg[20]  ( .D(n831), .CP(clk), .CD(n1275), .Q(out1_p1[20])
         );
  CFD2QXL \out1_p1_reg[19]  ( .D(n829), .CP(clk), .CD(n1276), .Q(out1_p1[19])
         );
  CFD2QXL \out1_p1_reg[18]  ( .D(n827), .CP(clk), .CD(n1276), .Q(out1_p1[18])
         );
  CFD2QXL \out1_p1_reg[17]  ( .D(n825), .CP(clk), .CD(n1276), .Q(out1_p1[17])
         );
  CFD2QXL \out1_p1_reg[16]  ( .D(n823), .CP(clk), .CD(n1276), .Q(out1_p1[16])
         );
  CFD2QXL \out1_p1_reg[15]  ( .D(n821), .CP(clk), .CD(n1276), .Q(out1_p1[15])
         );
  CFD2QXL \out1_p1_reg[14]  ( .D(n819), .CP(clk), .CD(n1276), .Q(out1_p1[14])
         );
  CFD2QXL \out1_p1_reg[13]  ( .D(n817), .CP(clk), .CD(n1276), .Q(out1_p1[13])
         );
  CFD2QXL \out1_p1_reg[12]  ( .D(n815), .CP(clk), .CD(n1277), .Q(out1_p1[12])
         );
  CFD2QXL \out1_p1_reg[11]  ( .D(n813), .CP(clk), .CD(n1277), .Q(out1_p1[11])
         );
  CFD2QXL \out1_p1_reg[10]  ( .D(n811), .CP(clk), .CD(n1277), .Q(out1_p1[10])
         );
  CFD2QXL \out1_p1_reg[9]  ( .D(n809), .CP(clk), .CD(n1277), .Q(out1_p1[9]) );
  CFD2QXL \out1_p1_reg[8]  ( .D(n807), .CP(clk), .CD(n1277), .Q(out1_p1[8]) );
  CFD2QXL \out1_p1_reg[7]  ( .D(n805), .CP(clk), .CD(n1277), .Q(out1_p1[7]) );
  CFD2QXL \out1_p1_reg[6]  ( .D(n803), .CP(clk), .CD(n1278), .Q(out1_p1[6]) );
  CFD2QXL \out1_p1_reg[5]  ( .D(n801), .CP(clk), .CD(n1278), .Q(out1_p1[5]) );
  CFD2QXL \out1_p1_reg[4]  ( .D(n799), .CP(clk), .CD(n1278), .Q(out1_p1[4]) );
  CFD2QXL \out1_p1_reg[3]  ( .D(n797), .CP(clk), .CD(n1278), .Q(out1_p1[3]) );
  CFD2QXL \out1_p1_reg[2]  ( .D(n795), .CP(clk), .CD(n1278), .Q(out1_p1[2]) );
  CFD2QXL \out1_p1_reg[1]  ( .D(n793), .CP(clk), .CD(n1278), .Q(out1_p1[1]) );
  CFD2QXL \out1_p1_reg[0]  ( .D(n791), .CP(clk), .CD(n1279), .Q(out1_p1[0]) );
  CFD2QXL \out0_p2_reg[0]  ( .D(n753), .CP(clk), .CD(n1300), .Q(out0_p2[0]) );
  CFD2QXL \out0_p2_reg[1]  ( .D(n752), .CP(clk), .CD(n1299), .Q(out0_p2[1]) );
  CFD2QXL \out0_p2_reg[2]  ( .D(n751), .CP(clk), .CD(n1299), .Q(out0_p2[2]) );
  CFD2QXL \out0_p2_reg[3]  ( .D(n750), .CP(clk), .CD(n1299), .Q(out0_p2[3]) );
  CFD2QXL \out0_p2_reg[4]  ( .D(n749), .CP(clk), .CD(n1298), .Q(out0_p2[4]) );
  CFD2QXL \out0_p2_reg[5]  ( .D(n748), .CP(clk), .CD(n1298), .Q(out0_p2[5]) );
  CFD2QXL \out0_p2_reg[6]  ( .D(n747), .CP(clk), .CD(n1297), .Q(out0_p2[6]) );
  CFD2QXL \out0_p2_reg[7]  ( .D(n746), .CP(clk), .CD(n1297), .Q(out0_p2[7]) );
  CFD2QXL \out0_p2_reg[8]  ( .D(n745), .CP(clk), .CD(n1297), .Q(out0_p2[8]) );
  CFD2QXL \out0_p2_reg[9]  ( .D(n744), .CP(clk), .CD(n1296), .Q(out0_p2[9]) );
  CFD2QXL \out0_p2_reg[10]  ( .D(n743), .CP(clk), .CD(n1296), .Q(out0_p2[10])
         );
  CFD2QXL \out0_p2_reg[11]  ( .D(n742), .CP(clk), .CD(n1295), .Q(out0_p2[11])
         );
  CFD2QXL \out0_p2_reg[12]  ( .D(n741), .CP(clk), .CD(n1295), .Q(out0_p2[12])
         );
  CFD2QXL \out0_p2_reg[13]  ( .D(n740), .CP(clk), .CD(n1295), .Q(out0_p2[13])
         );
  CFD2QXL \out0_p2_reg[14]  ( .D(n739), .CP(clk), .CD(n1294), .Q(out0_p2[14])
         );
  CFD2QXL \out0_p2_reg[15]  ( .D(n738), .CP(clk), .CD(n1294), .Q(out0_p2[15])
         );
  CFD2QXL \out0_p2_reg[16]  ( .D(n737), .CP(clk), .CD(n1294), .Q(out0_p2[16])
         );
  CFD2QXL \out0_p2_reg[17]  ( .D(n736), .CP(clk), .CD(n1293), .Q(out0_p2[17])
         );
  CFD2QXL \out0_p2_reg[18]  ( .D(n735), .CP(clk), .CD(n1293), .Q(out0_p2[18])
         );
  CFD2QXL \out0_p2_reg[19]  ( .D(n734), .CP(clk), .CD(n1292), .Q(out0_p2[19])
         );
  CFD2QXL \out0_p2_reg[20]  ( .D(n733), .CP(clk), .CD(n1317), .Q(out0_p2[20])
         );
  CFD2QXL \out0_p2_reg[21]  ( .D(n732), .CP(clk), .CD(n1316), .Q(out0_p2[21])
         );
  CFD2QXL \out0_p2_reg[22]  ( .D(n731), .CP(clk), .CD(n1316), .Q(out0_p2[22])
         );
  CFD2QXL \out0_p2_reg[23]  ( .D(n730), .CP(clk), .CD(n1316), .Q(out0_p2[23])
         );
  CFD2QXL \out0_p2_reg[24]  ( .D(n729), .CP(clk), .CD(n1315), .Q(out0_p2[24])
         );
  CFD2QXL \out0_p2_reg[25]  ( .D(n728), .CP(clk), .CD(n1315), .Q(out0_p2[25])
         );
  CFD2QXL \out0_p2_reg[26]  ( .D(n727), .CP(clk), .CD(n1313), .Q(out0_p2[26])
         );
  CFD2QXL \out0_p2_reg[27]  ( .D(n726), .CP(clk), .CD(n1314), .Q(out0_p2[27])
         );
  CFD2QXL \out0_p2_reg[28]  ( .D(n725), .CP(clk), .CD(n1314), .Q(out0_p2[28])
         );
  CFD2QXL \out0_p2_reg[29]  ( .D(n724), .CP(clk), .CD(n1313), .Q(out0_p2[29])
         );
  CFD2QXL \out0_p2_reg[30]  ( .D(n723), .CP(clk), .CD(n1313), .Q(out0_p2[30])
         );
  CFD2QXL \out0_p2_reg[31]  ( .D(n722), .CP(clk), .CD(n1313), .Q(out0_p2[31])
         );
  CFD2QXL \out0_p2_reg[32]  ( .D(n721), .CP(clk), .CD(n1312), .Q(out0_p2[32])
         );
  CFD2QXL \out0_p2_reg[33]  ( .D(n720), .CP(clk), .CD(n1312), .Q(out0_p2[33])
         );
  CFD2QXL \out0_p2_reg[34]  ( .D(n719), .CP(clk), .CD(n1311), .Q(out0_p2[34])
         );
  CFD2QXL \out0_p2_reg[35]  ( .D(n718), .CP(clk), .CD(n1311), .Q(out0_p2[35])
         );
  CFD2QXL \out0_p2_reg[36]  ( .D(n717), .CP(clk), .CD(n1311), .Q(out0_p2[36])
         );
  CFD2QXL \out0_p2_reg[37]  ( .D(n716), .CP(clk), .CD(n1310), .Q(out0_p2[37])
         );
  CFD2QXL \out0_p2_reg[38]  ( .D(n715), .CP(clk), .CD(n1310), .Q(out0_p2[38])
         );
  CFD2QXL \out0_p2_reg[39]  ( .D(n714), .CP(clk), .CD(n1309), .Q(out0_p2[39])
         );
  CFD2QXL \out0_p2_reg[40]  ( .D(n713), .CP(clk), .CD(n1309), .Q(out0_p2[40])
         );
  CFD2QXL \out0_p2_reg[41]  ( .D(n712), .CP(clk), .CD(n1309), .Q(out0_p2[41])
         );
  CFD2QXL \out0_p2_reg[42]  ( .D(n711), .CP(clk), .CD(n1308), .Q(out0_p2[42])
         );
  CFD2QXL \out0_p2_reg[43]  ( .D(n710), .CP(clk), .CD(n1308), .Q(out0_p2[43])
         );
  CFD2QXL \out0_p2_reg[44]  ( .D(n709), .CP(clk), .CD(n1307), .Q(out0_p2[44])
         );
  CFD2QXL \out0_p2_reg[45]  ( .D(n708), .CP(clk), .CD(n1307), .Q(out0_p2[45])
         );
  CFD2QXL \out0_p2_reg[46]  ( .D(n707), .CP(clk), .CD(n1307), .Q(out0_p2[46])
         );
  CFD2QXL \out0_p2_reg[47]  ( .D(n706), .CP(clk), .CD(n1306), .Q(out0_p2[47])
         );
  CFD2QXL \out0_p2_reg[48]  ( .D(n705), .CP(clk), .CD(n1306), .Q(out0_p2[48])
         );
  CFD2QXL \out0_p2_reg[49]  ( .D(n704), .CP(clk), .CD(n1306), .Q(out0_p2[49])
         );
  CFD2QXL \out0_p2_reg[50]  ( .D(n703), .CP(clk), .CD(n1305), .Q(out0_p2[50])
         );
  CFD2QXL \out0_p2_reg[51]  ( .D(n702), .CP(clk), .CD(n1305), .Q(out0_p2[51])
         );
  CFD2QXL \out0_p2_reg[52]  ( .D(n701), .CP(clk), .CD(n1283), .Q(out0_p2[52])
         );
  CFD2QXL \out0_p2_reg[53]  ( .D(n700), .CP(clk), .CD(n1283), .Q(out0_p2[53])
         );
  CFD2QXL \out0_p2_reg[54]  ( .D(n699), .CP(clk), .CD(n1282), .Q(out0_p2[54])
         );
  CFD2QXL \out0_p2_reg[55]  ( .D(n698), .CP(clk), .CD(n1282), .Q(out0_p2[55])
         );
  CFD2QXL \out0_p2_reg[56]  ( .D(n697), .CP(clk), .CD(n1281), .Q(out0_p2[56])
         );
  CFD2QXL \out0_p2_reg[57]  ( .D(n696), .CP(clk), .CD(n1281), .Q(out0_p2[57])
         );
  CFD2QXL \out0_p2_reg[58]  ( .D(n695), .CP(clk), .CD(n1281), .Q(out0_p2[58])
         );
  CFD2QXL \out0_p2_reg[59]  ( .D(n694), .CP(clk), .CD(n1280), .Q(out0_p2[59])
         );
  CFD2QXL \out0_p2_reg[60]  ( .D(n693), .CP(clk), .CD(n1280), .Q(out0_p2[60])
         );
  CFD2QXL \out0_p2_reg[61]  ( .D(n692), .CP(clk), .CD(n1279), .Q(out0_p2[61])
         );
  CFD2QXL \out0_p2_reg[62]  ( .D(n691), .CP(clk), .CD(n1279), .Q(out0_p2[62])
         );
  CFD2QXL \out1_p2_reg[0]  ( .D(n545), .CP(clk), .CD(n1300), .Q(out1_p2[0]) );
  CFD2QXL \out1_p2_reg[1]  ( .D(n543), .CP(clk), .CD(n1299), .Q(out1_p2[1]) );
  CFD2QXL \out1_p2_reg[2]  ( .D(n541), .CP(clk), .CD(n1299), .Q(out1_p2[2]) );
  CFD2QXL \out1_p2_reg[3]  ( .D(n539), .CP(clk), .CD(n1299), .Q(out1_p2[3]) );
  CFD2QXL \out1_p2_reg[4]  ( .D(n537), .CP(clk), .CD(n1298), .Q(out1_p2[4]) );
  CFD2QXL \out1_p2_reg[5]  ( .D(n535), .CP(clk), .CD(n1298), .Q(out1_p2[5]) );
  CFD2QXL \out1_p2_reg[6]  ( .D(n533), .CP(clk), .CD(n1297), .Q(out1_p2[6]) );
  CFD2QXL \out1_p2_reg[7]  ( .D(n531), .CP(clk), .CD(n1297), .Q(out1_p2[7]) );
  CFD2QXL \out1_p2_reg[8]  ( .D(n529), .CP(clk), .CD(n1297), .Q(out1_p2[8]) );
  CFD2QXL \out1_p2_reg[9]  ( .D(n527), .CP(clk), .CD(n1296), .Q(out1_p2[9]) );
  CFD2QXL \out1_p2_reg[16]  ( .D(n513), .CP(clk), .CD(n1294), .Q(out1_p2[16])
         );
  CFD2QXL \acc_reg[0]  ( .D(n544), .CP(clk), .CD(n1300), .Q(acc[0]) );
  CFD2QXL \acc_reg[1]  ( .D(n542), .CP(clk), .CD(n1299), .Q(acc[1]) );
  CFD2QXL \acc_reg[2]  ( .D(n540), .CP(clk), .CD(n1299), .Q(acc[2]) );
  CFD2QXL \acc_reg[3]  ( .D(n538), .CP(clk), .CD(n1299), .Q(acc[3]) );
  CFD2QXL \acc_reg[4]  ( .D(n536), .CP(clk), .CD(n1298), .Q(acc[4]) );
  CFD2QXL \acc_reg[5]  ( .D(n534), .CP(clk), .CD(n1298), .Q(acc[5]) );
  CFD2QXL \acc_reg[6]  ( .D(n532), .CP(clk), .CD(n1298), .Q(acc[6]) );
  CFD2QXL \acc_reg[7]  ( .D(n530), .CP(clk), .CD(n1297), .Q(acc[7]) );
  CFD2QXL \acc_reg[8]  ( .D(n528), .CP(clk), .CD(n1297), .Q(acc[8]) );
  CFD2QXL \acc_reg[9]  ( .D(n526), .CP(clk), .CD(n1296), .Q(acc[9]) );
  CFD2QXL \acc_reg[10]  ( .D(n524), .CP(clk), .CD(n1296), .Q(acc[10]) );
  CFD2QXL \acc_reg[11]  ( .D(n522), .CP(clk), .CD(n1296), .Q(acc[11]) );
  CFD2QXL \acc_reg[12]  ( .D(n520), .CP(clk), .CD(n1295), .Q(acc[12]) );
  CFD2QXL \acc_reg[13]  ( .D(n518), .CP(clk), .CD(n1295), .Q(acc[13]) );
  CFD2QXL \acc_reg[14]  ( .D(n516), .CP(clk), .CD(n1294), .Q(acc[14]) );
  CFD2QXL \acc_reg[15]  ( .D(n514), .CP(clk), .CD(n1294), .Q(acc[15]) );
  CFD2QXL \acc_reg[16]  ( .D(n512), .CP(clk), .CD(n1294), .Q(acc[16]) );
  CFD2QXL \acc_reg[17]  ( .D(n510), .CP(clk), .CD(n1293), .Q(acc[17]) );
  CFD2QXL \acc_reg[18]  ( .D(n508), .CP(clk), .CD(n1293), .Q(acc[18]) );
  CFD2QXL \acc_reg[19]  ( .D(n506), .CP(clk), .CD(n1293), .Q(acc[19]) );
  CFD2QXL \acc_reg[20]  ( .D(n504), .CP(clk), .CD(n1316), .Q(acc[20]) );
  CFD2QXL \acc_reg[21]  ( .D(n502), .CP(clk), .CD(n1317), .Q(acc[21]) );
  CFD2QXL \acc_reg[22]  ( .D(n500), .CP(clk), .CD(n1316), .Q(acc[22]) );
  CFD2QXL \acc_reg[23]  ( .D(n498), .CP(clk), .CD(n1316), .Q(acc[23]) );
  CFD2QXL \acc_reg[24]  ( .D(n496), .CP(clk), .CD(n1315), .Q(acc[24]) );
  CFD2QXL \acc_reg[25]  ( .D(n494), .CP(clk), .CD(n1315), .Q(acc[25]) );
  CFD2QXL \acc_reg[26]  ( .D(n492), .CP(clk), .CD(n1315), .Q(acc[26]) );
  CFD2QXL \acc_reg[27]  ( .D(n490), .CP(clk), .CD(n1314), .Q(acc[27]) );
  CFD2QXL \acc_reg[28]  ( .D(n488), .CP(clk), .CD(n1314), .Q(acc[28]) );
  CFD2QXL \acc_reg[29]  ( .D(n486), .CP(clk), .CD(n1314), .Q(acc[29]) );
  CFD2QXL \acc_reg[30]  ( .D(n484), .CP(clk), .CD(n1313), .Q(acc[30]) );
  CFD2QXL \acc_reg[31]  ( .D(n482), .CP(clk), .CD(n1313), .Q(acc[31]) );
  CFD2QXL en1_p1_reg ( .D(en1_p0), .CP(clk), .CD(n1279), .Q(en1_p1) );
  CFD2QXL en0_p1_reg ( .D(en0_p0), .CP(clk), .CD(n1288), .Q(en0_p1) );
  CFD2QXL _pushout_reg ( .D(n789), .CP(clk), .CD(n1301), .Q(pushout) );
  CFD2QXL \out0_p0_reg[63]  ( .D(N77), .CP(clk), .CD(n1287), .Q(out0_p0[63])
         );
  CFD2QXL \out0_p0_reg[41]  ( .D(N55), .CP(clk), .CD(n1308), .Q(out0_p0[41])
         );
  CFD2QXL \out0_p0_reg[40]  ( .D(N54), .CP(clk), .CD(n1309), .Q(out0_p0[40])
         );
  CFD2QXL \out0_p0_reg[39]  ( .D(N53), .CP(clk), .CD(n1309), .Q(out0_p0[39])
         );
  CFD2QXL \out0_p0_reg[38]  ( .D(N52), .CP(clk), .CD(n1310), .Q(out0_p0[38])
         );
  CFD2QXL \out0_p0_reg[37]  ( .D(N51), .CP(clk), .CD(n1310), .Q(out0_p0[37])
         );
  CFD2QXL \out0_p0_reg[36]  ( .D(N50), .CP(clk), .CD(n1310), .Q(out0_p0[36])
         );
  CFD2QXL \out0_p0_reg[35]  ( .D(N49), .CP(clk), .CD(n1311), .Q(out0_p0[35])
         );
  CFD2QXL \out0_p0_reg[34]  ( .D(N48), .CP(clk), .CD(n1311), .Q(out0_p0[34])
         );
  CFD2QXL \out0_p0_reg[33]  ( .D(N47), .CP(clk), .CD(n1312), .Q(out0_p0[33])
         );
  CFD2QXL \out0_p0_reg[32]  ( .D(N46), .CP(clk), .CD(n1311), .Q(out0_p0[32])
         );
  CFD2QXL \out0_p0_reg[31]  ( .D(N45), .CP(clk), .CD(n1312), .Q(out0_p0[31])
         );
  CFD2QXL \out0_p0_reg[30]  ( .D(N44), .CP(clk), .CD(n1313), .Q(out0_p0[30])
         );
  CFD2QXL \out0_p0_reg[29]  ( .D(N43), .CP(clk), .CD(n1313), .Q(out0_p0[29])
         );
  CFD2QXL \out0_p0_reg[27]  ( .D(N41), .CP(clk), .CD(n1314), .Q(out0_p0[27])
         );
  CFD2QXL \out0_p0_reg[26]  ( .D(N40), .CP(clk), .CD(n1314), .Q(out0_p0[26])
         );
  CFD2QXL \out0_p0_reg[25]  ( .D(N39), .CP(clk), .CD(n1315), .Q(out0_p0[25])
         );
  CFD2QXL \out0_p0_reg[24]  ( .D(N38), .CP(clk), .CD(n1315), .Q(out0_p0[24])
         );
  CFD2QXL \out0_p0_reg[23]  ( .D(N37), .CP(clk), .CD(n1316), .Q(out0_p0[23])
         );
  CFD2QXL \out0_p0_reg[22]  ( .D(N36), .CP(clk), .CD(n1316), .Q(out0_p0[22])
         );
  CFD2QXL \out0_p0_reg[17]  ( .D(N31), .CP(clk), .CD(n1293), .Q(out0_p0[17])
         );
  CFD2QXL \out0_p0_reg[16]  ( .D(N30), .CP(clk), .CD(n1293), .Q(out0_p0[16])
         );
  CFD2QXL \out0_p0_reg[9]  ( .D(N23), .CP(clk), .CD(n1296), .Q(out0_p0[9]) );
  CFD2QXL \out0_p0_reg[8]  ( .D(N22), .CP(clk), .CD(n1296), .Q(out0_p0[8]) );
  CFD2QXL \out0_p0_reg[7]  ( .D(N21), .CP(clk), .CD(n1297), .Q(out0_p0[7]) );
  CFD2QXL \out0_p0_reg[6]  ( .D(N20), .CP(clk), .CD(n1297), .Q(out0_p0[6]) );
  CFD2QXL \out0_p0_reg[5]  ( .D(N19), .CP(clk), .CD(n1298), .Q(out0_p0[5]) );
  CFD2QXL \out0_p0_reg[4]  ( .D(N18), .CP(clk), .CD(n1298), .Q(out0_p0[4]) );
  CFD2QXL \out0_p0_reg[3]  ( .D(N17), .CP(clk), .CD(n1298), .Q(out0_p0[3]) );
  CFD2QXL \out0_p0_reg[2]  ( .D(N16), .CP(clk), .CD(n1299), .Q(out0_p0[2]) );
  CFD2QXL \out0_p0_reg[1]  ( .D(N15), .CP(clk), .CD(n1299), .Q(out0_p0[1]) );
  CFD2QXL \out0_p0_reg[0]  ( .D(N14), .CP(clk), .CD(n1300), .Q(out0_p0[0]) );
  CFD2QXL \out1_p0_reg[63]  ( .D(N77), .CP(clk), .CD(n1290), .Q(out1_p0[63])
         );
  CFD2QXL \out1_p0_reg[40]  ( .D(N54), .CP(clk), .CD(n1272), .Q(out1_p0[40])
         );
  CFD2QXL \out1_p0_reg[39]  ( .D(N53), .CP(clk), .CD(n1273), .Q(out1_p0[39])
         );
  CFD2QXL \out1_p0_reg[38]  ( .D(N52), .CP(clk), .CD(n1272), .Q(out1_p0[38])
         );
  CFD2QXL \out1_p0_reg[37]  ( .D(N51), .CP(clk), .CD(n1273), .Q(out1_p0[37])
         );
  CFD2QXL \out1_p0_reg[36]  ( .D(N50), .CP(clk), .CD(n1273), .Q(out1_p0[36])
         );
  CFD2QXL \out1_p0_reg[35]  ( .D(N49), .CP(clk), .CD(n1273), .Q(out1_p0[35])
         );
  CFD2QXL \out1_p0_reg[34]  ( .D(N48), .CP(clk), .CD(n1273), .Q(out1_p0[34])
         );
  CFD2QXL \out1_p0_reg[33]  ( .D(N47), .CP(clk), .CD(n1273), .Q(out1_p0[33])
         );
  CFD2QXL \out1_p0_reg[32]  ( .D(N46), .CP(clk), .CD(n1273), .Q(out1_p0[32])
         );
  CFD2QXL \out1_p0_reg[31]  ( .D(N45), .CP(clk), .CD(n1274), .Q(out1_p0[31])
         );
  CFD2QXL \out1_p0_reg[30]  ( .D(N44), .CP(clk), .CD(n1274), .Q(out1_p0[30])
         );
  CFD2QXL \out1_p0_reg[29]  ( .D(N43), .CP(clk), .CD(n1274), .Q(out1_p0[29])
         );
  CFD2QXL \out1_p0_reg[27]  ( .D(N41), .CP(clk), .CD(n1274), .Q(out1_p0[27])
         );
  CFD2QXL \out1_p0_reg[26]  ( .D(N40), .CP(clk), .CD(n1274), .Q(out1_p0[26])
         );
  CFD2QXL \out1_p0_reg[25]  ( .D(N39), .CP(clk), .CD(n1275), .Q(out1_p0[25])
         );
  CFD2QXL \out1_p0_reg[24]  ( .D(N38), .CP(clk), .CD(n1275), .Q(out1_p0[24])
         );
  CFD2QXL \out1_p0_reg[23]  ( .D(N37), .CP(clk), .CD(n1275), .Q(out1_p0[23])
         );
  CFD2QXL \out1_p0_reg[22]  ( .D(N36), .CP(clk), .CD(n1275), .Q(out1_p0[22])
         );
  CFD2QXL \out1_p0_reg[17]  ( .D(N31), .CP(clk), .CD(n1276), .Q(out1_p0[17])
         );
  CFD2QXL \out1_p0_reg[16]  ( .D(N30), .CP(clk), .CD(n1276), .Q(out1_p0[16])
         );
  CFD2QXL \out1_p0_reg[9]  ( .D(N23), .CP(clk), .CD(n1277), .Q(out1_p0[9]) );
  CFD2QXL \out1_p0_reg[8]  ( .D(N22), .CP(clk), .CD(n1277), .Q(out1_p0[8]) );
  CFD2QXL \out1_p0_reg[7]  ( .D(N21), .CP(clk), .CD(n1277), .Q(out1_p0[7]) );
  CFD2QXL \out1_p0_reg[6]  ( .D(N20), .CP(clk), .CD(n1278), .Q(out1_p0[6]) );
  CFD2QXL \out1_p0_reg[5]  ( .D(N19), .CP(clk), .CD(n1278), .Q(out1_p0[5]) );
  CFD2QXL \out1_p0_reg[4]  ( .D(N18), .CP(clk), .CD(n1278), .Q(out1_p0[4]) );
  CFD2QXL \out1_p0_reg[3]  ( .D(N17), .CP(clk), .CD(n1278), .Q(out1_p0[3]) );
  CFD2QXL \out1_p0_reg[2]  ( .D(N16), .CP(clk), .CD(n1278), .Q(out1_p0[2]) );
  CFD2QXL \out1_p0_reg[1]  ( .D(N15), .CP(clk), .CD(n1278), .Q(out1_p0[1]) );
  CFD2QXL \out1_p0_reg[0]  ( .D(N14), .CP(clk), .CD(n1278), .Q(out1_p0[0]) );
  CFD2QXL \cmd0_p0_reg[1]  ( .D(n1063), .CP(clk), .CD(n1301), .Q(cmd0_p0[1])
         );
  CFD2QXL \cmd0_p1_reg[1]  ( .D(n1064), .CP(clk), .CD(n1301), .Q(cmd0_p1[1])
         );
  CFD2QXL \cmd0_p0_reg[0]  ( .D(n1066), .CP(clk), .CD(n1301), .Q(cmd0_p0[0])
         );
  CFD2QXL \cmd0_p1_reg[0]  ( .D(n1067), .CP(clk), .CD(n1301), .Q(cmd0_p1[0])
         );
  CFD2QXL push0_p0_reg ( .D(n1069), .CP(clk), .CD(n1301), .Q(push0_p0) );
  CFD2QXL push0_p1_reg ( .D(n1071), .CP(clk), .CD(n1301), .Q(push0_p1) );
  CFD2QX1 \h0_reg[0]  ( .D(n614), .CP(clk), .CD(n1287), .Q(h0[0]) );
  CFD2QX2 \q0_reg[1]  ( .D(n659), .CP(clk), .CD(n1271), .Q(q0[1]) );
  CFD2QX1 \q0_reg[21]  ( .D(n679), .CP(clk), .CD(n1271), .Q(q0[21]) );
  CFD2QXL en1_p2_d1_reg ( .D(n1261), .CP(clk), .CD(n1279), .Q(en1_p2_d1) );
  CFD2QXL en0_p2_d1_reg ( .D(n1256), .CP(clk), .CD(n1279), .Q(en0_p2_d1) );
  CFD2QXL en2_p2_reg ( .D(en2_p1), .CP(clk), .CD(n1288), .Q(en2_p2) );
  CFD2QX1 \q0_reg[31]  ( .D(n790), .CP(clk), .CD(n1292), .Q(q0[31]) );
  CFD2QX1 \q0_reg[17]  ( .D(n675), .CP(clk), .CD(n1284), .Q(q0[17]) );
  CFD2QX2 \h0_reg[5]  ( .D(n629), .CP(clk), .CD(n1287), .Q(h0[5]) );
  CFD2QX1 \h0_reg[1]  ( .D(n617), .CP(clk), .CD(n1287), .Q(h0[1]) );
  CFD2QX2 \h0_reg[2]  ( .D(n620), .CP(clk), .CD(n1287), .Q(h0[2]) );
  CFD2QX4 \h0_reg[3]  ( .D(n623), .CP(clk), .CD(n1287), .Q(h0[3]) );
  CFD2QX1 \h0_reg[4]  ( .D(n626), .CP(clk), .CD(n1287), .Q(h0[4]) );
  CFD2QX4 \h0_reg[20]  ( .D(n646), .CP(clk), .CD(n1286), .Q(h0[20]) );
  CFD2QX4 \h0_reg[29]  ( .D(n655), .CP(clk), .CD(n1285), .Q(h0[29]) );
  CFD2QX4 \h0_reg[28]  ( .D(n654), .CP(clk), .CD(n1285), .Q(h0[28]) );
  CFD2QX4 \h0_reg[30]  ( .D(n656), .CP(clk), .CD(n1285), .Q(h0[30]) );
  CFD2QX4 \h0_reg[17]  ( .D(n643), .CP(clk), .CD(n1286), .Q(h0[17]) );
  CFD2QX1 \h0_reg[12]  ( .D(n1074), .CP(clk), .CD(n1286), .Q(h0[12]) );
  CFD2QX1 \h0_reg[21]  ( .D(n1083), .CP(clk), .CD(n1286), .Q(h0[21]) );
  CFD2QX4 \h0_reg[27]  ( .D(n653), .CP(clk), .CD(n1285), .Q(h0[27]) );
  CFD2QX4 \h0_reg[19]  ( .D(n645), .CP(clk), .CD(n1286), .Q(h0[19]) );
  CFD2QX4 \h0_reg[22]  ( .D(n648), .CP(clk), .CD(n1286), .Q(h0[22]) );
  CFD2QX1 \h0_reg[15]  ( .D(n1080), .CP(clk), .CD(n1286), .Q(h0[15]) );
  CFD2QX4 \h0_reg[18]  ( .D(n644), .CP(clk), .CD(n1286), .Q(h0[18]) );
  CFD2QX1 \h0_reg[24]  ( .D(n1079), .CP(clk), .CD(n1286), .Q(h0[24]) );
  CFD2QX1 \h0_reg[13]  ( .D(n1077), .CP(clk), .CD(n1286), .Q(h0[13]) );
  CFD2QX4 \h0_reg[7]  ( .D(n633), .CP(clk), .CD(n1287), .Q(h0[7]) );
  CFD2QX1 \h0_reg[26]  ( .D(n1062), .CP(clk), .CD(n1285), .Q(h0[26]) );
  CFD2QX1 \h0_reg[10]  ( .D(n1081), .CP(clk), .CD(n1287), .Q(h0[10]) );
  CFD2QX1 \h0_reg[11]  ( .D(n1082), .CP(clk), .CD(n1287), .Q(h0[11]) );
  CFD2QX1 \q0_reg[22]  ( .D(n1078), .CP(clk), .CD(n1283), .Q(q0[22]) );
  CFD2QX4 \q0_reg[16]  ( .D(n674), .CP(clk), .CD(n1284), .Q(q0[16]) );
  CFD2QX1 \h0_reg[14]  ( .D(n1086), .CP(clk), .CD(n1286), .Q(h0[14]) );
  CFD2QX1 \h0_reg[16]  ( .D(n1085), .CP(clk), .CD(n1286), .Q(h0[16]) );
  CFD2QX1 \h0_reg[8]  ( .D(n1084), .CP(clk), .CD(n1287), .Q(h0[8]) );
  CFD2QX1 \h0_reg[9]  ( .D(n1154), .CP(clk), .CD(n1287), .Q(h0[9]) );
  CFD2QX1 \q0_reg[9]  ( .D(n667), .CP(clk), .CD(n1284), .Q(q0[9]) );
  CFD2QX1 \h0_reg[23]  ( .D(n1144), .CP(clk), .CD(n1286), .Q(h0[23]) );
  CFD2QX1 \q0_reg[23]  ( .D(n681), .CP(clk), .CD(n1271), .Q(q0[23]) );
  CFD2QX1 \h0_reg[25]  ( .D(n1157), .CP(clk), .CD(n1285), .Q(h0[25]) );
  CFD2QX1 \h0_reg[31]  ( .D(n1156), .CP(clk), .CD(n1285), .Q(h0[31]) );
  CFD2QX1 \q0_reg[6]  ( .D(n664), .CP(clk), .CD(n1285), .Q(q0[6]) );
  CFD2QX4 \q0_reg[28]  ( .D(n686), .CP(clk), .CD(n1289), .Q(q0[28]) );
  CFD2QX2 \q0_reg[11]  ( .D(n669), .CP(clk), .CD(n1284), .Q(q0[11]) );
  CFD2QX2 \q0_reg[26]  ( .D(n684), .CP(clk), .CD(n1283), .Q(q0[26]) );
  CFD2QX2 \q0_reg[10]  ( .D(n668), .CP(clk), .CD(n1284), .Q(q0[10]) );
  CFD2QX2 \q0_reg[18]  ( .D(n676), .CP(clk), .CD(n1284), .Q(q0[18]) );
  CFD2XL \out1_p2_reg[14]  ( .D(n517), .CP(clk), .CD(n1937), .Q(out1_p2[14]), 
        .QN(n1663) );
  CFD2XL \out1_p2_reg[12]  ( .D(n521), .CP(clk), .CD(n1937), .Q(out1_p2[12]), 
        .QN(n1671) );
  CFD2XL \out1_p2_reg[10]  ( .D(n525), .CP(clk), .CD(n1937), .Q(out1_p2[10]), 
        .QN(n1679) );
  CFD2XL \out1_p0_reg[11]  ( .D(N25), .CP(clk), .CD(n1937), .Q(out1_p0[11]) );
  CFD2XL \out0_p0_reg[11]  ( .D(N25), .CP(clk), .CD(n1937), .Q(out0_p0[11]) );
  CFD2XL \out2_p2_reg[55]  ( .D(n1143), .CP(clk), .CD(n1937), .Q(out2_p2[55]), 
        .QN(n1346) );
  CFD2XL \out1_p0_reg[10]  ( .D(N24), .CP(clk), .CD(n1937), .Q(out1_p0[10]) );
  CFD2XL \out0_p0_reg[10]  ( .D(N24), .CP(clk), .CD(n1937), .Q(out0_p0[10]) );
  CFD2XL \out2_p2_reg[49]  ( .D(n1146), .CP(clk), .CD(n1937), .Q(out2_p2[49]), 
        .QN(n1358) );
  CFD2XL \out2_p2_reg[53]  ( .D(n1150), .CP(clk), .CD(n1937), .Q(out2_p2[53]), 
        .QN(n1350) );
  CFD2XL \out1_p2_reg[32]  ( .D(n481), .CP(clk), .CD(n1937), .Q(out1_p2[32]), 
        .QN(n1591) );
  CFD2XL \out2_p2_reg[23]  ( .D(n1149), .CP(clk), .CD(n1937), .Q(out2_p2[23]), 
        .QN(n1413) );
  CFD2XL \out2_p2_reg[47]  ( .D(n1153), .CP(clk), .CD(n1937), .Q(out2_p2[47]), 
        .QN(n1362) );
  CFD2XL \out2_p2_reg[39]  ( .D(n1148), .CP(clk), .CD(n1937), .Q(out2_p2[39]), 
        .QN(n1378) );
  CFD2XL \out2_p2_reg[31]  ( .D(n1147), .CP(clk), .CD(n1937), .Q(out2_p2[31]), 
        .QN(n1397) );
  CFD2XL \out2_p2_reg[21]  ( .D(n1145), .CP(clk), .CD(n1937), .Q(out2_p2[21]), 
        .QN(n1417) );
  CFD2XL \out2_p2_reg[17]  ( .D(n1151), .CP(clk), .CD(n1937), .Q(out2_p2[17]), 
        .QN(n1425) );
  CFD2XL \out2_p2_reg[15]  ( .D(n1152), .CP(clk), .CD(n1937), .Q(out2_p2[15]), 
        .QN(n1429) );
  CFD2XL \out1_p2_reg[31]  ( .D(n483), .CP(clk), .CD(n1937), .Q(out1_p2[31]), 
        .QN(n1595) );
  CFD2XL \out1_p2_reg[30]  ( .D(n485), .CP(clk), .CD(n1937), .Q(out1_p2[30]), 
        .QN(n1599) );
  CFD2XL \out1_p2_reg[29]  ( .D(n487), .CP(clk), .CD(n1937), .Q(out1_p2[29]), 
        .QN(n1603) );
  CFD2XL \out1_p2_reg[28]  ( .D(n489), .CP(clk), .CD(n1937), .Q(out1_p2[28]), 
        .QN(n1607) );
  CFD2XL \out1_p2_reg[27]  ( .D(n491), .CP(clk), .CD(n1937), .Q(out1_p2[27]), 
        .QN(n1611) );
  CFD2XL \out1_p2_reg[26]  ( .D(n493), .CP(clk), .CD(n1937), .Q(out1_p2[26]), 
        .QN(n1615) );
  CFD2XL \out1_p2_reg[25]  ( .D(n495), .CP(clk), .CD(n1937), .Q(out1_p2[25]), 
        .QN(n1619) );
  CFD2XL \out1_p2_reg[24]  ( .D(n497), .CP(clk), .CD(n1937), .Q(out1_p2[24]), 
        .QN(n1623) );
  CFD2XL \out1_p2_reg[23]  ( .D(n499), .CP(clk), .CD(n1937), .Q(out1_p2[23]), 
        .QN(n1627) );
  CFD2XL \out1_p2_reg[22]  ( .D(n501), .CP(clk), .CD(n1937), .Q(out1_p2[22]), 
        .QN(n1631) );
  CFD2XL \out1_p2_reg[21]  ( .D(n503), .CP(clk), .CD(n1937), .Q(out1_p2[21]), 
        .QN(n1635) );
  CFD2XL \out1_p2_reg[20]  ( .D(n505), .CP(clk), .CD(n1937), .Q(out1_p2[20]), 
        .QN(n1639) );
  CFD2XL \out1_p2_reg[19]  ( .D(n507), .CP(clk), .CD(n1937), .Q(out1_p2[19]), 
        .QN(n1643) );
  CFD2XL \out1_p2_reg[18]  ( .D(n509), .CP(clk), .CD(n1937), .Q(out1_p2[18]), 
        .QN(n1647) );
  CFD2XL \out1_p2_reg[17]  ( .D(n511), .CP(clk), .CD(n1937), .Q(out1_p2[17]), 
        .QN(n1651) );
  CFD2XL \out2_p2_reg[7]  ( .D(n1142), .CP(clk), .CD(n1937), .Q(out2_p2[7]), 
        .QN(n1445) );
  CFD2XL \out2_p2_reg[33]  ( .D(n1140), .CP(clk), .CD(n1937), .Q(out2_p2[33]), 
        .QN(n1390) );
  CFD2XL \out2_p2_reg[45]  ( .D(n1139), .CP(clk), .CD(n1937), .Q(out2_p2[45]), 
        .QN(n1366) );
  CFD2XL \out2_p2_reg[41]  ( .D(n1141), .CP(clk), .CD(n1937), .Q(out2_p2[41]), 
        .QN(n1374) );
  CFD2XL \out2_p2_reg[37]  ( .D(n1089), .CP(clk), .CD(n1937), .Q(out2_p2[37]), 
        .QN(n1382) );
  CFD2XL \out2_p2_reg[29]  ( .D(n1090), .CP(clk), .CD(n1937), .Q(out2_p2[29]), 
        .QN(n1401) );
  CFD2XL \out2_p2_reg[25]  ( .D(n1092), .CP(clk), .CD(n1937), .Q(out2_p2[25]), 
        .QN(n1409) );
  CFD2XL \out1_p2_reg[15]  ( .D(n515), .CP(clk), .CD(n1937), .Q(out1_p2[15]), 
        .QN(n1659) );
  CFD2XL \out1_p2_reg[13]  ( .D(n519), .CP(clk), .CD(n1937), .Q(out1_p2[13]), 
        .QN(n1667) );
  CFD2XL \out1_p2_reg[11]  ( .D(n523), .CP(clk), .CD(n1937), .Q(out1_p2[11]), 
        .QN(n1675) );
  CFD2XL \out2_p2_reg[1]  ( .D(n1087), .CP(clk), .CD(n1937), .Q(out2_p2[1]), 
        .QN(n1457) );
  CFD2XL \out2_p2_reg[13]  ( .D(n1110), .CP(clk), .CD(n1937), .Q(out2_p2[13]), 
        .QN(n1433) );
  CFD2XL \out2_p2_reg[9]  ( .D(n1109), .CP(clk), .CD(n1937), .Q(out2_p2[9]), 
        .QN(n1441) );
  CFD2XL \out2_p2_reg[5]  ( .D(n1105), .CP(clk), .CD(n1937), .Q(out2_p2[5]), 
        .QN(n1449) );
  CFD2XL \out2_p2_reg[51]  ( .D(n1088), .CP(clk), .CD(n1937), .Q(out2_p2[51]), 
        .QN(n1354) );
  CFD2XL \out2_p2_reg[52]  ( .D(n1091), .CP(clk), .CD(n1937), .Q(out2_p2[52]), 
        .QN(n1352) );
  CFD2XL \out2_p2_reg[48]  ( .D(n1102), .CP(clk), .CD(n1937), .Q(out2_p2[48]), 
        .QN(n1360) );
  CFD2XL \out2_p2_reg[50]  ( .D(n1103), .CP(clk), .CD(n1937), .Q(out2_p2[50]), 
        .QN(n1356) );
  CFD2XL \out2_p2_reg[54]  ( .D(n1101), .CP(clk), .CD(n1937), .Q(out2_p2[54]), 
        .QN(n1348) );
  CFD2XL \out2_p2_reg[19]  ( .D(n1099), .CP(clk), .CD(n1937), .Q(out2_p2[19]), 
        .QN(n1421) );
  CFD2XL \out2_p2_reg[63]  ( .D(n547), .CP(clk), .CD(n1937), .Q(out2_p2[63])
         );
  CFD2XL \out1_p0_reg[13]  ( .D(N27), .CP(clk), .CD(n1937), .Q(out1_p0[13]) );
  CFD2XL \out0_p0_reg[13]  ( .D(N27), .CP(clk), .CD(n1937), .Q(out0_p0[13]) );
  CFD2XL \out2_p2_reg[27]  ( .D(n1100), .CP(clk), .CD(n1937), .Q(out2_p2[27]), 
        .QN(n1405) );
  CFD2XL \out2_p2_reg[32]  ( .D(n1097), .CP(clk), .CD(n1937), .Q(out2_p2[32]), 
        .QN(n1392) );
  CFD2XL \out2_p2_reg[43]  ( .D(n1098), .CP(clk), .CD(n1937), .Q(out2_p2[43]), 
        .QN(n1370) );
  CFD2XL \out2_p2_reg[22]  ( .D(n1095), .CP(clk), .CD(n1937), .Q(out2_p2[22]), 
        .QN(n1415) );
  CFD2XL \out2_p2_reg[20]  ( .D(n1094), .CP(clk), .CD(n1937), .Q(out2_p2[20]), 
        .QN(n1419) );
  CFD2XL \out2_p2_reg[18]  ( .D(n1096), .CP(clk), .CD(n1937), .Q(out2_p2[18]), 
        .QN(n1423) );
  CFD2XL \out2_p2_reg[16]  ( .D(n1093), .CP(clk), .CD(n1937), .Q(out2_p2[16]), 
        .QN(n1427) );
  CFD2XL \out2_p2_reg[35]  ( .D(n1104), .CP(clk), .CD(n1937), .Q(out2_p2[35]), 
        .QN(n1386) );
  CFD2XL \out2_p2_reg[61]  ( .D(n549), .CP(clk), .CD(n1937), .Q(out2_p2[61])
         );
  CFD2XL \out2_p2_reg[60]  ( .D(n550), .CP(clk), .CD(n1937), .Q(out2_p2[60])
         );
  CFD2XL \out2_p2_reg[36]  ( .D(n1155), .CP(clk), .CD(n1937), .Q(out2_p2[36]), 
        .QN(n1384) );
  CFD2XL \out2_p2_reg[46]  ( .D(n1137), .CP(clk), .CD(n1937), .Q(out2_p2[46]), 
        .QN(n1364) );
  CFD2XL \out2_p2_reg[44]  ( .D(n1138), .CP(clk), .CD(n1937), .Q(out2_p2[44]), 
        .QN(n1368) );
  CFD2XL \out2_p2_reg[42]  ( .D(n1129), .CP(clk), .CD(n1937), .Q(out2_p2[42]), 
        .QN(n1372) );
  CFD2XL \out2_p2_reg[40]  ( .D(n1133), .CP(clk), .CD(n1937), .Q(out2_p2[40]), 
        .QN(n1376) );
  CFD2XL \out2_p2_reg[34]  ( .D(n1132), .CP(clk), .CD(n1937), .Q(out2_p2[34]), 
        .QN(n1388) );
  CFD2XL \out2_p2_reg[38]  ( .D(n1134), .CP(clk), .CD(n1937), .Q(out2_p2[38]), 
        .QN(n1380) );
  CFD2XL \out2_p2_reg[11]  ( .D(n1135), .CP(clk), .CD(n1937), .Q(out2_p2[11]), 
        .QN(n1437) );
  CFD2XL \out2_p2_reg[3]  ( .D(n1136), .CP(clk), .CD(n1937), .Q(out2_p2[3]), 
        .QN(n1453) );
  CFD2XL \out2_p2_reg[30]  ( .D(n1119), .CP(clk), .CD(n1937), .Q(out2_p2[30]), 
        .QN(n1399) );
  CFD2XL \out2_p2_reg[28]  ( .D(n1117), .CP(clk), .CD(n1937), .Q(out2_p2[28]), 
        .QN(n1403) );
  CFD2XL \out2_p2_reg[26]  ( .D(n1127), .CP(clk), .CD(n1937), .Q(out2_p2[26]), 
        .QN(n1407) );
  CFD2XL \out2_p2_reg[24]  ( .D(n1121), .CP(clk), .CD(n1937), .Q(out2_p2[24]), 
        .QN(n1411) );
  CFD2XL \out2_p2_reg[4]  ( .D(n1125), .CP(clk), .CD(n1937), .Q(out2_p2[4]), 
        .QN(n1451) );
  CFD2XL \out2_p2_reg[0]  ( .D(n1126), .CP(clk), .CD(n1937), .Q(out2_p2[0]), 
        .QN(n1459) );
  CFD2XL \out2_p2_reg[14]  ( .D(n1124), .CP(clk), .CD(n1937), .Q(out2_p2[14]), 
        .QN(n1431) );
  CFD2XL \out2_p2_reg[12]  ( .D(n1118), .CP(clk), .CD(n1937), .Q(out2_p2[12]), 
        .QN(n1435) );
  CFD2XL \out2_p2_reg[10]  ( .D(n1120), .CP(clk), .CD(n1937), .Q(out2_p2[10]), 
        .QN(n1439) );
  CFD2XL \out2_p2_reg[8]  ( .D(n1123), .CP(clk), .CD(n1937), .Q(out2_p2[8]), 
        .QN(n1443) );
  CFD2XL \out2_p2_reg[2]  ( .D(n1122), .CP(clk), .CD(n1937), .Q(out2_p2[2]), 
        .QN(n1455) );
  CFD2XL \out2_p2_reg[6]  ( .D(n1106), .CP(clk), .CD(n1937), .Q(out2_p2[6]), 
        .QN(n1447) );
  CFD2XL \out2_p2_reg[58]  ( .D(n552), .CP(clk), .CD(n1937), .Q(out2_p2[58])
         );
  CFD2XL \out1_p0_reg[12]  ( .D(N26), .CP(clk), .CD(n1937), .Q(out1_p0[12]) );
  CFD2XL \out0_p0_reg[12]  ( .D(N26), .CP(clk), .CD(n1937), .Q(out0_p0[12]) );
  CFD2XL \out2_p2_reg[59]  ( .D(n551), .CP(clk), .CD(n1937), .Q(out2_p2[59])
         );
  CFD2XL \out2_p2_reg[57]  ( .D(n553), .CP(clk), .CD(n1937), .Q(out2_p2[57])
         );
  CFD2XL \out2_p2_reg[62]  ( .D(n548), .CP(clk), .CD(n1937), .Q(out2_p2[62])
         );
  CFD2XL \out1_p2_reg[48]  ( .D(n449), .CP(clk), .CD(n1937), .Q(out1_p2[48]), 
        .QN(n1527) );
  CFD2XL \out1_p2_reg[47]  ( .D(n451), .CP(clk), .CD(n1937), .Q(out1_p2[47]), 
        .QN(n1531) );
  CFD2XL \out1_p2_reg[46]  ( .D(n453), .CP(clk), .CD(n1937), .Q(out1_p2[46]), 
        .QN(n1535) );
  CFD2XL \out1_p2_reg[45]  ( .D(n455), .CP(clk), .CD(n1937), .Q(out1_p2[45]), 
        .QN(n1539) );
  CFD2XL \out1_p2_reg[44]  ( .D(n457), .CP(clk), .CD(n1937), .Q(out1_p2[44]), 
        .QN(n1543) );
  CFD2XL \out1_p2_reg[43]  ( .D(n459), .CP(clk), .CD(n1937), .Q(out1_p2[43]), 
        .QN(n1547) );
  CFD2XL \out1_p2_reg[42]  ( .D(n461), .CP(clk), .CD(n1937), .Q(out1_p2[42]), 
        .QN(n1551) );
  CFD2XL \out1_p2_reg[41]  ( .D(n463), .CP(clk), .CD(n1937), .Q(out1_p2[41]), 
        .QN(n1555) );
  CFD2XL \out1_p2_reg[40]  ( .D(n465), .CP(clk), .CD(n1937), .Q(out1_p2[40]), 
        .QN(n1559) );
  CFD2XL \out1_p2_reg[39]  ( .D(n467), .CP(clk), .CD(n1937), .Q(out1_p2[39]), 
        .QN(n1563) );
  CFD2XL \out1_p2_reg[38]  ( .D(n469), .CP(clk), .CD(n1937), .Q(out1_p2[38]), 
        .QN(n1567) );
  CFD2XL \out1_p2_reg[37]  ( .D(n471), .CP(clk), .CD(n1937), .Q(out1_p2[37]), 
        .QN(n1571) );
  CFD2XL \out1_p2_reg[36]  ( .D(n473), .CP(clk), .CD(n1937), .Q(out1_p2[36]), 
        .QN(n1575) );
  CFD2XL \out1_p2_reg[35]  ( .D(n475), .CP(clk), .CD(n1937), .Q(out1_p2[35]), 
        .QN(n1579) );
  CFD2XL \out1_p2_reg[34]  ( .D(n477), .CP(clk), .CD(n1937), .Q(out1_p2[34]), 
        .QN(n1583) );
  CFD2XL \out1_p2_reg[33]  ( .D(n479), .CP(clk), .CD(n1937), .Q(out1_p2[33]), 
        .QN(n1587) );
  CFD2XL \out2_p2_reg[56]  ( .D(n554), .CP(clk), .CD(n1937), .Q(out2_p2[56])
         );
  CFD2XL \out1_p2_reg[63]  ( .D(n419), .CP(clk), .CD(n1937), .Q(out1_p2[63]), 
        .QN(n1465) );
  CFD2XL \out1_p2_reg[62]  ( .D(n421), .CP(clk), .CD(n1937), .Q(out1_p2[62]), 
        .QN(n1471) );
  CFD2XL \out1_p2_reg[61]  ( .D(n423), .CP(clk), .CD(n1937), .Q(out1_p2[61]), 
        .QN(n1475) );
  CFD2XL \out1_p2_reg[60]  ( .D(n425), .CP(clk), .CD(n1937), .Q(out1_p2[60]), 
        .QN(n1479) );
  CFD2XL \out1_p2_reg[59]  ( .D(n427), .CP(clk), .CD(n1937), .Q(out1_p2[59]), 
        .QN(n1483) );
  CFD2XL \out1_p2_reg[58]  ( .D(n429), .CP(clk), .CD(n1937), .Q(out1_p2[58]), 
        .QN(n1487) );
  CFD2XL \out1_p2_reg[57]  ( .D(n431), .CP(clk), .CD(n1937), .Q(out1_p2[57]), 
        .QN(n1491) );
  CFD2XL \out1_p2_reg[56]  ( .D(n433), .CP(clk), .CD(n1937), .Q(out1_p2[56]), 
        .QN(n1495) );
  CFD2XL \out1_p2_reg[55]  ( .D(n435), .CP(clk), .CD(n1937), .Q(out1_p2[55]), 
        .QN(n1499) );
  CFD2XL \out1_p2_reg[54]  ( .D(n437), .CP(clk), .CD(n1937), .Q(out1_p2[54]), 
        .QN(n1503) );
  CFD2XL \out1_p2_reg[53]  ( .D(n439), .CP(clk), .CD(n1937), .Q(out1_p2[53]), 
        .QN(n1507) );
  CFD2XL \out1_p2_reg[52]  ( .D(n441), .CP(clk), .CD(n1937), .Q(out1_p2[52]), 
        .QN(n1511) );
  CFD2XL \out1_p2_reg[51]  ( .D(n443), .CP(clk), .CD(n1937), .Q(out1_p2[51]), 
        .QN(n1515) );
  CFD2XL \out1_p2_reg[50]  ( .D(n445), .CP(clk), .CD(n1937), .Q(out1_p2[50]), 
        .QN(n1519) );
  CFD2XL \out1_p2_reg[49]  ( .D(n447), .CP(clk), .CD(n1937), .Q(out1_p2[49]), 
        .QN(n1523) );
  CFD2XL \out1_p0_reg[14]  ( .D(N28), .CP(clk), .CD(n1937), .Q(out1_p0[14]) );
  CFD2XL \out0_p0_reg[14]  ( .D(N28), .CP(clk), .CD(n1937), .Q(out0_p0[14]) );
  CFD2XL \out1_p0_reg[18]  ( .D(N32), .CP(clk), .CD(n1937), .Q(out1_p0[18]) );
  CFD2XL \out0_p0_reg[18]  ( .D(N32), .CP(clk), .CD(n1937), .Q(out0_p0[18]) );
  CFD2XL \out1_p0_reg[21]  ( .D(N35), .CP(clk), .CD(n1937), .Q(out1_p0[21]) );
  CFD2XL \out0_p0_reg[21]  ( .D(N35), .CP(clk), .CD(n1937), .Q(out0_p0[21]) );
  CFD2XL \out1_p0_reg[15]  ( .D(N29), .CP(clk), .CD(n1937), .Q(out1_p0[15]) );
  CFD2XL \out0_p0_reg[15]  ( .D(N29), .CP(clk), .CD(n1937), .Q(out0_p0[15]) );
  CFD2XL \out1_p0_reg[19]  ( .D(N33), .CP(clk), .CD(n1937), .Q(out1_p0[19]) );
  CFD2XL \out0_p0_reg[19]  ( .D(N33), .CP(clk), .CD(n1937), .Q(out0_p0[19]) );
  CFD2XL \out1_p0_reg[28]  ( .D(N42), .CP(clk), .CD(n1937), .Q(out1_p0[28]) );
  CFD2XL \out0_p0_reg[28]  ( .D(N42), .CP(clk), .CD(n1937), .Q(out0_p0[28]) );
  CFD2XL \out1_p0_reg[20]  ( .D(N34), .CP(clk), .CD(n1937), .Q(out1_p0[20]) );
  CFD2XL \out0_p0_reg[20]  ( .D(N34), .CP(clk), .CD(n1937), .Q(out0_p0[20]) );
  CFD2X1 push0_p2_reg ( .D(n1107), .CP(clk), .CD(n1937), .Q(push0_p2), .QN(
        n1936) );
  CFD2QX1 \q0_reg[8]  ( .D(n1114), .CP(clk), .CD(n1284), .Q(q0[8]) );
  CFD2QX1 \q0_reg[5]  ( .D(n663), .CP(clk), .CD(n1285), .Q(q0[5]) );
  CFD2QX1 en1_p2_reg ( .D(n1130), .CP(clk), .CD(n1279), .Q(en1_p2) );
  CFD2QX1 \q0_reg[12]  ( .D(n1115), .CP(clk), .CD(n1284), .Q(q0[12]) );
  CFD2QX1 \h0_reg[6]  ( .D(n632), .CP(clk), .CD(n1287), .Q(h0[6]) );
  CFD2QX1 \q0_reg[24]  ( .D(n682), .CP(clk), .CD(n1283), .Q(q0[24]) );
  CMX2XL U918 ( .A0(q0[16]), .A1(q[16]), .S(n1340), .Z(n674) );
  CNIVX2 U919 ( .A(en2_p2), .Z(n1253) );
  CAN3X2 U920 ( .A(cmd0[1]), .B(n1940), .C(push0), .Z(n787) );
  CAN4X1 U921 ( .A(n1879), .B(push0_p2), .C(n1878), .D(n1877), .Z(n788) );
  CMX2XL U922 ( .A0(q0[31]), .A1(q[31]), .S(n1339), .Z(n689) );
  CMX2XL U923 ( .A0(h0[18]), .A1(h[18]), .S(n1342), .Z(n644) );
  CNIVX1 U924 ( .A(_pushout_d), .Z(n789) );
  CNIVX1 U925 ( .A(n689), .Z(n790) );
  CMX2X2 U926 ( .A0(out0_p2[62]), .A1(out0_p1[62]), .S(n1258), .Z(n691) );
  CMX2X2 U927 ( .A0(out0_p2[61]), .A1(out0_p1[61]), .S(n1259), .Z(n692) );
  CMX2X2 U928 ( .A0(out0_p2[60]), .A1(out0_p1[60]), .S(n1257), .Z(n693) );
  CMX2X2 U929 ( .A0(out0_p2[59]), .A1(out0_p1[59]), .S(n1256), .Z(n694) );
  CMX2X2 U930 ( .A0(out0_p2[58]), .A1(out0_p1[58]), .S(n1257), .Z(n695) );
  CMX2X2 U931 ( .A0(out0_p2[57]), .A1(out0_p1[57]), .S(n1258), .Z(n696) );
  CMX2X2 U932 ( .A0(out0_p2[56]), .A1(out0_p1[56]), .S(n1258), .Z(n697) );
  CMX2X2 U933 ( .A0(out0_p2[55]), .A1(out0_p1[55]), .S(n1259), .Z(n698) );
  CMX2X2 U934 ( .A0(out0_p2[54]), .A1(out0_p1[54]), .S(n1256), .Z(n699) );
  CMX2X2 U935 ( .A0(out0_p2[53]), .A1(out0_p1[53]), .S(n1257), .Z(n700) );
  CMX2X2 U936 ( .A0(out0_p2[52]), .A1(out0_p1[52]), .S(n1259), .Z(n701) );
  CMX2X2 U937 ( .A0(out0_p2[51]), .A1(out0_p1[51]), .S(n1258), .Z(n702) );
  CMX2X2 U938 ( .A0(out0_p2[50]), .A1(out0_p1[50]), .S(n1259), .Z(n703) );
  CMX2X2 U939 ( .A0(out0_p2[49]), .A1(out0_p1[49]), .S(n1256), .Z(n704) );
  CMX2X2 U940 ( .A0(out0_p2[48]), .A1(out0_p1[48]), .S(n1256), .Z(n705) );
  CMX2X2 U941 ( .A0(out0_p2[47]), .A1(out0_p1[47]), .S(n1257), .Z(n706) );
  CMX2X2 U942 ( .A0(out0_p2[46]), .A1(out0_p1[46]), .S(n1258), .Z(n707) );
  CMX2X2 U943 ( .A0(out0_p2[45]), .A1(out0_p1[45]), .S(n1259), .Z(n708) );
  CMX2X2 U944 ( .A0(out0_p2[44]), .A1(out0_p1[44]), .S(n1257), .Z(n709) );
  CMX2X2 U945 ( .A0(out0_p2[43]), .A1(out0_p1[43]), .S(n1256), .Z(n710) );
  CMX2X2 U946 ( .A0(out0_p2[42]), .A1(out0_p1[42]), .S(n1257), .Z(n711) );
  CMX2X2 U947 ( .A0(out0_p2[41]), .A1(out0_p1[41]), .S(n1258), .Z(n712) );
  CMX2X2 U948 ( .A0(out0_p2[40]), .A1(out0_p1[40]), .S(n1258), .Z(n713) );
  CMX2X2 U949 ( .A0(out0_p2[39]), .A1(out0_p1[39]), .S(n1259), .Z(n714) );
  CMX2X2 U950 ( .A0(out0_p2[38]), .A1(out0_p1[38]), .S(n1256), .Z(n715) );
  CMX2X2 U951 ( .A0(out0_p2[37]), .A1(out0_p1[37]), .S(n1257), .Z(n716) );
  CMX2X2 U952 ( .A0(out0_p2[36]), .A1(out0_p1[36]), .S(n1259), .Z(n717) );
  CMX2X2 U953 ( .A0(out0_p2[35]), .A1(out0_p1[35]), .S(n1258), .Z(n718) );
  CMX2X2 U954 ( .A0(out0_p2[34]), .A1(out0_p1[34]), .S(n1259), .Z(n719) );
  CMX2X2 U955 ( .A0(out0_p2[33]), .A1(out0_p1[33]), .S(n1256), .Z(n720) );
  CMX2X2 U956 ( .A0(out0_p2[32]), .A1(out0_p1[32]), .S(n1256), .Z(n721) );
  CMX2X2 U957 ( .A0(out0_p2[31]), .A1(out0_p1[31]), .S(n1257), .Z(n722) );
  CMX2X2 U958 ( .A0(out0_p2[30]), .A1(out0_p1[30]), .S(n1258), .Z(n723) );
  CMX2X2 U959 ( .A0(out0_p2[29]), .A1(out0_p1[29]), .S(n1259), .Z(n724) );
  CMX2X2 U960 ( .A0(out0_p2[28]), .A1(out0_p1[28]), .S(n1257), .Z(n725) );
  CMX2X2 U961 ( .A0(out0_p2[27]), .A1(out0_p1[27]), .S(n1256), .Z(n726) );
  CMX2X2 U962 ( .A0(out0_p2[26]), .A1(out0_p1[26]), .S(n1257), .Z(n727) );
  CMX2X2 U963 ( .A0(out0_p2[25]), .A1(out0_p1[25]), .S(n1258), .Z(n728) );
  CMX2X2 U964 ( .A0(out0_p2[24]), .A1(out0_p1[24]), .S(n1258), .Z(n729) );
  CMX2X2 U965 ( .A0(out0_p2[23]), .A1(out0_p1[23]), .S(n1259), .Z(n730) );
  CMX2X2 U966 ( .A0(out0_p2[22]), .A1(out0_p1[22]), .S(n1256), .Z(n731) );
  CMX2X2 U967 ( .A0(out0_p2[21]), .A1(out0_p1[21]), .S(n1257), .Z(n732) );
  CMX2X2 U968 ( .A0(out0_p2[20]), .A1(out0_p1[20]), .S(n1259), .Z(n733) );
  CMX2X2 U969 ( .A0(out0_p2[19]), .A1(out0_p1[19]), .S(n1258), .Z(n734) );
  CMX2X2 U970 ( .A0(out0_p2[18]), .A1(out0_p1[18]), .S(n1259), .Z(n735) );
  CMX2X2 U971 ( .A0(out0_p2[17]), .A1(out0_p1[17]), .S(n1256), .Z(n736) );
  CMX2X2 U972 ( .A0(out0_p2[16]), .A1(out0_p1[16]), .S(n1256), .Z(n737) );
  CMX2X2 U973 ( .A0(out0_p2[15]), .A1(out0_p1[15]), .S(n1257), .Z(n738) );
  CMX2X2 U974 ( .A0(out0_p2[14]), .A1(out0_p1[14]), .S(n1258), .Z(n739) );
  CMX2X2 U975 ( .A0(out0_p2[13]), .A1(out0_p1[13]), .S(n1259), .Z(n740) );
  CMX2X2 U976 ( .A0(out0_p2[12]), .A1(out0_p1[12]), .S(n1257), .Z(n741) );
  CMX2X2 U977 ( .A0(out0_p2[11]), .A1(out0_p1[11]), .S(n1256), .Z(n742) );
  CMX2X2 U978 ( .A0(out0_p2[10]), .A1(out0_p1[10]), .S(n1257), .Z(n743) );
  CMX2X2 U979 ( .A0(out0_p2[9]), .A1(out0_p1[9]), .S(n1258), .Z(n744) );
  CMX2X2 U980 ( .A0(out0_p2[8]), .A1(out0_p1[8]), .S(n1258), .Z(n745) );
  CMX2X2 U981 ( .A0(out0_p2[7]), .A1(out0_p1[7]), .S(n1259), .Z(n746) );
  CMX2X2 U982 ( .A0(out0_p2[6]), .A1(out0_p1[6]), .S(n1256), .Z(n747) );
  CMX2X2 U983 ( .A0(out0_p2[5]), .A1(out0_p1[5]), .S(n1257), .Z(n748) );
  CMX2X2 U984 ( .A0(out0_p2[4]), .A1(out0_p1[4]), .S(n1259), .Z(n749) );
  CMX2X2 U985 ( .A0(out0_p2[3]), .A1(out0_p1[3]), .S(n1258), .Z(n750) );
  CMX2X2 U986 ( .A0(out0_p2[2]), .A1(out0_p1[2]), .S(n1259), .Z(n751) );
  CMX2X2 U987 ( .A0(out0_p2[1]), .A1(out0_p1[1]), .S(n1256), .Z(n752) );
  CMX2X2 U988 ( .A0(out0_p2[0]), .A1(out0_p1[0]), .S(n1256), .Z(n753) );
  CIVDX1 U989 ( .A(out1_p0[0]), .Z1(n792) );
  CNIVX1 U990 ( .A(n792), .Z(n791) );
  CIVDX1 U991 ( .A(out1_p0[1]), .Z1(n794) );
  CNIVX1 U992 ( .A(n794), .Z(n793) );
  CIVDX1 U993 ( .A(out1_p0[2]), .Z1(n796) );
  CNIVX1 U994 ( .A(n796), .Z(n795) );
  CIVDX1 U995 ( .A(out1_p0[3]), .Z1(n798) );
  CNIVX1 U996 ( .A(n798), .Z(n797) );
  CIVDX1 U997 ( .A(out1_p0[4]), .Z1(n800) );
  CNIVX1 U998 ( .A(n800), .Z(n799) );
  CIVDX1 U999 ( .A(out1_p0[5]), .Z1(n802) );
  CNIVX1 U1000 ( .A(n802), .Z(n801) );
  CIVDX1 U1001 ( .A(out1_p0[6]), .Z1(n804) );
  CNIVX1 U1002 ( .A(n804), .Z(n803) );
  CIVDX1 U1003 ( .A(out1_p0[7]), .Z1(n806) );
  CNIVX1 U1004 ( .A(n806), .Z(n805) );
  CIVDX1 U1005 ( .A(out1_p0[8]), .Z1(n808) );
  CNIVX1 U1006 ( .A(n808), .Z(n807) );
  CIVDX1 U1007 ( .A(out1_p0[9]), .Z1(n810) );
  CNIVX1 U1008 ( .A(n810), .Z(n809) );
  CIVDX1 U1009 ( .A(out1_p0[10]), .Z1(n812) );
  CNIVX1 U1010 ( .A(n812), .Z(n811) );
  CIVDX1 U1011 ( .A(out1_p0[11]), .Z1(n814) );
  CNIVX1 U1012 ( .A(n814), .Z(n813) );
  CIVDX1 U1013 ( .A(out1_p0[12]), .Z1(n816) );
  CNIVX1 U1014 ( .A(n816), .Z(n815) );
  CIVDX1 U1015 ( .A(out1_p0[13]), .Z1(n818) );
  CNIVX1 U1016 ( .A(n818), .Z(n817) );
  CIVDX1 U1017 ( .A(out1_p0[14]), .Z1(n820) );
  CNIVX1 U1018 ( .A(n820), .Z(n819) );
  CIVDX1 U1019 ( .A(out1_p0[15]), .Z1(n822) );
  CNIVX1 U1020 ( .A(n822), .Z(n821) );
  CIVDX1 U1021 ( .A(out1_p0[16]), .Z1(n824) );
  CNIVX1 U1022 ( .A(n824), .Z(n823) );
  CIVDX1 U1023 ( .A(out1_p0[17]), .Z1(n826) );
  CNIVX1 U1024 ( .A(n826), .Z(n825) );
  CIVDX1 U1025 ( .A(out1_p0[18]), .Z1(n828) );
  CNIVX1 U1026 ( .A(n828), .Z(n827) );
  CIVDX1 U1027 ( .A(out1_p0[19]), .Z1(n830) );
  CNIVX1 U1028 ( .A(n830), .Z(n829) );
  CIVDX1 U1029 ( .A(out1_p0[20]), .Z1(n832) );
  CNIVX1 U1030 ( .A(n832), .Z(n831) );
  CIVDX1 U1031 ( .A(out1_p0[21]), .Z1(n834) );
  CNIVX1 U1032 ( .A(n834), .Z(n833) );
  CIVDX1 U1033 ( .A(out1_p0[22]), .Z1(n836) );
  CNIVX1 U1034 ( .A(n836), .Z(n835) );
  CIVDX1 U1035 ( .A(out1_p0[23]), .Z1(n838) );
  CNIVX1 U1036 ( .A(n838), .Z(n837) );
  CIVDX1 U1037 ( .A(out1_p0[24]), .Z1(n840) );
  CNIVX1 U1038 ( .A(n840), .Z(n839) );
  CIVDX1 U1039 ( .A(out1_p0[25]), .Z1(n842) );
  CNIVX1 U1040 ( .A(n842), .Z(n841) );
  CIVDX1 U1041 ( .A(out1_p0[26]), .Z1(n844) );
  CNIVX1 U1042 ( .A(n844), .Z(n843) );
  CIVDX1 U1043 ( .A(out1_p0[27]), .Z1(n846) );
  CNIVX1 U1044 ( .A(n846), .Z(n845) );
  CIVDX1 U1045 ( .A(out1_p0[28]), .Z1(n848) );
  CNIVX1 U1046 ( .A(n848), .Z(n847) );
  CIVDX1 U1047 ( .A(out1_p0[29]), .Z1(n850) );
  CNIVX1 U1048 ( .A(n850), .Z(n849) );
  CIVDX1 U1049 ( .A(out1_p0[30]), .Z1(n852) );
  CNIVX1 U1050 ( .A(n852), .Z(n851) );
  CIVDX1 U1051 ( .A(out1_p0[31]), .Z1(n854) );
  CNIVX1 U1052 ( .A(n854), .Z(n853) );
  CIVDX1 U1053 ( .A(out1_p0[32]), .Z1(n856) );
  CNIVX1 U1054 ( .A(n856), .Z(n855) );
  CIVDX1 U1055 ( .A(out1_p0[33]), .Z1(n858) );
  CNIVX1 U1056 ( .A(n858), .Z(n857) );
  CIVDX1 U1057 ( .A(out1_p0[34]), .Z1(n860) );
  CNIVX1 U1058 ( .A(n860), .Z(n859) );
  CIVDX1 U1059 ( .A(out1_p0[35]), .Z1(n862) );
  CNIVX1 U1060 ( .A(n862), .Z(n861) );
  CIVDX1 U1061 ( .A(out1_p0[36]), .Z1(n864) );
  CNIVX1 U1062 ( .A(n864), .Z(n863) );
  CIVDX1 U1063 ( .A(out1_p0[37]), .Z1(n866) );
  CNIVX1 U1064 ( .A(n866), .Z(n865) );
  CIVDX1 U1065 ( .A(out1_p0[38]), .Z1(n868) );
  CNIVX1 U1066 ( .A(n868), .Z(n867) );
  CIVDX1 U1067 ( .A(out1_p0[39]), .Z1(n870) );
  CNIVX1 U1068 ( .A(n870), .Z(n869) );
  CIVDX1 U1069 ( .A(out1_p0[40]), .Z1(n872) );
  CNIVX1 U1070 ( .A(n872), .Z(n871) );
  CIVDX1 U1071 ( .A(out1_p0[42]), .Z1(n874) );
  CNIVX1 U1072 ( .A(n874), .Z(n873) );
  CIVDX1 U1073 ( .A(out1_p0[43]), .Z1(n876) );
  CNIVX1 U1074 ( .A(n876), .Z(n875) );
  CIVDX1 U1075 ( .A(out1_p0[44]), .Z1(n878) );
  CNIVX1 U1076 ( .A(n878), .Z(n877) );
  CIVDX1 U1077 ( .A(out1_p0[45]), .Z1(n880) );
  CNIVX1 U1078 ( .A(n880), .Z(n879) );
  CIVDX1 U1079 ( .A(out1_p0[46]), .Z1(n882) );
  CNIVX1 U1080 ( .A(n882), .Z(n881) );
  CIVDX1 U1081 ( .A(out1_p0[47]), .Z1(n884) );
  CNIVX1 U1082 ( .A(n884), .Z(n883) );
  CIVDX1 U1083 ( .A(out1_p0[48]), .Z1(n886) );
  CNIVX1 U1084 ( .A(n886), .Z(n885) );
  CIVDX1 U1085 ( .A(out1_p0[49]), .Z1(n888) );
  CNIVX1 U1086 ( .A(n888), .Z(n887) );
  CIVDX1 U1087 ( .A(out1_p0[50]), .Z1(n890) );
  CNIVX1 U1088 ( .A(n890), .Z(n889) );
  CIVDX1 U1089 ( .A(out1_p0[51]), .Z1(n892) );
  CNIVX1 U1090 ( .A(n892), .Z(n891) );
  CIVDX1 U1091 ( .A(out1_p0[52]), .Z1(n894) );
  CNIVX1 U1092 ( .A(n894), .Z(n893) );
  CIVDX1 U1093 ( .A(out1_p0[53]), .Z1(n896) );
  CNIVX1 U1094 ( .A(n896), .Z(n895) );
  CIVDX1 U1095 ( .A(out1_p0[55]), .Z1(n898) );
  CNIVX1 U1096 ( .A(n898), .Z(n897) );
  CIVDX1 U1097 ( .A(out1_p0[56]), .Z1(n900) );
  CNIVX1 U1098 ( .A(n900), .Z(n899) );
  CIVDX1 U1099 ( .A(out1_p0[57]), .Z1(n902) );
  CNIVX1 U1100 ( .A(n902), .Z(n901) );
  CIVDX1 U1101 ( .A(out1_p0[58]), .Z1(n904) );
  CNIVX1 U1102 ( .A(n904), .Z(n903) );
  CIVDX1 U1103 ( .A(out1_p0[59]), .Z1(n906) );
  CNIVX1 U1104 ( .A(n906), .Z(n905) );
  CIVDX1 U1105 ( .A(en0_p1), .Z1(n908) );
  CNIVX1 U1106 ( .A(n908), .Z(n907) );
  CIVDX1 U1107 ( .A(cmd0_p1[1]), .Z1(n910) );
  CNIVX1 U1108 ( .A(n910), .Z(n909) );
  CIVDX1 U1109 ( .A(cmd0_p1[0]), .Z1(n912) );
  CNIVX1 U1110 ( .A(n912), .Z(n911) );
  CMX2X2 U1111 ( .A0(out0_p2[63]), .A1(out0_p1[63]), .S(n1257), .Z(n690) );
  CIVDX1 U1112 ( .A(out1_p0[54]), .Z1(n914) );
  CNIVX1 U1113 ( .A(n914), .Z(n913) );
  CIVDX1 U1114 ( .A(out1_p0[60]), .Z1(n916) );
  CNIVX1 U1115 ( .A(n916), .Z(n915) );
  CIVDX1 U1116 ( .A(out1_p0[61]), .Z1(n918) );
  CNIVX1 U1117 ( .A(n918), .Z(n917) );
  CIVDX1 U1118 ( .A(out1_p0[62]), .Z1(n920) );
  CNIVX1 U1119 ( .A(n920), .Z(n919) );
  CIVDX1 U1120 ( .A(out1_p0[63]), .Z1(n922) );
  CNIVX1 U1121 ( .A(n922), .Z(n921) );
  CNIVX1 U1122 ( .A(n613), .Z(n923) );
  CNIVX1 U1123 ( .A(n616), .Z(n924) );
  CNIVX1 U1124 ( .A(h0[1]), .Z(n925) );
  CNIVX1 U1125 ( .A(n619), .Z(n926) );
  CNIVX1 U1126 ( .A(h0[2]), .Z(n927) );
  CNIVX1 U1127 ( .A(n622), .Z(n928) );
  CNIVX1 U1128 ( .A(n625), .Z(n929) );
  CNIVX1 U1129 ( .A(n628), .Z(n930) );
  CNIVX1 U1130 ( .A(h0[5]), .Z(n931) );
  CNIVX1 U1131 ( .A(n631), .Z(n932) );
  CNIVX1 U1132 ( .A(h0[6]), .Z(n933) );
  CMXI2X2 U1133 ( .A0(n1881), .A1(n1880), .S(n788), .Z(n755) );
  CMX2X2 U1134 ( .A0(z[1]), .A1(acc[1]), .S(n788), .Z(n756) );
  CMXI2X2 U1135 ( .A0(n1883), .A1(n1882), .S(n788), .Z(n757) );
  CMX2X2 U1136 ( .A0(z[3]), .A1(acc[3]), .S(n788), .Z(n758) );
  CMXI2X2 U1137 ( .A0(n1885), .A1(n1884), .S(n788), .Z(n759) );
  CMXI2X2 U1138 ( .A0(n1887), .A1(n1886), .S(n788), .Z(n760) );
  CMXI2X2 U1139 ( .A0(n1889), .A1(n1888), .S(n788), .Z(n761) );
  CMXI2X2 U1140 ( .A0(n1891), .A1(n1890), .S(n788), .Z(n762) );
  CMXI2X2 U1141 ( .A0(n1893), .A1(n1892), .S(n788), .Z(n763) );
  CMX2X2 U1142 ( .A0(z[9]), .A1(acc[9]), .S(n788), .Z(n764) );
  CMXI2X2 U1143 ( .A0(n1895), .A1(n1894), .S(n788), .Z(n765) );
  CMX2X2 U1144 ( .A0(z[11]), .A1(acc[11]), .S(n788), .Z(n766) );
  CMXI2X2 U1145 ( .A0(n1897), .A1(n1896), .S(n788), .Z(n767) );
  CMXI2X2 U1146 ( .A0(n1899), .A1(n1898), .S(n788), .Z(n768) );
  CMXI2X2 U1147 ( .A0(n1901), .A1(n1900), .S(n788), .Z(n769) );
  CMXI2X2 U1148 ( .A0(n1903), .A1(n1902), .S(n788), .Z(n770) );
  CMXI2X2 U1149 ( .A0(n1905), .A1(n1904), .S(n788), .Z(n771) );
  CMXI2X2 U1150 ( .A0(n1907), .A1(n1906), .S(n788), .Z(n772) );
  CMXI2X2 U1151 ( .A0(n1909), .A1(n1908), .S(n788), .Z(n773) );
  CMXI2X2 U1152 ( .A0(n1911), .A1(n1910), .S(n788), .Z(n774) );
  CMXI2X2 U1153 ( .A0(n1913), .A1(n1912), .S(n788), .Z(n775) );
  CMXI2X2 U1154 ( .A0(n1915), .A1(n1914), .S(n788), .Z(n776) );
  CMXI2X2 U1155 ( .A0(n1917), .A1(n1916), .S(n788), .Z(n777) );
  CMXI2X2 U1156 ( .A0(n1919), .A1(n1918), .S(n788), .Z(n778) );
  CMXI2X2 U1157 ( .A0(n1921), .A1(n1920), .S(n788), .Z(n779) );
  CMXI2X2 U1158 ( .A0(n1923), .A1(n1922), .S(n788), .Z(n780) );
  CMXI2X2 U1159 ( .A0(n1925), .A1(n1924), .S(n788), .Z(n781) );
  CMXI2X2 U1160 ( .A0(n1927), .A1(n1926), .S(n788), .Z(n782) );
  CMXI2X2 U1161 ( .A0(n1929), .A1(n1928), .S(n788), .Z(n783) );
  CMXI2X2 U1162 ( .A0(n1931), .A1(n1930), .S(n788), .Z(n784) );
  CMXI2X2 U1163 ( .A0(n1933), .A1(n1932), .S(n788), .Z(n785) );
  CMXI2X2 U1164 ( .A0(n1935), .A1(n1934), .S(n788), .Z(n786) );
  CIVDX1 U1165 ( .A(out0_p0[0]), .Z1(n935) );
  CNIVX1 U1166 ( .A(n935), .Z(n934) );
  CIVDX1 U1167 ( .A(out0_p0[1]), .Z1(n937) );
  CNIVX1 U1168 ( .A(n937), .Z(n936) );
  CIVDX1 U1169 ( .A(out0_p0[2]), .Z1(n939) );
  CNIVX1 U1170 ( .A(n939), .Z(n938) );
  CIVDX1 U1171 ( .A(out0_p0[3]), .Z1(n941) );
  CNIVX1 U1172 ( .A(n941), .Z(n940) );
  CIVDX1 U1173 ( .A(out0_p0[4]), .Z1(n943) );
  CNIVX1 U1174 ( .A(n943), .Z(n942) );
  CIVDX1 U1175 ( .A(out0_p0[5]), .Z1(n945) );
  CNIVX1 U1176 ( .A(n945), .Z(n944) );
  CIVDX1 U1177 ( .A(out0_p0[6]), .Z1(n947) );
  CNIVX1 U1178 ( .A(n947), .Z(n946) );
  CIVDX1 U1179 ( .A(out0_p0[7]), .Z1(n949) );
  CNIVX1 U1180 ( .A(n949), .Z(n948) );
  CIVDX1 U1181 ( .A(out0_p0[8]), .Z1(n951) );
  CNIVX1 U1182 ( .A(n951), .Z(n950) );
  CIVDX1 U1183 ( .A(out0_p0[9]), .Z1(n953) );
  CNIVX1 U1184 ( .A(n953), .Z(n952) );
  CIVDX1 U1185 ( .A(out0_p0[10]), .Z1(n955) );
  CNIVX1 U1186 ( .A(n955), .Z(n954) );
  CIVDX1 U1187 ( .A(out0_p0[11]), .Z1(n957) );
  CNIVX1 U1188 ( .A(n957), .Z(n956) );
  CIVDX1 U1189 ( .A(out0_p0[12]), .Z1(n959) );
  CNIVX1 U1190 ( .A(n959), .Z(n958) );
  CIVDX1 U1191 ( .A(out0_p0[13]), .Z1(n961) );
  CNIVX1 U1192 ( .A(n961), .Z(n960) );
  CIVDX1 U1193 ( .A(out0_p0[14]), .Z1(n963) );
  CNIVX1 U1194 ( .A(n963), .Z(n962) );
  CIVDX1 U1195 ( .A(out0_p0[15]), .Z1(n965) );
  CNIVX1 U1196 ( .A(n965), .Z(n964) );
  CIVDX1 U1197 ( .A(out0_p0[16]), .Z1(n967) );
  CNIVX1 U1198 ( .A(n967), .Z(n966) );
  CIVDX1 U1199 ( .A(out0_p0[17]), .Z1(n969) );
  CNIVX1 U1200 ( .A(n969), .Z(n968) );
  CIVDX1 U1201 ( .A(out0_p0[18]), .Z1(n971) );
  CNIVX1 U1202 ( .A(n971), .Z(n970) );
  CIVDX1 U1203 ( .A(out0_p0[19]), .Z1(n973) );
  CNIVX1 U1204 ( .A(n973), .Z(n972) );
  CIVDX1 U1205 ( .A(out0_p0[20]), .Z1(n975) );
  CNIVX1 U1206 ( .A(n975), .Z(n974) );
  CIVDX1 U1207 ( .A(out0_p0[21]), .Z1(n977) );
  CNIVX1 U1208 ( .A(n977), .Z(n976) );
  CIVDX1 U1209 ( .A(out0_p0[22]), .Z1(n979) );
  CNIVX1 U1210 ( .A(n979), .Z(n978) );
  CIVDX1 U1211 ( .A(out0_p0[23]), .Z1(n981) );
  CNIVX1 U1212 ( .A(n981), .Z(n980) );
  CIVDX1 U1213 ( .A(out0_p0[24]), .Z1(n983) );
  CNIVX1 U1214 ( .A(n983), .Z(n982) );
  CIVDX1 U1215 ( .A(out0_p0[25]), .Z1(n985) );
  CNIVX1 U1216 ( .A(n985), .Z(n984) );
  CIVDX1 U1217 ( .A(out0_p0[26]), .Z1(n987) );
  CNIVX1 U1218 ( .A(n987), .Z(n986) );
  CIVDX1 U1219 ( .A(out0_p0[27]), .Z1(n989) );
  CNIVX1 U1220 ( .A(n989), .Z(n988) );
  CIVDX1 U1221 ( .A(out0_p0[28]), .Z1(n991) );
  CNIVX1 U1222 ( .A(n991), .Z(n990) );
  CIVDX1 U1223 ( .A(out0_p0[29]), .Z1(n993) );
  CNIVX1 U1224 ( .A(n993), .Z(n992) );
  CIVDX1 U1225 ( .A(out0_p0[30]), .Z1(n995) );
  CNIVX1 U1226 ( .A(n995), .Z(n994) );
  CIVDX1 U1227 ( .A(out0_p0[31]), .Z1(n997) );
  CNIVX1 U1228 ( .A(n997), .Z(n996) );
  CIVDX1 U1229 ( .A(out0_p0[32]), .Z1(n999) );
  CNIVX1 U1230 ( .A(n999), .Z(n998) );
  CIVDX1 U1231 ( .A(out0_p0[33]), .Z1(n1001) );
  CNIVX1 U1232 ( .A(n1001), .Z(n1000) );
  CIVDX1 U1233 ( .A(out0_p0[34]), .Z1(n1003) );
  CNIVX1 U1234 ( .A(n1003), .Z(n1002) );
  CIVDX1 U1235 ( .A(out0_p0[35]), .Z1(n1005) );
  CNIVX1 U1236 ( .A(n1005), .Z(n1004) );
  CIVDX1 U1237 ( .A(out0_p0[36]), .Z1(n1007) );
  CNIVX1 U1238 ( .A(n1007), .Z(n1006) );
  CIVDX1 U1239 ( .A(out0_p0[37]), .Z1(n1009) );
  CNIVX1 U1240 ( .A(n1009), .Z(n1008) );
  CIVDX1 U1241 ( .A(out0_p0[38]), .Z1(n1011) );
  CNIVX1 U1242 ( .A(n1011), .Z(n1010) );
  CIVDX1 U1243 ( .A(out0_p0[39]), .Z1(n1013) );
  CNIVX1 U1244 ( .A(n1013), .Z(n1012) );
  CIVDX1 U1245 ( .A(out0_p0[40]), .Z1(n1015) );
  CNIVX1 U1246 ( .A(n1015), .Z(n1014) );
  CIVDX1 U1247 ( .A(out0_p0[41]), .Z1(n1017) );
  CNIVX1 U1248 ( .A(n1017), .Z(n1016) );
  CIVDX1 U1249 ( .A(out0_p0[42]), .Z1(n1019) );
  CNIVX1 U1250 ( .A(n1019), .Z(n1018) );
  CIVDX1 U1251 ( .A(out0_p0[43]), .Z1(n1021) );
  CNIVX1 U1252 ( .A(n1021), .Z(n1020) );
  CIVDX1 U1253 ( .A(out0_p0[44]), .Z1(n1023) );
  CNIVX1 U1254 ( .A(n1023), .Z(n1022) );
  CIVDX1 U1255 ( .A(out0_p0[45]), .Z1(n1025) );
  CNIVX1 U1256 ( .A(n1025), .Z(n1024) );
  CIVDX1 U1257 ( .A(out0_p0[46]), .Z1(n1027) );
  CNIVX1 U1258 ( .A(n1027), .Z(n1026) );
  CIVDX1 U1259 ( .A(out0_p0[47]), .Z1(n1029) );
  CNIVX1 U1260 ( .A(n1029), .Z(n1028) );
  CIVDX1 U1261 ( .A(out0_p0[48]), .Z1(n1031) );
  CNIVX1 U1262 ( .A(n1031), .Z(n1030) );
  CIVDX1 U1263 ( .A(out0_p0[49]), .Z1(n1033) );
  CNIVX1 U1264 ( .A(n1033), .Z(n1032) );
  CIVDX1 U1265 ( .A(out0_p0[50]), .Z1(n1035) );
  CNIVX1 U1266 ( .A(n1035), .Z(n1034) );
  CIVDX1 U1267 ( .A(out0_p0[51]), .Z1(n1037) );
  CNIVX1 U1268 ( .A(n1037), .Z(n1036) );
  CIVDX1 U1269 ( .A(out0_p0[52]), .Z1(n1039) );
  CNIVX1 U1270 ( .A(n1039), .Z(n1038) );
  CIVDX1 U1271 ( .A(out0_p0[53]), .Z1(n1041) );
  CNIVX1 U1272 ( .A(n1041), .Z(n1040) );
  CIVDX1 U1273 ( .A(out0_p0[54]), .Z1(n1043) );
  CNIVX1 U1274 ( .A(n1043), .Z(n1042) );
  CIVDX1 U1275 ( .A(out0_p0[55]), .Z1(n1045) );
  CNIVX1 U1276 ( .A(n1045), .Z(n1044) );
  CIVDX1 U1277 ( .A(out0_p0[56]), .Z1(n1047) );
  CNIVX1 U1278 ( .A(n1047), .Z(n1046) );
  CIVDX1 U1279 ( .A(out0_p0[57]), .Z1(n1049) );
  CNIVX1 U1280 ( .A(n1049), .Z(n1048) );
  CIVDX1 U1281 ( .A(out0_p0[58]), .Z1(n1051) );
  CNIVX1 U1282 ( .A(n1051), .Z(n1050) );
  CIVDX1 U1283 ( .A(out0_p0[59]), .Z1(n1053) );
  CNIVX1 U1284 ( .A(n1053), .Z(n1052) );
  CIVDX1 U1285 ( .A(out0_p0[60]), .Z1(n1055) );
  CNIVX1 U1286 ( .A(n1055), .Z(n1054) );
  CIVDX1 U1287 ( .A(out0_p0[61]), .Z1(n1057) );
  CNIVX1 U1288 ( .A(n1057), .Z(n1056) );
  CIVDX1 U1289 ( .A(out0_p0[62]), .Z1(n1059) );
  CNIVX1 U1290 ( .A(n1059), .Z(n1058) );
  CIVDX1 U1291 ( .A(out0_p0[63]), .Z1(n1061) );
  CNIVX1 U1292 ( .A(n1061), .Z(n1060) );
  CNIVX1 U1293 ( .A(n652), .Z(n1062) );
  CIVDX1 U1294 ( .A(cmd0[1]), .Z1(n1063) );
  CIVDX1 U1295 ( .A(cmd0_p0[1]), .Z1(n1065) );
  CNIVX1 U1296 ( .A(n1065), .Z(n1064) );
  CIVDX1 U1297 ( .A(cmd0[0]), .Z1(n1066) );
  CIVDX1 U1298 ( .A(cmd0_p0[0]), .Z1(n1068) );
  CNIVX1 U1299 ( .A(n1068), .Z(n1067) );
  CNIVX1 U1300 ( .A(n1070), .Z(n1069) );
  CNIVX1 U1301 ( .A(push0), .Z(n1070) );
  CIVDX1 U1302 ( .A(push0_p0), .Z1(n1072) );
  CNIVX1 U1303 ( .A(n1072), .Z(n1071) );
  CNIVX1 U1304 ( .A(h0[4]), .Z(n1073) );
  CNIVX1 U1305 ( .A(n638), .Z(n1074) );
  CIVDX1 U1306 ( .A(out1_p0[41]), .Z1(n1076) );
  CNIVX1 U1307 ( .A(n1076), .Z(n1075) );
  CNIVX1 U1308 ( .A(n639), .Z(n1077) );
  CNIVX1 U1309 ( .A(n680), .Z(n1078) );
  CNIVX1 U1310 ( .A(n650), .Z(n1079) );
  CNIVX1 U1311 ( .A(n641), .Z(n1080) );
  CNIVX1 U1312 ( .A(n636), .Z(n1081) );
  CNIVX1 U1313 ( .A(n637), .Z(n1082) );
  CNIVX1 U1314 ( .A(n647), .Z(n1083) );
  CNIVX1 U1315 ( .A(n634), .Z(n1084) );
  CNIVX1 U1316 ( .A(n642), .Z(n1085) );
  CNIVX1 U1317 ( .A(n640), .Z(n1086) );
  CNIVX1 U1318 ( .A(n609), .Z(n1087) );
  CNIVX1 U1319 ( .A(n559), .Z(n1088) );
  CNIVX1 U1320 ( .A(n573), .Z(n1089) );
  CNIVX1 U1321 ( .A(n581), .Z(n1090) );
  CNIVX1 U1322 ( .A(n558), .Z(n1091) );
  CNIVX1 U1323 ( .A(n585), .Z(n1092) );
  CNIVX1 U1324 ( .A(n594), .Z(n1093) );
  CNIVX1 U1325 ( .A(n590), .Z(n1094) );
  CNIVX1 U1326 ( .A(n588), .Z(n1095) );
  CNIVX1 U1327 ( .A(n592), .Z(n1096) );
  CNIVX1 U1328 ( .A(n578), .Z(n1097) );
  CNIVX1 U1329 ( .A(n567), .Z(n1098) );
  CNIVX1 U1330 ( .A(n591), .Z(n1099) );
  CNIVX1 U1331 ( .A(n583), .Z(n1100) );
  CNIVX1 U1332 ( .A(n556), .Z(n1101) );
  CNIVX1 U1333 ( .A(n562), .Z(n1102) );
  CNIVX1 U1334 ( .A(n560), .Z(n1103) );
  CNIVX1 U1335 ( .A(n575), .Z(n1104) );
  CNIVX1 U1336 ( .A(n605), .Z(n1105) );
  CNIVX1 U1337 ( .A(n604), .Z(n1106) );
  CNIVX1 U1338 ( .A(n1108), .Z(n1107) );
  CNIVX1 U1339 ( .A(push0_p1), .Z(n1108) );
  CNIVX1 U1340 ( .A(n601), .Z(n1109) );
  CNIVX1 U1341 ( .A(n597), .Z(n1110) );
  CNIVX1 U1342 ( .A(n658), .Z(n1111) );
  CNIVX1 U1343 ( .A(n660), .Z(n1112) );
  CNIVX1 U1344 ( .A(n662), .Z(n1113) );
  CNIVX1 U1345 ( .A(n666), .Z(n1114) );
  CNIVX1 U1346 ( .A(n670), .Z(n1115) );
  CNIVX1 U1347 ( .A(n678), .Z(n1116) );
  CMX2XL U1348 ( .A0(q0[20]), .A1(q[20]), .S(n1339), .Z(n678) );
  CNIVX1 U1349 ( .A(n582), .Z(n1117) );
  CNIVX1 U1350 ( .A(n598), .Z(n1118) );
  CNIVX1 U1351 ( .A(n580), .Z(n1119) );
  CNIVX1 U1352 ( .A(n600), .Z(n1120) );
  CNIVX1 U1353 ( .A(n586), .Z(n1121) );
  CNIVX1 U1354 ( .A(n608), .Z(n1122) );
  CNIVX1 U1355 ( .A(n602), .Z(n1123) );
  CNIVX1 U1356 ( .A(n596), .Z(n1124) );
  CNIVX1 U1357 ( .A(n606), .Z(n1125) );
  CNIVX1 U1358 ( .A(n610), .Z(n1126) );
  CNIVX1 U1359 ( .A(n584), .Z(n1127) );
  CNIVX1 U1360 ( .A(h0[0]), .Z(n1128) );
  CNIVX1 U1361 ( .A(n568), .Z(n1129) );
  CNIVX1 U1362 ( .A(n1131), .Z(n1130) );
  CNIVX1 U1363 ( .A(en1_p1), .Z(n1131) );
  CNIVX1 U1364 ( .A(n576), .Z(n1132) );
  CNIVX1 U1365 ( .A(n570), .Z(n1133) );
  CNIVX1 U1366 ( .A(n572), .Z(n1134) );
  CNIVX1 U1367 ( .A(n599), .Z(n1135) );
  CNIVX1 U1368 ( .A(n607), .Z(n1136) );
  CNIVX1 U1369 ( .A(n564), .Z(n1137) );
  CNIVX1 U1370 ( .A(n566), .Z(n1138) );
  CNIVX1 U1371 ( .A(n565), .Z(n1139) );
  CNIVX1 U1372 ( .A(n577), .Z(n1140) );
  CNIVX1 U1373 ( .A(n569), .Z(n1141) );
  CNIVX1 U1374 ( .A(n603), .Z(n1142) );
  CNIVX1 U1375 ( .A(n555), .Z(n1143) );
  CNIVX1 U1376 ( .A(n649), .Z(n1144) );
  CNIVX1 U1377 ( .A(n589), .Z(n1145) );
  CNIVX1 U1378 ( .A(n561), .Z(n1146) );
  CNIVX1 U1379 ( .A(n579), .Z(n1147) );
  CNIVX1 U1380 ( .A(n571), .Z(n1148) );
  CNIVX1 U1381 ( .A(n587), .Z(n1149) );
  CNIVX1 U1382 ( .A(n557), .Z(n1150) );
  CNIVX1 U1383 ( .A(n593), .Z(n1151) );
  CNIVX1 U1384 ( .A(n595), .Z(n1152) );
  CNIVX1 U1385 ( .A(n563), .Z(n1153) );
  CNIVX1 U1386 ( .A(n635), .Z(n1154) );
  CNIVX1 U1387 ( .A(n574), .Z(n1155) );
  CNIVX1 U1388 ( .A(n657), .Z(n1156) );
  CNIVX1 U1389 ( .A(n651), .Z(n1157) );
  CIVX4 U1390 ( .A(rst), .Z(n1937) );
  CDLY1XL U1391 ( .A(q0[29]), .Z(n1158) );
  CDLY1XL U1392 ( .A(q0[25]), .Z(n1159) );
  CDLY1XL U1393 ( .A(q0[10]), .Z(n1160) );
  CDLY1XL U1394 ( .A(q0[21]), .Z(n1161) );
  CMX2XL U1395 ( .A0(n1160), .A1(q[10]), .S(n1340), .Z(n668) );
  CDLY1XL U1396 ( .A(q0[19]), .Z(n1162) );
  CDLY1XL U1397 ( .A(q0[1]), .Z(n1163) );
  CMX2XL U1398 ( .A0(q0[28]), .A1(q[28]), .S(n1339), .Z(n686) );
  CDLY1XL U1399 ( .A(q0[9]), .Z(n1164) );
  CDLY1XL U1400 ( .A(q0[17]), .Z(n1165) );
  CDLY1XL U1401 ( .A(q0[6]), .Z(n1171) );
  CDLY1XL U1402 ( .A(q0[15]), .Z(n1166) );
  CMX2XL U1403 ( .A0(q0[18]), .A1(q[18]), .S(n1340), .Z(n676) );
  CMX2XL U1404 ( .A0(n1236), .A1(q[14]), .S(n1340), .Z(n672) );
  CDLY1XL U1405 ( .A(q0[3]), .Z(n1167) );
  CDLY1XL U1406 ( .A(q0[11]), .Z(n1168) );
  CMX2XL U1407 ( .A0(h0[25]), .A1(h[25]), .S(n1342), .Z(n651) );
  CDLY1XL U1408 ( .A(q0[23]), .Z(n1169) );
  CMX2XL U1409 ( .A0(n1164), .A1(q[9]), .S(n1340), .Z(n667) );
  CDLY1XL U1410 ( .A(q0[7]), .Z(n1170) );
  CMX2XL U1411 ( .A0(n1159), .A1(q[25]), .S(n1339), .Z(n683) );
  CMX2XL U1412 ( .A0(h0[8]), .A1(h[8]), .S(n1343), .Z(n634) );
  CMX2XL U1413 ( .A0(h0[16]), .A1(h[16]), .S(n1342), .Z(n642) );
  CDLY1XL U1414 ( .A(q0[5]), .Z(n1172) );
  CMX2XL U1415 ( .A0(h0[11]), .A1(h[11]), .S(n1343), .Z(n637) );
  CMX2XL U1416 ( .A0(h0[13]), .A1(h[13]), .S(n1343), .Z(n639) );
  CDLY1XL U1417 ( .A(q0[13]), .Z(n1173) );
  CMX2XL U1418 ( .A0(n1168), .A1(q[11]), .S(n1340), .Z(n669) );
  CMX2XL U1419 ( .A0(h0[12]), .A1(h[12]), .S(n1343), .Z(n638) );
  CDLY1XL U1420 ( .A(q0[27]), .Z(n1237) );
  CIVXL U1421 ( .A(n1073), .Z(n1867) );
  CMX2XL U1422 ( .A0(n1073), .A1(h[4]), .S(n1343), .Z(n626) );
  CMX2XL U1423 ( .A0(n927), .A1(h[2]), .S(n1344), .Z(n620) );
  CIVXL U1424 ( .A(n927), .Z(n1871) );
  CMX2XL U1425 ( .A0(n925), .A1(h[1]), .S(n1344), .Z(n617) );
  CIVXL U1426 ( .A(n925), .Z(n1873) );
  CMX2XL U1427 ( .A0(n933), .A1(h[6]), .S(n1343), .Z(n632) );
  CIVXL U1428 ( .A(n933), .Z(n1863) );
  CMX2XL U1429 ( .A0(n931), .A1(h[5]), .S(n1343), .Z(n629) );
  CIVXL U1430 ( .A(n931), .Z(n1865) );
  CMX2XL U1431 ( .A0(n1165), .A1(q[17]), .S(n1340), .Z(n675) );
  CMXI2XL U1432 ( .A0(n2258), .A1(n2257), .S(n1239), .Z(n2260) );
  CMXI2XL U1433 ( .A0(n2237), .A1(n2236), .S(n1243), .Z(n2239) );
  CNR2XL U1434 ( .A(n2060), .B(n1239), .Z(n2129) );
  CNIVX1 U1435 ( .A(en2_p2), .Z(n1255) );
  CND3X1 U1436 ( .A(n1252), .B(n1394), .C(n1345), .Z(n1395) );
  CANR2X1 U1437 ( .A(acc[57]), .B(n1856), .C(out1_p2[57]), .D(n1855), .Z(n1843) );
  CANR2XL U1438 ( .A(n1719), .B(acc[24]), .C(n1718), .D(out0_p2[24]), .Z(n1622) );
  CNR2X1 U1439 ( .A(n2151), .B(n1248), .Z(n2235) );
  CNR2X1 U1440 ( .A(n2147), .B(n1244), .Z(n2234) );
  CNR2X1 U1441 ( .A(n2155), .B(n1244), .Z(n2244) );
  CNR2X1 U1442 ( .A(n2208), .B(n1245), .Z(n2233) );
  CNR2X1 U1443 ( .A(n2179), .B(n1247), .Z(n2247) );
  CNR2X1 U1444 ( .A(n2159), .B(n1249), .Z(n2245) );
  CNR2X1 U1445 ( .A(n2175), .B(n1248), .Z(n2246) );
  COND1XL U1446 ( .A(n1269), .B(n1844), .C(n1843), .Z(acc_cmd2[57]) );
  COND1XL U1447 ( .A(n1265), .B(n1730), .C(n1729), .Z(acc_cmd2[63]) );
  CMXI2X1 U1448 ( .A0(n1955), .A1(n2248), .S(n1251), .Z(n1231) );
  CNR3XL U1449 ( .A(n1945), .B(n1251), .C(n1250), .Z(N401) );
  CNR3XL U1450 ( .A(n1942), .B(n1251), .C(n1250), .Z(N398) );
  CMXI2XL U1451 ( .A0(n2025), .A1(n2028), .S(n1328), .Z(n2059) );
  CMXI2XL U1452 ( .A0(n1978), .A1(n1977), .S(n1327), .Z(n2041) );
  CMXI2XL U1453 ( .A0(n1980), .A1(n1979), .S(n1327), .Z(n2044) );
  CMXI2XL U1454 ( .A0(n1976), .A1(n1975), .S(n1327), .Z(n2042) );
  CMXI2XL U1455 ( .A0(n1974), .A1(n1973), .S(n1327), .Z(n2038) );
  CMXI2XL U1456 ( .A0(n1971), .A1(n1970), .S(n1326), .Z(n2039) );
  CMXI2XL U1457 ( .A0(n1969), .A1(n1968), .S(n1326), .Z(n2036) );
  CMXI2XL U1458 ( .A0(n2135), .A1(n2134), .S(n1335), .Z(n2207) );
  CMXI2XL U1459 ( .A0(n1967), .A1(n1966), .S(n1326), .Z(n2037) );
  CMXI2XL U1460 ( .A0(n1965), .A1(n1964), .S(n1326), .Z(n2034) );
  CMXI2XL U1461 ( .A0(n1963), .A1(n1962), .S(n1326), .Z(n2035) );
  CMXI2XL U1462 ( .A0(n1961), .A1(n1960), .S(n1326), .Z(n2032) );
  CMXI2XL U1463 ( .A0(n2125), .A1(n2128), .S(n1333), .Z(n2178) );
  CMXI2XL U1464 ( .A0(n2118), .A1(n2121), .S(n1333), .Z(n2174) );
  CMXI2XL U1465 ( .A0(n2111), .A1(n2114), .S(n1333), .Z(n2158) );
  CMXI2XL U1466 ( .A0(n2087), .A1(n2090), .S(n1332), .Z(n2150) );
  CMXI2XL U1467 ( .A0(n2080), .A1(n2083), .S(n1332), .Z(n2146) );
  CMXI2XL U1468 ( .A0(n2140), .A1(n2139), .S(n1335), .Z(n2273) );
  CMXI2XL U1469 ( .A0(n2133), .A1(n2132), .S(n1335), .Z(n2267) );
  CMXI2XL U1470 ( .A0(n1959), .A1(n1958), .S(n1326), .Z(n2033) );
  CMXI2XL U1471 ( .A0(n1957), .A1(n1956), .S(n1326), .Z(n2249) );
  CMXI2XL U1472 ( .A0(n2164), .A1(n2163), .S(n1330), .Z(n2250) );
  CMXI2XL U1473 ( .A0(n2259), .A1(n2126), .S(n1333), .Z(n2055) );
  CMXI2XL U1474 ( .A0(n2251), .A1(n2119), .S(n1333), .Z(n2040) );
  CMXI2XL U1475 ( .A0(n2238), .A1(n2112), .S(n1333), .Z(n2020) );
  CMXI2XL U1476 ( .A0(n2200), .A1(n2088), .S(n1332), .Z(n1986) );
  CMXI2XL U1477 ( .A0(n2166), .A1(n2081), .S(n1332), .Z(n1972) );
  CMXI2XL U1478 ( .A0(n2272), .A1(n2271), .S(n1336), .Z(n2274) );
  CMXI2XL U1479 ( .A0(n2266), .A1(n2265), .S(n1336), .Z(n2268) );
  CNR2X1 U1480 ( .A(n2077), .B(n1241), .Z(n2115) );
  CNR2X1 U1481 ( .A(n2045), .B(n1240), .Z(n2122) );
  CMXI2XL U1482 ( .A0(n1180), .A1(n1181), .S(n1318), .Z(n2023) );
  CMXI2XL U1483 ( .A0(n2000), .A1(n1999), .S(n1239), .Z(n2109) );
  CMXI2XL U1484 ( .A0(n1178), .A1(n1179), .S(n1318), .Z(n2024) );
  CMXI2XL U1485 ( .A0(n1182), .A1(n1183), .S(n1318), .Z(n2026) );
  CMXI2XL U1486 ( .A0(n1194), .A1(n1177), .S(n1319), .Z(n2021) );
  CMXI2XL U1487 ( .A0(n1184), .A1(n1175), .S(n1318), .Z(n2025) );
  CMXI2XL U1488 ( .A0(n1195), .A1(n1196), .S(n1319), .Z(n2022) );
  CMXI2XL U1489 ( .A0(n1998), .A1(n1997), .S(n1243), .Z(n2106) );
  CMXI2XL U1490 ( .A0(n1200), .A1(n1199), .S(n1320), .Z(n2018) );
  CMXI2XL U1491 ( .A0(n1197), .A1(n1198), .S(n1319), .Z(n2019) );
  CMXI2XL U1492 ( .A0(n1187), .A1(n1186), .S(n1319), .Z(n2016) );
  CMXI2XL U1493 ( .A0(n1188), .A1(n1189), .S(n1319), .Z(n2017) );
  CMXI2XL U1494 ( .A0(n1191), .A1(n1190), .S(n1319), .Z(n2014) );
  CMXI2XL U1495 ( .A0(n1192), .A1(n1193), .S(n1319), .Z(n2015) );
  CMXI2XL U1496 ( .A0(n1995), .A1(n1994), .S(n1242), .Z(n2107) );
  CMXI2XL U1497 ( .A0(n1202), .A1(n1201), .S(n1319), .Z(n2012) );
  CMXI2XL U1498 ( .A0(n1203), .A1(n1204), .S(n1319), .Z(n2013) );
  CMXI2XL U1499 ( .A0(n1206), .A1(n1205), .S(n1319), .Z(n2010) );
  CMXI2XL U1500 ( .A0(n1207), .A1(n1208), .S(n1319), .Z(n2011) );
  CMXI2XL U1501 ( .A0(n1210), .A1(n1209), .S(n1320), .Z(n2008) );
  CMXI2XL U1502 ( .A0(n1211), .A1(n1212), .S(n1320), .Z(n2009) );
  CMXI2XL U1503 ( .A0(n1214), .A1(n1213), .S(n1320), .Z(n2006) );
  CMXI2XL U1504 ( .A0(n1215), .A1(n1216), .S(n1320), .Z(n2007) );
  CMXI2XL U1505 ( .A0(n1993), .A1(n1992), .S(n1239), .Z(n2104) );
  CMXI2XL U1506 ( .A0(n1991), .A1(n1990), .S(n1242), .Z(n2105) );
  CMXI2XL U1507 ( .A0(n1218), .A1(n1217), .S(n1320), .Z(n2004) );
  CMXI2XL U1508 ( .A0(n1219), .A1(n1220), .S(n1320), .Z(n2005) );
  CMXI2XL U1509 ( .A0(n1222), .A1(n1221), .S(n1320), .Z(n2096) );
  CMXI2XL U1510 ( .A0(n1223), .A1(n1224), .S(n1318), .Z(n2197) );
  CMXI2XL U1511 ( .A0(n1989), .A1(n1988), .S(n1241), .Z(n2220) );
  CMXI2XL U1512 ( .A0(n1226), .A1(n1225), .S(n1318), .Z(n2198) );
  CMXI2XL U1513 ( .A0(n1227), .A1(n1228), .S(n1318), .Z(n2195) );
  CMXI2XL U1514 ( .A0(n1185), .A1(n1229), .S(n1318), .Z(n2196) );
  CMXI2XL U1515 ( .A0(n2260), .A1(n2259), .S(n1336), .Z(n2262) );
  CMXI2XL U1516 ( .A0(n2252), .A1(n2251), .S(n1336), .Z(n2254) );
  CMXI2XL U1517 ( .A0(n2250), .A1(n2249), .S(n1241), .Z(n2252) );
  CMXI2XL U1518 ( .A0(n2239), .A1(n2238), .S(n1336), .Z(n2241) );
  CMXI2XL U1519 ( .A0(n2221), .A1(n2220), .S(n1336), .Z(n2223) );
  CMXI2XL U1520 ( .A0(n2219), .A1(n2218), .S(n1242), .Z(n2221) );
  CMXI2XL U1521 ( .A0(n2201), .A1(n2200), .S(n1336), .Z(n2203) );
  CMXI2XL U1522 ( .A0(n2196), .A1(n2195), .S(n1330), .Z(n2199) );
  CMXI2XL U1523 ( .A0(n2167), .A1(n2166), .S(n1336), .Z(n2169) );
  CMXI2XL U1524 ( .A0(n2162), .A1(n2161), .S(n1329), .Z(n2165) );
  CMXI2XL U1525 ( .A0(n2098), .A1(n2272), .S(n1334), .Z(n2100) );
  CMXI2XL U1526 ( .A0(n1862), .A1(n1230), .S(n1318), .Z(n2094) );
  CND2XL U1527 ( .A(n1983), .B(n1331), .Z(n2001) );
  CIVXL U1528 ( .A(n1861), .Z(n1862) );
  CANR2XL U1529 ( .A(n1719), .B(acc[28]), .C(n1718), .D(out0_p2[28]), .Z(n1606) );
  CANR2XL U1530 ( .A(n1719), .B(acc[16]), .C(n1718), .D(out0_p2[16]), .Z(n1654) );
  CANR2XL U1531 ( .A(n1719), .B(acc[40]), .C(n1718), .D(out0_p2[40]), .Z(n1558) );
  CANR2XL U1532 ( .A(n1719), .B(acc[48]), .C(n1718), .D(out0_p2[48]), .Z(n1526) );
  CANR2XL U1533 ( .A(n1719), .B(acc[52]), .C(n1718), .D(out0_p2[52]), .Z(n1510) );
  CANR2XL U1534 ( .A(n1719), .B(acc[36]), .C(n1718), .D(out0_p2[36]), .Z(n1574) );
  CANR2XL U1535 ( .A(n1719), .B(acc[60]), .C(n1718), .D(out0_p2[60]), .Z(n1478) );
  CANR2XL U1536 ( .A(n1719), .B(acc[20]), .C(n1718), .D(out0_p2[20]), .Z(n1638) );
  CANR2XL U1537 ( .A(acc[56]), .B(n1856), .C(out1_p2[56]), .D(n1855), .Z(n1847) );
  CANR2XL U1538 ( .A(acc[55]), .B(n1856), .C(out1_p2[55]), .D(n1855), .Z(n1845) );
  CANR2XL U1539 ( .A(acc[31]), .B(n1856), .C(out1_p2[31]), .D(n1855), .Z(n1793) );
  CANR2XL U1540 ( .A(acc[32]), .B(n1856), .C(out1_p2[32]), .D(n1855), .Z(n1795) );
  CANR2XL U1541 ( .A(acc[35]), .B(n1856), .C(out1_p2[35]), .D(n1855), .Z(n1801) );
  CANR2XL U1542 ( .A(acc[47]), .B(n1856), .C(out1_p2[47]), .D(n1855), .Z(n1825) );
  CANR2XL U1543 ( .A(acc[36]), .B(n1856), .C(out1_p2[36]), .D(n1855), .Z(n1803) );
  CANR2XL U1544 ( .A(acc[48]), .B(n1856), .C(out1_p2[48]), .D(n1855), .Z(n1827) );
  CANR2XL U1545 ( .A(acc[51]), .B(n1856), .C(out1_p2[51]), .D(n1855), .Z(n1833) );
  CANR2XL U1546 ( .A(acc[52]), .B(n1856), .C(out1_p2[52]), .D(n1855), .Z(n1835) );
  CANR2XL U1547 ( .A(acc[39]), .B(n1856), .C(out1_p2[39]), .D(n1855), .Z(n1809) );
  CANR2XL U1548 ( .A(acc[33]), .B(n1856), .C(out1_p2[33]), .D(n1855), .Z(n1797) );
  CANR2XL U1549 ( .A(acc[40]), .B(n1856), .C(out1_p2[40]), .D(n1855), .Z(n1811) );
  CANR2XL U1550 ( .A(acc[34]), .B(n1856), .C(out1_p2[34]), .D(n1855), .Z(n1799) );
  CANR2XL U1551 ( .A(acc[43]), .B(n1856), .C(out1_p2[43]), .D(n1855), .Z(n1817) );
  CANR2XL U1552 ( .A(acc[37]), .B(n1856), .C(out1_p2[37]), .D(n1855), .Z(n1805) );
  CANR2XL U1553 ( .A(acc[49]), .B(n1856), .C(out1_p2[49]), .D(n1855), .Z(n1829) );
  CANR2XL U1554 ( .A(acc[44]), .B(n1856), .C(out1_p2[44]), .D(n1855), .Z(n1819) );
  CANR2XL U1555 ( .A(acc[38]), .B(n1856), .C(out1_p2[38]), .D(n1855), .Z(n1807) );
  CANR2XL U1556 ( .A(acc[50]), .B(n1856), .C(out1_p2[50]), .D(n1855), .Z(n1831) );
  CANR2XL U1557 ( .A(acc[53]), .B(n1856), .C(out1_p2[53]), .D(n1855), .Z(n1837) );
  CANR2XL U1558 ( .A(acc[54]), .B(n1856), .C(out1_p2[54]), .D(n1855), .Z(n1839) );
  CANR2XL U1559 ( .A(acc[41]), .B(n1856), .C(out1_p2[41]), .D(n1855), .Z(n1813) );
  CANR2XL U1560 ( .A(acc[42]), .B(n1856), .C(out1_p2[42]), .D(n1855), .Z(n1815) );
  CANR2XL U1561 ( .A(acc[45]), .B(n1856), .C(out1_p2[45]), .D(n1855), .Z(n1821) );
  CANR2XL U1562 ( .A(acc[46]), .B(n1856), .C(out1_p2[46]), .D(n1855), .Z(n1823) );
  CANR2XL U1563 ( .A(acc[15]), .B(n1856), .C(out1_p2[15]), .D(n1855), .Z(n1761) );
  CANR2XL U1564 ( .A(acc[16]), .B(n1856), .C(out1_p2[16]), .D(n1855), .Z(n1763) );
  CANR2XL U1565 ( .A(acc[19]), .B(n1856), .C(out1_p2[19]), .D(n1855), .Z(n1769) );
  CANR2XL U1566 ( .A(acc[20]), .B(n1856), .C(out1_p2[20]), .D(n1855), .Z(n1771) );
  CANR2XL U1567 ( .A(acc[23]), .B(n1856), .C(out1_p2[23]), .D(n1855), .Z(n1777) );
  CANR2XL U1568 ( .A(acc[17]), .B(n1856), .C(out1_p2[17]), .D(n1855), .Z(n1765) );
  CANR2XL U1569 ( .A(acc[24]), .B(n1856), .C(out1_p2[24]), .D(n1855), .Z(n1779) );
  CANR2XL U1570 ( .A(acc[18]), .B(n1856), .C(out1_p2[18]), .D(n1855), .Z(n1767) );
  CANR2XL U1571 ( .A(acc[27]), .B(n1856), .C(out1_p2[27]), .D(n1855), .Z(n1785) );
  CANR2XL U1572 ( .A(acc[21]), .B(n1856), .C(out1_p2[21]), .D(n1855), .Z(n1773) );
  CANR2XL U1573 ( .A(acc[28]), .B(n1856), .C(out1_p2[28]), .D(n1855), .Z(n1787) );
  CANR2XL U1574 ( .A(acc[22]), .B(n1856), .C(out1_p2[22]), .D(n1855), .Z(n1775) );
  CANR2XL U1575 ( .A(acc[25]), .B(n1856), .C(out1_p2[25]), .D(n1855), .Z(n1781) );
  CANR2XL U1576 ( .A(acc[26]), .B(n1856), .C(out1_p2[26]), .D(n1855), .Z(n1783) );
  CANR2XL U1577 ( .A(acc[29]), .B(n1856), .C(out1_p2[29]), .D(n1855), .Z(n1789) );
  CANR2XL U1578 ( .A(acc[30]), .B(n1856), .C(out1_p2[30]), .D(n1855), .Z(n1791) );
  CANR2XL U1579 ( .A(acc[7]), .B(n1856), .C(out1_p2[7]), .D(n1855), .Z(n1745)
         );
  CANR2XL U1580 ( .A(acc[8]), .B(n1856), .C(out1_p2[8]), .D(n1855), .Z(n1747)
         );
  CANR2XL U1581 ( .A(acc[11]), .B(n1856), .C(out1_p2[11]), .D(n1855), .Z(n1753) );
  CANR2XL U1582 ( .A(acc[12]), .B(n1856), .C(out1_p2[12]), .D(n1855), .Z(n1755) );
  CANR2XL U1583 ( .A(acc[9]), .B(n1856), .C(out1_p2[9]), .D(n1855), .Z(n1749)
         );
  CANR2XL U1584 ( .A(acc[10]), .B(n1856), .C(out1_p2[10]), .D(n1855), .Z(n1751) );
  CANR2XL U1585 ( .A(acc[13]), .B(n1856), .C(out1_p2[13]), .D(n1855), .Z(n1757) );
  CANR2XL U1586 ( .A(acc[14]), .B(n1856), .C(out1_p2[14]), .D(n1855), .Z(n1759) );
  CANR2XL U1587 ( .A(acc[3]), .B(n1856), .C(out1_p2[3]), .D(n1855), .Z(n1737)
         );
  CANR2XL U1588 ( .A(acc[4]), .B(n1856), .C(out1_p2[4]), .D(n1855), .Z(n1739)
         );
  CANR2XL U1589 ( .A(acc[5]), .B(n1856), .C(out1_p2[5]), .D(n1855), .Z(n1741)
         );
  CANR2XL U1590 ( .A(acc[6]), .B(n1856), .C(out1_p2[6]), .D(n1855), .Z(n1743)
         );
  CANR2XL U1591 ( .A(acc[1]), .B(n1856), .C(out1_p2[1]), .D(n1855), .Z(n1733)
         );
  CANR2XL U1592 ( .A(acc[2]), .B(n1856), .C(out1_p2[2]), .D(n1855), .Z(n1735)
         );
  CANR2XL U1593 ( .A(acc[63]), .B(n1856), .C(out1_p2[63]), .D(n1855), .Z(n1729) );
  CANR2XL U1594 ( .A(acc[61]), .B(n1856), .C(out1_p2[61]), .D(n1855), .Z(n1857) );
  CANR2XL U1595 ( .A(acc[60]), .B(n1856), .C(out1_p2[60]), .D(n1855), .Z(n1849) );
  CANR2XL U1596 ( .A(n1719), .B(acc[18]), .C(n1718), .D(out0_p2[18]), .Z(n1646) );
  CANR2XL U1597 ( .A(acc[59]), .B(n1856), .C(out1_p2[59]), .D(n1855), .Z(n1851) );
  CANR2XL U1598 ( .A(n1719), .B(acc[11]), .C(n1718), .D(out0_p2[11]), .Z(n1674) );
  CANR2XL U1599 ( .A(n1719), .B(acc[10]), .C(n1718), .D(out0_p2[10]), .Z(n1678) );
  CANR2XL U1600 ( .A(n1719), .B(acc[2]), .C(n1718), .D(out0_p2[2]), .Z(n1710)
         );
  CANR2XL U1601 ( .A(n1719), .B(acc[23]), .C(n1718), .D(out0_p2[23]), .Z(n1626) );
  CANR2XL U1602 ( .A(n1719), .B(acc[17]), .C(n1718), .D(out0_p2[17]), .Z(n1650) );
  CANR2XL U1603 ( .A(n1719), .B(acc[22]), .C(n1718), .D(out0_p2[22]), .Z(n1630) );
  CANR2XL U1604 ( .A(n1719), .B(acc[25]), .C(n1718), .D(out0_p2[25]), .Z(n1618) );
  CANR2XL U1605 ( .A(n1719), .B(acc[8]), .C(n1718), .D(out0_p2[8]), .Z(n1686)
         );
  CANR2XL U1606 ( .A(n1719), .B(acc[19]), .C(n1718), .D(out0_p2[19]), .Z(n1642) );
  CANR2XL U1607 ( .A(n1719), .B(acc[26]), .C(n1718), .D(out0_p2[26]), .Z(n1614) );
  CANR2XL U1608 ( .A(n1719), .B(acc[6]), .C(n1718), .D(out0_p2[6]), .Z(n1694)
         );
  CANR2XL U1609 ( .A(n1719), .B(acc[27]), .C(n1718), .D(out0_p2[27]), .Z(n1610) );
  CANR2XL U1610 ( .A(n1719), .B(acc[1]), .C(n1718), .D(out0_p2[1]), .Z(n1714)
         );
  CANR2XL U1611 ( .A(n1719), .B(acc[29]), .C(n1718), .D(out0_p2[29]), .Z(n1602) );
  CANR2XL U1612 ( .A(n1719), .B(acc[14]), .C(n1718), .D(out0_p2[14]), .Z(n1662) );
  CANR2XL U1613 ( .A(n1719), .B(acc[35]), .C(n1718), .D(out0_p2[35]), .Z(n1578) );
  CANR2XL U1614 ( .A(n1719), .B(acc[15]), .C(n1718), .D(out0_p2[15]), .Z(n1658) );
  CANR2XL U1615 ( .A(n1719), .B(acc[3]), .C(n1718), .D(out0_p2[3]), .Z(n1706)
         );
  CANR2XL U1616 ( .A(n1719), .B(acc[7]), .C(n1718), .D(out0_p2[7]), .Z(n1690)
         );
  CANR2XL U1617 ( .A(n1719), .B(acc[13]), .C(n1718), .D(out0_p2[13]), .Z(n1666) );
  CANR2XL U1618 ( .A(acc[0]), .B(n1856), .C(out1_p2[0]), .D(n1855), .Z(n1731)
         );
  CANR2XL U1619 ( .A(n1719), .B(acc[41]), .C(n1718), .D(out0_p2[41]), .Z(n1554) );
  CANR2XL U1620 ( .A(n1719), .B(acc[21]), .C(n1718), .D(out0_p2[21]), .Z(n1634) );
  CANR2XL U1621 ( .A(n1719), .B(acc[5]), .C(n1718), .D(out0_p2[5]), .Z(n1698)
         );
  CANR2XL U1622 ( .A(n1719), .B(acc[12]), .C(n1718), .D(out0_p2[12]), .Z(n1670) );
  CANR2XL U1623 ( .A(n1719), .B(acc[30]), .C(n1718), .D(out0_p2[30]), .Z(n1598) );
  CANR2XL U1624 ( .A(n1719), .B(acc[31]), .C(n1718), .D(out0_p2[31]), .Z(n1594) );
  CANR2XL U1625 ( .A(n1719), .B(acc[33]), .C(n1718), .D(out0_p2[33]), .Z(n1586) );
  CANR2XL U1626 ( .A(n1719), .B(acc[49]), .C(n1718), .D(out0_p2[49]), .Z(n1522) );
  CANR2XL U1627 ( .A(n1719), .B(acc[0]), .C(n1718), .D(out0_p2[0]), .Z(n1720)
         );
  CANR2XL U1628 ( .A(n1719), .B(acc[34]), .C(n1718), .D(out0_p2[34]), .Z(n1582) );
  CANR2XL U1629 ( .A(n1719), .B(acc[42]), .C(n1718), .D(out0_p2[42]), .Z(n1550) );
  CANR2XL U1630 ( .A(n1719), .B(acc[43]), .C(n1718), .D(out0_p2[43]), .Z(n1546) );
  CANR2XL U1631 ( .A(n1719), .B(acc[4]), .C(n1718), .D(out0_p2[4]), .Z(n1702)
         );
  CANR2XL U1632 ( .A(n1719), .B(acc[58]), .C(n1718), .D(out0_p2[58]), .Z(n1486) );
  CANR2XL U1633 ( .A(n1719), .B(acc[57]), .C(n1718), .D(out0_p2[57]), .Z(n1490) );
  CANR2XL U1634 ( .A(n1719), .B(acc[50]), .C(n1718), .D(out0_p2[50]), .Z(n1518) );
  CANR2XL U1635 ( .A(n1719), .B(acc[51]), .C(n1718), .D(out0_p2[51]), .Z(n1514) );
  CANR2XL U1636 ( .A(n1719), .B(acc[56]), .C(n1718), .D(out0_p2[56]), .Z(n1494) );
  CANR2XL U1637 ( .A(n1719), .B(acc[32]), .C(n1718), .D(out0_p2[32]), .Z(n1590) );
  CANR2XL U1638 ( .A(n1719), .B(acc[59]), .C(n1718), .D(out0_p2[59]), .Z(n1482) );
  CANR2XL U1639 ( .A(n1719), .B(acc[44]), .C(n1718), .D(out0_p2[44]), .Z(n1542) );
  CANR2XL U1640 ( .A(n1719), .B(acc[45]), .C(n1718), .D(out0_p2[45]), .Z(n1538) );
  CMXI2XL U1641 ( .A0(n2063), .A1(n2062), .S(n1248), .Z(n2066) );
  CANR2XL U1642 ( .A(n2181), .B(n1174), .C(n2182), .D(n1264), .Z(n1396) );
  CANR2XL U1643 ( .A(n1719), .B(acc[47]), .C(n1718), .D(out0_p2[47]), .Z(n1530) );
  CANR2XL U1644 ( .A(n1719), .B(acc[53]), .C(n1718), .D(out0_p2[53]), .Z(n1506) );
  CANR2XL U1645 ( .A(n1719), .B(acc[38]), .C(n1718), .D(out0_p2[38]), .Z(n1566) );
  CANR2XL U1646 ( .A(n1719), .B(acc[55]), .C(n1718), .D(out0_p2[55]), .Z(n1498) );
  CANR2XL U1647 ( .A(n1719), .B(acc[39]), .C(n1718), .D(out0_p2[39]), .Z(n1562) );
  CANR2XL U1648 ( .A(n1719), .B(acc[46]), .C(n1718), .D(out0_p2[46]), .Z(n1534) );
  CANR2XL U1649 ( .A(n1719), .B(acc[54]), .C(n1718), .D(out0_p2[54]), .Z(n1502) );
  CANR2XL U1650 ( .A(n1719), .B(acc[37]), .C(n1718), .D(out0_p2[37]), .Z(n1570) );
  CANR2XL U1651 ( .A(n1719), .B(acc[61]), .C(n1718), .D(out0_p2[61]), .Z(n1474) );
  CANR2XL U1652 ( .A(n1719), .B(acc[62]), .C(n1718), .D(out0_p2[62]), .Z(n1470) );
  CANR2XL U1653 ( .A(n1719), .B(acc[63]), .C(n1718), .D(out0_p2[63]), .Z(n1464) );
  CANR2XL U1654 ( .A(n1234), .B(out0_p2[11]), .C(N429), .D(n1233), .Z(n1673)
         );
  CANR2XL U1655 ( .A(n1234), .B(out0_p2[9]), .C(N427), .D(n1233), .Z(n1681) );
  CANR2XL U1656 ( .A(n1234), .B(out0_p2[3]), .C(N421), .D(n1233), .Z(n1705) );
  CANR2XL U1657 ( .A(n1234), .B(out0_p2[1]), .C(N419), .D(n1233), .Z(n1713) );
  CIVXL U1658 ( .A(n2233), .Z(n1942) );
  CIVXL U1659 ( .A(n2234), .Z(n1943) );
  CIVXL U1660 ( .A(n2235), .Z(n1944) );
  CIVXL U1661 ( .A(n2244), .Z(n1945) );
  CNR2XL U1662 ( .A(n1251), .B(n2248), .Z(N405) );
  CIVXL U1663 ( .A(n2246), .Z(n1947) );
  CIVXL U1664 ( .A(n2245), .Z(n1946) );
  CIVXL U1665 ( .A(n2247), .Z(n1948) );
  CIVX2 U1666 ( .A(n1395), .Z(n1264) );
  CIVX4 U1667 ( .A(n1461), .Z(n1722) );
  CIVX4 U1668 ( .A(n1462), .Z(n1719) );
  CIVX2 U1669 ( .A(n1331), .Z(n1327) );
  CIVX2 U1670 ( .A(n1331), .Z(n1326) );
  CIVX2 U1671 ( .A(n1331), .Z(n1328) );
  CIVX2 U1672 ( .A(n1331), .Z(n1329) );
  CIVX2 U1673 ( .A(n1324), .Z(n1318) );
  CIVX2 U1674 ( .A(n1324), .Z(n1320) );
  CIVX2 U1675 ( .A(n1324), .Z(n1321) );
  CIVX2 U1676 ( .A(n1324), .Z(n1322) );
  CIVX2 U1677 ( .A(n1324), .Z(n1319) );
  CNR2X1 U1678 ( .A(n2001), .B(n1242), .Z(n2136) );
  CNR2IX1 U1679 ( .B(acc_cmd2[63]), .A(n1318), .Z(n1983) );
  CNR2X1 U1680 ( .A(n2206), .B(n1246), .Z(n2232) );
  CNR2X1 U1681 ( .A(n2193), .B(n1247), .Z(n2231) );
  CNR2X1 U1682 ( .A(n2191), .B(n1248), .Z(n2230) );
  CNR2X1 U1683 ( .A(n2189), .B(n1249), .Z(n2229) );
  CNR2X1 U1684 ( .A(n2187), .B(n1245), .Z(n2228) );
  CNR2X1 U1685 ( .A(n2185), .B(n1249), .Z(n2227) );
  CNR2X1 U1686 ( .A(n2101), .B(n1245), .Z(n2217) );
  CNR2X1 U1687 ( .A(n2170), .B(n1244), .Z(n2226) );
  CND3XL U1688 ( .A(n1253), .B(n1725), .C(n1727), .Z(n1726) );
  CNR2X1 U1689 ( .A(n2064), .B(n1246), .Z(n2181) );
  CNIVX1 U1690 ( .A(n1859), .Z(n1268) );
  CNIVX1 U1691 ( .A(n1859), .Z(n1267) );
  CNIVX1 U1692 ( .A(n1859), .Z(n1266) );
  CNIVX1 U1693 ( .A(n1859), .Z(n1269) );
  CNIVX1 U1694 ( .A(n1859), .Z(n1265) );
  CIVX2 U1695 ( .A(n1331), .Z(n1325) );
  CNIVX1 U1696 ( .A(n1859), .Z(n1270) );
  CND2XL U1697 ( .A(n2029), .B(n1331), .Z(n2060) );
  CND2X1 U1698 ( .A(n2129), .B(n1337), .Z(n2179) );
  CND2X1 U1699 ( .A(n2122), .B(n1337), .Z(n2175) );
  CND2X1 U1700 ( .A(n2115), .B(n1337), .Z(n2159) );
  CND2X1 U1701 ( .A(n2108), .B(n1337), .Z(n2155) );
  CND2X1 U1702 ( .A(n2091), .B(n1337), .Z(n2151) );
  CND2X1 U1703 ( .A(n2084), .B(n1337), .Z(n2147) );
  CND2X1 U1704 ( .A(n2143), .B(n1337), .Z(n2208) );
  CND2X1 U1705 ( .A(n2136), .B(n1337), .Z(n2064) );
  CAN3X2 U1706 ( .A(n1250), .B(n1252), .C(n1394), .Z(n1174) );
  CIVX2 U1707 ( .A(n1337), .Z(n1335) );
  CIVX2 U1708 ( .A(n1337), .Z(n1333) );
  CIVX2 U1709 ( .A(n1337), .Z(n1334) );
  CND3XL U1710 ( .A(n1252), .B(n1394), .C(n1345), .Z(n1238) );
  CNR3XL U1711 ( .A(n1936), .B(n1938), .C(n1939), .Z(_pushout_d) );
  CIVX2 U1712 ( .A(n1337), .Z(n1336) );
  CIVX2 U1713 ( .A(n1337), .Z(n1332) );
  CNIVX1 U1714 ( .A(n1937), .Z(n1303) );
  CNIVX1 U1715 ( .A(n1937), .Z(n1304) );
  CNIVX1 U1716 ( .A(n1937), .Z(n1286) );
  CNIVX1 U1717 ( .A(n1937), .Z(n1289) );
  CNIVX1 U1718 ( .A(n1937), .Z(n1301) );
  CNIVX1 U1719 ( .A(n1937), .Z(n1302) );
  CNIVX1 U1720 ( .A(n1937), .Z(n1278) );
  CNIVX1 U1721 ( .A(n1937), .Z(n1277) );
  CNIVX1 U1722 ( .A(n1937), .Z(n1276) );
  CNIVX1 U1723 ( .A(n1937), .Z(n1275) );
  CNIVX1 U1724 ( .A(n1937), .Z(n1274) );
  CNIVX1 U1725 ( .A(n1937), .Z(n1273) );
  CNIVX1 U1726 ( .A(n1937), .Z(n1288) );
  CNIVX1 U1727 ( .A(n1937), .Z(n1300) );
  CNIVX1 U1728 ( .A(n1937), .Z(n1299) );
  CNIVX1 U1729 ( .A(n1937), .Z(n1297) );
  CNIVX1 U1730 ( .A(n1937), .Z(n1296) );
  CNIVX1 U1731 ( .A(n1937), .Z(n1295) );
  CNIVX1 U1732 ( .A(n1937), .Z(n1294) );
  CNIVX1 U1733 ( .A(n1937), .Z(n1293) );
  CNIVX1 U1734 ( .A(n1937), .Z(n1298) );
  CNIVX1 U1735 ( .A(n1937), .Z(n1316) );
  CNIVX1 U1736 ( .A(n1937), .Z(n1315) );
  CNIVX1 U1737 ( .A(n1937), .Z(n1314) );
  CNIVX1 U1738 ( .A(n1937), .Z(n1313) );
  CNIVX1 U1739 ( .A(n1937), .Z(n1312) );
  CNIVX1 U1740 ( .A(n1937), .Z(n1310) );
  CNIVX1 U1741 ( .A(n1937), .Z(n1309) );
  CNIVX1 U1742 ( .A(n1937), .Z(n1287) );
  CNIVX1 U1743 ( .A(n1937), .Z(n1285) );
  CNIVX1 U1744 ( .A(n1937), .Z(n1284) );
  CNIVX1 U1745 ( .A(n1937), .Z(n1283) );
  CNIVX1 U1746 ( .A(n1937), .Z(n1311) );
  CNIVX1 U1747 ( .A(n1937), .Z(n1306) );
  CNIVX1 U1748 ( .A(n1937), .Z(n1305) );
  CNIVX1 U1749 ( .A(n1937), .Z(n1281) );
  CNIVX1 U1750 ( .A(n1937), .Z(n1279) );
  CNIVX1 U1751 ( .A(n1937), .Z(n1308) );
  CNIVX1 U1752 ( .A(n1937), .Z(n1290) );
  CNIVX1 U1753 ( .A(n1937), .Z(n1307) );
  CNIVX1 U1754 ( .A(n1937), .Z(n1282) );
  CNIVX1 U1755 ( .A(n1937), .Z(n1280) );
  CNIVX1 U1756 ( .A(n1937), .Z(n1271) );
  CNIVX1 U1757 ( .A(n1937), .Z(n1292) );
  CNIVX1 U1758 ( .A(n1937), .Z(n1291) );
  CNIVX1 U1759 ( .A(n1937), .Z(n1272) );
  CNIVX1 U1760 ( .A(n1937), .Z(n1317) );
  COND1XL U1761 ( .A(n1722), .B(n1531), .C(n1530), .Z(acc_cmd1[47]) );
  COND1XL U1762 ( .A(n1722), .B(n1527), .C(n1526), .Z(acc_cmd1[48]) );
  COND1XL U1763 ( .A(n1722), .B(n1631), .C(n1630), .Z(acc_cmd1[22]) );
  COND1XL U1764 ( .A(n1722), .B(n1627), .C(n1626), .Z(acc_cmd1[23]) );
  COND1XL U1765 ( .A(n1722), .B(n1639), .C(n1638), .Z(acc_cmd1[20]) );
  COND1XL U1766 ( .A(n1722), .B(n1623), .C(n1622), .Z(acc_cmd1[24]) );
  COND1XL U1767 ( .A(n1722), .B(n1543), .C(n1542), .Z(acc_cmd1[44]) );
  COND1XL U1768 ( .A(n1722), .B(n1607), .C(n1606), .Z(acc_cmd1[28]) );
  COND1XL U1769 ( .A(n1722), .B(n1511), .C(n1510), .Z(acc_cmd1[52]) );
  COND1XL U1770 ( .A(n1722), .B(n1615), .C(n1614), .Z(acc_cmd1[26]) );
  COND1XL U1771 ( .A(n1722), .B(n1523), .C(n1522), .Z(acc_cmd1[49]) );
  COND1XL U1772 ( .A(n1722), .B(n1519), .C(n1518), .Z(acc_cmd1[50]) );
  COND1XL U1773 ( .A(n1722), .B(n1655), .C(n1654), .Z(acc_cmd1[16]) );
  COND1XL U1774 ( .A(n1722), .B(n1635), .C(n1634), .Z(acc_cmd1[21]) );
  COND1XL U1775 ( .A(n1722), .B(n1603), .C(n1602), .Z(acc_cmd1[29]) );
  COND1XL U1776 ( .A(n1722), .B(n1507), .C(n1506), .Z(acc_cmd1[53]) );
  COND1XL U1777 ( .A(n1722), .B(n1711), .C(n1710), .Z(acc_cmd1[2]) );
  COND1XL U1778 ( .A(n1722), .B(n1595), .C(n1594), .Z(acc_cmd1[31]) );
  COND1XL U1779 ( .A(n1722), .B(n1663), .C(n1662), .Z(acc_cmd1[14]) );
  COND1XL U1780 ( .A(n1722), .B(n1503), .C(n1502), .Z(acc_cmd1[54]) );
  COND1XL U1781 ( .A(n1722), .B(n1515), .C(n1514), .Z(acc_cmd1[51]) );
  COND1XL U1782 ( .A(n1722), .B(n1671), .C(n1670), .Z(acc_cmd1[12]) );
  COND1XL U1783 ( .A(n1722), .B(n1721), .C(n1720), .Z(acc_cmd1[0]) );
  COND1XL U1784 ( .A(n1722), .B(n1495), .C(n1494), .Z(acc_cmd1[56]) );
  COND1XL U1785 ( .A(n1722), .B(n1703), .C(n1702), .Z(acc_cmd1[4]) );
  COND1XL U1786 ( .A(n1722), .B(n1499), .C(n1498), .Z(acc_cmd1[55]) );
  COND1XL U1787 ( .A(n1722), .B(n1491), .C(n1490), .Z(acc_cmd1[57]) );
  COND1XL U1788 ( .A(n1722), .B(n1487), .C(n1486), .Z(acc_cmd1[58]) );
  COND1XL U1789 ( .A(n1722), .B(n1483), .C(n1482), .Z(acc_cmd1[59]) );
  COND1XL U1790 ( .A(n1722), .B(n1475), .C(n1474), .Z(acc_cmd1[61]) );
  COND1XL U1791 ( .A(n1722), .B(n1479), .C(n1478), .Z(acc_cmd1[60]) );
  COND1XL U1792 ( .A(n1722), .B(n1471), .C(n1470), .Z(acc_cmd1[62]) );
  COND1XL U1793 ( .A(n1722), .B(n1465), .C(n1464), .Z(acc_cmd1[63]) );
  CIVX4 U1794 ( .A(n1463), .Z(n1718) );
  COND1XL U1795 ( .A(n1265), .B(n1732), .C(n1731), .Z(n1861) );
  COND1XL U1796 ( .A(n1722), .B(n1583), .C(n1582), .Z(acc_cmd1[34]) );
  COND1XL U1797 ( .A(n1722), .B(n1535), .C(n1534), .Z(acc_cmd1[46]) );
  COND1XL U1798 ( .A(n1722), .B(n1647), .C(n1646), .Z(acc_cmd1[18]) );
  COND1XL U1799 ( .A(n1722), .B(n1551), .C(n1550), .Z(acc_cmd1[42]) );
  COND1XL U1800 ( .A(n1722), .B(n1555), .C(n1554), .Z(acc_cmd1[41]) );
  COND1XL U1801 ( .A(n1722), .B(n1539), .C(n1538), .Z(acc_cmd1[45]) );
  COND1XL U1802 ( .A(n1722), .B(n1567), .C(n1566), .Z(acc_cmd1[38]) );
  COND1XL U1803 ( .A(n1722), .B(n1651), .C(n1650), .Z(acc_cmd1[17]) );
  COND1XL U1804 ( .A(n1722), .B(n1619), .C(n1618), .Z(acc_cmd1[25]) );
  COND1XL U1805 ( .A(n1722), .B(n1675), .C(n1674), .Z(acc_cmd1[11]) );
  COND1XL U1806 ( .A(n1722), .B(n1559), .C(n1558), .Z(acc_cmd1[40]) );
  COND1XL U1807 ( .A(n1722), .B(n1579), .C(n1578), .Z(acc_cmd1[35]) );
  COND1XL U1808 ( .A(n1722), .B(n1587), .C(n1586), .Z(acc_cmd1[33]) );
  COND1XL U1809 ( .A(n1722), .B(n1563), .C(n1562), .Z(acc_cmd1[39]) );
  COND1XL U1810 ( .A(n1722), .B(n1547), .C(n1546), .Z(acc_cmd1[43]) );
  COND1XL U1811 ( .A(n1722), .B(n1643), .C(n1642), .Z(acc_cmd1[19]) );
  COND1XL U1812 ( .A(n1722), .B(n1575), .C(n1574), .Z(acc_cmd1[36]) );
  COND1XL U1813 ( .A(n1722), .B(n1679), .C(n1678), .Z(acc_cmd1[10]) );
  COND1XL U1814 ( .A(n1722), .B(n1659), .C(n1658), .Z(acc_cmd1[15]) );
  COND1XL U1815 ( .A(n1722), .B(n1611), .C(n1610), .Z(acc_cmd1[27]) );
  COND1XL U1816 ( .A(n1722), .B(n1599), .C(n1598), .Z(acc_cmd1[30]) );
  COND1XL U1817 ( .A(n1722), .B(n1683), .C(n1682), .Z(acc_cmd1[9]) );
  COND1XL U1818 ( .A(n1722), .B(n1667), .C(n1666), .Z(acc_cmd1[13]) );
  COND1XL U1819 ( .A(n1722), .B(n1571), .C(n1570), .Z(acc_cmd1[37]) );
  COND1XL U1820 ( .A(n1722), .B(n1695), .C(n1694), .Z(acc_cmd1[6]) );
  COND1XL U1821 ( .A(n1722), .B(n1691), .C(n1690), .Z(acc_cmd1[7]) );
  COND1XL U1822 ( .A(n1722), .B(n1687), .C(n1686), .Z(acc_cmd1[8]) );
  COND1XL U1823 ( .A(n1722), .B(n1699), .C(n1698), .Z(acc_cmd1[5]) );
  COND1XL U1824 ( .A(n1722), .B(n1591), .C(n1590), .Z(acc_cmd1[32]) );
  COND1XL U1825 ( .A(n1722), .B(n1707), .C(n1706), .Z(acc_cmd1[3]) );
  COND1XL U1826 ( .A(n1722), .B(n1715), .C(n1714), .Z(acc_cmd1[1]) );
  COAN1X1 U1827 ( .A(n1269), .B(n1846), .C(n1845), .Z(n1175) );
  COAN1X1 U1828 ( .A(n1269), .B(n1848), .C(n1847), .Z(n1176) );
  COAN1X1 U1829 ( .A(n1269), .B(n1826), .C(n1825), .Z(n1177) );
  COAN1X1 U1830 ( .A(n1269), .B(n1828), .C(n1827), .Z(n1178) );
  COAN1X1 U1831 ( .A(n1269), .B(n1830), .C(n1829), .Z(n1179) );
  COAN1X1 U1832 ( .A(n1269), .B(n1832), .C(n1831), .Z(n1180) );
  COAN1X1 U1833 ( .A(n1269), .B(n1834), .C(n1833), .Z(n1181) );
  COAN1X1 U1834 ( .A(n1269), .B(n1836), .C(n1835), .Z(n1182) );
  COAN1X1 U1835 ( .A(n1269), .B(n1838), .C(n1837), .Z(n1183) );
  COAN1X1 U1836 ( .A(n1269), .B(n1840), .C(n1839), .Z(n1184) );
  COAN1X1 U1837 ( .A(n1265), .B(n1736), .C(n1735), .Z(n1185) );
  COAN1X1 U1838 ( .A(n1268), .B(n1810), .C(n1809), .Z(n1186) );
  COAN1X1 U1839 ( .A(n1268), .B(n1808), .C(n1807), .Z(n1187) );
  COAN1X1 U1840 ( .A(n1268), .B(n1804), .C(n1803), .Z(n1188) );
  COAN1X1 U1841 ( .A(n1268), .B(n1806), .C(n1805), .Z(n1189) );
  COAN1X1 U1842 ( .A(n1268), .B(n1802), .C(n1801), .Z(n1190) );
  COAN1X1 U1843 ( .A(n1267), .B(n1800), .C(n1799), .Z(n1191) );
  COAN1X1 U1844 ( .A(n1267), .B(n1796), .C(n1795), .Z(n1192) );
  COAN1X1 U1845 ( .A(n1267), .B(n1798), .C(n1797), .Z(n1193) );
  COAN1X1 U1846 ( .A(n1268), .B(n1824), .C(n1823), .Z(n1194) );
  COAN1X1 U1847 ( .A(n1268), .B(n1820), .C(n1819), .Z(n1195) );
  COAN1X1 U1848 ( .A(n1268), .B(n1822), .C(n1821), .Z(n1196) );
  COAN1X1 U1849 ( .A(n1268), .B(n1812), .C(n1811), .Z(n1197) );
  COAN1X1 U1850 ( .A(n1268), .B(n1814), .C(n1813), .Z(n1198) );
  COAN1X1 U1851 ( .A(n1268), .B(n1818), .C(n1817), .Z(n1199) );
  COAN1X1 U1852 ( .A(n1268), .B(n1816), .C(n1815), .Z(n1200) );
  COAN1X1 U1853 ( .A(n1267), .B(n1794), .C(n1793), .Z(n1201) );
  COAN1X1 U1854 ( .A(n1267), .B(n1792), .C(n1791), .Z(n1202) );
  COAN1X1 U1855 ( .A(n1267), .B(n1788), .C(n1787), .Z(n1203) );
  COAN1X1 U1856 ( .A(n1267), .B(n1790), .C(n1789), .Z(n1204) );
  COAN1X1 U1857 ( .A(n1267), .B(n1786), .C(n1785), .Z(n1205) );
  COAN1X1 U1858 ( .A(n1267), .B(n1784), .C(n1783), .Z(n1206) );
  COAN1X1 U1859 ( .A(n1267), .B(n1780), .C(n1779), .Z(n1207) );
  COAN1X1 U1860 ( .A(n1267), .B(n1782), .C(n1781), .Z(n1208) );
  COAN1X1 U1861 ( .A(n1267), .B(n1778), .C(n1777), .Z(n1209) );
  COAN1X1 U1862 ( .A(n1266), .B(n1776), .C(n1775), .Z(n1210) );
  COAN1X1 U1863 ( .A(n1266), .B(n1772), .C(n1771), .Z(n1211) );
  COAN1X1 U1864 ( .A(n1266), .B(n1774), .C(n1773), .Z(n1212) );
  COAN1X1 U1865 ( .A(n1266), .B(n1770), .C(n1769), .Z(n1213) );
  COAN1X1 U1866 ( .A(n1266), .B(n1768), .C(n1767), .Z(n1214) );
  COAN1X1 U1867 ( .A(n1266), .B(n1764), .C(n1763), .Z(n1215) );
  COAN1X1 U1868 ( .A(n1266), .B(n1766), .C(n1765), .Z(n1216) );
  COAN1X1 U1869 ( .A(n1266), .B(n1762), .C(n1761), .Z(n1217) );
  COAN1X1 U1870 ( .A(n1266), .B(n1760), .C(n1759), .Z(n1218) );
  COAN1X1 U1871 ( .A(n1266), .B(n1756), .C(n1755), .Z(n1219) );
  COAN1X1 U1872 ( .A(n1266), .B(n1758), .C(n1757), .Z(n1220) );
  COAN1X1 U1873 ( .A(n1266), .B(n1754), .C(n1753), .Z(n1221) );
  COAN1X1 U1874 ( .A(n1265), .B(n1752), .C(n1751), .Z(n1222) );
  COAN1X1 U1875 ( .A(n1265), .B(n1748), .C(n1747), .Z(n1223) );
  COAN1X1 U1876 ( .A(n1265), .B(n1750), .C(n1749), .Z(n1224) );
  COAN1X1 U1877 ( .A(n1265), .B(n1746), .C(n1745), .Z(n1225) );
  COAN1X1 U1878 ( .A(n1265), .B(n1744), .C(n1743), .Z(n1226) );
  COAN1X1 U1879 ( .A(n1265), .B(n1740), .C(n1739), .Z(n1227) );
  COAN1X1 U1880 ( .A(n1265), .B(n1742), .C(n1741), .Z(n1228) );
  COAN1X1 U1881 ( .A(n1265), .B(n1738), .C(n1737), .Z(n1229) );
  COAN1X1 U1882 ( .A(n1265), .B(n1734), .C(n1733), .Z(n1230) );
  COND1XL U1883 ( .A(n1270), .B(n1854), .C(n1853), .Z(acc_cmd2[62]) );
  COND1XL U1884 ( .A(n1270), .B(n1852), .C(n1851), .Z(acc_cmd2[59]) );
  COND1XL U1885 ( .A(n1270), .B(n1858), .C(n1857), .Z(acc_cmd2[61]) );
  COND1XL U1886 ( .A(n1270), .B(n1850), .C(n1849), .Z(acc_cmd2[60]) );
  COND1XL U1887 ( .A(n1269), .B(n1842), .C(n1841), .Z(acc_cmd2[58]) );
  CMX2X1 U1888 ( .A0(n1231), .A1(roundit), .S(n1232), .Z(n611) );
  CND2X1 U1889 ( .A(n1254), .B(n1317), .Z(n1232) );
  COND1XL U1890 ( .A(n1253), .B(n1405), .C(n1404), .Z(n583) );
  COND1XL U1891 ( .A(n1252), .B(n1407), .C(n1406), .Z(n584) );
  COND1XL U1892 ( .A(n1254), .B(n1409), .C(n1408), .Z(n585) );
  COND1XL U1893 ( .A(n1255), .B(n1411), .C(n1410), .Z(n586) );
  COND1XL U1894 ( .A(n1254), .B(n1413), .C(n1412), .Z(n587) );
  COND1XL U1895 ( .A(n1253), .B(n1415), .C(n1414), .Z(n588) );
  COND1XL U1896 ( .A(n1255), .B(n1417), .C(n1416), .Z(n589) );
  COND1XL U1897 ( .A(n1252), .B(n1419), .C(n1418), .Z(n590) );
  COND1XL U1898 ( .A(n1255), .B(n1421), .C(n1420), .Z(n591) );
  COND1XL U1899 ( .A(n1254), .B(n1423), .C(n1422), .Z(n592) );
  COND1XL U1900 ( .A(n1253), .B(n1459), .C(n1458), .Z(n610) );
  COND1XL U1901 ( .A(n1252), .B(n1457), .C(n1456), .Z(n609) );
  COND1XL U1902 ( .A(n1255), .B(n1453), .C(n1452), .Z(n607) );
  COND1XL U1903 ( .A(n1254), .B(n1455), .C(n1454), .Z(n608) );
  COND1XL U1904 ( .A(n1252), .B(n1397), .C(n1396), .Z(n579) );
  COND1XL U1905 ( .A(n1254), .B(n1445), .C(n1444), .Z(n603) );
  COND1XL U1906 ( .A(n1253), .B(n1447), .C(n1446), .Z(n604) );
  COND1XL U1907 ( .A(n1255), .B(n1449), .C(n1448), .Z(n605) );
  COND1XL U1908 ( .A(n1252), .B(n1451), .C(n1450), .Z(n606) );
  COND1XL U1909 ( .A(n1255), .B(n1443), .C(n1442), .Z(n602) );
  COND1XL U1910 ( .A(n1255), .B(n1399), .C(n1398), .Z(n580) );
  COND1XL U1911 ( .A(n1253), .B(n1401), .C(n1400), .Z(n581) );
  COND1XL U1912 ( .A(n1254), .B(n1403), .C(n1402), .Z(n582) );
  COND1XL U1913 ( .A(n1253), .B(n1427), .C(n1426), .Z(n594) );
  COND1XL U1914 ( .A(n1254), .B(n1441), .C(n1440), .Z(n601) );
  COND1XL U1915 ( .A(n1252), .B(n1425), .C(n1424), .Z(n593) );
  COND1XL U1916 ( .A(n1253), .B(n1437), .C(n1436), .Z(n599) );
  COND1XL U1917 ( .A(n1252), .B(n1439), .C(n1438), .Z(n600) );
  COND1XL U1918 ( .A(n1252), .B(n1429), .C(n1428), .Z(n595) );
  COND1XL U1919 ( .A(n1255), .B(n1431), .C(n1430), .Z(n596) );
  COND1XL U1920 ( .A(n1253), .B(n1433), .C(n1432), .Z(n597) );
  COND1XL U1921 ( .A(n1254), .B(n1435), .C(n1434), .Z(n598) );
  CNIVX1 U1922 ( .A(pushin), .Z(n1344) );
  CND3XL U1923 ( .A(en1_p2_d1), .B(n1255), .C(n1727), .Z(n1728) );
  CNR3XL U1924 ( .A(n1948), .B(n1251), .C(n1250), .Z(N404) );
  CNR3XL U1925 ( .A(n1947), .B(n1251), .C(n1250), .Z(N403) );
  CNR3XL U1926 ( .A(n1946), .B(n1251), .C(n1250), .Z(N402) );
  CNR3XL U1927 ( .A(n1943), .B(n1251), .C(n1250), .Z(N399) );
  CNR3XL U1928 ( .A(n1944), .B(n1251), .C(n1250), .Z(N400) );
  CAN2X1 U1929 ( .A(n1466), .B(push0_p2), .Z(n1233) );
  CAN2X1 U1930 ( .A(n12), .B(push0_p2), .Z(n1234) );
  CAN2X1 U1931 ( .A(n1467), .B(push0_p2), .Z(n1235) );
  CNIVXL U1932 ( .A(en2_p2), .Z(n1252) );
  CNIVX1 U1933 ( .A(en0_p2), .Z(n1256) );
  CNIVXL U1934 ( .A(en1_p2), .Z(n1261) );
  CNIVXL U1935 ( .A(en1_p2), .Z(n1262) );
  CNIVXL U1936 ( .A(en1_p2), .Z(n1263) );
  CNIVX1 U1937 ( .A(en0_p2), .Z(n1257) );
  CNIVX1 U1938 ( .A(en0_p2), .Z(n1258) );
  CNIVX1 U1939 ( .A(en0_p2), .Z(n1259) );
  CNIVX1 U1940 ( .A(h0_p1[2]), .Z(n1239) );
  CNIVX1 U1941 ( .A(h0_p1[2]), .Z(n1242) );
  CNIVX1 U1942 ( .A(h0_p1[2]), .Z(n1241) );
  CNIVX1 U1943 ( .A(h0_p1[2]), .Z(n1240) );
  CNIVX1 U1944 ( .A(h0_p1[2]), .Z(n1243) );
  CNIVX1 U1945 ( .A(h0_p1[4]), .Z(n1249) );
  CNIVX1 U1946 ( .A(h0_p1[4]), .Z(n1248) );
  CNIVX1 U1947 ( .A(h0_p1[4]), .Z(n1245) );
  CNIVX1 U1948 ( .A(h0_p1[4]), .Z(n1247) );
  CNIVX1 U1949 ( .A(h0_p1[4]), .Z(n1246) );
  CNIVX1 U1950 ( .A(h0_p1[4]), .Z(n1244) );
  CNIVX1 U1951 ( .A(pushin), .Z(n1343) );
  CNIVX1 U1952 ( .A(pushin), .Z(n1342) );
  CNIVXL U1953 ( .A(en2_p2), .Z(n1254) );
  CNIVX1 U1954 ( .A(pushin), .Z(n1340) );
  CNIVX1 U1955 ( .A(pushin), .Z(n1341) );
  CNIVX1 U1956 ( .A(pushin), .Z(n1339) );
  CNR2X1 U1957 ( .A(cmd0_p2[0]), .B(cmd0_p2[1]), .Z(n12) );
  CNIVX1 U1958 ( .A(h0_p1[5]), .Z(n1250) );
  CNIVX1 U1959 ( .A(h0_p1[6]), .Z(n1251) );
  CNR3XL U1960 ( .A(n1941), .B(cmd0[1]), .C(cmd0[0]), .Z(en0_p0) );
  CNIVX4 U1961 ( .A(q0[14]), .Z(n1236) );
  CMX2XL U1962 ( .A0(n1162), .A1(q[19]), .S(n1340), .Z(n677) );
  CMX2XL U1963 ( .A0(n1172), .A1(q[5]), .S(n1341), .Z(n663) );
  CMX2XL U1964 ( .A0(n1166), .A1(q[15]), .S(n1340), .Z(n673) );
  CMX2XL U1965 ( .A0(n1167), .A1(q[3]), .S(n1341), .Z(n661) );
  CMX2XL U1966 ( .A0(n1169), .A1(q[23]), .S(n1339), .Z(n681) );
  CMX2XL U1967 ( .A0(n1170), .A1(q[7]), .S(n1341), .Z(n665) );
  CMX2XL U1968 ( .A0(n1161), .A1(q[21]), .S(n1339), .Z(n679) );
  CMX2XL U1969 ( .A0(n1158), .A1(q[29]), .S(n1339), .Z(n687) );
  CMX2XL U1970 ( .A0(n1237), .A1(q[27]), .S(n1339), .Z(n685) );
  CMX2XL U1971 ( .A0(n1163), .A1(q[1]), .S(n1341), .Z(n659) );
  CMX2XL U1972 ( .A0(n1173), .A1(q[13]), .S(n1340), .Z(n671) );
  CNIVX4 U1973 ( .A(en1_p2), .Z(n1260) );
  CIVXL U1974 ( .A(n1324), .Z(n1323) );
  CIVX1 U1975 ( .A(h0_p1[0]), .Z(n1324) );
  CIVXL U1976 ( .A(n1331), .Z(n1330) );
  CIVX2 U1977 ( .A(h0_p1[1]), .Z(n1331) );
  CIVX2 U1978 ( .A(h0_p1[3]), .Z(n1337) );
  CIVXL U1979 ( .A(n1128), .Z(n1338) );
  CMX2X1 U1980 ( .A0(q0[30]), .A1(q[30]), .S(n1339), .Z(n688) );
  CMX2X1 U1981 ( .A0(q0[26]), .A1(q[26]), .S(n1339), .Z(n684) );
  CMX2X1 U1982 ( .A0(q0[24]), .A1(q[24]), .S(n1339), .Z(n682) );
  CMX2X1 U1983 ( .A0(q0[22]), .A1(q[22]), .S(n1339), .Z(n680) );
  CMX2X1 U1984 ( .A0(q0[12]), .A1(q[12]), .S(n1340), .Z(n670) );
  CMX2X1 U1985 ( .A0(q0[8]), .A1(q[8]), .S(n1340), .Z(n666) );
  CMX2X1 U1986 ( .A0(n1171), .A1(q[6]), .S(n1341), .Z(n664) );
  CMX2X1 U1987 ( .A0(q0[4]), .A1(q[4]), .S(n1341), .Z(n662) );
  CMX2X1 U1988 ( .A0(q0[2]), .A1(q[2]), .S(n1341), .Z(n660) );
  CMX2X1 U1989 ( .A0(q0[0]), .A1(q[0]), .S(n1341), .Z(n658) );
  CMX2X1 U1990 ( .A0(h0[31]), .A1(h[31]), .S(n1341), .Z(n657) );
  CMX2X1 U1991 ( .A0(h0[30]), .A1(h[30]), .S(n1341), .Z(n656) );
  CMX2X1 U1992 ( .A0(h0[29]), .A1(h[29]), .S(n1341), .Z(n655) );
  CMX2X1 U1993 ( .A0(h0[28]), .A1(h[28]), .S(n1341), .Z(n654) );
  CMX2X1 U1994 ( .A0(h0[27]), .A1(h[27]), .S(n1342), .Z(n653) );
  CMX2X1 U1995 ( .A0(h0[26]), .A1(h[26]), .S(n1342), .Z(n652) );
  CMX2X1 U1996 ( .A0(h0[24]), .A1(h[24]), .S(n1342), .Z(n650) );
  CMX2X1 U1997 ( .A0(h0[23]), .A1(h[23]), .S(n1342), .Z(n649) );
  CMX2X1 U1998 ( .A0(h0[22]), .A1(h[22]), .S(n1342), .Z(n648) );
  CMX2X1 U1999 ( .A0(h0[21]), .A1(h[21]), .S(n1342), .Z(n647) );
  CMX2X1 U2000 ( .A0(h0[20]), .A1(h[20]), .S(n1342), .Z(n646) );
  CMX2X1 U2001 ( .A0(h0[19]), .A1(h[19]), .S(n1342), .Z(n645) );
  CMX2X1 U2002 ( .A0(h0[17]), .A1(h[17]), .S(n1342), .Z(n643) );
  CMX2X1 U2003 ( .A0(h0[15]), .A1(h[15]), .S(n1343), .Z(n641) );
  CMX2X1 U2004 ( .A0(h0[14]), .A1(h[14]), .S(n1343), .Z(n640) );
  CMX2X1 U2005 ( .A0(h0[10]), .A1(h[10]), .S(n1343), .Z(n636) );
  CMX2X1 U2006 ( .A0(h0[9]), .A1(h[9]), .S(n1343), .Z(n635) );
  CMX2X1 U2007 ( .A0(h0[7]), .A1(h[7]), .S(n1343), .Z(n633) );
  CMX2X1 U2008 ( .A0(h0[3]), .A1(h[3]), .S(n1344), .Z(n623) );
  CMX2X1 U2009 ( .A0(n1128), .A1(h[0]), .S(n1344), .Z(n614) );
  CMX2X1 U2010 ( .A0(out2_p2[63]), .A1(N405), .S(n1252), .Z(n547) );
  CMX2X1 U2011 ( .A0(out2_p2[62]), .A1(N404), .S(n1255), .Z(n548) );
  CMX2X1 U2012 ( .A0(out2_p2[61]), .A1(N403), .S(n1254), .Z(n549) );
  CMX2X1 U2013 ( .A0(out2_p2[60]), .A1(N402), .S(n1252), .Z(n550) );
  CMX2X1 U2014 ( .A0(out2_p2[59]), .A1(N401), .S(n1253), .Z(n551) );
  CMX2X1 U2015 ( .A0(out2_p2[58]), .A1(N400), .S(n1252), .Z(n552) );
  CMX2X1 U2016 ( .A0(out2_p2[57]), .A1(N399), .S(n1255), .Z(n553) );
  CMX2X1 U2017 ( .A0(out2_p2[56]), .A1(N398), .S(n1253), .Z(n554) );
  CIVX2 U2018 ( .A(n1251), .Z(n1394) );
  CIVX2 U2019 ( .A(n1250), .Z(n1345) );
  CIVX2 U2020 ( .A(n2232), .Z(n1347) );
  COND2X1 U2021 ( .A(n1238), .B(n1347), .C(n1253), .D(n1346), .Z(n555) );
  CIVX2 U2022 ( .A(n2231), .Z(n1349) );
  COND2X1 U2023 ( .A(n1238), .B(n1349), .C(n1254), .D(n1348), .Z(n556) );
  CIVX2 U2024 ( .A(n2230), .Z(n1351) );
  COND2X1 U2025 ( .A(n1395), .B(n1351), .C(n1253), .D(n1350), .Z(n557) );
  CIVX2 U2026 ( .A(n2229), .Z(n1353) );
  COND2X1 U2027 ( .A(n1238), .B(n1353), .C(n1252), .D(n1352), .Z(n558) );
  CIVX2 U2028 ( .A(n2228), .Z(n1355) );
  COND2X1 U2029 ( .A(n1395), .B(n1355), .C(n1254), .D(n1354), .Z(n559) );
  CIVX2 U2030 ( .A(n2227), .Z(n1357) );
  COND2X1 U2031 ( .A(n1238), .B(n1357), .C(n1255), .D(n1356), .Z(n560) );
  CIVX2 U2032 ( .A(n2226), .Z(n1359) );
  COND2X1 U2033 ( .A(n1395), .B(n1359), .C(n1254), .D(n1358), .Z(n561) );
  CIVX2 U2034 ( .A(n2217), .Z(n1361) );
  COND2X1 U2035 ( .A(n1238), .B(n1361), .C(n1253), .D(n1360), .Z(n562) );
  CIVX2 U2036 ( .A(n2216), .Z(n1363) );
  COND2X1 U2037 ( .A(n1395), .B(n1363), .C(n1255), .D(n1362), .Z(n563) );
  CIVX2 U2038 ( .A(n2215), .Z(n1365) );
  COND2X1 U2039 ( .A(n1238), .B(n1365), .C(n1252), .D(n1364), .Z(n564) );
  CIVX2 U2040 ( .A(n2214), .Z(n1367) );
  COND2X1 U2041 ( .A(n1395), .B(n1367), .C(n1255), .D(n1366), .Z(n565) );
  CIVX2 U2042 ( .A(n2213), .Z(n1369) );
  COND2X1 U2043 ( .A(n1238), .B(n1369), .C(n1254), .D(n1368), .Z(n566) );
  CIVX2 U2044 ( .A(n2212), .Z(n1371) );
  COND2X1 U2045 ( .A(n1395), .B(n1371), .C(n1252), .D(n1370), .Z(n567) );
  CIVX2 U2046 ( .A(n2211), .Z(n1373) );
  COND2X1 U2047 ( .A(n1238), .B(n1373), .C(n1253), .D(n1372), .Z(n568) );
  CIVX2 U2048 ( .A(n2210), .Z(n1375) );
  COND2X1 U2049 ( .A(n1395), .B(n1375), .C(n1252), .D(n1374), .Z(n569) );
  CIVX2 U2050 ( .A(n2275), .Z(n1377) );
  COND2X1 U2051 ( .A(n1238), .B(n1377), .C(n1255), .D(n1376), .Z(n570) );
  CIVX2 U2052 ( .A(n2269), .Z(n1379) );
  COND2X1 U2053 ( .A(n1395), .B(n1379), .C(n1253), .D(n1378), .Z(n571) );
  CIVX2 U2054 ( .A(n2263), .Z(n1381) );
  COND2X1 U2055 ( .A(n1238), .B(n1381), .C(n1254), .D(n1380), .Z(n572) );
  CIVX2 U2056 ( .A(n2255), .Z(n1383) );
  COND2X1 U2057 ( .A(n1395), .B(n1383), .C(n1253), .D(n1382), .Z(n573) );
  CIVX2 U2058 ( .A(n2242), .Z(n1385) );
  COND2X1 U2059 ( .A(n1238), .B(n1385), .C(n1252), .D(n1384), .Z(n574) );
  CIVX2 U2060 ( .A(n2224), .Z(n1387) );
  COND2X1 U2061 ( .A(n1395), .B(n1387), .C(n1254), .D(n1386), .Z(n575) );
  CIVX2 U2062 ( .A(n2204), .Z(n1389) );
  COND2X1 U2063 ( .A(n1238), .B(n1389), .C(n1255), .D(n1388), .Z(n576) );
  CIVX2 U2064 ( .A(n2184), .Z(n1391) );
  COND2X1 U2065 ( .A(n1395), .B(n1391), .C(n1254), .D(n1390), .Z(n577) );
  CIVX2 U2066 ( .A(n2183), .Z(n1393) );
  COND2X1 U2067 ( .A(n1393), .B(n1238), .C(n1253), .D(n1392), .Z(n578) );
  CANR2X1 U2068 ( .A(n2247), .B(n1174), .C(n2180), .D(n1264), .Z(n1398) );
  CANR2X1 U2069 ( .A(n2246), .B(n1174), .C(n2176), .D(n1264), .Z(n1400) );
  CANR2X1 U2070 ( .A(n2245), .B(n1174), .C(n2160), .D(n1264), .Z(n1402) );
  CANR2X1 U2071 ( .A(n2244), .B(n1174), .C(n2156), .D(n1264), .Z(n1404) );
  CANR2X1 U2072 ( .A(n2235), .B(n1174), .C(n2152), .D(n1264), .Z(n1406) );
  CANR2X1 U2073 ( .A(n2234), .B(n1174), .C(n2148), .D(n1264), .Z(n1408) );
  CANR2X1 U2074 ( .A(n2233), .B(n1174), .C(n2144), .D(n1264), .Z(n1410) );
  CANR2X1 U2075 ( .A(n2232), .B(n1174), .C(n2138), .D(n1264), .Z(n1412) );
  CANR2X1 U2076 ( .A(n2231), .B(n1174), .C(n2131), .D(n1264), .Z(n1414) );
  CANR2X1 U2077 ( .A(n2230), .B(n1174), .C(n2124), .D(n1264), .Z(n1416) );
  CANR2X1 U2078 ( .A(n2229), .B(n1174), .C(n2117), .D(n1264), .Z(n1418) );
  CANR2X1 U2079 ( .A(n2228), .B(n1174), .C(n2110), .D(n1264), .Z(n1420) );
  CANR2X1 U2080 ( .A(n2227), .B(n1174), .C(n2093), .D(n1264), .Z(n1422) );
  CANR2X1 U2081 ( .A(n2226), .B(n1174), .C(n2086), .D(n1264), .Z(n1424) );
  CANR2X1 U2082 ( .A(n2217), .B(n1174), .C(n2079), .D(n1264), .Z(n1426) );
  CANR2X1 U2083 ( .A(n2216), .B(n1174), .C(n2066), .D(n1264), .Z(n1428) );
  CANR2X1 U2084 ( .A(n2215), .B(n1174), .C(n2061), .D(n1264), .Z(n1430) );
  CANR2X1 U2085 ( .A(n2214), .B(n1174), .C(n2046), .D(n1264), .Z(n1432) );
  CANR2X1 U2086 ( .A(n2213), .B(n1174), .C(n2031), .D(n1264), .Z(n1434) );
  CANR2X1 U2087 ( .A(n2212), .B(n1174), .C(n2003), .D(n1264), .Z(n1436) );
  CANR2X1 U2088 ( .A(n2211), .B(n1174), .C(n1987), .D(n1264), .Z(n1438) );
  CANR2X1 U2089 ( .A(n2210), .B(n1174), .C(n1985), .D(n1264), .Z(n1440) );
  CANR2X1 U2090 ( .A(n2275), .B(n1174), .C(n2276), .D(n1264), .Z(n1442) );
  CANR2X1 U2091 ( .A(n2269), .B(n1174), .C(n2270), .D(n1264), .Z(n1444) );
  CANR2X1 U2092 ( .A(n2263), .B(n1174), .C(n2264), .D(n1264), .Z(n1446) );
  CANR2X1 U2093 ( .A(n2255), .B(n1174), .C(n2256), .D(n1264), .Z(n1448) );
  CANR2X1 U2094 ( .A(n2242), .B(n1174), .C(n2243), .D(n1264), .Z(n1450) );
  CANR2X1 U2095 ( .A(n2224), .B(n1174), .C(n2225), .D(n1264), .Z(n1452) );
  CANR2X1 U2096 ( .A(n2204), .B(n1174), .C(n2205), .D(n1264), .Z(n1454) );
  CANR2X1 U2097 ( .A(n2184), .B(n1174), .C(n2172), .D(n1264), .Z(n1456) );
  CANR2X1 U2098 ( .A(n2183), .B(n1174), .C(n2103), .D(n1264), .Z(n1458) );
  CIVX2 U2099 ( .A(cmd0[1]), .Z(n1460) );
  CAN3X2 U2100 ( .A(n1070), .B(cmd0[0]), .C(n1460), .Z(en1_p0) );
  CIVX2 U2101 ( .A(en1_p2_d1), .Z(n1725) );
  CND2X1 U2102 ( .A(n1260), .B(n1725), .Z(n1461) );
  CIVX2 U2103 ( .A(en0_p2_d1), .Z(n1727) );
  CND2X1 U2104 ( .A(n1722), .B(n1727), .Z(n1462) );
  CND2X1 U2105 ( .A(n1722), .B(en0_p2_d1), .Z(n1463) );
  CMX2X1 U2106 ( .A0(out1_p2[62]), .A1(N270), .S(n1262), .Z(n421) );
  CIVX2 U2107 ( .A(cmd0_p2[0]), .Z(n1939) );
  CND2X1 U2108 ( .A(cmd0_p2[1]), .B(n1939), .Z(n1879) );
  CIVX2 U2109 ( .A(n1879), .Z(n1466) );
  CANR2X1 U2110 ( .A(n1234), .B(out0_p2[62]), .C(N480), .D(n1233), .Z(n1469)
         );
  CIVX2 U2111 ( .A(cmd0_p2[1]), .Z(n1938) );
  CND2X1 U2112 ( .A(cmd0_p2[0]), .B(n1938), .Z(n1878) );
  CIVX2 U2113 ( .A(n1878), .Z(n1467) );
  CANR2X1 U2114 ( .A(n1235), .B(out1_p2[62]), .C(acc[62]), .D(n1936), .Z(n1468) );
  CND2X1 U2115 ( .A(n1469), .B(n1468), .Z(n420) );
  CMX2X1 U2116 ( .A0(out1_p2[61]), .A1(N269), .S(n1263), .Z(n423) );
  CANR2X1 U2117 ( .A(n1234), .B(out0_p2[61]), .C(N479), .D(n1233), .Z(n1473)
         );
  CANR2X1 U2118 ( .A(n1235), .B(out1_p2[61]), .C(acc[61]), .D(n1936), .Z(n1472) );
  CND2X1 U2119 ( .A(n1473), .B(n1472), .Z(n422) );
  CMX2X1 U2120 ( .A0(out1_p2[60]), .A1(N268), .S(n1262), .Z(n425) );
  CANR2X1 U2121 ( .A(n1234), .B(out0_p2[60]), .C(N478), .D(n1233), .Z(n1477)
         );
  CANR2X1 U2122 ( .A(n1235), .B(out1_p2[60]), .C(acc[60]), .D(n1936), .Z(n1476) );
  CND2X1 U2123 ( .A(n1477), .B(n1476), .Z(n424) );
  CMX2X1 U2124 ( .A0(out1_p2[59]), .A1(N267), .S(n1261), .Z(n427) );
  CANR2X1 U2125 ( .A(n1234), .B(out0_p2[59]), .C(N477), .D(n1233), .Z(n1481)
         );
  CANR2X1 U2126 ( .A(n1235), .B(out1_p2[59]), .C(acc[59]), .D(n1936), .Z(n1480) );
  CND2X1 U2127 ( .A(n1481), .B(n1480), .Z(n426) );
  CMX2X1 U2128 ( .A0(out1_p2[58]), .A1(N266), .S(n1260), .Z(n429) );
  CANR2X1 U2129 ( .A(n1234), .B(out0_p2[58]), .C(N476), .D(n1233), .Z(n1485)
         );
  CANR2X1 U2130 ( .A(n1235), .B(out1_p2[58]), .C(acc[58]), .D(n1936), .Z(n1484) );
  CND2X1 U2131 ( .A(n1485), .B(n1484), .Z(n428) );
  CMX2X1 U2132 ( .A0(out1_p2[57]), .A1(N265), .S(n1261), .Z(n431) );
  CANR2X1 U2133 ( .A(n1234), .B(out0_p2[57]), .C(N475), .D(n1233), .Z(n1489)
         );
  CANR2X1 U2134 ( .A(n1235), .B(out1_p2[57]), .C(acc[57]), .D(n1936), .Z(n1488) );
  CND2X1 U2135 ( .A(n1489), .B(n1488), .Z(n430) );
  CMX2X1 U2136 ( .A0(out1_p2[56]), .A1(N264), .S(n1263), .Z(n433) );
  CANR2X1 U2137 ( .A(n1234), .B(out0_p2[56]), .C(N474), .D(n1233), .Z(n1493)
         );
  CANR2X1 U2138 ( .A(n1235), .B(out1_p2[56]), .C(acc[56]), .D(n1936), .Z(n1492) );
  CND2X1 U2139 ( .A(n1493), .B(n1492), .Z(n432) );
  CMX2X1 U2140 ( .A0(out1_p2[55]), .A1(N263), .S(n1262), .Z(n435) );
  CANR2X1 U2141 ( .A(n1234), .B(out0_p2[55]), .C(N473), .D(n1233), .Z(n1497)
         );
  CANR2X1 U2142 ( .A(n1235), .B(out1_p2[55]), .C(acc[55]), .D(n1936), .Z(n1496) );
  CND2X1 U2143 ( .A(n1497), .B(n1496), .Z(n434) );
  CMX2X1 U2144 ( .A0(out1_p2[54]), .A1(N262), .S(n1262), .Z(n437) );
  CANR2X1 U2145 ( .A(n1234), .B(out0_p2[54]), .C(N472), .D(n1233), .Z(n1501)
         );
  CANR2X1 U2146 ( .A(n1235), .B(out1_p2[54]), .C(acc[54]), .D(n1936), .Z(n1500) );
  CND2X1 U2147 ( .A(n1501), .B(n1500), .Z(n436) );
  CMX2X1 U2148 ( .A0(out1_p2[53]), .A1(N261), .S(n1263), .Z(n439) );
  CANR2X1 U2149 ( .A(n1234), .B(out0_p2[53]), .C(N471), .D(n1233), .Z(n1505)
         );
  CANR2X1 U2150 ( .A(n1235), .B(out1_p2[53]), .C(acc[53]), .D(n1936), .Z(n1504) );
  CND2X1 U2151 ( .A(n1505), .B(n1504), .Z(n438) );
  CMX2X1 U2152 ( .A0(out1_p2[52]), .A1(N260), .S(n1260), .Z(n441) );
  CANR2X1 U2153 ( .A(n1234), .B(out0_p2[52]), .C(N470), .D(n1233), .Z(n1509)
         );
  CANR2X1 U2154 ( .A(n1235), .B(out1_p2[52]), .C(acc[52]), .D(n1936), .Z(n1508) );
  CND2X1 U2155 ( .A(n1509), .B(n1508), .Z(n440) );
  CMX2X1 U2156 ( .A0(out1_p2[51]), .A1(N259), .S(n1263), .Z(n443) );
  CANR2X1 U2157 ( .A(n1234), .B(out0_p2[51]), .C(N469), .D(n1233), .Z(n1513)
         );
  CANR2X1 U2158 ( .A(n1235), .B(out1_p2[51]), .C(acc[51]), .D(n1936), .Z(n1512) );
  CND2X1 U2159 ( .A(n1513), .B(n1512), .Z(n442) );
  CMX2X1 U2160 ( .A0(out1_p2[50]), .A1(N258), .S(n1260), .Z(n445) );
  CANR2X1 U2161 ( .A(n1234), .B(out0_p2[50]), .C(N468), .D(n1233), .Z(n1517)
         );
  CANR2X1 U2162 ( .A(n1235), .B(out1_p2[50]), .C(acc[50]), .D(n1936), .Z(n1516) );
  CND2X1 U2163 ( .A(n1517), .B(n1516), .Z(n444) );
  CMX2X1 U2164 ( .A0(out1_p2[49]), .A1(N257), .S(n1261), .Z(n447) );
  CANR2X1 U2165 ( .A(n1234), .B(out0_p2[49]), .C(N467), .D(n1233), .Z(n1521)
         );
  CANR2X1 U2166 ( .A(n1235), .B(out1_p2[49]), .C(acc[49]), .D(n1936), .Z(n1520) );
  CND2X1 U2167 ( .A(n1521), .B(n1520), .Z(n446) );
  CMX2X1 U2168 ( .A0(out1_p2[48]), .A1(N256), .S(n1261), .Z(n449) );
  CANR2X1 U2169 ( .A(n1234), .B(out0_p2[48]), .C(N466), .D(n1233), .Z(n1525)
         );
  CANR2X1 U2170 ( .A(n1235), .B(out1_p2[48]), .C(acc[48]), .D(n1936), .Z(n1524) );
  CND2X1 U2171 ( .A(n1525), .B(n1524), .Z(n448) );
  CMX2X1 U2172 ( .A0(out1_p2[47]), .A1(N255), .S(n1260), .Z(n451) );
  CANR2X1 U2173 ( .A(n1234), .B(out0_p2[47]), .C(N465), .D(n1233), .Z(n1529)
         );
  CANR2X1 U2174 ( .A(n1235), .B(out1_p2[47]), .C(acc[47]), .D(n1936), .Z(n1528) );
  CND2X1 U2175 ( .A(n1529), .B(n1528), .Z(n450) );
  CMX2X1 U2176 ( .A0(out1_p2[46]), .A1(N254), .S(n1262), .Z(n453) );
  CANR2X1 U2177 ( .A(n1234), .B(out0_p2[46]), .C(N464), .D(n1233), .Z(n1533)
         );
  CANR2X1 U2178 ( .A(n1235), .B(out1_p2[46]), .C(acc[46]), .D(n1936), .Z(n1532) );
  CND2X1 U2179 ( .A(n1533), .B(n1532), .Z(n452) );
  CMX2X1 U2180 ( .A0(out1_p2[45]), .A1(N253), .S(n1263), .Z(n455) );
  CANR2X1 U2181 ( .A(n1234), .B(out0_p2[45]), .C(N463), .D(n1233), .Z(n1537)
         );
  CANR2X1 U2182 ( .A(n1235), .B(out1_p2[45]), .C(acc[45]), .D(n1936), .Z(n1536) );
  CND2X1 U2183 ( .A(n1537), .B(n1536), .Z(n454) );
  CMX2X1 U2184 ( .A0(out1_p2[44]), .A1(N252), .S(n1262), .Z(n457) );
  CANR2X1 U2185 ( .A(n1234), .B(out0_p2[44]), .C(N462), .D(n1233), .Z(n1541)
         );
  CANR2X1 U2186 ( .A(n1235), .B(out1_p2[44]), .C(acc[44]), .D(n1936), .Z(n1540) );
  CND2X1 U2187 ( .A(n1541), .B(n1540), .Z(n456) );
  CMX2X1 U2188 ( .A0(out1_p2[43]), .A1(N251), .S(n1261), .Z(n459) );
  CANR2X1 U2189 ( .A(n1234), .B(out0_p2[43]), .C(N461), .D(n1233), .Z(n1545)
         );
  CANR2X1 U2190 ( .A(n1235), .B(out1_p2[43]), .C(acc[43]), .D(n1936), .Z(n1544) );
  CND2X1 U2191 ( .A(n1545), .B(n1544), .Z(n458) );
  CMX2X1 U2192 ( .A0(out1_p2[42]), .A1(N250), .S(n1260), .Z(n461) );
  CANR2X1 U2193 ( .A(n1234), .B(out0_p2[42]), .C(N460), .D(n1233), .Z(n1549)
         );
  CANR2X1 U2194 ( .A(n1235), .B(out1_p2[42]), .C(acc[42]), .D(n1936), .Z(n1548) );
  CND2X1 U2195 ( .A(n1549), .B(n1548), .Z(n460) );
  CMX2X1 U2196 ( .A0(out1_p2[41]), .A1(N249), .S(n1261), .Z(n463) );
  CANR2X1 U2197 ( .A(n1234), .B(out0_p2[41]), .C(N459), .D(n1233), .Z(n1553)
         );
  CANR2X1 U2198 ( .A(n1235), .B(out1_p2[41]), .C(acc[41]), .D(n1936), .Z(n1552) );
  CND2X1 U2199 ( .A(n1553), .B(n1552), .Z(n462) );
  CMX2X1 U2200 ( .A0(out1_p2[40]), .A1(N248), .S(n1263), .Z(n465) );
  CANR2X1 U2201 ( .A(n1234), .B(out0_p2[40]), .C(N458), .D(n1233), .Z(n1557)
         );
  CANR2X1 U2202 ( .A(n1235), .B(out1_p2[40]), .C(acc[40]), .D(n1936), .Z(n1556) );
  CND2X1 U2203 ( .A(n1557), .B(n1556), .Z(n464) );
  CMX2X1 U2204 ( .A0(out1_p2[39]), .A1(N247), .S(n1262), .Z(n467) );
  CANR2X1 U2205 ( .A(n1234), .B(out0_p2[39]), .C(N457), .D(n1233), .Z(n1561)
         );
  CANR2X1 U2206 ( .A(n1235), .B(out1_p2[39]), .C(acc[39]), .D(n1936), .Z(n1560) );
  CND2X1 U2207 ( .A(n1561), .B(n1560), .Z(n466) );
  CMX2X1 U2208 ( .A0(out1_p2[38]), .A1(N246), .S(n1262), .Z(n469) );
  CANR2X1 U2209 ( .A(n1234), .B(out0_p2[38]), .C(N456), .D(n1233), .Z(n1565)
         );
  CANR2X1 U2210 ( .A(n1235), .B(out1_p2[38]), .C(acc[38]), .D(n1936), .Z(n1564) );
  CND2X1 U2211 ( .A(n1565), .B(n1564), .Z(n468) );
  CMX2X1 U2212 ( .A0(out1_p2[37]), .A1(N245), .S(n1263), .Z(n471) );
  CANR2X1 U2213 ( .A(n1234), .B(out0_p2[37]), .C(N455), .D(n1233), .Z(n1569)
         );
  CANR2X1 U2214 ( .A(n1235), .B(out1_p2[37]), .C(acc[37]), .D(n1936), .Z(n1568) );
  CND2X1 U2215 ( .A(n1569), .B(n1568), .Z(n470) );
  CMX2X1 U2216 ( .A0(out1_p2[36]), .A1(N244), .S(n1260), .Z(n473) );
  CANR2X1 U2217 ( .A(n1234), .B(out0_p2[36]), .C(N454), .D(n1233), .Z(n1573)
         );
  CANR2X1 U2218 ( .A(n1235), .B(out1_p2[36]), .C(acc[36]), .D(n1936), .Z(n1572) );
  CND2X1 U2219 ( .A(n1573), .B(n1572), .Z(n472) );
  CMX2X1 U2220 ( .A0(out1_p2[35]), .A1(N243), .S(n1263), .Z(n475) );
  CANR2X1 U2221 ( .A(n1234), .B(out0_p2[35]), .C(N453), .D(n1233), .Z(n1577)
         );
  CANR2X1 U2222 ( .A(n1235), .B(out1_p2[35]), .C(acc[35]), .D(n1936), .Z(n1576) );
  CND2X1 U2223 ( .A(n1577), .B(n1576), .Z(n474) );
  CMX2X1 U2224 ( .A0(out1_p2[34]), .A1(N242), .S(n1260), .Z(n477) );
  CANR2X1 U2225 ( .A(n1234), .B(out0_p2[34]), .C(N452), .D(n1233), .Z(n1581)
         );
  CANR2X1 U2226 ( .A(n1235), .B(out1_p2[34]), .C(acc[34]), .D(n1936), .Z(n1580) );
  CND2X1 U2227 ( .A(n1581), .B(n1580), .Z(n476) );
  CMX2X1 U2228 ( .A0(out1_p2[33]), .A1(N241), .S(n1261), .Z(n479) );
  CANR2X1 U2229 ( .A(n1234), .B(out0_p2[33]), .C(N451), .D(n1233), .Z(n1585)
         );
  CANR2X1 U2230 ( .A(n1235), .B(out1_p2[33]), .C(acc[33]), .D(n1936), .Z(n1584) );
  CND2X1 U2231 ( .A(n1585), .B(n1584), .Z(n478) );
  CMX2X1 U2232 ( .A0(out1_p2[32]), .A1(N240), .S(n1261), .Z(n481) );
  CANR2X1 U2233 ( .A(n1234), .B(out0_p2[32]), .C(N450), .D(n1233), .Z(n1589)
         );
  CANR2X1 U2234 ( .A(n1235), .B(out1_p2[32]), .C(acc[32]), .D(n1936), .Z(n1588) );
  CND2X1 U2235 ( .A(n1589), .B(n1588), .Z(n480) );
  CMX2X1 U2236 ( .A0(out1_p2[31]), .A1(N239), .S(n1260), .Z(n483) );
  CANR2X1 U2237 ( .A(n1234), .B(out0_p2[31]), .C(N449), .D(n1233), .Z(n1593)
         );
  CANR2X1 U2238 ( .A(n1235), .B(out1_p2[31]), .C(acc[31]), .D(n1936), .Z(n1592) );
  CND2X1 U2239 ( .A(n1593), .B(n1592), .Z(n482) );
  CMX2X1 U2240 ( .A0(out1_p2[30]), .A1(N238), .S(n1262), .Z(n485) );
  CANR2X1 U2241 ( .A(n1234), .B(out0_p2[30]), .C(N448), .D(n1233), .Z(n1597)
         );
  CANR2X1 U2242 ( .A(n1235), .B(out1_p2[30]), .C(acc[30]), .D(n1936), .Z(n1596) );
  CND2X1 U2243 ( .A(n1597), .B(n1596), .Z(n484) );
  CMX2X1 U2244 ( .A0(out1_p2[29]), .A1(N237), .S(n1263), .Z(n487) );
  CANR2X1 U2245 ( .A(n1234), .B(out0_p2[29]), .C(N447), .D(n1233), .Z(n1601)
         );
  CANR2X1 U2246 ( .A(n1235), .B(out1_p2[29]), .C(acc[29]), .D(n1936), .Z(n1600) );
  CND2X1 U2247 ( .A(n1601), .B(n1600), .Z(n486) );
  CMX2X1 U2248 ( .A0(out1_p2[28]), .A1(N236), .S(n1262), .Z(n489) );
  CANR2X1 U2249 ( .A(n1234), .B(out0_p2[28]), .C(N446), .D(n1233), .Z(n1605)
         );
  CANR2X1 U2250 ( .A(n1235), .B(out1_p2[28]), .C(acc[28]), .D(n1936), .Z(n1604) );
  CND2X1 U2251 ( .A(n1605), .B(n1604), .Z(n488) );
  CMX2X1 U2252 ( .A0(out1_p2[27]), .A1(N235), .S(n1261), .Z(n491) );
  CANR2X1 U2253 ( .A(n1234), .B(out0_p2[27]), .C(N445), .D(n1233), .Z(n1609)
         );
  CANR2X1 U2254 ( .A(n1235), .B(out1_p2[27]), .C(acc[27]), .D(n1936), .Z(n1608) );
  CND2X1 U2255 ( .A(n1609), .B(n1608), .Z(n490) );
  CMX2X1 U2256 ( .A0(out1_p2[26]), .A1(N234), .S(n1260), .Z(n493) );
  CANR2X1 U2257 ( .A(n1234), .B(out0_p2[26]), .C(N444), .D(n1233), .Z(n1613)
         );
  CANR2X1 U2258 ( .A(n1235), .B(out1_p2[26]), .C(acc[26]), .D(n1936), .Z(n1612) );
  CND2X1 U2259 ( .A(n1613), .B(n1612), .Z(n492) );
  CMX2X1 U2260 ( .A0(out1_p2[25]), .A1(N233), .S(n1261), .Z(n495) );
  CANR2X1 U2261 ( .A(n1234), .B(out0_p2[25]), .C(N443), .D(n1233), .Z(n1617)
         );
  CANR2X1 U2262 ( .A(n1235), .B(out1_p2[25]), .C(acc[25]), .D(n1936), .Z(n1616) );
  CND2X1 U2263 ( .A(n1617), .B(n1616), .Z(n494) );
  CMX2X1 U2264 ( .A0(out1_p2[24]), .A1(N232), .S(n1263), .Z(n497) );
  CANR2X1 U2265 ( .A(n1234), .B(out0_p2[24]), .C(N442), .D(n1233), .Z(n1621)
         );
  CANR2X1 U2266 ( .A(n1235), .B(out1_p2[24]), .C(acc[24]), .D(n1936), .Z(n1620) );
  CND2X1 U2267 ( .A(n1621), .B(n1620), .Z(n496) );
  CMX2X1 U2268 ( .A0(out1_p2[23]), .A1(N231), .S(n1262), .Z(n499) );
  CANR2X1 U2269 ( .A(n1234), .B(out0_p2[23]), .C(N441), .D(n1233), .Z(n1625)
         );
  CANR2X1 U2270 ( .A(n1235), .B(out1_p2[23]), .C(acc[23]), .D(n1936), .Z(n1624) );
  CND2X1 U2271 ( .A(n1625), .B(n1624), .Z(n498) );
  CMX2X1 U2272 ( .A0(out1_p2[22]), .A1(N230), .S(n1262), .Z(n501) );
  CANR2X1 U2273 ( .A(n1234), .B(out0_p2[22]), .C(N440), .D(n1233), .Z(n1629)
         );
  CANR2X1 U2274 ( .A(n1235), .B(out1_p2[22]), .C(acc[22]), .D(n1936), .Z(n1628) );
  CND2X1 U2275 ( .A(n1629), .B(n1628), .Z(n500) );
  CMX2X1 U2276 ( .A0(out1_p2[21]), .A1(N229), .S(n1263), .Z(n503) );
  CANR2X1 U2277 ( .A(n1234), .B(out0_p2[21]), .C(N439), .D(n1233), .Z(n1633)
         );
  CANR2X1 U2278 ( .A(n1235), .B(out1_p2[21]), .C(acc[21]), .D(n1936), .Z(n1632) );
  CND2X1 U2279 ( .A(n1633), .B(n1632), .Z(n502) );
  CMX2X1 U2280 ( .A0(out1_p2[20]), .A1(N228), .S(n1260), .Z(n505) );
  CANR2X1 U2281 ( .A(n1234), .B(out0_p2[20]), .C(N438), .D(n1233), .Z(n1637)
         );
  CANR2X1 U2282 ( .A(n1235), .B(out1_p2[20]), .C(acc[20]), .D(n1936), .Z(n1636) );
  CND2X1 U2283 ( .A(n1637), .B(n1636), .Z(n504) );
  CMX2X1 U2284 ( .A0(out1_p2[19]), .A1(N227), .S(n1263), .Z(n507) );
  CANR2X1 U2285 ( .A(n1234), .B(out0_p2[19]), .C(N437), .D(n1233), .Z(n1641)
         );
  CANR2X1 U2286 ( .A(n1235), .B(out1_p2[19]), .C(acc[19]), .D(n1936), .Z(n1640) );
  CND2X1 U2287 ( .A(n1641), .B(n1640), .Z(n506) );
  CMX2X1 U2288 ( .A0(out1_p2[18]), .A1(N226), .S(n1260), .Z(n509) );
  CANR2X1 U2289 ( .A(n1234), .B(out0_p2[18]), .C(N436), .D(n1233), .Z(n1645)
         );
  CANR2X1 U2290 ( .A(n1235), .B(out1_p2[18]), .C(acc[18]), .D(n1936), .Z(n1644) );
  CND2X1 U2291 ( .A(n1645), .B(n1644), .Z(n508) );
  CMX2X1 U2292 ( .A0(out1_p2[17]), .A1(N225), .S(n1261), .Z(n511) );
  CANR2X1 U2293 ( .A(n1234), .B(out0_p2[17]), .C(N435), .D(n1233), .Z(n1649)
         );
  CANR2X1 U2294 ( .A(n1235), .B(out1_p2[17]), .C(acc[17]), .D(n1936), .Z(n1648) );
  CND2X1 U2295 ( .A(n1649), .B(n1648), .Z(n510) );
  CMX2X1 U2296 ( .A0(out1_p2[16]), .A1(N224), .S(n1261), .Z(n513) );
  CANR2X1 U2297 ( .A(n1234), .B(out0_p2[16]), .C(N434), .D(n1233), .Z(n1653)
         );
  CANR2X1 U2298 ( .A(n1235), .B(out1_p2[16]), .C(acc[16]), .D(n1936), .Z(n1652) );
  CND2X1 U2299 ( .A(n1653), .B(n1652), .Z(n512) );
  CIVX2 U2300 ( .A(out1_p2[16]), .Z(n1655) );
  CMX2X1 U2301 ( .A0(out1_p2[15]), .A1(N223), .S(n1260), .Z(n515) );
  CANR2X1 U2302 ( .A(n1234), .B(out0_p2[15]), .C(N433), .D(n1233), .Z(n1657)
         );
  CANR2X1 U2303 ( .A(n1235), .B(out1_p2[15]), .C(acc[15]), .D(n1936), .Z(n1656) );
  CND2X1 U2304 ( .A(n1657), .B(n1656), .Z(n514) );
  CMX2X1 U2305 ( .A0(out1_p2[14]), .A1(N222), .S(n1262), .Z(n517) );
  CANR2X1 U2306 ( .A(n1234), .B(out0_p2[14]), .C(N432), .D(n1233), .Z(n1661)
         );
  CANR2X1 U2307 ( .A(n1235), .B(out1_p2[14]), .C(acc[14]), .D(n1936), .Z(n1660) );
  CND2X1 U2308 ( .A(n1661), .B(n1660), .Z(n516) );
  CMX2X1 U2309 ( .A0(out1_p2[13]), .A1(N221), .S(n1263), .Z(n519) );
  CANR2X1 U2310 ( .A(n1234), .B(out0_p2[13]), .C(N431), .D(n1233), .Z(n1665)
         );
  CANR2X1 U2311 ( .A(n1235), .B(out1_p2[13]), .C(acc[13]), .D(n1936), .Z(n1664) );
  CND2X1 U2312 ( .A(n1665), .B(n1664), .Z(n518) );
  CMX2X1 U2313 ( .A0(out1_p2[12]), .A1(N220), .S(n1262), .Z(n521) );
  CANR2X1 U2314 ( .A(n1234), .B(out0_p2[12]), .C(N430), .D(n1233), .Z(n1669)
         );
  CANR2X1 U2315 ( .A(n1235), .B(out1_p2[12]), .C(acc[12]), .D(n1936), .Z(n1668) );
  CND2X1 U2316 ( .A(n1669), .B(n1668), .Z(n520) );
  CMX2X1 U2317 ( .A0(out1_p2[11]), .A1(N219), .S(n1261), .Z(n523) );
  CANR2X1 U2318 ( .A(n1235), .B(out1_p2[11]), .C(acc[11]), .D(n1936), .Z(n1672) );
  CND2X1 U2319 ( .A(n1673), .B(n1672), .Z(n522) );
  CMX2X1 U2320 ( .A0(out1_p2[10]), .A1(N218), .S(n1260), .Z(n525) );
  CANR2X1 U2321 ( .A(n1234), .B(out0_p2[10]), .C(N428), .D(n1233), .Z(n1677)
         );
  CANR2X1 U2322 ( .A(n1235), .B(out1_p2[10]), .C(acc[10]), .D(n1936), .Z(n1676) );
  CND2X1 U2323 ( .A(n1677), .B(n1676), .Z(n524) );
  CMX2X1 U2324 ( .A0(out1_p2[9]), .A1(N217), .S(n1261), .Z(n527) );
  CANR2X1 U2325 ( .A(n1235), .B(out1_p2[9]), .C(acc[9]), .D(n1936), .Z(n1680)
         );
  CND2X1 U2326 ( .A(n1681), .B(n1680), .Z(n526) );
  CIVX2 U2327 ( .A(out1_p2[9]), .Z(n1683) );
  CANR2X1 U2328 ( .A(n1719), .B(acc[9]), .C(n1718), .D(out0_p2[9]), .Z(n1682)
         );
  CMX2X1 U2329 ( .A0(out1_p2[8]), .A1(N216), .S(n1263), .Z(n529) );
  CANR2X1 U2330 ( .A(n1234), .B(out0_p2[8]), .C(N426), .D(n1233), .Z(n1685) );
  CANR2X1 U2331 ( .A(n1235), .B(out1_p2[8]), .C(acc[8]), .D(n1936), .Z(n1684)
         );
  CND2X1 U2332 ( .A(n1685), .B(n1684), .Z(n528) );
  CIVX2 U2333 ( .A(out1_p2[8]), .Z(n1687) );
  CMX2X1 U2334 ( .A0(out1_p2[7]), .A1(N215), .S(n1262), .Z(n531) );
  CANR2X1 U2335 ( .A(n1234), .B(out0_p2[7]), .C(N425), .D(n1233), .Z(n1689) );
  CANR2X1 U2336 ( .A(n1235), .B(out1_p2[7]), .C(acc[7]), .D(n1936), .Z(n1688)
         );
  CND2X1 U2337 ( .A(n1689), .B(n1688), .Z(n530) );
  CIVX2 U2338 ( .A(out1_p2[7]), .Z(n1691) );
  CMX2X1 U2339 ( .A0(out1_p2[6]), .A1(N214), .S(n1262), .Z(n533) );
  CANR2X1 U2340 ( .A(n1234), .B(out0_p2[6]), .C(N424), .D(n1233), .Z(n1693) );
  CANR2X1 U2341 ( .A(n1235), .B(out1_p2[6]), .C(acc[6]), .D(n1936), .Z(n1692)
         );
  CND2X1 U2342 ( .A(n1693), .B(n1692), .Z(n532) );
  CIVX2 U2343 ( .A(out1_p2[6]), .Z(n1695) );
  CMX2X1 U2344 ( .A0(out1_p2[5]), .A1(N213), .S(n1263), .Z(n535) );
  CANR2X1 U2345 ( .A(n1234), .B(out0_p2[5]), .C(N423), .D(n1233), .Z(n1697) );
  CANR2X1 U2346 ( .A(n1235), .B(out1_p2[5]), .C(acc[5]), .D(n1936), .Z(n1696)
         );
  CND2X1 U2347 ( .A(n1697), .B(n1696), .Z(n534) );
  CIVX2 U2348 ( .A(out1_p2[5]), .Z(n1699) );
  CMX2X1 U2349 ( .A0(out1_p2[4]), .A1(N212), .S(n1260), .Z(n537) );
  CANR2X1 U2350 ( .A(n1234), .B(out0_p2[4]), .C(N422), .D(n1233), .Z(n1701) );
  CANR2X1 U2351 ( .A(n1235), .B(out1_p2[4]), .C(acc[4]), .D(n1936), .Z(n1700)
         );
  CND2X1 U2352 ( .A(n1701), .B(n1700), .Z(n536) );
  CIVX2 U2353 ( .A(out1_p2[4]), .Z(n1703) );
  CMX2X1 U2354 ( .A0(out1_p2[3]), .A1(N211), .S(n1263), .Z(n539) );
  CANR2X1 U2355 ( .A(n1235), .B(out1_p2[3]), .C(acc[3]), .D(n1936), .Z(n1704)
         );
  CND2X1 U2356 ( .A(n1705), .B(n1704), .Z(n538) );
  CIVX2 U2357 ( .A(out1_p2[3]), .Z(n1707) );
  CMX2X1 U2358 ( .A0(out1_p2[2]), .A1(N210), .S(n1260), .Z(n541) );
  CANR2X1 U2359 ( .A(n1234), .B(out0_p2[2]), .C(N420), .D(n1233), .Z(n1709) );
  CANR2X1 U2360 ( .A(n1235), .B(out1_p2[2]), .C(acc[2]), .D(n1936), .Z(n1708)
         );
  CND2X1 U2361 ( .A(n1709), .B(n1708), .Z(n540) );
  CIVX2 U2362 ( .A(out1_p2[2]), .Z(n1711) );
  CMX2X1 U2363 ( .A0(out1_p2[1]), .A1(N209), .S(n1261), .Z(n543) );
  CANR2X1 U2364 ( .A(n1235), .B(out1_p2[1]), .C(acc[1]), .D(n1936), .Z(n1712)
         );
  CND2X1 U2365 ( .A(n1713), .B(n1712), .Z(n542) );
  CIVX2 U2366 ( .A(out1_p2[1]), .Z(n1715) );
  CMX2X1 U2367 ( .A0(out1_p2[0]), .A1(N208), .S(n1261), .Z(n545) );
  CANR2X1 U2368 ( .A(n1234), .B(out0_p2[0]), .C(N418), .D(n1233), .Z(n1717) );
  CANR2X1 U2369 ( .A(n1235), .B(out1_p2[0]), .C(acc[0]), .D(n1936), .Z(n1716)
         );
  CND2X1 U2370 ( .A(n1717), .B(n1716), .Z(n544) );
  CIVX2 U2371 ( .A(out1_p2[0]), .Z(n1721) );
  CMX2X1 U2372 ( .A0(out1_p2[63]), .A1(N271), .S(n1260), .Z(n419) );
  CANR2X1 U2373 ( .A(n1234), .B(out0_p2[63]), .C(N481), .D(n1233), .Z(n1724)
         );
  CANR2X1 U2374 ( .A(n1235), .B(out1_p2[63]), .C(acc[63]), .D(n1936), .Z(n1723) );
  CND2X1 U2375 ( .A(n1724), .B(n1723), .Z(n546) );
  CND2X1 U2376 ( .A(en0_p2_d1), .B(n1255), .Z(n1859) );
  CIVX2 U2377 ( .A(out0_p2[63]), .Z(n1730) );
  CIVX2 U2378 ( .A(n1726), .Z(n1856) );
  CIVX2 U2379 ( .A(n1728), .Z(n1855) );
  CIVX2 U2380 ( .A(n1070), .Z(n1941) );
  CIVX2 U2381 ( .A(cmd0[0]), .Z(n1940) );
  CIVX2 U2382 ( .A(out0_p2[0]), .Z(n1732) );
  CAN2X1 U2383 ( .A(n1861), .B(n1323), .Z(n1950) );
  CIVX2 U2384 ( .A(out0_p2[1]), .Z(n1734) );
  CIVX2 U2385 ( .A(out0_p2[2]), .Z(n1736) );
  CMXI2X1 U2386 ( .A0(n1230), .A1(n1185), .S(n1323), .Z(n2162) );
  CIVX2 U2387 ( .A(out0_p2[3]), .Z(n1738) );
  CIVX2 U2388 ( .A(out0_p2[4]), .Z(n1740) );
  CMXI2X1 U2389 ( .A0(n1229), .A1(n1227), .S(n1323), .Z(n2161) );
  CIVX2 U2390 ( .A(out0_p2[5]), .Z(n1742) );
  CIVX2 U2391 ( .A(out0_p2[6]), .Z(n1744) );
  CMXI2X1 U2392 ( .A0(n1228), .A1(n1226), .S(n1323), .Z(n2164) );
  CIVX2 U2393 ( .A(out0_p2[7]), .Z(n1746) );
  CIVX2 U2394 ( .A(out0_p2[8]), .Z(n1748) );
  CMXI2X1 U2395 ( .A0(n1225), .A1(n1223), .S(n1322), .Z(n2163) );
  CIVX2 U2396 ( .A(out0_p2[9]), .Z(n1750) );
  CIVX2 U2397 ( .A(out0_p2[10]), .Z(n1752) );
  CMXI2X1 U2398 ( .A0(n1224), .A1(n1222), .S(n1322), .Z(n1957) );
  CIVX2 U2399 ( .A(out0_p2[11]), .Z(n1754) );
  CIVX2 U2400 ( .A(out0_p2[12]), .Z(n1756) );
  CMXI2X1 U2401 ( .A0(n1221), .A1(n1219), .S(n1322), .Z(n1956) );
  CIVX2 U2402 ( .A(out0_p2[13]), .Z(n1758) );
  CIVX2 U2403 ( .A(out0_p2[14]), .Z(n1760) );
  CMXI2X1 U2404 ( .A0(n1220), .A1(n1218), .S(n1322), .Z(n1959) );
  CIVX2 U2405 ( .A(out0_p2[15]), .Z(n1762) );
  CIVX2 U2406 ( .A(out0_p2[16]), .Z(n1764) );
  CMXI2X1 U2407 ( .A0(n1217), .A1(n1215), .S(n1322), .Z(n1958) );
  CIVX2 U2408 ( .A(out0_p2[17]), .Z(n1766) );
  CIVX2 U2409 ( .A(out0_p2[18]), .Z(n1768) );
  CMXI2X1 U2410 ( .A0(n1216), .A1(n1214), .S(n1322), .Z(n1961) );
  CIVX2 U2411 ( .A(out0_p2[19]), .Z(n1770) );
  CIVX2 U2412 ( .A(out0_p2[20]), .Z(n1772) );
  CMXI2X1 U2413 ( .A0(n1213), .A1(n1211), .S(n1322), .Z(n1960) );
  CIVX2 U2414 ( .A(out0_p2[21]), .Z(n1774) );
  CIVX2 U2415 ( .A(out0_p2[22]), .Z(n1776) );
  CMXI2X1 U2416 ( .A0(n1212), .A1(n1210), .S(n1322), .Z(n1963) );
  CIVX2 U2417 ( .A(out0_p2[23]), .Z(n1778) );
  CIVX2 U2418 ( .A(out0_p2[24]), .Z(n1780) );
  CMXI2X1 U2419 ( .A0(n1209), .A1(n1207), .S(n1322), .Z(n1962) );
  CIVX2 U2420 ( .A(out0_p2[25]), .Z(n1782) );
  CIVX2 U2421 ( .A(out0_p2[26]), .Z(n1784) );
  CMXI2X1 U2422 ( .A0(n1208), .A1(n1206), .S(n1322), .Z(n1965) );
  CIVX2 U2423 ( .A(out0_p2[27]), .Z(n1786) );
  CIVX2 U2424 ( .A(out0_p2[28]), .Z(n1788) );
  CMXI2X1 U2425 ( .A0(n1205), .A1(n1203), .S(n1322), .Z(n1964) );
  CIVX2 U2426 ( .A(out0_p2[29]), .Z(n1790) );
  CIVX2 U2427 ( .A(out0_p2[30]), .Z(n1792) );
  CMXI2X1 U2428 ( .A0(n1204), .A1(n1202), .S(n1321), .Z(n1967) );
  CIVX2 U2429 ( .A(out0_p2[31]), .Z(n1794) );
  CIVX2 U2430 ( .A(out0_p2[32]), .Z(n1796) );
  CMXI2X1 U2431 ( .A0(n1201), .A1(n1192), .S(n1321), .Z(n1966) );
  CIVX2 U2432 ( .A(out0_p2[33]), .Z(n1798) );
  CIVX2 U2433 ( .A(out0_p2[34]), .Z(n1800) );
  CMXI2X1 U2434 ( .A0(n1193), .A1(n1191), .S(n1321), .Z(n1969) );
  CIVX2 U2435 ( .A(out0_p2[35]), .Z(n1802) );
  CIVX2 U2436 ( .A(out0_p2[36]), .Z(n1804) );
  CMXI2X1 U2437 ( .A0(n1190), .A1(n1188), .S(n1321), .Z(n1968) );
  CIVX2 U2438 ( .A(out0_p2[37]), .Z(n1806) );
  CIVX2 U2439 ( .A(out0_p2[38]), .Z(n1808) );
  CMXI2X1 U2440 ( .A0(n1189), .A1(n1187), .S(n1321), .Z(n1971) );
  CIVX2 U2441 ( .A(out0_p2[39]), .Z(n1810) );
  CIVX2 U2442 ( .A(out0_p2[40]), .Z(n1812) );
  CMXI2X1 U2443 ( .A0(n1186), .A1(n1197), .S(n1321), .Z(n1970) );
  CIVX2 U2444 ( .A(out0_p2[41]), .Z(n1814) );
  CIVX2 U2445 ( .A(out0_p2[42]), .Z(n1816) );
  CMXI2X1 U2446 ( .A0(n1198), .A1(n1200), .S(n1321), .Z(n1974) );
  CIVX2 U2447 ( .A(out0_p2[43]), .Z(n1818) );
  CIVX2 U2448 ( .A(out0_p2[44]), .Z(n1820) );
  CMXI2X1 U2449 ( .A0(n1199), .A1(n1195), .S(n1321), .Z(n1973) );
  CIVX2 U2450 ( .A(out0_p2[45]), .Z(n1822) );
  CIVX2 U2451 ( .A(out0_p2[46]), .Z(n1824) );
  CMXI2X1 U2452 ( .A0(n1196), .A1(n1194), .S(n1321), .Z(n1976) );
  CIVX2 U2453 ( .A(out0_p2[47]), .Z(n1826) );
  CIVX2 U2454 ( .A(out0_p2[48]), .Z(n1828) );
  CMXI2X1 U2455 ( .A0(n1177), .A1(n1178), .S(n1321), .Z(n1975) );
  CIVX2 U2456 ( .A(out0_p2[49]), .Z(n1830) );
  CIVX2 U2457 ( .A(out0_p2[50]), .Z(n1832) );
  CMXI2X1 U2458 ( .A0(n1179), .A1(n1180), .S(n1321), .Z(n1978) );
  CIVX2 U2459 ( .A(out0_p2[51]), .Z(n1834) );
  CIVX2 U2460 ( .A(out0_p2[52]), .Z(n1836) );
  CMXI2X1 U2461 ( .A0(n1181), .A1(n1182), .S(n1320), .Z(n1977) );
  CIVX2 U2462 ( .A(out0_p2[53]), .Z(n1838) );
  CIVX2 U2463 ( .A(out0_p2[54]), .Z(n1840) );
  CMXI2X1 U2464 ( .A0(n1183), .A1(n1184), .S(n1320), .Z(n1980) );
  CIVX2 U2465 ( .A(out0_p2[58]), .Z(n1842) );
  CANR2X1 U2466 ( .A(acc[58]), .B(n1856), .C(out1_p2[58]), .D(n1855), .Z(n1841) );
  CIVX2 U2467 ( .A(out0_p2[57]), .Z(n1844) );
  CIVX2 U2468 ( .A(out0_p2[55]), .Z(n1846) );
  CIVX2 U2469 ( .A(out0_p2[56]), .Z(n1848) );
  CMXI2X1 U2470 ( .A0(n1175), .A1(n1176), .S(n1320), .Z(n1979) );
  CIVX2 U2471 ( .A(out0_p2[60]), .Z(n1850) );
  CIVX2 U2472 ( .A(out0_p2[59]), .Z(n1852) );
  CIVX2 U2473 ( .A(out0_p2[62]), .Z(n1854) );
  CANR2X1 U2474 ( .A(acc[62]), .B(n1856), .C(out1_p2[62]), .D(n1855), .Z(n1853) );
  CIVX2 U2475 ( .A(out0_p2[61]), .Z(n1858) );
  CIVX2 U2476 ( .A(acc_cmd2[57]), .Z(n1860) );
  CMXI2X1 U2477 ( .A0(n1176), .A1(n1860), .S(n1318), .Z(n2028) );
  CIVX2 U2478 ( .A(h0_p0[6]), .Z(n1864) );
  CIVX2 U2479 ( .A(n787), .Z(n1875) );
  COND2X1 U2480 ( .A(n787), .B(n1864), .C(n1875), .D(n1863), .Z(n631) );
  CIVX2 U2481 ( .A(h0_p0[5]), .Z(n1866) );
  COND2X1 U2482 ( .A(n787), .B(n1866), .C(n1875), .D(n1865), .Z(n628) );
  CIVX2 U2483 ( .A(h0_p0[4]), .Z(n1868) );
  COND2X1 U2484 ( .A(n787), .B(n1868), .C(n1875), .D(n1867), .Z(n625) );
  CIVX2 U2485 ( .A(h0_p0[3]), .Z(n1870) );
  CIVX2 U2486 ( .A(h0[3]), .Z(n1869) );
  COND2X1 U2487 ( .A(n787), .B(n1870), .C(n1875), .D(n1869), .Z(n622) );
  CIVX2 U2488 ( .A(h0_p0[2]), .Z(n1872) );
  COND2X1 U2489 ( .A(n787), .B(n1872), .C(n1875), .D(n1871), .Z(n619) );
  CIVX2 U2490 ( .A(h0_p0[1]), .Z(n1874) );
  COND2X1 U2491 ( .A(n787), .B(n1874), .C(n1875), .D(n1873), .Z(n616) );
  CIVX2 U2492 ( .A(h0_p0[0]), .Z(n1876) );
  COND2X1 U2493 ( .A(n787), .B(n1876), .C(n1338), .D(n1875), .Z(n613) );
  CIVX2 U2494 ( .A(z[0]), .Z(n1881) );
  CIVX2 U2495 ( .A(acc[0]), .Z(n1880) );
  CIVX2 U2496 ( .A(n12), .Z(n1877) );
  CIVX2 U2497 ( .A(z[2]), .Z(n1883) );
  CIVX2 U2498 ( .A(acc[2]), .Z(n1882) );
  CIVX2 U2499 ( .A(z[4]), .Z(n1885) );
  CIVX2 U2500 ( .A(acc[4]), .Z(n1884) );
  CIVX2 U2501 ( .A(z[5]), .Z(n1887) );
  CIVX2 U2502 ( .A(acc[5]), .Z(n1886) );
  CIVX2 U2503 ( .A(z[6]), .Z(n1889) );
  CIVX2 U2504 ( .A(acc[6]), .Z(n1888) );
  CIVX2 U2505 ( .A(z[7]), .Z(n1891) );
  CIVX2 U2506 ( .A(acc[7]), .Z(n1890) );
  CIVX2 U2507 ( .A(z[8]), .Z(n1893) );
  CIVX2 U2508 ( .A(acc[8]), .Z(n1892) );
  CIVX2 U2509 ( .A(z[10]), .Z(n1895) );
  CIVX2 U2510 ( .A(acc[10]), .Z(n1894) );
  CIVX2 U2511 ( .A(z[12]), .Z(n1897) );
  CIVX2 U2512 ( .A(acc[12]), .Z(n1896) );
  CIVX2 U2513 ( .A(z[13]), .Z(n1899) );
  CIVX2 U2514 ( .A(acc[13]), .Z(n1898) );
  CIVX2 U2515 ( .A(z[14]), .Z(n1901) );
  CIVX2 U2516 ( .A(acc[14]), .Z(n1900) );
  CIVX2 U2517 ( .A(z[15]), .Z(n1903) );
  CIVX2 U2518 ( .A(acc[15]), .Z(n1902) );
  CIVX2 U2519 ( .A(z[16]), .Z(n1905) );
  CIVX2 U2520 ( .A(acc[16]), .Z(n1904) );
  CIVX2 U2521 ( .A(z[17]), .Z(n1907) );
  CIVX2 U2522 ( .A(acc[17]), .Z(n1906) );
  CIVX2 U2523 ( .A(z[18]), .Z(n1909) );
  CIVX2 U2524 ( .A(acc[18]), .Z(n1908) );
  CIVX2 U2525 ( .A(z[19]), .Z(n1911) );
  CIVX2 U2526 ( .A(acc[19]), .Z(n1910) );
  CIVX2 U2527 ( .A(z[20]), .Z(n1913) );
  CIVX2 U2528 ( .A(acc[20]), .Z(n1912) );
  CIVX2 U2529 ( .A(z[21]), .Z(n1915) );
  CIVX2 U2530 ( .A(acc[21]), .Z(n1914) );
  CIVX2 U2531 ( .A(z[22]), .Z(n1917) );
  CIVX2 U2532 ( .A(acc[22]), .Z(n1916) );
  CIVX2 U2533 ( .A(z[23]), .Z(n1919) );
  CIVX2 U2534 ( .A(acc[23]), .Z(n1918) );
  CIVX2 U2535 ( .A(z[24]), .Z(n1921) );
  CIVX2 U2536 ( .A(acc[24]), .Z(n1920) );
  CIVX2 U2537 ( .A(z[25]), .Z(n1923) );
  CIVX2 U2538 ( .A(acc[25]), .Z(n1922) );
  CIVX2 U2539 ( .A(z[26]), .Z(n1925) );
  CIVX2 U2540 ( .A(acc[26]), .Z(n1924) );
  CIVX2 U2541 ( .A(z[27]), .Z(n1927) );
  CIVX2 U2542 ( .A(acc[27]), .Z(n1926) );
  CIVX2 U2543 ( .A(z[28]), .Z(n1929) );
  CIVX2 U2544 ( .A(acc[28]), .Z(n1928) );
  CIVX2 U2545 ( .A(z[29]), .Z(n1931) );
  CIVX2 U2546 ( .A(acc[29]), .Z(n1930) );
  CIVX2 U2547 ( .A(z[30]), .Z(n1933) );
  CIVX2 U2548 ( .A(acc[30]), .Z(n1932) );
  CIVX2 U2549 ( .A(z[31]), .Z(n1935) );
  CIVX2 U2550 ( .A(acc[31]), .Z(n1934) );
  CIVX2 U2551 ( .A(en2_p1), .Z(n1949) );
  CMXI2X1 U2552 ( .A0(n1950), .A1(n2162), .S(n1325), .Z(n1951) );
  CMXI2X1 U2553 ( .A0(n2161), .A1(n2164), .S(n1325), .Z(n2219) );
  CMXI2X1 U2554 ( .A0(n1951), .A1(n2219), .S(n1242), .Z(n1952) );
  CMXI2X1 U2555 ( .A0(n2163), .A1(n1957), .S(n1325), .Z(n2218) );
  CMXI2X1 U2556 ( .A0(n1956), .A1(n1959), .S(n1325), .Z(n1989) );
  CMXI2X1 U2557 ( .A0(n2218), .A1(n1989), .S(n1243), .Z(n2266) );
  CMXI2X1 U2558 ( .A0(n1952), .A1(n2266), .S(n1332), .Z(n1953) );
  CMXI2X1 U2559 ( .A0(n1958), .A1(n1961), .S(n1325), .Z(n1988) );
  CMXI2X1 U2560 ( .A0(n1960), .A1(n1963), .S(n1325), .Z(n1991) );
  CMXI2X1 U2561 ( .A0(n1988), .A1(n1991), .S(n1239), .Z(n2265) );
  CMXI2X1 U2562 ( .A0(n1962), .A1(n1965), .S(n1325), .Z(n1990) );
  CMXI2X1 U2563 ( .A0(n1964), .A1(n1967), .S(n1325), .Z(n1993) );
  CMXI2X1 U2564 ( .A0(n1990), .A1(n1993), .S(n1240), .Z(n2133) );
  CMXI2X1 U2565 ( .A0(n2265), .A1(n2133), .S(n1332), .Z(n2063) );
  CMXI2X1 U2566 ( .A0(n1953), .A1(n2063), .S(n1247), .Z(n1954) );
  CMXI2X1 U2567 ( .A0(n1966), .A1(n1969), .S(n1325), .Z(n1992) );
  CMXI2X1 U2568 ( .A0(n1968), .A1(n1971), .S(n1325), .Z(n1995) );
  CMXI2X1 U2569 ( .A0(n1992), .A1(n1995), .S(n1240), .Z(n2132) );
  CMXI2X1 U2570 ( .A0(n1970), .A1(n1974), .S(n1325), .Z(n1994) );
  CMXI2X1 U2571 ( .A0(n1973), .A1(n1976), .S(n1325), .Z(n1998) );
  CMXI2X1 U2572 ( .A0(n1994), .A1(n1998), .S(n1243), .Z(n2135) );
  CMXI2X1 U2573 ( .A0(n2132), .A1(n2135), .S(n1332), .Z(n2062) );
  CMXI2X1 U2574 ( .A0(n1975), .A1(n1978), .S(n1326), .Z(n1997) );
  CMXI2X1 U2575 ( .A0(n1977), .A1(n1980), .S(n1326), .Z(n2000) );
  CMXI2X1 U2576 ( .A0(n1997), .A1(n2000), .S(n1241), .Z(n2134) );
  CMX2X1 U2577 ( .A0(acc_cmd2[58]), .A1(acc_cmd2[57]), .S(n1324), .Z(n1982) );
  CMXI2X1 U2578 ( .A0(n1979), .A1(n1982), .S(n1326), .Z(n1999) );
  CMX2X1 U2579 ( .A0(acc_cmd2[60]), .A1(acc_cmd2[59]), .S(n1324), .Z(n1981) );
  CMX2X1 U2580 ( .A0(acc_cmd2[62]), .A1(acc_cmd2[61]), .S(n1324), .Z(n1984) );
  CMXI2X1 U2581 ( .A0(n1981), .A1(n1984), .S(n1326), .Z(n2002) );
  CMXI2X1 U2582 ( .A0(n1999), .A1(n2002), .S(n1242), .Z(n2137) );
  CMXI2X1 U2583 ( .A0(n2134), .A1(n2137), .S(n1332), .Z(n2065) );
  CMXI2X1 U2584 ( .A0(n2062), .A1(n2065), .S(n1245), .Z(n2182) );
  CMXI2X1 U2585 ( .A0(n1954), .A1(n2182), .S(n1250), .Z(n1955) );
  CND2IX1 U2586 ( .B(n1250), .A(n2181), .Z(n2248) );
  CMXI2X1 U2587 ( .A0(n2249), .A1(n2033), .S(n1243), .Z(n2166) );
  CMXI2X1 U2588 ( .A0(n2032), .A1(n2035), .S(n1241), .Z(n2081) );
  CMXI2X1 U2589 ( .A0(n2034), .A1(n2037), .S(n1239), .Z(n2080) );
  CMXI2X1 U2590 ( .A0(n2036), .A1(n2039), .S(n1239), .Z(n2083) );
  CMXI2X1 U2591 ( .A0(n1972), .A1(n2146), .S(n1246), .Z(n1985) );
  CMXI2X1 U2592 ( .A0(n2038), .A1(n2042), .S(n1240), .Z(n2082) );
  CMXI2X1 U2593 ( .A0(n2041), .A1(n2044), .S(n1241), .Z(n2085) );
  CMXI2X1 U2594 ( .A0(n2082), .A1(n2085), .S(n1332), .Z(n2145) );
  CMXI2X1 U2595 ( .A0(n1982), .A1(n1981), .S(n1327), .Z(n2043) );
  CMXI2X1 U2596 ( .A0(n1984), .A1(n1983), .S(n1327), .Z(n2045) );
  CMXI2X1 U2597 ( .A0(n2043), .A1(n2045), .S(n1242), .Z(n2084) );
  CMXI2X1 U2598 ( .A0(n2145), .A1(n2147), .S(n1247), .Z(n2210) );
  CMXI2X1 U2599 ( .A0(n2096), .A1(n2005), .S(n1327), .Z(n2257) );
  CMXI2X1 U2600 ( .A0(n2004), .A1(n2007), .S(n1327), .Z(n2048) );
  CMXI2X1 U2601 ( .A0(n2257), .A1(n2048), .S(n1240), .Z(n2200) );
  CMXI2X1 U2602 ( .A0(n2006), .A1(n2009), .S(n1327), .Z(n2047) );
  CMXI2X1 U2603 ( .A0(n2008), .A1(n2011), .S(n1327), .Z(n2050) );
  CMXI2X1 U2604 ( .A0(n2047), .A1(n2050), .S(n1242), .Z(n2088) );
  CMXI2X1 U2605 ( .A0(n2010), .A1(n2013), .S(n1327), .Z(n2049) );
  CMXI2X1 U2606 ( .A0(n2012), .A1(n2015), .S(n1327), .Z(n2052) );
  CMXI2X1 U2607 ( .A0(n2049), .A1(n2052), .S(n1243), .Z(n2087) );
  CMXI2X1 U2608 ( .A0(n2014), .A1(n2017), .S(n1328), .Z(n2051) );
  CMXI2X1 U2609 ( .A0(n2016), .A1(n2019), .S(n1328), .Z(n2054) );
  CMXI2X1 U2610 ( .A0(n2051), .A1(n2054), .S(n1239), .Z(n2090) );
  CMXI2X1 U2611 ( .A0(n1986), .A1(n2150), .S(n1248), .Z(n1987) );
  CMXI2X1 U2612 ( .A0(n2018), .A1(n2022), .S(n1328), .Z(n2053) );
  CMXI2X1 U2613 ( .A0(n2021), .A1(n2024), .S(n1328), .Z(n2057) );
  CMXI2X1 U2614 ( .A0(n2053), .A1(n2057), .S(n1243), .Z(n2089) );
  CMXI2X1 U2615 ( .A0(n2023), .A1(n2026), .S(n1328), .Z(n2056) );
  CMXI2X1 U2616 ( .A0(n2056), .A1(n2059), .S(n1241), .Z(n2092) );
  CMXI2X1 U2617 ( .A0(n2089), .A1(n2092), .S(n1332), .Z(n2149) );
  CMX2X1 U2618 ( .A0(acc_cmd2[59]), .A1(acc_cmd2[58]), .S(n1324), .Z(n2027) );
  CMX2X1 U2619 ( .A0(acc_cmd2[61]), .A1(acc_cmd2[60]), .S(n1324), .Z(n2030) );
  CMXI2X1 U2620 ( .A0(n2027), .A1(n2030), .S(n1328), .Z(n2058) );
  CMX2X1 U2621 ( .A0(acc_cmd2[63]), .A1(acc_cmd2[62]), .S(n1324), .Z(n2029) );
  CMXI2X1 U2622 ( .A0(n2058), .A1(n2060), .S(n1240), .Z(n2091) );
  CMXI2X1 U2623 ( .A0(n2149), .A1(n2151), .S(n1246), .Z(n2211) );
  CMXI2X1 U2624 ( .A0(n2220), .A1(n2105), .S(n1332), .Z(n1996) );
  CMXI2X1 U2625 ( .A0(n2104), .A1(n2107), .S(n1332), .Z(n2154) );
  CMXI2X1 U2626 ( .A0(n1996), .A1(n2154), .S(n1248), .Z(n2003) );
  CMXI2X1 U2627 ( .A0(n2106), .A1(n2109), .S(n1333), .Z(n2153) );
  CMXI2X1 U2628 ( .A0(n2002), .A1(n2001), .S(n1240), .Z(n2108) );
  CMXI2X1 U2629 ( .A0(n2153), .A1(n2155), .S(n1249), .Z(n2212) );
  CMXI2X1 U2630 ( .A0(n2005), .A1(n2004), .S(n1328), .Z(n2097) );
  CMXI2X1 U2631 ( .A0(n2007), .A1(n2006), .S(n1328), .Z(n2068) );
  CMXI2X1 U2632 ( .A0(n2097), .A1(n2068), .S(n1240), .Z(n2238) );
  CMXI2X1 U2633 ( .A0(n2009), .A1(n2008), .S(n1328), .Z(n2067) );
  CMXI2X1 U2634 ( .A0(n2011), .A1(n2010), .S(n1328), .Z(n2070) );
  CMXI2X1 U2635 ( .A0(n2067), .A1(n2070), .S(n1243), .Z(n2112) );
  CMXI2X1 U2636 ( .A0(n2013), .A1(n2012), .S(n1328), .Z(n2069) );
  CMXI2X1 U2637 ( .A0(n2015), .A1(n2014), .S(n1329), .Z(n2072) );
  CMXI2X1 U2638 ( .A0(n2069), .A1(n2072), .S(n1241), .Z(n2111) );
  CMXI2X1 U2639 ( .A0(n2017), .A1(n2016), .S(n1329), .Z(n2071) );
  CMXI2X1 U2640 ( .A0(n2019), .A1(n2018), .S(n1329), .Z(n2074) );
  CMXI2X1 U2641 ( .A0(n2071), .A1(n2074), .S(n1242), .Z(n2114) );
  CMXI2X1 U2642 ( .A0(n2020), .A1(n2158), .S(n1244), .Z(n2031) );
  CMXI2X1 U2643 ( .A0(n2022), .A1(n2021), .S(n1329), .Z(n2073) );
  CMXI2X1 U2644 ( .A0(n2024), .A1(n2023), .S(n1329), .Z(n2076) );
  CMXI2X1 U2645 ( .A0(n2073), .A1(n2076), .S(n1243), .Z(n2113) );
  CMXI2X1 U2646 ( .A0(n2026), .A1(n2025), .S(n1329), .Z(n2075) );
  CMXI2X1 U2647 ( .A0(n2028), .A1(n2027), .S(n1329), .Z(n2078) );
  CMXI2X1 U2648 ( .A0(n2075), .A1(n2078), .S(n1241), .Z(n2116) );
  CMXI2X1 U2649 ( .A0(n2113), .A1(n2116), .S(n1333), .Z(n2157) );
  CMXI2X1 U2650 ( .A0(n2030), .A1(n2029), .S(n1329), .Z(n2077) );
  CMXI2X1 U2651 ( .A0(n2157), .A1(n2159), .S(n1245), .Z(n2213) );
  CMXI2X1 U2652 ( .A0(n2033), .A1(n2032), .S(n1239), .Z(n2251) );
  CMXI2X1 U2653 ( .A0(n2035), .A1(n2034), .S(n1239), .Z(n2119) );
  CMXI2X1 U2654 ( .A0(n2037), .A1(n2036), .S(n1240), .Z(n2118) );
  CMXI2X1 U2655 ( .A0(n2039), .A1(n2038), .S(n1241), .Z(n2121) );
  CMXI2X1 U2656 ( .A0(n2040), .A1(n2174), .S(n1246), .Z(n2046) );
  CMXI2X1 U2657 ( .A0(n2042), .A1(n2041), .S(n1242), .Z(n2120) );
  CMXI2X1 U2658 ( .A0(n2044), .A1(n2043), .S(n1240), .Z(n2123) );
  CMXI2X1 U2659 ( .A0(n2120), .A1(n2123), .S(n1333), .Z(n2173) );
  CMXI2X1 U2660 ( .A0(n2173), .A1(n2175), .S(n1247), .Z(n2214) );
  CMXI2X1 U2661 ( .A0(n2048), .A1(n2047), .S(n1242), .Z(n2259) );
  CMXI2X1 U2662 ( .A0(n2050), .A1(n2049), .S(n1243), .Z(n2126) );
  CMXI2X1 U2663 ( .A0(n2052), .A1(n2051), .S(n1239), .Z(n2125) );
  CMXI2X1 U2664 ( .A0(n2054), .A1(n2053), .S(n1243), .Z(n2128) );
  CMXI2X1 U2665 ( .A0(n2055), .A1(n2178), .S(n1249), .Z(n2061) );
  CMXI2X1 U2666 ( .A0(n2057), .A1(n2056), .S(n1241), .Z(n2127) );
  CMXI2X1 U2667 ( .A0(n2059), .A1(n2058), .S(n1240), .Z(n2130) );
  CMXI2X1 U2668 ( .A0(n2127), .A1(n2130), .S(n1333), .Z(n2177) );
  CMXI2X1 U2669 ( .A0(n2177), .A1(n2179), .S(n1247), .Z(n2215) );
  CMXI2X1 U2670 ( .A0(n2065), .A1(n2064), .S(n1249), .Z(n2216) );
  CMXI2X1 U2671 ( .A0(n2068), .A1(n2067), .S(n1241), .Z(n2271) );
  CMXI2X1 U2672 ( .A0(n2070), .A1(n2069), .S(n1242), .Z(n2140) );
  CMXI2X1 U2673 ( .A0(n2271), .A1(n2140), .S(n1333), .Z(n2099) );
  CMXI2X1 U2674 ( .A0(n2072), .A1(n2071), .S(n1239), .Z(n2139) );
  CMXI2X1 U2675 ( .A0(n2074), .A1(n2073), .S(n1242), .Z(n2142) );
  CMXI2X1 U2676 ( .A0(n2139), .A1(n2142), .S(n1333), .Z(n2102) );
  CMXI2X1 U2677 ( .A0(n2099), .A1(n2102), .S(n1244), .Z(n2079) );
  CMXI2X1 U2678 ( .A0(n2076), .A1(n2075), .S(n1243), .Z(n2141) );
  CMXI2X1 U2679 ( .A0(n2078), .A1(n2077), .S(n1239), .Z(n2143) );
  CMXI2X1 U2680 ( .A0(n2141), .A1(n2143), .S(n1334), .Z(n2101) );
  CMXI2X1 U2681 ( .A0(n2081), .A1(n2080), .S(n1334), .Z(n2168) );
  CMXI2X1 U2682 ( .A0(n2083), .A1(n2082), .S(n1334), .Z(n2171) );
  CMXI2X1 U2683 ( .A0(n2168), .A1(n2171), .S(n1248), .Z(n2086) );
  CMXI2X1 U2684 ( .A0(n2085), .A1(n2084), .S(n1334), .Z(n2170) );
  CMXI2X1 U2685 ( .A0(n2088), .A1(n2087), .S(n1334), .Z(n2202) );
  CMXI2X1 U2686 ( .A0(n2090), .A1(n2089), .S(n1334), .Z(n2186) );
  CMXI2X1 U2687 ( .A0(n2202), .A1(n2186), .S(n1244), .Z(n2093) );
  CMXI2X1 U2688 ( .A0(n2092), .A1(n2091), .S(n1334), .Z(n2185) );
  CMXI2X1 U2689 ( .A0(n2094), .A1(n2196), .S(n1329), .Z(n2095) );
  CMXI2X1 U2690 ( .A0(n2195), .A1(n2198), .S(n1329), .Z(n2237) );
  CMXI2X1 U2691 ( .A0(n2095), .A1(n2237), .S(n1240), .Z(n2098) );
  CMXI2X1 U2692 ( .A0(n2197), .A1(n2096), .S(n1329), .Z(n2236) );
  CMXI2X1 U2693 ( .A0(n2236), .A1(n2097), .S(n1240), .Z(n2272) );
  CMXI2X1 U2694 ( .A0(n2100), .A1(n2099), .S(n1245), .Z(n2103) );
  CMXI2X1 U2695 ( .A0(n2102), .A1(n2101), .S(n1246), .Z(n2183) );
  CMXI2X1 U2696 ( .A0(n2105), .A1(n2104), .S(n1334), .Z(n2222) );
  CMXI2X1 U2697 ( .A0(n2107), .A1(n2106), .S(n1334), .Z(n2188) );
  CMXI2X1 U2698 ( .A0(n2222), .A1(n2188), .S(n1247), .Z(n2110) );
  CMXI2X1 U2699 ( .A0(n2109), .A1(n2108), .S(n1334), .Z(n2187) );
  CMXI2X1 U2700 ( .A0(n2112), .A1(n2111), .S(n1334), .Z(n2240) );
  CMXI2X1 U2701 ( .A0(n2114), .A1(n2113), .S(n1335), .Z(n2190) );
  CMXI2X1 U2702 ( .A0(n2240), .A1(n2190), .S(n1248), .Z(n2117) );
  CMXI2X1 U2703 ( .A0(n2116), .A1(n2115), .S(n1335), .Z(n2189) );
  CMXI2X1 U2704 ( .A0(n2119), .A1(n2118), .S(n1335), .Z(n2253) );
  CMXI2X1 U2705 ( .A0(n2121), .A1(n2120), .S(n1335), .Z(n2192) );
  CMXI2X1 U2706 ( .A0(n2253), .A1(n2192), .S(n1249), .Z(n2124) );
  CMXI2X1 U2707 ( .A0(n2123), .A1(n2122), .S(n1335), .Z(n2191) );
  CMXI2X1 U2708 ( .A0(n2126), .A1(n2125), .S(n1335), .Z(n2261) );
  CMXI2X1 U2709 ( .A0(n2128), .A1(n2127), .S(n1335), .Z(n2194) );
  CMXI2X1 U2710 ( .A0(n2261), .A1(n2194), .S(n1245), .Z(n2131) );
  CMXI2X1 U2711 ( .A0(n2130), .A1(n2129), .S(n1335), .Z(n2193) );
  CMXI2X1 U2712 ( .A0(n2267), .A1(n2207), .S(n1249), .Z(n2138) );
  CMXI2X1 U2713 ( .A0(n2137), .A1(n2136), .S(n1335), .Z(n2206) );
  CMXI2X1 U2714 ( .A0(n2142), .A1(n2141), .S(n1336), .Z(n2209) );
  CMXI2X1 U2715 ( .A0(n2273), .A1(n2209), .S(n1244), .Z(n2144) );
  CMXI2X1 U2716 ( .A0(n2146), .A1(n2145), .S(n1245), .Z(n2148) );
  CMXI2X1 U2717 ( .A0(n2150), .A1(n2149), .S(n1246), .Z(n2152) );
  CMXI2X1 U2718 ( .A0(n2154), .A1(n2153), .S(n1244), .Z(n2156) );
  CMXI2X1 U2719 ( .A0(n2158), .A1(n2157), .S(n1246), .Z(n2160) );
  CMXI2X1 U2720 ( .A0(n2165), .A1(n2250), .S(n1243), .Z(n2167) );
  CMXI2X1 U2721 ( .A0(n2169), .A1(n2168), .S(n1247), .Z(n2172) );
  CMXI2X1 U2722 ( .A0(n2171), .A1(n2170), .S(n1248), .Z(n2184) );
  CMXI2X1 U2723 ( .A0(n2174), .A1(n2173), .S(n1249), .Z(n2176) );
  CMXI2X1 U2724 ( .A0(n2178), .A1(n2177), .S(n1244), .Z(n2180) );
  CMXI2X1 U2725 ( .A0(n2186), .A1(n2185), .S(n1245), .Z(n2204) );
  CMXI2X1 U2726 ( .A0(n2188), .A1(n2187), .S(n1247), .Z(n2224) );
  CMXI2X1 U2727 ( .A0(n2190), .A1(n2189), .S(n1245), .Z(n2242) );
  CMXI2X1 U2728 ( .A0(n2192), .A1(n2191), .S(n1246), .Z(n2255) );
  CMXI2X1 U2729 ( .A0(n2194), .A1(n2193), .S(n1247), .Z(n2263) );
  CMXI2X1 U2730 ( .A0(n2198), .A1(n2197), .S(n1330), .Z(n2258) );
  CMXI2X1 U2731 ( .A0(n2199), .A1(n2258), .S(n1241), .Z(n2201) );
  CMXI2X1 U2732 ( .A0(n2203), .A1(n2202), .S(n1248), .Z(n2205) );
  CMXI2X1 U2733 ( .A0(n2207), .A1(n2206), .S(n1246), .Z(n2269) );
  CMXI2X1 U2734 ( .A0(n2209), .A1(n2208), .S(n1248), .Z(n2275) );
  CMXI2X1 U2735 ( .A0(n2223), .A1(n2222), .S(n1249), .Z(n2225) );
  CMXI2X1 U2736 ( .A0(n2241), .A1(n2240), .S(n1244), .Z(n2243) );
  CMXI2X1 U2737 ( .A0(n2254), .A1(n2253), .S(n1245), .Z(n2256) );
  CMXI2X1 U2738 ( .A0(n2262), .A1(n2261), .S(n1246), .Z(n2264) );
  CMXI2X1 U2739 ( .A0(n2268), .A1(n2267), .S(n1247), .Z(n2270) );
  CMXI2X1 U2740 ( .A0(n2274), .A1(n2273), .S(n1249), .Z(n2276) );
endmodule

