
module sfilt_DW02_mult_3_stage_J1_0 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, \A_extended[32] , \B_extended[32] , \mult_x_1/n1740 ,
         \mult_x_1/n1692 , \mult_x_1/n1685 , \mult_x_1/n1684 ,
         \mult_x_1/n1676 , \mult_x_1/n1675 , \mult_x_1/n1674 ,
         \mult_x_1/n1669 , \mult_x_1/n1667 , \mult_x_1/n1666 ,
         \mult_x_1/n1657 , \mult_x_1/n1655 , \mult_x_1/n1654 ,
         \mult_x_1/n1645 , \mult_x_1/n1643 , \mult_x_1/n1642 ,
         \mult_x_1/n1631 , \mult_x_1/n1629 , \mult_x_1/n1628 ,
         \mult_x_1/n1617 , \mult_x_1/n1615 , \mult_x_1/n1614 ,
         \mult_x_1/n1601 , \mult_x_1/n1600 , \mult_x_1/n1599 ,
         \mult_x_1/n1598 , \mult_x_1/n1589 , \mult_x_1/n1587 ,
         \mult_x_1/n1585 , \mult_x_1/n1584 , \mult_x_1/n1571 ,
         \mult_x_1/n1569 , \mult_x_1/n1567 , \mult_x_1/n1566 ,
         \mult_x_1/n1553 , \mult_x_1/n1551 , \mult_x_1/n1549 ,
         \mult_x_1/n1548 , \mult_x_1/n1533 , \mult_x_1/n1531 ,
         \mult_x_1/n1529 , \mult_x_1/n1528 , \mult_x_1/n1513 ,
         \mult_x_1/n1511 , \mult_x_1/n1509 , \mult_x_1/n1508 ,
         \mult_x_1/n1491 , \mult_x_1/n1490 , \mult_x_1/n1489 ,
         \mult_x_1/n1488 , \mult_x_1/n1487 , \mult_x_1/n1486 ,
         \mult_x_1/n1471 , \mult_x_1/n1469 , \mult_x_1/n1468 ,
         \mult_x_1/n1467 , \mult_x_1/n1466 , \mult_x_1/n1447 ,
         \mult_x_1/n1445 , \mult_x_1/n1444 , \mult_x_1/n1443 ,
         \mult_x_1/n1442 , \mult_x_1/n1423 , \mult_x_1/n1421 ,
         \mult_x_1/n1420 , \mult_x_1/n1419 , \mult_x_1/n1418 ,
         \mult_x_1/n1397 , \mult_x_1/n1395 , \mult_x_1/n1394 ,
         \mult_x_1/n1393 , \mult_x_1/n1392 , \mult_x_1/n1371 ,
         \mult_x_1/n1369 , \mult_x_1/n1368 , \mult_x_1/n1367 ,
         \mult_x_1/n1366 , \mult_x_1/n1343 , \mult_x_1/n1341 ,
         \mult_x_1/n1340 , \mult_x_1/n1339 , \mult_x_1/n1338 ,
         \mult_x_1/n1315 , \mult_x_1/n1314 , \mult_x_1/n1313 ,
         \mult_x_1/n1312 , \mult_x_1/n1311 , \mult_x_1/n1310 ,
         \mult_x_1/n1289 , \mult_x_1/n1287 , \mult_x_1/n1285 ,
         \mult_x_1/n1284 , \mult_x_1/n1283 , \mult_x_1/n1282 ,
         \mult_x_1/n1259 , \mult_x_1/n1257 , \mult_x_1/n1255 ,
         \mult_x_1/n1254 , \mult_x_1/n1253 , \mult_x_1/n1252 ,
         \mult_x_1/n1229 , \mult_x_1/n1227 , \mult_x_1/n1226 ,
         \mult_x_1/n1225 , \mult_x_1/n1224 , \mult_x_1/n1223 ,
         \mult_x_1/n1222 , \mult_x_1/n1199 , \mult_x_1/n1197 ,
         \mult_x_1/n1196 , \mult_x_1/n1195 , \mult_x_1/n1194 ,
         \mult_x_1/n1173 , \mult_x_1/n1171 , \mult_x_1/n1169 ,
         \mult_x_1/n1168 , \mult_x_1/n1167 , \mult_x_1/n1166 ,
         \mult_x_1/n1147 , \mult_x_1/n1145 , \mult_x_1/n1143 ,
         \mult_x_1/n1141 , \mult_x_1/n1140 , \mult_x_1/n1117 ,
         \mult_x_1/n1115 , \mult_x_1/n1114 , \mult_x_1/n1113 ,
         \mult_x_1/n1112 , \mult_x_1/n1093 , \mult_x_1/n1091 ,
         \mult_x_1/n1090 , \mult_x_1/n1089 , \mult_x_1/n1088 ,
         \mult_x_1/n1069 , \mult_x_1/n1067 , \mult_x_1/n1066 ,
         \mult_x_1/n1065 , \mult_x_1/n1064 , \mult_x_1/n1047 ,
         \mult_x_1/n1045 , \mult_x_1/n1044 , \mult_x_1/n1043 ,
         \mult_x_1/n1042 , \mult_x_1/n1025 , \mult_x_1/n1023 ,
         \mult_x_1/n1022 , \mult_x_1/n1021 , \mult_x_1/n1020 ,
         \mult_x_1/n1005 , \mult_x_1/n1003 , \mult_x_1/n1002 ,
         \mult_x_1/n1001 , \mult_x_1/n1000 , \mult_x_1/n985 , \mult_x_1/n983 ,
         \mult_x_1/n981 , \mult_x_1/n980 , \mult_x_1/n963 , \mult_x_1/n962 ,
         \mult_x_1/n961 , \mult_x_1/n960 , \mult_x_1/n945 , \mult_x_1/n944 ,
         \mult_x_1/n943 , \mult_x_1/n942 , \mult_x_1/n929 , \mult_x_1/n928 ,
         \mult_x_1/n927 , \mult_x_1/n926 , \mult_x_1/n913 , \mult_x_1/n912 ,
         \mult_x_1/n911 , \mult_x_1/n910 , \mult_x_1/n899 , \mult_x_1/n897 ,
         \mult_x_1/n883 , \mult_x_1/n881 , \mult_x_1/n880 , \mult_x_1/n872 ,
         \mult_x_1/n871 , \mult_x_1/n870 , \mult_x_1/n869 , \mult_x_1/n868 ,
         \mult_x_1/n861 , \mult_x_1/n859 , \mult_x_1/n858 , \mult_x_1/n853 ,
         \mult_x_1/n851 , \mult_x_1/n850 , \mult_x_1/n849 , \mult_x_1/n848 ,
         \mult_x_1/n841 , \mult_x_1/n839 , \mult_x_1/n838 , \mult_x_1/n829 ,
         \mult_x_1/n828 , \mult_x_1/n823 , \mult_x_1/n821 , \mult_x_1/n820 ,
         \mult_x_1/n817 , \mult_x_1/n815 , \mult_x_1/n807 , \mult_x_1/n806 ,
         \mult_x_1/n803 , \mult_x_1/n796 , \mult_x_1/n794 , \mult_x_1/n739 ,
         \mult_x_1/n702 , \mult_x_1/n701 , \mult_x_1/n700 , \mult_x_1/n697 ,
         \mult_x_1/n696 , \mult_x_1/n542 , \mult_x_1/n531 , \mult_x_1/n524 ,
         \mult_x_1/n513 , \mult_x_1/n506 , \mult_x_1/n495 , \mult_x_1/n486 ,
         \mult_x_1/n472 , \mult_x_1/n471 , \mult_x_1/n461 , \mult_x_1/n460 ,
         \mult_x_1/n452 , \mult_x_1/n451 , \mult_x_1/n441 , \mult_x_1/n440 ,
         \mult_x_1/n428 , \mult_x_1/n427 , \mult_x_1/n413 , \mult_x_1/n412 ,
         \mult_x_1/n406 , \mult_x_1/n405 , \mult_x_1/n395 , \mult_x_1/n394 ,
         \mult_x_1/n382 , \mult_x_1/n381 , \mult_x_1/n373 , \mult_x_1/n372 ,
         \mult_x_1/n354 , \mult_x_1/n353 , \mult_x_1/n349 , \mult_x_1/n332 ,
         \mult_x_1/n331 , \mult_x_1/n323 , \mult_x_1/n320 , \mult_x_1/n308 ,
         \mult_x_1/n307 , \mult_x_1/n303 , \mult_x_1/n286 , \mult_x_1/n283 ,
         \mult_x_1/n273 , \mult_x_1/n272 , \mult_x_1/n255 , \mult_x_1/n246 ,
         \mult_x_1/n236 , \mult_x_1/n233 , \mult_x_1/n179 , \mult_x_1/n178 ,
         \mult_x_1/n177 , \mult_x_1/n176 , \mult_x_1/n175 , \mult_x_1/n174 ,
         \mult_x_1/n173 , \mult_x_1/n172 , \mult_x_1/n171 , \mult_x_1/n170 ,
         \mult_x_1/n169 , \mult_x_1/n168 , \mult_x_1/n167 , \mult_x_1/n166 ,
         \mult_x_1/n165 , \mult_x_1/n164 , \mult_x_1/n163 , \mult_x_1/n162 ,
         \mult_x_1/n161 , \mult_x_1/n160 , \mult_x_1/n159 , \mult_x_1/n158 ,
         \mult_x_1/n156 , \mult_x_1/n153 , \mult_x_1/n149 , n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2847,
         n2849, n2851, n2853, n2855, n2857, n2859, n2861;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  CFD1QX1 clk_r_REG211_S2 ( .D(n2891), .CP(CLK), .Q(PRODUCT[28]) );
  CFD1QX1 clk_r_REG216_S2 ( .D(n2892), .CP(CLK), .Q(PRODUCT[27]) );
  CFD1QX1 clk_r_REG225_S2 ( .D(n2893), .CP(CLK), .Q(PRODUCT[26]) );
  CFD1QX1 clk_r_REG228_S2 ( .D(n2894), .CP(CLK), .Q(PRODUCT[25]) );
  CFD1QX1 clk_r_REG236_S2 ( .D(n2895), .CP(CLK), .Q(PRODUCT[24]) );
  CFD1QX1 clk_r_REG239_S2 ( .D(n2896), .CP(CLK), .Q(PRODUCT[23]) );
  CFD1QX1 clk_r_REG247_S2 ( .D(n2897), .CP(CLK), .Q(PRODUCT[22]) );
  CFD1QX1 clk_r_REG252_S2 ( .D(n2898), .CP(CLK), .Q(PRODUCT[21]) );
  CFD1QX1 clk_r_REG260_S2 ( .D(n2899), .CP(CLK), .Q(PRODUCT[20]) );
  CFD1QX1 clk_r_REG262_S2 ( .D(n2900), .CP(CLK), .Q(PRODUCT[19]) );
  CFD1QX1 clk_r_REG270_S2 ( .D(n2901), .CP(CLK), .Q(PRODUCT[18]) );
  CFD1QX1 clk_r_REG275_S2 ( .D(n2902), .CP(CLK), .Q(PRODUCT[17]) );
  CFD1QX1 clk_r_REG282_S2 ( .D(n2903), .CP(CLK), .Q(PRODUCT[16]) );
  CFD1QX1 clk_r_REG285_S2 ( .D(n2904), .CP(CLK), .Q(PRODUCT[15]) );
  CFD1QX1 clk_r_REG291_S2 ( .D(n2905), .CP(CLK), .Q(PRODUCT[14]) );
  CFD1QX1 clk_r_REG293_S2 ( .D(n2906), .CP(CLK), .Q(PRODUCT[13]) );
  CFD1QX1 clk_r_REG300_S2 ( .D(n2907), .CP(CLK), .Q(PRODUCT[12]) );
  CFD1QX1 clk_r_REG303_S2 ( .D(n2908), .CP(CLK), .Q(PRODUCT[11]) );
  CFD1QX1 clk_r_REG309_S2 ( .D(n58), .CP(CLK), .Q(PRODUCT[10]) );
  CFD1QX1 clk_r_REG313_S2 ( .D(n2910), .CP(CLK), .Q(PRODUCT[9]) );
  CFD1QX1 clk_r_REG316_S2 ( .D(n59), .CP(CLK), .Q(PRODUCT[8]) );
  CFD1QX1 clk_r_REG319_S2 ( .D(n50), .CP(CLK), .Q(PRODUCT[7]) );
  CFD1QX1 clk_r_REG322_S2 ( .D(n54), .CP(CLK), .Q(PRODUCT[6]) );
  CFD1QX1 clk_r_REG324_S2 ( .D(n44), .CP(CLK), .Q(PRODUCT[5]) );
  CFD1QX1 clk_r_REG326_S2 ( .D(n46), .CP(CLK), .Q(PRODUCT[4]) );
  CFD1QX1 clk_r_REG328_S2 ( .D(n48), .CP(CLK), .Q(PRODUCT[3]) );
  CFD1QX1 clk_r_REG330_S2 ( .D(n40), .CP(CLK), .Q(PRODUCT[2]) );
  CFD1QX1 clk_r_REG332_S2 ( .D(n42), .CP(CLK), .Q(PRODUCT[1]) );
  CFD1QX1 clk_r_REG334_S2 ( .D(n38), .CP(CLK), .Q(PRODUCT[0]) );
  CFD1QXL clk_r_REG323_S1 ( .D(n2913), .CP(CLK), .Q(n2857) );
  CFD1QXL clk_r_REG325_S1 ( .D(n2914), .CP(CLK), .Q(n2855) );
  CFD1QXL clk_r_REG327_S1 ( .D(n2915), .CP(CLK), .Q(n2853) );
  CFD1QXL clk_r_REG329_S1 ( .D(n2916), .CP(CLK), .Q(n2851) );
  CFD1QXL clk_r_REG331_S1 ( .D(n2917), .CP(CLK), .Q(n2849) );
  CFD1QXL clk_r_REG333_S1 ( .D(n2918), .CP(CLK), .Q(n2847) );
  CFD1QXL \mult_x_1/clk_r_REG175_S1  ( .D(\mult_x_1/n1145 ), .CP(CLK), .Q(
        n2722) );
  CFD1QXL \mult_x_1/clk_r_REG117_S2  ( .D(\mult_x_1/n233 ), .CP(CLK), .Q(n2567) );
  CFD1QXL \mult_x_1/clk_r_REG320_S1  ( .D(\mult_x_1/n702 ), .CP(CLK), .Q(n2634) );
  CFD1QXL \mult_x_1/clk_r_REG311_S1  ( .D(\mult_x_1/n1692 ), .CP(CLK), .Q(
        n2840) );
  CFD1QXL \mult_x_1/clk_r_REG301_S1  ( .D(\mult_x_1/n1674 ), .CP(CLK), .Q(
        n2835) );
  CFD1QXL \mult_x_1/clk_r_REG144_S2  ( .D(n23), .CP(CLK), .Q(n2637) );
  CFD1QXL \mult_x_1/clk_r_REG289_S1  ( .D(\mult_x_1/n1601 ), .CP(CLK), .Q(
        n2819) );
  CFD1QXL \mult_x_1/clk_r_REG277_S1  ( .D(\mult_x_1/n1585 ), .CP(CLK), .Q(
        n2813) );
  CFD1QXL \mult_x_1/clk_r_REG272_S1  ( .D(\mult_x_1/n1567 ), .CP(CLK), .Q(
        n2809) );
  CFD1QXL \mult_x_1/clk_r_REG264_S1  ( .D(\mult_x_1/n1549 ), .CP(CLK), .Q(
        n2805) );
  CFD1QXL \mult_x_1/clk_r_REG251_S1  ( .D(\mult_x_1/n1529 ), .CP(CLK), .Q(
        n2801) );
  CFD1QXL \mult_x_1/clk_r_REG249_S1  ( .D(\mult_x_1/n1487 ), .CP(CLK), .Q(
        n2791) );
  CFD1QXL \mult_x_1/clk_r_REG214_S1  ( .D(\mult_x_1/n1392 ), .CP(CLK), .Q(
        n2770) );
  CFD1QXL \mult_x_1/clk_r_REG185_S1  ( .D(\mult_x_1/n1341 ), .CP(CLK), .Q(
        n2763) );
  CFD1QXL \mult_x_1/clk_r_REG190_S1  ( .D(\mult_x_1/n1313 ), .CP(CLK), .Q(
        n2757) );
  CFD1QXL \mult_x_1/clk_r_REG1_S1  ( .D(\mult_x_1/n1283 ), .CP(CLK), .Q(n2749)
         );
  CFD1QXL \mult_x_1/clk_r_REG197_S1  ( .D(\mult_x_1/n1169 ), .CP(CLK), .Q(
        n2727) );
  CFD1QXL \mult_x_1/clk_r_REG196_S1  ( .D(\mult_x_1/n1168 ), .CP(CLK), .Q(
        n2726) );
  CFD1QXL \mult_x_1/clk_r_REG201_S1  ( .D(\mult_x_1/n1117 ), .CP(CLK), .Q(
        n2718) );
  CFD1QXL \mult_x_1/clk_r_REG176_S1  ( .D(\mult_x_1/n1112 ), .CP(CLK), .Q(
        n2714) );
  CFD1QXL \mult_x_1/clk_r_REG202_S1  ( .D(\mult_x_1/n1088 ), .CP(CLK), .Q(
        n2709) );
  CFD1QXL \mult_x_1/clk_r_REG62_S1  ( .D(\mult_x_1/n1064 ), .CP(CLK), .Q(n2704) );
  CFD1QXL \mult_x_1/clk_r_REG64_S1  ( .D(\mult_x_1/n1042 ), .CP(CLK), .Q(n2699) );
  CFD1QXL \mult_x_1/clk_r_REG74_S1  ( .D(\mult_x_1/n1020 ), .CP(CLK), .Q(n2694) );
  CFD1QXL \mult_x_1/clk_r_REG76_S1  ( .D(\mult_x_1/n1000 ), .CP(CLK), .Q(n2689) );
  CFD1QXL \mult_x_1/clk_r_REG204_S1  ( .D(\mult_x_1/n980 ), .CP(CLK), .Q(n2685) );
  CFD1QXL \mult_x_1/clk_r_REG169_S1  ( .D(\mult_x_1/n945 ), .CP(CLK), .Q(n2680) );
  CFD1QXL \mult_x_1/clk_r_REG168_S1  ( .D(\mult_x_1/n944 ), .CP(CLK), .Q(n2679) );
  CFD1QXL \mult_x_1/clk_r_REG95_S1  ( .D(\mult_x_1/n943 ), .CP(CLK), .Q(n2678)
         );
  CFD1QXL \mult_x_1/clk_r_REG161_S1  ( .D(\mult_x_1/n928 ), .CP(CLK), .Q(n2675) );
  CFD1QXL \mult_x_1/clk_r_REG98_S1  ( .D(\mult_x_1/n927 ), .CP(CLK), .Q(n2674)
         );
  CFD1QXL \mult_x_1/clk_r_REG170_S1  ( .D(\mult_x_1/n912 ), .CP(CLK), .Q(n2671) );
  CFD1QXL \mult_x_1/clk_r_REG164_S1  ( .D(\mult_x_1/n911 ), .CP(CLK), .Q(n2670) );
  CFD1QXL \mult_x_1/clk_r_REG165_S1  ( .D(\mult_x_1/n897 ), .CP(CLK), .Q(n2667) );
  CFD1QXL \mult_x_1/clk_r_REG195_S1  ( .D(\mult_x_1/n883 ), .CP(CLK), .Q(n2666) );
  CFD1QXL \mult_x_1/clk_r_REG104_S1  ( .D(\mult_x_1/n871 ), .CP(CLK), .Q(n2662) );
  CFD1QXL \mult_x_1/clk_r_REG129_S1  ( .D(\mult_x_1/n861 ), .CP(CLK), .Q(n2658) );
  CFD1QXL \mult_x_1/clk_r_REG122_S1  ( .D(\mult_x_1/n859 ), .CP(CLK), .Q(n2657) );
  CFD1QXL \mult_x_1/clk_r_REG133_S1  ( .D(\mult_x_1/n851 ), .CP(CLK), .Q(n2654) );
  CFD1QXL \mult_x_1/clk_r_REG132_S1  ( .D(\mult_x_1/n850 ), .CP(CLK), .Q(n2653) );
  CFD1QXL \mult_x_1/clk_r_REG131_S1  ( .D(\mult_x_1/n849 ), .CP(CLK), .Q(n2652) );
  CFD1QXL \mult_x_1/clk_r_REG126_S1  ( .D(\mult_x_1/n839 ), .CP(CLK), .Q(n2649) );
  CFD1QXL \mult_x_1/clk_r_REG125_S1  ( .D(\mult_x_1/n838 ), .CP(CLK), .Q(n2648) );
  CFD1QXL \mult_x_1/clk_r_REG193_S1  ( .D(\mult_x_1/n823 ), .CP(CLK), .Q(n2645) );
  CFD1QXL \mult_x_1/clk_r_REG147_S1  ( .D(\mult_x_1/n817 ), .CP(CLK), .Q(n2642) );
  CFD1QXL \mult_x_1/clk_r_REG294_S1  ( .D(\mult_x_1/n1642 ), .CP(CLK), .Q(
        n2826) );
  CFD1QXL \mult_x_1/clk_r_REG283_S1  ( .D(\mult_x_1/n1628 ), .CP(CLK), .Q(
        n2823) );
  CFD1QXL \mult_x_1/clk_r_REG286_S1  ( .D(\mult_x_1/n1614 ), .CP(CLK), .Q(
        n2820) );
  CFD1QXL \mult_x_1/clk_r_REG273_S1  ( .D(\mult_x_1/n1598 ), .CP(CLK), .Q(
        n2816) );
  CFD1QXL \mult_x_1/clk_r_REG24_S1  ( .D(\mult_x_1/n1252 ), .CP(CLK), .Q(n2742) );
  CFD1QXL \mult_x_1/clk_r_REG19_S1  ( .D(\mult_x_1/n1194 ), .CP(CLK), .Q(n2730) );
  CFD1QXL \mult_x_1/clk_r_REG83_S1  ( .D(\mult_x_1/n1166 ), .CP(CLK), .Q(n2724) );
  CFD1QXL \mult_x_1/clk_r_REG85_S1  ( .D(\mult_x_1/n1140 ), .CP(CLK), .Q(n2719) );
  CFD1QXL \mult_x_1/clk_r_REG203_S1  ( .D(\mult_x_1/n1089 ), .CP(CLK), .Q(
        n2710) );
  CFD1QXL \mult_x_1/clk_r_REG65_S1  ( .D(\mult_x_1/n1043 ), .CP(CLK), .Q(n2700) );
  CFD1QXL \mult_x_1/clk_r_REG75_S1  ( .D(\mult_x_1/n1021 ), .CP(CLK), .Q(n2695) );
  CFD1QXL \mult_x_1/clk_r_REG77_S1  ( .D(\mult_x_1/n1001 ), .CP(CLK), .Q(n2690) );
  CFD1QXL \mult_x_1/clk_r_REG205_S1  ( .D(\mult_x_1/n981 ), .CP(CLK), .Q(n2686) );
  CFD1QXL \mult_x_1/clk_r_REG92_S1  ( .D(\mult_x_1/n963 ), .CP(CLK), .Q(n2684)
         );
  CFD1QXL \mult_x_1/clk_r_REG91_S1  ( .D(\mult_x_1/n962 ), .CP(CLK), .Q(n2683)
         );
  CFD1QXL \mult_x_1/clk_r_REG162_S1  ( .D(\mult_x_1/n929 ), .CP(CLK), .Q(n2676) );
  CFD1QXL \mult_x_1/clk_r_REG171_S1  ( .D(\mult_x_1/n913 ), .CP(CLK), .Q(n2672) );
  CFD1QXL \mult_x_1/clk_r_REG180_S1  ( .D(\mult_x_1/n899 ), .CP(CLK), .Q(n2668) );
  CFD1QXL \mult_x_1/clk_r_REG166_S1  ( .D(\mult_x_1/n880 ), .CP(CLK), .Q(n2664) );
  CFD1QXL \mult_x_1/clk_r_REG219_S1  ( .D(\mult_x_1/n872 ), .CP(CLK), .Q(n2663) );
  CFD1QXL \mult_x_1/clk_r_REG178_S1  ( .D(\mult_x_1/n868 ), .CP(CLK), .Q(n2659) );
  CFD1QXL \mult_x_1/clk_r_REG124_S1  ( .D(\mult_x_1/n853 ), .CP(CLK), .Q(n2655) );
  CFD1QXL \mult_x_1/clk_r_REG194_S1  ( .D(\mult_x_1/n841 ), .CP(CLK), .Q(n2650) );
  CFD1QXL \mult_x_1/clk_r_REG135_S1  ( .D(\mult_x_1/n829 ), .CP(CLK), .Q(n2647) );
  CFD1QXL \mult_x_1/clk_r_REG138_S1  ( .D(\mult_x_1/n821 ), .CP(CLK), .Q(n2644) );
  CFD1QXL \mult_x_1/clk_r_REG137_S1  ( .D(\mult_x_1/n820 ), .CP(CLK), .Q(n2643) );
  CFD1QXL \mult_x_1/clk_r_REG315_S1  ( .D(\mult_x_1/n701 ), .CP(CLK), .Q(n2612) );
  CFD1QXL \mult_x_1/clk_r_REG158_S2  ( .D(n25), .CP(CLK), .Q(n2551) );
  CFD1QXL \mult_x_1/clk_r_REG307_S1  ( .D(\mult_x_1/n1684 ), .CP(CLK), .Q(
        n2838) );
  CFD1QXL \mult_x_1/clk_r_REG317_S1  ( .D(\mult_x_1/n700 ), .CP(CLK), .Q(n2611) );
  CFD1QXL \mult_x_1/clk_r_REG306_S1  ( .D(\mult_x_1/n1655 ), .CP(CLK), .Q(
        n2830) );
  CFD1QXL \mult_x_1/clk_r_REG287_S1  ( .D(\mult_x_1/n1615 ), .CP(CLK), .Q(
        n2821) );
  CFD1QXL \mult_x_1/clk_r_REG220_S1  ( .D(\mult_x_1/n1143 ), .CP(CLK), .Q(
        n2721) );
  CFD1QXL \mult_x_1/clk_r_REG86_S1  ( .D(\mult_x_1/n1141 ), .CP(CLK), .Q(n2720) );
  CFD1QXL \mult_x_1/clk_r_REG68_S1  ( .D(\mult_x_1/n1115 ), .CP(CLK), .Q(n2717) );
  CFD1QXL \mult_x_1/clk_r_REG159_S1  ( .D(\mult_x_1/n960 ), .CP(CLK), .Q(n2681) );
  CFD1QXL \mult_x_1/clk_r_REG94_S1  ( .D(\mult_x_1/n942 ), .CP(CLK), .Q(n2677)
         );
  CFD1QXL \mult_x_1/clk_r_REG97_S1  ( .D(\mult_x_1/n926 ), .CP(CLK), .Q(n2673)
         );
  CFD1QXL \mult_x_1/clk_r_REG163_S1  ( .D(\mult_x_1/n910 ), .CP(CLK), .Q(n2669) );
  CFD1QXL \mult_x_1/clk_r_REG103_S1  ( .D(\mult_x_1/n870 ), .CP(CLK), .Q(n2661) );
  CFD1QXL \mult_x_1/clk_r_REG179_S1  ( .D(\mult_x_1/n869 ), .CP(CLK), .Q(n2660) );
  CFD1QXL \mult_x_1/clk_r_REG121_S1  ( .D(\mult_x_1/n858 ), .CP(CLK), .Q(n2656) );
  CFD1QXL \mult_x_1/clk_r_REG130_S1  ( .D(\mult_x_1/n848 ), .CP(CLK), .Q(n2651) );
  CFD1QXL \mult_x_1/clk_r_REG134_S1  ( .D(\mult_x_1/n828 ), .CP(CLK), .Q(n2646) );
  CFD1QXL \mult_x_1/clk_r_REG152_S1  ( .D(\mult_x_1/n815 ), .CP(CLK), .Q(n2641) );
  CFD1QXL \mult_x_1/clk_r_REG174_S2  ( .D(n26), .CP(CLK), .Q(n2633) );
  CFD1QXL \mult_x_1/clk_r_REG111_S2  ( .D(\mult_x_1/n236 ), .CP(CLK), .Q(n2614) );
  CFD1QXL \mult_x_1/clk_r_REG61_S2  ( .D(\mult_x_1/n170 ), .CP(CLK), .Q(n2597)
         );
  CFD1QXL \mult_x_1/clk_r_REG73_S2  ( .D(\mult_x_1/n168 ), .CP(CLK), .Q(n2594)
         );
  CFD1QXL \mult_x_1/clk_r_REG78_S2  ( .D(\mult_x_1/n167 ), .CP(CLK), .Q(n2592)
         );
  CFD1QXL \mult_x_1/clk_r_REG90_S2  ( .D(\mult_x_1/n166 ), .CP(CLK), .Q(n2591)
         );
  CFD1QXL \mult_x_1/clk_r_REG93_S2  ( .D(\mult_x_1/n165 ), .CP(CLK), .Q(n2589)
         );
  CFD1QXL \mult_x_1/clk_r_REG96_S2  ( .D(\mult_x_1/n164 ), .CP(CLK), .Q(n2587)
         );
  CFD1QXL \mult_x_1/clk_r_REG99_S2  ( .D(\mult_x_1/n163 ), .CP(CLK), .Q(n2586)
         );
  CFD1QXL \mult_x_1/clk_r_REG106_S2  ( .D(\mult_x_1/n161 ), .CP(CLK), .Q(n2582) );
  CFD1QXL \mult_x_1/clk_r_REG119_S2  ( .D(\mult_x_1/n160 ), .CP(CLK), .Q(n2581) );
  CFD1QXL \mult_x_1/clk_r_REG120_S2  ( .D(\mult_x_1/n159 ), .CP(CLK), .Q(n2580) );
  CFD1QXL \mult_x_1/clk_r_REG123_S2  ( .D(\mult_x_1/n158 ), .CP(CLK), .Q(n2578) );
  CFD1QXL \mult_x_1/clk_r_REG136_S2  ( .D(\mult_x_1/n156 ), .CP(CLK), .Q(n2575) );
  CFD1QXL \mult_x_1/clk_r_REG156_S2  ( .D(n30), .CP(CLK), .Q(n2570) );
  CFD1QXL \mult_x_1/clk_r_REG142_S2  ( .D(n29), .CP(CLK), .Q(n2568) );
  CFD1QXL \mult_x_1/clk_r_REG40_S2  ( .D(\mult_x_1/n406 ), .CP(CLK), .Q(n2621)
         );
  CFD1QXL \mult_x_1/clk_r_REG43_S2  ( .D(\mult_x_1/n373 ), .CP(CLK), .Q(n2619)
         );
  CFD1QXL \mult_x_1/clk_r_REG42_S2  ( .D(\mult_x_1/n413 ), .CP(CLK), .Q(n2564)
         );
  CFD1QXL \mult_x_1/clk_r_REG44_S2  ( .D(\mult_x_1/n382 ), .CP(CLK), .Q(n2562)
         );
  CFD1QXL \mult_x_1/clk_r_REG155_S2  ( .D(n33), .CP(CLK), .Q(n2552) );
  CFD1QXL \mult_x_1/clk_r_REG139_S2  ( .D(n32), .CP(CLK), .Q(n2573) );
  CFD1QXL \mult_x_1/clk_r_REG143_S1  ( .D(n2844), .CP(CLK), .Q(n2549) );
  CFD1QXL \mult_x_1/clk_r_REG157_S1  ( .D(n2843), .CP(CLK), .Q(n2550) );
  CFD1QXL \mult_x_1/clk_r_REG153_S1  ( .D(\mult_x_1/n803 ), .CP(CLK), .Q(n2638) );
  CFD1QXL \mult_x_1/clk_r_REG148_S1  ( .D(\mult_x_1/n806 ), .CP(CLK), .Q(n2639) );
  CFD1QXL \mult_x_1/clk_r_REG154_S1  ( .D(\mult_x_1/n255 ), .CP(CLK), .Q(n2571) );
  CFD1QXL \mult_x_1/clk_r_REG141_S1  ( .D(\mult_x_1/n246 ), .CP(CLK), .Q(n2569) );
  CFD1QXL \mult_x_1/clk_r_REG149_S1  ( .D(\mult_x_1/n807 ), .CP(CLK), .Q(n2640) );
  CFD1QXL \mult_x_1/clk_r_REG145_S1  ( .D(\mult_x_1/n794 ), .CP(CLK), .Q(n2841) );
  CFD1QXL \mult_x_1/clk_r_REG140_S1  ( .D(\mult_x_1/n796 ), .CP(CLK), .Q(n2636) );
  CFD1QXL \mult_x_1/clk_r_REG173_S1  ( .D(\mult_x_1/n1740 ), .CP(CLK), .Q(
        n2632) );
  CFD1QX1 \mult_x_1/clk_r_REG146_S2  ( .D(n34), .CP(CLK), .Q(n2842) );
  CFD1QX1 \mult_x_1/clk_r_REG310_S1  ( .D(\mult_x_1/n1676 ), .CP(CLK), .Q(
        n2837) );
  CFD1QX1 \mult_x_1/clk_r_REG304_S1  ( .D(\mult_x_1/n1669 ), .CP(CLK), .Q(
        n2834) );
  CFD1QX1 \mult_x_1/clk_r_REG299_S1  ( .D(\mult_x_1/n1667 ), .CP(CLK), .Q(
        n2833) );
  CFD1QX1 \mult_x_1/clk_r_REG298_S1  ( .D(\mult_x_1/n1666 ), .CP(CLK), .Q(
        n2832) );
  CFD1QX1 \mult_x_1/clk_r_REG292_S1  ( .D(\mult_x_1/n1657 ), .CP(CLK), .Q(
        n2831) );
  CFD1QX1 \mult_x_1/clk_r_REG305_S1  ( .D(\mult_x_1/n1654 ), .CP(CLK), .Q(
        n2829) );
  CFD1QX1 \mult_x_1/clk_r_REG290_S1  ( .D(\mult_x_1/n1645 ), .CP(CLK), .Q(
        n2828) );
  CFD1QX1 \mult_x_1/clk_r_REG295_S1  ( .D(\mult_x_1/n1643 ), .CP(CLK), .Q(
        n2827) );
  CFD1QX1 \mult_x_1/clk_r_REG296_S1  ( .D(\mult_x_1/n1631 ), .CP(CLK), .Q(
        n2825) );
  CFD1QX1 \mult_x_1/clk_r_REG281_S1  ( .D(\mult_x_1/n1617 ), .CP(CLK), .Q(
        n2822) );
  CFD1QX1 \mult_x_1/clk_r_REG288_S1  ( .D(\mult_x_1/n1600 ), .CP(CLK), .Q(
        n2818) );
  CFD1QX1 \mult_x_1/clk_r_REG276_S1  ( .D(\mult_x_1/n1584 ), .CP(CLK), .Q(
        n2812) );
  CFD1QX1 \mult_x_1/clk_r_REG261_S1  ( .D(\mult_x_1/n1571 ), .CP(CLK), .Q(
        n2811) );
  CFD1QX1 \mult_x_1/clk_r_REG297_S1  ( .D(\mult_x_1/n1569 ), .CP(CLK), .Q(
        n2810) );
  CFD1QX1 \mult_x_1/clk_r_REG271_S1  ( .D(\mult_x_1/n1566 ), .CP(CLK), .Q(
        n2808) );
  CFD1QX1 \mult_x_1/clk_r_REG280_S1  ( .D(\mult_x_1/n1553 ), .CP(CLK), .Q(
        n2807) );
  CFD1QX1 \mult_x_1/clk_r_REG259_S1  ( .D(\mult_x_1/n1551 ), .CP(CLK), .Q(
        n2806) );
  CFD1QX1 \mult_x_1/clk_r_REG263_S1  ( .D(\mult_x_1/n1548 ), .CP(CLK), .Q(
        n2804) );
  CFD1QX1 \mult_x_1/clk_r_REG265_S1  ( .D(\mult_x_1/n1533 ), .CP(CLK), .Q(
        n2803) );
  CFD1QX1 \mult_x_1/clk_r_REG268_S1  ( .D(\mult_x_1/n1531 ), .CP(CLK), .Q(
        n2802) );
  CFD1QX1 \mult_x_1/clk_r_REG250_S1  ( .D(\mult_x_1/n1528 ), .CP(CLK), .Q(
        n2800) );
  CFD1QX1 \mult_x_1/clk_r_REG246_S1  ( .D(\mult_x_1/n1513 ), .CP(CLK), .Q(
        n2799) );
  CFD1QX1 \mult_x_1/clk_r_REG253_S1  ( .D(\mult_x_1/n1511 ), .CP(CLK), .Q(
        n2798) );
  CFD1QX1 \mult_x_1/clk_r_REG254_S1  ( .D(\mult_x_1/n1508 ), .CP(CLK), .Q(
        n2796) );
  CFD1QX1 \mult_x_1/clk_r_REG257_S1  ( .D(\mult_x_1/n1491 ), .CP(CLK), .Q(
        n2795) );
  CFD1QX1 \mult_x_1/clk_r_REG238_S1  ( .D(\mult_x_1/n1489 ), .CP(CLK), .Q(
        n2793) );
  CFD1QX1 \mult_x_1/clk_r_REG237_S1  ( .D(\mult_x_1/n1488 ), .CP(CLK), .Q(
        n2792) );
  CFD1QX1 \mult_x_1/clk_r_REG248_S1  ( .D(\mult_x_1/n1486 ), .CP(CLK), .Q(
        n2790) );
  CFD1QX1 \mult_x_1/clk_r_REG245_S1  ( .D(\mult_x_1/n1469 ), .CP(CLK), .Q(
        n2788) );
  CFD1QX1 \mult_x_1/clk_r_REG241_S1  ( .D(\mult_x_1/n1467 ), .CP(CLK), .Q(
        n2786) );
  CFD1QX1 \mult_x_1/clk_r_REG240_S1  ( .D(\mult_x_1/n1466 ), .CP(CLK), .Q(
        n2785) );
  CFD1QX1 \mult_x_1/clk_r_REG243_S1  ( .D(\mult_x_1/n1445 ), .CP(CLK), .Q(
        n2783) );
  CFD1QX1 \mult_x_1/clk_r_REG227_S1  ( .D(\mult_x_1/n1443 ), .CP(CLK), .Q(
        n2781) );
  CFD1QX1 \mult_x_1/clk_r_REG226_S1  ( .D(\mult_x_1/n1442 ), .CP(CLK), .Q(
        n2780) );
  CFD1QX1 \mult_x_1/clk_r_REG232_S1  ( .D(\mult_x_1/n1421 ), .CP(CLK), .Q(
        n2778) );
  CFD1QX1 \mult_x_1/clk_r_REG231_S1  ( .D(\mult_x_1/n1420 ), .CP(CLK), .Q(
        n2777) );
  CFD1QX1 \mult_x_1/clk_r_REG229_S1  ( .D(\mult_x_1/n1418 ), .CP(CLK), .Q(
        n2775) );
  CFD1QX1 \mult_x_1/clk_r_REG233_S1  ( .D(\mult_x_1/n1397 ), .CP(CLK), .Q(
        n2774) );
  CFD1QX1 \mult_x_1/clk_r_REG267_S1  ( .D(\mult_x_1/n1395 ), .CP(CLK), .Q(
        n2773) );
  CFD1QX1 \mult_x_1/clk_r_REG266_S1  ( .D(\mult_x_1/n1394 ), .CP(CLK), .Q(
        n2772) );
  CFD1QX1 \mult_x_1/clk_r_REG215_S1  ( .D(\mult_x_1/n1393 ), .CP(CLK), .Q(
        n2771) );
  CFD1QX1 \mult_x_1/clk_r_REG223_S1  ( .D(\mult_x_1/n1371 ), .CP(CLK), .Q(
        n2769) );
  CFD1QX1 \mult_x_1/clk_r_REG218_S1  ( .D(\mult_x_1/n1369 ), .CP(CLK), .Q(
        n2768) );
  CFD1QX1 \mult_x_1/clk_r_REG217_S1  ( .D(\mult_x_1/n1368 ), .CP(CLK), .Q(
        n2767) );
  CFD1QX1 \mult_x_1/clk_r_REG209_S1  ( .D(\mult_x_1/n1366 ), .CP(CLK), .Q(
        n2765) );
  CFD1QX1 \mult_x_1/clk_r_REG222_S1  ( .D(\mult_x_1/n1343 ), .CP(CLK), .Q(
        n2764) );
  CFD1QX1 \mult_x_1/clk_r_REG184_S1  ( .D(\mult_x_1/n1340 ), .CP(CLK), .Q(
        n2762) );
  CFD1QX1 \mult_x_1/clk_r_REG212_S1  ( .D(\mult_x_1/n1338 ), .CP(CLK), .Q(
        n2760) );
  CFD1QX1 \mult_x_1/clk_r_REG188_S1  ( .D(\mult_x_1/n1315 ), .CP(CLK), .Q(
        n2759) );
  CFD1QX1 \mult_x_1/clk_r_REG187_S1  ( .D(\mult_x_1/n1314 ), .CP(CLK), .Q(
        n2758) );
  CFD1QX1 \mult_x_1/clk_r_REG189_S1  ( .D(\mult_x_1/n1312 ), .CP(CLK), .Q(
        n2756) );
  CFD1QX1 \mult_x_1/clk_r_REG181_S1  ( .D(\mult_x_1/n1310 ), .CP(CLK), .Q(
        n2754) );
  CFD1QX1 \mult_x_1/clk_r_REG200_S1  ( .D(\mult_x_1/n1289 ), .CP(CLK), .Q(
        n2753) );
  CFD1QX1 \mult_x_1/clk_r_REG23_S1  ( .D(\mult_x_1/n1287 ), .CP(CLK), .Q(n2752) );
  CFD1QX1 \mult_x_1/clk_r_REG192_S1  ( .D(\mult_x_1/n1285 ), .CP(CLK), .Q(
        n2751) );
  CFD1QX1 \mult_x_1/clk_r_REG191_S1  ( .D(\mult_x_1/n1284 ), .CP(CLK), .Q(
        n2750) );
  CFD1QX1 \mult_x_1/clk_r_REG0_S1  ( .D(\mult_x_1/n1282 ), .CP(CLK), .Q(n2748)
         );
  CFD1QX1 \mult_x_1/clk_r_REG258_S1  ( .D(\mult_x_1/n1259 ), .CP(CLK), .Q(
        n2747) );
  CFD1QX1 \mult_x_1/clk_r_REG199_S1  ( .D(\mult_x_1/n1257 ), .CP(CLK), .Q(
        n2746) );
  CFD1QX1 \mult_x_1/clk_r_REG16_S1  ( .D(\mult_x_1/n1255 ), .CP(CLK), .Q(n2745) );
  CFD1QX1 \mult_x_1/clk_r_REG15_S1  ( .D(\mult_x_1/n1254 ), .CP(CLK), .Q(n2744) );
  CFD1QX1 \mult_x_1/clk_r_REG18_S1  ( .D(\mult_x_1/n1229 ), .CP(CLK), .Q(n2741) );
  CFD1QX1 \mult_x_1/clk_r_REG88_S1  ( .D(\mult_x_1/n1227 ), .CP(CLK), .Q(n2740) );
  CFD1QX1 \mult_x_1/clk_r_REG27_S1  ( .D(\mult_x_1/n1225 ), .CP(CLK), .Q(n2738) );
  CFD1QX1 \mult_x_1/clk_r_REG26_S1  ( .D(\mult_x_1/n1224 ), .CP(CLK), .Q(n2737) );
  CFD1QX1 \mult_x_1/clk_r_REG28_S1  ( .D(\mult_x_1/n1222 ), .CP(CLK), .Q(n2735) );
  CFD1QX1 \mult_x_1/clk_r_REG82_S1  ( .D(\mult_x_1/n1199 ), .CP(CLK), .Q(n2734) );
  CFD1QX1 \mult_x_1/clk_r_REG31_S1  ( .D(\mult_x_1/n1197 ), .CP(CLK), .Q(n2733) );
  CFD1QX1 \mult_x_1/clk_r_REG30_S1  ( .D(\mult_x_1/n1196 ), .CP(CLK), .Q(n2732) );
  CFD1QX1 \mult_x_1/clk_r_REG20_S1  ( .D(\mult_x_1/n1195 ), .CP(CLK), .Q(n2731) );
  CFD1QX1 \mult_x_1/clk_r_REG172_S1  ( .D(\mult_x_1/n1173 ), .CP(CLK), .Q(
        n2729) );
  CFD1QX1 \mult_x_1/clk_r_REG221_S1  ( .D(\mult_x_1/n1171 ), .CP(CLK), .Q(
        n2728) );
  CFD1QX1 \mult_x_1/clk_r_REG198_S1  ( .D(\mult_x_1/n1147 ), .CP(CLK), .Q(
        n2723) );
  CFD1QX1 \mult_x_1/clk_r_REG67_S1  ( .D(\mult_x_1/n1114 ), .CP(CLK), .Q(n2716) );
  CFD1QX1 \mult_x_1/clk_r_REG69_S1  ( .D(\mult_x_1/n1093 ), .CP(CLK), .Q(n2713) );
  CFD1QX1 \mult_x_1/clk_r_REG33_S1  ( .D(\mult_x_1/n1091 ), .CP(CLK), .Q(n2712) );
  CFD1QX1 \mult_x_1/clk_r_REG32_S1  ( .D(\mult_x_1/n1090 ), .CP(CLK), .Q(n2711) );
  CFD1QX1 \mult_x_1/clk_r_REG70_S1  ( .D(\mult_x_1/n1069 ), .CP(CLK), .Q(n2708) );
  CFD1QX1 \mult_x_1/clk_r_REG80_S1  ( .D(\mult_x_1/n1067 ), .CP(CLK), .Q(n2707) );
  CFD1QX1 \mult_x_1/clk_r_REG79_S1  ( .D(\mult_x_1/n1066 ), .CP(CLK), .Q(n2706) );
  CFD1QX1 \mult_x_1/clk_r_REG81_S1  ( .D(\mult_x_1/n1047 ), .CP(CLK), .Q(n2703) );
  CFD1QX1 \mult_x_1/clk_r_REG72_S1  ( .D(\mult_x_1/n1045 ), .CP(CLK), .Q(n2702) );
  CFD1QX1 \mult_x_1/clk_r_REG71_S1  ( .D(\mult_x_1/n1044 ), .CP(CLK), .Q(n2701) );
  CFD1QX1 \mult_x_1/clk_r_REG102_S1  ( .D(\mult_x_1/n1025 ), .CP(CLK), .Q(
        n2698) );
  CFD1QX1 \mult_x_1/clk_r_REG207_S1  ( .D(\mult_x_1/n1023 ), .CP(CLK), .Q(
        n2697) );
  CFD1QX1 \mult_x_1/clk_r_REG206_S1  ( .D(\mult_x_1/n1022 ), .CP(CLK), .Q(
        n2696) );
  CFD1QX1 \mult_x_1/clk_r_REG208_S1  ( .D(\mult_x_1/n1005 ), .CP(CLK), .Q(
        n2693) );
  CFD1QX1 \mult_x_1/clk_r_REG101_S1  ( .D(\mult_x_1/n1003 ), .CP(CLK), .Q(
        n2692) );
  CFD1QX1 \mult_x_1/clk_r_REG100_S1  ( .D(\mult_x_1/n1002 ), .CP(CLK), .Q(
        n2691) );
  CFD1QX1 \mult_x_1/clk_r_REG89_S1  ( .D(\mult_x_1/n985 ), .CP(CLK), .Q(n2688)
         );
  CFD1QX1 \mult_x_1/clk_r_REG234_S1  ( .D(\mult_x_1/n983 ), .CP(CLK), .Q(n2687) );
  CFD1QX1 \mult_x_1/clk_r_REG3_S2  ( .D(\mult_x_1/n542 ), .CP(CLK), .Q(n2631)
         );
  CFD1QX1 \mult_x_1/clk_r_REG5_S2  ( .D(\mult_x_1/n531 ), .CP(CLK), .Q(n2630)
         );
  CFD1QX1 \mult_x_1/clk_r_REG6_S2  ( .D(\mult_x_1/n524 ), .CP(CLK), .Q(n2629)
         );
  CFD1QX1 \mult_x_1/clk_r_REG7_S2  ( .D(\mult_x_1/n513 ), .CP(CLK), .Q(n2628)
         );
  CFD1QX1 \mult_x_1/clk_r_REG36_S2  ( .D(\mult_x_1/n461 ), .CP(CLK), .Q(n2624)
         );
  CFD1QX1 \mult_x_1/clk_r_REG37_S2  ( .D(\mult_x_1/n452 ), .CP(CLK), .Q(n2623)
         );
  CFD1QX1 \mult_x_1/clk_r_REG38_S2  ( .D(\mult_x_1/n428 ), .CP(CLK), .Q(n2622)
         );
  CFD1QX1 \mult_x_1/clk_r_REG41_S2  ( .D(\mult_x_1/n395 ), .CP(CLK), .Q(n2620)
         );
  CFD1QX1 \mult_x_1/clk_r_REG45_S2  ( .D(\mult_x_1/n354 ), .CP(CLK), .Q(n2618)
         );
  CFD1QX1 \mult_x_1/clk_r_REG108_S2  ( .D(\mult_x_1/n323 ), .CP(CLK), .Q(n2617) );
  CFD1QX1 \mult_x_1/clk_r_REG46_S2  ( .D(\mult_x_1/n308 ), .CP(CLK), .Q(n2616)
         );
  CFD1QX1 \mult_x_1/clk_r_REG110_S2  ( .D(\mult_x_1/n286 ), .CP(CLK), .Q(n2615) );
  CFD1QX1 \mult_x_1/clk_r_REG12_S2  ( .D(\mult_x_1/n179 ), .CP(CLK), .Q(n2613)
         );
  CFD1QX1 \mult_x_1/clk_r_REG13_S2  ( .D(\mult_x_1/n178 ), .CP(CLK), .Q(n2608)
         );
  CFD1QX1 \mult_x_1/clk_r_REG14_S2  ( .D(\mult_x_1/n177 ), .CP(CLK), .Q(n2607)
         );
  CFD1QX1 \mult_x_1/clk_r_REG17_S2  ( .D(\mult_x_1/n176 ), .CP(CLK), .Q(n2606)
         );
  CFD1QX1 \mult_x_1/clk_r_REG21_S2  ( .D(\mult_x_1/n175 ), .CP(CLK), .Q(n2605)
         );
  CFD1QX1 \mult_x_1/clk_r_REG22_S2  ( .D(\mult_x_1/n174 ), .CP(CLK), .Q(n2604)
         );
  CFD1QX1 \mult_x_1/clk_r_REG34_S2  ( .D(\mult_x_1/n173 ), .CP(CLK), .Q(n2603)
         );
  CFD1QX1 \mult_x_1/clk_r_REG35_S2  ( .D(\mult_x_1/n472 ), .CP(CLK), .Q(n2602)
         );
  CFD1QX1 \mult_x_1/clk_r_REG48_S2  ( .D(\mult_x_1/n471 ), .CP(CLK), .Q(n2601)
         );
  CFD1QX1 \mult_x_1/clk_r_REG47_S2  ( .D(\mult_x_1/n172 ), .CP(CLK), .Q(n2600)
         );
  CFD1QX1 \mult_x_1/clk_r_REG60_S2  ( .D(\mult_x_1/n171 ), .CP(CLK), .Q(n2599)
         );
  CFD1QX1 \mult_x_1/clk_r_REG49_S2  ( .D(\mult_x_1/n460 ), .CP(CLK), .Q(n2598)
         );
  CFD1QX1 \mult_x_1/clk_r_REG50_S2  ( .D(\mult_x_1/n451 ), .CP(CLK), .Q(n2596)
         );
  CFD1QX1 \mult_x_1/clk_r_REG66_S2  ( .D(\mult_x_1/n169 ), .CP(CLK), .Q(n2595)
         );
  CFD1QX1 \mult_x_1/clk_r_REG51_S2  ( .D(\mult_x_1/n427 ), .CP(CLK), .Q(n2593)
         );
  CFD1QX1 \mult_x_1/clk_r_REG53_S2  ( .D(\mult_x_1/n405 ), .CP(CLK), .Q(n2590)
         );
  CFD1QX1 \mult_x_1/clk_r_REG54_S2  ( .D(\mult_x_1/n394 ), .CP(CLK), .Q(n2588)
         );
  CFD1QX1 \mult_x_1/clk_r_REG56_S2  ( .D(\mult_x_1/n372 ), .CP(CLK), .Q(n2585)
         );
  CFD1QX1 \mult_x_1/clk_r_REG58_S2  ( .D(\mult_x_1/n353 ), .CP(CLK), .Q(n2583)
         );
  CFD1QX1 \mult_x_1/clk_r_REG114_S2  ( .D(\mult_x_1/n320 ), .CP(CLK), .Q(n2579) );
  CFD1QX1 \mult_x_1/clk_r_REG59_S2  ( .D(\mult_x_1/n307 ), .CP(CLK), .Q(n2577)
         );
  CFD1QX1 \mult_x_1/clk_r_REG127_S2  ( .D(\mult_x_1/n303 ), .CP(CLK), .Q(n2576) );
  CFD1QX1 \mult_x_1/clk_r_REG151_S2  ( .D(n36), .CP(CLK), .Q(n2572) );
  CFD1QX1 \mult_x_1/clk_r_REG39_S2  ( .D(\mult_x_1/n441 ), .CP(CLK), .Q(n2566)
         );
  CFD1QX1 \mult_x_1/clk_r_REG52_S2  ( .D(\mult_x_1/n440 ), .CP(CLK), .Q(n2565)
         );
  CFD1QX1 \mult_x_1/clk_r_REG55_S2  ( .D(\mult_x_1/n412 ), .CP(CLK), .Q(n2563)
         );
  CFD1QX1 \mult_x_1/clk_r_REG57_S2  ( .D(\mult_x_1/n381 ), .CP(CLK), .Q(n2561)
         );
  CFD1QX1 \mult_x_1/clk_r_REG107_S2  ( .D(\mult_x_1/n349 ), .CP(CLK), .Q(n2560) );
  CFD1QX1 \mult_x_1/clk_r_REG113_S2  ( .D(n2845), .CP(CLK), .Q(n2559) );
  CFD1QX1 \mult_x_1/clk_r_REG109_S2  ( .D(\mult_x_1/n332 ), .CP(CLK), .Q(n2558) );
  CFD1QX1 \mult_x_1/clk_r_REG115_S2  ( .D(\mult_x_1/n331 ), .CP(CLK), .Q(n2557) );
  CFD1QX1 \mult_x_1/clk_r_REG128_S2  ( .D(\mult_x_1/n739 ), .CP(CLK), .Q(n2556) );
  CFD1QX1 \mult_x_1/clk_r_REG112_S2  ( .D(\mult_x_1/n273 ), .CP(CLK), .Q(n2555) );
  CFD1QX1 \mult_x_1/clk_r_REG118_S2  ( .D(\mult_x_1/n272 ), .CP(CLK), .Q(n2554) );
  CFD1QX1 \mult_x_1/clk_r_REG150_S2  ( .D(n37), .CP(CLK), .Q(n2553) );
  CFD1QX1 \mult_x_1/clk_r_REG213_S1  ( .D(\mult_x_1/n1339 ), .CP(CLK), .Q(
        n2761) );
  CFD1QX2 clk_r_REG183_S2 ( .D(n2889), .CP(CLK), .Q(PRODUCT[30]) );
  CFD1QX1 \mult_x_1/clk_r_REG160_S1  ( .D(\mult_x_1/n961 ), .CP(CLK), .Q(n2682) );
  CFD1QX2 clk_r_REG2_S2 ( .D(n2888), .CP(CLK), .Q(PRODUCT[31]) );
  CFD1QX2 clk_r_REG186_S2 ( .D(n2890), .CP(CLK), .Q(PRODUCT[29]) );
  CFD1QX1 \mult_x_1/clk_r_REG302_S1  ( .D(\mult_x_1/n1675 ), .CP(CLK), .Q(
        n2836) );
  CFD1QX4 \mult_x_1/clk_r_REG11_S2  ( .D(\mult_x_1/n149 ), .CP(CLK), .Q(n2635)
         );
  CFD1QX2 clk_r_REG4_S2 ( .D(n2887), .CP(CLK), .Q(PRODUCT[32]) );
  CFD1QX2 clk_r_REG321_S1 ( .D(n2912), .CP(CLK), .Q(n2859) );
  CFD1QX2 clk_r_REG318_S1 ( .D(n2911), .CP(CLK), .Q(n2861) );
  CFD1QX2 \mult_x_1/clk_r_REG167_S1  ( .D(\mult_x_1/n881 ), .CP(CLK), .Q(n2665) );
  CFD1QX2 \mult_x_1/clk_r_REG279_S1  ( .D(\mult_x_1/n1447 ), .CP(CLK), .Q(
        n2784) );
  CFD1QX2 \mult_x_1/clk_r_REG224_S1  ( .D(\mult_x_1/n1423 ), .CP(CLK), .Q(
        n2779) );
  CFD1QX2 \mult_x_1/clk_r_REG308_S1  ( .D(\mult_x_1/n1685 ), .CP(CLK), .Q(
        n2839) );
  CFD1QX2 \mult_x_1/clk_r_REG177_S1  ( .D(\mult_x_1/n1113 ), .CP(CLK), .Q(
        n2715) );
  CFD1QX2 \mult_x_1/clk_r_REG210_S1  ( .D(\mult_x_1/n1367 ), .CP(CLK), .Q(
        n2766) );
  CFD1QX2 \mult_x_1/clk_r_REG87_S1  ( .D(\mult_x_1/n1226 ), .CP(CLK), .Q(n2739) );
  CFD1QX2 \mult_x_1/clk_r_REG269_S1  ( .D(\mult_x_1/n1587 ), .CP(CLK), .Q(
        n2814) );
  CFD1QXL \mult_x_1/clk_r_REG116_S2  ( .D(\mult_x_1/n283 ), .CP(CLK), .Q(n2574) );
  CFD1QX1 \mult_x_1/clk_r_REG182_S1  ( .D(\mult_x_1/n1311 ), .CP(CLK), .Q(
        n2755) );
  CFD1QX2 \mult_x_1/clk_r_REG244_S1  ( .D(\mult_x_1/n1468 ), .CP(CLK), .Q(
        n2787) );
  CFD1QX2 \mult_x_1/clk_r_REG242_S1  ( .D(\mult_x_1/n1444 ), .CP(CLK), .Q(
        n2782) );
  CFD1QX1 \mult_x_1/clk_r_REG63_S1  ( .D(\mult_x_1/n1065 ), .CP(CLK), .Q(n2705) );
  CFD1QXL \mult_x_1/clk_r_REG105_S2  ( .D(\mult_x_1/n162 ), .CP(CLK), .Q(n2584) );
  CFD1QX2 \mult_x_1/clk_r_REG278_S1  ( .D(\mult_x_1/n1589 ), .CP(CLK), .Q(
        n2815) );
  CFD1QX2 \mult_x_1/clk_r_REG255_S1  ( .D(\mult_x_1/n1509 ), .CP(CLK), .Q(
        n2797) );
  CFD1QX2 \mult_x_1/clk_r_REG274_S1  ( .D(\mult_x_1/n1599 ), .CP(CLK), .Q(
        n2817) );
  CFD1QX2 \mult_x_1/clk_r_REG25_S1  ( .D(\mult_x_1/n1253 ), .CP(CLK), .Q(n2743) );
  CFD1QX2 \mult_x_1/clk_r_REG29_S1  ( .D(\mult_x_1/n1223 ), .CP(CLK), .Q(n2736) );
  CFD1QX2 \mult_x_1/clk_r_REG84_S1  ( .D(\mult_x_1/n1167 ), .CP(CLK), .Q(n2725) );
  CFD1QX2 \mult_x_1/clk_r_REG235_S1  ( .D(\mult_x_1/n1471 ), .CP(CLK), .Q(
        n2789) );
  CFD1QX4 \mult_x_1/clk_r_REG256_S1  ( .D(\mult_x_1/n1490 ), .CP(CLK), .Q(
        n2794) );
  CFD1QX2 \mult_x_1/clk_r_REG314_S1  ( .D(\mult_x_1/n696 ), .CP(CLK), .Q(n2609) );
  CFD1QX2 \mult_x_1/clk_r_REG284_S1  ( .D(\mult_x_1/n1629 ), .CP(CLK), .Q(
        n2824) );
  CFD1QX2 \mult_x_1/clk_r_REG10_S2  ( .D(\mult_x_1/n486 ), .CP(CLK), .Q(n2625)
         );
  CFD1QX2 \mult_x_1/clk_r_REG9_S2  ( .D(\mult_x_1/n495 ), .CP(CLK), .Q(n2626)
         );
  CFD1QX2 \mult_x_1/clk_r_REG8_S2  ( .D(\mult_x_1/n506 ), .CP(CLK), .Q(n2627)
         );
  CFD1QX1 \mult_x_1/clk_r_REG312_S1  ( .D(\mult_x_1/n697 ), .CP(CLK), .Q(n2610) );
  CFD1QX2 \mult_x_1/clk_r_REG230_S1  ( .D(\mult_x_1/n1419 ), .CP(CLK), .Q(
        n2776) );
  CIVX3 U1 ( .A(n1829), .Z(n5) );
  CND2X1 U2 ( .A(n1434), .B(n1433), .Z(\mult_x_1/n697 ) );
  CENXL U3 ( .A(n1289), .B(n1965), .Z(n634) );
  CENXL U4 ( .A(n1289), .B(n1630), .Z(n1572) );
  CENXL U5 ( .A(n1289), .B(n1847), .Z(n1221) );
  CENXL U6 ( .A(n1289), .B(n1969), .Z(n1505) );
  CENXL U7 ( .A(n1289), .B(n1712), .Z(n1251) );
  CENXL U8 ( .A(n1289), .B(n1707), .Z(n1640) );
  CENXL U9 ( .A(n1289), .B(n1466), .Z(n472) );
  CENXL U10 ( .A(n1289), .B(n1699), .Z(n1222) );
  CENXL U11 ( .A(n1289), .B(n1720), .Z(n1392) );
  CND2X4 U12 ( .A(n299), .B(n298), .Z(n6) );
  CND2X2 U13 ( .A(n299), .B(n298), .Z(n1926) );
  CENXL U14 ( .A(n1289), .B(n1687), .Z(n588) );
  CNIVX8 U15 ( .A(n404), .Z(n2434) );
  CENX2 U16 ( .A(n2470), .B(n1811), .Z(n1508) );
  CENX2 U17 ( .A(n2470), .B(n1961), .Z(n1509) );
  CAOR1XL U18 ( .A(n2051), .B(n2050), .C(n2049), .Z(n2351) );
  COND2XL U19 ( .A(n2050), .B(n344), .C(n1967), .D(n708), .Z(n719) );
  CND2X4 U20 ( .A(n284), .B(n1834), .Z(n7) );
  CIVX12 U21 ( .A(n552), .Z(n1973) );
  CIVX4 U22 ( .A(n550), .Z(n552) );
  CEOX2 U23 ( .A(n183), .B(n184), .Z(n1901) );
  CIVX2 U24 ( .A(n953), .Z(n10) );
  CEOX4 U25 ( .A(A[10]), .B(n1704), .Z(n297) );
  CENX2 U26 ( .A(n1838), .B(A[10]), .Z(n296) );
  CENX2 U27 ( .A(n540), .B(n539), .Z(n587) );
  CENX1 U28 ( .A(n1040), .B(n126), .Z(n2887) );
  CENXL U29 ( .A(n1966), .B(n1965), .Z(n2049) );
  CENXL U30 ( .A(n1966), .B(n1699), .Z(n1473) );
  CENXL U31 ( .A(n1966), .B(n1630), .Z(n1524) );
  CNIVX2 U32 ( .A(n2434), .Z(n243) );
  CND2X2 U33 ( .A(n312), .B(n311), .Z(n8) );
  CND2X2 U34 ( .A(n312), .B(n311), .Z(n9) );
  CND2XL U35 ( .A(n312), .B(n311), .Z(n2524) );
  COAN1XL U36 ( .A(n952), .B(n12), .C(n10), .Z(n954) );
  CIVXL U37 ( .A(n952), .Z(n1914) );
  CIVX8 U38 ( .A(n264), .Z(n1924) );
  CNR2X1 U39 ( .A(n1434), .B(n1433), .Z(\mult_x_1/n696 ) );
  CNIVX4 U40 ( .A(B[28]), .Z(n2469) );
  CNR2IX4 U41 ( .B(n1714), .A(n2406), .Z(n1379) );
  COND2X2 U42 ( .A(n2436), .B(n405), .C(n2434), .D(n1500), .Z(n1421) );
  COND2XL U43 ( .A(n8), .B(n2442), .C(n2522), .D(n740), .Z(n688) );
  COND2XL U44 ( .A(n8), .B(n2005), .C(n2522), .D(n1980), .Z(n2267) );
  COND2X2 U45 ( .A(n255), .B(n1865), .C(n2388), .D(n1364), .Z(n2322) );
  CIVX8 U46 ( .A(n270), .Z(n11) );
  CIVX3 U47 ( .A(n270), .Z(n1832) );
  COND2X2 U48 ( .A(n2004), .B(n1558), .C(n2002), .D(n1223), .Z(n1240) );
  CANR1X2 U49 ( .A(n2029), .B(n75), .C(n76), .Z(n12) );
  CANR1X1 U50 ( .A(n2029), .B(n75), .C(n76), .Z(n266) );
  CIVX4 U51 ( .A(A[3]), .Z(n579) );
  CND2X2 U52 ( .A(n310), .B(n1842), .Z(n13) );
  CND2X2 U53 ( .A(n310), .B(n1842), .Z(n14) );
  CNIVXL U54 ( .A(n388), .Z(n15) );
  CND2X2 U55 ( .A(n310), .B(n1842), .Z(n2055) );
  CIVX12 U56 ( .A(n921), .Z(n1829) );
  CIVX8 U57 ( .A(n1716), .Z(n2395) );
  CIVX4 U58 ( .A(n1716), .Z(n1970) );
  CNIVX4 U59 ( .A(n313), .Z(n2522) );
  CENX2 U60 ( .A(A[23]), .B(A[24]), .Z(n313) );
  COND2XL U61 ( .A(n1815), .B(n1415), .C(n2002), .D(n1504), .Z(n2056) );
  CIVDX3 U62 ( .A(n371), .Z0(n1692) );
  CENXL U63 ( .A(n1738), .B(n151), .Z(n153) );
  CANR5CX1 U64 ( .A(n1376), .B(n80), .C(n81), .Z(n82) );
  COND2X1 U65 ( .A(n2398), .B(n1351), .C(n2392), .D(n1352), .Z(n81) );
  CENX2 U66 ( .A(n1387), .B(n1707), .Z(n640) );
  CIVXL U67 ( .A(n260), .Z(n16) );
  COND2X1 U68 ( .A(n2406), .B(n1565), .C(n2436), .D(n1393), .Z(n187) );
  CIVX2 U69 ( .A(n188), .Z(n1810) );
  CEOX2 U70 ( .A(A[22]), .B(A[23]), .Z(n320) );
  CEOX2 U71 ( .A(A[14]), .B(n1848), .Z(n17) );
  CENXL U72 ( .A(n136), .B(n123), .Z(n497) );
  CIVX3 U73 ( .A(n343), .Z(n18) );
  CIVX4 U74 ( .A(n343), .Z(n1880) );
  CENXL U75 ( .A(n186), .B(n79), .Z(n2285) );
  CIVXL U76 ( .A(n361), .Z(n19) );
  CIVXL U77 ( .A(n19), .Z(n20) );
  CANR1X2 U78 ( .A(n268), .B(n275), .C(n945), .Z(n2535) );
  CENXL U79 ( .A(n1387), .B(n1965), .Z(n244) );
  CAN2XL U80 ( .A(n147), .B(n148), .Z(n2179) );
  CENX2 U81 ( .A(n1387), .B(n1965), .Z(n1818) );
  CNIVX2 U82 ( .A(n1692), .Z(n21) );
  CNIVX2 U83 ( .A(n1692), .Z(n22) );
  CNIVX1 U84 ( .A(n1692), .Z(n1690) );
  CEOX4 U85 ( .A(A[8]), .B(n1838), .Z(n299) );
  COND2X1 U86 ( .A(n2233), .B(n1444), .C(n1834), .D(n1747), .Z(n1538) );
  CNIVX3 U87 ( .A(n2636), .Z(n24) );
  CNIVX1 U88 ( .A(n24), .Z(n23) );
  CNIVX1 U89 ( .A(n31), .Z(n25) );
  CNIVX3 U90 ( .A(n2632), .Z(n27) );
  CNIVX1 U91 ( .A(n27), .Z(n26) );
  CNIVX1 U92 ( .A(n2569), .Z(n28) );
  CNIVX1 U93 ( .A(n278), .Z(n29) );
  CNIVX1 U94 ( .A(\mult_x_1/n153 ), .Z(n30) );
  CNIVX1 U95 ( .A(n2550), .Z(n31) );
  CNIVX1 U96 ( .A(n280), .Z(n32) );
  CNIVX1 U97 ( .A(n1107), .Z(n33) );
  CNIVX3 U98 ( .A(n2841), .Z(n35) );
  CNIVX1 U99 ( .A(n35), .Z(n34) );
  CNIVX1 U100 ( .A(n1109), .Z(n36) );
  CNIVX1 U101 ( .A(n281), .Z(n37) );
  CNIVX3 U102 ( .A(n2847), .Z(n39) );
  CNIVX1 U103 ( .A(n39), .Z(n38) );
  CNIVX3 U104 ( .A(n2851), .Z(n41) );
  CNIVX1 U105 ( .A(n41), .Z(n40) );
  CNIVX3 U106 ( .A(n2849), .Z(n43) );
  CNIVX1 U107 ( .A(n43), .Z(n42) );
  CNIVX3 U108 ( .A(n2857), .Z(n45) );
  CNIVX1 U109 ( .A(n45), .Z(n44) );
  CNIVX3 U110 ( .A(n2855), .Z(n47) );
  CNIVX1 U111 ( .A(n47), .Z(n46) );
  CNIVX3 U112 ( .A(n2853), .Z(n49) );
  CNIVX1 U113 ( .A(n49), .Z(n48) );
  CNIVX1 U114 ( .A(n51), .Z(n50) );
  CNIVX1 U115 ( .A(n52), .Z(n51) );
  CNIVX1 U116 ( .A(n53), .Z(n52) );
  CNIVX1 U117 ( .A(n2861), .Z(n53) );
  CNIVX1 U118 ( .A(n55), .Z(n54) );
  CNIVX1 U119 ( .A(n56), .Z(n55) );
  CNIVX1 U120 ( .A(n57), .Z(n56) );
  CNIVX1 U121 ( .A(n2859), .Z(n57) );
  CNIVX1 U122 ( .A(n2909), .Z(n58) );
  CNIVX1 U123 ( .A(n282), .Z(n59) );
  CENX1 U124 ( .A(n1387), .B(n1464), .Z(n654) );
  CENX1 U125 ( .A(n1387), .B(n1466), .Z(n933) );
  COND1XL U126 ( .A(n2483), .B(n893), .C(n2482), .Z(n1011) );
  COAN1X1 U127 ( .A(n2537), .B(n823), .C(n2033), .Z(n2030) );
  CNR2X1 U128 ( .A(n947), .B(n946), .Z(n2532) );
  CIVX4 U129 ( .A(n238), .Z(n239) );
  CIVX2 U130 ( .A(n2509), .Z(n238) );
  CND2X1 U131 ( .A(n1426), .B(n1425), .Z(n1427) );
  CND2X1 U132 ( .A(n273), .B(n2412), .Z(n137) );
  CANR5CXL U133 ( .A(n342), .B(n340), .C(n339), .Z(n167) );
  CND2XL U134 ( .A(n574), .B(n572), .Z(n433) );
  COND1XL U135 ( .A(n572), .B(n574), .C(n571), .Z(n434) );
  CND2XL U136 ( .A(n366), .B(n365), .Z(\mult_x_1/n1674 ) );
  CND2XL U137 ( .A(n370), .B(n367), .Z(n365) );
  COND1XL U138 ( .A(n367), .B(n370), .C(n368), .Z(n366) );
  CND2XL U139 ( .A(n1003), .B(n2557), .Z(n60) );
  CANR1XL U140 ( .A(n1004), .B(n2557), .C(n2558), .Z(n61) );
  COND1XL U141 ( .A(n2635), .B(n60), .C(n61), .Z(n62) );
  CENX1 U142 ( .A(n2580), .B(n62), .Z(PRODUCT[53]) );
  CANR5CXL U143 ( .A(n95), .B(n96), .C(n939), .Z(n63) );
  CIVX1 U144 ( .A(n63), .Z(n946) );
  CNR2X1 U145 ( .A(n2511), .B(n2609), .Z(n64) );
  COND1XL U146 ( .A(n2511), .B(n2610), .C(n2512), .Z(n65) );
  CANR1X1 U147 ( .A(n2513), .B(n64), .C(n65), .Z(n728) );
  CENX1 U148 ( .A(n809), .B(n807), .Z(n66) );
  CENXL U149 ( .A(n808), .B(n66), .Z(n825) );
  COND2X1 U150 ( .A(n1603), .B(n2510), .C(n2509), .D(n591), .Z(n67) );
  COND2XL U151 ( .A(n2430), .B(n590), .C(n2432), .D(n588), .Z(n68) );
  CENX1 U152 ( .A(n1186), .B(n67), .Z(n69) );
  CENX1 U153 ( .A(n68), .B(n69), .Z(n1197) );
  CANR5CX1 U154 ( .A(n1186), .B(n67), .C(n68), .Z(n70) );
  CIVX1 U155 ( .A(n70), .Z(n1517) );
  CIVXL U156 ( .A(n431), .Z(n71) );
  CIVXL U157 ( .A(n432), .Z(n72) );
  CANR5CX1 U158 ( .A(n2418), .B(n71), .C(n72), .Z(n340) );
  CANR5CX1 U159 ( .A(n316), .B(n318), .C(n315), .Z(n73) );
  CIVXL U160 ( .A(n73), .Z(\mult_x_1/n1088 ) );
  CENXL U161 ( .A(n254), .B(n1711), .Z(n74) );
  COND2X1 U162 ( .A(n2434), .B(n1682), .C(n245), .D(n74), .Z(n147) );
  CNR2X1 U163 ( .A(n830), .B(n2543), .Z(n75) );
  COND1X2 U164 ( .A(n830), .B(n2030), .C(n829), .Z(n76) );
  CIVXL U165 ( .A(n1533), .Z(n77) );
  CANR4CXL U166 ( .A(n18), .B(n1714), .C(n248), .D(n77), .Z(n580) );
  CANR5CXL U167 ( .A(n114), .B(n805), .C(n804), .Z(n78) );
  CIVX1 U168 ( .A(n78), .Z(n831) );
  CENXL U169 ( .A(n2284), .B(n187), .Z(n79) );
  COND2X1 U170 ( .A(n1884), .B(n1349), .C(n1886), .D(n1350), .Z(n80) );
  CIVX1 U171 ( .A(n82), .Z(n1953) );
  CENXL U172 ( .A(n1376), .B(n81), .Z(n83) );
  CENX1 U173 ( .A(n80), .B(n83), .Z(n1374) );
  CEOX1 U174 ( .A(n431), .B(n2418), .Z(n84) );
  CENX1 U175 ( .A(n432), .B(n84), .Z(n571) );
  CENXL U176 ( .A(n129), .B(n924), .Z(n85) );
  CENXL U177 ( .A(n925), .B(n85), .Z(n947) );
  CANR5CX1 U178 ( .A(n865), .B(n867), .C(n866), .Z(n86) );
  CIVX2 U179 ( .A(n86), .Z(n891) );
  COND2XL U180 ( .A(n1884), .B(n936), .C(n1886), .D(n578), .Z(n87) );
  CENX1 U181 ( .A(n1711), .B(n1533), .Z(n88) );
  COND2XL U182 ( .A(n1857), .B(n88), .C(n1880), .D(n934), .Z(n89) );
  CEOXL U183 ( .A(n87), .B(n89), .Z(n581) );
  CAN2XL U184 ( .A(n87), .B(n89), .Z(n937) );
  CIVXL U185 ( .A(n2635), .Z(n90) );
  CANR1XL U186 ( .A(n991), .B(n90), .C(n992), .Z(n91) );
  CEOX1 U187 ( .A(n2570), .B(n91), .Z(PRODUCT[59]) );
  CNR2IXL U188 ( .B(n1017), .A(n2467), .Z(n1021) );
  CENX1 U189 ( .A(n120), .B(n121), .Z(n92) );
  CENX1 U190 ( .A(n418), .B(n92), .Z(n1133) );
  CAN2X1 U191 ( .A(n824), .B(n825), .Z(n2544) );
  CENXL U192 ( .A(n1711), .B(n1973), .Z(n93) );
  COND2X1 U193 ( .A(n2004), .B(n93), .C(n2002), .D(n1439), .Z(n183) );
  COND1X1 U194 ( .A(n870), .B(n869), .C(n868), .Z(n94) );
  CND2X1 U195 ( .A(n94), .B(n693), .Z(n694) );
  COND2XL U196 ( .A(n18), .B(n929), .C(n1857), .D(n933), .Z(n95) );
  COND2XL U197 ( .A(n1884), .B(n926), .C(n1886), .D(n935), .Z(n96) );
  CENX1 U198 ( .A(n939), .B(n95), .Z(n97) );
  CENX1 U199 ( .A(n96), .B(n97), .Z(n944) );
  CND2X1 U200 ( .A(n676), .B(n678), .Z(n98) );
  CND2XL U201 ( .A(n676), .B(n677), .Z(n99) );
  COND3X1 U202 ( .A(n674), .B(n98), .C(n675), .D(n99), .Z(n682) );
  CIVXL U203 ( .A(n2635), .Z(n100) );
  CND2XL U204 ( .A(n1207), .B(n1206), .Z(n101) );
  CND2X1 U205 ( .A(n101), .B(n1205), .Z(n102) );
  CANR11X1 U206 ( .A(n1204), .B(n1207), .C(n100), .D(n102), .Z(PRODUCT[63]) );
  CNR2XL U207 ( .A(n1035), .B(n2481), .Z(n103) );
  CND2XL U208 ( .A(n1036), .B(n103), .Z(n1034) );
  COR2X1 U209 ( .A(n825), .B(n824), .Z(n2545) );
  COND1XL U210 ( .A(n2635), .B(n2585), .C(n2619), .Z(n104) );
  CENX1 U211 ( .A(n2584), .B(n104), .Z(PRODUCT[50]) );
  CENX1 U212 ( .A(n879), .B(n880), .Z(n105) );
  CENX1 U213 ( .A(n878), .B(n105), .Z(n695) );
  CENX1 U214 ( .A(n866), .B(n867), .Z(n106) );
  CENX1 U215 ( .A(n865), .B(n106), .Z(n890) );
  COND2X1 U216 ( .A(n8), .B(n1344), .C(n2522), .D(n1343), .Z(n107) );
  COND2X1 U217 ( .A(n8), .B(n1346), .C(n2522), .D(n1345), .Z(n108) );
  CAN2X1 U218 ( .A(n107), .B(n108), .Z(n2320) );
  CEOX1 U219 ( .A(n107), .B(n108), .Z(n1852) );
  CNR2IXL U220 ( .B(n1057), .A(n1059), .Z(n1061) );
  CANR5CXL U221 ( .A(n129), .B(n925), .C(n924), .Z(n109) );
  CIVXL U222 ( .A(n109), .Z(n922) );
  CND2X1 U223 ( .A(n2505), .B(n727), .Z(n110) );
  CND2XL U224 ( .A(n727), .B(n729), .Z(n111) );
  COND3X1 U225 ( .A(n728), .B(n110), .C(n726), .D(n111), .Z(n697) );
  CANR5CXL U226 ( .A(n2809), .B(n521), .C(n520), .Z(n112) );
  CIVX1 U227 ( .A(n112), .Z(n528) );
  CENX1 U228 ( .A(n2773), .B(n2771), .Z(n113) );
  CENX1 U229 ( .A(n792), .B(n113), .Z(n114) );
  CENX1 U230 ( .A(n804), .B(n805), .Z(n115) );
  CENX1 U231 ( .A(n114), .B(n115), .Z(n827) );
  CIVXL U232 ( .A(n2635), .Z(n116) );
  CANR1XL U233 ( .A(n1204), .B(n116), .C(n1206), .Z(n117) );
  CND2X1 U234 ( .A(n1207), .B(n1205), .Z(n118) );
  CEOX1 U235 ( .A(n117), .B(n118), .Z(PRODUCT[62]) );
  CANR5CXL U236 ( .A(n133), .B(n132), .C(n1739), .Z(n119) );
  CIVX1 U237 ( .A(n119), .Z(n1484) );
  COND2X1 U238 ( .A(n329), .B(n2510), .C(n2509), .D(n332), .Z(n120) );
  COND2X1 U239 ( .A(n2398), .B(n330), .C(n2392), .D(n419), .Z(n121) );
  CANR5CXL U240 ( .A(n418), .B(n120), .C(n121), .Z(n122) );
  CIVXL U241 ( .A(n122), .Z(n432) );
  CANR5CX1 U242 ( .A(n538), .B(n537), .C(n540), .Z(n123) );
  CIVXL U243 ( .A(n123), .Z(n495) );
  CND2XL U244 ( .A(n1171), .B(n1169), .Z(n124) );
  CND3X1 U245 ( .A(n124), .B(n259), .C(n258), .Z(n201) );
  CIVX1 U246 ( .A(n2500), .Z(n125) );
  CANR1X1 U247 ( .A(n2501), .B(n2502), .C(n125), .Z(n932) );
  CNR2IXL U248 ( .B(n1029), .A(n1030), .Z(n126) );
  CND2IXL U249 ( .B(n2467), .A(n2468), .Z(\mult_x_1/n174 ) );
  COND1XL U250 ( .A(n2032), .B(n2542), .C(n2537), .Z(n127) );
  CND2XL U251 ( .A(n2033), .B(n2034), .Z(n128) );
  CENX1 U252 ( .A(n127), .B(n128), .Z(n2894) );
  CND2IX1 U253 ( .B(n1052), .A(n1061), .Z(n1064) );
  COND2XL U254 ( .A(n1861), .B(n914), .C(n1893), .D(n918), .Z(n129) );
  COND1XL U255 ( .A(n2635), .B(n2588), .C(n2620), .Z(n130) );
  CENXL U256 ( .A(n2587), .B(n130), .Z(PRODUCT[48]) );
  CIVXL U257 ( .A(n960), .Z(n131) );
  COND1X1 U258 ( .A(n962), .B(n131), .C(n961), .Z(n963) );
  COND2X1 U259 ( .A(n1893), .B(n1521), .C(n241), .D(n1474), .Z(n132) );
  COND2XL U260 ( .A(n246), .B(n1524), .C(n2051), .D(n1473), .Z(n133) );
  CENX1 U261 ( .A(n1739), .B(n132), .Z(n134) );
  CENX1 U262 ( .A(n133), .B(n134), .Z(n1754) );
  CENXL U263 ( .A(n158), .B(n427), .Z(n135) );
  CENX1 U264 ( .A(n1589), .B(n135), .Z(n1593) );
  CANR5CXL U265 ( .A(n536), .B(n534), .C(n535), .Z(n136) );
  CIVXL U266 ( .A(n136), .Z(n496) );
  CND2X2 U267 ( .A(n137), .B(n2411), .Z(n268) );
  CND2IXL U268 ( .B(n897), .A(n896), .Z(\mult_x_1/n175 ) );
  CND2XL U269 ( .A(n1023), .B(n1021), .Z(n138) );
  CANR1XL U270 ( .A(n1025), .B(n1021), .C(n1020), .Z(n139) );
  COND1XL U271 ( .A(n1028), .B(n138), .C(n139), .Z(\mult_x_1/n486 ) );
  CANR5CXL U272 ( .A(n201), .B(n1182), .C(n1181), .Z(n140) );
  CIVXL U273 ( .A(n140), .Z(\mult_x_1/n1486 ) );
  COND1XL U274 ( .A(n2491), .B(n2490), .C(n2489), .Z(n141) );
  CND2IX1 U275 ( .B(n2492), .A(n2493), .Z(n142) );
  CENX1 U276 ( .A(n141), .B(n142), .Z(n2905) );
  COND1XL U277 ( .A(n2464), .B(n2463), .C(n2462), .Z(n143) );
  CND2IXL U278 ( .B(n2465), .A(n2466), .Z(n144) );
  CENX1 U279 ( .A(n143), .B(n144), .Z(n2899) );
  COND1XL U280 ( .A(n2542), .B(n2543), .C(n2541), .Z(n145) );
  CND2IXL U281 ( .B(n2544), .A(n2545), .Z(n146) );
  CENX1 U282 ( .A(n145), .B(n146), .Z(n2893) );
  COND2X1 U283 ( .A(n1684), .B(n245), .C(n2434), .D(n1683), .Z(n148) );
  CEOX1 U284 ( .A(n147), .B(n148), .Z(n2246) );
  COND1X1 U285 ( .A(n2635), .B(n2563), .C(n2564), .Z(n149) );
  CENX1 U286 ( .A(n2591), .B(n149), .Z(PRODUCT[46]) );
  COND1XL U287 ( .A(n2635), .B(n2583), .C(n2618), .Z(n150) );
  CENX1 U288 ( .A(n2582), .B(n150), .Z(PRODUCT[51]) );
  CNR2IXL U289 ( .B(n959), .A(n962), .Z(n964) );
  COND2XL U290 ( .A(n1884), .B(n1471), .C(n1886), .D(n1526), .Z(n151) );
  COND2XL U291 ( .A(n1842), .B(n1469), .C(n14), .D(n1744), .Z(n152) );
  CENX1 U292 ( .A(n152), .B(n153), .Z(n1755) );
  CANR5CXL U293 ( .A(n1738), .B(n151), .C(n152), .Z(n154) );
  CIVX1 U294 ( .A(n154), .Z(n1485) );
  CANR5CXL U295 ( .A(n219), .B(n220), .C(n2331), .Z(n155) );
  CIVXL U296 ( .A(n155), .Z(n2336) );
  CNR2X1 U297 ( .A(n263), .B(n1497), .Z(n156) );
  CNR2XL U298 ( .A(n2522), .B(n424), .Z(n157) );
  CNR2X1 U299 ( .A(n156), .B(n157), .Z(n158) );
  CIVX2 U300 ( .A(n1589), .Z(n159) );
  CANR5CX1 U301 ( .A(n427), .B(n158), .C(n159), .Z(n1136) );
  CENX1 U302 ( .A(n218), .B(n1590), .Z(n160) );
  CENX1 U303 ( .A(n1591), .B(n160), .Z(n1513) );
  COR2X1 U304 ( .A(n922), .B(n923), .Z(n1015) );
  CANR1XL U305 ( .A(n1025), .B(n1017), .C(n1018), .Z(n161) );
  CND2XL U306 ( .A(n1017), .B(n1023), .Z(n162) );
  COND1XL U307 ( .A(n1028), .B(n162), .C(n161), .Z(\mult_x_1/n495 ) );
  CANR5CX1 U308 ( .A(n585), .B(n587), .C(n584), .Z(n163) );
  CIVXL U309 ( .A(n163), .Z(\mult_x_1/n1310 ) );
  CIVXL U310 ( .A(n1056), .Z(n164) );
  CANR1XL U311 ( .A(n1067), .B(n1053), .C(n164), .Z(\mult_x_1/n406 ) );
  CNR2X1 U312 ( .A(n1108), .B(n1109), .Z(n165) );
  CANR1XL U313 ( .A(n2549), .B(n1107), .C(n165), .Z(n166) );
  COND3XL U314 ( .A(n1110), .B(n1112), .C(n166), .D(n28), .Z(\mult_x_1/n236 )
         );
  CIVXL U315 ( .A(n167), .Z(\mult_x_1/n868 ) );
  CENX1 U316 ( .A(n1181), .B(n1182), .Z(n168) );
  CENXL U317 ( .A(n201), .B(n168), .Z(\mult_x_1/n1487 ) );
  CNR2IXL U318 ( .B(n2610), .A(n2609), .Z(n169) );
  CENX1 U319 ( .A(n2514), .B(n169), .Z(n2910) );
  CANR1XL U320 ( .A(n2505), .B(n2507), .C(n729), .Z(n170) );
  CND2XL U321 ( .A(n727), .B(n726), .Z(n171) );
  CEOX1 U322 ( .A(n170), .B(n171), .Z(n2907) );
  CND2XL U323 ( .A(n2495), .B(n2494), .Z(n172) );
  CENX1 U324 ( .A(n2496), .B(n172), .Z(n2904) );
  CND2XL U325 ( .A(n2547), .B(n2546), .Z(n173) );
  CENX1 U326 ( .A(n2548), .B(n173), .Z(n2898) );
  CANR1XL U327 ( .A(n2540), .B(n2545), .C(n2544), .Z(n174) );
  CND2XL U328 ( .A(n2545), .B(n2028), .Z(n175) );
  COND1XL U329 ( .A(n2542), .B(n175), .C(n174), .Z(n176) );
  CND2XL U330 ( .A(n828), .B(n267), .Z(n177) );
  CENX1 U331 ( .A(n176), .B(n177), .Z(n2892) );
  CANR1XL U332 ( .A(n1004), .B(n2579), .C(n2617), .Z(n178) );
  CND2XL U333 ( .A(n1003), .B(n2579), .Z(n179) );
  COND1XL U334 ( .A(n2635), .B(n179), .C(n178), .Z(n180) );
  CENX1 U335 ( .A(n2578), .B(n180), .Z(PRODUCT[54]) );
  CIVXL U336 ( .A(n2576), .Z(n181) );
  CANR1XL U337 ( .A(n2616), .B(n2556), .C(n181), .Z(n978) );
  CANR5CXL U338 ( .A(n879), .B(n880), .C(n878), .Z(n182) );
  CIVXL U339 ( .A(n182), .Z(n898) );
  COND2X1 U340 ( .A(n2002), .B(n551), .C(n552), .D(n1815), .Z(n184) );
  CAN2X1 U341 ( .A(n183), .B(n184), .Z(n2086) );
  CIVX1 U342 ( .A(n1050), .Z(n185) );
  CANR1X1 U343 ( .A(n1051), .B(n1113), .C(n185), .Z(n1080) );
  COND2X1 U344 ( .A(n2430), .B(n1573), .C(n2310), .D(n1392), .Z(n186) );
  CANR5CX1 U345 ( .A(n2284), .B(n186), .C(n187), .Z(n188) );
  CNR2IX1 U346 ( .B(n1714), .A(n1967), .Z(n189) );
  COND2XL U347 ( .A(n1884), .B(n350), .C(n1886), .D(n658), .Z(n190) );
  CENX1 U348 ( .A(n189), .B(n361), .Z(n191) );
  CENX1 U349 ( .A(n190), .B(n191), .Z(n1148) );
  CANR5CXL U350 ( .A(n189), .B(n20), .C(n190), .Z(n192) );
  CIVX1 U351 ( .A(n192), .Z(n1143) );
  CANR5CXL U352 ( .A(n218), .B(n1591), .C(n1590), .Z(n193) );
  CIVX1 U353 ( .A(n193), .Z(n1592) );
  CIVXL U354 ( .A(n2058), .Z(n194) );
  COND1XL U355 ( .A(n2059), .B(n194), .C(n1417), .Z(n195) );
  CENX1 U356 ( .A(n1510), .B(n1511), .Z(n196) );
  CENX1 U357 ( .A(n195), .B(n196), .Z(n1431) );
  CANR5CXL U358 ( .A(n1510), .B(n1511), .C(n195), .Z(n197) );
  CIVX1 U359 ( .A(n197), .Z(n1512) );
  CIVXL U360 ( .A(n21), .Z(n198) );
  COND1XL U361 ( .A(n1714), .B(n198), .C(n1886), .Z(n997) );
  CANR5CXL U362 ( .A(n498), .B(n496), .C(n495), .Z(n199) );
  CIVXL U363 ( .A(n199), .Z(\mult_x_1/n1282 ) );
  CANR5CXL U364 ( .A(n225), .B(n1686), .C(n1685), .Z(n200) );
  CIVXL U365 ( .A(n200), .Z(\mult_x_1/n1312 ) );
  CND2IXL U366 ( .B(n1055), .A(n1054), .Z(\mult_x_1/n165 ) );
  CND2XL U367 ( .A(n273), .B(n2411), .Z(n202) );
  CENX1 U368 ( .A(n2412), .B(n202), .Z(n2914) );
  CNR2IXL U369 ( .B(n2612), .A(n2611), .Z(n203) );
  CENX1 U370 ( .A(n2634), .B(n203), .Z(n282) );
  COND1XL U371 ( .A(n2609), .B(n2514), .C(n2610), .Z(n204) );
  CND2IXL U372 ( .B(n2511), .A(n2512), .Z(n205) );
  CENX1 U373 ( .A(n204), .B(n205), .Z(n2909) );
  CNR2IXL U374 ( .B(n2489), .A(n2491), .Z(n206) );
  CENX1 U375 ( .A(n2490), .B(n206), .Z(n2906) );
  CND2X1 U376 ( .A(n2495), .B(n2496), .Z(n207) );
  CND2XL U377 ( .A(n207), .B(n2494), .Z(n208) );
  CND2IXL U378 ( .B(n671), .A(n672), .Z(n209) );
  CENX1 U379 ( .A(n208), .B(n209), .Z(n2903) );
  CND2XL U380 ( .A(n2547), .B(n2548), .Z(n210) );
  CND2X1 U381 ( .A(n210), .B(n2546), .Z(n211) );
  CND2IXL U382 ( .B(n797), .A(n796), .Z(n212) );
  CENX1 U383 ( .A(n211), .B(n212), .Z(n2897) );
  COND1XL U384 ( .A(n2635), .B(n2593), .C(n2622), .Z(n213) );
  CENX1 U385 ( .A(n2592), .B(n213), .Z(PRODUCT[45]) );
  CENX1 U386 ( .A(n535), .B(n534), .Z(n214) );
  CENX1 U387 ( .A(n536), .B(n214), .Z(n585) );
  CEOX1 U388 ( .A(n2041), .B(n2037), .Z(n215) );
  CENX1 U389 ( .A(n2042), .B(n215), .Z(n1791) );
  CANR5CXL U390 ( .A(n216), .B(n2041), .C(n2042), .Z(n217) );
  CIVX1 U391 ( .A(n2037), .Z(n216) );
  CIVX1 U392 ( .A(n217), .Z(n2043) );
  COND2X1 U393 ( .A(n2398), .B(n1499), .C(n2392), .D(n1506), .Z(n218) );
  COND2X1 U394 ( .A(n1920), .B(n349), .C(n1877), .D(n707), .Z(n219) );
  COND2X1 U395 ( .A(n18), .B(n706), .C(n253), .D(n353), .Z(n220) );
  CENX1 U396 ( .A(n2331), .B(n219), .Z(n221) );
  CENX1 U397 ( .A(n220), .B(n221), .Z(n367) );
  CENX1 U398 ( .A(n409), .B(n411), .Z(n222) );
  CENX1 U399 ( .A(n410), .B(n222), .Z(\mult_x_1/n961 ) );
  CND2IX1 U400 ( .B(\mult_x_1/n460 ), .A(n1117), .Z(\mult_x_1/n451 ) );
  CND2IX1 U401 ( .B(n2487), .A(n2488), .Z(\mult_x_1/n173 ) );
  CND2IX1 U402 ( .B(n2481), .A(n2482), .Z(\mult_x_1/n177 ) );
  CND2IX1 U403 ( .B(n888), .A(n887), .Z(\mult_x_1/n179 ) );
  CND2IX1 U404 ( .B(n1095), .A(n1094), .Z(\mult_x_1/n156 ) );
  CND2IX1 U405 ( .B(n1086), .A(n1101), .Z(\mult_x_1/n159 ) );
  CND2IX1 U406 ( .B(n1059), .A(n1074), .Z(\mult_x_1/n164 ) );
  CANR5CXL U407 ( .A(n773), .B(n775), .C(n774), .Z(n223) );
  CIVX1 U408 ( .A(n223), .Z(\mult_x_1/n1042 ) );
  COND1XL U409 ( .A(n1673), .B(n1675), .C(n1674), .Z(n224) );
  CND2X1 U410 ( .A(n224), .B(n1676), .Z(n225) );
  CENX1 U411 ( .A(n1686), .B(n225), .Z(n226) );
  CENX1 U412 ( .A(n1685), .B(n226), .Z(\mult_x_1/n1313 ) );
  COND1XL U413 ( .A(n1489), .B(n1488), .C(n1487), .Z(n227) );
  CND2X1 U414 ( .A(n227), .B(n235), .Z(n228) );
  CENX1 U415 ( .A(n1494), .B(n228), .Z(n229) );
  CENX1 U416 ( .A(n1493), .B(n229), .Z(\mult_x_1/n1529 ) );
  CANR5CXL U417 ( .A(n1493), .B(n1494), .C(n228), .Z(n230) );
  CIVX1 U418 ( .A(n230), .Z(\mult_x_1/n1528 ) );
  COAN1X1 U419 ( .A(n998), .B(n997), .C(n999), .Z(n2917) );
  CEO3X2 U420 ( .A(n1483), .B(n1482), .C(n1481), .Z(n1487) );
  CEOXL U421 ( .A(n1489), .B(n1488), .Z(n231) );
  CEOXL U422 ( .A(n231), .B(n1487), .Z(\mult_x_1/n1551 ) );
  CND2XL U423 ( .A(n1483), .B(n1482), .Z(n232) );
  CND2XL U424 ( .A(n1483), .B(n1481), .Z(n233) );
  CND2X1 U425 ( .A(n1482), .B(n1481), .Z(n234) );
  CND3X1 U426 ( .A(n232), .B(n233), .C(n234), .Z(n1326) );
  CND2X1 U427 ( .A(n1489), .B(n1488), .Z(n235) );
  COR2X1 U428 ( .A(n14), .B(n1469), .Z(n236) );
  COR2XL U429 ( .A(n1842), .B(n1309), .Z(n237) );
  CND2X2 U430 ( .A(n236), .B(n237), .Z(n1481) );
  CENXL U431 ( .A(n1975), .B(n1701), .Z(n1469) );
  CENXL U432 ( .A(n1975), .B(n1630), .Z(n1309) );
  COND2XL U433 ( .A(n1857), .B(n485), .C(n18), .D(n1283), .Z(n1798) );
  CNIVXL U434 ( .A(n1891), .Z(n240) );
  CNIVX4 U435 ( .A(n1891), .Z(n241) );
  CNIVX2 U436 ( .A(n1891), .Z(n242) );
  CENX1 U437 ( .A(n354), .B(A[4]), .Z(n1891) );
  COND2X2 U438 ( .A(n1886), .B(n1282), .C(n1884), .D(n1288), .Z(n1647) );
  CIVX4 U439 ( .A(A[1]), .Z(n371) );
  CANR1X1 U440 ( .A(n960), .B(n840), .C(n839), .Z(n841) );
  CHA1XL U441 ( .A(n1538), .B(n1537), .CO(n1545), .S(n2076) );
  CNIVX20 U442 ( .A(n354), .Z(n1387) );
  CIVX2 U443 ( .A(n2532), .Z(n2534) );
  CENX2 U444 ( .A(n291), .B(A[16]), .Z(n283) );
  CND2X2 U445 ( .A(n286), .B(n404), .Z(n245) );
  CND2X2 U446 ( .A(n286), .B(n404), .Z(n2436) );
  CND2X2 U447 ( .A(n297), .B(n296), .Z(n246) );
  CND2X2 U448 ( .A(n297), .B(n296), .Z(n2050) );
  CNIVX4 U449 ( .A(A[5]), .Z(n247) );
  CNIVX1 U450 ( .A(n1857), .Z(n248) );
  CENX1 U451 ( .A(A[24]), .B(n319), .Z(n312) );
  CIVX8 U452 ( .A(n319), .Z(n1632) );
  CENX2 U453 ( .A(n1161), .B(A[22]), .Z(n249) );
  CIVX8 U454 ( .A(n249), .Z(n292) );
  CIVDX3 U455 ( .A(A[21]), .Z0(n1161), .Z1(n2390) );
  CIVX8 U456 ( .A(n579), .Z(n354) );
  CENX2 U457 ( .A(n354), .B(A[4]), .Z(n351) );
  CNIVX3 U458 ( .A(n354), .Z(n1533) );
  CANR1X1 U459 ( .A(n682), .B(n531), .C(n530), .Z(n802) );
  COND1X1 U460 ( .A(n2465), .B(n2462), .C(n2466), .Z(n530) );
  CND2XL U461 ( .A(n808), .B(n807), .Z(n250) );
  CND2X1 U462 ( .A(n808), .B(n809), .Z(n251) );
  CND2XL U463 ( .A(n807), .B(n809), .Z(n252) );
  CND3XL U464 ( .A(n250), .B(n251), .C(n252), .Z(n826) );
  CANR1X1 U465 ( .A(n2544), .B(n267), .C(n2031), .Z(n829) );
  CNIVXL U466 ( .A(n248), .Z(n253) );
  CEOX2 U467 ( .A(n319), .B(A[26]), .Z(n314) );
  CNIVX4 U468 ( .A(n313), .Z(n311) );
  CIVXL U469 ( .A(n1786), .Z(n1574) );
  CAOR1X1 U470 ( .A(n1834), .B(n7), .C(n417), .Z(n423) );
  CEOX4 U471 ( .A(A[16]), .B(n1977), .Z(n284) );
  CIVX8 U472 ( .A(n1684), .Z(n254) );
  CEOX2 U473 ( .A(A[14]), .B(n1848), .Z(n398) );
  CND2X4 U474 ( .A(n288), .B(n265), .Z(n255) );
  CND2X4 U475 ( .A(n288), .B(n265), .Z(n256) );
  CND2X2 U476 ( .A(n288), .B(n265), .Z(n2387) );
  CEOX4 U477 ( .A(A[18]), .B(n276), .Z(n288) );
  CND2X1 U478 ( .A(n2534), .B(n2533), .Z(n2536) );
  CEOX1 U479 ( .A(n1169), .B(n1171), .Z(n257) );
  CEOX1 U480 ( .A(n257), .B(n1170), .Z(\mult_x_1/n1511 ) );
  CND2X1 U481 ( .A(n1170), .B(n1171), .Z(n258) );
  CND2X1 U482 ( .A(n1170), .B(n1169), .Z(n259) );
  CIVX2 U483 ( .A(n245), .Z(n260) );
  CIVX3 U484 ( .A(n260), .Z(n261) );
  CND2X1 U485 ( .A(n853), .B(n852), .Z(n854) );
  CENX1 U486 ( .A(n853), .B(n720), .Z(n857) );
  CEOX4 U487 ( .A(A[4]), .B(n247), .Z(n352) );
  CENX4 U488 ( .A(n1829), .B(A[6]), .Z(n347) );
  CIVX2 U489 ( .A(n8), .Z(n262) );
  CIVX2 U490 ( .A(n262), .Z(n263) );
  COND2X1 U491 ( .A(n1209), .B(n270), .C(n642), .D(n1244), .Z(n648) );
  COND2X2 U492 ( .A(n2436), .B(n1768), .C(n2434), .D(n1213), .Z(n1781) );
  COND2X2 U493 ( .A(n2436), .B(n1643), .C(n2434), .D(n1642), .Z(n1664) );
  CIVX8 U494 ( .A(n1346), .Z(n2470) );
  CFA1X2 U495 ( .A(n664), .B(n663), .CI(n662), .CO(n1150), .S(n668) );
  CENX4 U496 ( .A(A[8]), .B(n270), .Z(n264) );
  CIVDX3 U497 ( .A(A[7]), .Z0(n270), .Z1(n271) );
  CENX4 U498 ( .A(n1600), .B(A[18]), .Z(n265) );
  COND1X1 U499 ( .A(n803), .B(n802), .C(n801), .Z(n2029) );
  CENX1 U500 ( .A(n948), .B(n1016), .Z(n2911) );
  CENX4 U501 ( .A(n354), .B(A[4]), .Z(n1861) );
  COR2X1 U502 ( .A(n827), .B(n826), .Z(n267) );
  CIVX8 U503 ( .A(n484), .Z(n1637) );
  CNIVX2 U504 ( .A(n1834), .Z(n269) );
  COND2X1 U505 ( .A(n13), .B(n597), .C(n1842), .D(n596), .Z(n598) );
  COR2X1 U506 ( .A(n525), .B(n524), .Z(n272) );
  COR2X1 U507 ( .A(n938), .B(n937), .Z(n273) );
  COR2X1 U508 ( .A(n731), .B(n730), .Z(n274) );
  COR2X1 U509 ( .A(n944), .B(n943), .Z(n275) );
  CIVDX4 U510 ( .A(n289), .Z0(n276), .Z1(n277) );
  CND2X1 U511 ( .A(n1106), .B(n1104), .Z(n280) );
  CIVX2 U512 ( .A(n2571), .Z(n1107) );
  CND2X1 U513 ( .A(n2549), .B(n28), .Z(n278) );
  COR2X1 U514 ( .A(n2640), .B(n279), .Z(n1106) );
  CND2X1 U515 ( .A(n2640), .B(n279), .Z(n1104) );
  CND2XL U516 ( .A(n2639), .B(n2638), .Z(n1109) );
  CNR2X1 U517 ( .A(n2639), .B(n2638), .Z(n623) );
  CIVXL U518 ( .A(n623), .Z(n281) );
  CIVX4 U519 ( .A(A[17]), .Z(n1446) );
  CIVX4 U520 ( .A(n1446), .Z(n1977) );
  CIVX4 U521 ( .A(A[15]), .Z(n291) );
  CIVX8 U522 ( .A(n283), .Z(n1834) );
  CND2X4 U523 ( .A(n284), .B(n1834), .Z(n2233) );
  CIVX8 U524 ( .A(n1446), .Z(n1600) );
  CNIVX2 U525 ( .A(B[21]), .Z(n1811) );
  CENX1 U526 ( .A(n1600), .B(n1811), .Z(n285) );
  CNIVX1 U527 ( .A(n1834), .Z(n2231) );
  CNIVX2 U528 ( .A(B[22]), .Z(n1717) );
  CENX1 U529 ( .A(n1600), .B(n1717), .Z(n1601) );
  COND2X1 U530 ( .A(n7), .B(n285), .C(n2231), .D(n1601), .Z(n2169) );
  CNIVX2 U531 ( .A(B[20]), .Z(n1961) );
  CENX1 U532 ( .A(n1600), .B(n1961), .Z(n1224) );
  COND2X1 U533 ( .A(n2233), .B(n1224), .C(n1834), .D(n285), .Z(n302) );
  CEOX1 U534 ( .A(A[28]), .B(A[29]), .Z(n286) );
  CIVX8 U535 ( .A(A[27]), .Z(n1254) );
  CIVX12 U536 ( .A(n1254), .Z(n1289) );
  CENX4 U537 ( .A(n1289), .B(A[28]), .Z(n404) );
  CIVX2 U538 ( .A(A[29]), .Z(n1684) );
  CNIVX2 U539 ( .A(B[8]), .Z(n1630) );
  CENX1 U540 ( .A(n254), .B(n1630), .Z(n1213) );
  CNIVX2 U541 ( .A(B[9]), .Z(n1699) );
  CENX1 U542 ( .A(n254), .B(n1699), .Z(n589) );
  COND2X1 U543 ( .A(n245), .B(n1213), .C(n2406), .D(n589), .Z(n301) );
  CEOX4 U544 ( .A(A[6]), .B(n1832), .Z(n348) );
  CIVX3 U545 ( .A(A[5]), .Z(n921) );
  CND2X2 U546 ( .A(n348), .B(n347), .Z(n1209) );
  CNIVX2 U547 ( .A(B[30]), .Z(n2389) );
  CENX1 U548 ( .A(n11), .B(n2389), .Z(n1208) );
  CENX4 U549 ( .A(n1829), .B(A[6]), .Z(n1877) );
  CNIVX4 U550 ( .A(\B_extended[32] ), .Z(n1965) );
  CENXL U551 ( .A(n1832), .B(n1965), .Z(n592) );
  COND2X1 U552 ( .A(n1209), .B(n1208), .C(n1877), .D(n592), .Z(n300) );
  CIVX4 U553 ( .A(A[19]), .Z(n289) );
  CENX2 U554 ( .A(n1600), .B(A[18]), .Z(n287) );
  CIVX4 U555 ( .A(n289), .Z(n1721) );
  CNIVX2 U556 ( .A(B[19]), .Z(n1697) );
  CENX1 U557 ( .A(n1721), .B(n1697), .Z(n293) );
  CENX2 U558 ( .A(n1600), .B(A[18]), .Z(n1722) );
  CENX1 U559 ( .A(n1721), .B(n1961), .Z(n610) );
  COND2X1 U560 ( .A(n255), .B(n293), .C(n1722), .D(n610), .Z(n2167) );
  CIVX8 U561 ( .A(n291), .Z(n1848) );
  CIVX4 U562 ( .A(A[13]), .Z(n565) );
  CENX2 U563 ( .A(n565), .B(A[14]), .Z(n290) );
  CIVX8 U564 ( .A(n290), .Z(n2002) );
  CND2X4 U565 ( .A(n398), .B(n2002), .Z(n1815) );
  CIVX2 U566 ( .A(n291), .Z(n550) );
  CENX1 U567 ( .A(n1973), .B(n1717), .Z(n1223) );
  CNIVX2 U568 ( .A(B[23]), .Z(n2426) );
  CENX1 U569 ( .A(n1973), .B(n2426), .Z(n602) );
  COND2X1 U570 ( .A(n1815), .B(n1223), .C(n2002), .D(n602), .Z(n308) );
  CIVX8 U571 ( .A(n1161), .Z(n1388) );
  CND2X4 U572 ( .A(n320), .B(n292), .Z(n1661) );
  CIVX2 U573 ( .A(A[23]), .Z(n1716) );
  CNIVX2 U574 ( .A(B[14]), .Z(n1703) );
  CENX1 U575 ( .A(n2395), .B(n1703), .Z(n1215) );
  CNIVX2 U576 ( .A(B[15]), .Z(n1981) );
  CENX1 U577 ( .A(n1970), .B(n1981), .Z(n604) );
  COND2X1 U578 ( .A(n1661), .B(n1215), .C(n292), .D(n604), .Z(n307) );
  CNIVX2 U579 ( .A(B[18]), .Z(n1969) );
  CENX1 U580 ( .A(n1721), .B(n1969), .Z(n1225) );
  COND2X1 U581 ( .A(n256), .B(n1225), .C(n2388), .D(n293), .Z(n306) );
  CIVX2 U582 ( .A(A[20]), .Z(n294) );
  CENX4 U583 ( .A(n1388), .B(n294), .Z(n395) );
  CENX2 U584 ( .A(A[19]), .B(A[20]), .Z(n295) );
  CNIVX4 U585 ( .A(n295), .Z(n396) );
  CND2X4 U586 ( .A(n395), .B(n396), .Z(n2392) );
  CNIVX2 U587 ( .A(B[16]), .Z(n1979) );
  CENX1 U588 ( .A(n1388), .B(n1979), .Z(n1216) );
  CNIVX8 U589 ( .A(n295), .Z(n2398) );
  CNIVX2 U590 ( .A(B[17]), .Z(n1831) );
  CENX1 U591 ( .A(n1388), .B(n1831), .Z(n605) );
  COND2X1 U592 ( .A(n2392), .B(n1216), .C(n2398), .D(n605), .Z(n305) );
  CIVX3 U593 ( .A(n346), .Z(n1704) );
  CIVX4 U594 ( .A(A[9]), .Z(n360) );
  CIVX8 U595 ( .A(n360), .Z(n1838) );
  CIVDX2 U596 ( .A(A[11]), .Z0(n346), .Z1(n1677) );
  CNIVX2 U597 ( .A(B[26]), .Z(n1972) );
  CENX1 U598 ( .A(n1677), .B(n1972), .Z(n1218) );
  CIVX8 U599 ( .A(n360), .Z(n1843) );
  CENX4 U600 ( .A(n1843), .B(A[10]), .Z(n2051) );
  CNIVX2 U601 ( .A(B[27]), .Z(n2393) );
  CENX1 U602 ( .A(n1677), .B(n2393), .Z(n595) );
  COND2X1 U603 ( .A(n2050), .B(n1218), .C(n2051), .D(n595), .Z(n304) );
  CENX2 U604 ( .A(n271), .B(A[8]), .Z(n298) );
  CENX1 U605 ( .A(n1843), .B(n2469), .Z(n1212) );
  CNIVX2 U606 ( .A(B[29]), .Z(n2441) );
  CENX1 U607 ( .A(n1843), .B(n2441), .Z(n593) );
  COND2X1 U608 ( .A(n6), .B(n1212), .C(n1924), .D(n593), .Z(n303) );
  CFA1X1 U609 ( .A(n302), .B(n301), .CI(n300), .CO(n2168), .S(n1266) );
  CFA1X1 U610 ( .A(n305), .B(n304), .CI(n303), .CO(n1194), .S(n1267) );
  CFA1X1 U611 ( .A(n308), .B(n307), .CI(n306), .CO(n1193), .S(n1268) );
  CIVX12 U612 ( .A(n565), .Z(n1975) );
  CEOX2 U613 ( .A(A[12]), .B(n1975), .Z(n310) );
  CENX2 U614 ( .A(n346), .B(A[12]), .Z(n309) );
  CIVX4 U615 ( .A(n309), .Z(n1842) );
  CNIVX2 U616 ( .A(B[24]), .Z(n1976) );
  CENX1 U617 ( .A(n1975), .B(n1976), .Z(n1214) );
  CNIVX2 U618 ( .A(B[25]), .Z(n1498) );
  CENX1 U619 ( .A(n1975), .B(n1498), .Z(n597) );
  COND2X1 U620 ( .A(n14), .B(n1214), .C(n1842), .D(n597), .Z(n1780) );
  CIVX4 U621 ( .A(A[25]), .Z(n319) );
  CNIVX2 U622 ( .A(B[12]), .Z(n1840) );
  CENX1 U623 ( .A(n1632), .B(n1840), .Z(n1219) );
  CNIVX2 U624 ( .A(B[13]), .Z(n1963) );
  CENX1 U625 ( .A(n1632), .B(n1963), .Z(n600) );
  COND2X1 U626 ( .A(n9), .B(n1219), .C(n2522), .D(n600), .Z(n1779) );
  CIVX8 U627 ( .A(n1254), .Z(n1982) );
  CEOX4 U628 ( .A(A[26]), .B(n1982), .Z(n323) );
  CNIVX4 U629 ( .A(n314), .Z(n322) );
  CND2X4 U630 ( .A(n323), .B(n322), .Z(n2432) );
  CNIVX2 U631 ( .A(B[10]), .Z(n1847) );
  CNIVX8 U632 ( .A(n314), .Z(n2430) );
  CNIVX2 U633 ( .A(B[11]), .Z(n1687) );
  COND2X1 U634 ( .A(n2432), .B(n1221), .C(n2430), .D(n588), .Z(n1778) );
  CENX1 U635 ( .A(n316), .B(n315), .Z(n317) );
  CENXL U636 ( .A(n318), .B(n317), .Z(\mult_x_1/n1089 ) );
  CNIVX2 U637 ( .A(n319), .Z(n1346) );
  CENX1 U638 ( .A(n2470), .B(n2426), .Z(n424) );
  CENX1 U639 ( .A(n2470), .B(n1976), .Z(n321) );
  COND2X1 U640 ( .A(n8), .B(n424), .C(n2522), .D(n321), .Z(n430) );
  CND2X4 U641 ( .A(n320), .B(n292), .Z(n2440) );
  CENX1 U642 ( .A(n2395), .B(n1498), .Z(n415) );
  CENX1 U643 ( .A(n2395), .B(n1972), .Z(n325) );
  COND2X1 U644 ( .A(n2440), .B(n415), .C(n292), .D(n325), .Z(n429) );
  CENX1 U645 ( .A(n1982), .B(n1811), .Z(n420) );
  CENX1 U646 ( .A(n1982), .B(n1717), .Z(n324) );
  COND2X1 U647 ( .A(n2432), .B(n420), .C(n2430), .D(n324), .Z(n428) );
  CENX1 U648 ( .A(n2470), .B(n1498), .Z(n334) );
  COND2X1 U649 ( .A(n8), .B(n321), .C(n2522), .D(n334), .Z(n337) );
  CENX1 U650 ( .A(n2390), .B(n2469), .Z(n330) );
  CENX1 U651 ( .A(n2390), .B(n2441), .Z(n2391) );
  COND2X1 U652 ( .A(n2392), .B(n330), .C(n2398), .D(n2391), .Z(n336) );
  CENX1 U653 ( .A(n1721), .B(n2389), .Z(n333) );
  CENX1 U654 ( .A(n1721), .B(n1965), .Z(n2386) );
  COND2X1 U655 ( .A(n256), .B(n333), .C(n287), .D(n2386), .Z(n335) );
  CND2X4 U656 ( .A(n323), .B(n322), .Z(n2310) );
  CENX1 U657 ( .A(n1982), .B(n2426), .Z(n338) );
  COND2X1 U658 ( .A(n2310), .B(n324), .C(n2430), .D(n338), .Z(n2415) );
  CENX1 U659 ( .A(n2395), .B(n2393), .Z(n2404) );
  COND2X1 U660 ( .A(n1661), .B(n325), .C(n292), .D(n2404), .Z(n2414) );
  CENX1 U661 ( .A(n254), .B(n1961), .Z(n331) );
  CNIVX4 U662 ( .A(n404), .Z(n2406) );
  CENX1 U663 ( .A(n254), .B(n1811), .Z(n2407) );
  COND2X1 U664 ( .A(n245), .B(n331), .C(n2406), .D(n2407), .Z(n2413) );
  CEOX1 U665 ( .A(A[30]), .B(\A_extended[32] ), .Z(n327) );
  CENX1 U666 ( .A(A[29]), .B(A[30]), .Z(n328) );
  CNIVX1 U667 ( .A(n328), .Z(n326) );
  CND2X4 U668 ( .A(n327), .B(n326), .Z(n2509) );
  CENX1 U669 ( .A(n1637), .B(n1969), .Z(n329) );
  CENX1 U670 ( .A(n1637), .B(n1697), .Z(n2402) );
  CNIVX4 U671 ( .A(n328), .Z(n2510) );
  COND2X1 U672 ( .A(n239), .B(n329), .C(n2402), .D(n2510), .Z(n2418) );
  CENX1 U673 ( .A(n1637), .B(n1831), .Z(n332) );
  CENX1 U674 ( .A(n2390), .B(n2393), .Z(n419) );
  CENX1 U675 ( .A(n254), .B(n1697), .Z(n421) );
  COND2X1 U676 ( .A(n245), .B(n421), .C(n2406), .D(n331), .Z(n418) );
  CENX1 U677 ( .A(n1637), .B(n1979), .Z(n2306) );
  COND2X1 U678 ( .A(n2509), .B(n2306), .C(n332), .D(n2510), .Z(n427) );
  CENX1 U679 ( .A(n1600), .B(n1965), .Z(n417) );
  CENX1 U680 ( .A(n1721), .B(n2441), .Z(n416) );
  CENX2 U681 ( .A(n1600), .B(A[18]), .Z(n2388) );
  COND2X1 U682 ( .A(n255), .B(n416), .C(n1722), .D(n333), .Z(n422) );
  CENX1 U683 ( .A(n2470), .B(n1972), .Z(n2394) );
  COND2X1 U684 ( .A(n263), .B(n334), .C(n2522), .D(n2394), .Z(n1277) );
  CFA1X1 U685 ( .A(n337), .B(n336), .CI(n335), .CO(n1276), .S(n1273) );
  CENX1 U686 ( .A(n1982), .B(n1976), .Z(n696) );
  COND2X1 U687 ( .A(n2432), .B(n338), .C(n2430), .D(n696), .Z(n1275) );
  CENX1 U688 ( .A(n340), .B(n339), .Z(n341) );
  CENXL U689 ( .A(n342), .B(n341), .Z(\mult_x_1/n869 ) );
  CEOX2 U690 ( .A(A[2]), .B(n354), .Z(n465) );
  CENX2 U691 ( .A(n371), .B(A[2]), .Z(n343) );
  CND2X2 U692 ( .A(n1880), .B(n465), .Z(n1857) );
  CENX1 U693 ( .A(n1533), .B(n1630), .Z(n353) );
  CENX1 U694 ( .A(n1387), .B(n1699), .Z(n706) );
  CNIVX1 U695 ( .A(B[0]), .Z(n1711) );
  CENXL U696 ( .A(n1711), .B(n1704), .Z(n344) );
  CENX4 U697 ( .A(n1843), .B(A[10]), .Z(n1967) );
  CIVX2 U698 ( .A(n346), .Z(n1966) );
  CNIVX2 U699 ( .A(B[1]), .Z(n1712) );
  CENX1 U700 ( .A(n1966), .B(n1712), .Z(n708) );
  CNIVX4 U701 ( .A(B[0]), .Z(n1714) );
  CND2IXL U702 ( .B(n1714), .A(n1704), .Z(n345) );
  COND2XL U703 ( .A(n246), .B(n346), .C(n345), .D(n2051), .Z(n718) );
  CND2X4 U704 ( .A(n348), .B(n347), .Z(n1920) );
  CNIVX2 U705 ( .A(B[4]), .Z(n1464) );
  CENX1 U706 ( .A(n11), .B(n1464), .Z(n349) );
  CNIVX2 U707 ( .A(B[5]), .Z(n1707) );
  CENXL U708 ( .A(n271), .B(n1707), .Z(n707) );
  CNIVX2 U709 ( .A(B[3]), .Z(n1694) );
  CENXL U710 ( .A(n1832), .B(n1694), .Z(n364) );
  CENX2 U711 ( .A(n1829), .B(A[6]), .Z(n1244) );
  COND2X1 U712 ( .A(n1209), .B(n364), .C(n1244), .D(n349), .Z(n361) );
  CIVX3 U713 ( .A(n371), .Z(n1470) );
  CIVX4 U714 ( .A(A[0]), .Z(n1884) );
  CND2X4 U715 ( .A(n1470), .B(n1884), .Z(n1886) );
  CENXL U716 ( .A(n1470), .B(n1699), .Z(n658) );
  CENX1 U717 ( .A(n1470), .B(n1847), .Z(n350) );
  CENX1 U718 ( .A(n1470), .B(n1687), .Z(n709) );
  COND2X1 U719 ( .A(n1886), .B(n350), .C(n1884), .D(n709), .Z(n717) );
  CND2X4 U720 ( .A(n352), .B(n351), .Z(n1893) );
  CNIVX2 U721 ( .A(B[6]), .Z(n1720) );
  CENX1 U722 ( .A(n1829), .B(n1720), .Z(n355) );
  CNIVX2 U723 ( .A(B[7]), .Z(n1701) );
  CENX1 U724 ( .A(n1829), .B(n1701), .Z(n714) );
  COND2X1 U725 ( .A(n1893), .B(n355), .C(n241), .D(n714), .Z(n716) );
  CNIVX2 U726 ( .A(B[2]), .Z(n1466) );
  CENX1 U727 ( .A(n1843), .B(n1466), .Z(n356) );
  CENX1 U728 ( .A(n1843), .B(n1694), .Z(n710) );
  COND2X1 U729 ( .A(n6), .B(n356), .C(n1924), .D(n710), .Z(n715) );
  CND2X2 U730 ( .A(n465), .B(n1880), .Z(n1882) );
  CIVX3 U731 ( .A(n579), .Z(n1718) );
  CENX1 U732 ( .A(n1718), .B(n1701), .Z(n363) );
  COND2X1 U733 ( .A(n1882), .B(n363), .C(n18), .D(n353), .Z(n1146) );
  CENX1 U734 ( .A(n1829), .B(n1707), .Z(n362) );
  COND2XL U735 ( .A(n1893), .B(n362), .C(n1861), .D(n355), .Z(n1145) );
  CENX1 U736 ( .A(n1843), .B(n1712), .Z(n357) );
  COND2X1 U737 ( .A(n6), .B(n357), .C(n1924), .D(n356), .Z(n1144) );
  CENXL U738 ( .A(n1711), .B(n1838), .Z(n358) );
  COND2X1 U739 ( .A(n6), .B(n358), .C(n1924), .D(n357), .Z(n661) );
  CND2IX1 U740 ( .B(n1714), .A(n1838), .Z(n359) );
  COND2XL U741 ( .A(n1926), .B(n360), .C(n359), .D(n1924), .Z(n660) );
  CENX1 U742 ( .A(n1829), .B(n1464), .Z(n645) );
  COND2X1 U743 ( .A(n1893), .B(n645), .C(n1861), .D(n362), .Z(n667) );
  CENX1 U744 ( .A(n1387), .B(n1720), .Z(n639) );
  COND2X1 U745 ( .A(n1882), .B(n639), .C(n18), .D(n363), .Z(n666) );
  CENXL U746 ( .A(n11), .B(n1466), .Z(n643) );
  COND2X1 U747 ( .A(n1920), .B(n643), .C(n1877), .D(n364), .Z(n665) );
  CENX1 U748 ( .A(n368), .B(n367), .Z(n369) );
  CENXL U749 ( .A(n370), .B(n369), .Z(\mult_x_1/n1675 ) );
  CENX1 U750 ( .A(n1632), .B(n1694), .Z(n1357) );
  CENX1 U751 ( .A(n1632), .B(n1464), .Z(n469) );
  COND2X1 U752 ( .A(n2524), .B(n1357), .C(n311), .D(n469), .Z(n1378) );
  CENX1 U753 ( .A(n1692), .B(n2393), .Z(n1349) );
  CENX1 U754 ( .A(n1692), .B(n2469), .Z(n482) );
  COND2X1 U755 ( .A(n1886), .B(n1349), .C(n1884), .D(n482), .Z(n1377) );
  CENX1 U756 ( .A(n11), .B(n1811), .Z(n1246) );
  CENX4 U757 ( .A(n1829), .B(A[6]), .Z(n1918) );
  CENX1 U758 ( .A(n11), .B(n1717), .Z(n475) );
  COND2X1 U759 ( .A(n1920), .B(n1246), .C(n1918), .D(n475), .Z(n377) );
  CENX1 U760 ( .A(n2390), .B(n1701), .Z(n1351) );
  CENX1 U761 ( .A(n1388), .B(n1630), .Z(n381) );
  COND2X1 U762 ( .A(n2392), .B(n1351), .C(n2398), .D(n381), .Z(n376) );
  CENX1 U763 ( .A(n1970), .B(n1707), .Z(n1355) );
  CENX1 U764 ( .A(n1970), .B(n1720), .Z(n470) );
  COND2X1 U765 ( .A(n1661), .B(n1355), .C(n292), .D(n470), .Z(n375) );
  CENX1 U766 ( .A(n1718), .B(n1498), .Z(n1365) );
  CENX1 U767 ( .A(n1718), .B(n1972), .Z(n480) );
  COND2X1 U768 ( .A(n1857), .B(n1365), .C(n1880), .D(n480), .Z(n374) );
  CENX1 U769 ( .A(n1829), .B(n2426), .Z(n1367) );
  CENX1 U770 ( .A(n1829), .B(n1976), .Z(n474) );
  COND2X1 U771 ( .A(n1893), .B(n1367), .C(n1861), .D(n474), .Z(n373) );
  COND2X1 U772 ( .A(n2310), .B(n1251), .C(n2430), .D(n472), .Z(n372) );
  CIVX2 U773 ( .A(n386), .Z(n378) );
  CFA1X1 U774 ( .A(n374), .B(n372), .CI(n373), .CO(n1670), .S(n1140) );
  CFA1X1 U775 ( .A(n376), .B(n377), .CI(n375), .CO(n1671), .S(n1139) );
  CENX1 U776 ( .A(n1975), .B(n1981), .Z(n1353) );
  CENX1 U777 ( .A(n1975), .B(n1979), .Z(n478) );
  COND2X1 U778 ( .A(n2055), .B(n1353), .C(n1842), .D(n478), .Z(n384) );
  CENX1 U779 ( .A(n1704), .B(n1831), .Z(n1347) );
  CENX1 U780 ( .A(n1966), .B(n1969), .Z(n1957) );
  COND2X1 U781 ( .A(n246), .B(n1347), .C(n1967), .D(n1957), .Z(n383) );
  CENX1 U782 ( .A(n1848), .B(n1963), .Z(n1371) );
  CENX1 U783 ( .A(n1973), .B(n1703), .Z(n1955) );
  COND2X1 U784 ( .A(n1815), .B(n1371), .C(n2002), .D(n1955), .Z(n382) );
  CENX2 U785 ( .A(n378), .B(n388), .Z(n385) );
  CENX1 U786 ( .A(n1843), .B(n1697), .Z(n1369) );
  CENX1 U787 ( .A(n1843), .B(n1961), .Z(n379) );
  COND2X1 U788 ( .A(n6), .B(n1369), .C(n1924), .D(n379), .Z(n2095) );
  CENX1 U789 ( .A(n1600), .B(n1687), .Z(n1361) );
  CENXL U790 ( .A(n1977), .B(n1840), .Z(n380) );
  COND2XL U791 ( .A(n7), .B(n1361), .C(n1834), .D(n380), .Z(n2094) );
  CENX1 U792 ( .A(n1721), .B(n1699), .Z(n1363) );
  CENX1 U793 ( .A(n1721), .B(n1847), .Z(n476) );
  COND2X1 U794 ( .A(n255), .B(n1363), .C(n1722), .D(n476), .Z(n2093) );
  CENX1 U795 ( .A(n1843), .B(n1811), .Z(n466) );
  COND2X1 U796 ( .A(n1926), .B(n379), .C(n1924), .D(n466), .Z(n1681) );
  CENXL U797 ( .A(n1977), .B(n1963), .Z(n1625) );
  COND2X1 U798 ( .A(n2233), .B(n380), .C(n1834), .D(n1625), .Z(n1680) );
  CND2X1 U799 ( .A(n396), .B(n395), .Z(n1163) );
  CENX1 U800 ( .A(n1388), .B(n1699), .Z(n1623) );
  COND2X1 U801 ( .A(n1163), .B(n381), .C(n2398), .D(n1623), .Z(n1679) );
  CFA1X1 U802 ( .A(n382), .B(n383), .CI(n384), .CO(n1674), .S(n1138) );
  CEO3X2 U803 ( .A(n1673), .B(n1675), .C(n1674), .Z(n387) );
  CEOX2 U804 ( .A(n387), .B(n385), .Z(\mult_x_1/n1339 ) );
  CND2XL U805 ( .A(n388), .B(n386), .Z(n391) );
  CND2X1 U806 ( .A(n386), .B(n387), .Z(n390) );
  CND2X1 U807 ( .A(n15), .B(n387), .Z(n389) );
  CND3X1 U808 ( .A(n391), .B(n390), .C(n389), .Z(\mult_x_1/n1338 ) );
  CENX1 U809 ( .A(n1632), .B(n1831), .Z(n1980) );
  CENX1 U810 ( .A(n1632), .B(n1969), .Z(n393) );
  COND2X1 U811 ( .A(n9), .B(n1980), .C(n2522), .D(n393), .Z(n2358) );
  CENX1 U812 ( .A(n2395), .B(n1697), .Z(n1971) );
  CENX1 U813 ( .A(n2395), .B(n1961), .Z(n392) );
  COND2X1 U814 ( .A(n2440), .B(n1971), .C(n292), .D(n392), .Z(n2357) );
  CENX1 U815 ( .A(n1973), .B(n2393), .Z(n1974) );
  CENX1 U816 ( .A(n1973), .B(n2469), .Z(n399) );
  COND2X1 U817 ( .A(n1815), .B(n1974), .C(n2002), .D(n399), .Z(n2356) );
  CENX1 U818 ( .A(n1721), .B(n1976), .Z(n394) );
  CENX1 U819 ( .A(n1721), .B(n1498), .Z(n400) );
  COND2X1 U820 ( .A(n256), .B(n394), .C(n287), .D(n400), .Z(n408) );
  CENX1 U821 ( .A(n2395), .B(n1811), .Z(n1420) );
  COND2X1 U822 ( .A(n2440), .B(n392), .C(n292), .D(n1420), .Z(n407) );
  CENX1 U823 ( .A(n2470), .B(n1697), .Z(n1418) );
  COND2X1 U824 ( .A(n9), .B(n393), .C(n2522), .D(n1418), .Z(n406) );
  CENXL U825 ( .A(n1977), .B(n1498), .Z(n1978) );
  CENXL U826 ( .A(n1977), .B(n1972), .Z(n402) );
  COND2XL U827 ( .A(n2233), .B(n1978), .C(n1834), .D(n402), .Z(n2355) );
  CENX1 U828 ( .A(n1721), .B(n2426), .Z(n1608) );
  COND2X1 U829 ( .A(n256), .B(n1608), .C(n2388), .D(n394), .Z(n2354) );
  CND2X4 U830 ( .A(n396), .B(n395), .Z(n2400) );
  CENX1 U831 ( .A(n2390), .B(n1811), .Z(n1962) );
  CENX1 U832 ( .A(n2390), .B(n1717), .Z(n397) );
  COND2X1 U833 ( .A(n2400), .B(n1962), .C(n2398), .D(n397), .Z(n2353) );
  CENXL U834 ( .A(n1977), .B(n2393), .Z(n401) );
  CENX1 U835 ( .A(n1600), .B(n2469), .Z(n2232) );
  COND2X1 U836 ( .A(n2233), .B(n401), .C(n2231), .D(n2232), .Z(n1412) );
  CENX1 U837 ( .A(n2390), .B(n2426), .Z(n1419) );
  COND2X1 U838 ( .A(n2400), .B(n397), .C(n2398), .D(n1419), .Z(n1992) );
  CND2X4 U839 ( .A(n17), .B(n2002), .Z(n2004) );
  CENX1 U840 ( .A(n1973), .B(n2441), .Z(n1415) );
  COND2X1 U841 ( .A(n2004), .B(n399), .C(n2002), .D(n1415), .Z(n1991) );
  CENX1 U842 ( .A(n1975), .B(n2389), .Z(n2052) );
  CENX1 U843 ( .A(n1975), .B(n1965), .Z(n1414) );
  COND2X1 U844 ( .A(n14), .B(n2052), .C(n1842), .D(n1414), .Z(n1990) );
  CENX1 U845 ( .A(n1721), .B(n1972), .Z(n2235) );
  COND2X1 U846 ( .A(n255), .B(n400), .C(n287), .D(n2235), .Z(n1410) );
  CENX1 U847 ( .A(n1982), .B(n1979), .Z(n2015) );
  CENX1 U848 ( .A(n1982), .B(n1831), .Z(n403) );
  COND2X1 U849 ( .A(n2432), .B(n2015), .C(n2430), .D(n403), .Z(n1986) );
  CENX1 U850 ( .A(n254), .B(n1703), .Z(n2017) );
  CENX1 U851 ( .A(n254), .B(n1981), .Z(n405) );
  COND2X1 U852 ( .A(n245), .B(n2017), .C(n2434), .D(n405), .Z(n1985) );
  COND2X1 U853 ( .A(n7), .B(n402), .C(n1834), .D(n401), .Z(n1984) );
  CENX1 U854 ( .A(n1637), .B(n1963), .Z(n1413) );
  CENX1 U855 ( .A(n1637), .B(n1703), .Z(n425) );
  COND2X1 U856 ( .A(n2509), .B(n1413), .C(n425), .D(n2510), .Z(n1423) );
  COND2X1 U857 ( .A(n2432), .B(n403), .C(n2430), .D(n1505), .Z(n1422) );
  CENX1 U858 ( .A(n254), .B(n1979), .Z(n1500) );
  CFA1X1 U859 ( .A(n408), .B(n407), .CI(n406), .CO(n1425), .S(n1184) );
  CEO3X2 U860 ( .A(n1424), .B(n1426), .C(n1425), .Z(n410) );
  CND2XL U861 ( .A(n409), .B(n411), .Z(n414) );
  CND2XL U862 ( .A(n409), .B(n410), .Z(n413) );
  CND2XL U863 ( .A(n411), .B(n410), .Z(n412) );
  CND3XL U864 ( .A(n414), .B(n413), .C(n412), .Z(\mult_x_1/n960 ) );
  CENX1 U865 ( .A(n2395), .B(n1976), .Z(n1496) );
  COND2X1 U866 ( .A(n2440), .B(n1496), .C(n292), .D(n415), .Z(n1588) );
  CENX1 U867 ( .A(n1721), .B(n2469), .Z(n1495) );
  COND2X1 U868 ( .A(n256), .B(n1495), .C(n287), .D(n416), .Z(n1587) );
  CENX1 U869 ( .A(n1600), .B(n2389), .Z(n426) );
  COND2X1 U870 ( .A(n2233), .B(n426), .C(n1834), .D(n417), .Z(n1586) );
  CENX1 U871 ( .A(n2390), .B(n1972), .Z(n1499) );
  COND2X1 U872 ( .A(n2400), .B(n1499), .C(n2398), .D(n419), .Z(n2379) );
  CENX1 U873 ( .A(n1982), .B(n1961), .Z(n2308) );
  COND2X1 U874 ( .A(n2432), .B(n2308), .C(n2430), .D(n420), .Z(n2378) );
  CENX1 U875 ( .A(n254), .B(n1969), .Z(n2311) );
  COND2X1 U876 ( .A(n245), .B(n2311), .C(n2434), .D(n421), .Z(n2377) );
  CFA1X1 U877 ( .A(n427), .B(n423), .CI(n422), .CO(n431), .S(n1137) );
  CENX1 U878 ( .A(n2470), .B(n1717), .Z(n1497) );
  CENX1 U879 ( .A(n1637), .B(n1981), .Z(n2307) );
  COND2X1 U880 ( .A(n2509), .B(n425), .C(n2307), .D(n2510), .Z(n2305) );
  CENX1 U881 ( .A(n1848), .B(n1965), .Z(n1503) );
  CAOR1X1 U882 ( .A(n2002), .B(n2004), .C(n1503), .Z(n2304) );
  CENX1 U883 ( .A(n1600), .B(n2441), .Z(n2230) );
  COND2X1 U884 ( .A(n7), .B(n2230), .C(n1834), .D(n426), .Z(n2303) );
  CFA1X1 U885 ( .A(n430), .B(n429), .CI(n428), .CO(n1274), .S(n1135) );
  CND2X1 U886 ( .A(n434), .B(n433), .Z(\mult_x_1/n880 ) );
  CFA1X1 U887 ( .A(n2708), .B(n2707), .CI(n2711), .CO(n436), .S(n883) );
  CFA1X1 U888 ( .A(n2709), .B(n435), .CI(n2705), .CO(n437), .S(n882) );
  CNR2X1 U889 ( .A(n735), .B(n734), .Z(\mult_x_1/n471 ) );
  CIVX1 U890 ( .A(\mult_x_1/n471 ), .Z(n736) );
  CFA1X1 U891 ( .A(n2703), .B(n2702), .CI(n2706), .CO(n441), .S(n439) );
  CFA1X1 U892 ( .A(n2704), .B(n436), .CI(n2700), .CO(n442), .S(n438) );
  CFA1X1 U893 ( .A(n439), .B(n438), .CI(n437), .CO(n732), .S(n735) );
  CNR2X1 U894 ( .A(n733), .B(n732), .Z(n440) );
  CIVX2 U895 ( .A(n440), .Z(n970) );
  CND2X1 U896 ( .A(n736), .B(n970), .Z(\mult_x_1/n460 ) );
  CFA1X1 U897 ( .A(n2701), .B(n2697), .CI(n2698), .CO(n445), .S(n444) );
  CFA1X1 U898 ( .A(n2699), .B(n441), .CI(n2695), .CO(n446), .S(n443) );
  CFA1X1 U899 ( .A(n444), .B(n443), .CI(n442), .CO(n749), .S(n733) );
  COR2X1 U900 ( .A(n750), .B(n749), .Z(n1117) );
  CFA1X1 U901 ( .A(n2693), .B(n2692), .CI(n2696), .CO(n457), .S(n448) );
  CFA1X1 U902 ( .A(n2694), .B(n445), .CI(n2690), .CO(n458), .S(n447) );
  CFA1X1 U903 ( .A(n448), .B(n447), .CI(n446), .CO(n730), .S(n750) );
  CND2X1 U904 ( .A(n1117), .B(n274), .Z(n1048) );
  CNR2X1 U905 ( .A(\mult_x_1/n460 ), .B(n1048), .Z(n1119) );
  CFA1X1 U906 ( .A(n2680), .B(n2681), .CI(n2683), .CO(n449), .S(n462) );
  CFA1X1 U907 ( .A(n2688), .B(n2687), .CI(n2691), .CO(n456), .S(n460) );
  CNR2X1 U908 ( .A(n744), .B(n743), .Z(n570) );
  CFA1X1 U909 ( .A(n2679), .B(n2677), .CI(n2676), .CO(n454), .S(n450) );
  CFA1X1 U910 ( .A(n2674), .B(n450), .CI(n449), .CO(n754), .S(n744) );
  CNR2X1 U911 ( .A(n755), .B(n754), .Z(n1055) );
  CNR2X1 U912 ( .A(n570), .B(n1055), .Z(n1057) );
  CFA1X1 U913 ( .A(n2671), .B(n2669), .CI(n2668), .CO(n451), .S(n453) );
  CFA1X1 U914 ( .A(n2675), .B(n2673), .CI(n2672), .CO(n452), .S(n455) );
  COR2X1 U915 ( .A(n759), .B(n758), .Z(n1066) );
  CFA1X1 U916 ( .A(n2666), .B(n2665), .CI(n451), .CO(n766), .S(n759) );
  COR2X1 U917 ( .A(n766), .B(n765), .Z(n1071) );
  CND2X1 U918 ( .A(n1066), .B(n1071), .Z(n1073) );
  CFA1X1 U919 ( .A(n2667), .B(n453), .CI(n452), .CO(n758), .S(n748) );
  CFA1X1 U920 ( .A(n2670), .B(n455), .CI(n454), .CO(n747), .S(n755) );
  CNR2X1 U921 ( .A(n748), .B(n747), .Z(n1059) );
  CNR2X1 U922 ( .A(n1073), .B(n1059), .Z(n1076) );
  CND2X1 U923 ( .A(n1057), .B(n1076), .Z(n1079) );
  CFA1X1 U924 ( .A(n2685), .B(n456), .CI(n2684), .CO(n461), .S(n464) );
  CFA1X1 U925 ( .A(n2689), .B(n457), .CI(n2686), .CO(n463), .S(n459) );
  CFA1X1 U926 ( .A(n460), .B(n459), .CI(n458), .CO(n737), .S(n731) );
  COR2X1 U927 ( .A(n738), .B(n737), .Z(n1118) );
  CFA1X1 U928 ( .A(n2678), .B(n462), .CI(n461), .CO(n743), .S(n746) );
  CFA1X1 U929 ( .A(n2682), .B(n464), .CI(n463), .CO(n745), .S(n738) );
  COR2X1 U930 ( .A(n746), .B(n745), .Z(n1051) );
  CND2X1 U931 ( .A(n1118), .B(n1051), .Z(n1052) );
  CNR2X1 U932 ( .A(n1079), .B(n1052), .Z(n1082) );
  CND2XL U933 ( .A(n1119), .B(n1082), .Z(\mult_x_1/n353 ) );
  CIVDX2 U934 ( .A(\A_extended[32] ), .Z0(n484), .Z1(n2427) );
  CENX1 U935 ( .A(n2427), .B(n1961), .Z(n2401) );
  CENX1 U936 ( .A(n2427), .B(n1811), .Z(n698) );
  COND2X1 U937 ( .A(n239), .B(n2401), .C(n698), .D(n2510), .Z(n2527) );
  CNIVX4 U938 ( .A(n1388), .Z(n1695) );
  CENX1 U939 ( .A(n1695), .B(n1965), .Z(n2397) );
  CAOR1X1 U940 ( .A(n2398), .B(n2400), .C(n2397), .Z(n2526) );
  CENX1 U941 ( .A(n2395), .B(n2441), .Z(n2396) );
  CENX1 U942 ( .A(n2395), .B(n2389), .Z(n713) );
  COND2X1 U943 ( .A(n2440), .B(n2396), .C(n292), .D(n713), .Z(n2525) );
  CND2X1 U944 ( .A(n465), .B(n1880), .Z(n1312) );
  CENX1 U945 ( .A(n1718), .B(n2393), .Z(n479) );
  CENX1 U946 ( .A(n1718), .B(n2469), .Z(n485) );
  COND2X1 U947 ( .A(n1312), .B(n479), .C(n18), .D(n485), .Z(n1636) );
  CENX1 U948 ( .A(n1829), .B(n1498), .Z(n473) );
  CENX1 U949 ( .A(n1829), .B(n1972), .Z(n1280) );
  COND2X1 U950 ( .A(n1893), .B(n473), .C(n1861), .D(n1280), .Z(n1635) );
  CENX1 U951 ( .A(n254), .B(n1712), .Z(n1682) );
  CENX1 U952 ( .A(n254), .B(n1466), .Z(n1643) );
  COND2X1 U953 ( .A(n245), .B(n1682), .C(n2406), .D(n1643), .Z(n1634) );
  CENX1 U954 ( .A(n1843), .B(n1717), .Z(n1279) );
  COND2X1 U955 ( .A(n1926), .B(n466), .C(n1924), .D(n1279), .Z(n488) );
  CENX1 U956 ( .A(n1975), .B(n1831), .Z(n477) );
  CENX1 U957 ( .A(n1975), .B(n1969), .Z(n1278) );
  COND2X1 U958 ( .A(n13), .B(n477), .C(n1842), .D(n1278), .Z(n487) );
  CENX1 U959 ( .A(n1973), .B(n1981), .Z(n1954) );
  CENX1 U960 ( .A(n1848), .B(n1979), .Z(n1281) );
  COND2X1 U961 ( .A(n1815), .B(n1954), .C(n2002), .D(n1281), .Z(n486) );
  CNR2IX1 U962 ( .B(n1714), .A(n2510), .Z(n489) );
  CENXL U963 ( .A(n1289), .B(n1694), .Z(n471) );
  COR2XL U964 ( .A(n2310), .B(n471), .Z(n468) );
  CENXL U965 ( .A(n1289), .B(n1464), .Z(n1641) );
  COR2XL U966 ( .A(n2430), .B(n1641), .Z(n467) );
  CND2X1 U967 ( .A(n468), .B(n467), .Z(n491) );
  CENX1 U968 ( .A(n1692), .B(n2441), .Z(n481) );
  CENX1 U969 ( .A(n21), .B(n2389), .Z(n1282) );
  COND2X1 U970 ( .A(n1886), .B(n481), .C(n1884), .D(n1282), .Z(n490) );
  CEO3X2 U971 ( .A(n489), .B(n491), .C(n490), .Z(n540) );
  CENX1 U972 ( .A(n1632), .B(n1707), .Z(n1633) );
  COND2X1 U973 ( .A(n9), .B(n469), .C(n2522), .D(n1633), .Z(n549) );
  CENX1 U974 ( .A(n2395), .B(n1701), .Z(n1631) );
  COND2X1 U975 ( .A(n1661), .B(n470), .C(n292), .D(n1631), .Z(n548) );
  COND2X1 U976 ( .A(n2310), .B(n472), .C(n2430), .D(n471), .Z(n547) );
  COND2X1 U977 ( .A(n1893), .B(n474), .C(n1861), .D(n473), .Z(n546) );
  CENX1 U978 ( .A(n11), .B(n2426), .Z(n1629) );
  COND2X1 U979 ( .A(n1920), .B(n475), .C(n1877), .D(n1629), .Z(n545) );
  CENX1 U980 ( .A(n1721), .B(n1687), .Z(n1627) );
  COND2X1 U981 ( .A(n2387), .B(n476), .C(n1722), .D(n1627), .Z(n544) );
  COND2X1 U982 ( .A(n2055), .B(n478), .C(n1842), .D(n477), .Z(n543) );
  COND2X1 U983 ( .A(n1857), .B(n480), .C(n18), .D(n479), .Z(n542) );
  COND2X1 U984 ( .A(n1886), .B(n482), .C(n1884), .D(n481), .Z(n541) );
  CND2IX1 U985 ( .B(n1714), .A(n1637), .Z(n483) );
  COND2X1 U986 ( .A(n2509), .B(n484), .C(n483), .D(n2510), .Z(n1799) );
  CENX1 U987 ( .A(n1718), .B(n2441), .Z(n1283) );
  CFA1X1 U988 ( .A(n488), .B(n487), .CI(n486), .CO(n2204), .S(n537) );
  CND2XL U989 ( .A(n489), .B(n491), .Z(n494) );
  CND2XL U990 ( .A(n489), .B(n490), .Z(n493) );
  CND2XL U991 ( .A(n491), .B(n490), .Z(n492) );
  CND3X1 U992 ( .A(n494), .B(n493), .C(n492), .Z(n2203) );
  CENXL U993 ( .A(n498), .B(n497), .Z(\mult_x_1/n1283 ) );
  CFA1X1 U994 ( .A(n2803), .B(n2804), .CI(n2802), .CO(n794), .S(n502) );
  CNR2X1 U995 ( .A(n500), .B(n499), .Z(n797) );
  CND2X1 U996 ( .A(n500), .B(n499), .Z(n796) );
  CFA1X1 U997 ( .A(n2801), .B(n502), .CI(n501), .CO(n499), .S(n533) );
  CFA1X1 U998 ( .A(n2807), .B(n2808), .CI(n2806), .CO(n501), .S(n519) );
  CNR2X1 U999 ( .A(n533), .B(n532), .Z(n793) );
  CIVX1 U1000 ( .A(n793), .Z(n2547) );
  CNR2X1 U1001 ( .A(n507), .B(n506), .Z(n2492) );
  CFA1X1 U1002 ( .A(n2831), .B(n2830), .CI(n2832), .CO(n506), .S(n505) );
  CNR2X1 U1003 ( .A(n505), .B(n504), .Z(n2491) );
  CNR2XL U1004 ( .A(n2492), .B(n2491), .Z(n509) );
  CFA1X1 U1005 ( .A(n2837), .B(n2833), .CI(n2834), .CO(n504), .S(n503) );
  COR2X1 U1006 ( .A(n503), .B(n2835), .Z(n727) );
  COR2X1 U1007 ( .A(n2836), .B(n2838), .Z(n2505) );
  COND1XL U1008 ( .A(n2611), .B(n2634), .C(n2612), .Z(n2513) );
  CNR2X1 U1009 ( .A(n2839), .B(n2840), .Z(n2511) );
  CND2XL U1010 ( .A(n2839), .B(n2840), .Z(n2512) );
  CND2XL U1011 ( .A(n2836), .B(n2838), .Z(n2504) );
  CIVX1 U1012 ( .A(n2504), .Z(n729) );
  CND2X1 U1013 ( .A(n503), .B(n2835), .Z(n726) );
  CND2X1 U1014 ( .A(n505), .B(n504), .Z(n2489) );
  CND2X1 U1015 ( .A(n507), .B(n506), .Z(n2493) );
  COND1XL U1016 ( .A(n2489), .B(n2492), .C(n2493), .Z(n508) );
  CANR1XL U1017 ( .A(n509), .B(n697), .C(n508), .Z(n674) );
  CNR2X1 U1018 ( .A(n513), .B(n512), .Z(n671) );
  CFA1X1 U1019 ( .A(n2825), .B(n2824), .CI(n2826), .CO(n512), .S(n511) );
  CFA1X1 U1020 ( .A(n2828), .B(n2827), .CI(n2829), .CO(n510), .S(n507) );
  CNR2X1 U1021 ( .A(n511), .B(n510), .Z(n673) );
  CNR2X1 U1022 ( .A(n671), .B(n673), .Z(n678) );
  CFA1X1 U1023 ( .A(n2822), .B(n2821), .CI(n2823), .CO(n514), .S(n513) );
  COR2X1 U1024 ( .A(n515), .B(n514), .Z(n676) );
  CND2X1 U1025 ( .A(n511), .B(n510), .Z(n2494) );
  CND2X1 U1026 ( .A(n513), .B(n512), .Z(n672) );
  COND1XL U1027 ( .A(n2494), .B(n671), .C(n672), .Z(n677) );
  CND2X1 U1028 ( .A(n515), .B(n514), .Z(n675) );
  CFA1X1 U1029 ( .A(n2819), .B(n2817), .CI(n2820), .CO(n522), .S(n515) );
  CNR2X1 U1030 ( .A(n523), .B(n522), .Z(n2458) );
  CIVX1 U1031 ( .A(n2458), .Z(n681) );
  CFA1X1 U1032 ( .A(n2811), .B(n2812), .CI(n2810), .CO(n518), .S(n521) );
  CFA1X1 U1033 ( .A(n2815), .B(n2818), .CI(n2814), .CO(n520), .S(n517) );
  CENX1 U1034 ( .A(n2809), .B(n520), .Z(n516) );
  CENX1 U1035 ( .A(n521), .B(n516), .Z(n525) );
  CFA1X1 U1036 ( .A(n2813), .B(n517), .CI(n2816), .CO(n524), .S(n523) );
  CND2X1 U1037 ( .A(n681), .B(n272), .Z(n2464) );
  CFA1X1 U1038 ( .A(n2805), .B(n519), .CI(n518), .CO(n532), .S(n529) );
  CNR2X1 U1039 ( .A(n529), .B(n528), .Z(n2465) );
  CNR2XL U1040 ( .A(n2464), .B(n2465), .Z(n531) );
  CND2X1 U1041 ( .A(n523), .B(n522), .Z(n2457) );
  CIVX1 U1042 ( .A(n2457), .Z(n527) );
  CND2X1 U1043 ( .A(n525), .B(n524), .Z(n2459) );
  CIVX1 U1044 ( .A(n2459), .Z(n526) );
  CANR1X1 U1045 ( .A(n527), .B(n272), .C(n526), .Z(n2462) );
  CND2X1 U1046 ( .A(n529), .B(n528), .Z(n2466) );
  CIVXL U1047 ( .A(n802), .Z(n2548) );
  CND2X1 U1048 ( .A(n533), .B(n532), .Z(n2546) );
  CENX1 U1049 ( .A(n538), .B(n537), .Z(n539) );
  CFA1X1 U1050 ( .A(n543), .B(n542), .CI(n541), .CO(n534), .S(n1131) );
  CFA1X1 U1051 ( .A(n546), .B(n545), .CI(n544), .CO(n535), .S(n1130) );
  CFA1X1 U1052 ( .A(n549), .B(n548), .CI(n547), .CO(n536), .S(n1129) );
  CENX1 U1053 ( .A(n1848), .B(n1712), .Z(n1439) );
  CND2IX1 U1054 ( .B(n1714), .A(n550), .Z(n551) );
  CENX1 U1055 ( .A(n1843), .B(n1720), .Z(n556) );
  CENX1 U1056 ( .A(n1843), .B(n1701), .Z(n1442) );
  COND2X1 U1057 ( .A(n6), .B(n556), .C(n1924), .D(n1442), .Z(n560) );
  CENX1 U1058 ( .A(n1829), .B(n1847), .Z(n561) );
  CENX1 U1059 ( .A(n1829), .B(n1687), .Z(n1440) );
  COND2X1 U1060 ( .A(n1893), .B(n561), .C(n242), .D(n1440), .Z(n559) );
  CENX1 U1061 ( .A(n1692), .B(n1703), .Z(n553) );
  CENX1 U1062 ( .A(n1692), .B(n1981), .Z(n1436) );
  COND2X1 U1063 ( .A(n1886), .B(n553), .C(n1884), .D(n1436), .Z(n558) );
  CENXL U1064 ( .A(n11), .B(n1630), .Z(n566) );
  CENXL U1065 ( .A(n11), .B(n1699), .Z(n1441) );
  COND2X1 U1066 ( .A(n1209), .B(n566), .C(n1244), .D(n1441), .Z(n1900) );
  CENX1 U1067 ( .A(n1966), .B(n1464), .Z(n554) );
  CENX1 U1068 ( .A(n1966), .B(n1707), .Z(n1438) );
  COND2X1 U1069 ( .A(n2050), .B(n554), .C(n1967), .D(n1438), .Z(n1899) );
  CENX1 U1070 ( .A(n1975), .B(n1466), .Z(n557) );
  CENX1 U1071 ( .A(n1975), .B(n1694), .Z(n1435) );
  COND2X1 U1072 ( .A(n14), .B(n557), .C(n1842), .D(n1435), .Z(n1898) );
  CENX1 U1073 ( .A(n1533), .B(n1840), .Z(n555) );
  CENX1 U1074 ( .A(n1718), .B(n1963), .Z(n1437) );
  COND2X1 U1075 ( .A(n1882), .B(n555), .C(n18), .D(n1437), .Z(n1903) );
  CNR2IX1 U1076 ( .B(n1714), .A(n2002), .Z(n1889) );
  CENX1 U1077 ( .A(n1690), .B(n1963), .Z(n1883) );
  COND2X1 U1078 ( .A(n1886), .B(n1883), .C(n1884), .D(n553), .Z(n1888) );
  CENX1 U1079 ( .A(n1966), .B(n1694), .Z(n1896) );
  COND2X1 U1080 ( .A(n246), .B(n1896), .C(n2051), .D(n554), .Z(n1887) );
  CNR2XL U1081 ( .A(n771), .B(n772), .Z(n569) );
  CENX1 U1082 ( .A(n1387), .B(n1687), .Z(n1879) );
  COND2X1 U1083 ( .A(n1882), .B(n1879), .C(n18), .D(n555), .Z(n2131) );
  CENX1 U1084 ( .A(n1843), .B(n1707), .Z(n1894) );
  COND2X1 U1085 ( .A(n6), .B(n1894), .C(n1924), .D(n556), .Z(n2130) );
  CENX1 U1086 ( .A(n1975), .B(n1712), .Z(n562) );
  CNIVX2 U1087 ( .A(n1842), .Z(n2053) );
  COND2X1 U1088 ( .A(n13), .B(n562), .C(n2053), .D(n557), .Z(n2129) );
  CFA1X1 U1089 ( .A(n560), .B(n559), .CI(n558), .CO(n2085), .S(n1620) );
  CENX1 U1090 ( .A(n1829), .B(n1699), .Z(n1890) );
  COND2X1 U1091 ( .A(n1893), .B(n1890), .C(n241), .D(n561), .Z(n2137) );
  CENX1 U1092 ( .A(n1714), .B(n1975), .Z(n563) );
  COND2XL U1093 ( .A(n13), .B(n563), .C(n1842), .D(n562), .Z(n705) );
  CND2IXL U1094 ( .B(n1714), .A(n1975), .Z(n564) );
  COND2XL U1095 ( .A(n13), .B(n565), .C(n564), .D(n1842), .Z(n704) );
  CENX1 U1096 ( .A(n11), .B(n1701), .Z(n1876) );
  COND2X1 U1097 ( .A(n1920), .B(n1876), .C(n1877), .D(n566), .Z(n2135) );
  CIVXL U1098 ( .A(n770), .Z(n568) );
  CND2XL U1099 ( .A(n771), .B(n772), .Z(n567) );
  COND1XL U1100 ( .A(n569), .B(n568), .C(n567), .Z(\mult_x_1/n1614 ) );
  CIVX1 U1101 ( .A(n1119), .Z(\mult_x_1/n440 ) );
  CNR2X1 U1102 ( .A(\mult_x_1/n440 ), .B(n1052), .Z(n1111) );
  CIVX1 U1103 ( .A(n570), .Z(n1053) );
  CND2XL U1104 ( .A(n1111), .B(n1053), .Z(\mult_x_1/n405 ) );
  CND2XL U1105 ( .A(n1111), .B(n1057), .Z(\mult_x_1/n394 ) );
  CENX1 U1106 ( .A(n572), .B(n571), .Z(n573) );
  CENX1 U1107 ( .A(n574), .B(n573), .Z(\mult_x_1/n881 ) );
  CENX1 U1108 ( .A(n1470), .B(n1712), .Z(n575) );
  COND2XL U1109 ( .A(n1886), .B(n1711), .C(n1884), .D(n575), .Z(n998) );
  CND2X1 U1110 ( .A(n998), .B(n997), .Z(n999) );
  CIVX1 U1111 ( .A(n999), .Z(n2502) );
  CENX1 U1112 ( .A(n1470), .B(n1466), .Z(n578) );
  COND2X1 U1113 ( .A(n1886), .B(n575), .C(n1884), .D(n578), .Z(n577) );
  CNR2IX1 U1114 ( .B(n1714), .A(n18), .Z(n576) );
  COR2X1 U1115 ( .A(n577), .B(n576), .Z(n2501) );
  CND2X1 U1116 ( .A(n577), .B(n576), .Z(n2500) );
  CENX1 U1117 ( .A(n1470), .B(n1694), .Z(n936) );
  CENX1 U1118 ( .A(n1387), .B(n1712), .Z(n934) );
  CNR2X1 U1119 ( .A(n581), .B(n580), .Z(n931) );
  CIVX1 U1120 ( .A(n931), .Z(n582) );
  CND2X1 U1121 ( .A(n581), .B(n580), .Z(n930) );
  CND2X1 U1122 ( .A(n582), .B(n930), .Z(n583) );
  CEOXL U1123 ( .A(n932), .B(n583), .Z(n2915) );
  CENX2 U1124 ( .A(n585), .B(n584), .Z(n586) );
  CENX1 U1125 ( .A(n587), .B(n586), .Z(\mult_x_1/n1311 ) );
  CENX1 U1126 ( .A(n1637), .B(n1701), .Z(n591) );
  CENX1 U1127 ( .A(n1637), .B(n1630), .Z(n1603) );
  CENX1 U1128 ( .A(n1982), .B(n1840), .Z(n590) );
  CENX1 U1129 ( .A(n254), .B(n1847), .Z(n611) );
  COND2X1 U1130 ( .A(n2436), .B(n589), .C(n2406), .D(n611), .Z(n1186) );
  CENX1 U1131 ( .A(n1975), .B(n1972), .Z(n596) );
  CENX1 U1132 ( .A(n1975), .B(n2393), .Z(n2000) );
  COND2X1 U1133 ( .A(n13), .B(n596), .C(n1842), .D(n2000), .Z(n608) );
  CENX1 U1134 ( .A(n2395), .B(n1979), .Z(n603) );
  CENX1 U1135 ( .A(n2395), .B(n1831), .Z(n2012) );
  COND2X1 U1136 ( .A(n1661), .B(n603), .C(n292), .D(n2012), .Z(n607) );
  CENX1 U1137 ( .A(n1677), .B(n2469), .Z(n594) );
  CENX1 U1138 ( .A(n1677), .B(n2441), .Z(n1611) );
  COND2X1 U1139 ( .A(n246), .B(n594), .C(n1967), .D(n1611), .Z(n606) );
  CENX1 U1140 ( .A(n1973), .B(n1976), .Z(n601) );
  CENX1 U1141 ( .A(n1973), .B(n1498), .Z(n2003) );
  COND2X1 U1142 ( .A(n2004), .B(n601), .C(n2002), .D(n2003), .Z(n1597) );
  CENX1 U1143 ( .A(n2470), .B(n1703), .Z(n599) );
  CENX1 U1144 ( .A(n2470), .B(n1981), .Z(n2006) );
  COND2X1 U1145 ( .A(n8), .B(n599), .C(n2522), .D(n2006), .Z(n1596) );
  CENX1 U1146 ( .A(n1982), .B(n1963), .Z(n1598) );
  COND2X1 U1147 ( .A(n2432), .B(n590), .C(n2430), .D(n1598), .Z(n1595) );
  CENX1 U1148 ( .A(n1637), .B(n1720), .Z(n1210) );
  COND2X1 U1149 ( .A(n2509), .B(n1210), .C(n591), .D(n2510), .Z(n2037) );
  CAOR1X1 U1150 ( .A(n1918), .B(n1209), .C(n592), .Z(n2036) );
  CENX1 U1151 ( .A(n1843), .B(n2389), .Z(n612) );
  COND2X1 U1152 ( .A(n1926), .B(n593), .C(n1924), .D(n612), .Z(n2035) );
  COND2X1 U1153 ( .A(n2050), .B(n595), .C(n2051), .D(n594), .Z(n1188) );
  COND2X1 U1154 ( .A(n8), .B(n600), .C(n2522), .D(n599), .Z(n1187) );
  COND2X1 U1155 ( .A(n2004), .B(n602), .C(n2002), .D(n601), .Z(n1191) );
  COND2X1 U1156 ( .A(n1661), .B(n604), .C(n292), .D(n603), .Z(n1190) );
  CENX1 U1157 ( .A(n1695), .B(n1969), .Z(n1604) );
  COND2X1 U1158 ( .A(n2392), .B(n605), .C(n2398), .D(n1604), .Z(n1189) );
  CENX1 U1159 ( .A(n1721), .B(n1811), .Z(n609) );
  CENX1 U1160 ( .A(n1721), .B(n1717), .Z(n1609) );
  COND2X1 U1161 ( .A(n256), .B(n609), .C(n2388), .D(n1609), .Z(n1607) );
  CFA1X1 U1162 ( .A(n608), .B(n607), .CI(n606), .CO(n1606), .S(n1516) );
  COND2X1 U1163 ( .A(n255), .B(n610), .C(n287), .D(n609), .Z(n2166) );
  CENX1 U1164 ( .A(n254), .B(n1687), .Z(n1599) );
  COND2X1 U1165 ( .A(n245), .B(n611), .C(n2406), .D(n1599), .Z(n2165) );
  CENX1 U1166 ( .A(n1843), .B(n1965), .Z(n1610) );
  COND2X1 U1167 ( .A(n1926), .B(n612), .C(n1924), .D(n1610), .Z(n2164) );
  CNR2X1 U1168 ( .A(\mult_x_1/n440 ), .B(n1064), .Z(n613) );
  CND2XL U1169 ( .A(n613), .B(n1066), .Z(\mult_x_1/n372 ) );
  CIVXL U1170 ( .A(n613), .Z(\mult_x_1/n381 ) );
  CENX1 U1171 ( .A(n254), .B(n2389), .Z(n614) );
  CENX1 U1172 ( .A(n254), .B(n1965), .Z(n615) );
  COND2X1 U1173 ( .A(n261), .B(n614), .C(n243), .D(n615), .Z(n629) );
  CENX1 U1174 ( .A(n2427), .B(n1972), .Z(n684) );
  CENX1 U1175 ( .A(n1637), .B(n2393), .Z(n631) );
  COND2X1 U1176 ( .A(n239), .B(n684), .C(n631), .D(n2510), .Z(n635) );
  CAOR1X1 U1177 ( .A(n2430), .B(n2310), .C(n634), .Z(n633) );
  CENX1 U1178 ( .A(n254), .B(n2441), .Z(n636) );
  COND2X1 U1179 ( .A(n245), .B(n636), .C(n2434), .D(n614), .Z(n632) );
  CENX1 U1180 ( .A(n1637), .B(n2469), .Z(n630) );
  CENX1 U1181 ( .A(n1637), .B(n2441), .Z(n616) );
  COND2X1 U1182 ( .A(n239), .B(n630), .C(n616), .D(n2510), .Z(n2499) );
  CIVX1 U1183 ( .A(n2499), .Z(n627) );
  CAOR1X1 U1184 ( .A(n243), .B(n261), .C(n615), .Z(n2498) );
  CENX1 U1185 ( .A(n2427), .B(n2389), .Z(n1121) );
  COND2X1 U1186 ( .A(n239), .B(n616), .C(n1121), .D(n2510), .Z(n2497) );
  CND2XL U1187 ( .A(n626), .B(n625), .Z(\mult_x_1/n246 ) );
  CFA1X1 U1188 ( .A(n2662), .B(n2660), .CI(n2664), .CO(n760), .S(n765) );
  COR2X1 U1189 ( .A(n761), .B(n760), .Z(n2845) );
  CFA1X1 U1190 ( .A(n2658), .B(n2661), .CI(n2663), .CO(n621), .S(n617) );
  CFA1X1 U1191 ( .A(n2657), .B(n617), .CI(n2659), .CO(n756), .S(n761) );
  COR2X1 U1192 ( .A(n757), .B(n756), .Z(n1085) );
  CND2X1 U1193 ( .A(n2845), .B(n1085), .Z(n751) );
  CNR2X1 U1194 ( .A(n1093), .B(n1092), .Z(n767) );
  CFA1X1 U1195 ( .A(n2642), .B(n2641), .CI(n2643), .CO(n279), .S(n769) );
  CFA1X1 U1196 ( .A(n2645), .B(n2646), .CI(n2644), .CO(n768), .S(n1092) );
  CNR2X1 U1197 ( .A(n769), .B(n768), .Z(n1095) );
  CNR2X1 U1198 ( .A(n767), .B(n1095), .Z(n1097) );
  CFA1X1 U1199 ( .A(n2648), .B(n618), .CI(n2647), .CO(n1093), .S(n764) );
  CFA1X1 U1200 ( .A(n2653), .B(n2651), .CI(n2650), .CO(n618), .S(n620) );
  CFA1X1 U1201 ( .A(n2654), .B(n2656), .CI(n2655), .CO(n619), .S(n622) );
  COR2X1 U1202 ( .A(n764), .B(n763), .Z(n1088) );
  CND2X1 U1203 ( .A(n1097), .B(n1088), .Z(n1100) );
  CFA1X1 U1204 ( .A(n2649), .B(n620), .CI(n619), .CO(n763), .S(n753) );
  CFA1X1 U1205 ( .A(n2652), .B(n622), .CI(n621), .CO(n752), .S(n757) );
  CNR2X1 U1206 ( .A(n753), .B(n752), .Z(n1086) );
  COR2X1 U1207 ( .A(n1100), .B(n1086), .Z(n1103) );
  CNR2X1 U1208 ( .A(n751), .B(n1103), .Z(\mult_x_1/n283 ) );
  CND2X1 U1209 ( .A(\mult_x_1/n283 ), .B(n1106), .Z(n624) );
  CIVXL U1210 ( .A(n624), .Z(\mult_x_1/n272 ) );
  CND2XL U1211 ( .A(n2550), .B(n2549), .Z(n1108) );
  COR2XL U1212 ( .A(n623), .B(n1108), .Z(n1110) );
  CNR2XL U1213 ( .A(n624), .B(n1110), .Z(\mult_x_1/n233 ) );
  CNR2X1 U1214 ( .A(n751), .B(n1086), .Z(\mult_x_1/n320 ) );
  CND2XL U1215 ( .A(\mult_x_1/n320 ), .B(n1088), .Z(n1090) );
  CNR2XL U1216 ( .A(\mult_x_1/n353 ), .B(n1090), .Z(\mult_x_1/n307 ) );
  COR2XL U1217 ( .A(n626), .B(n625), .Z(n2844) );
  CFA1X1 U1218 ( .A(n629), .B(n628), .CI(n627), .CO(n626), .S(n638) );
  COND2X1 U1219 ( .A(n239), .B(n631), .C(n630), .D(n2510), .Z(n2226) );
  CFA1X1 U1220 ( .A(n635), .B(n633), .CI(n632), .CO(n628), .S(n2225) );
  CENX1 U1221 ( .A(n1982), .B(n2389), .Z(n685) );
  COND2X1 U1222 ( .A(n2432), .B(n685), .C(n2430), .D(n634), .Z(n2160) );
  CIVX1 U1223 ( .A(n635), .Z(n2159) );
  CENX1 U1224 ( .A(n254), .B(n2469), .Z(n741) );
  COND2X1 U1225 ( .A(n16), .B(n741), .C(n243), .D(n636), .Z(n2158) );
  CND2XL U1226 ( .A(n638), .B(n637), .Z(\mult_x_1/n255 ) );
  COR2XL U1227 ( .A(n638), .B(n637), .Z(n2843) );
  CENX1 U1228 ( .A(n1470), .B(n1720), .Z(n653) );
  CENX1 U1229 ( .A(n1692), .B(n1701), .Z(n647) );
  COND2X1 U1230 ( .A(n1886), .B(n653), .C(n1884), .D(n647), .Z(n652) );
  COND2X1 U1231 ( .A(n1312), .B(n654), .C(n1880), .D(n640), .Z(n651) );
  CENX1 U1232 ( .A(n1829), .B(n1466), .Z(n914) );
  CENX1 U1233 ( .A(n1829), .B(n1694), .Z(n646) );
  COND2X1 U1234 ( .A(n1893), .B(n914), .C(n1861), .D(n646), .Z(n650) );
  COND2X1 U1235 ( .A(n248), .B(n640), .C(n18), .D(n639), .Z(n657) );
  CENXL U1236 ( .A(n1711), .B(n11), .Z(n641) );
  CENXL U1237 ( .A(n11), .B(n1712), .Z(n644) );
  COND2X1 U1238 ( .A(n1920), .B(n641), .C(n1918), .D(n644), .Z(n649) );
  CND2IXL U1239 ( .B(n1714), .A(n11), .Z(n642) );
  COND2X1 U1240 ( .A(n1920), .B(n644), .C(n1918), .D(n643), .Z(n655) );
  CNR2IX1 U1241 ( .B(n1714), .A(n1924), .Z(n664) );
  COND2X1 U1242 ( .A(n1893), .B(n646), .C(n1861), .D(n645), .Z(n663) );
  CENX1 U1243 ( .A(n1470), .B(n1630), .Z(n659) );
  COND2X1 U1244 ( .A(n1886), .B(n647), .C(n1884), .D(n659), .Z(n662) );
  CHA1X1 U1245 ( .A(n649), .B(n648), .CO(n656), .S(n913) );
  CFA1X1 U1246 ( .A(n652), .B(n650), .CI(n651), .CO(n670), .S(n912) );
  CENX1 U1247 ( .A(n1470), .B(n1707), .Z(n926) );
  COND2X1 U1248 ( .A(n1886), .B(n926), .C(n1884), .D(n653), .Z(n917) );
  CENX1 U1249 ( .A(n1387), .B(n1694), .Z(n929) );
  COND2X1 U1250 ( .A(n1312), .B(n929), .C(n18), .D(n654), .Z(n916) );
  CNR2IX1 U1251 ( .B(n1714), .A(n1244), .Z(n915) );
  CND2XL U1252 ( .A(n1911), .B(n1910), .Z(\mult_x_1/n701 ) );
  CFA1X1 U1253 ( .A(n657), .B(n656), .CI(n655), .CO(n1271), .S(n669) );
  COND2X1 U1254 ( .A(n1886), .B(n659), .C(n1884), .D(n658), .Z(n1152) );
  CHA1XL U1255 ( .A(n661), .B(n660), .CO(n1149), .S(n1151) );
  CFA1X1 U1256 ( .A(n667), .B(n666), .CI(n665), .CO(n1147), .S(n1269) );
  CFA1X1 U1257 ( .A(n670), .B(n669), .CI(n668), .CO(n1433), .S(n1911) );
  CIVX1 U1258 ( .A(n673), .Z(n2495) );
  CIVXL U1259 ( .A(n674), .Z(n2496) );
  CND2X1 U1260 ( .A(n676), .B(n675), .Z(n680) );
  CANR1XL U1261 ( .A(n678), .B(n2496), .C(n677), .Z(n679) );
  CEOXL U1262 ( .A(n680), .B(n679), .Z(n2902) );
  CND2X1 U1263 ( .A(n681), .B(n2457), .Z(n683) );
  CIVXL U1264 ( .A(n682), .Z(n2463) );
  CEOXL U1265 ( .A(n683), .B(n2463), .Z(n2901) );
  CENX1 U1266 ( .A(n2427), .B(n1498), .Z(n739) );
  COND2X1 U1267 ( .A(n239), .B(n739), .C(n684), .D(n2510), .Z(n2157) );
  CENX1 U1268 ( .A(n1982), .B(n2469), .Z(n2429) );
  CENX1 U1269 ( .A(n1982), .B(n2441), .Z(n686) );
  COND2X1 U1270 ( .A(n2432), .B(n2429), .C(n2430), .D(n686), .Z(n689) );
  CENX1 U1271 ( .A(n2470), .B(n2389), .Z(n2442) );
  CENX1 U1272 ( .A(n1632), .B(n1965), .Z(n740) );
  CENX1 U1273 ( .A(n254), .B(n1972), .Z(n2433) );
  CENX1 U1274 ( .A(n254), .B(n2393), .Z(n742) );
  COND2X1 U1275 ( .A(n245), .B(n2433), .C(n2434), .D(n742), .Z(n687) );
  COND2X1 U1276 ( .A(n2432), .B(n686), .C(n2430), .D(n685), .Z(n2155) );
  CFA1X1 U1277 ( .A(n689), .B(n688), .CI(n687), .CO(n2156), .S(\mult_x_1/n823 ) );
  CFA1X1 U1278 ( .A(n2718), .B(n2717), .CI(n2719), .CO(n875), .S(n879) );
  CFA1X1 U1279 ( .A(n2723), .B(n2721), .CI(n2722), .CO(n877), .S(n690) );
  CFA1X1 U1280 ( .A(n692), .B(n691), .CI(n690), .CO(n880), .S(n870) );
  CFA1X1 U1281 ( .A(n2729), .B(n2732), .CI(n2728), .CO(n692), .S(n859) );
  CFA1X1 U1282 ( .A(n2726), .B(n2720), .CI(n2724), .CO(n876), .S(n869) );
  CND2XL U1283 ( .A(n870), .B(n869), .Z(n693) );
  CNR2X1 U1284 ( .A(n695), .B(n694), .Z(n897) );
  CND2X1 U1285 ( .A(n695), .B(n694), .Z(n896) );
  CENX1 U1286 ( .A(n1982), .B(n1498), .Z(n699) );
  COND2X1 U1287 ( .A(n2310), .B(n696), .C(n2430), .D(n699), .Z(n2474) );
  CIVX1 U1288 ( .A(n2527), .Z(n2473) );
  CENX1 U1289 ( .A(n254), .B(n1717), .Z(n2405) );
  CENX1 U1290 ( .A(n254), .B(n2426), .Z(n700) );
  COND2X1 U1291 ( .A(n261), .B(n2405), .C(n2434), .D(n700), .Z(n2472) );
  CIVXL U1292 ( .A(n697), .Z(n2490) );
  CENX1 U1293 ( .A(n2427), .B(n1717), .Z(n2438) );
  COND2X1 U1294 ( .A(n239), .B(n698), .C(n2438), .D(n2510), .Z(n703) );
  CENX1 U1295 ( .A(n1982), .B(n1972), .Z(n711) );
  COND2XL U1296 ( .A(n2310), .B(n699), .C(n2430), .D(n711), .Z(n702) );
  CENX1 U1297 ( .A(n254), .B(n1976), .Z(n712) );
  COND2X1 U1298 ( .A(n261), .B(n700), .C(n2434), .D(n712), .Z(n701) );
  CFA1XL U1299 ( .A(n703), .B(n702), .CI(n701), .CO(\mult_x_1/n850 ), .S(
        \mult_x_1/n851 ) );
  CHA1XL U1300 ( .A(n705), .B(n704), .CO(n2136), .S(n2134) );
  CENX1 U1301 ( .A(n1387), .B(n1847), .Z(n1881) );
  COND2X1 U1302 ( .A(n1882), .B(n706), .C(n18), .D(n1881), .Z(n2334) );
  CENXL U1303 ( .A(n271), .B(n1720), .Z(n1878) );
  COND2X1 U1304 ( .A(n1920), .B(n707), .C(n1877), .D(n1878), .Z(n2333) );
  CENX1 U1305 ( .A(n1966), .B(n1466), .Z(n1897) );
  COND2X1 U1306 ( .A(n2050), .B(n708), .C(n2051), .D(n1897), .Z(n2332) );
  CNR2IX1 U1307 ( .B(n1714), .A(n2053), .Z(n2330) );
  CENX1 U1308 ( .A(n22), .B(n1840), .Z(n1885) );
  COND2X1 U1309 ( .A(n1886), .B(n709), .C(n1884), .D(n1885), .Z(n2329) );
  CENX1 U1310 ( .A(n1843), .B(n1464), .Z(n1895) );
  COND2X1 U1311 ( .A(n6), .B(n710), .C(n1924), .D(n1895), .Z(n2328) );
  CENX1 U1312 ( .A(n1982), .B(n2393), .Z(n2431) );
  COND2X1 U1313 ( .A(n2310), .B(n711), .C(n2430), .D(n2431), .Z(n2448) );
  CENX1 U1314 ( .A(n254), .B(n1498), .Z(n2435) );
  COND2X1 U1315 ( .A(n261), .B(n712), .C(n243), .D(n2435), .Z(n2447) );
  CENX1 U1316 ( .A(n1970), .B(n1965), .Z(n2439) );
  COND2X1 U1317 ( .A(n2440), .B(n713), .C(n292), .D(n2439), .Z(n2446) );
  CENX1 U1318 ( .A(n247), .B(n1630), .Z(n1892) );
  COND2XL U1319 ( .A(n1893), .B(n714), .C(n241), .D(n1892), .Z(n2193) );
  CFA1X1 U1320 ( .A(n717), .B(n716), .CI(n715), .CO(n2192), .S(n1142) );
  CHA1XL U1321 ( .A(n719), .B(n718), .CO(n2191), .S(n2331) );
  CENX1 U1322 ( .A(n852), .B(n851), .Z(n720) );
  CFA1X1 U1323 ( .A(n2747), .B(n2746), .CI(n2750), .CO(n852), .S(n722) );
  CFA1X1 U1324 ( .A(n2745), .B(n721), .CI(n2748), .CO(n853), .S(n845) );
  CFA1X1 U1325 ( .A(n2743), .B(n723), .CI(n722), .CO(n856), .S(n844) );
  CFA1X1 U1326 ( .A(n2753), .B(n2752), .CI(n2758), .CO(n721), .S(n776) );
  CNR2X2 U1327 ( .A(n725), .B(n724), .Z(n888) );
  CND2X1 U1328 ( .A(n725), .B(n724), .Z(n887) );
  CIVX1 U1329 ( .A(n728), .Z(n2507) );
  CND2X1 U1330 ( .A(n731), .B(n730), .Z(n1045) );
  CND2XL U1331 ( .A(n274), .B(n1045), .Z(\mult_x_1/n169 ) );
  CND2X1 U1332 ( .A(n733), .B(n732), .Z(n967) );
  CND2XL U1333 ( .A(n970), .B(n967), .Z(\mult_x_1/n171 ) );
  CND2X1 U1334 ( .A(n735), .B(n734), .Z(\mult_x_1/n472 ) );
  CND2XL U1335 ( .A(n736), .B(\mult_x_1/n472 ), .Z(\mult_x_1/n172 ) );
  CND2X1 U1336 ( .A(n738), .B(n737), .Z(n1049) );
  CND2XL U1337 ( .A(n1118), .B(n1049), .Z(\mult_x_1/n168 ) );
  CENX1 U1338 ( .A(n2427), .B(n1976), .Z(n2428) );
  COND2X1 U1339 ( .A(n239), .B(n2428), .C(n739), .D(n2510), .Z(n2425) );
  CAOR1X1 U1340 ( .A(n2522), .B(n263), .C(n740), .Z(n2154) );
  COND2X1 U1341 ( .A(n261), .B(n742), .C(n2434), .D(n741), .Z(n2153) );
  CND2X1 U1342 ( .A(n744), .B(n743), .Z(n1056) );
  CND2XL U1343 ( .A(n1053), .B(n1056), .Z(\mult_x_1/n166 ) );
  CND2X1 U1344 ( .A(n746), .B(n745), .Z(n1050) );
  CND2XL U1345 ( .A(n1051), .B(n1050), .Z(\mult_x_1/n167 ) );
  CND2X1 U1346 ( .A(n748), .B(n747), .Z(n1074) );
  CND2X1 U1347 ( .A(n750), .B(n749), .Z(n1044) );
  CND2XL U1348 ( .A(n1117), .B(n1044), .Z(\mult_x_1/n170 ) );
  CIVXL U1349 ( .A(n751), .Z(\mult_x_1/n331 ) );
  CND2X1 U1350 ( .A(n753), .B(n752), .Z(n1101) );
  CND2X1 U1351 ( .A(n755), .B(n754), .Z(n1054) );
  CND2X1 U1352 ( .A(n757), .B(n756), .Z(n1083) );
  CND2XL U1353 ( .A(n1085), .B(n1083), .Z(\mult_x_1/n160 ) );
  CND2X1 U1354 ( .A(n759), .B(n758), .Z(n1065) );
  CND2XL U1355 ( .A(n1066), .B(n1065), .Z(\mult_x_1/n163 ) );
  CND2X1 U1356 ( .A(n761), .B(n760), .Z(n762) );
  CND2XL U1357 ( .A(n2845), .B(n762), .Z(\mult_x_1/n161 ) );
  CIVX1 U1358 ( .A(n762), .Z(\mult_x_1/n349 ) );
  CND2X1 U1359 ( .A(n764), .B(n763), .Z(n1087) );
  CND2XL U1360 ( .A(n1088), .B(n1087), .Z(\mult_x_1/n158 ) );
  CND2X1 U1361 ( .A(n766), .B(n765), .Z(n1068) );
  CND2XL U1362 ( .A(n1071), .B(n1068), .Z(\mult_x_1/n162 ) );
  CIVXL U1363 ( .A(n767), .Z(\mult_x_1/n739 ) );
  CND2X1 U1364 ( .A(n769), .B(n768), .Z(n1094) );
  CNR2IXL U1365 ( .B(n1714), .A(n1884), .Z(n2918) );
  CEO3X1 U1366 ( .A(n772), .B(n771), .C(n770), .Z(\mult_x_1/n1615 ) );
  CEO3X1 U1367 ( .A(n775), .B(n774), .C(n773), .Z(\mult_x_1/n1043 ) );
  CFA1X1 U1368 ( .A(n2751), .B(n2754), .CI(n2756), .CO(n723), .S(n848) );
  CFA1X1 U1369 ( .A(n2749), .B(n777), .CI(n776), .CO(n843), .S(n847) );
  CFA1X1 U1370 ( .A(n2759), .B(n2760), .CI(n2762), .CO(n777), .S(n781) );
  CFA1X1 U1371 ( .A(n2757), .B(n778), .CI(n2755), .CO(n846), .S(n780) );
  CNR2X1 U1372 ( .A(n838), .B(n837), .Z(n956) );
  CFA1X1 U1373 ( .A(n781), .B(n780), .CI(n779), .CO(n837), .S(n836) );
  CFA1X1 U1374 ( .A(n2764), .B(n2765), .CI(n2767), .CO(n778), .S(n785) );
  CFA1X1 U1375 ( .A(n2763), .B(n782), .CI(n2761), .CO(n779), .S(n784) );
  CNR2X1 U1376 ( .A(n836), .B(n835), .Z(n962) );
  CNR2X1 U1377 ( .A(n956), .B(n962), .Z(n840) );
  CFA1X1 U1378 ( .A(n785), .B(n784), .CI(n783), .CO(n835), .S(n834) );
  CFA1X1 U1379 ( .A(n2769), .B(n2768), .CI(n2772), .CO(n782), .S(n791) );
  CFA1X1 U1380 ( .A(n2770), .B(n786), .CI(n2766), .CO(n783), .S(n790) );
  COND1X1 U1381 ( .A(n2773), .B(n792), .C(n2771), .Z(n788) );
  CND2X1 U1382 ( .A(n792), .B(n2773), .Z(n787) );
  CND2X1 U1383 ( .A(n788), .B(n787), .Z(n789) );
  CNR2X1 U1384 ( .A(n834), .B(n833), .Z(n949) );
  CFA1X1 U1385 ( .A(n791), .B(n790), .CI(n789), .CO(n833), .S(n832) );
  CFA1X1 U1386 ( .A(n2777), .B(n2775), .CI(n2774), .CO(n786), .S(n805) );
  CNR2X1 U1387 ( .A(n832), .B(n831), .Z(n952) );
  CNR2X1 U1388 ( .A(n949), .B(n952), .Z(n959) );
  CND2X1 U1389 ( .A(n840), .B(n959), .Z(n842) );
  CNR2X1 U1390 ( .A(n793), .B(n797), .Z(n2518) );
  CFA1X1 U1391 ( .A(n2799), .B(n2800), .CI(n2798), .CO(n817), .S(n795) );
  CFA1X1 U1392 ( .A(n2797), .B(n795), .CI(n794), .CO(n798), .S(n500) );
  COR2X1 U1393 ( .A(n799), .B(n798), .Z(n2516) );
  CND2XL U1394 ( .A(n2518), .B(n2516), .Z(n803) );
  COND1XL U1395 ( .A(n2546), .B(n797), .C(n796), .Z(n2517) );
  CND2X1 U1396 ( .A(n799), .B(n798), .Z(n2515) );
  CIVXL U1397 ( .A(n2515), .Z(n800) );
  CANR1XL U1398 ( .A(n2516), .B(n2517), .C(n800), .Z(n801) );
  CFA1X1 U1399 ( .A(n2782), .B(n2778), .CI(n2779), .CO(n792), .S(n809) );
  CFA1X1 U1400 ( .A(n2780), .B(n2776), .CI(n806), .CO(n804), .S(n808) );
  CFA1X1 U1401 ( .A(n2787), .B(n2783), .CI(n2784), .CO(n806), .S(n813) );
  CFA1X1 U1402 ( .A(n2785), .B(n810), .CI(n2781), .CO(n807), .S(n812) );
  CND2X1 U1403 ( .A(n267), .B(n2545), .Z(n830) );
  CFA1X1 U1404 ( .A(n813), .B(n812), .CI(n811), .CO(n824), .S(n822) );
  CFA1X1 U1405 ( .A(n2794), .B(n2788), .CI(n2789), .CO(n810), .S(n816) );
  CFA1X1 U1406 ( .A(n2792), .B(n2790), .CI(n2786), .CO(n811), .S(n815) );
  CFA1X1 U1407 ( .A(n2795), .B(n2793), .CI(n2796), .CO(n814), .S(n818) );
  CNR2X2 U1408 ( .A(n822), .B(n821), .Z(n823) );
  CIVX2 U1409 ( .A(n823), .Z(n2034) );
  CFA1X1 U1410 ( .A(n816), .B(n815), .CI(n814), .CO(n821), .S(n820) );
  CFA1X1 U1411 ( .A(n2791), .B(n818), .CI(n817), .CO(n819), .S(n799) );
  CNR2X1 U1412 ( .A(n820), .B(n819), .Z(n2032) );
  CIVX1 U1413 ( .A(n2032), .Z(n2538) );
  CND2X1 U1414 ( .A(n2034), .B(n2538), .Z(n2543) );
  CND2X1 U1415 ( .A(n820), .B(n819), .Z(n2537) );
  CND2X1 U1416 ( .A(n822), .B(n821), .Z(n2033) );
  CND2X1 U1417 ( .A(n827), .B(n826), .Z(n828) );
  CIVX2 U1418 ( .A(n828), .Z(n2031) );
  CND2X1 U1419 ( .A(n832), .B(n831), .Z(n1913) );
  CND2X1 U1420 ( .A(n834), .B(n833), .Z(n950) );
  COND1XL U1421 ( .A(n1913), .B(n949), .C(n950), .Z(n960) );
  CND2X1 U1422 ( .A(n836), .B(n835), .Z(n961) );
  CND2X1 U1423 ( .A(n838), .B(n837), .Z(n957) );
  COND1XL U1424 ( .A(n961), .B(n956), .C(n957), .Z(n839) );
  COND1X1 U1425 ( .A(n842), .B(n266), .C(n841), .Z(n1010) );
  CIVX2 U1426 ( .A(n1010), .Z(n1040) );
  CFA1X1 U1427 ( .A(n845), .B(n844), .CI(n843), .CO(n724), .S(n850) );
  CFA1X1 U1428 ( .A(n848), .B(n847), .CI(n846), .CO(n849), .S(n838) );
  CNR2X1 U1429 ( .A(n850), .B(n849), .Z(n1030) );
  CND2X1 U1430 ( .A(n850), .B(n849), .Z(n1029) );
  CFA1X1 U1431 ( .A(n2733), .B(n2731), .CI(n2735), .CO(n860), .S(n866) );
  COND1X2 U1432 ( .A(n852), .B(n853), .C(n851), .Z(n855) );
  CND2X2 U1433 ( .A(n855), .B(n854), .Z(n867) );
  CFA1X1 U1434 ( .A(n2741), .B(n2740), .CI(n2744), .CO(n864), .S(n851) );
  CFA1X1 U1435 ( .A(n2738), .B(n2736), .CI(n2742), .CO(n863), .S(n858) );
  CFA1X1 U1436 ( .A(n2739), .B(n2737), .CI(n2734), .CO(n861), .S(n862) );
  CFA1X1 U1437 ( .A(n858), .B(n857), .CI(n856), .CO(n889), .S(n725) );
  CNR2X1 U1438 ( .A(n890), .B(n889), .Z(n1035) );
  CFA1X1 U1439 ( .A(n2727), .B(n2725), .CI(n2730), .CO(n691), .S(n874) );
  CFA1X1 U1440 ( .A(n861), .B(n860), .CI(n859), .CO(n868), .S(n873) );
  CFA1X1 U1441 ( .A(n864), .B(n863), .CI(n862), .CO(n872), .S(n865) );
  CNR2X1 U1442 ( .A(n892), .B(n891), .Z(n2481) );
  CNR2X1 U1443 ( .A(n888), .B(n1030), .Z(n1036) );
  CEOX1 U1444 ( .A(n869), .B(n868), .Z(n871) );
  CEOX1 U1445 ( .A(n871), .B(n870), .Z(n895) );
  CFA1X1 U1446 ( .A(n874), .B(n873), .CI(n872), .CO(n894), .S(n892) );
  CNR2X1 U1447 ( .A(n895), .B(n894), .Z(n1022) );
  CNR2X1 U1448 ( .A(n1022), .B(n897), .Z(n1017) );
  CFA1X1 U1449 ( .A(n2713), .B(n2712), .CI(n2716), .CO(n435), .S(n886) );
  CFA1X1 U1450 ( .A(n2714), .B(n875), .CI(n2710), .CO(n881), .S(n885) );
  CFA1X1 U1451 ( .A(n877), .B(n876), .CI(n2715), .CO(n884), .S(n878) );
  CNR2X1 U1452 ( .A(n899), .B(n898), .Z(n2467) );
  CFA1X1 U1453 ( .A(n883), .B(n882), .CI(n881), .CO(n734), .S(n901) );
  CFA1X1 U1454 ( .A(n886), .B(n885), .CI(n884), .CO(n900), .S(n899) );
  CNR2X1 U1455 ( .A(n901), .B(n900), .Z(n2487) );
  CNR2X1 U1456 ( .A(n2467), .B(n2487), .Z(n903) );
  CND2X1 U1457 ( .A(n1017), .B(n903), .Z(n905) );
  CNR2XL U1458 ( .A(n1034), .B(n905), .Z(n907) );
  COND1X1 U1459 ( .A(n1029), .B(n888), .C(n887), .Z(n1038) );
  CNR2X1 U1460 ( .A(n1035), .B(n2481), .Z(n1012) );
  CND2X1 U1461 ( .A(n890), .B(n889), .Z(n2483) );
  CNR2XL U1462 ( .A(n892), .B(n891), .Z(n893) );
  CND2X1 U1463 ( .A(n892), .B(n891), .Z(n2482) );
  CANR1XL U1464 ( .A(n1038), .B(n1012), .C(n1011), .Z(n1033) );
  CND2X1 U1465 ( .A(n895), .B(n894), .Z(n2485) );
  COND1X1 U1466 ( .A(n2485), .B(n897), .C(n896), .Z(n1018) );
  CND2X1 U1467 ( .A(n899), .B(n898), .Z(n2468) );
  CND2X1 U1468 ( .A(n901), .B(n900), .Z(n2488) );
  COND1XL U1469 ( .A(n2487), .B(n2468), .C(n2488), .Z(n902) );
  CANR1XL U1470 ( .A(n1018), .B(n903), .C(n902), .Z(n904) );
  COND1XL U1471 ( .A(n905), .B(n1033), .C(n904), .Z(n906) );
  CANR1XL U1472 ( .A(n907), .B(n1010), .C(n906), .Z(\mult_x_1/n149 ) );
  CIVXL U1473 ( .A(n962), .Z(n908) );
  CAN2XL U1474 ( .A(n908), .B(n961), .Z(n910) );
  CIVX2 U1475 ( .A(n12), .Z(n1912) );
  CANR1X1 U1476 ( .A(n959), .B(n1912), .C(n960), .Z(n909) );
  CENXL U1477 ( .A(n910), .B(n909), .Z(n2889) );
  CFA1X1 U1478 ( .A(n913), .B(n912), .CI(n911), .CO(n1910), .S(n923) );
  CENX1 U1479 ( .A(n1829), .B(n1712), .Z(n918) );
  CFA1X1 U1480 ( .A(n917), .B(n916), .CI(n915), .CO(n911), .S(n925) );
  CENX1 U1481 ( .A(n1714), .B(n247), .Z(n919) );
  COND2X1 U1482 ( .A(n1893), .B(n919), .C(n1861), .D(n918), .Z(n928) );
  CND2IX1 U1483 ( .B(n1714), .A(n247), .Z(n920) );
  COND2X1 U1484 ( .A(n1893), .B(n5), .C(n920), .D(n1861), .Z(n927) );
  CND2X1 U1485 ( .A(n923), .B(n922), .Z(n1013) );
  CND2X2 U1486 ( .A(n1015), .B(n1013), .Z(n948) );
  CENX1 U1487 ( .A(n1470), .B(n1464), .Z(n935) );
  CHA1X1 U1488 ( .A(n928), .B(n927), .CO(n924), .S(n939) );
  COND1X1 U1489 ( .A(n932), .B(n931), .C(n930), .Z(n2412) );
  CNR2IX1 U1490 ( .B(n1714), .A(n241), .Z(n942) );
  COND2X1 U1491 ( .A(n1312), .B(n934), .C(n18), .D(n933), .Z(n941) );
  COND2X1 U1492 ( .A(n1886), .B(n936), .C(n1884), .D(n935), .Z(n940) );
  CND2X1 U1493 ( .A(n938), .B(n937), .Z(n2411) );
  CFA1X1 U1494 ( .A(n942), .B(n941), .CI(n940), .CO(n943), .S(n938) );
  CND2X1 U1495 ( .A(n944), .B(n943), .Z(n1042) );
  CIVX1 U1496 ( .A(n1042), .Z(n945) );
  CND2X1 U1497 ( .A(n947), .B(n946), .Z(n2533) );
  COND1X1 U1498 ( .A(n2532), .B(n2535), .C(n2533), .Z(n1016) );
  CIVXL U1499 ( .A(n949), .Z(n951) );
  CAN2XL U1500 ( .A(n951), .B(n950), .Z(n955) );
  CIVX1 U1501 ( .A(n1913), .Z(n953) );
  CENXL U1502 ( .A(n955), .B(n954), .Z(n2890) );
  CIVXL U1503 ( .A(n956), .Z(n958) );
  CAN2XL U1504 ( .A(n958), .B(n957), .Z(n966) );
  CANR1X1 U1505 ( .A(n964), .B(n1912), .C(n963), .Z(n965) );
  CENXL U1506 ( .A(n966), .B(n965), .Z(n2888) );
  CIVXL U1507 ( .A(\mult_x_1/n472 ), .Z(n969) );
  CIVX1 U1508 ( .A(n967), .Z(n968) );
  CANR1X1 U1509 ( .A(n970), .B(n969), .C(n968), .Z(\mult_x_1/n461 ) );
  CIVX2 U1510 ( .A(n2583), .Z(n1003) );
  CND2XL U1511 ( .A(n1003), .B(n2554), .Z(n972) );
  CIVX1 U1512 ( .A(n2618), .Z(n1004) );
  CANR1XL U1513 ( .A(n2554), .B(n1004), .C(n2555), .Z(n971) );
  COND1XL U1514 ( .A(n972), .B(n2635), .C(n971), .Z(n974) );
  CND2X1 U1515 ( .A(n2553), .B(n2572), .Z(n973) );
  CENX1 U1516 ( .A(n974), .B(n973), .Z(PRODUCT[58]) );
  COND1X1 U1517 ( .A(n2601), .B(n2635), .C(n2602), .Z(n975) );
  CENX1 U1518 ( .A(n975), .B(n2599), .Z(PRODUCT[41]) );
  COND1X1 U1519 ( .A(n2598), .B(n2635), .C(n2624), .Z(n976) );
  CENX1 U1520 ( .A(n976), .B(n2597), .Z(PRODUCT[42]) );
  COND1X1 U1521 ( .A(n2561), .B(n2635), .C(n2562), .Z(n977) );
  CENX1 U1522 ( .A(n977), .B(n2586), .Z(PRODUCT[49]) );
  CND2XL U1523 ( .A(n2577), .B(n2556), .Z(n979) );
  COND1XL U1524 ( .A(n979), .B(n2635), .C(n978), .Z(n980) );
  CENX1 U1525 ( .A(n980), .B(n2575), .Z(PRODUCT[56]) );
  CND2X1 U1526 ( .A(n2554), .B(n2553), .Z(n983) );
  CNR2X1 U1527 ( .A(n2583), .B(n983), .Z(n991) );
  CIVXL U1528 ( .A(n2572), .Z(n981) );
  CANR1XL U1529 ( .A(n2553), .B(n2555), .C(n981), .Z(n982) );
  COND1XL U1530 ( .A(n983), .B(n2618), .C(n982), .Z(n992) );
  CND2X1 U1531 ( .A(n1003), .B(n2559), .Z(n985) );
  CANR1XL U1532 ( .A(n2559), .B(n1004), .C(n2560), .Z(n984) );
  COND1X1 U1533 ( .A(n985), .B(n2635), .C(n984), .Z(n986) );
  CENX1 U1534 ( .A(n986), .B(n2581), .Z(PRODUCT[52]) );
  CIVXL U1535 ( .A(n2577), .Z(n988) );
  CIVXL U1536 ( .A(n2616), .Z(n987) );
  COND1XL U1537 ( .A(n988), .B(n2635), .C(n987), .Z(n990) );
  CND2X1 U1538 ( .A(n2556), .B(n2576), .Z(n989) );
  CENX1 U1539 ( .A(n990), .B(n989), .Z(PRODUCT[55]) );
  CND2XL U1540 ( .A(n991), .B(n2551), .Z(n994) );
  CANR1XL U1541 ( .A(n2551), .B(n992), .C(n2552), .Z(n993) );
  COND1XL U1542 ( .A(n994), .B(n2635), .C(n993), .Z(n995) );
  CENX1 U1543 ( .A(n995), .B(n2568), .Z(PRODUCT[60]) );
  COND1X1 U1544 ( .A(n2565), .B(n2635), .C(n2566), .Z(n996) );
  CENX1 U1545 ( .A(n996), .B(n2594), .Z(PRODUCT[44]) );
  CENX1 U1546 ( .A(n2628), .B(n2606), .Z(PRODUCT[36]) );
  CENX1 U1547 ( .A(n2627), .B(n2605), .Z(PRODUCT[37]) );
  CENX1 U1548 ( .A(n2626), .B(n2604), .Z(PRODUCT[38]) );
  CENX1 U1549 ( .A(n2625), .B(n2603), .Z(PRODUCT[39]) );
  CENX1 U1550 ( .A(n2630), .B(n2608), .Z(PRODUCT[34]) );
  CENX1 U1551 ( .A(n2629), .B(n2607), .Z(PRODUCT[35]) );
  CENX1 U1552 ( .A(n2631), .B(n2613), .Z(PRODUCT[33]) );
  CND2XL U1553 ( .A(n1003), .B(n2574), .Z(n1001) );
  CANR1XL U1554 ( .A(n2574), .B(n1004), .C(n2615), .Z(n1000) );
  COND1XL U1555 ( .A(n1001), .B(n2635), .C(n1000), .Z(n1002) );
  CENX1 U1556 ( .A(n1002), .B(n2573), .Z(PRODUCT[57]) );
  CND2XL U1557 ( .A(n1003), .B(n2567), .Z(n1006) );
  CANR1XL U1558 ( .A(n2567), .B(n1004), .C(n2614), .Z(n1005) );
  COND1XL U1559 ( .A(n1006), .B(n2635), .C(n1005), .Z(n1009) );
  CIVX1 U1560 ( .A(n2842), .Z(n1007) );
  COR2X1 U1561 ( .A(n2637), .B(n1007), .Z(n1126) );
  CND2X1 U1562 ( .A(n2637), .B(n1007), .Z(n1124) );
  CND2X1 U1563 ( .A(n1126), .B(n1124), .Z(n1008) );
  CENX1 U1564 ( .A(n1009), .B(n1008), .Z(PRODUCT[61]) );
  CIVXL U1565 ( .A(n1010), .Z(n1028) );
  CIVX1 U1566 ( .A(n1034), .Z(n1023) );
  CAOR1X1 U1567 ( .A(n1038), .B(n1012), .C(n1011), .Z(n1025) );
  CIVXL U1568 ( .A(n1013), .Z(n1014) );
  CANR1XL U1569 ( .A(n1016), .B(n1015), .C(n1014), .Z(\mult_x_1/n702 ) );
  CIVXL U1570 ( .A(n1018), .Z(n1019) );
  COND1XL U1571 ( .A(n2467), .B(n1019), .C(n2468), .Z(n1020) );
  CIVX1 U1572 ( .A(n1022), .Z(n2486) );
  CND2XL U1573 ( .A(n1023), .B(n2486), .Z(n1027) );
  CIVXL U1574 ( .A(n2485), .Z(n1024) );
  CANR1XL U1575 ( .A(n2486), .B(n1025), .C(n1024), .Z(n1026) );
  COND1XL U1576 ( .A(n1028), .B(n1027), .C(n1026), .Z(\mult_x_1/n506 ) );
  COND1XL U1577 ( .A(n1030), .B(n1040), .C(n1029), .Z(\mult_x_1/n542 ) );
  CIVXL U1578 ( .A(n1036), .Z(n1032) );
  CIVXL U1579 ( .A(n1038), .Z(n1031) );
  COND1XL U1580 ( .A(n1032), .B(n1040), .C(n1031), .Z(\mult_x_1/n531 ) );
  COND1XL U1581 ( .A(n1034), .B(n1040), .C(n1033), .Z(\mult_x_1/n513 ) );
  CIVX2 U1582 ( .A(n1035), .Z(n2484) );
  CND2XL U1583 ( .A(n1036), .B(n2484), .Z(n1041) );
  CIVX2 U1584 ( .A(n2483), .Z(n1037) );
  CANR1XL U1585 ( .A(n2484), .B(n1038), .C(n1037), .Z(n1039) );
  COND1XL U1586 ( .A(n1041), .B(n1040), .C(n1039), .Z(\mult_x_1/n524 ) );
  CND2X1 U1587 ( .A(n275), .B(n1042), .Z(n1043) );
  CENX1 U1588 ( .A(n1043), .B(n268), .Z(n2913) );
  CIVX1 U1589 ( .A(n1044), .Z(n1115) );
  CIVXL U1590 ( .A(n1045), .Z(n1046) );
  CANR1XL U1591 ( .A(n1115), .B(n274), .C(n1046), .Z(n1047) );
  COND1XL U1592 ( .A(n1048), .B(\mult_x_1/n461 ), .C(n1047), .Z(n1114) );
  CIVXL U1593 ( .A(n1114), .Z(\mult_x_1/n441 ) );
  CIVX1 U1594 ( .A(n1049), .Z(n1113) );
  COND1XL U1595 ( .A(n1052), .B(\mult_x_1/n441 ), .C(n1080), .Z(n1067) );
  COND1XL U1596 ( .A(n1056), .B(n1055), .C(n1054), .Z(n1077) );
  CANR1XL U1597 ( .A(n1057), .B(n1067), .C(n1077), .Z(\mult_x_1/n395 ) );
  CIVXL U1598 ( .A(n1080), .Z(n1062) );
  CIVXL U1599 ( .A(n1077), .Z(n1058) );
  COND1XL U1600 ( .A(n1059), .B(n1058), .C(n1074), .Z(n1060) );
  CANR1XL U1601 ( .A(n1062), .B(n1061), .C(n1060), .Z(n1063) );
  COND1XL U1602 ( .A(n1064), .B(\mult_x_1/n441 ), .C(n1063), .Z(n1091) );
  CIVX1 U1603 ( .A(n1065), .Z(n1070) );
  CANR1XL U1604 ( .A(n1066), .B(n1091), .C(n1070), .Z(\mult_x_1/n373 ) );
  CIVXL U1605 ( .A(n1067), .Z(\mult_x_1/n413 ) );
  CIVXL U1606 ( .A(n1068), .Z(n1069) );
  CANR1XL U1607 ( .A(n1071), .B(n1070), .C(n1069), .Z(n1072) );
  COND1XL U1608 ( .A(n1074), .B(n1073), .C(n1072), .Z(n1075) );
  CANR1XL U1609 ( .A(n1077), .B(n1076), .C(n1075), .Z(n1078) );
  COND1XL U1610 ( .A(n1080), .B(n1079), .C(n1078), .Z(n1081) );
  CANR1XL U1611 ( .A(n1082), .B(n1114), .C(n1081), .Z(\mult_x_1/n354 ) );
  CIVX1 U1612 ( .A(n1083), .Z(n1084) );
  CANR1X1 U1613 ( .A(\mult_x_1/n349 ), .B(n1085), .C(n1084), .Z(n1120) );
  COND1XL U1614 ( .A(n1086), .B(n1120), .C(n1101), .Z(\mult_x_1/n323 ) );
  CIVXL U1615 ( .A(n1087), .Z(n1098) );
  CANR1XL U1616 ( .A(n1088), .B(\mult_x_1/n323 ), .C(n1098), .Z(n1089) );
  COND1XL U1617 ( .A(n1090), .B(\mult_x_1/n354 ), .C(n1089), .Z(
        \mult_x_1/n308 ) );
  CIVXL U1618 ( .A(n1091), .Z(\mult_x_1/n382 ) );
  CND2X1 U1619 ( .A(n1093), .B(n1092), .Z(\mult_x_1/n303 ) );
  COND1XL U1620 ( .A(n1095), .B(\mult_x_1/n303 ), .C(n1094), .Z(n1096) );
  CANR1XL U1621 ( .A(n1098), .B(n1097), .C(n1096), .Z(n1099) );
  COAN1XL U1622 ( .A(n1101), .B(n1100), .C(n1099), .Z(n1102) );
  COND1X1 U1623 ( .A(n1103), .B(n1120), .C(n1102), .Z(\mult_x_1/n286 ) );
  CIVXL U1624 ( .A(n1104), .Z(n1105) );
  CANR1XL U1625 ( .A(n1106), .B(\mult_x_1/n286 ), .C(n1105), .Z(n1112) );
  CIVXL U1626 ( .A(n1111), .Z(\mult_x_1/n412 ) );
  CIVXL U1627 ( .A(n1112), .Z(\mult_x_1/n273 ) );
  CANR1XL U1628 ( .A(n1118), .B(n1114), .C(n1113), .Z(\mult_x_1/n428 ) );
  CIVXL U1629 ( .A(\mult_x_1/n461 ), .Z(n1116) );
  CANR1XL U1630 ( .A(n1117), .B(n1116), .C(n1115), .Z(\mult_x_1/n452 ) );
  CND2XL U1631 ( .A(n1119), .B(n1118), .Z(\mult_x_1/n427 ) );
  CIVXL U1632 ( .A(n1120), .Z(\mult_x_1/n332 ) );
  CENX1 U1633 ( .A(n2427), .B(n1965), .Z(n2508) );
  COND2XL U1634 ( .A(n239), .B(n1121), .C(n2508), .D(n2510), .Z(
        \mult_x_1/n794 ) );
  COND1X1 U1635 ( .A(n2596), .B(n2635), .C(n2623), .Z(n1122) );
  CENX1 U1636 ( .A(n1122), .B(n2595), .Z(PRODUCT[43]) );
  COND1X1 U1637 ( .A(n2590), .B(n2635), .C(n2621), .Z(n1123) );
  CENX1 U1638 ( .A(n1123), .B(n2589), .Z(PRODUCT[47]) );
  CND2X1 U1639 ( .A(n2567), .B(n1126), .Z(n1128) );
  CNR2X1 U1640 ( .A(n2583), .B(n1128), .Z(n1204) );
  CIVXL U1641 ( .A(n1124), .Z(n1125) );
  CANR1XL U1642 ( .A(n1126), .B(n2614), .C(n1125), .Z(n1127) );
  COND1XL U1643 ( .A(n1128), .B(n2618), .C(n1127), .Z(n1206) );
  COR2X1 U1644 ( .A(n2633), .B(n2842), .Z(n1207) );
  CND2X1 U1645 ( .A(n2633), .B(n2842), .Z(n1205) );
  CEOX1 U1646 ( .A(n2600), .B(n2635), .Z(PRODUCT[40]) );
  CFA1X1 U1647 ( .A(n1131), .B(n1130), .CI(n1129), .CO(n584), .S(
        \mult_x_1/n1343 ) );
  CFA1X1 U1648 ( .A(n1134), .B(n1133), .CI(n1132), .CO(n572), .S(
        \mult_x_1/n899 ) );
  CFA1X1 U1649 ( .A(n1137), .B(n1136), .CI(n1135), .CO(n574), .S(
        \mult_x_1/n897 ) );
  CFA1X1 U1650 ( .A(n1140), .B(n1139), .CI(n1138), .CO(n388), .S(
        \mult_x_1/n1371 ) );
  CFA1X1 U1651 ( .A(n1143), .B(n1142), .CI(n1141), .CO(\mult_x_1/n1676 ), .S(
        n370) );
  CFA1X1 U1652 ( .A(n1146), .B(n1145), .CI(n1144), .CO(n1141), .S(n1155) );
  CFA1X1 U1653 ( .A(n1149), .B(n1148), .CI(n1147), .CO(n368), .S(n1154) );
  CFA1X1 U1654 ( .A(n1152), .B(n1151), .CI(n1150), .CO(n1153), .S(n1270) );
  CFA1X1 U1655 ( .A(n1155), .B(n1154), .CI(n1153), .CO(\mult_x_1/n1684 ), .S(
        \mult_x_1/n1685 ) );
  CENX1 U1656 ( .A(n1838), .B(n1840), .Z(n1308) );
  CENX1 U1657 ( .A(n1838), .B(n1963), .Z(n1156) );
  COND2X1 U1658 ( .A(n1926), .B(n1308), .C(n1924), .D(n1156), .Z(n1325) );
  CENX1 U1659 ( .A(n1600), .B(n1464), .Z(n1159) );
  CENX1 U1660 ( .A(n1600), .B(n1707), .Z(n1164) );
  COND2X1 U1661 ( .A(n2233), .B(n1159), .C(n1834), .D(n1164), .Z(n1324) );
  CENX1 U1662 ( .A(n1721), .B(n1466), .Z(n1304) );
  CENX1 U1663 ( .A(n1721), .B(n1694), .Z(n1157) );
  COND2X1 U1664 ( .A(n2387), .B(n1304), .C(n2388), .D(n1157), .Z(n1323) );
  CENX1 U1665 ( .A(n11), .B(n1981), .Z(n1319) );
  CENX1 U1666 ( .A(n11), .B(n1979), .Z(n1919) );
  COND2X1 U1667 ( .A(n1209), .B(n1319), .C(n1244), .D(n1919), .Z(n1180) );
  CENX1 U1668 ( .A(n1966), .B(n1687), .Z(n1313) );
  CENX1 U1669 ( .A(n1704), .B(n1840), .Z(n1706) );
  COND2X1 U1670 ( .A(n246), .B(n1313), .C(n1967), .D(n1706), .Z(n1179) );
  CENX1 U1671 ( .A(n1838), .B(n1703), .Z(n1925) );
  COND2X1 U1672 ( .A(n6), .B(n1156), .C(n1924), .D(n1925), .Z(n1178) );
  CNR2IX1 U1673 ( .B(n1714), .A(n292), .Z(n1174) );
  CENX1 U1674 ( .A(n1721), .B(n1464), .Z(n1708) );
  COND2X1 U1675 ( .A(n2387), .B(n1157), .C(n287), .D(n1708), .Z(n1173) );
  CENX1 U1676 ( .A(n1692), .B(n1811), .Z(n1315) );
  CENX1 U1677 ( .A(n1692), .B(n1717), .Z(n1691) );
  COND2X1 U1678 ( .A(n1886), .B(n1315), .C(n1884), .D(n1691), .Z(n1172) );
  CENX1 U1679 ( .A(n247), .B(n1831), .Z(n1321) );
  CENX1 U1680 ( .A(n247), .B(n1969), .Z(n1698) );
  COND2X1 U1681 ( .A(n1893), .B(n1321), .C(n242), .D(n1698), .Z(n1177) );
  CENX1 U1682 ( .A(n1975), .B(n1699), .Z(n1158) );
  CENX1 U1683 ( .A(n1975), .B(n1847), .Z(n1688) );
  COND2X1 U1684 ( .A(n13), .B(n1158), .C(n1842), .D(n1688), .Z(n1176) );
  CENX1 U1685 ( .A(n1973), .B(n1701), .Z(n1317) );
  CENX1 U1686 ( .A(n1848), .B(n1630), .Z(n1700) );
  COND2X1 U1687 ( .A(n2004), .B(n1317), .C(n2002), .D(n1700), .Z(n1175) );
  COND2XL U1688 ( .A(n13), .B(n1309), .C(n1842), .D(n1158), .Z(n1492) );
  CNR2IX1 U1689 ( .B(n1714), .A(n2398), .Z(n1477) );
  CENX1 U1690 ( .A(n1600), .B(n1694), .Z(n1467) );
  COND2X1 U1691 ( .A(n2233), .B(n1467), .C(n1834), .D(n1159), .Z(n1476) );
  CENX1 U1692 ( .A(n1692), .B(n1697), .Z(n1471) );
  CENX1 U1693 ( .A(n1692), .B(n1961), .Z(n1316) );
  COND2X1 U1694 ( .A(n1886), .B(n1471), .C(n1884), .D(n1316), .Z(n1475) );
  CND2IXL U1695 ( .B(n1714), .A(n1388), .Z(n1160) );
  COND2X1 U1696 ( .A(n1163), .B(n1161), .C(n1160), .D(n2398), .Z(n1333) );
  CENXL U1697 ( .A(n1711), .B(n1388), .Z(n1162) );
  CENX1 U1698 ( .A(n1388), .B(n1712), .Z(n1165) );
  COND2X1 U1699 ( .A(n1163), .B(n1162), .C(n2398), .D(n1165), .Z(n1332) );
  CENX1 U1700 ( .A(n1718), .B(n1697), .Z(n1310) );
  CENX1 U1701 ( .A(n1718), .B(n1961), .Z(n1689) );
  COND2X1 U1702 ( .A(n1857), .B(n1310), .C(n18), .D(n1689), .Z(n2340) );
  CENX1 U1703 ( .A(n1600), .B(n1720), .Z(n1702) );
  COND2X1 U1704 ( .A(n7), .B(n1164), .C(n1834), .D(n1702), .Z(n2339) );
  CENX1 U1705 ( .A(n1695), .B(n1466), .Z(n1710) );
  COND2X1 U1706 ( .A(n2392), .B(n1165), .C(n2398), .D(n1710), .Z(n2338) );
  CFA1X1 U1707 ( .A(n1168), .B(n1167), .CI(n1166), .CO(n1182), .S(
        \mult_x_1/n1513 ) );
  CFA1X1 U1708 ( .A(n1174), .B(n1173), .CI(n1172), .CO(n1932), .S(n1166) );
  CFA1X1 U1709 ( .A(n1177), .B(n1176), .CI(n1175), .CO(n1931), .S(n1171) );
  CFA1X1 U1710 ( .A(n1180), .B(n1179), .CI(n1178), .CO(n1930), .S(n1167) );
  CFA1X1 U1711 ( .A(n1185), .B(n1184), .CI(n1183), .CO(n409), .S(
        \mult_x_1/n983 ) );
  CFA1X1 U1712 ( .A(n598), .B(n1188), .CI(n1187), .CO(n1199), .S(n1196) );
  CFA1X1 U1713 ( .A(n1191), .B(n1190), .CI(n1189), .CO(n1198), .S(n1195) );
  CFA1X1 U1714 ( .A(n1194), .B(n1193), .CI(n1192), .CO(n1203), .S(n315) );
  CFA1X1 U1715 ( .A(n1197), .B(n1196), .CI(n1195), .CO(n1202), .S(
        \mult_x_1/n1093 ) );
  CFA1X1 U1716 ( .A(n1200), .B(n1199), .CI(n1198), .CO(n775), .S(n1201) );
  CFA1X1 U1717 ( .A(n1203), .B(n1202), .CI(n1201), .CO(\mult_x_1/n1064 ), .S(
        \mult_x_1/n1065 ) );
  COND2X1 U1718 ( .A(n2432), .B(n1572), .C(n2430), .D(n1222), .Z(n1562) );
  CENX1 U1719 ( .A(n1388), .B(n1703), .Z(n1389) );
  CENX1 U1720 ( .A(n1388), .B(n1981), .Z(n1217) );
  COND2X1 U1721 ( .A(n2392), .B(n1389), .C(n2398), .D(n1217), .Z(n1561) );
  CENX1 U1722 ( .A(n1632), .B(n1847), .Z(n1571) );
  CENX1 U1723 ( .A(n1632), .B(n1687), .Z(n1220) );
  COND2X1 U1724 ( .A(n2524), .B(n1571), .C(n2522), .D(n1220), .Z(n1560) );
  CENX1 U1725 ( .A(n1637), .B(n1464), .Z(n1563) );
  CENX1 U1726 ( .A(n2427), .B(n1707), .Z(n1211) );
  COND2X1 U1727 ( .A(n2509), .B(n1563), .C(n1211), .D(n2510), .Z(n1786) );
  CENX1 U1728 ( .A(n1829), .B(n1965), .Z(n1776) );
  CAOR1X1 U1729 ( .A(n1861), .B(n1893), .C(n1776), .Z(n1785) );
  CENX1 U1730 ( .A(n11), .B(n2441), .Z(n1774) );
  COND2X1 U1731 ( .A(n1209), .B(n1774), .C(n1918), .D(n1208), .Z(n1784) );
  COND2X1 U1732 ( .A(n2509), .B(n1211), .C(n1210), .D(n2510), .Z(n1783) );
  CENX1 U1733 ( .A(n1843), .B(n2393), .Z(n1770) );
  COND2X1 U1734 ( .A(n1926), .B(n1770), .C(n1924), .D(n1212), .Z(n1782) );
  CENX1 U1735 ( .A(n254), .B(n1701), .Z(n1768) );
  CENX1 U1736 ( .A(n1975), .B(n2426), .Z(n1403) );
  COND2X1 U1737 ( .A(n2055), .B(n1403), .C(n1842), .D(n1214), .Z(n1234) );
  CENX1 U1738 ( .A(n2395), .B(n1963), .Z(n1766) );
  COND2X1 U1739 ( .A(n1661), .B(n1766), .C(n292), .D(n1215), .Z(n1233) );
  COND2X1 U1740 ( .A(n2400), .B(n1217), .C(n2398), .D(n1216), .Z(n1232) );
  CENX1 U1741 ( .A(n1677), .B(n1498), .Z(n1556) );
  COND2X1 U1742 ( .A(n2050), .B(n1556), .C(n1967), .D(n1218), .Z(n1237) );
  COND2X1 U1743 ( .A(n9), .B(n1220), .C(n2522), .D(n1219), .Z(n1236) );
  COND2X1 U1744 ( .A(n2310), .B(n1222), .C(n2430), .D(n1221), .Z(n1235) );
  CENX1 U1745 ( .A(n1973), .B(n1811), .Z(n1558) );
  CENX1 U1746 ( .A(n1600), .B(n1697), .Z(n1772) );
  COND2X1 U1747 ( .A(n7), .B(n1772), .C(n1834), .D(n1224), .Z(n1239) );
  CENX1 U1748 ( .A(n276), .B(n1831), .Z(n1554) );
  COND2X1 U1749 ( .A(n2387), .B(n1554), .C(n2388), .D(n1225), .Z(n1238) );
  CFA1X1 U1750 ( .A(n1228), .B(n1227), .CI(n1226), .CO(n1243), .S(
        \mult_x_1/n1145 ) );
  CFA1X1 U1751 ( .A(n1229), .B(n1230), .CI(n1231), .CO(n1242), .S(
        \mult_x_1/n1143 ) );
  CFA1X1 U1752 ( .A(n1232), .B(n1233), .CI(n1234), .CO(n2040), .S(n1231) );
  CFA1X1 U1753 ( .A(n1236), .B(n1237), .CI(n1235), .CO(n2039), .S(n1230) );
  CFA1X1 U1754 ( .A(n1240), .B(n1239), .CI(n1238), .CO(n2038), .S(n1229) );
  CFA1X1 U1755 ( .A(n1241), .B(n1242), .CI(n1243), .CO(\mult_x_1/n1112 ), .S(
        \mult_x_1/n1113 ) );
  CENX1 U1756 ( .A(n1600), .B(n1630), .Z(n1833) );
  CENX1 U1757 ( .A(n1600), .B(n1699), .Z(n1262) );
  COND2X1 U1758 ( .A(n2233), .B(n1833), .C(n269), .D(n1262), .Z(n2259) );
  CENX1 U1759 ( .A(n1695), .B(n1464), .Z(n1696) );
  CENX1 U1760 ( .A(n1695), .B(n1707), .Z(n1261) );
  COND2X1 U1761 ( .A(n2392), .B(n1696), .C(n2398), .D(n1261), .Z(n2258) );
  CENX1 U1762 ( .A(n1970), .B(n1466), .Z(n1724) );
  CENX1 U1763 ( .A(n1970), .B(n1694), .Z(n1245) );
  COND2X1 U1764 ( .A(n2440), .B(n1724), .C(n292), .D(n1245), .Z(n2257) );
  CENX1 U1765 ( .A(n11), .B(n1697), .Z(n1836) );
  CENX1 U1766 ( .A(n11), .B(n1961), .Z(n1247) );
  COND2X1 U1767 ( .A(n1920), .B(n1836), .C(n1244), .D(n1247), .Z(n1260) );
  CENX1 U1768 ( .A(n1975), .B(n1963), .Z(n1841) );
  CENX1 U1769 ( .A(n1975), .B(n1703), .Z(n1354) );
  COND2X1 U1770 ( .A(n14), .B(n1841), .C(n1842), .D(n1354), .Z(n1259) );
  CENX1 U1771 ( .A(n1848), .B(n1687), .Z(n1863) );
  CENX1 U1772 ( .A(n1848), .B(n1840), .Z(n1372) );
  COND2X1 U1773 ( .A(n2004), .B(n1863), .C(n2002), .D(n1372), .Z(n1258) );
  CNR2IX1 U1774 ( .B(n1714), .A(n2430), .Z(n1250) );
  CENX1 U1775 ( .A(n1970), .B(n1464), .Z(n1356) );
  COND2X1 U1776 ( .A(n2440), .B(n1245), .C(n292), .D(n1356), .Z(n1249) );
  CENX1 U1777 ( .A(n1692), .B(n1498), .Z(n1858) );
  CENX1 U1778 ( .A(n1692), .B(n1972), .Z(n1350) );
  COND2X1 U1779 ( .A(n1886), .B(n1858), .C(n1884), .D(n1350), .Z(n1248) );
  COND2X1 U1780 ( .A(n1920), .B(n1247), .C(n1918), .D(n1246), .Z(n2101) );
  CFA1X1 U1781 ( .A(n1250), .B(n1249), .CI(n1248), .CO(n2100), .S(n1255) );
  CENXL U1782 ( .A(n1711), .B(n1982), .Z(n1252) );
  COND2X1 U1783 ( .A(n2310), .B(n1252), .C(n2430), .D(n1251), .Z(n1360) );
  CND2IX1 U1784 ( .B(n1714), .A(n1982), .Z(n1253) );
  COND2X1 U1785 ( .A(n2432), .B(n1254), .C(n1253), .D(n2430), .Z(n1359) );
  CFA1X1 U1786 ( .A(n1257), .B(n1256), .CI(n1255), .CO(n1264), .S(
        \mult_x_1/n1423 ) );
  CFA1X1 U1787 ( .A(n1258), .B(n1259), .CI(n1260), .CO(n2098), .S(n1256) );
  CENX1 U1788 ( .A(n1718), .B(n2426), .Z(n1855) );
  CENX1 U1789 ( .A(n1718), .B(n1976), .Z(n1366) );
  COND2X1 U1790 ( .A(n1882), .B(n1855), .C(n18), .D(n1366), .Z(n2318) );
  CENX1 U1791 ( .A(n1388), .B(n1720), .Z(n1352) );
  COND2X1 U1792 ( .A(n2392), .B(n1261), .C(n2398), .D(n1352), .Z(n2317) );
  CENX1 U1793 ( .A(n1632), .B(n1712), .Z(n1343) );
  CENX1 U1794 ( .A(n1632), .B(n1466), .Z(n1358) );
  COND2X1 U1795 ( .A(n8), .B(n1343), .C(n2522), .D(n1358), .Z(n2316) );
  CENX1 U1796 ( .A(n1829), .B(n1811), .Z(n1860) );
  CENX1 U1797 ( .A(n1829), .B(n1717), .Z(n1368) );
  COND2X1 U1798 ( .A(n1893), .B(n1860), .C(n1861), .D(n1368), .Z(n2324) );
  CENX1 U1799 ( .A(n1600), .B(n1847), .Z(n1362) );
  COND2X1 U1800 ( .A(n7), .B(n1262), .C(n1834), .D(n1362), .Z(n2323) );
  CENX1 U1801 ( .A(n1721), .B(n1701), .Z(n1865) );
  CENX1 U1802 ( .A(n1721), .B(n1630), .Z(n1364) );
  CFA1X1 U1803 ( .A(n1265), .B(n1264), .CI(n1263), .CO(\mult_x_1/n1392 ), .S(
        \mult_x_1/n1393 ) );
  CFA1X1 U1804 ( .A(n1268), .B(n1267), .CI(n1266), .CO(n318), .S(
        \mult_x_1/n1117 ) );
  CFA1X1 U1805 ( .A(n1271), .B(n1270), .CI(n1269), .CO(\mult_x_1/n1692 ), .S(
        n1434) );
  CFA1X1 U1806 ( .A(n1274), .B(n1273), .CI(n1272), .CO(n342), .S(
        \mult_x_1/n883 ) );
  CFA1X1 U1807 ( .A(n1277), .B(n1276), .CI(n1275), .CO(\mult_x_1/n872 ), .S(
        n339) );
  CENX1 U1808 ( .A(n1695), .B(n1847), .Z(n1622) );
  CENX1 U1809 ( .A(n1388), .B(n1687), .Z(n1297) );
  COND2X1 U1810 ( .A(n2400), .B(n1622), .C(n2398), .D(n1297), .Z(n2178) );
  CENXL U1811 ( .A(n1977), .B(n1703), .Z(n1624) );
  CENXL U1812 ( .A(n1977), .B(n1981), .Z(n1287) );
  COND2X1 U1813 ( .A(n7), .B(n1624), .C(n269), .D(n1287), .Z(n2177) );
  CENX1 U1814 ( .A(n1975), .B(n1697), .Z(n1296) );
  COND2X1 U1815 ( .A(n14), .B(n1278), .C(n1842), .D(n1296), .Z(n2176) );
  CENX1 U1816 ( .A(n276), .B(n1840), .Z(n1626) );
  CENX1 U1817 ( .A(n276), .B(n1963), .Z(n1284) );
  COND2X1 U1818 ( .A(n255), .B(n1626), .C(n2388), .D(n1284), .Z(n1646) );
  CENX1 U1819 ( .A(n1843), .B(n2426), .Z(n1797) );
  COND2X1 U1820 ( .A(n6), .B(n1279), .C(n1924), .D(n1797), .Z(n1645) );
  CENX1 U1821 ( .A(n11), .B(n1976), .Z(n1628) );
  CENX1 U1822 ( .A(n11), .B(n1498), .Z(n1801) );
  COND2X1 U1823 ( .A(n1920), .B(n1628), .C(n1918), .D(n1801), .Z(n1644) );
  CENX1 U1824 ( .A(n1829), .B(n2393), .Z(n1286) );
  COND2X1 U1825 ( .A(n1893), .B(n1280), .C(n241), .D(n1286), .Z(n1649) );
  CENX1 U1826 ( .A(n1848), .B(n1831), .Z(n1285) );
  COND2X1 U1827 ( .A(n2004), .B(n1281), .C(n2002), .D(n1285), .Z(n1648) );
  CENXL U1828 ( .A(n1470), .B(n1965), .Z(n1288) );
  CENX1 U1829 ( .A(n1718), .B(n2389), .Z(n1819) );
  COND2X1 U1830 ( .A(n1882), .B(n1283), .C(n1880), .D(n1819), .Z(n1795) );
  CENX1 U1831 ( .A(n254), .B(n1694), .Z(n1642) );
  CENX1 U1832 ( .A(n254), .B(n1464), .Z(n1393) );
  COND2X1 U1833 ( .A(n245), .B(n1642), .C(n2406), .D(n1393), .Z(n1794) );
  CENX1 U1834 ( .A(n276), .B(n1703), .Z(n1397) );
  COND2X1 U1835 ( .A(n2387), .B(n1284), .C(n1722), .D(n1397), .Z(n1793) );
  CENX1 U1836 ( .A(n1677), .B(n1811), .Z(n1658) );
  CENX1 U1837 ( .A(n1677), .B(n1717), .Z(n1823) );
  COND2X1 U1838 ( .A(n246), .B(n1658), .C(n1967), .D(n1823), .Z(n1300) );
  CENX1 U1839 ( .A(n1848), .B(n1969), .Z(n1814) );
  COND2X1 U1840 ( .A(n1815), .B(n1285), .C(n2002), .D(n1814), .Z(n1299) );
  CENX1 U1841 ( .A(n1829), .B(n2469), .Z(n1821) );
  COND2X1 U1842 ( .A(n1893), .B(n1286), .C(n240), .D(n1821), .Z(n1298) );
  CENXL U1843 ( .A(n1977), .B(n1979), .Z(n1391) );
  COND2X1 U1844 ( .A(n2233), .B(n1287), .C(n1834), .D(n1391), .Z(n1804) );
  CAOR1X1 U1845 ( .A(n1884), .B(n1886), .C(n1288), .Z(n1803) );
  COND2X1 U1846 ( .A(n2310), .B(n1640), .C(n2430), .D(n1392), .Z(n1802) );
  CFA1X1 U1847 ( .A(n1292), .B(n1291), .CI(n1290), .CO(n1303), .S(
        \mult_x_1/n1259 ) );
  CFA1X1 U1848 ( .A(n1295), .B(n1294), .CI(n1293), .CO(n1302), .S(
        \mult_x_1/n1257 ) );
  CENX1 U1849 ( .A(n1637), .B(n1712), .Z(n1638) );
  CENX1 U1850 ( .A(n1637), .B(n1466), .Z(n1386) );
  COND2X1 U1851 ( .A(n2509), .B(n1638), .C(n1386), .D(n2510), .Z(n1657) );
  CENX1 U1852 ( .A(n1975), .B(n1961), .Z(n1825) );
  COND2X1 U1853 ( .A(n14), .B(n1296), .C(n1842), .D(n1825), .Z(n1656) );
  COR2X1 U1854 ( .A(n1657), .B(n1656), .Z(n2146) );
  CENX1 U1855 ( .A(n1388), .B(n1840), .Z(n1395) );
  COND2X1 U1856 ( .A(n2400), .B(n1297), .C(n2398), .D(n1395), .Z(n2202) );
  CENX1 U1857 ( .A(n1970), .B(n1699), .Z(n1659) );
  CENX1 U1858 ( .A(n1970), .B(n1847), .Z(n1399) );
  COND2X1 U1859 ( .A(n2440), .B(n1659), .C(n292), .D(n1399), .Z(n2201) );
  CENX1 U1860 ( .A(n2470), .B(n1701), .Z(n1662) );
  CENX1 U1861 ( .A(n1632), .B(n1630), .Z(n1817) );
  COND2X1 U1862 ( .A(n1662), .B(n8), .C(n2522), .D(n1817), .Z(n2200) );
  CFA1X1 U1863 ( .A(n1298), .B(n1299), .CI(n1300), .CO(n2144), .S(n1294) );
  CFA1X1 U1864 ( .A(n1303), .B(n1302), .CI(n1301), .CO(\mult_x_1/n1222 ), .S(
        \mult_x_1/n1223 ) );
  CENX1 U1865 ( .A(n1533), .B(n1831), .Z(n1472) );
  CENX1 U1866 ( .A(n1387), .B(n1969), .Z(n1311) );
  COND2X1 U1867 ( .A(n1857), .B(n1472), .C(n18), .D(n1311), .Z(n1480) );
  CENX1 U1868 ( .A(n1848), .B(n1707), .Z(n1465) );
  CENX1 U1869 ( .A(n1848), .B(n1720), .Z(n1318) );
  COND2X1 U1870 ( .A(n1815), .B(n1465), .C(n2002), .D(n1318), .Z(n1479) );
  CENX1 U1871 ( .A(n1721), .B(n1712), .Z(n1305) );
  COND2X1 U1872 ( .A(n255), .B(n1305), .C(n1722), .D(n1304), .Z(n1478) );
  CENX1 U1873 ( .A(n11), .B(n1963), .Z(n1468) );
  CENX1 U1874 ( .A(n11), .B(n1703), .Z(n1320) );
  COND2X1 U1875 ( .A(n1920), .B(n1468), .C(n1918), .D(n1320), .Z(n1753) );
  CENXL U1876 ( .A(n1711), .B(n276), .Z(n1306) );
  COND2X1 U1877 ( .A(n255), .B(n1306), .C(n1722), .D(n1305), .Z(n1741) );
  CND2IXL U1878 ( .B(n1714), .A(n276), .Z(n1307) );
  COND2X1 U1879 ( .A(n255), .B(n277), .C(n1307), .D(n1722), .Z(n1740) );
  CENX1 U1880 ( .A(n1843), .B(n1687), .Z(n1463) );
  COND2X1 U1881 ( .A(n6), .B(n1463), .C(n1924), .D(n1308), .Z(n1751) );
  CENX1 U1882 ( .A(n247), .B(n1981), .Z(n1474) );
  CENX1 U1883 ( .A(n247), .B(n1979), .Z(n1322) );
  COND2X1 U1884 ( .A(n1893), .B(n1474), .C(n1861), .D(n1322), .Z(n1483) );
  CENX1 U1885 ( .A(n1966), .B(n1847), .Z(n1314) );
  COND2X1 U1886 ( .A(n2050), .B(n1473), .C(n2051), .D(n1314), .Z(n1482) );
  COND2X1 U1887 ( .A(n1312), .B(n1311), .C(n1880), .D(n1310), .Z(n1339) );
  COND2X1 U1888 ( .A(n246), .B(n1314), .C(n1967), .D(n1313), .Z(n1338) );
  COND2X1 U1889 ( .A(n1886), .B(n1316), .C(n1884), .D(n1315), .Z(n1337) );
  COND2X1 U1890 ( .A(n2004), .B(n1318), .C(n2002), .D(n1317), .Z(n1336) );
  COND2X1 U1891 ( .A(n1920), .B(n1320), .C(n1877), .D(n1319), .Z(n1335) );
  COND2X1 U1892 ( .A(n1893), .B(n1322), .C(n1861), .D(n1321), .Z(n1334) );
  CFA1X1 U1893 ( .A(n1325), .B(n1324), .CI(n1323), .CO(n1168), .S(n1329) );
  CFA1X1 U1894 ( .A(n1328), .B(n1327), .CI(n1326), .CO(n1342), .S(
        \mult_x_1/n1533 ) );
  CFA1X1 U1895 ( .A(n1331), .B(n1330), .CI(n1329), .CO(n1341), .S(
        \mult_x_1/n1531 ) );
  CHA1X1 U1896 ( .A(n1333), .B(n1332), .CO(n1944), .S(n1490) );
  CFA1X1 U1897 ( .A(n1336), .B(n1335), .CI(n1334), .CO(n1943), .S(n1330) );
  CFA1X1 U1898 ( .A(n1337), .B(n1338), .CI(n1339), .CO(n1942), .S(n1331) );
  CFA1X1 U1899 ( .A(n1342), .B(n1341), .CI(n1340), .CO(\mult_x_1/n1508 ), .S(
        \mult_x_1/n1509 ) );
  CENX1 U1900 ( .A(n1838), .B(n1831), .Z(n1839) );
  CENX1 U1901 ( .A(n1843), .B(n1969), .Z(n1370) );
  COND2X1 U1902 ( .A(n6), .B(n1839), .C(n1924), .D(n1370), .Z(n2321) );
  CENXL U1903 ( .A(n1711), .B(n2470), .Z(n1344) );
  CND2IX1 U1904 ( .B(n1714), .A(n2470), .Z(n1345) );
  CENX1 U1905 ( .A(n1704), .B(n1981), .Z(n1853) );
  CENX1 U1906 ( .A(n1704), .B(n1979), .Z(n1348) );
  COND2X1 U1907 ( .A(n2050), .B(n1853), .C(n1967), .D(n1348), .Z(n2319) );
  COND2X1 U1908 ( .A(n2050), .B(n1348), .C(n2051), .D(n1347), .Z(n1376) );
  COND2X1 U1909 ( .A(n2055), .B(n1354), .C(n1842), .D(n1353), .Z(n1382) );
  COND2X1 U1910 ( .A(n1661), .B(n1356), .C(n292), .D(n1355), .Z(n1381) );
  COND2X1 U1911 ( .A(n9), .B(n1358), .C(n2522), .D(n1357), .Z(n1380) );
  CHA1X1 U1912 ( .A(n1360), .B(n1359), .CO(n1950), .S(n2099) );
  COND2X1 U1913 ( .A(n7), .B(n1362), .C(n1834), .D(n1361), .Z(n2119) );
  COND2X1 U1914 ( .A(n256), .B(n1364), .C(n2388), .D(n1363), .Z(n2118) );
  COND2X1 U1915 ( .A(n1882), .B(n1366), .C(n18), .D(n1365), .Z(n2117) );
  COND2X1 U1916 ( .A(n1893), .B(n1368), .C(n241), .D(n1367), .Z(n2125) );
  COND2X1 U1917 ( .A(n6), .B(n1370), .C(n1924), .D(n1369), .Z(n2124) );
  COND2X1 U1918 ( .A(n2004), .B(n1372), .C(n2002), .D(n1371), .Z(n2123) );
  CFA1X1 U1919 ( .A(n1375), .B(n1374), .CI(n1373), .CO(n1384), .S(
        \mult_x_1/n1397 ) );
  CFA1X1 U1920 ( .A(n1379), .B(n1378), .CI(n1377), .CO(n1672), .S(n1952) );
  CFA1X1 U1921 ( .A(n1382), .B(n1381), .CI(n1380), .CO(n1951), .S(n1373) );
  CFA1X1 U1922 ( .A(n1385), .B(n1384), .CI(n1383), .CO(\mult_x_1/n1366 ), .S(
        \mult_x_1/n1367 ) );
  CENX1 U1923 ( .A(n1637), .B(n1694), .Z(n1564) );
  COND2X1 U1924 ( .A(n2509), .B(n1386), .C(n1564), .D(n2510), .Z(n1406) );
  CAOR1X1 U1925 ( .A(n1880), .B(n1857), .C(n1818), .Z(n1405) );
  CENX1 U1926 ( .A(n1829), .B(n2441), .Z(n1820) );
  CENX1 U1927 ( .A(n1829), .B(n2389), .Z(n1777) );
  COND2X1 U1928 ( .A(n1893), .B(n1820), .C(n241), .D(n1777), .Z(n1404) );
  CENX1 U1929 ( .A(n1677), .B(n2426), .Z(n1822) );
  CENX1 U1930 ( .A(n1677), .B(n1976), .Z(n1557) );
  COND2X1 U1931 ( .A(n246), .B(n1822), .C(n2051), .D(n1557), .Z(n1569) );
  CENX1 U1932 ( .A(n1973), .B(n1697), .Z(n1813) );
  CENX1 U1933 ( .A(n1973), .B(n1961), .Z(n1559) );
  COND2X1 U1934 ( .A(n2004), .B(n1813), .C(n2002), .D(n1559), .Z(n1568) );
  CENXL U1935 ( .A(n1977), .B(n1831), .Z(n1390) );
  CENX1 U1936 ( .A(n1600), .B(n1969), .Z(n1773) );
  COND2X1 U1937 ( .A(n7), .B(n1390), .C(n1834), .D(n1773), .Z(n1567) );
  CENX1 U1938 ( .A(n276), .B(n1981), .Z(n1396) );
  CENX1 U1939 ( .A(n276), .B(n1979), .Z(n1555) );
  COND2X1 U1940 ( .A(n2387), .B(n1396), .C(n2388), .D(n1555), .Z(n1553) );
  CENX1 U1941 ( .A(n1970), .B(n1687), .Z(n1398) );
  CENX1 U1942 ( .A(n1970), .B(n1840), .Z(n1767) );
  COND2X1 U1943 ( .A(n1661), .B(n1398), .C(n292), .D(n1767), .Z(n1552) );
  CENX1 U1944 ( .A(n1388), .B(n1963), .Z(n1394) );
  COND2X1 U1945 ( .A(n2392), .B(n1394), .C(n2398), .D(n1389), .Z(n1551) );
  COND2X1 U1946 ( .A(n7), .B(n1391), .C(n1834), .D(n1390), .Z(n2284) );
  CENX1 U1947 ( .A(n1982), .B(n1701), .Z(n1573) );
  CENX1 U1948 ( .A(n254), .B(n1707), .Z(n1565) );
  CENX1 U1949 ( .A(n1843), .B(n1976), .Z(n1796) );
  CENX1 U1950 ( .A(n1843), .B(n1498), .Z(n1570) );
  COND2X1 U1951 ( .A(n6), .B(n1796), .C(n1924), .D(n1570), .Z(n2283) );
  CIVX2 U1952 ( .A(n1406), .Z(n2282) );
  CENX1 U1953 ( .A(n11), .B(n1972), .Z(n1800) );
  CENX1 U1954 ( .A(n11), .B(n2393), .Z(n1566) );
  COND2X1 U1955 ( .A(n1920), .B(n1800), .C(n1877), .D(n1566), .Z(n2281) );
  COND2X1 U1956 ( .A(n2400), .B(n1395), .C(n2398), .D(n1394), .Z(n2220) );
  COND2X1 U1957 ( .A(n255), .B(n1397), .C(n1722), .D(n1396), .Z(n2219) );
  COND2X1 U1958 ( .A(n1661), .B(n1399), .C(n292), .D(n1398), .Z(n2218) );
  CFA1X1 U1959 ( .A(n1400), .B(n1401), .CI(n1402), .CO(n1408), .S(
        \mult_x_1/n1199 ) );
  CENX1 U1960 ( .A(n1975), .B(n1717), .Z(n1812) );
  COND2X1 U1961 ( .A(n14), .B(n1812), .C(n2053), .D(n1403), .Z(n1576) );
  CFA1X1 U1962 ( .A(n1404), .B(n1406), .CI(n1405), .CO(n1575), .S(n1402) );
  CFA1X1 U1963 ( .A(n1409), .B(n1408), .CI(n1407), .CO(\mult_x_1/n1166 ), .S(
        \mult_x_1/n1167 ) );
  CFA1X1 U1964 ( .A(n1412), .B(n1411), .CI(n1410), .CO(n1432), .S(n411) );
  CENX1 U1965 ( .A(n1637), .B(n1840), .Z(n2013) );
  COND2X1 U1966 ( .A(n2509), .B(n2013), .C(n1413), .D(n2510), .Z(n2058) );
  CANR1X1 U1967 ( .A(n1842), .B(n13), .C(n1414), .Z(n2059) );
  CND2IXL U1968 ( .B(n2058), .A(n2059), .Z(n1416) );
  CENX1 U1969 ( .A(n1973), .B(n2389), .Z(n1504) );
  CND2X1 U1970 ( .A(n1416), .B(n2056), .Z(n1417) );
  COND2X1 U1971 ( .A(n9), .B(n1418), .C(n2522), .D(n1509), .Z(n2065) );
  CENX1 U1972 ( .A(n2390), .B(n1976), .Z(n1507) );
  COND2X1 U1973 ( .A(n2400), .B(n1419), .C(n2398), .D(n1507), .Z(n2064) );
  CENX1 U1974 ( .A(n2395), .B(n1717), .Z(n1502) );
  COND2X1 U1975 ( .A(n1661), .B(n1420), .C(n292), .D(n1502), .Z(n2063) );
  CFA1X1 U1976 ( .A(n1423), .B(n1422), .CI(n1421), .CO(n1510), .S(n1426) );
  CND2X1 U1977 ( .A(n1424), .B(n1426), .Z(n1429) );
  CND2X1 U1978 ( .A(n1424), .B(n1425), .Z(n1428) );
  CND3X2 U1979 ( .A(n1429), .B(n1428), .C(n1427), .Z(n1430) );
  CFA1X1 U1980 ( .A(n1432), .B(n1431), .CI(n1430), .CO(\mult_x_1/n942 ), .S(
        \mult_x_1/n943 ) );
  CNR2IX1 U1981 ( .B(n1714), .A(n1834), .Z(n1453) );
  CENX1 U1982 ( .A(n1975), .B(n1464), .Z(n1518) );
  COND2X1 U1983 ( .A(n2055), .B(n1435), .C(n1842), .D(n1518), .Z(n1452) );
  CENX1 U1984 ( .A(n1692), .B(n1979), .Z(n1536) );
  COND2X1 U1985 ( .A(n1886), .B(n1436), .C(n1884), .D(n1536), .Z(n1451) );
  CENX1 U1986 ( .A(n1718), .B(n1703), .Z(n1534) );
  COND2X1 U1987 ( .A(n1882), .B(n1437), .C(n18), .D(n1534), .Z(n1456) );
  CENX1 U1988 ( .A(n1966), .B(n1720), .Z(n1519) );
  COND2X1 U1989 ( .A(n2050), .B(n1438), .C(n2051), .D(n1519), .Z(n1455) );
  CENX1 U1990 ( .A(n1848), .B(n1466), .Z(n1520) );
  COND2X1 U1991 ( .A(n1815), .B(n1439), .C(n2002), .D(n1520), .Z(n1454) );
  CENX1 U1992 ( .A(n247), .B(n1840), .Z(n1443) );
  COND2X1 U1993 ( .A(n1893), .B(n1440), .C(n1861), .D(n1443), .Z(n1459) );
  CENXL U1994 ( .A(n11), .B(n1847), .Z(n1447) );
  COND2X1 U1995 ( .A(n1920), .B(n1441), .C(n1918), .D(n1447), .Z(n1458) );
  CENX1 U1996 ( .A(n1843), .B(n1630), .Z(n1532) );
  COND2X1 U1997 ( .A(n1926), .B(n1442), .C(n1924), .D(n1532), .Z(n1457) );
  CENX1 U1998 ( .A(n247), .B(n1963), .Z(n1522) );
  COND2X1 U1999 ( .A(n1893), .B(n1443), .C(n242), .D(n1522), .Z(n2077) );
  CENXL U2000 ( .A(n1714), .B(n1977), .Z(n1444) );
  CENX1 U2001 ( .A(n1600), .B(n1712), .Z(n1747) );
  CND2IXL U2002 ( .B(n1714), .A(n1977), .Z(n1445) );
  COND2X1 U2003 ( .A(n2233), .B(n1446), .C(n1445), .D(n1834), .Z(n1537) );
  CENXL U2004 ( .A(n11), .B(n1687), .Z(n1530) );
  COND2X1 U2005 ( .A(n1920), .B(n1447), .C(n1877), .D(n1530), .Z(n2075) );
  CFA1X1 U2006 ( .A(n1450), .B(n1449), .CI(n1448), .CO(n1461), .S(
        \mult_x_1/n1617 ) );
  CFA1X1 U2007 ( .A(n1453), .B(n1452), .CI(n1451), .CO(n2074), .S(n1450) );
  CFA1X1 U2008 ( .A(n1454), .B(n1455), .CI(n1456), .CO(n2073), .S(n1449) );
  CFA1X1 U2009 ( .A(n1459), .B(n1458), .CI(n1457), .CO(n2072), .S(n1448) );
  CFA1X1 U2010 ( .A(n1462), .B(n1461), .CI(n1460), .CO(\mult_x_1/n1598 ), .S(
        \mult_x_1/n1599 ) );
  CENX1 U2011 ( .A(n1843), .B(n1847), .Z(n1523) );
  COND2X1 U2012 ( .A(n6), .B(n1523), .C(n1924), .D(n1463), .Z(n1541) );
  CENX1 U2013 ( .A(n1848), .B(n1464), .Z(n1527) );
  COND2X1 U2014 ( .A(n2004), .B(n1527), .C(n2002), .D(n1465), .Z(n1540) );
  CENX1 U2015 ( .A(n1600), .B(n1466), .Z(n1746) );
  COND2X1 U2016 ( .A(n7), .B(n1746), .C(n1834), .D(n1467), .Z(n1539) );
  CENX1 U2017 ( .A(n11), .B(n1840), .Z(n1529) );
  COND2X1 U2018 ( .A(n1920), .B(n1529), .C(n1918), .D(n1468), .Z(n1738) );
  CENX1 U2019 ( .A(n1975), .B(n1720), .Z(n1744) );
  CENXL U2020 ( .A(n1470), .B(n1969), .Z(n1526) );
  CENX1 U2021 ( .A(n1533), .B(n1979), .Z(n1742) );
  COND2X1 U2022 ( .A(n1857), .B(n1742), .C(n18), .D(n1472), .Z(n1739) );
  CENX1 U2023 ( .A(n247), .B(n1703), .Z(n1521) );
  CFA1X1 U2024 ( .A(n1477), .B(n1476), .CI(n1475), .CO(n1491), .S(n1489) );
  CFA1X1 U2025 ( .A(n1480), .B(n1479), .CI(n1478), .CO(n1328), .S(n1488) );
  CFA1X1 U2026 ( .A(n1486), .B(n1485), .CI(n1484), .CO(n1494), .S(
        \mult_x_1/n1553 ) );
  CFA1X1 U2027 ( .A(n1492), .B(n1491), .CI(n1490), .CO(n1170), .S(n1493) );
  CENX1 U2028 ( .A(n1721), .B(n2393), .Z(n2234) );
  COND2X1 U2029 ( .A(n256), .B(n2234), .C(n2388), .D(n1495), .Z(n2382) );
  CENX1 U2030 ( .A(n2395), .B(n2426), .Z(n1501) );
  COND2X1 U2031 ( .A(n2440), .B(n1501), .C(n292), .D(n1496), .Z(n2381) );
  COND2X1 U2032 ( .A(n263), .B(n1508), .C(n2522), .D(n1497), .Z(n2380) );
  CENX1 U2033 ( .A(n2390), .B(n1498), .Z(n1506) );
  CENX1 U2034 ( .A(n254), .B(n1831), .Z(n2312) );
  COND2X1 U2035 ( .A(n2436), .B(n1500), .C(n2406), .D(n2312), .Z(n2238) );
  COND2X1 U2036 ( .A(n2440), .B(n1502), .C(n292), .D(n1501), .Z(n2237) );
  COND2X1 U2037 ( .A(n1815), .B(n1504), .C(n2002), .D(n1503), .Z(n2236) );
  CENX1 U2038 ( .A(n1982), .B(n1697), .Z(n2309) );
  COND2X1 U2039 ( .A(n2310), .B(n1505), .C(n2430), .D(n2309), .Z(n2229) );
  COND2X1 U2040 ( .A(n2400), .B(n1507), .C(n2398), .D(n1506), .Z(n2228) );
  COND2X1 U2041 ( .A(n9), .B(n1509), .C(n2522), .D(n1508), .Z(n2227) );
  CFA1X1 U2042 ( .A(n1514), .B(n1512), .CI(n1513), .CO(\mult_x_1/n926 ), .S(
        \mult_x_1/n927 ) );
  CFA1X1 U2043 ( .A(n1517), .B(n1516), .CI(n1515), .CO(n773), .S(
        \mult_x_1/n1069 ) );
  CENX1 U2044 ( .A(n1975), .B(n1707), .Z(n1745) );
  COND2X1 U2045 ( .A(n13), .B(n1518), .C(n2053), .D(n1745), .Z(n2083) );
  CENX1 U2046 ( .A(n1677), .B(n1701), .Z(n1525) );
  COND2X1 U2047 ( .A(n246), .B(n1519), .C(n2051), .D(n1525), .Z(n2082) );
  CENX1 U2048 ( .A(n1848), .B(n1694), .Z(n1528) );
  COND2X1 U2049 ( .A(n2004), .B(n1520), .C(n2002), .D(n1528), .Z(n2081) );
  COND2X1 U2050 ( .A(n1893), .B(n1522), .C(n241), .D(n1521), .Z(n1737) );
  CENX1 U2051 ( .A(n1843), .B(n1699), .Z(n1531) );
  COND2X1 U2052 ( .A(n6), .B(n1531), .C(n1924), .D(n1523), .Z(n1736) );
  COND2X1 U2053 ( .A(n246), .B(n1525), .C(n2051), .D(n1524), .Z(n1735) );
  CNR2IX1 U2054 ( .B(n1714), .A(n287), .Z(n1750) );
  CENX1 U2055 ( .A(n22), .B(n1831), .Z(n1535) );
  COND2X1 U2056 ( .A(n1886), .B(n1535), .C(n1884), .D(n1526), .Z(n1749) );
  COND2X1 U2057 ( .A(n1815), .B(n1528), .C(n2002), .D(n1527), .Z(n1748) );
  COND2X1 U2058 ( .A(n1920), .B(n1530), .C(n1877), .D(n1529), .Z(n1547) );
  COND2X1 U2059 ( .A(n6), .B(n1532), .C(n1924), .D(n1531), .Z(n2089) );
  CENX1 U2060 ( .A(n1533), .B(n1981), .Z(n1743) );
  COND2X1 U2061 ( .A(n1882), .B(n1534), .C(n18), .D(n1743), .Z(n2088) );
  COND2X1 U2062 ( .A(n1886), .B(n1536), .C(n1884), .D(n1535), .Z(n2087) );
  CFA1X1 U2063 ( .A(n1541), .B(n1540), .CI(n1539), .CO(n1486), .S(n1550) );
  CFA1X1 U2064 ( .A(n1544), .B(n1543), .CI(n1542), .CO(n1549), .S(
        \mult_x_1/n1587 ) );
  CFA1X1 U2065 ( .A(n1547), .B(n1546), .CI(n1545), .CO(n1548), .S(
        \mult_x_1/n1589 ) );
  CFA1X1 U2066 ( .A(n1550), .B(n1549), .CI(n1548), .CO(\mult_x_1/n1566 ), .S(
        \mult_x_1/n1567 ) );
  CFA1X1 U2067 ( .A(n1553), .B(n1552), .CI(n1551), .CO(n1579), .S(n1400) );
  COND2X1 U2068 ( .A(n256), .B(n1555), .C(n1722), .D(n1554), .Z(n1765) );
  COND2X1 U2069 ( .A(n246), .B(n1557), .C(n2051), .D(n1556), .Z(n1764) );
  COND2X1 U2070 ( .A(n2004), .B(n1559), .C(n2002), .D(n1558), .Z(n1763) );
  CFA1X1 U2071 ( .A(n1561), .B(n1562), .CI(n1560), .CO(n1228), .S(n1577) );
  COND2X1 U2072 ( .A(n2509), .B(n1564), .C(n1563), .D(n2510), .Z(n2143) );
  CENX1 U2073 ( .A(n254), .B(n1720), .Z(n1769) );
  COND2X1 U2074 ( .A(n245), .B(n1565), .C(n2434), .D(n1769), .Z(n2142) );
  CENX1 U2075 ( .A(n11), .B(n2469), .Z(n1775) );
  COND2X1 U2076 ( .A(n1920), .B(n1566), .C(n1918), .D(n1775), .Z(n2141) );
  CFA1X1 U2077 ( .A(n1569), .B(n1568), .CI(n1567), .CO(n1581), .S(n1401) );
  CENX1 U2078 ( .A(n1843), .B(n1972), .Z(n1771) );
  COND2X1 U2079 ( .A(n6), .B(n1570), .C(n1924), .D(n1771), .Z(n2149) );
  CENX1 U2080 ( .A(n1632), .B(n1699), .Z(n1816) );
  COND2X1 U2081 ( .A(n8), .B(n1816), .C(n2522), .D(n1571), .Z(n2148) );
  COND2X1 U2082 ( .A(n2310), .B(n1573), .C(n2430), .D(n1572), .Z(n2147) );
  CFA1X1 U2083 ( .A(n1576), .B(n1575), .CI(n1574), .CO(n1585), .S(n1407) );
  CFA1X1 U2084 ( .A(n1579), .B(n1578), .CI(n1577), .CO(n1584), .S(
        \mult_x_1/n1171 ) );
  CFA1X1 U2085 ( .A(n1582), .B(n1581), .CI(n1580), .CO(n1583), .S(
        \mult_x_1/n1173 ) );
  CFA1X1 U2086 ( .A(n1585), .B(n1584), .CI(n1583), .CO(\mult_x_1/n1140 ), .S(
        \mult_x_1/n1141 ) );
  CFA1X1 U2087 ( .A(n1588), .B(n1587), .CI(n1586), .CO(n1134), .S(n1594) );
  CFA1X1 U2088 ( .A(n1594), .B(n1593), .CI(n1592), .CO(\mult_x_1/n910 ), .S(
        \mult_x_1/n911 ) );
  CFA1X1 U2089 ( .A(n1597), .B(n1596), .CI(n1595), .CO(n1615), .S(n1515) );
  CENX1 U2090 ( .A(n1637), .B(n1699), .Z(n1602) );
  CENX1 U2091 ( .A(n2427), .B(n1847), .Z(n1612) );
  COND2X1 U2092 ( .A(n2509), .B(n1602), .C(n1612), .D(n2510), .Z(n1998) );
  CENX1 U2093 ( .A(n1982), .B(n1703), .Z(n1983) );
  COND2X1 U2094 ( .A(n2432), .B(n1598), .C(n2430), .D(n1983), .Z(n1997) );
  CENX1 U2095 ( .A(n254), .B(n1840), .Z(n1964) );
  COND2X1 U2096 ( .A(n245), .B(n1599), .C(n2406), .D(n1964), .Z(n1996) );
  CENX1 U2097 ( .A(n1600), .B(n2426), .Z(n2008) );
  COND2X1 U2098 ( .A(n2233), .B(n1601), .C(n1834), .D(n2008), .Z(n2172) );
  COND2X1 U2099 ( .A(n2509), .B(n1603), .C(n1602), .D(n2510), .Z(n2364) );
  CIVX2 U2100 ( .A(n2364), .Z(n2171) );
  CENX1 U2101 ( .A(n2390), .B(n1697), .Z(n2010) );
  COND2X1 U2102 ( .A(n2400), .B(n1604), .C(n2398), .D(n2010), .Z(n2170) );
  CFA1X1 U2103 ( .A(n1607), .B(n1606), .CI(n1605), .CO(n1618), .S(n774) );
  COND2X1 U2104 ( .A(n255), .B(n1609), .C(n287), .D(n1608), .Z(n2024) );
  CAOR1X1 U2105 ( .A(n1924), .B(n1926), .C(n1610), .Z(n2363) );
  CENX1 U2106 ( .A(n1677), .B(n2389), .Z(n1968) );
  COND2X1 U2107 ( .A(n2050), .B(n1611), .C(n1967), .D(n1968), .Z(n2362) );
  CENX1 U2108 ( .A(n1637), .B(n1687), .Z(n2014) );
  COND2X1 U2109 ( .A(n239), .B(n1612), .C(n2014), .D(n2510), .Z(n2352) );
  CIVX1 U2110 ( .A(n2352), .Z(n2022) );
  CFA1X1 U2111 ( .A(n1615), .B(n1614), .CI(n1613), .CO(n1616), .S(
        \mult_x_1/n1047 ) );
  CFA1X1 U2112 ( .A(n1618), .B(n1617), .CI(n1616), .CO(\mult_x_1/n1020 ), .S(
        \mult_x_1/n1021 ) );
  CFA1X1 U2113 ( .A(n1621), .B(n1620), .CI(n1619), .CO(n770), .S(
        \mult_x_1/n1631 ) );
  COND2X1 U2114 ( .A(n2400), .B(n1623), .C(n2398), .D(n1622), .Z(n2244) );
  COND2X1 U2115 ( .A(n2233), .B(n1625), .C(n269), .D(n1624), .Z(n2243) );
  COND2X1 U2116 ( .A(n255), .B(n1627), .C(n2388), .D(n1626), .Z(n2242) );
  COND2X1 U2117 ( .A(n1920), .B(n1629), .C(n1877), .D(n1628), .Z(n2250) );
  CENX1 U2118 ( .A(n1970), .B(n1630), .Z(n1660) );
  COND2X1 U2119 ( .A(n2440), .B(n1631), .C(n292), .D(n1660), .Z(n2249) );
  CENX1 U2120 ( .A(n1632), .B(n1720), .Z(n1663) );
  COND2X1 U2121 ( .A(n9), .B(n1633), .C(n2522), .D(n1663), .Z(n2248) );
  CFA1X1 U2122 ( .A(n1636), .B(n1635), .CI(n1634), .CO(n1650), .S(n538) );
  CENXL U2123 ( .A(n1711), .B(n1637), .Z(n1639) );
  COND2X1 U2124 ( .A(n2509), .B(n1639), .C(n1638), .D(n2510), .Z(n1666) );
  COND2X1 U2125 ( .A(n2310), .B(n1641), .C(n2430), .D(n1640), .Z(n1665) );
  CFA1X1 U2126 ( .A(n1646), .B(n1645), .CI(n1644), .CO(n1291), .S(n1654) );
  CFA1X1 U2127 ( .A(n1649), .B(n1648), .CI(n1647), .CO(n1290), .S(n1653) );
  CFA1X1 U2128 ( .A(n1652), .B(n1651), .CI(n1650), .CO(n1669), .S(
        \mult_x_1/n1289 ) );
  CFA1X1 U2129 ( .A(n1655), .B(n1654), .CI(n1653), .CO(n1668), .S(
        \mult_x_1/n1287 ) );
  CENX1 U2130 ( .A(n1657), .B(n1656), .Z(n2217) );
  CENX1 U2131 ( .A(n1677), .B(n1961), .Z(n1678) );
  COND2X1 U2132 ( .A(n2050), .B(n1678), .C(n2051), .D(n1658), .Z(n2184) );
  COND2X1 U2133 ( .A(n1661), .B(n1660), .C(n292), .D(n1659), .Z(n2183) );
  COND2X1 U2134 ( .A(n8), .B(n1663), .C(n2522), .D(n1662), .Z(n2182) );
  CFA1X1 U2135 ( .A(n1666), .B(n1665), .CI(n1664), .CO(n2215), .S(n1655) );
  CFA1X1 U2136 ( .A(n1669), .B(n1668), .CI(n1667), .CO(\mult_x_1/n1252 ), .S(
        \mult_x_1/n1253 ) );
  CFA1X1 U2137 ( .A(n1672), .B(n1671), .CI(n1670), .CO(n1686), .S(n386) );
  CND2X1 U2138 ( .A(n1673), .B(n1675), .Z(n1676) );
  CENX1 U2139 ( .A(n1677), .B(n1697), .Z(n1956) );
  COND2X1 U2140 ( .A(n246), .B(n1956), .C(n2051), .D(n1678), .Z(n2181) );
  CFA1X1 U2141 ( .A(n1681), .B(n1680), .CI(n1679), .CO(n2180), .S(n1675) );
  CND2IX1 U2142 ( .B(n1714), .A(n254), .Z(n1683) );
  CENX1 U2143 ( .A(n1975), .B(n1687), .Z(n1846) );
  COND2X1 U2144 ( .A(n14), .B(n1688), .C(n1842), .D(n1846), .Z(n2343) );
  CENX1 U2145 ( .A(n1718), .B(n1811), .Z(n1719) );
  COND2X1 U2146 ( .A(n1882), .B(n1689), .C(n18), .D(n1719), .Z(n2342) );
  CENX1 U2147 ( .A(n21), .B(n2426), .Z(n1693) );
  COND2X1 U2148 ( .A(n1886), .B(n1691), .C(n1884), .D(n1693), .Z(n2341) );
  CNR2IX1 U2149 ( .B(n1714), .A(n2522), .Z(n1728) );
  CENX1 U2150 ( .A(n1692), .B(n1976), .Z(n1859) );
  COND2X1 U2151 ( .A(n1886), .B(n1693), .C(n1884), .D(n1859), .Z(n1727) );
  CENX1 U2152 ( .A(n1695), .B(n1694), .Z(n1709) );
  COND2X1 U2153 ( .A(n2392), .B(n1709), .C(n2398), .D(n1696), .Z(n1726) );
  CENX1 U2154 ( .A(n1829), .B(n1697), .Z(n1830) );
  COND2X1 U2155 ( .A(n1893), .B(n1698), .C(n1861), .D(n1830), .Z(n2346) );
  CENX1 U2156 ( .A(n1848), .B(n1699), .Z(n1849) );
  COND2X1 U2157 ( .A(n1815), .B(n1700), .C(n2002), .D(n1849), .Z(n2345) );
  CENXL U2158 ( .A(n1977), .B(n1701), .Z(n1835) );
  COND2X1 U2159 ( .A(n7), .B(n1702), .C(n269), .D(n1835), .Z(n2344) );
  CENX1 U2160 ( .A(n1704), .B(n1963), .Z(n1705) );
  CENX1 U2161 ( .A(n1704), .B(n1703), .Z(n1854) );
  COND2X1 U2162 ( .A(n246), .B(n1705), .C(n1967), .D(n1854), .Z(n1929) );
  COND2X1 U2163 ( .A(n2050), .B(n1706), .C(n1967), .D(n1705), .Z(n1938) );
  CENX1 U2164 ( .A(n1721), .B(n1707), .Z(n1723) );
  COND2X1 U2165 ( .A(n255), .B(n1708), .C(n287), .D(n1723), .Z(n1937) );
  COND2X1 U2166 ( .A(n2400), .B(n1710), .C(n2398), .D(n1709), .Z(n1936) );
  CENXL U2167 ( .A(n1711), .B(n2395), .Z(n1713) );
  CENX1 U2168 ( .A(n1970), .B(n1712), .Z(n1725) );
  COND2X1 U2169 ( .A(n2440), .B(n1713), .C(n292), .D(n1725), .Z(n1922) );
  CND2IX1 U2170 ( .B(n1714), .A(n1970), .Z(n1715) );
  COND2X1 U2171 ( .A(n2440), .B(n1716), .C(n1715), .D(n292), .Z(n1921) );
  CENX1 U2172 ( .A(n1718), .B(n1717), .Z(n1856) );
  COND2X1 U2173 ( .A(n1857), .B(n1719), .C(n18), .D(n1856), .Z(n2296) );
  CENX1 U2174 ( .A(n1721), .B(n1720), .Z(n1866) );
  COND2X1 U2175 ( .A(n255), .B(n1723), .C(n1722), .D(n1866), .Z(n2295) );
  COND2X1 U2176 ( .A(n2440), .B(n1725), .C(n292), .D(n1724), .Z(n2294) );
  CFA1X1 U2177 ( .A(n1728), .B(n1727), .CI(n1726), .CO(n1850), .S(n1730) );
  CFA1X1 U2178 ( .A(n1731), .B(n1730), .CI(n1729), .CO(n1732), .S(
        \mult_x_1/n1471 ) );
  CFA1X1 U2179 ( .A(n1734), .B(n1733), .CI(n1732), .CO(\mult_x_1/n1442 ), .S(
        \mult_x_1/n1443 ) );
  CFA1X1 U2180 ( .A(n1737), .B(n1736), .CI(n1735), .CO(n1756), .S(n1543) );
  CHA1X1 U2181 ( .A(n1741), .B(n1740), .CO(n1752), .S(n1759) );
  COND2X1 U2182 ( .A(n1882), .B(n1743), .C(n18), .D(n1742), .Z(n2071) );
  COND2XL U2183 ( .A(n13), .B(n1745), .C(n1842), .D(n1744), .Z(n2070) );
  COND2X1 U2184 ( .A(n2233), .B(n1747), .C(n269), .D(n1746), .Z(n2069) );
  CFA1X1 U2185 ( .A(n1750), .B(n1749), .CI(n1748), .CO(n1757), .S(n1542) );
  CFA1X1 U2186 ( .A(n1753), .B(n1752), .CI(n1751), .CO(n1327), .S(n1762) );
  CFA1X1 U2187 ( .A(n1756), .B(n1755), .CI(n1754), .CO(n1761), .S(
        \mult_x_1/n1569 ) );
  CFA1X1 U2188 ( .A(n1759), .B(n1758), .CI(n1757), .CO(n1760), .S(
        \mult_x_1/n1571 ) );
  CFA1X1 U2189 ( .A(n1762), .B(n1761), .CI(n1760), .CO(\mult_x_1/n1548 ), .S(
        \mult_x_1/n1549 ) );
  CFA1X1 U2190 ( .A(n1765), .B(n1764), .CI(n1763), .CO(n1789), .S(n1578) );
  COND2X1 U2191 ( .A(n2440), .B(n1767), .C(n292), .D(n1766), .Z(n2107) );
  COND2X1 U2192 ( .A(n245), .B(n1769), .C(n2434), .D(n1768), .Z(n2106) );
  COND2X1 U2193 ( .A(n6), .B(n1771), .C(n1924), .D(n1770), .Z(n2105) );
  COND2X1 U2194 ( .A(n7), .B(n1773), .C(n1834), .D(n1772), .Z(n2113) );
  COND2X1 U2195 ( .A(n1920), .B(n1775), .C(n1918), .D(n1774), .Z(n2112) );
  COND2X1 U2196 ( .A(n1893), .B(n1777), .C(n241), .D(n1776), .Z(n2111) );
  CFA1X1 U2197 ( .A(n1780), .B(n1779), .CI(n1778), .CO(n1192), .S(n1792) );
  CFA1X1 U2198 ( .A(n1783), .B(n1782), .CI(n1781), .CO(n2042), .S(n1226) );
  CFA1X1 U2199 ( .A(n1786), .B(n1785), .CI(n1784), .CO(n2041), .S(n1227) );
  CFA1X1 U2200 ( .A(n1789), .B(n1788), .CI(n1787), .CO(n1790), .S(
        \mult_x_1/n1147 ) );
  CFA1X1 U2201 ( .A(n1792), .B(n1791), .CI(n1790), .CO(\mult_x_1/n1114 ), .S(
        \mult_x_1/n1115 ) );
  CFA1X1 U2202 ( .A(n1795), .B(n1794), .CI(n1793), .CO(n1807), .S(n1295) );
  COND2X1 U2203 ( .A(n6), .B(n1797), .C(n1924), .D(n1796), .Z(n2208) );
  CHA1X1 U2204 ( .A(n1799), .B(n1798), .CO(n2207), .S(n2205) );
  COND2X1 U2205 ( .A(n1920), .B(n1801), .C(n1918), .D(n1800), .Z(n2206) );
  CFA1X1 U2206 ( .A(n1804), .B(n1803), .CI(n1802), .CO(n1805), .S(n1293) );
  CFA1X1 U2207 ( .A(n1807), .B(n1806), .CI(n1805), .CO(n1828), .S(
        \mult_x_1/n1229 ) );
  CFA1X1 U2208 ( .A(n1810), .B(n1809), .CI(n1808), .CO(n1409), .S(n1827) );
  CENX1 U2209 ( .A(n1975), .B(n1811), .Z(n1824) );
  COND2XL U2210 ( .A(n13), .B(n1824), .C(n1842), .D(n1812), .Z(n2110) );
  COND2X1 U2211 ( .A(n1815), .B(n1814), .C(n2002), .D(n1813), .Z(n2280) );
  COND2X1 U2212 ( .A(n9), .B(n1817), .C(n2522), .D(n1816), .Z(n2279) );
  COND2X1 U2213 ( .A(n1882), .B(n1819), .C(n18), .D(n244), .Z(n2278) );
  COND2X1 U2214 ( .A(n1893), .B(n1821), .C(n1861), .D(n1820), .Z(n2214) );
  COND2X1 U2215 ( .A(n2050), .B(n1823), .C(n2051), .D(n1822), .Z(n2213) );
  COND2X1 U2216 ( .A(n2055), .B(n1825), .C(n1842), .D(n1824), .Z(n2212) );
  CFA1X1 U2217 ( .A(n1828), .B(n1827), .CI(n1826), .CO(\mult_x_1/n1194 ), .S(
        \mult_x_1/n1195 ) );
  CENX1 U2218 ( .A(n1829), .B(n1961), .Z(n1862) );
  COND2X1 U2219 ( .A(n1893), .B(n1830), .C(n241), .D(n1862), .Z(n2293) );
  CENX1 U2220 ( .A(n11), .B(n1831), .Z(n1917) );
  CENXL U2221 ( .A(n11), .B(n1969), .Z(n1837) );
  COND2X1 U2222 ( .A(n1920), .B(n1917), .C(n1877), .D(n1837), .Z(n2292) );
  COND2X1 U2223 ( .A(n2233), .B(n1835), .C(n1834), .D(n1833), .Z(n2291) );
  COND2X1 U2224 ( .A(n1920), .B(n1837), .C(n1877), .D(n1836), .Z(n1869) );
  CENX1 U2225 ( .A(n1838), .B(n1979), .Z(n1844) );
  COND2X1 U2226 ( .A(n1926), .B(n1844), .C(n1924), .D(n1839), .Z(n1868) );
  CENX1 U2227 ( .A(n1975), .B(n1840), .Z(n1845) );
  COND2X1 U2228 ( .A(n13), .B(n1845), .C(n1842), .D(n1841), .Z(n1867) );
  CENX1 U2229 ( .A(n1843), .B(n1981), .Z(n1923) );
  COND2X1 U2230 ( .A(n6), .B(n1923), .C(n1924), .D(n1844), .Z(n2290) );
  COND2X1 U2231 ( .A(n14), .B(n1846), .C(n2053), .D(n1845), .Z(n2289) );
  CENX1 U2232 ( .A(n1848), .B(n1847), .Z(n1864) );
  COND2X1 U2233 ( .A(n1815), .B(n1849), .C(n2002), .D(n1864), .Z(n2288) );
  CFA1X1 U2234 ( .A(n1852), .B(n1851), .CI(n1850), .CO(n1875), .S(n1733) );
  COND2X1 U2235 ( .A(n2050), .B(n1854), .C(n2051), .D(n1853), .Z(n2262) );
  COND2X1 U2236 ( .A(n1857), .B(n1856), .C(n18), .D(n1855), .Z(n2261) );
  COND2X1 U2237 ( .A(n1886), .B(n1859), .C(n1884), .D(n1858), .Z(n2260) );
  COND2X1 U2238 ( .A(n1893), .B(n1862), .C(n1861), .D(n1860), .Z(n2256) );
  COND2X1 U2239 ( .A(n1815), .B(n1864), .C(n2002), .D(n1863), .Z(n2255) );
  COND2X1 U2240 ( .A(n256), .B(n1866), .C(n287), .D(n1865), .Z(n2254) );
  CFA1X1 U2241 ( .A(n1868), .B(n1869), .CI(n1867), .CO(n2120), .S(n1871) );
  CFA1X1 U2242 ( .A(n1872), .B(n1871), .CI(n1870), .CO(n1873), .S(
        \mult_x_1/n1447 ) );
  CFA1X1 U2243 ( .A(n1875), .B(n1874), .CI(n1873), .CO(\mult_x_1/n1418 ), .S(
        \mult_x_1/n1419 ) );
  COND2X1 U2244 ( .A(n1920), .B(n1878), .C(n1877), .D(n1876), .Z(n2196) );
  COND2X1 U2245 ( .A(n1882), .B(n1881), .C(n18), .D(n1879), .Z(n2195) );
  COND2X1 U2246 ( .A(n1886), .B(n1885), .C(n1884), .D(n1883), .Z(n2194) );
  CFA1X1 U2247 ( .A(n1889), .B(n1888), .CI(n1887), .CO(n1902), .S(n1905) );
  COND2X1 U2248 ( .A(n1893), .B(n1892), .C(n242), .D(n1890), .Z(n2190) );
  COND2X1 U2249 ( .A(n6), .B(n1895), .C(n1924), .D(n1894), .Z(n2189) );
  COND2X1 U2250 ( .A(n2050), .B(n1897), .C(n1967), .D(n1896), .Z(n2188) );
  CFA1X1 U2251 ( .A(n1900), .B(n1899), .CI(n1898), .CO(n2084), .S(n1909) );
  CFA1X1 U2252 ( .A(n1903), .B(n1902), .CI(n1901), .CO(n772), .S(n1908) );
  CFA1X1 U2253 ( .A(n1906), .B(n1905), .CI(n1904), .CO(n1907), .S(
        \mult_x_1/n1645 ) );
  CFA1X1 U2254 ( .A(n1909), .B(n1907), .CI(n1908), .CO(\mult_x_1/n1628 ), .S(
        \mult_x_1/n1629 ) );
  CNR2X1 U2255 ( .A(n1911), .B(n1910), .Z(\mult_x_1/n700 ) );
  CNIVX1 U2256 ( .A(n1912), .Z(n1916) );
  CND2X1 U2257 ( .A(n1914), .B(n1913), .Z(n1915) );
  CENX1 U2258 ( .A(n1916), .B(n1915), .Z(n2891) );
  COND2X1 U2259 ( .A(n1920), .B(n1919), .C(n1918), .D(n1917), .Z(n1941) );
  CHA1X1 U2260 ( .A(n1922), .B(n1921), .CO(n1927), .S(n1940) );
  COND2X1 U2261 ( .A(n6), .B(n1925), .C(n1924), .D(n1923), .Z(n1939) );
  CFA1X1 U2262 ( .A(n1929), .B(n1928), .CI(n1927), .CO(n1734), .S(n1934) );
  CFA1X1 U2263 ( .A(n1932), .B(n1931), .CI(n1930), .CO(n1933), .S(n1181) );
  CFA1X1 U2264 ( .A(n1935), .B(n1934), .CI(n1933), .CO(\mult_x_1/n1466 ), .S(
        \mult_x_1/n1467 ) );
  CFA1X1 U2265 ( .A(n1938), .B(n1937), .CI(n1936), .CO(n1928), .S(n1947) );
  CFA1X1 U2266 ( .A(n1941), .B(n1940), .CI(n1939), .CO(n1935), .S(n1946) );
  CFA1X1 U2267 ( .A(n1944), .B(n1943), .CI(n1942), .CO(n1945), .S(n1340) );
  CFA1X1 U2268 ( .A(n1947), .B(n1946), .CI(n1945), .CO(\mult_x_1/n1488 ), .S(
        \mult_x_1/n1489 ) );
  CFA1X1 U2269 ( .A(n1950), .B(n1948), .CI(n1949), .CO(n1960), .S(n1385) );
  CFA1X1 U2270 ( .A(n1953), .B(n1952), .CI(n1951), .CO(n1959), .S(n1383) );
  COND2X1 U2271 ( .A(n2004), .B(n1955), .C(n2002), .D(n1954), .Z(n2247) );
  COND2X1 U2272 ( .A(n2050), .B(n1957), .C(n1967), .D(n1956), .Z(n2245) );
  CFA1X1 U2273 ( .A(n1960), .B(n1958), .CI(n1959), .CO(\mult_x_1/n1340 ), .S(
        \mult_x_1/n1341 ) );
  CENX1 U2274 ( .A(n2390), .B(n1961), .Z(n2009) );
  COND2X1 U2275 ( .A(n2400), .B(n2009), .C(n2398), .D(n1962), .Z(n2274) );
  CENX1 U2276 ( .A(n254), .B(n1963), .Z(n2018) );
  COND2X1 U2277 ( .A(n245), .B(n1964), .C(n2434), .D(n2018), .Z(n2273) );
  COND2X1 U2278 ( .A(n246), .B(n1968), .C(n1967), .D(n2049), .Z(n2272) );
  CENX1 U2279 ( .A(n1970), .B(n1969), .Z(n2011) );
  COND2X1 U2280 ( .A(n2440), .B(n2011), .C(n292), .D(n1971), .Z(n2271) );
  CENX1 U2281 ( .A(n1973), .B(n1972), .Z(n2001) );
  COND2X1 U2282 ( .A(n1815), .B(n2001), .C(n2002), .D(n1974), .Z(n2270) );
  CENX1 U2283 ( .A(n1975), .B(n2469), .Z(n1999) );
  CENX1 U2284 ( .A(n1975), .B(n2441), .Z(n2054) );
  COND2X1 U2285 ( .A(n14), .B(n1999), .C(n2053), .D(n2054), .Z(n2269) );
  CENXL U2286 ( .A(n1977), .B(n1976), .Z(n2007) );
  COND2X1 U2287 ( .A(n2233), .B(n2007), .C(n269), .D(n1978), .Z(n2268) );
  CENX1 U2288 ( .A(n2470), .B(n1979), .Z(n2005) );
  CENX1 U2289 ( .A(n1982), .B(n1981), .Z(n2016) );
  COND2X1 U2290 ( .A(n2310), .B(n1983), .C(n2430), .D(n2016), .Z(n2266) );
  CFA1X1 U2291 ( .A(n1986), .B(n1985), .CI(n1984), .CO(n1424), .S(n1995) );
  CFA1X1 U2292 ( .A(n1989), .B(n1988), .CI(n1987), .CO(n1994), .S(
        \mult_x_1/n1005 ) );
  CFA1X1 U2293 ( .A(n1992), .B(n1991), .CI(n1990), .CO(n1411), .S(n1993) );
  CFA1X1 U2294 ( .A(n1995), .B(n1994), .CI(n1993), .CO(\mult_x_1/n980 ), .S(
        \mult_x_1/n981 ) );
  CFA1X1 U2295 ( .A(n1998), .B(n1996), .CI(n1997), .CO(n2021), .S(n1614) );
  COND2X1 U2296 ( .A(n14), .B(n2000), .C(n2053), .D(n1999), .Z(n2370) );
  COND2X1 U2297 ( .A(n2004), .B(n2003), .C(n2002), .D(n2001), .Z(n2369) );
  COND2X1 U2298 ( .A(n8), .B(n2006), .C(n2522), .D(n2005), .Z(n2368) );
  COND2X1 U2299 ( .A(n7), .B(n2008), .C(n269), .D(n2007), .Z(n2367) );
  COND2X1 U2300 ( .A(n2400), .B(n2010), .C(n2398), .D(n2009), .Z(n2366) );
  COND2X1 U2301 ( .A(n2440), .B(n2012), .C(n292), .D(n2011), .Z(n2365) );
  COND2X1 U2302 ( .A(n239), .B(n2014), .C(n2013), .D(n2510), .Z(n2048) );
  COND2X1 U2303 ( .A(n2432), .B(n2016), .C(n2430), .D(n2015), .Z(n2047) );
  COND2X1 U2304 ( .A(n245), .B(n2018), .C(n2434), .D(n2017), .Z(n2046) );
  CFA1X1 U2305 ( .A(n2021), .B(n2020), .CI(n2019), .CO(n2026), .S(
        \mult_x_1/n1025 ) );
  CFA1X1 U2306 ( .A(n2024), .B(n2023), .CI(n2022), .CO(n2025), .S(n1617) );
  CFA1X1 U2307 ( .A(n2027), .B(n2026), .CI(n2025), .CO(\mult_x_1/n1000 ), .S(
        \mult_x_1/n1001 ) );
  CIVXL U2308 ( .A(n2543), .Z(n2028) );
  CIVXL U2309 ( .A(n2029), .Z(n2542) );
  CIVXL U2310 ( .A(n2030), .Z(n2540) );
  CFA1X1 U2311 ( .A(n2037), .B(n2036), .CI(n2035), .CO(n1200), .S(n2045) );
  CFA1X1 U2312 ( .A(n2040), .B(n2039), .CI(n2038), .CO(n2044), .S(n1241) );
  CFA1X1 U2313 ( .A(n2045), .B(n2044), .CI(n2043), .CO(\mult_x_1/n1090 ), .S(
        \mult_x_1/n1091 ) );
  CIVX1 U2314 ( .A(n2058), .Z(n2062) );
  CFA1X1 U2315 ( .A(n2048), .B(n2047), .CI(n2046), .CO(n2061), .S(n2027) );
  COND2X1 U2316 ( .A(n14), .B(n2054), .C(n2053), .D(n2052), .Z(n2350) );
  CIVXL U2317 ( .A(n2056), .Z(n2057) );
  CEO3XL U2318 ( .A(n2059), .B(n2058), .C(n2057), .Z(n2068) );
  CFA1X1 U2319 ( .A(n2062), .B(n2061), .CI(n2060), .CO(n2067), .S(
        \mult_x_1/n985 ) );
  CFA1X1 U2320 ( .A(n2065), .B(n2064), .CI(n2063), .CO(n1511), .S(n2066) );
  CFA1X1 U2321 ( .A(n2068), .B(n2067), .CI(n2066), .CO(\mult_x_1/n962 ), .S(
        \mult_x_1/n963 ) );
  CFA1X1 U2322 ( .A(n2071), .B(n2070), .CI(n2069), .CO(n1758), .S(n2080) );
  CFA1X1 U2323 ( .A(n2074), .B(n2073), .CI(n2072), .CO(n2079), .S(n1460) );
  CFA1X1 U2324 ( .A(n2077), .B(n2076), .CI(n2075), .CO(n2078), .S(n1462) );
  CFA1X1 U2325 ( .A(n2080), .B(n2079), .CI(n2078), .CO(\mult_x_1/n1584 ), .S(
        \mult_x_1/n1585 ) );
  CFA1X1 U2326 ( .A(n2083), .B(n2082), .CI(n2081), .CO(n1544), .S(n2092) );
  CFA1X1 U2327 ( .A(n2086), .B(n2085), .CI(n2084), .CO(n2091), .S(n771) );
  CFA1X1 U2328 ( .A(n2089), .B(n2088), .CI(n2087), .CO(n1546), .S(n2090) );
  CFA1X1 U2329 ( .A(n2092), .B(n2091), .CI(n2090), .CO(\mult_x_1/n1600 ), .S(
        \mult_x_1/n1601 ) );
  CFA1X1 U2330 ( .A(n2095), .B(n2094), .CI(n2093), .CO(n1673), .S(n2104) );
  CFA1X1 U2331 ( .A(n2096), .B(n2098), .CI(n2097), .CO(n2103), .S(n1263) );
  CFA1X1 U2332 ( .A(n2101), .B(n2100), .CI(n2099), .CO(n2102), .S(n1265) );
  CFA1X1 U2333 ( .A(n2104), .B(n2103), .CI(n2102), .CO(\mult_x_1/n1368 ), .S(
        \mult_x_1/n1369 ) );
  CFA1X1 U2334 ( .A(n2107), .B(n2106), .CI(n2105), .CO(n1788), .S(n2116) );
  CFA1X1 U2335 ( .A(n2110), .B(n2109), .CI(n2108), .CO(n2115), .S(n1826) );
  CFA1X1 U2336 ( .A(n2113), .B(n2112), .CI(n2111), .CO(n1787), .S(n2114) );
  CFA1X1 U2337 ( .A(n2116), .B(n2115), .CI(n2114), .CO(\mult_x_1/n1168 ), .S(
        \mult_x_1/n1169 ) );
  CFA1X1 U2338 ( .A(n2119), .B(n2118), .CI(n2117), .CO(n1949), .S(n2128) );
  CFA1X1 U2339 ( .A(n2122), .B(n2121), .CI(n2120), .CO(n2127), .S(n1874) );
  CFA1X1 U2340 ( .A(n2125), .B(n2123), .CI(n2124), .CO(n1948), .S(n2126) );
  CFA1X1 U2341 ( .A(n2128), .B(n2127), .CI(n2126), .CO(\mult_x_1/n1394 ), .S(
        \mult_x_1/n1395 ) );
  CFA1X1 U2342 ( .A(n2131), .B(n2130), .CI(n2129), .CO(n1621), .S(n2140) );
  CFA1X1 U2343 ( .A(n2134), .B(n2133), .CI(n2132), .CO(n2139), .S(
        \mult_x_1/n1657 ) );
  CFA1X1 U2344 ( .A(n2137), .B(n2136), .CI(n2135), .CO(n1619), .S(n2138) );
  CFA1X1 U2345 ( .A(n2140), .B(n2139), .CI(n2138), .CO(\mult_x_1/n1642 ), .S(
        \mult_x_1/n1643 ) );
  CFA1X1 U2346 ( .A(n2143), .B(n2142), .CI(n2141), .CO(n1582), .S(n2152) );
  CFA1X1 U2347 ( .A(n2146), .B(n2145), .CI(n2144), .CO(n2151), .S(n1301) );
  CFA1X1 U2348 ( .A(n2149), .B(n2148), .CI(n2147), .CO(n1580), .S(n2150) );
  CFA1X1 U2349 ( .A(n2152), .B(n2151), .CI(n2150), .CO(\mult_x_1/n1196 ), .S(
        \mult_x_1/n1197 ) );
  CFA1X1 U2350 ( .A(n2425), .B(n2154), .CI(n2153), .CO(n2163), .S(
        \mult_x_1/n817 ) );
  CFA1X1 U2351 ( .A(n2157), .B(n2156), .CI(n2155), .CO(n2162), .S(
        \mult_x_1/n815 ) );
  CFA1X1 U2352 ( .A(n2160), .B(n2159), .CI(n2158), .CO(n2224), .S(n2161) );
  CFA1X1 U2353 ( .A(n2163), .B(n2162), .CI(n2161), .CO(\mult_x_1/n806 ), .S(
        \mult_x_1/n807 ) );
  CFA1X1 U2354 ( .A(n2166), .B(n2165), .CI(n2164), .CO(n1605), .S(n2175) );
  CFA1X1 U2355 ( .A(n2169), .B(n2168), .CI(n2167), .CO(n2174), .S(n316) );
  CFA1X1 U2356 ( .A(n2172), .B(n2171), .CI(n2170), .CO(n1613), .S(n2173) );
  CFA1X1 U2357 ( .A(n2175), .B(n2174), .CI(n2173), .CO(\mult_x_1/n1066 ), .S(
        \mult_x_1/n1067 ) );
  CFA1X1 U2358 ( .A(n2178), .B(n2177), .CI(n2176), .CO(n1292), .S(n2187) );
  CFA1X1 U2359 ( .A(n2181), .B(n2180), .CI(n2179), .CO(n2186), .S(n1685) );
  CFA1X1 U2360 ( .A(n2183), .B(n2184), .CI(n2182), .CO(n2216), .S(n2185) );
  CFA1X1 U2361 ( .A(n2187), .B(n2186), .CI(n2185), .CO(\mult_x_1/n1284 ), .S(
        \mult_x_1/n1285 ) );
  CFA1X1 U2362 ( .A(n2190), .B(n2189), .CI(n2188), .CO(n1904), .S(n2199) );
  CFA1X1 U2363 ( .A(n2193), .B(n2192), .CI(n2191), .CO(n2198), .S(
        \mult_x_1/n1669 ) );
  CFA1X1 U2364 ( .A(n2196), .B(n2195), .CI(n2194), .CO(n1906), .S(n2197) );
  CFA1X1 U2365 ( .A(n2199), .B(n2198), .CI(n2197), .CO(\mult_x_1/n1654 ), .S(
        \mult_x_1/n1655 ) );
  CFA1X1 U2366 ( .A(n2202), .B(n2201), .CI(n2200), .CO(n2145), .S(n2211) );
  CFA1X1 U2367 ( .A(n2205), .B(n2204), .CI(n2203), .CO(n2210), .S(n498) );
  CFA1X1 U2368 ( .A(n2208), .B(n2207), .CI(n2206), .CO(n1806), .S(n2209) );
  CFA1X1 U2369 ( .A(n2211), .B(n2210), .CI(n2209), .CO(\mult_x_1/n1254 ), .S(
        \mult_x_1/n1255 ) );
  CFA1X1 U2370 ( .A(n2214), .B(n2213), .CI(n2212), .CO(n2108), .S(n2223) );
  CFA1X1 U2371 ( .A(n2217), .B(n2216), .CI(n2215), .CO(n2222), .S(n1667) );
  CFA1X1 U2372 ( .A(n2220), .B(n2219), .CI(n2218), .CO(n1808), .S(n2221) );
  CFA1X1 U2373 ( .A(n2223), .B(n2222), .CI(n2221), .CO(\mult_x_1/n1224 ), .S(
        \mult_x_1/n1225 ) );
  CFA1X1 U2374 ( .A(n2226), .B(n2225), .CI(n2224), .CO(n637), .S(
        \mult_x_1/n803 ) );
  CFA1X1 U2375 ( .A(n2229), .B(n2227), .CI(n2228), .CO(n1590), .S(n2241) );
  COND2X1 U2376 ( .A(n2233), .B(n2232), .C(n2231), .D(n2230), .Z(n2302) );
  CIVX1 U2377 ( .A(n2305), .Z(n2301) );
  COND2X1 U2378 ( .A(n256), .B(n2235), .C(n2388), .D(n2234), .Z(n2300) );
  CFA1X1 U2379 ( .A(n2238), .B(n2237), .CI(n2236), .CO(n1591), .S(n2239) );
  CFA1X1 U2380 ( .A(n2241), .B(n2240), .CI(n2239), .CO(\mult_x_1/n944 ), .S(
        \mult_x_1/n945 ) );
  CFA1X1 U2381 ( .A(n2244), .B(n2243), .CI(n2242), .CO(n1652), .S(n2253) );
  CFA1X1 U2382 ( .A(n2247), .B(n2246), .CI(n2245), .CO(n2252), .S(n1958) );
  CFA1X1 U2383 ( .A(n2250), .B(n2249), .CI(n2248), .CO(n1651), .S(n2251) );
  CFA1X1 U2384 ( .A(n2253), .B(n2252), .CI(n2251), .CO(\mult_x_1/n1314 ), .S(
        \mult_x_1/n1315 ) );
  CFA1X1 U2385 ( .A(n2256), .B(n2255), .CI(n2254), .CO(n2121), .S(n2265) );
  CFA1X1 U2386 ( .A(n2259), .B(n2258), .CI(n2257), .CO(n1257), .S(n2264) );
  CFA1X1 U2387 ( .A(n2261), .B(n2262), .CI(n2260), .CO(n2122), .S(n2263) );
  CFA1X1 U2388 ( .A(n2265), .B(n2264), .CI(n2263), .CO(\mult_x_1/n1444 ), .S(
        \mult_x_1/n1445 ) );
  CFA1X1 U2389 ( .A(n2268), .B(n2267), .CI(n2266), .CO(n1987), .S(n2277) );
  CFA1X1 U2390 ( .A(n2271), .B(n2270), .CI(n2269), .CO(n1988), .S(n2276) );
  CFA1X1 U2391 ( .A(n2274), .B(n2273), .CI(n2272), .CO(n1989), .S(n2275) );
  CFA1X1 U2392 ( .A(n2277), .B(n2276), .CI(n2275), .CO(\mult_x_1/n1022 ), .S(
        \mult_x_1/n1023 ) );
  CFA1X1 U2393 ( .A(n2280), .B(n2279), .CI(n2278), .CO(n2109), .S(n2287) );
  CFA1X1 U2394 ( .A(n2283), .B(n2282), .CI(n2281), .CO(n1809), .S(n2286) );
  CFA1X1 U2395 ( .A(n2287), .B(n2286), .CI(n2285), .CO(\mult_x_1/n1226 ), .S(
        \mult_x_1/n1227 ) );
  CFA1X1 U2396 ( .A(n2290), .B(n2289), .CI(n2288), .CO(n1870), .S(n2299) );
  CFA1X1 U2397 ( .A(n2293), .B(n2292), .CI(n2291), .CO(n1872), .S(n2298) );
  CFA1X1 U2398 ( .A(n2296), .B(n2295), .CI(n2294), .CO(n1851), .S(n2297) );
  CFA1X1 U2399 ( .A(n2299), .B(n2298), .CI(n2297), .CO(\mult_x_1/n1468 ), .S(
        \mult_x_1/n1469 ) );
  CFA1X1 U2400 ( .A(n2302), .B(n2301), .CI(n2300), .CO(n2315), .S(n2240) );
  CFA1X1 U2401 ( .A(n2305), .B(n2304), .CI(n2303), .CO(n1589), .S(n2314) );
  COND2X1 U2402 ( .A(n239), .B(n2307), .C(n2306), .D(n2510), .Z(n2376) );
  COND2X1 U2403 ( .A(n2310), .B(n2309), .C(n2430), .D(n2308), .Z(n2375) );
  COND2X1 U2404 ( .A(n261), .B(n2312), .C(n2434), .D(n2311), .Z(n2374) );
  CFA1X1 U2405 ( .A(n2315), .B(n2314), .CI(n2313), .CO(\mult_x_1/n928 ), .S(
        \mult_x_1/n929 ) );
  CFA1X1 U2406 ( .A(n2318), .B(n2317), .CI(n2316), .CO(n2097), .S(n2327) );
  CFA1X1 U2407 ( .A(n2321), .B(n2320), .CI(n2319), .CO(n1375), .S(n2326) );
  CFA1X1 U2408 ( .A(n2324), .B(n2322), .CI(n2323), .CO(n2096), .S(n2325) );
  CFA1X1 U2409 ( .A(n2327), .B(n2326), .CI(n2325), .CO(\mult_x_1/n1420 ), .S(
        \mult_x_1/n1421 ) );
  CFA1X1 U2410 ( .A(n2330), .B(n2329), .CI(n2328), .CO(n2132), .S(n2337) );
  CFA1X1 U2411 ( .A(n2334), .B(n2333), .CI(n2332), .CO(n2133), .S(n2335) );
  CFA1X1 U2412 ( .A(n2337), .B(n2336), .CI(n2335), .CO(\mult_x_1/n1666 ), .S(
        \mult_x_1/n1667 ) );
  CFA1X1 U2413 ( .A(n2340), .B(n2339), .CI(n2338), .CO(n2349), .S(n1169) );
  CFA1X1 U2414 ( .A(n2343), .B(n2342), .CI(n2341), .CO(n1731), .S(n2348) );
  CFA1X1 U2415 ( .A(n2346), .B(n2345), .CI(n2344), .CO(n1729), .S(n2347) );
  CFA1X1 U2416 ( .A(n2349), .B(n2348), .CI(n2347), .CO(\mult_x_1/n1490 ), .S(
        \mult_x_1/n1491 ) );
  CFA1X1 U2417 ( .A(n2352), .B(n2351), .CI(n2350), .CO(n2060), .S(n2361) );
  CFA1X1 U2418 ( .A(n2355), .B(n2354), .CI(n2353), .CO(n1183), .S(n2360) );
  CFA1X1 U2419 ( .A(n2358), .B(n2357), .CI(n2356), .CO(n1185), .S(n2359) );
  CFA1X1 U2420 ( .A(n2361), .B(n2360), .CI(n2359), .CO(\mult_x_1/n1002 ), .S(
        \mult_x_1/n1003 ) );
  CFA1X1 U2421 ( .A(n2364), .B(n2363), .CI(n2362), .CO(n2023), .S(n2373) );
  CFA1X1 U2422 ( .A(n2367), .B(n2366), .CI(n2365), .CO(n2019), .S(n2372) );
  CFA1X1 U2423 ( .A(n2370), .B(n2369), .CI(n2368), .CO(n2020), .S(n2371) );
  CFA1X1 U2424 ( .A(n2373), .B(n2372), .CI(n2371), .CO(\mult_x_1/n1044 ), .S(
        \mult_x_1/n1045 ) );
  CFA1X1 U2425 ( .A(n2376), .B(n2375), .CI(n2374), .CO(n2385), .S(n2313) );
  CFA1X1 U2426 ( .A(n2379), .B(n2378), .CI(n2377), .CO(n1132), .S(n2384) );
  CFA1X1 U2427 ( .A(n2382), .B(n2381), .CI(n2380), .CO(n2383), .S(n1514) );
  CFA1X1 U2428 ( .A(n2385), .B(n2384), .CI(n2383), .CO(\mult_x_1/n912 ), .S(
        \mult_x_1/n913 ) );
  CAOR1X1 U2429 ( .A(n1722), .B(n256), .C(n2386), .Z(n2417) );
  CENX1 U2430 ( .A(n2390), .B(n2389), .Z(n2399) );
  COND2X1 U2431 ( .A(n2392), .B(n2391), .C(n2398), .D(n2399), .Z(n2416) );
  CENX1 U2432 ( .A(n2470), .B(n2393), .Z(n2471) );
  COND2X1 U2433 ( .A(n263), .B(n2394), .C(n2522), .D(n2471), .Z(n2477) );
  CENX1 U2434 ( .A(n2395), .B(n2469), .Z(n2403) );
  COND2X1 U2435 ( .A(n2440), .B(n2403), .C(n292), .D(n2396), .Z(n2476) );
  COND2X1 U2436 ( .A(n2400), .B(n2399), .C(n2398), .D(n2397), .Z(n2475) );
  COND2X1 U2437 ( .A(n239), .B(n2402), .C(n2401), .D(n2510), .Z(n2421) );
  COND2X1 U2438 ( .A(n2440), .B(n2404), .C(n292), .D(n2403), .Z(n2420) );
  COND2X1 U2439 ( .A(n261), .B(n2407), .C(n243), .D(n2405), .Z(n2419) );
  CFA1X1 U2440 ( .A(n2410), .B(n2409), .CI(n2408), .CO(\mult_x_1/n858 ), .S(
        \mult_x_1/n859 ) );
  CFA1X1 U2441 ( .A(n2415), .B(n2414), .CI(n2413), .CO(n2424), .S(n1272) );
  CFA1X1 U2442 ( .A(n2418), .B(n2417), .CI(n2416), .CO(n2410), .S(n2423) );
  CFA1X1 U2443 ( .A(n2421), .B(n2420), .CI(n2419), .CO(n2408), .S(n2422) );
  CFA1X1 U2444 ( .A(n2424), .B(n2423), .CI(n2422), .CO(\mult_x_1/n870 ), .S(
        \mult_x_1/n871 ) );
  CIVX1 U2445 ( .A(n2425), .Z(n2445) );
  CENX1 U2446 ( .A(n2427), .B(n2426), .Z(n2437) );
  COND2X1 U2447 ( .A(n239), .B(n2437), .C(n2428), .D(n2510), .Z(n2453) );
  COND2X1 U2448 ( .A(n2432), .B(n2431), .C(n2430), .D(n2429), .Z(n2452) );
  COND2X1 U2449 ( .A(n261), .B(n2435), .C(n2434), .D(n2433), .Z(n2451) );
  COND2X1 U2450 ( .A(n239), .B(n2438), .C(n2437), .D(n2510), .Z(n2528) );
  CAOR1X1 U2451 ( .A(n292), .B(n2440), .C(n2439), .Z(n2450) );
  CENX1 U2452 ( .A(n2470), .B(n2441), .Z(n2521) );
  COND2X1 U2453 ( .A(n263), .B(n2521), .C(n2522), .D(n2442), .Z(n2449) );
  CFA1X1 U2454 ( .A(n2445), .B(n2444), .CI(n2443), .CO(\mult_x_1/n820 ), .S(
        \mult_x_1/n821 ) );
  CFA1X1 U2455 ( .A(n2448), .B(n2447), .CI(n2446), .CO(n2456), .S(
        \mult_x_1/n841 ) );
  CFA1X1 U2456 ( .A(n2528), .B(n2450), .CI(n2449), .CO(n2443), .S(n2455) );
  CFA1X1 U2457 ( .A(n2453), .B(n2452), .CI(n2451), .CO(n2444), .S(n2454) );
  CFA1X1 U2458 ( .A(n2456), .B(n2455), .CI(n2454), .CO(\mult_x_1/n828 ), .S(
        \mult_x_1/n829 ) );
  COND1XL U2459 ( .A(n2458), .B(n2463), .C(n2457), .Z(n2461) );
  CND2X1 U2460 ( .A(n272), .B(n2459), .Z(n2460) );
  CENX1 U2461 ( .A(n2461), .B(n2460), .Z(n2900) );
  CENX1 U2462 ( .A(n2470), .B(n2469), .Z(n2523) );
  COND2X1 U2463 ( .A(n263), .B(n2471), .C(n2522), .D(n2523), .Z(n2480) );
  CFA1X1 U2464 ( .A(n2474), .B(n2473), .CI(n2472), .CO(n2479), .S(
        \mult_x_1/n861 ) );
  CFA1X1 U2465 ( .A(n2477), .B(n2476), .CI(n2475), .CO(n2478), .S(n2409) );
  CFA1X1 U2466 ( .A(n2480), .B(n2479), .CI(n2478), .CO(\mult_x_1/n848 ), .S(
        \mult_x_1/n849 ) );
  CND2X1 U2467 ( .A(n2484), .B(n2483), .Z(\mult_x_1/n178 ) );
  CND2X1 U2468 ( .A(n2486), .B(n2485), .Z(\mult_x_1/n176 ) );
  CFA1X1 U2469 ( .A(n2499), .B(n2498), .CI(n2497), .CO(\mult_x_1/n796 ), .S(
        n625) );
  CND2X1 U2470 ( .A(n2501), .B(n2500), .Z(n2503) );
  CENX1 U2471 ( .A(n2503), .B(n2502), .Z(n2916) );
  CND2XL U2472 ( .A(n2505), .B(n2504), .Z(n2506) );
  CENX1 U2473 ( .A(n2507), .B(n2506), .Z(n2908) );
  CAOR1X1 U2474 ( .A(n2510), .B(n239), .C(n2508), .Z(\mult_x_1/n1740 ) );
  CIVX1 U2475 ( .A(n2513), .Z(n2514) );
  CND2XL U2476 ( .A(n2516), .B(n2515), .Z(n2520) );
  CANR1XL U2477 ( .A(n2518), .B(n2548), .C(n2517), .Z(n2519) );
  CEOXL U2478 ( .A(n2520), .B(n2519), .Z(n2896) );
  COND2X1 U2479 ( .A(n263), .B(n2523), .C(n2522), .D(n2521), .Z(n2531) );
  CFA1X1 U2480 ( .A(n2527), .B(n2526), .CI(n2525), .CO(n2530), .S(
        \mult_x_1/n853 ) );
  CIVX1 U2481 ( .A(n2528), .Z(n2529) );
  CFA1X1 U2482 ( .A(n2531), .B(n2530), .CI(n2529), .CO(\mult_x_1/n838 ), .S(
        \mult_x_1/n839 ) );
  CND2XL U2483 ( .A(n31), .B(n2571), .Z(\mult_x_1/n153 ) );
  CEOXL U2484 ( .A(n2536), .B(n2535), .Z(n2912) );
  CND2X1 U2485 ( .A(n2538), .B(n2537), .Z(n2539) );
  CEOXL U2486 ( .A(n2539), .B(n2542), .Z(n2895) );
  CIVXL U2487 ( .A(n2540), .Z(n2541) );
endmodule


module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push_2, push_0, push_1, n498, n499, n500, n502, n503, n504, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n572, n574, n576, n577, n578, n579, n580,
         n582, n584, n586, n588, n596, n599, n602, n603, n604, n605, n606,
         n607, n608, n634, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] mulout;
  wire   [63:0] acc;
  wire   [1:0] cmd_2;
  wire   [6:0] h2;
  wire   [1:0] cmd0;
  wire   [6:0] h1;
  wire   [1:0] cmd_1;

  CFD2QX1 \h0_reg[31]  ( .D(n774), .CP(clk), .CD(n3633), .Q(h0[31]) );
  CFD2QX1 \h0_reg[30]  ( .D(n773), .CP(clk), .CD(n3629), .Q(h0[30]) );
  CFD2QX1 \h0_reg[29]  ( .D(n772), .CP(clk), .CD(n3629), .Q(h0[29]) );
  CFD2QX1 \h0_reg[28]  ( .D(n771), .CP(clk), .CD(n3629), .Q(h0[28]) );
  CFD2QX1 \h0_reg[27]  ( .D(n770), .CP(clk), .CD(n3629), .Q(h0[27]) );
  CFD2QX1 \h0_reg[26]  ( .D(n769), .CP(clk), .CD(n3629), .Q(h0[26]) );
  CFD2QX1 \h0_reg[25]  ( .D(n768), .CP(clk), .CD(n3633), .Q(h0[25]) );
  CFD2QX1 \h0_reg[24]  ( .D(n767), .CP(clk), .CD(n3629), .Q(h0[24]) );
  CFD2QX1 \h0_reg[23]  ( .D(n765), .CP(clk), .CD(n3633), .Q(h0[23]) );
  CFD2QX1 \h0_reg[22]  ( .D(n763), .CP(clk), .CD(n3629), .Q(h0[22]) );
  CFD2QX1 \h0_reg[21]  ( .D(n761), .CP(clk), .CD(n3633), .Q(h0[21]) );
  CFD2QX1 \h0_reg[20]  ( .D(n759), .CP(clk), .CD(n3629), .Q(h0[20]) );
  CFD2QX1 \h0_reg[19]  ( .D(n757), .CP(clk), .CD(n3633), .Q(h0[19]) );
  CFD2QX1 \h0_reg[18]  ( .D(n755), .CP(clk), .CD(n3629), .Q(h0[18]) );
  CFD2QX1 \h0_reg[17]  ( .D(n753), .CP(clk), .CD(n3633), .Q(h0[17]) );
  CFD2QX1 \h0_reg[16]  ( .D(n751), .CP(clk), .CD(n3629), .Q(h0[16]) );
  CFD2QX1 \h0_reg[15]  ( .D(n749), .CP(clk), .CD(n3633), .Q(h0[15]) );
  CFD2QX1 \h0_reg[14]  ( .D(n747), .CP(clk), .CD(n3629), .Q(h0[14]) );
  CFD2QX1 \h0_reg[13]  ( .D(n745), .CP(clk), .CD(n3629), .Q(h0[13]) );
  CFD2QX1 \h0_reg[12]  ( .D(n743), .CP(clk), .CD(n3629), .Q(h0[12]) );
  CFD2QX1 \h0_reg[11]  ( .D(n741), .CP(clk), .CD(n3633), .Q(h0[11]) );
  CFD2QX1 \h0_reg[10]  ( .D(n739), .CP(clk), .CD(n3629), .Q(h0[10]) );
  CFD2QX1 \h0_reg[9]  ( .D(n737), .CP(clk), .CD(n3629), .Q(h0[9]) );
  CFD2QX1 \h0_reg[8]  ( .D(n735), .CP(clk), .CD(n3633), .Q(h0[8]) );
  CFD2QX1 \h0_reg[7]  ( .D(n733), .CP(clk), .CD(n3633), .Q(h0[7]) );
  CFD2QX1 \h0_reg[6]  ( .D(n608), .CP(clk), .CD(n3629), .Q(h0[6]) );
  CFD2QX1 \h0_reg[5]  ( .D(n607), .CP(clk), .CD(n3633), .Q(h0[5]) );
  CFD2QX1 \h0_reg[4]  ( .D(n606), .CP(clk), .CD(n3629), .Q(h0[4]) );
  CFD2QX1 \h0_reg[3]  ( .D(n605), .CP(clk), .CD(n3633), .Q(h0[3]) );
  CFD2QX1 \h0_reg[2]  ( .D(n604), .CP(clk), .CD(n3633), .Q(h0[2]) );
  CFD2QX1 \h0_reg[1]  ( .D(n603), .CP(clk), .CD(n3633), .Q(h0[1]) );
  CFD2QX1 \h0_reg[0]  ( .D(n602), .CP(clk), .CD(n3629), .Q(h0[0]) );
  CFD2QX1 \q0_reg[30]  ( .D(n731), .CP(clk), .CD(n3629), .Q(q0[30]) );
  CFD2QX1 \q0_reg[24]  ( .D(n729), .CP(clk), .CD(n3629), .Q(q0[24]) );
  CFD2QX1 \q0_reg[22]  ( .D(n727), .CP(clk), .CD(n3629), .Q(q0[22]) );
  CFD2QX1 \q0_reg[21]  ( .D(n726), .CP(clk), .CD(n3629), .Q(q0[21]) );
  CFD2QX1 \q0_reg[20]  ( .D(n725), .CP(clk), .CD(n3629), .Q(q0[20]) );
  CFD2QX1 \q0_reg[17]  ( .D(n724), .CP(clk), .CD(n3629), .Q(q0[17]) );
  CFD2QX1 \q0_reg[12]  ( .D(n582), .CP(clk), .CD(n3633), .Q(q0[12]) );
  CFD2QX1 \q0_reg[11]  ( .D(n723), .CP(clk), .CD(n3629), .Q(q0[11]) );
  CFD2QX1 \q0_reg[9]  ( .D(n579), .CP(clk), .CD(n3629), .Q(q0[9]) );
  CFD2QX1 \q0_reg[7]  ( .D(n577), .CP(clk), .CD(n3629), .Q(q0[7]) );
  CFD2QX1 \q0_reg[3]  ( .D(n1708), .CP(clk), .CD(n3633), .Q(q0[3]) );
  CFD2QX1 \q0_reg[2]  ( .D(n572), .CP(clk), .CD(n3629), .Q(q0[2]) );
  CFD2QX1 \acc_reg[3]  ( .D(n1706), .CP(clk), .CD(n3629), .Q(acc[3]) );
  CFD2QX1 \acc_reg[4]  ( .D(n565), .CP(clk), .CD(n3629), .Q(acc[4]) );
  CFD2QX1 \acc_reg[5]  ( .D(n564), .CP(clk), .CD(n3633), .Q(acc[5]) );
  CFD2QX1 \acc_reg[6]  ( .D(n563), .CP(clk), .CD(n3633), .Q(acc[6]) );
  CFD2QX1 \acc_reg[7]  ( .D(n562), .CP(clk), .CD(n3629), .Q(acc[7]) );
  CFD2QX1 \acc_reg[9]  ( .D(n560), .CP(clk), .CD(n3629), .Q(acc[9]) );
  CFD2QX1 \acc_reg[12]  ( .D(n557), .CP(clk), .CD(n3629), .Q(acc[12]) );
  CFD2QX1 \acc_reg[13]  ( .D(n556), .CP(clk), .CD(n3629), .Q(acc[13]) );
  CFD2QX1 \acc_reg[14]  ( .D(n555), .CP(clk), .CD(n3629), .Q(acc[14]) );
  CFD2QX1 \acc_reg[15]  ( .D(n554), .CP(clk), .CD(n3629), .Q(acc[15]) );
  CFD2QX1 \acc_reg[21]  ( .D(n548), .CP(clk), .CD(n3633), .Q(acc[21]) );
  CFD2QX1 \acc_reg[22]  ( .D(n547), .CP(clk), .CD(n3629), .Q(acc[22]) );
  CFD2QX1 \acc_reg[23]  ( .D(n546), .CP(clk), .CD(n3629), .Q(acc[23]) );
  CFD2QX1 \acc_reg[24]  ( .D(n545), .CP(clk), .CD(n3629), .Q(acc[24]) );
  CFD2QX1 \acc_reg[25]  ( .D(n544), .CP(clk), .CD(n3633), .Q(acc[25]) );
  CFD2QX1 \acc_reg[27]  ( .D(n542), .CP(clk), .CD(n3633), .Q(acc[27]) );
  CFD2QX1 \acc_reg[28]  ( .D(n541), .CP(clk), .CD(n3629), .Q(acc[28]) );
  sfilt_DW02_mult_3_stage_J1_0 pipe ( .A(q0), .B(h0), .TC(1'b1), .CLK(clk), 
        .PRODUCT(mulout) );
  CFD1QX4 \h2_reg[5]  ( .D(n779), .CP(clk), .Q(h2[5]) );
  CFD1QX4 \h2_reg[3]  ( .D(n720), .CP(clk), .Q(h2[3]) );
  CFD1QX4 \h2_reg[4]  ( .D(n502), .CP(clk), .Q(h2[4]) );
  CFD2QX2 \q0_reg[29]  ( .D(n599), .CP(clk), .CD(n3629), .Q(q0[29]) );
  CFD2QX2 \q0_reg[23]  ( .D(n730), .CP(clk), .CD(n3629), .Q(q0[23]) );
  CFD2QX2 \q0_reg[31]  ( .D(n728), .CP(clk), .CD(n3629), .Q(q0[31]) );
  CFD2QX2 \q0_reg[27]  ( .D(n732), .CP(clk), .CD(n3629), .Q(q0[27]) );
  CFD2QX4 \q0_reg[10]  ( .D(n580), .CP(clk), .CD(n3629), .Q(q0[10]) );
  CFD2QX4 \q0_reg[18]  ( .D(n588), .CP(clk), .CD(n3629), .Q(q0[18]) );
  CFD2QX4 \q0_reg[4]  ( .D(n574), .CP(clk), .CD(n3629), .Q(q0[4]) );
  CFD1QX4 \h2_reg[0]  ( .D(n498), .CP(clk), .Q(h2[0]) );
  CFD1QX4 \h2_reg[1]  ( .D(n499), .CP(clk), .Q(h2[1]) );
  CFD2QX2 \acc_reg[53]  ( .D(n516), .CP(clk), .CD(n3629), .Q(acc[53]) );
  CFD2QX2 \acc_reg[52]  ( .D(n517), .CP(clk), .CD(n3629), .Q(acc[52]) );
  CFD2QX2 \acc_reg[33]  ( .D(n536), .CP(clk), .CD(n3633), .Q(acc[33]) );
  CFD2QX2 \acc_reg[51]  ( .D(n518), .CP(clk), .CD(n3629), .Q(acc[51]) );
  CFD2QX2 \acc_reg[41]  ( .D(n528), .CP(clk), .CD(n3629), .Q(acc[41]) );
  CFD2QX2 \q0_reg[15]  ( .D(n849), .CP(clk), .CD(n3629), .Q(q0[15]) );
  CFD2QX2 \q0_reg[13]  ( .D(n847), .CP(clk), .CD(n3629), .Q(q0[13]) );
  CFD2QX2 \q0_reg[19]  ( .D(n848), .CP(clk), .CD(n3629), .Q(q0[19]) );
  CFD2QX2 \acc_reg[58]  ( .D(n511), .CP(clk), .CD(n3633), .Q(acc[58]) );
  CFD2QX2 \acc_reg[20]  ( .D(n549), .CP(clk), .CD(n3629), .Q(acc[20]) );
  CFD2QX2 \acc_reg[46]  ( .D(n523), .CP(clk), .CD(n3629), .Q(acc[46]) );
  CFD2QX2 \acc_reg[47]  ( .D(n522), .CP(clk), .CD(n3629), .Q(acc[47]) );
  CFD2QX2 \q0_reg[8]  ( .D(n578), .CP(clk), .CD(n3629), .Q(q0[8]) );
  CFD2QX2 \acc_reg[43]  ( .D(n526), .CP(clk), .CD(n3629), .Q(acc[43]) );
  CFD2QX2 \acc_reg[36]  ( .D(n533), .CP(clk), .CD(n3629), .Q(acc[36]) );
  CFD2QX2 \acc_reg[57]  ( .D(n512), .CP(clk), .CD(n3629), .Q(acc[57]) );
  CFD2QX2 \acc_reg[48]  ( .D(n521), .CP(clk), .CD(n3629), .Q(acc[48]) );
  CFD2QX2 \acc_reg[38]  ( .D(n531), .CP(clk), .CD(n3629), .Q(acc[38]) );
  CFD2QX2 \acc_reg[55]  ( .D(n514), .CP(clk), .CD(n3629), .Q(acc[55]) );
  CFD2QX4 \q0_reg[6]  ( .D(n576), .CP(clk), .CD(n3629), .Q(q0[6]) );
  CFD2QX2 \acc_reg[30]  ( .D(n539), .CP(clk), .CD(n3629), .Q(acc[30]) );
  CFD2QX2 \acc_reg[11]  ( .D(n558), .CP(clk), .CD(n3629), .Q(acc[11]) );
  CFD2QX2 \acc_reg[8]  ( .D(n561), .CP(clk), .CD(n3629), .Q(acc[8]) );
  CFD2QX2 \acc_reg[10]  ( .D(n559), .CP(clk), .CD(n3629), .Q(acc[10]) );
  CFD2X2 \acc_reg[62]  ( .D(n507), .CP(clk), .CD(n3629), .Q(acc[62]), .QN(
        n3630) );
  CFD2QX2 \q0_reg[28]  ( .D(n843), .CP(clk), .CD(n3629), .Q(q0[28]) );
  CFD2QX2 \acc_reg[17]  ( .D(n552), .CP(clk), .CD(n3629), .Q(acc[17]) );
  CFD2X1 \acc_reg[44]  ( .D(n525), .CP(clk), .CD(n3629), .Q(acc[44]), .QN(
        n3632) );
  CFD2QXL \h1_reg[6]  ( .D(n840), .CP(clk), .CD(n3629), .Q(h1[6]) );
  CFD2QXL \h1_reg[5]  ( .D(n827), .CP(clk), .CD(n3629), .Q(h1[5]) );
  CFD2QXL push_2_reg ( .D(n830), .CP(clk), .CD(n3629), .Q(push_2) );
  CFD2QXL \cmd_2_reg[1]  ( .D(n832), .CP(clk), .CD(n3629), .Q(cmd_2[1]) );
  CFD2QXL \h1_reg[4]  ( .D(n834), .CP(clk), .CD(n3629), .Q(h1[4]) );
  CFD2QXL \h1_reg[3]  ( .D(n837), .CP(clk), .CD(n3629), .Q(h1[3]) );
  CFD2QXL \h1_reg[2]  ( .D(n815), .CP(clk), .CD(n3629), .Q(h1[2]) );
  CFD2QXL \h1_reg[1]  ( .D(n818), .CP(clk), .CD(n3629), .Q(h1[1]) );
  CFD2QXL push_1_reg ( .D(n821), .CP(clk), .CD(n3629), .Q(push_1) );
  CFD2QXL \cmd_2_reg[0]  ( .D(n823), .CP(clk), .CD(n3629), .Q(cmd_2[0]) );
  CFD2QXL \cmd_1_reg[1]  ( .D(n825), .CP(clk), .CD(n3629), .Q(cmd_1[1]) );
  CFD2QXL \cmd_1_reg[0]  ( .D(n810), .CP(clk), .CD(n3629), .Q(cmd_1[0]) );
  CFD2QXL \h1_reg[0]  ( .D(n812), .CP(clk), .CD(n3629), .Q(h1[0]) );
  CFD2QXL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n3629), .Q(cmd0[1]) );
  CFD2QXL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n3629), .Q(cmd0[0]) );
  CFD2QXL _pushout_reg ( .D(n3628), .CP(clk), .CD(n3629), .Q(pushout) );
  CFD2QXL push_0_reg ( .D(pushin), .CP(clk), .CD(n3629), .Q(push_0) );
  CFD2QXL \dout_reg[31]  ( .D(n807), .CP(clk), .CD(n3629), .Q(z[31]) );
  CFD2QXL \dout_reg[30]  ( .D(n808), .CP(clk), .CD(n3629), .Q(z[30]) );
  CFD2QXL \dout_reg[29]  ( .D(n637), .CP(clk), .CD(n3629), .Q(z[29]) );
  CFD2QXL \dout_reg[28]  ( .D(n809), .CP(clk), .CD(n3629), .Q(z[28]) );
  CFD2QXL \dout_reg[1]  ( .D(n802), .CP(clk), .CD(n3629), .Q(z[1]) );
  CFD2QXL \dout_reg[0]  ( .D(n666), .CP(clk), .CD(n3629), .Q(z[0]) );
  CFD2QXL \dout_reg[27]  ( .D(n804), .CP(clk), .CD(n3629), .Q(z[27]) );
  CFD2QXL \dout_reg[26]  ( .D(n805), .CP(clk), .CD(n3629), .Q(z[26]) );
  CFD2QXL \dout_reg[25]  ( .D(n806), .CP(clk), .CD(n3629), .Q(z[25]) );
  CFD2QXL \dout_reg[24]  ( .D(n797), .CP(clk), .CD(n3629), .Q(z[24]) );
  CFD2QXL \dout_reg[23]  ( .D(n798), .CP(clk), .CD(n3629), .Q(z[23]) );
  CFD2QXL \dout_reg[22]  ( .D(n799), .CP(clk), .CD(n3629), .Q(z[22]) );
  CFD2QXL \dout_reg[21]  ( .D(n800), .CP(clk), .CD(n3629), .Q(z[21]) );
  CFD2QXL \dout_reg[20]  ( .D(n801), .CP(clk), .CD(n3629), .Q(z[20]) );
  CFD2QXL \dout_reg[19]  ( .D(n793), .CP(clk), .CD(n3629), .Q(z[19]) );
  CFD2QXL \dout_reg[18]  ( .D(n715), .CP(clk), .CD(n3629), .Q(z[18]) );
  CFD2QXL \dout_reg[17]  ( .D(n794), .CP(clk), .CD(n3629), .Q(z[17]) );
  CFD2QXL \dout_reg[16]  ( .D(n795), .CP(clk), .CD(n3629), .Q(z[16]) );
  CFD2QXL \dout_reg[15]  ( .D(n796), .CP(clk), .CD(n3629), .Q(z[15]) );
  CFD2QXL \dout_reg[14]  ( .D(n789), .CP(clk), .CD(n3629), .Q(z[14]) );
  CFD2QXL \dout_reg[13]  ( .D(n716), .CP(clk), .CD(n3629), .Q(z[13]) );
  CFD2QXL \dout_reg[12]  ( .D(n790), .CP(clk), .CD(n3629), .Q(z[12]) );
  CFD2QXL \dout_reg[11]  ( .D(n791), .CP(clk), .CD(n3629), .Q(z[11]) );
  CFD2QXL \dout_reg[10]  ( .D(n792), .CP(clk), .CD(n3629), .Q(z[10]) );
  CFD2QXL \dout_reg[9]  ( .D(n785), .CP(clk), .CD(n3629), .Q(z[9]) );
  CFD2QXL \dout_reg[8]  ( .D(n717), .CP(clk), .CD(n3629), .Q(z[8]) );
  CFD2QXL \dout_reg[7]  ( .D(n786), .CP(clk), .CD(n3629), .Q(z[7]) );
  CFD2QXL \dout_reg[6]  ( .D(n787), .CP(clk), .CD(n3629), .Q(z[6]) );
  CFD2QXL \dout_reg[5]  ( .D(n788), .CP(clk), .CD(n3629), .Q(z[5]) );
  CFD2QXL \dout_reg[4]  ( .D(n783), .CP(clk), .CD(n3629), .Q(z[4]) );
  CFD2QXL \dout_reg[3]  ( .D(n718), .CP(clk), .CD(n3629), .Q(z[3]) );
  CFD2QXL \dout_reg[2]  ( .D(n784), .CP(clk), .CD(n3629), .Q(z[2]) );
  CFD4X2 \acc_reg[0]  ( .D(n782), .CP(clk), .SD(n3629), .QN(acc[0]) );
  CFD4X2 \acc_reg[2]  ( .D(n781), .CP(clk), .SD(n3629), .QN(acc[2]) );
  CFD1QX4 \h2_reg[6]  ( .D(n780), .CP(clk), .Q(h2[6]) );
  CFD2X1 \acc_reg[63]  ( .D(n506), .CP(clk), .CD(n3629), .Q(acc[63]), .QN(
        n3631) );
  CFD1QX4 \h2_reg[2]  ( .D(n778), .CP(clk), .Q(h2[2]) );
  CFD2QX2 \q0_reg[16]  ( .D(n586), .CP(clk), .CD(n3629), .Q(q0[16]) );
  CFD2X2 \acc_reg[60]  ( .D(n509), .CP(clk), .CD(n3629), .Q(n1180), .QN(n1181)
         );
  CFD2QX2 \q0_reg[1]  ( .D(n777), .CP(clk), .CD(n3629), .Q(q0[1]) );
  CFD2XL \acc_reg[40]  ( .D(n529), .CP(clk), .CD(n3629), .Q(n1166), .QN(n1167)
         );
  CFD2X2 \acc_reg[56]  ( .D(n513), .CP(clk), .CD(n3633), .Q(n1108), .QN(n1109)
         );
  CFD2QX2 \q0_reg[5]  ( .D(n776), .CP(clk), .CD(n3633), .Q(q0[5]) );
  CFD2X1 \acc_reg[49]  ( .D(n520), .CP(clk), .CD(n3629), .Q(n1162), .QN(n1163)
         );
  CFD2XL \acc_reg[50]  ( .D(n519), .CP(clk), .CD(n3633), .Q(n1126), .QN(n1125)
         );
  CFD2X2 \acc_reg[54]  ( .D(n515), .CP(clk), .CD(n3629), .Q(n1088), .QN(n1089)
         );
  CFD2QX4 \acc_reg[31]  ( .D(n538), .CP(clk), .CD(n3629), .Q(acc[31]) );
  CFD2QX2 \q0_reg[26]  ( .D(n596), .CP(clk), .CD(n3629), .Q(q0[26]) );
  CFD2X2 \acc_reg[61]  ( .D(n508), .CP(clk), .CD(n3629), .Q(n1080), .QN(n1081)
         );
  CFD2QX2 \q0_reg[25]  ( .D(n1717), .CP(clk), .CD(n3629), .Q(q0[25]) );
  CFD2X2 \acc_reg[42]  ( .D(n527), .CP(clk), .CD(n3629), .Q(n1072), .QN(n1073)
         );
  CFD2X4 \acc_reg[59]  ( .D(n510), .CP(clk), .CD(n3629), .Q(n1065), .QN(n1066)
         );
  CFD2QX1 \acc_reg[35]  ( .D(n534), .CP(clk), .CD(n3629), .Q(acc[35]) );
  CFD2QX1 \q0_reg[0]  ( .D(n775), .CP(clk), .CD(n3629), .Q(q0[0]) );
  CFD4X1 \acc_reg[1]  ( .D(n719), .CP(clk), .SD(n3629), .QN(acc[1]) );
  CFD2X1 \acc_reg[29]  ( .D(n540), .CP(clk), .CD(n3629), .Q(n1139), .QN(n1138)
         );
  CFD2X2 \acc_reg[45]  ( .D(n524), .CP(clk), .CD(n3633), .Q(n858) );
  CFD2QX4 \acc_reg[34]  ( .D(n535), .CP(clk), .CD(n3633), .Q(acc[34]) );
  CFD2QX2 \acc_reg[26]  ( .D(n543), .CP(clk), .CD(n3633), .Q(acc[26]) );
  CFD2QX2 \acc_reg[16]  ( .D(n553), .CP(clk), .CD(n3633), .Q(acc[16]) );
  CFD2QX4 \acc_reg[19]  ( .D(n550), .CP(clk), .CD(n3629), .Q(acc[19]) );
  CFD2QX2 \acc_reg[18]  ( .D(n551), .CP(clk), .CD(n3629), .Q(acc[18]) );
  CFD2QX2 \q0_reg[14]  ( .D(n584), .CP(clk), .CD(n3629), .Q(q0[14]) );
  CFD2QX2 \acc_reg[37]  ( .D(n532), .CP(clk), .CD(n3629), .Q(acc[37]) );
  CFD2QX2 \acc_reg[39]  ( .D(n530), .CP(clk), .CD(n3629), .Q(acc[39]) );
  CFD2QX2 \acc_reg[32]  ( .D(n537), .CP(clk), .CD(n3629), .Q(acc[32]) );
  CIVXL U737 ( .A(n669), .Z(n1201) );
  CND3XL U738 ( .A(n2686), .B(n3513), .C(n1141), .Z(n669) );
  CNR2XL U739 ( .A(n3319), .B(n3318), .Z(n3324) );
  CND2XL U740 ( .A(n3324), .B(n3323), .Z(n520) );
  CNR2X2 U741 ( .A(n1617), .B(n1242), .Z(n1244) );
  CIVX3 U742 ( .A(n1558), .Z(n1648) );
  CIVX3 U743 ( .A(n3025), .Z(n3255) );
  CANR2X1 U744 ( .A(n2058), .B(n2007), .C(n2151), .D(n2052), .Z(n2008) );
  CND3X2 U745 ( .A(n2010), .B(n2009), .C(n2008), .Z(n2022) );
  CND2IX1 U746 ( .B(n2978), .A(n2979), .Z(n2996) );
  CND2IXL U747 ( .B(n2996), .A(n3269), .Z(n2982) );
  CND2IXL U748 ( .B(n670), .A(n2680), .Z(n2682) );
  CIVXL U749 ( .A(n3162), .Z(n670) );
  COND1X1 U750 ( .A(n3605), .B(n672), .C(n671), .Z(n3550) );
  CIVX2 U751 ( .A(n3527), .Z(n671) );
  CIVX2 U752 ( .A(n3608), .Z(n672) );
  CND2X1 U753 ( .A(n1517), .B(acc[16]), .Z(n1373) );
  CND2IX2 U754 ( .B(n2155), .A(n2052), .Z(n1792) );
  CND2X1 U755 ( .A(n1981), .B(n2373), .Z(n1827) );
  CAN3X2 U756 ( .A(n1850), .B(n1848), .C(n1849), .Z(n2660) );
  CND2X2 U757 ( .A(n673), .B(n2060), .Z(n2062) );
  CIVX2 U758 ( .A(n2061), .Z(n673) );
  CND3X1 U759 ( .A(n3039), .B(n3038), .C(n674), .Z(n509) );
  CANR1X2 U760 ( .A(n3029), .B(n3168), .C(n3028), .Z(n674) );
  CNR2X2 U761 ( .A(n1446), .B(n1080), .Z(n1023) );
  CND2IX2 U762 ( .B(n2768), .A(n2774), .Z(n2773) );
  CND2X2 U763 ( .A(n2015), .B(n2368), .Z(n1788) );
  CANR1X2 U764 ( .A(n676), .B(n675), .C(n2577), .Z(n2578) );
  CIVX2 U765 ( .A(n2774), .Z(n675) );
  CIVX2 U766 ( .A(n1031), .Z(n676) );
  COND1X2 U767 ( .A(n3325), .B(n679), .C(n677), .Z(n561) );
  CNR2IX2 U768 ( .B(n3378), .A(n678), .Z(n677) );
  CIVX2 U769 ( .A(n845), .Z(n678) );
  CENX2 U770 ( .A(n3373), .B(n3372), .Z(n679) );
  CND3X2 U771 ( .A(n3255), .B(n692), .C(n691), .Z(n3168) );
  COND1X1 U772 ( .A(n680), .B(n688), .C(n2268), .Z(n2188) );
  CND2X1 U773 ( .A(n1790), .B(n1791), .Z(n680) );
  CND2X2 U774 ( .A(n1508), .B(n1089), .Z(n1359) );
  CIVX2 U775 ( .A(n2629), .Z(n1083) );
  CANR2X1 U776 ( .A(n2707), .B(n2014), .C(n2137), .D(n1831), .Z(n2321) );
  CNR2X1 U777 ( .A(n1756), .B(n1755), .Z(n2707) );
  CND4X2 U778 ( .A(n1449), .B(n1450), .C(n1448), .D(n681), .Z(n2100) );
  CND2IX1 U779 ( .B(n1447), .A(n682), .Z(n681) );
  CIVX2 U780 ( .A(n1633), .Z(n682) );
  CNR2XL U781 ( .A(n684), .B(n683), .Z(n1406) );
  CIVXL U782 ( .A(n1390), .Z(n683) );
  CND2XL U783 ( .A(n685), .B(n2121), .Z(n684) );
  CND2IXL U784 ( .B(n686), .A(n1681), .Z(n685) );
  CIVX3 U785 ( .A(n1922), .Z(n686) );
  CNIVX3 U786 ( .A(n2820), .Z(n1186) );
  CND2IXL U787 ( .B(n687), .A(n2422), .Z(n2356) );
  CIVX2 U788 ( .A(n2344), .Z(n687) );
  CNR2X2 U789 ( .A(n1806), .B(n1805), .Z(n2190) );
  CANR1X2 U790 ( .A(n2349), .B(n2190), .C(n2507), .Z(n3127) );
  CND2X1 U791 ( .A(n1789), .B(n1788), .Z(n688) );
  CND2IX1 U792 ( .B(n3143), .A(n689), .Z(n543) );
  CANR1X2 U793 ( .A(n3144), .B(n3229), .C(n690), .Z(n689) );
  CIVX2 U794 ( .A(n3153), .Z(n690) );
  CND2IX1 U795 ( .B(n1625), .A(acc[38]), .Z(n1417) );
  CND3X2 U796 ( .A(n1417), .B(n1416), .C(n1415), .Z(n2103) );
  CNR2X1 U797 ( .A(n3022), .B(n3023), .Z(n691) );
  CIVXL U798 ( .A(n3024), .Z(n692) );
  CND2XL U799 ( .A(n694), .B(n693), .Z(n2633) );
  COND11X1 U800 ( .A(n1210), .B(n3015), .C(n1105), .D(n2632), .Z(n693) );
  CND3X1 U801 ( .A(n2630), .B(n2629), .C(n695), .Z(n694) );
  CIVX3 U802 ( .A(n2766), .Z(n695) );
  CND2X2 U803 ( .A(n2589), .B(n1199), .Z(n698) );
  CND2XL U804 ( .A(n696), .B(n953), .Z(n2595) );
  CND3X1 U805 ( .A(n2589), .B(n1199), .C(n697), .Z(n696) );
  CIVXL U806 ( .A(n952), .Z(n697) );
  CIVX2 U807 ( .A(n698), .Z(n3519) );
  CND2X2 U808 ( .A(n698), .B(n3511), .Z(n3040) );
  CIVX2 U809 ( .A(n2508), .Z(n2448) );
  CND2X2 U810 ( .A(n701), .B(n699), .Z(n2508) );
  CNR2IX2 U811 ( .B(n2087), .A(n700), .Z(n699) );
  CNR2XL U812 ( .A(n2088), .B(n2089), .Z(n700) );
  CIVX2 U813 ( .A(n2092), .Z(n701) );
  CND2X2 U814 ( .A(n2448), .B(n2435), .Z(n2390) );
  COND1X1 U815 ( .A(n2761), .B(n2762), .C(n2760), .Z(n511) );
  CNR2X2 U816 ( .A(n2744), .B(n1193), .Z(n2762) );
  CANR1X1 U817 ( .A(n3595), .B(n966), .C(n965), .Z(n3627) );
  CND2XL U818 ( .A(n2904), .B(n702), .Z(n528) );
  CANR1XL U819 ( .A(n2902), .B(n1105), .C(n2898), .Z(n702) );
  CNR2XL U820 ( .A(n3555), .B(n1204), .Z(n2499) );
  CDLY1XL U821 ( .A(q0[13]), .Z(n708) );
  COND1XL U822 ( .A(n1953), .B(n1952), .C(h2[5]), .Z(n703) );
  CNR2X2 U823 ( .A(n1949), .B(n1948), .Z(n2852) );
  COR2XL U824 ( .A(n1204), .B(n3551), .Z(n2501) );
  COR2XL U825 ( .A(n3335), .B(n3551), .Z(n3336) );
  CNR2X1 U826 ( .A(n3390), .B(n3389), .Z(n3391) );
  CND2XL U827 ( .A(n3391), .B(n3392), .Z(n555) );
  CND2XL U828 ( .A(n3443), .B(n3464), .Z(n1144) );
  COND1X1 U829 ( .A(n3325), .B(n3499), .C(n3498), .Z(n542) );
  CND2IXL U830 ( .B(n704), .A(n3575), .Z(n2819) );
  CND2XL U831 ( .A(n2812), .B(n2791), .Z(n704) );
  CND2IXL U832 ( .B(n705), .A(n3575), .Z(n3601) );
  CND3XL U833 ( .A(n3578), .B(n3576), .C(n3269), .Z(n705) );
  CDLY1XL U834 ( .A(q0[3]), .Z(n1094) );
  CND2XL U835 ( .A(n2933), .B(n2932), .Z(n2934) );
  CIVX2 U836 ( .A(n2177), .Z(n706) );
  CNR2IXL U837 ( .B(n1361), .A(n707), .Z(n1362) );
  CND2X1 U838 ( .A(n2411), .B(n706), .Z(n707) );
  CDLY1XL U839 ( .A(q0[1]), .Z(n710) );
  COND1X1 U840 ( .A(n3325), .B(n2738), .C(n2737), .Z(n550) );
  CND2X2 U841 ( .A(n2588), .B(n2549), .Z(n1105) );
  CND2X2 U842 ( .A(n2588), .B(n2549), .Z(n3002) );
  CND3XL U843 ( .A(n2846), .B(n2840), .C(n2845), .Z(n563) );
  COND3XL U844 ( .A(n3295), .B(n2839), .C(n2838), .D(n2837), .Z(n2846) );
  CND2X1 U845 ( .A(n3551), .B(n3555), .Z(n3276) );
  CND3X1 U846 ( .A(n2623), .B(n2622), .C(n2621), .Z(n559) );
  CND2IX1 U847 ( .B(n2606), .A(n3288), .Z(n2623) );
  CND4X2 U848 ( .A(n2387), .B(n2386), .C(n2385), .D(n2384), .Z(n2388) );
  CIVXL U849 ( .A(n1632), .Z(n709) );
  CNR2XL U850 ( .A(n2940), .B(n3431), .Z(n2941) );
  CNR2XL U851 ( .A(n2937), .B(n3431), .Z(n2812) );
  CNR2XL U852 ( .A(n3431), .B(n3325), .Z(n3430) );
  CND2X1 U853 ( .A(n2580), .B(n3060), .Z(n714) );
  CIVX3 U854 ( .A(n1341), .Z(n1395) );
  CND3X1 U855 ( .A(n2030), .B(n2029), .C(n2028), .Z(n711) );
  CND3X1 U856 ( .A(n2030), .B(n2029), .C(n2028), .Z(n2522) );
  CND3X1 U857 ( .A(n2197), .B(n1869), .C(n999), .Z(n1852) );
  CND2X1 U858 ( .A(n2138), .B(n1922), .Z(n2197) );
  CIVXL U859 ( .A(n2321), .Z(n2661) );
  CND3X1 U860 ( .A(n1871), .B(n1868), .C(n2018), .Z(n1854) );
  CNR2X2 U861 ( .A(n2032), .B(n2033), .Z(n1155) );
  CANR1X1 U862 ( .A(n2180), .B(n2179), .C(n2178), .Z(n712) );
  CIVX2 U863 ( .A(n2370), .Z(n2175) );
  CNR2X1 U864 ( .A(n2434), .B(n2177), .Z(n2178) );
  CIVX2 U865 ( .A(n3030), .Z(n2745) );
  CNR3X1 U866 ( .A(n2605), .B(n2604), .C(n2603), .Z(n713) );
  CND2X2 U867 ( .A(n2013), .B(n2368), .Z(n1909) );
  CNIVX1 U868 ( .A(n648), .Z(n715) );
  CNIVX1 U869 ( .A(n653), .Z(n716) );
  CNIVX1 U870 ( .A(n658), .Z(n717) );
  CNIVX1 U871 ( .A(n663), .Z(n718) );
  CNIVX1 U872 ( .A(n3627), .Z(n719) );
  CNIVX1 U873 ( .A(n2539), .Z(n720) );
  CNIVX1 U874 ( .A(n2524), .Z(n721) );
  CNIVX1 U875 ( .A(n1017), .Z(n722) );
  CNIVX1 U876 ( .A(n1710), .Z(n723) );
  CNIVX1 U877 ( .A(n1711), .Z(n724) );
  CNIVX1 U878 ( .A(n1712), .Z(n725) );
  CNIVX1 U879 ( .A(n1713), .Z(n726) );
  CNIVX1 U880 ( .A(n1714), .Z(n727) );
  CNIVX1 U881 ( .A(n1715), .Z(n728) );
  CNIVX1 U882 ( .A(n1716), .Z(n729) );
  CNIVX1 U883 ( .A(n1718), .Z(n730) );
  CNIVX1 U884 ( .A(n1719), .Z(n731) );
  CNIVX1 U885 ( .A(n1720), .Z(n732) );
  CNIVX1 U886 ( .A(n734), .Z(n733) );
  CNIVX1 U887 ( .A(n1721), .Z(n734) );
  CNIVX1 U888 ( .A(n736), .Z(n735) );
  CNIVX1 U889 ( .A(n1722), .Z(n736) );
  CNIVX1 U890 ( .A(n738), .Z(n737) );
  CNIVX1 U891 ( .A(n1723), .Z(n738) );
  CNIVX1 U892 ( .A(n740), .Z(n739) );
  CNIVX1 U893 ( .A(n1724), .Z(n740) );
  CNIVX1 U894 ( .A(n742), .Z(n741) );
  CNIVX1 U895 ( .A(n1725), .Z(n742) );
  CNIVX1 U896 ( .A(n744), .Z(n743) );
  CNIVX1 U897 ( .A(n1726), .Z(n744) );
  CNIVX1 U898 ( .A(n746), .Z(n745) );
  CNIVX1 U899 ( .A(n1727), .Z(n746) );
  CNIVX1 U900 ( .A(n748), .Z(n747) );
  CNIVX1 U901 ( .A(n1728), .Z(n748) );
  CNIVX1 U902 ( .A(n750), .Z(n749) );
  CNIVX1 U903 ( .A(n1729), .Z(n750) );
  CNIVX1 U904 ( .A(n752), .Z(n751) );
  CNIVX1 U905 ( .A(n1730), .Z(n752) );
  CNIVX1 U906 ( .A(n754), .Z(n753) );
  CNIVX1 U907 ( .A(n1731), .Z(n754) );
  CNIVX1 U908 ( .A(n756), .Z(n755) );
  CNIVX1 U909 ( .A(n1732), .Z(n756) );
  CNIVX1 U910 ( .A(n758), .Z(n757) );
  CNIVX1 U911 ( .A(n1733), .Z(n758) );
  CNIVX1 U912 ( .A(n760), .Z(n759) );
  CNIVX1 U913 ( .A(n1734), .Z(n760) );
  CNIVX1 U914 ( .A(n762), .Z(n761) );
  CNIVX1 U915 ( .A(n1735), .Z(n762) );
  CNIVX1 U916 ( .A(n764), .Z(n763) );
  CNIVX1 U917 ( .A(n1736), .Z(n764) );
  CNIVX1 U918 ( .A(n766), .Z(n765) );
  CNIVX1 U919 ( .A(n1737), .Z(n766) );
  CNIVX3 U920 ( .A(n1738), .Z(n767) );
  CNIVX3 U921 ( .A(n1739), .Z(n768) );
  CNIVX3 U922 ( .A(n1740), .Z(n769) );
  CNIVX3 U923 ( .A(n1741), .Z(n770) );
  CNIVX3 U924 ( .A(n1742), .Z(n771) );
  CNIVX3 U925 ( .A(n1743), .Z(n772) );
  CNIVX3 U926 ( .A(n1744), .Z(n773) );
  CNIVX1 U927 ( .A(n1745), .Z(n774) );
  CNIVX1 U928 ( .A(n1747), .Z(n775) );
  CNIVX1 U929 ( .A(n1709), .Z(n776) );
  CNIVX1 U930 ( .A(n1707), .Z(n777) );
  CNIVX1 U931 ( .A(n500), .Z(n778) );
  CMX2XL U932 ( .A0(h1[5]), .A1(h2[5]), .S(rst), .Z(n503) );
  CNIVX1 U933 ( .A(n503), .Z(n779) );
  CNIVX1 U934 ( .A(n504), .Z(n780) );
  CNIVX1 U935 ( .A(n3626), .Z(n781) );
  CNIVX1 U936 ( .A(n1211), .Z(n782) );
  CNIVX1 U937 ( .A(n662), .Z(n783) );
  CNIVX1 U938 ( .A(n664), .Z(n784) );
  CNIVX1 U939 ( .A(n657), .Z(n785) );
  CNIVX1 U940 ( .A(n659), .Z(n786) );
  CNIVX1 U941 ( .A(n660), .Z(n787) );
  CNIVX1 U942 ( .A(n661), .Z(n788) );
  CNIVX1 U943 ( .A(n652), .Z(n789) );
  CNIVX1 U944 ( .A(n654), .Z(n790) );
  CNIVX1 U945 ( .A(n655), .Z(n791) );
  CNIVX1 U946 ( .A(n656), .Z(n792) );
  CNIVX1 U947 ( .A(n647), .Z(n793) );
  CNIVX1 U948 ( .A(n649), .Z(n794) );
  CNIVX1 U949 ( .A(n650), .Z(n795) );
  CNIVX1 U950 ( .A(n651), .Z(n796) );
  CNIVX1 U951 ( .A(n642), .Z(n797) );
  CNIVX1 U952 ( .A(n643), .Z(n798) );
  CNIVX1 U953 ( .A(n644), .Z(n799) );
  CNIVX1 U954 ( .A(n645), .Z(n800) );
  CNIVX1 U955 ( .A(n646), .Z(n801) );
  CNIVX1 U956 ( .A(n665), .Z(n802) );
  CMX2X2 U957 ( .A0(n803), .A1(z[0]), .S(n3435), .Z(n666) );
  CNIVXL U958 ( .A(acc[0]), .Z(n803) );
  CNIVX1 U959 ( .A(n639), .Z(n804) );
  CNIVX1 U960 ( .A(n640), .Z(n805) );
  CNIVX1 U961 ( .A(n641), .Z(n806) );
  CNIVX1 U962 ( .A(n634), .Z(n807) );
  CNIVX1 U963 ( .A(n636), .Z(n808) );
  CMX2X2 U964 ( .A0(n1140), .A1(z[29]), .S(n3435), .Z(n637) );
  CNIVX1 U965 ( .A(n638), .Z(n809) );
  CNIVX3 U966 ( .A(cmd0[0]), .Z(n811) );
  CNIVX1 U967 ( .A(n811), .Z(n810) );
  CNIVX1 U968 ( .A(n813), .Z(n812) );
  CNIVX1 U969 ( .A(n814), .Z(n813) );
  CNIVX1 U970 ( .A(h0[0]), .Z(n814) );
  CNIVX1 U971 ( .A(n816), .Z(n815) );
  CNIVX1 U972 ( .A(n817), .Z(n816) );
  CNIVX1 U973 ( .A(h0[2]), .Z(n817) );
  CNIVX1 U974 ( .A(n819), .Z(n818) );
  CNIVX1 U975 ( .A(n820), .Z(n819) );
  CNIVX1 U976 ( .A(h0[1]), .Z(n820) );
  CNIVX3 U977 ( .A(push_0), .Z(n822) );
  CNIVX1 U978 ( .A(n822), .Z(n821) );
  CNIVX3 U979 ( .A(cmd_1[0]), .Z(n824) );
  CNIVX1 U980 ( .A(n824), .Z(n823) );
  CNIVX3 U981 ( .A(cmd0[1]), .Z(n826) );
  CNIVX1 U982 ( .A(n826), .Z(n825) );
  CNIVX1 U983 ( .A(n828), .Z(n827) );
  CNIVX1 U984 ( .A(n829), .Z(n828) );
  CNIVX1 U985 ( .A(h0[5]), .Z(n829) );
  CNIVX3 U986 ( .A(push_1), .Z(n831) );
  CNIVX1 U987 ( .A(n831), .Z(n830) );
  CNIVX3 U988 ( .A(cmd_1[1]), .Z(n833) );
  CNIVX1 U989 ( .A(n833), .Z(n832) );
  CNIVX1 U990 ( .A(n835), .Z(n834) );
  CNIVX1 U991 ( .A(n836), .Z(n835) );
  CNIVX1 U992 ( .A(h0[4]), .Z(n836) );
  CNIVX1 U993 ( .A(n838), .Z(n837) );
  CNIVX1 U994 ( .A(n839), .Z(n838) );
  CNIVX1 U995 ( .A(h0[3]), .Z(n839) );
  CNIVX1 U996 ( .A(n841), .Z(n840) );
  CNIVX1 U997 ( .A(n842), .Z(n841) );
  CNIVX1 U998 ( .A(h0[6]), .Z(n842) );
  CNIVX1 U999 ( .A(n1746), .Z(n843) );
  CNIVX1 U1000 ( .A(n2907), .Z(n844) );
  CNIVXL U1001 ( .A(n3374), .Z(n845) );
  CNIVX1 U1002 ( .A(n1058), .Z(n846) );
  CANR2XL U1003 ( .A(n3617), .B(acc[47]), .C(n1659), .D(mulout[47]), .Z(n1058)
         );
  CNIVX1 U1004 ( .A(n1748), .Z(n847) );
  CNIVX1 U1005 ( .A(n1749), .Z(n848) );
  CNIVX1 U1006 ( .A(n1750), .Z(n849) );
  CND4X2 U1007 ( .A(n2581), .B(n2590), .C(n2873), .D(n2379), .Z(n1069) );
  COND1X2 U1008 ( .A(n2396), .B(n2402), .C(n850), .Z(n2590) );
  CND2X2 U1009 ( .A(n2363), .B(n3573), .Z(n850) );
  CND2X2 U1010 ( .A(n852), .B(n851), .Z(n2402) );
  CIVX2 U1011 ( .A(n1953), .Z(n851) );
  CIVX2 U1012 ( .A(n1952), .Z(n852) );
  CND2X2 U1013 ( .A(n855), .B(n853), .Z(n2873) );
  CND2IX1 U1014 ( .B(n854), .A(n3574), .Z(n853) );
  CIVX2 U1015 ( .A(n2435), .Z(n854) );
  CND2X1 U1016 ( .A(n2376), .B(n2671), .Z(n855) );
  CND2X2 U1017 ( .A(n2583), .B(n2584), .Z(n2379) );
  CND2X2 U1018 ( .A(n2375), .B(n3573), .Z(n2584) );
  CND2IX1 U1019 ( .B(n2374), .A(n2413), .Z(n2583) );
  CND2X2 U1020 ( .A(n2367), .B(n2366), .Z(n2581) );
  CND2XL U1021 ( .A(n2365), .B(n2979), .Z(n2366) );
  COR2X1 U1022 ( .A(n2396), .B(n2364), .Z(n2367) );
  CNR2X2 U1023 ( .A(n1844), .B(n856), .Z(n2136) );
  CIVX2 U1024 ( .A(n1845), .Z(n856) );
  CIVX2 U1025 ( .A(n1845), .Z(n1323) );
  CNR2X2 U1026 ( .A(n1322), .B(n1321), .Z(n1845) );
  CND2X2 U1027 ( .A(n857), .B(n2099), .Z(n1926) );
  CND2X2 U1028 ( .A(n857), .B(n1922), .Z(n1425) );
  CIVX2 U1029 ( .A(n2103), .Z(n857) );
  CAN2X2 U1030 ( .A(n2102), .B(n2101), .Z(n2108) );
  CANR1X2 U1031 ( .A(n2007), .B(n2040), .C(n2763), .Z(n1985) );
  CIVXL U1032 ( .A(n2208), .Z(n859) );
  CND2X1 U1033 ( .A(n1813), .B(n1812), .Z(n1817) );
  COND1X1 U1034 ( .A(n2068), .B(n1821), .C(n2337), .Z(n1822) );
  CND2X1 U1035 ( .A(n1403), .B(n1402), .Z(n1840) );
  CIVX2 U1036 ( .A(n2172), .Z(n2122) );
  CNIVXL U1037 ( .A(n2417), .Z(n3387) );
  CNIVX1 U1038 ( .A(push_2), .Z(n3580) );
  CNR2X1 U1039 ( .A(n1632), .B(acc[33]), .Z(n1321) );
  CND2X1 U1040 ( .A(n1200), .B(n2983), .Z(n1352) );
  CND2X1 U1041 ( .A(n2025), .B(n2024), .Z(n2027) );
  CND2X1 U1042 ( .A(n1891), .B(n2368), .Z(n1542) );
  CNR2X1 U1043 ( .A(n2119), .B(n2118), .Z(n2120) );
  COND1XL U1044 ( .A(n2117), .B(n2155), .C(n2116), .Z(n2118) );
  CNR2X1 U1045 ( .A(n919), .B(n920), .Z(n1843) );
  CND2X1 U1046 ( .A(n1383), .B(n1382), .Z(n1838) );
  COND1X1 U1047 ( .A(n1862), .B(n1861), .C(n2161), .Z(n1863) );
  CND3XL U1048 ( .A(n1623), .B(n1622), .C(n1621), .Z(n1078) );
  CAN2X1 U1049 ( .A(n1629), .B(n1628), .Z(n1630) );
  CNIVX1 U1050 ( .A(n2402), .Z(n2978) );
  CND2IX1 U1051 ( .B(n1762), .A(n1761), .Z(n1763) );
  COND1X1 U1052 ( .A(n2636), .B(n3588), .C(n3262), .Z(n2491) );
  COND1XL U1053 ( .A(n2473), .B(n2779), .C(n2472), .Z(n3064) );
  CND2X1 U1054 ( .A(n1776), .B(n2099), .Z(n2204) );
  CAN2X1 U1055 ( .A(n1773), .B(n1772), .Z(n1774) );
  CND2X1 U1056 ( .A(n2369), .B(n2122), .Z(n1699) );
  CND2X1 U1057 ( .A(n2319), .B(n2086), .Z(n1835) );
  COND1X1 U1058 ( .A(n1841), .B(n1840), .C(n2007), .Z(n1865) );
  COND1XL U1059 ( .A(n1937), .B(n1936), .C(n2125), .Z(n1938) );
  COND1XL U1060 ( .A(n1935), .B(n1934), .C(n2122), .Z(n1939) );
  CIVDX1 U1061 ( .A(n1757), .Z0(n2312), .Z1(n2176) );
  COND1XL U1062 ( .A(n2427), .B(n2426), .C(n2268), .Z(n1178) );
  CNIVX1 U1063 ( .A(n2552), .Z(n2572) );
  COND1XL U1064 ( .A(n2533), .B(n3452), .C(n2532), .Z(n3381) );
  CNIVX1 U1065 ( .A(n1070), .Z(n1192) );
  CIVX2 U1066 ( .A(n3620), .Z(n1085) );
  CNIVX1 U1067 ( .A(pushin), .Z(n3624) );
  CANR1XL U1068 ( .A(n3595), .B(n3056), .C(n3055), .Z(n3057) );
  CENX1 U1069 ( .A(n1186), .B(n1133), .Z(n1664) );
  CND3XL U1070 ( .A(n2311), .B(n2310), .C(n2309), .Z(n556) );
  CIVXL U1071 ( .A(n2151), .Z(n860) );
  COR3X1 U1072 ( .A(n1525), .B(n1524), .C(n860), .Z(n2112) );
  CNR2XL U1073 ( .A(n1632), .B(n1384), .Z(n861) );
  CNR2XL U1074 ( .A(n1625), .B(n1616), .Z(n862) );
  CNR2X1 U1075 ( .A(n861), .B(n862), .Z(n1836) );
  CNR2XL U1076 ( .A(acc[38]), .B(n1611), .Z(n863) );
  CNR2X1 U1077 ( .A(n1547), .B(acc[35]), .Z(n864) );
  CNR2X2 U1078 ( .A(n863), .B(n864), .Z(n1842) );
  CIVX1 U1079 ( .A(n3068), .Z(n865) );
  CANR1X1 U1080 ( .A(n3063), .B(n3069), .C(n865), .Z(n2870) );
  CANR11X1 U1081 ( .A(n1308), .B(n1310), .C(n1309), .D(n2129), .Z(n866) );
  CND2XL U1082 ( .A(n2337), .B(n1291), .Z(n867) );
  CNR2X2 U1083 ( .A(n866), .B(n867), .Z(n2024) );
  CND2IX1 U1084 ( .B(cmd_2[0]), .A(cmd_2[1]), .Z(n3247) );
  CND2XL U1085 ( .A(n2625), .B(n2624), .Z(n868) );
  CENX1 U1086 ( .A(n3591), .B(n868), .Z(n869) );
  CND2X1 U1087 ( .A(n3595), .B(n869), .Z(n2628) );
  CANR2XL U1088 ( .A(acc[32]), .B(n3617), .C(mulout[32]), .D(n1659), .Z(n870)
         );
  CND2X1 U1089 ( .A(n3515), .B(n3514), .Z(n871) );
  CEOXL U1090 ( .A(n3614), .B(n871), .Z(n872) );
  CND2X1 U1091 ( .A(n3595), .B(n872), .Z(n873) );
  COND3XL U1092 ( .A(n3513), .B(n3520), .C(n870), .D(n873), .Z(n3516) );
  CNR2IXL U1093 ( .B(n3376), .A(n3375), .Z(n874) );
  CENX1 U1094 ( .A(n3452), .B(n874), .Z(n3377) );
  CANR1XL U1095 ( .A(n2456), .B(n3504), .C(n2465), .Z(n875) );
  CNR2IXL U1096 ( .B(n3214), .A(n3215), .Z(n876) );
  CENX1 U1097 ( .A(n875), .B(n876), .Z(n877) );
  CND2X1 U1098 ( .A(n3595), .B(n877), .Z(n2283) );
  CNR2XL U1099 ( .A(n1633), .B(acc[0]), .Z(n878) );
  CNR2XL U1100 ( .A(n1634), .B(acc[3]), .Z(n879) );
  CNR2X1 U1101 ( .A(n878), .B(n879), .Z(n1635) );
  CND2XL U1102 ( .A(n1899), .B(n2137), .Z(n880) );
  COND1XL U1103 ( .A(n1810), .B(n1811), .C(n2371), .Z(n881) );
  CND2X1 U1104 ( .A(n880), .B(n881), .Z(n1979) );
  COND1XL U1105 ( .A(n3169), .B(n3174), .C(n3170), .Z(n882) );
  CANR1X1 U1106 ( .A(n2724), .B(n3173), .C(n882), .Z(n3237) );
  CND2XL U1107 ( .A(h2[5]), .B(n3353), .Z(n883) );
  CND4XL U1108 ( .A(n3354), .B(n3356), .C(n3355), .D(n883), .Z(n3402) );
  CNR3X1 U1109 ( .A(n3297), .B(n2836), .C(n2835), .Z(n884) );
  CND3XL U1110 ( .A(n2822), .B(n2823), .C(n884), .Z(n2838) );
  CND3XL U1111 ( .A(n3529), .B(n3604), .C(n3530), .Z(n885) );
  CEOXL U1112 ( .A(n3528), .B(n885), .Z(n886) );
  CNR2XL U1113 ( .A(n3531), .B(n886), .Z(n3535) );
  CND2X1 U1114 ( .A(n2912), .B(n2911), .Z(n887) );
  CND2XL U1115 ( .A(n887), .B(n2910), .Z(n888) );
  CND2IXL U1116 ( .B(n2908), .A(n2909), .Z(n889) );
  CENX1 U1117 ( .A(n888), .B(n889), .Z(n2913) );
  CNR2IXL U1118 ( .B(n2575), .A(n2574), .Z(n890) );
  CND2XL U1119 ( .A(n2625), .B(n3591), .Z(n891) );
  CND2XL U1120 ( .A(n891), .B(n2624), .Z(n892) );
  COND1XL U1121 ( .A(n890), .B(n892), .C(n3595), .Z(n893) );
  CANR1XL U1122 ( .A(n890), .B(n892), .C(n893), .Z(n2577) );
  CIVXL U1123 ( .A(n3614), .Z(n894) );
  CANR1XL U1124 ( .A(n3610), .B(n894), .C(n3612), .Z(n895) );
  CND2XL U1125 ( .A(n2872), .B(n3613), .Z(n896) );
  COND1XL U1126 ( .A(n895), .B(n896), .C(n3595), .Z(n897) );
  CANR1XL U1127 ( .A(n895), .B(n896), .C(n897), .Z(n2876) );
  CNR2XL U1128 ( .A(n3398), .B(n3400), .Z(n898) );
  COND1XL U1129 ( .A(n3398), .B(n3401), .C(n3399), .Z(n899) );
  CANR1XL U1130 ( .A(n3504), .B(n898), .C(n899), .Z(n900) );
  CNR2IXL U1131 ( .B(n3090), .A(n3089), .Z(n901) );
  CENX1 U1132 ( .A(n900), .B(n901), .Z(n3096) );
  CND2IXL U1133 ( .B(n858), .A(n1196), .Z(n1537) );
  CNR2X1 U1134 ( .A(n2747), .B(n2750), .Z(n902) );
  CND3X1 U1135 ( .A(n2748), .B(n2664), .C(n902), .Z(n2665) );
  CND3X2 U1136 ( .A(n2042), .B(n2050), .C(n2041), .Z(n903) );
  CND2X2 U1137 ( .A(n1067), .B(n2059), .Z(n904) );
  CND3X2 U1138 ( .A(n904), .B(n2337), .C(n903), .Z(n2825) );
  CANR11XL U1139 ( .A(n2967), .B(n3060), .C(n1097), .D(n2877), .Z(n905) );
  CNR2XL U1140 ( .A(n1560), .B(n3580), .Z(n906) );
  CANR1XL U1141 ( .A(n1659), .B(mulout[38]), .C(n906), .Z(n907) );
  CND2IX1 U1142 ( .B(n905), .A(n907), .Z(n2875) );
  CANR1XL U1143 ( .A(n3333), .B(n3591), .C(n3332), .Z(n908) );
  CNR2IXL U1144 ( .B(n3331), .A(n3330), .Z(n909) );
  CENX1 U1145 ( .A(n908), .B(n909), .Z(n3334) );
  COND1XL U1146 ( .A(n2971), .B(n3614), .C(n2970), .Z(n910) );
  CND2XL U1147 ( .A(n2972), .B(n3065), .Z(n911) );
  CENX1 U1148 ( .A(n910), .B(n911), .Z(n2973) );
  CIVX1 U1149 ( .A(n3504), .Z(n912) );
  COND1XL U1150 ( .A(n3400), .B(n912), .C(n3401), .Z(n913) );
  CND2IXL U1151 ( .B(n3398), .A(n3399), .Z(n914) );
  CENX1 U1152 ( .A(n913), .B(n914), .Z(n915) );
  CND2X1 U1153 ( .A(n3595), .B(n915), .Z(n3408) );
  CND2X1 U1154 ( .A(n3380), .B(n3381), .Z(n916) );
  CND2XL U1155 ( .A(n916), .B(n3379), .Z(n917) );
  CND2IXL U1156 ( .B(n2525), .A(n2526), .Z(n918) );
  CENX1 U1157 ( .A(n917), .B(n918), .Z(n2534) );
  CNR2IX1 U1158 ( .B(acc[18]), .A(n1611), .Z(n1369) );
  CNR2XL U1159 ( .A(n1632), .B(acc[37]), .Z(n919) );
  CNR2XL U1160 ( .A(n1195), .B(acc[36]), .Z(n920) );
  CND3X2 U1161 ( .A(n1646), .B(n1644), .C(n1645), .Z(n921) );
  CNR2XL U1162 ( .A(n2069), .B(n1818), .Z(n922) );
  CNR2X2 U1163 ( .A(n921), .B(n922), .Z(n1666) );
  CND3XL U1164 ( .A(n2411), .B(n2412), .C(n2413), .Z(n923) );
  CND2XL U1165 ( .A(n3250), .B(n2435), .Z(n924) );
  CND2X1 U1166 ( .A(n924), .B(n923), .Z(n3348) );
  CAN3XL U1167 ( .A(n3394), .B(n3393), .C(n3395), .Z(n3403) );
  CIVXL U1168 ( .A(n3346), .Z(n925) );
  CIVXL U1169 ( .A(n3344), .Z(n926) );
  COND1XL U1170 ( .A(n3346), .B(n926), .C(n3345), .Z(n927) );
  CANR11XL U1171 ( .A(n3343), .B(n3591), .C(n925), .D(n927), .Z(n928) );
  CNR2IXL U1172 ( .B(n3342), .A(n3341), .Z(n929) );
  CENX1 U1173 ( .A(n928), .B(n929), .Z(n3347) );
  CND2XL U1174 ( .A(n3613), .B(n3610), .Z(n930) );
  CANR1XL U1175 ( .A(n3613), .B(n3612), .C(n3611), .Z(n931) );
  COND1XL U1176 ( .A(n3614), .B(n930), .C(n931), .Z(n932) );
  CND2XL U1177 ( .A(n3615), .B(n3616), .Z(n933) );
  CENX1 U1178 ( .A(n932), .B(n933), .Z(n3619) );
  COND1XL U1179 ( .A(n3365), .B(n3366), .C(n3364), .Z(n934) );
  CNR2XL U1180 ( .A(n3363), .B(n3366), .Z(n935) );
  CANR1XL U1181 ( .A(n3504), .B(n935), .C(n934), .Z(n936) );
  CNR2IXL U1182 ( .B(n3362), .A(n3361), .Z(n937) );
  CENX1 U1183 ( .A(n936), .B(n937), .Z(n3367) );
  CNR2X1 U1184 ( .A(n3386), .B(n3580), .Z(n938) );
  CANR1XL U1185 ( .A(mulout[14]), .B(n1659), .C(n938), .Z(n939) );
  COND4CXL U1186 ( .A(n3387), .B(n3445), .C(n3388), .D(n939), .Z(n3389) );
  CND2X1 U1187 ( .A(n2528), .B(n3455), .Z(n940) );
  CND2X1 U1188 ( .A(n2530), .B(n3455), .Z(n941) );
  COND3XL U1189 ( .A(n3452), .B(n940), .C(n3454), .D(n941), .Z(n942) );
  CND2IXL U1190 ( .B(n2304), .A(n2305), .Z(n943) );
  CENX1 U1191 ( .A(n942), .B(n943), .Z(n2307) );
  CIVXL U1192 ( .A(n3297), .Z(n944) );
  CANR11XL U1193 ( .A(n3269), .B(n1124), .C(n944), .D(n3298), .Z(n945) );
  COND3XL U1194 ( .A(n1086), .B(n1085), .C(n945), .D(n1087), .Z(n564) );
  COND2XL U1195 ( .A(n2155), .B(n1783), .C(n2003), .D(n2117), .Z(n946) );
  CNR2IXL U1196 ( .B(n2113), .A(n1128), .Z(n947) );
  COND1X1 U1197 ( .A(n946), .B(n947), .C(n2018), .Z(n1784) );
  CND2XL U1198 ( .A(n1196), .B(n1163), .Z(n948) );
  CND2XL U1199 ( .A(n1595), .B(n2983), .Z(n949) );
  CND3X2 U1200 ( .A(n948), .B(n1579), .C(n949), .Z(n1892) );
  CNR2XL U1201 ( .A(n3569), .B(n2747), .Z(n950) );
  CND2X1 U1202 ( .A(n3572), .B(n950), .Z(n2937) );
  CNR2IXL U1203 ( .B(n2916), .A(n2918), .Z(n2931) );
  CANR2XL U1204 ( .A(n3617), .B(acc[10]), .C(n1659), .D(mulout[10]), .Z(n951)
         );
  COND1XL U1205 ( .A(n3281), .B(n2618), .C(n951), .Z(n2619) );
  CNR3XL U1206 ( .A(n3531), .B(n2786), .C(n1097), .Z(n2776) );
  COR3X1 U1207 ( .A(n3360), .B(n3325), .C(n3357), .Z(n2519) );
  CND3XL U1208 ( .A(n2688), .B(n1176), .C(n3513), .Z(n952) );
  CND2XL U1209 ( .A(n1110), .B(n3269), .Z(n953) );
  CIVXL U1210 ( .A(n2924), .Z(n954) );
  CIVXL U1211 ( .A(n2926), .Z(n955) );
  COND1XL U1212 ( .A(n2924), .B(n955), .C(n2925), .Z(n956) );
  CANR11XL U1213 ( .A(n2927), .B(n3504), .C(n954), .D(n956), .Z(n957) );
  CNR2IXL U1214 ( .B(n2733), .A(n2732), .Z(n958) );
  CENX1 U1215 ( .A(n957), .B(n958), .Z(n2736) );
  CND2XL U1216 ( .A(n3445), .B(n3387), .Z(n959) );
  CNR3XL U1217 ( .A(n1151), .B(n3325), .C(n959), .Z(n3383) );
  COND1XL U1218 ( .A(n3453), .B(n3452), .C(n3451), .Z(n960) );
  CND2XL U1219 ( .A(n3454), .B(n3455), .Z(n961) );
  CENX1 U1220 ( .A(n960), .B(n961), .Z(n3459) );
  CND2IXL U1221 ( .B(n2224), .A(n2223), .Z(n1704) );
  CNR2XL U1222 ( .A(n1532), .B(n1531), .Z(n962) );
  CEOXL U1223 ( .A(n962), .B(n1673), .Z(n963) );
  CANR2XL U1224 ( .A(n3617), .B(acc[1]), .C(mulout[1]), .D(n1659), .Z(n964) );
  COND1XL U1225 ( .A(n963), .B(n3325), .C(n964), .Z(n965) );
  CEOX1 U1226 ( .A(n1672), .B(n1674), .Z(n966) );
  CNR2IXL U1227 ( .B(acc[15]), .A(n1459), .Z(n1370) );
  CNR2XL U1228 ( .A(n2129), .B(n2344), .Z(n967) );
  CND3XL U1229 ( .A(n1962), .B(n1961), .C(n967), .Z(n1965) );
  CAN2XL U1230 ( .A(n2552), .B(n2568), .Z(n2550) );
  CNR2X1 U1231 ( .A(n3580), .B(n2454), .Z(n968) );
  CANR1XL U1232 ( .A(mulout[53]), .B(n1659), .C(n968), .Z(n969) );
  COND3X1 U1233 ( .A(n2452), .B(n3261), .C(n2453), .D(n969), .Z(n2498) );
  CND2IXL U1234 ( .B(n2222), .A(n2225), .Z(n1660) );
  CNR2XL U1235 ( .A(n3554), .B(n3325), .Z(n970) );
  CND3XL U1236 ( .A(n3432), .B(n3431), .C(n970), .Z(n3433) );
  CANR2XL U1237 ( .A(mulout[35]), .B(n1659), .C(acc[35]), .D(n3617), .Z(n971)
         );
  CANR1XL U1238 ( .A(n2782), .B(n2781), .C(n2780), .Z(n972) );
  CND2XL U1239 ( .A(n2782), .B(n2778), .Z(n973) );
  COND1XL U1240 ( .A(n3614), .B(n973), .C(n972), .Z(n974) );
  CND2X1 U1241 ( .A(n2784), .B(n2783), .Z(n975) );
  CENX1 U1242 ( .A(n974), .B(n975), .Z(n976) );
  CND2X1 U1243 ( .A(n3620), .B(n976), .Z(n977) );
  CND2X1 U1244 ( .A(n971), .B(n977), .Z(n2785) );
  CANR1XL U1245 ( .A(n3591), .B(n3343), .C(n3344), .Z(n978) );
  CND2XL U1246 ( .A(n3345), .B(n2770), .Z(n979) );
  COND1XL U1247 ( .A(n978), .B(n979), .C(n3620), .Z(n980) );
  CANR1XL U1248 ( .A(n978), .B(n979), .C(n980), .Z(n1207) );
  CND2XL U1249 ( .A(mulout[27]), .B(n1659), .Z(n981) );
  COND1XL U1250 ( .A(n3495), .B(n3580), .C(n981), .Z(n3496) );
  CNR2X1 U1251 ( .A(n2507), .B(n2506), .Z(n982) );
  CND2XL U1252 ( .A(n2508), .B(h2[5]), .Z(n983) );
  CND2X1 U1253 ( .A(n982), .B(n983), .Z(n3360) );
  CANR1XL U1254 ( .A(n2927), .B(n3504), .C(n2926), .Z(n984) );
  CNR2IXL U1255 ( .B(n2925), .A(n2924), .Z(n985) );
  CENX1 U1256 ( .A(n984), .B(n985), .Z(n2928) );
  CANR2XL U1257 ( .A(acc[9]), .B(n3617), .C(mulout[9]), .D(n1659), .Z(n986) );
  COND1XL U1258 ( .A(n3375), .B(n3452), .C(n3376), .Z(n987) );
  CNR2IX1 U1259 ( .B(n3283), .A(n3282), .Z(n988) );
  COND1XL U1260 ( .A(n987), .B(n988), .C(n3595), .Z(n989) );
  COND4CX1 U1261 ( .A(n988), .B(n987), .C(n989), .D(n986), .Z(n3284) );
  CND2IX1 U1262 ( .B(n3247), .A(push_2), .Z(n3531) );
  CANR2X1 U1263 ( .A(n803), .B(n3617), .C(mulout[0]), .D(n1659), .Z(n990) );
  COND3XL U1264 ( .A(n2181), .B(n2028), .C(n1673), .D(n3269), .Z(n991) );
  COND3XL U1265 ( .A(n803), .B(mulout[0]), .C(n3595), .D(n1674), .Z(n992) );
  CAN3XL U1266 ( .A(n990), .B(n991), .C(n992), .Z(n1211) );
  CND2XL U1267 ( .A(n3439), .B(n3438), .Z(n993) );
  CENX1 U1268 ( .A(n3440), .B(n993), .Z(n994) );
  COND1XL U1269 ( .A(n3580), .B(n3442), .C(n3441), .Z(n995) );
  CANR1XL U1270 ( .A(n994), .B(n3595), .C(n995), .Z(n996) );
  CEOXL U1271 ( .A(n3437), .B(n1124), .Z(n997) );
  COND1XL U1272 ( .A(n3325), .B(n997), .C(n996), .Z(n565) );
  CND2XL U1273 ( .A(n1553), .B(acc[8]), .Z(n1629) );
  CNR2IX1 U1274 ( .B(acc[28]), .A(n1617), .Z(n1604) );
  COND1XL U1275 ( .A(n2427), .B(n2426), .C(n2268), .Z(n998) );
  CND3X1 U1276 ( .A(n2439), .B(n2552), .C(n998), .Z(n2440) );
  CNR2IXL U1277 ( .B(n2151), .A(n2152), .Z(n2157) );
  CND3XL U1278 ( .A(n1845), .B(n2368), .C(n1846), .Z(n999) );
  CND2IXL U1279 ( .B(n2072), .A(n1501), .Z(n2075) );
  CND2IXL U1280 ( .B(n2458), .A(n2457), .Z(n2255) );
  CNR3XL U1281 ( .A(n3554), .B(n3326), .C(n3325), .Z(n1000) );
  CND2XL U1282 ( .A(n3329), .B(n1000), .Z(n3339) );
  CND2XL U1283 ( .A(n2549), .B(n2550), .Z(n1001) );
  CNR2XL U1284 ( .A(n1001), .B(n2551), .Z(n1002) );
  CMXI2XL U1285 ( .A0(n1002), .A1(n2563), .S(n3015), .Z(n2565) );
  CANR1XL U1286 ( .A(n2946), .B(n3240), .C(n2758), .Z(n1003) );
  CND2XL U1287 ( .A(n2757), .B(n2756), .Z(n1004) );
  CEOXL U1288 ( .A(n1003), .B(n1004), .Z(n2759) );
  COND1XL U1289 ( .A(n2777), .B(n3614), .C(n2779), .Z(n1005) );
  CND2XL U1290 ( .A(n2596), .B(n2782), .Z(n1006) );
  CENX1 U1291 ( .A(n1005), .B(n1006), .Z(n2599) );
  CNR2XL U1292 ( .A(n2507), .B(n2509), .Z(n1007) );
  CND2XL U1293 ( .A(n2380), .B(h2[5]), .Z(n1008) );
  CND2X1 U1294 ( .A(n1007), .B(n1008), .Z(n3359) );
  CND2XL U1295 ( .A(n3503), .B(n3502), .Z(n1009) );
  CENX1 U1296 ( .A(n3504), .B(n1009), .Z(n3508) );
  CND2XL U1297 ( .A(n3380), .B(n3379), .Z(n1010) );
  CENX1 U1298 ( .A(n3381), .B(n1010), .Z(n1011) );
  CAN2X1 U1299 ( .A(n3595), .B(n1011), .Z(n3382) );
  CND2X1 U1300 ( .A(n3440), .B(n3439), .Z(n1012) );
  CNR2IXL U1301 ( .B(n3293), .A(n3292), .Z(n1013) );
  CND2XL U1302 ( .A(n3438), .B(n1012), .Z(n1014) );
  CENX1 U1303 ( .A(n1013), .B(n1014), .Z(n1086) );
  CND2XL U1304 ( .A(n2823), .B(n2290), .Z(n1015) );
  CENX1 U1305 ( .A(n1082), .B(n1015), .Z(n1016) );
  CANR2XL U1306 ( .A(n3617), .B(acc[3]), .C(mulout[3]), .D(n1659), .Z(n1017)
         );
  CENX1 U1307 ( .A(n1705), .B(n1704), .Z(n1018) );
  CND2X1 U1308 ( .A(n1018), .B(n3595), .Z(n1019) );
  COND3XL U1309 ( .A(n3531), .B(n1016), .C(n722), .D(n1019), .Z(n1706) );
  CNR2XL U1310 ( .A(n1391), .B(n1634), .Z(n1020) );
  CNR2XL U1311 ( .A(n1633), .B(n3473), .Z(n1021) );
  CNR2XL U1312 ( .A(n1020), .B(n1021), .Z(n1394) );
  CND2XL U1313 ( .A(n1995), .B(n2368), .Z(n1022) );
  CND2X1 U1314 ( .A(n1917), .B(n1022), .Z(n1120) );
  CIVX1 U1315 ( .A(n1120), .Z(n1121) );
  CNR2XL U1316 ( .A(n1459), .B(acc[58]), .Z(n1024) );
  CNR2X2 U1317 ( .A(n1023), .B(n1024), .Z(n1271) );
  CND2XL U1318 ( .A(n3250), .B(n2582), .Z(n1025) );
  CND3XL U1319 ( .A(n1025), .B(n2584), .C(n2583), .Z(n3513) );
  CNR2XL U1320 ( .A(n2507), .B(n2282), .Z(n1026) );
  CND2XL U1321 ( .A(n2189), .B(n2349), .Z(n1027) );
  CND2X1 U1322 ( .A(n1026), .B(n1027), .Z(n3225) );
  CND2X1 U1323 ( .A(n1659), .B(mulout[59]), .Z(n1028) );
  COND1XL U1324 ( .A(n3580), .B(n1066), .C(n1028), .Z(n2656) );
  CND2XL U1325 ( .A(mulout[31]), .B(n1659), .Z(n1029) );
  COND1XL U1326 ( .A(n3580), .B(n3054), .C(n1029), .Z(n3055) );
  CIVX1 U1327 ( .A(n2270), .Z(n1030) );
  COND1XL U1328 ( .A(n3101), .B(n3207), .C(n1030), .Z(n2274) );
  CND2IX1 U1329 ( .B(n1670), .A(n1671), .Z(n1672) );
  CNR2IXL U1330 ( .B(n2863), .A(n3325), .Z(n2930) );
  CND4XL U1331 ( .A(n2572), .B(n3269), .C(n2765), .D(n2631), .Z(n1031) );
  CNR2XL U1332 ( .A(n3542), .B(n2541), .Z(n1032) );
  COND1XL U1333 ( .A(n3542), .B(n2542), .C(n3543), .Z(n1033) );
  CANR1XL U1334 ( .A(n3538), .B(n1032), .C(n1033), .Z(n1034) );
  CND2X1 U1335 ( .A(n3536), .B(n1032), .Z(n1035) );
  COND1XL U1336 ( .A(n3614), .B(n1035), .C(n1034), .Z(n1036) );
  CND2IXL U1337 ( .B(n2543), .A(n2544), .Z(n1037) );
  CENX1 U1338 ( .A(n1036), .B(n1037), .Z(n1038) );
  CND2X1 U1339 ( .A(n3620), .B(n1038), .Z(n2547) );
  CND3X1 U1340 ( .A(n3575), .B(n3269), .C(n3340), .Z(n3352) );
  CIVXL U1341 ( .A(n3359), .Z(n1039) );
  CNR3XL U1342 ( .A(n3325), .B(n3360), .C(n1039), .Z(n2517) );
  COND1XL U1343 ( .A(n3563), .B(n3562), .C(n3561), .Z(n1040) );
  CNR2XL U1344 ( .A(n3563), .B(n3560), .Z(n1041) );
  CANR1XL U1345 ( .A(n3591), .B(n1041), .C(n1040), .Z(n1042) );
  CNR2IXL U1346 ( .B(n3559), .A(n3558), .Z(n1043) );
  CENX1 U1347 ( .A(n1042), .B(n1043), .Z(n3565) );
  CND2XL U1348 ( .A(mulout[34]), .B(n1659), .Z(n1044) );
  COND1XL U1349 ( .A(n3580), .B(n2597), .C(n1044), .Z(n2598) );
  CND2XL U1350 ( .A(mulout[19]), .B(n1659), .Z(n1045) );
  COND1XL U1351 ( .A(n3580), .B(n2734), .C(n1045), .Z(n2735) );
  CND2XL U1352 ( .A(n2905), .B(n3444), .Z(n1046) );
  CNR2X1 U1353 ( .A(n3463), .B(n1046), .Z(n3385) );
  CNR2IXL U1354 ( .B(n3465), .A(n3467), .Z(n1047) );
  CENX1 U1355 ( .A(n3466), .B(n1047), .Z(n2844) );
  CANR2XL U1356 ( .A(n3554), .B(n3430), .C(n3595), .D(n3429), .Z(n1048) );
  CND3XL U1357 ( .A(n3433), .B(n3434), .C(n1048), .Z(n514) );
  CND2IX1 U1358 ( .B(n2058), .A(n2137), .Z(n1262) );
  CAN3X1 U1359 ( .A(n1623), .B(n1621), .C(n1622), .Z(n1983) );
  CAOR2X1 U1360 ( .A(n1401), .B(acc[11]), .C(n1455), .D(acc[14]), .Z(n1841) );
  CNR2IX1 U1361 ( .B(n2983), .A(n1547), .Z(n1277) );
  CNR2IX1 U1362 ( .B(n2410), .A(n3248), .Z(n2412) );
  CNR2IX1 U1363 ( .B(n3172), .A(n3176), .Z(n3178) );
  CND2X1 U1364 ( .A(n3529), .B(n3528), .Z(n1049) );
  CNR2X1 U1365 ( .A(n2548), .B(n1049), .Z(n2568) );
  CND2IX1 U1366 ( .B(n2891), .A(n2892), .Z(n2893) );
  CNR2X1 U1367 ( .A(n3076), .B(n3075), .Z(n1050) );
  CND2X1 U1368 ( .A(n3083), .B(n3269), .Z(n1051) );
  CNR2X1 U1369 ( .A(n1050), .B(n1051), .Z(n3077) );
  CND2IX1 U1370 ( .B(n3212), .A(n3213), .Z(n3219) );
  CNR2X1 U1371 ( .A(n2521), .B(n2520), .Z(n2849) );
  CND2IX1 U1372 ( .B(n2824), .A(n1115), .Z(n2835) );
  CNR3XL U1373 ( .A(n3015), .B(n3530), .C(n3325), .Z(n3017) );
  CND2X1 U1374 ( .A(n2719), .B(n3236), .Z(n1052) );
  CEOX1 U1375 ( .A(n2727), .B(n1052), .Z(n1053) );
  CND2X1 U1376 ( .A(n3595), .B(n1053), .Z(n2730) );
  CANR2X1 U1377 ( .A(mulout[46]), .B(n1659), .C(n3617), .D(acc[46]), .Z(n1054)
         );
  CND2X1 U1378 ( .A(n2769), .B(n1054), .Z(n1055) );
  CND2X1 U1379 ( .A(n2768), .B(n1054), .Z(n1056) );
  COND1XL U1380 ( .A(n2766), .B(n1055), .C(n1056), .Z(n2771) );
  CNR2IX1 U1381 ( .B(n2930), .A(n2931), .Z(n2932) );
  CNR3XL U1382 ( .A(n3325), .B(n1102), .C(n3387), .Z(n2308) );
  CND3XL U1383 ( .A(n3443), .B(n3464), .C(n3281), .Z(n3285) );
  CND2IX1 U1384 ( .B(n3468), .A(n3469), .Z(n3470) );
  CND3XL U1385 ( .A(n2277), .B(n3206), .C(n2276), .Z(n1057) );
  CND3XL U1386 ( .A(n2273), .B(n2274), .C(n1057), .Z(n540) );
  CND2X1 U1387 ( .A(n3595), .B(n3347), .Z(n1059) );
  CND4X1 U1388 ( .A(n3352), .B(n3351), .C(n846), .D(n1059), .Z(n522) );
  CND3XL U1389 ( .A(n3357), .B(n2518), .C(n3360), .Z(n1060) );
  CNR2X1 U1390 ( .A(n2517), .B(n2516), .Z(n1061) );
  CND3XL U1391 ( .A(n2519), .B(n1060), .C(n1061), .Z(n549) );
  CIVX2 U1392 ( .A(n3132), .Z(n1062) );
  COR2X1 U1393 ( .A(n2147), .B(n2004), .Z(n1794) );
  CND2XL U1394 ( .A(n2004), .B(n2169), .Z(n1248) );
  CIVXL U1395 ( .A(n2604), .Z(n1063) );
  CIVXL U1396 ( .A(n1063), .Z(n1064) );
  CND3X2 U1397 ( .A(n1873), .B(n1872), .C(n2337), .Z(n2603) );
  CND2X1 U1398 ( .A(n1200), .B(n1066), .Z(n1585) );
  CND2IXL U1399 ( .B(n3321), .A(n2998), .Z(n2999) );
  CND2X2 U1400 ( .A(n1998), .B(n1997), .Z(n1999) );
  CND2IX1 U1401 ( .B(n2001), .A(n2368), .Z(n2345) );
  CND2IX1 U1402 ( .B(n3554), .A(n3329), .Z(n3321) );
  CND2X1 U1403 ( .A(n1122), .B(n2631), .Z(n2318) );
  CND2X1 U1404 ( .A(n1991), .B(n2344), .Z(n1761) );
  CNR2X2 U1405 ( .A(n1614), .B(n1613), .Z(n1067) );
  CNR2X1 U1406 ( .A(n1614), .B(n1613), .Z(n2040) );
  CIVXL U1407 ( .A(n3129), .Z(n1068) );
  CND2IXL U1408 ( .B(n2301), .A(n2300), .Z(n2311) );
  CNR2XL U1409 ( .A(n3385), .B(n3388), .Z(n3390) );
  CIVXL U1410 ( .A(n1098), .Z(n1070) );
  CNR2X2 U1411 ( .A(n2832), .B(n2830), .Z(n1071) );
  CNR2X2 U1412 ( .A(n2832), .B(n2830), .Z(n2097) );
  CIVX3 U1413 ( .A(n2553), .Z(n2585) );
  CANR1X1 U1414 ( .A(n2349), .B(n2189), .C(n2507), .Z(n1074) );
  CNR2XL U1415 ( .A(n1219), .B(n1218), .Z(n1075) );
  CND2IX1 U1416 ( .B(n2195), .A(n1076), .Z(n2322) );
  COAN1XL U1417 ( .A(n2172), .B(n1860), .C(n1859), .Z(n1076) );
  CND2XL U1418 ( .A(n1878), .B(n2371), .Z(n1765) );
  CNIVXL U1419 ( .A(q0[25]), .Z(n1077) );
  CND3XL U1420 ( .A(n1623), .B(n1622), .C(n1621), .Z(n1079) );
  CNR2IX1 U1421 ( .B(n1980), .A(n1979), .Z(n1989) );
  CND2XL U1422 ( .A(n2690), .B(n2688), .Z(n2705) );
  CNIVXL U1423 ( .A(n2821), .Z(n1082) );
  CND2X2 U1424 ( .A(n1903), .B(n1902), .Z(n2506) );
  CND2X1 U1425 ( .A(n2388), .B(n2344), .Z(n1903) );
  CMX2XL U1426 ( .A0(h1[2]), .A1(h2[2]), .S(rst), .Z(n500) );
  CNR2IX1 U1427 ( .B(n1109), .A(n1625), .Z(n1344) );
  CND2XL U1428 ( .A(n2173), .B(n2371), .Z(n1698) );
  CNR2XL U1429 ( .A(n2173), .B(n2172), .Z(n2174) );
  CND2XL U1430 ( .A(n1580), .B(acc[3]), .Z(n1386) );
  COND1XL U1431 ( .A(n2172), .B(n1860), .C(n1859), .Z(n2194) );
  CNR2X2 U1432 ( .A(n2316), .B(n2763), .Z(n2631) );
  CND3X1 U1433 ( .A(n1253), .B(n1252), .C(n1251), .Z(n1254) );
  CNR2X2 U1434 ( .A(n1214), .B(h2[0]), .Z(n1084) );
  CNR2X2 U1435 ( .A(n1214), .B(h2[0]), .Z(n1312) );
  CND4XL U1436 ( .A(n3295), .B(n3437), .C(n3269), .D(n3297), .Z(n1087) );
  COAN1XL U1437 ( .A(n2121), .B(n2363), .C(n703), .Z(n1090) );
  CND2X2 U1438 ( .A(n1149), .B(n2099), .Z(n2198) );
  CND3XL U1439 ( .A(n2999), .B(n3001), .C(n3000), .Z(n519) );
  CNR3X2 U1440 ( .A(n3431), .B(n2949), .C(n2943), .Z(n2748) );
  CND2XL U1441 ( .A(n3385), .B(n2308), .Z(n2309) );
  CND2XL U1442 ( .A(n3385), .B(n3445), .Z(n2300) );
  COND1X1 U1443 ( .A(n3287), .B(n1144), .C(n2610), .Z(n2622) );
  CND2X2 U1444 ( .A(n3529), .B(n3528), .Z(n1091) );
  CNR2IX2 U1445 ( .B(n1092), .A(n2831), .Z(n3437) );
  COAN1XL U1446 ( .A(n1160), .B(n2828), .C(n2827), .Z(n1092) );
  CNR2X2 U1447 ( .A(n2063), .B(n2062), .Z(n1115) );
  CIVX2 U1448 ( .A(n2443), .Z(n1093) );
  CND2X2 U1449 ( .A(n2350), .B(n2349), .Z(n2355) );
  CND3X1 U1450 ( .A(n1271), .B(n1270), .C(n1269), .Z(n1095) );
  CND3X1 U1451 ( .A(n1271), .B(n1270), .C(n1269), .Z(n2011) );
  CND2X1 U1452 ( .A(n2188), .B(n2187), .Z(n3126) );
  CND4X2 U1453 ( .A(n2346), .B(n2347), .C(n2268), .D(n2345), .Z(n2010) );
  CND2X1 U1454 ( .A(n1967), .B(n2034), .Z(n1970) );
  CIVXL U1455 ( .A(n2874), .Z(n1096) );
  CIVX2 U1456 ( .A(n1096), .Z(n1097) );
  CIVX3 U1457 ( .A(h2[1]), .Z(n1098) );
  CIVX4 U1458 ( .A(h2[1]), .Z(n1214) );
  CNR2IX2 U1459 ( .B(n1194), .A(n1819), .Z(n1823) );
  CNIVXL U1460 ( .A(n2607), .Z(n1099) );
  COND1X1 U1461 ( .A(n2706), .B(n1864), .C(n1698), .Z(n1876) );
  CND3X2 U1462 ( .A(n3395), .B(n3393), .C(n1921), .Z(n1943) );
  CANR1X2 U1463 ( .A(n1121), .B(n1920), .C(n2507), .Z(n3393) );
  CND4X2 U1464 ( .A(n2581), .B(n2590), .C(n2379), .D(n2873), .Z(n1100) );
  CND2X1 U1465 ( .A(n1569), .B(n1568), .Z(n1756) );
  CIVXL U1466 ( .A(n1595), .Z(n1101) );
  CNR2X2 U1467 ( .A(n1477), .B(acc[46]), .Z(n1213) );
  CND3X2 U1468 ( .A(n1062), .B(n2209), .C(n2210), .Z(n1103) );
  CND3X1 U1469 ( .A(n2211), .B(n2209), .C(n2210), .Z(n1104) );
  CND3XL U1470 ( .A(n859), .B(n2211), .C(n2210), .Z(n2674) );
  CANR1X1 U1471 ( .A(n2703), .B(n3058), .C(n2702), .Z(n2704) );
  COND1X1 U1472 ( .A(n2087), .B(n1249), .C(n1248), .Z(n1264) );
  CND2XL U1473 ( .A(n1456), .B(acc[21]), .Z(n1457) );
  CND2XL U1474 ( .A(n1456), .B(acc[18]), .Z(n1253) );
  CND2X2 U1475 ( .A(h2[0]), .B(h2[1]), .Z(n1106) );
  CND2X2 U1476 ( .A(h2[1]), .B(h2[0]), .Z(n1341) );
  CND2XL U1477 ( .A(n2123), .B(n2122), .Z(n2216) );
  CND2X1 U1478 ( .A(n2123), .B(n2368), .Z(n1772) );
  CND2X2 U1479 ( .A(n1481), .B(n1480), .Z(n2123) );
  COND1XL U1480 ( .A(n1838), .B(n1837), .C(n2113), .Z(n1107) );
  CNR2X2 U1481 ( .A(n2087), .B(h2[4]), .Z(n2113) );
  CND2X2 U1482 ( .A(n1437), .B(n1173), .Z(n2104) );
  CNIVXL U1483 ( .A(n2590), .Z(n1110) );
  CND2X2 U1484 ( .A(n1197), .B(n3631), .Z(n1572) );
  CND3X4 U1485 ( .A(n1768), .B(n1767), .C(n1766), .Z(n3101) );
  CND2X2 U1486 ( .A(n2039), .B(n2038), .Z(n2826) );
  CIVXL U1487 ( .A(n3353), .Z(n1111) );
  CND2XL U1488 ( .A(n1183), .B(n2096), .Z(n2821) );
  CND2X1 U1489 ( .A(n1752), .B(n2122), .Z(n1562) );
  CND2X2 U1490 ( .A(n2416), .B(n2415), .Z(n2676) );
  CNR2X2 U1491 ( .A(n2282), .B(n3126), .Z(n2416) );
  CND2XL U1492 ( .A(n2321), .B(h2[5]), .Z(n2185) );
  CND2X1 U1493 ( .A(n1643), .B(acc[8]), .Z(n1306) );
  CND2X2 U1494 ( .A(n2221), .B(n2349), .Z(n2439) );
  CIVX2 U1495 ( .A(n2609), .Z(n1112) );
  CIVX2 U1496 ( .A(n2745), .Z(n1168) );
  CNR2X1 U1497 ( .A(n2049), .B(n2336), .Z(n1920) );
  CANR1XL U1498 ( .A(n2349), .B(n2190), .C(n2507), .Z(n1113) );
  CIVXL U1499 ( .A(n3443), .Z(n1114) );
  CND2X1 U1500 ( .A(n2104), .B(n1893), .Z(n1438) );
  CND2XL U1501 ( .A(n3232), .B(n3231), .Z(n544) );
  COND1X1 U1502 ( .A(n2087), .B(n1864), .C(n1863), .Z(n2195) );
  CNR3X1 U1503 ( .A(n1100), .B(n714), .C(n2401), .Z(n1116) );
  CNR3X1 U1504 ( .A(n1100), .B(n2401), .C(n714), .Z(n1171) );
  CND3X1 U1505 ( .A(n2347), .B(n2346), .C(n2345), .Z(n2348) );
  CNR2X2 U1506 ( .A(n2200), .B(n2199), .Z(n2278) );
  CNR2X2 U1507 ( .A(n1617), .B(n2597), .Z(n1226) );
  CIVXL U1508 ( .A(n3102), .Z(n1117) );
  CND3X2 U1509 ( .A(n1071), .B(n2096), .C(n2095), .Z(n1118) );
  CND3X1 U1510 ( .A(n2097), .B(n2096), .C(n2095), .Z(n2444) );
  CND2X1 U1511 ( .A(n2123), .B(n2371), .Z(n1923) );
  CND2X1 U1512 ( .A(n1894), .B(n2373), .Z(n1760) );
  COAN1XL U1513 ( .A(n3416), .B(n3432), .C(n3415), .Z(n3434) );
  CND3X2 U1514 ( .A(n2356), .B(n2355), .C(n2354), .Z(n1184) );
  CAN3XL U1515 ( .A(n1075), .B(n1221), .C(n1220), .Z(n1119) );
  CND2XL U1516 ( .A(n1570), .B(n1473), .Z(n1358) );
  CNR3X2 U1517 ( .A(n1904), .B(n2509), .C(n2506), .Z(n1122) );
  CND2X1 U1518 ( .A(n2104), .B(n2099), .Z(n1769) );
  CND2X1 U1519 ( .A(n1475), .B(n1474), .Z(n1476) );
  CND2IXL U1520 ( .B(n3002), .A(n2776), .Z(n2790) );
  CND3XL U1521 ( .A(n3020), .B(n3019), .C(n3018), .Z(n529) );
  CND4X1 U1522 ( .A(n2407), .B(n2404), .C(n2405), .D(n2406), .Z(n1592) );
  CNR2IX1 U1523 ( .B(n2344), .A(n2365), .Z(n1948) );
  CND2XL U1524 ( .A(n2100), .B(n2371), .Z(n1451) );
  CND2XL U1525 ( .A(n2100), .B(n2099), .Z(n2101) );
  CND2X1 U1526 ( .A(n2098), .B(n2122), .Z(n2102) );
  CND2IX1 U1527 ( .B(n1123), .A(n2571), .Z(n2579) );
  CAOR2XL U1528 ( .A(mulout[45]), .B(n1659), .C(n858), .D(n3617), .Z(n1123) );
  CND2X1 U1529 ( .A(n2823), .B(n2822), .Z(n1124) );
  CANR1XL U1530 ( .A(n2787), .B(n2786), .C(n2785), .Z(n2789) );
  CIVX2 U1531 ( .A(n1125), .Z(n1127) );
  CIVXL U1532 ( .A(n2110), .Z(n1128) );
  CNR2X2 U1533 ( .A(n1936), .B(n1937), .Z(n2110) );
  CND4X1 U1534 ( .A(n1789), .B(n1791), .C(n1790), .D(n1788), .Z(n1129) );
  CND4XL U1535 ( .A(n1790), .B(n1791), .C(n1789), .D(n1788), .Z(n1130) );
  CIVXL U1536 ( .A(n2323), .Z(n1131) );
  CND2XL U1537 ( .A(n1517), .B(acc[10]), .Z(n1511) );
  CND2XL U1538 ( .A(n1517), .B(acc[12]), .Z(n1403) );
  CND2XL U1539 ( .A(n1517), .B(acc[8]), .Z(n1392) );
  CND2XL U1540 ( .A(n1517), .B(acc[18]), .Z(n1461) );
  CND2X1 U1541 ( .A(n2201), .B(n2349), .Z(n2206) );
  COR2X1 U1542 ( .A(n2183), .B(n2184), .Z(n1132) );
  CNR2X2 U1543 ( .A(n1617), .B(n1597), .Z(n1598) );
  CND2IX2 U1544 ( .B(n1887), .A(n1886), .Z(n1888) );
  CIVX2 U1545 ( .A(n2823), .Z(n1133) );
  CND2X1 U1546 ( .A(n2124), .B(n2125), .Z(n1914) );
  CIVXL U1547 ( .A(n2207), .Z(n1134) );
  CNR2X1 U1548 ( .A(n1547), .B(acc[41]), .Z(n1135) );
  CIVXL U1549 ( .A(n2943), .Z(n1136) );
  CIVX2 U1550 ( .A(n1136), .Z(n1137) );
  CIVX2 U1551 ( .A(n1138), .Z(n1140) );
  CNR2X2 U1552 ( .A(n2561), .B(n2560), .Z(n1141) );
  CNR2X2 U1553 ( .A(n2561), .B(n2560), .Z(n3522) );
  CND2IXL U1554 ( .B(n1547), .A(acc[32]), .Z(n1551) );
  CIVXL U1555 ( .A(n3384), .Z(n1142) );
  CIVXL U1556 ( .A(n1142), .Z(n1143) );
  CND2X2 U1557 ( .A(n3443), .B(n3464), .Z(n3372) );
  CNR2X1 U1558 ( .A(acc[32]), .B(n1625), .Z(n1322) );
  CND2X2 U1559 ( .A(n1156), .B(n2275), .Z(n3207) );
  CIVXL U1560 ( .A(n2277), .Z(n1145) );
  CND4X1 U1561 ( .A(n1912), .B(n1911), .C(n1910), .D(n1909), .Z(n1146) );
  CIVDX2 U1562 ( .A(n1502), .Z0(n1555), .Z1(n1200) );
  CND4X1 U1563 ( .A(n1912), .B(n1911), .C(n1910), .D(n1909), .Z(n2045) );
  CNR2XL U1564 ( .A(n1883), .B(n1882), .Z(n1147) );
  CANR1X2 U1565 ( .A(h2[5]), .B(n2380), .C(n2507), .Z(n1148) );
  CND2X1 U1566 ( .A(n1078), .B(n2176), .Z(n1898) );
  CND2XL U1567 ( .A(n1078), .B(n1922), .Z(n1944) );
  CND2X2 U1568 ( .A(n1381), .B(n1380), .Z(n1149) );
  CND2X2 U1569 ( .A(n1381), .B(n1380), .Z(n2148) );
  CAN2X2 U1570 ( .A(n1702), .B(n1701), .Z(n2096) );
  CNR2X1 U1571 ( .A(n1885), .B(n1884), .Z(n1886) );
  CNR2X1 U1572 ( .A(n1596), .B(n1167), .Z(n1412) );
  CND2X1 U1573 ( .A(n1235), .B(n1234), .Z(n1905) );
  CAN2X1 U1574 ( .A(n2496), .B(n3620), .Z(n2497) );
  CEOX1 U1575 ( .A(n2494), .B(n2493), .Z(n2496) );
  COND1XL U1576 ( .A(n2087), .B(n1864), .C(n1863), .Z(n1150) );
  CND2IX1 U1577 ( .B(n2687), .A(n1201), .Z(n2690) );
  CNIVXL U1578 ( .A(n1143), .Z(n1151) );
  CND2X2 U1579 ( .A(n1519), .B(n1518), .Z(n1525) );
  CND3XL U1580 ( .A(n1846), .B(n1845), .C(n2368), .Z(n1152) );
  CIVX2 U1581 ( .A(n1844), .Z(n1846) );
  CND2X1 U1582 ( .A(n1437), .B(n1173), .Z(n1153) );
  COND1X1 U1583 ( .A(n3325), .B(n3510), .C(n3509), .Z(n553) );
  CND2IXL U1584 ( .B(n1624), .A(acc[14]), .Z(n1654) );
  CIVXL U1585 ( .A(n2795), .Z(n1154) );
  CNIVX1 U1586 ( .A(n3060), .Z(n3083) );
  CNR2X2 U1587 ( .A(n2032), .B(n2033), .Z(n1156) );
  CIVXL U1588 ( .A(n1090), .Z(n1157) );
  CANR1X1 U1589 ( .A(n2090), .B(n2339), .C(n1782), .Z(n1785) );
  CND3X1 U1590 ( .A(n2742), .B(n1168), .C(n2741), .Z(n2744) );
  CND3X2 U1591 ( .A(n2593), .B(n1171), .C(n3522), .Z(n3015) );
  CIVXL U1592 ( .A(n3500), .Z(n1158) );
  CIVXL U1593 ( .A(n1158), .Z(n1159) );
  CND3XL U1594 ( .A(n1896), .B(n1897), .C(n1898), .Z(n1160) );
  CNR3X2 U1595 ( .A(n3022), .B(n2977), .C(n3340), .Z(n3329) );
  CND2XL U1596 ( .A(n2339), .B(h2[5]), .Z(n2192) );
  CND2X1 U1597 ( .A(n1361), .B(n2411), .Z(n1161) );
  CND2X1 U1598 ( .A(n2372), .B(n2137), .Z(n1361) );
  CND2X2 U1599 ( .A(n2168), .B(n2169), .Z(n2411) );
  CND3X1 U1600 ( .A(n1230), .B(n1228), .C(n1229), .Z(n1164) );
  CND3X1 U1601 ( .A(n1229), .B(n1230), .C(n1228), .Z(n1996) );
  CND2X2 U1602 ( .A(n1165), .B(n1612), .Z(n1613) );
  COR2X1 U1603 ( .A(n2734), .B(n1611), .Z(n1165) );
  CND2XL U1604 ( .A(n1164), .B(n1893), .Z(n1804) );
  CND2X1 U1605 ( .A(n1996), .B(n2169), .Z(n1997) );
  CND2X2 U1606 ( .A(n1424), .B(n1425), .Z(n1441) );
  CND2XL U1607 ( .A(n3529), .B(n3269), .Z(n2886) );
  CNR2X1 U1608 ( .A(n2500), .B(n2499), .Z(n2502) );
  COND3XL U1609 ( .A(n3414), .B(n3413), .C(n3412), .D(n3411), .Z(n547) );
  CND2XL U1610 ( .A(n3413), .B(n3410), .Z(n3411) );
  CND2XL U1611 ( .A(n3413), .B(n3397), .Z(n3368) );
  CND2X1 U1612 ( .A(n2372), .B(n2169), .Z(n2431) );
  CND2XL U1613 ( .A(n1981), .B(n1893), .Z(n1609) );
  CND2XL U1614 ( .A(n1981), .B(n2014), .Z(n1896) );
  CND2XL U1615 ( .A(n1753), .B(n1751), .Z(n1561) );
  CND2IX1 U1616 ( .B(n2147), .A(n1982), .Z(n1987) );
  CND3X1 U1617 ( .A(n1850), .B(n1849), .C(n1848), .Z(n1169) );
  CND3XL U1618 ( .A(n1850), .B(n1849), .C(n1848), .Z(n2324) );
  CND2X1 U1619 ( .A(n1995), .B(n2125), .Z(n1998) );
  CND2X1 U1620 ( .A(n1677), .B(n1676), .Z(n1887) );
  CND3X1 U1621 ( .A(n2433), .B(n2432), .C(n2431), .Z(n2438) );
  CND2XL U1622 ( .A(n1570), .B(n1181), .Z(n1571) );
  CND2X1 U1623 ( .A(n2015), .B(n2371), .Z(n1912) );
  CIVXL U1624 ( .A(n1196), .Z(n1170) );
  CNR3X2 U1625 ( .A(n1069), .B(n2401), .C(n2400), .Z(n3521) );
  CND2X1 U1626 ( .A(n2138), .B(n2368), .Z(n1678) );
  CND2XL U1627 ( .A(n2138), .B(n2371), .Z(n1961) );
  CND2X1 U1628 ( .A(n1895), .B(n2371), .Z(n1897) );
  CND3X1 U1629 ( .A(n3567), .B(n3568), .C(n3566), .Z(n518) );
  CIVXL U1630 ( .A(n1968), .Z(n1363) );
  CND2X1 U1631 ( .A(n1274), .B(n1273), .Z(n1275) );
  CND2X2 U1632 ( .A(n1357), .B(n1356), .Z(n1697) );
  COAN1X1 U1633 ( .A(n1800), .B(n1095), .C(n1799), .Z(n2332) );
  CND2X2 U1634 ( .A(n2162), .B(n1893), .Z(n1694) );
  CND2X2 U1635 ( .A(n1314), .B(n1313), .Z(n1856) );
  CNR2X1 U1636 ( .A(n1447), .B(n1555), .Z(n1256) );
  CNR2X1 U1637 ( .A(n1555), .B(n1554), .Z(n1556) );
  CNR2X1 U1638 ( .A(n3054), .B(n1555), .Z(n1603) );
  CND2X1 U1639 ( .A(n1435), .B(n1436), .Z(n1172) );
  CIVX2 U1640 ( .A(n1172), .Z(n1173) );
  CND2XL U1641 ( .A(n2568), .B(n1174), .Z(n1210) );
  CNR2XL U1642 ( .A(n2563), .B(n3325), .Z(n1174) );
  COND1X2 U1643 ( .A(n2438), .B(n2437), .C(n2436), .Z(n2552) );
  CNR2IX1 U1644 ( .B(n1355), .A(n1555), .Z(n1479) );
  CIVX2 U1645 ( .A(acc[52]), .Z(n1355) );
  CANR1XL U1646 ( .A(n1990), .B(n1989), .C(n1988), .Z(n1175) );
  CANR1X1 U1647 ( .A(n1990), .B(n1989), .C(n1988), .Z(n2298) );
  CND2XL U1648 ( .A(n3102), .B(n3269), .Z(n3104) );
  CIVX2 U1649 ( .A(n1578), .Z(n1579) );
  CND2XL U1650 ( .A(n2367), .B(n2366), .Z(n1176) );
  CANR2X1 U1651 ( .A(n2015), .B(n2014), .C(n2137), .D(n2013), .Z(n1177) );
  CANR2XL U1652 ( .A(n2015), .B(n2014), .C(n2137), .D(n2013), .Z(n2343) );
  CND2X2 U1653 ( .A(n1594), .B(n1593), .Z(n1669) );
  CND2X1 U1654 ( .A(n2364), .B(n2090), .Z(n1593) );
  CND2XL U1655 ( .A(n2433), .B(n2264), .Z(n2267) );
  COND1X2 U1656 ( .A(n2166), .B(n2165), .C(n2371), .Z(n2265) );
  CND2XL U1657 ( .A(n2136), .B(n2169), .Z(n1179) );
  CNIVXL U1658 ( .A(n2557), .Z(n1182) );
  CND2XL U1659 ( .A(n2852), .B(n2851), .Z(n3501) );
  CNR2XL U1660 ( .A(n1459), .B(n1364), .Z(n1238) );
  CND2XL U1661 ( .A(n2145), .B(n1922), .Z(n1962) );
  CNR2IXL U1662 ( .B(n2146), .A(n2145), .Z(n2150) );
  CND3X1 U1663 ( .A(n3550), .B(n3549), .C(n3548), .Z(n527) );
  CANR11X1 U1664 ( .A(n3608), .B(n3535), .C(n3534), .D(n3533), .Z(n3549) );
  CNR2IX1 U1665 ( .B(n3630), .A(n1634), .Z(n1337) );
  COND11XL U1666 ( .A(n3325), .B(n3437), .C(n3297), .D(n3296), .Z(n3298) );
  CANR1XL U1667 ( .A(n2034), .B(n1690), .C(n1689), .Z(n1183) );
  COND1X1 U1668 ( .A(n3058), .B(n3059), .C(n3057), .Z(n538) );
  CND2X1 U1669 ( .A(n1899), .B(n1922), .Z(n1825) );
  CND3X1 U1670 ( .A(n1607), .B(n1606), .C(n1605), .Z(n1899) );
  CIVXL U1671 ( .A(n1124), .Z(n3295) );
  CNR2X2 U1672 ( .A(n2397), .B(n2396), .Z(n2398) );
  CND2X1 U1673 ( .A(n2439), .B(n2351), .Z(n2557) );
  CNR2IX2 U1674 ( .B(n1654), .A(n1653), .Z(n2037) );
  CND2XL U1675 ( .A(n2126), .B(n2125), .Z(n2217) );
  CDLY1XL U1676 ( .A(h2[0]), .Z(n1185) );
  CND2X2 U1677 ( .A(n1592), .B(h2[5]), .Z(n1955) );
  CND2XL U1678 ( .A(n1508), .B(acc[12]), .Z(n1513) );
  CND2XL U1679 ( .A(n1508), .B(acc[17]), .Z(n1295) );
  CANR2X2 U1680 ( .A(n2322), .B(n2344), .C(n2279), .D(n2278), .Z(n2210) );
  CNR2X2 U1681 ( .A(n1187), .B(n1272), .Z(n1953) );
  COAN1X1 U1682 ( .A(n1268), .B(n1267), .C(n1223), .Z(n1187) );
  CND2XL U1683 ( .A(n2874), .B(n3269), .Z(n3061) );
  CND2X2 U1684 ( .A(n1148), .B(n1881), .Z(n1904) );
  CND2IX1 U1685 ( .B(n1632), .A(acc[15]), .Z(n1518) );
  CNR2XL U1686 ( .A(n2669), .B(n2670), .Z(n1188) );
  CNR2XL U1687 ( .A(n2670), .B(n2669), .Z(n3021) );
  CND2X2 U1688 ( .A(n1445), .B(n1444), .Z(n1935) );
  COR2X1 U1689 ( .A(n2121), .B(n2381), .Z(n1189) );
  COND1X1 U1690 ( .A(n2194), .B(n1150), .C(n2086), .Z(n1873) );
  COND1X2 U1691 ( .A(n2092), .B(n2091), .C(n2090), .Z(n2093) );
  CNR2X1 U1692 ( .A(n3025), .B(n3245), .Z(n2714) );
  CNR2XL U1693 ( .A(n2847), .B(n2848), .Z(n2863) );
  CND2X2 U1694 ( .A(n1955), .B(n3355), .Z(n2850) );
  CND2X1 U1695 ( .A(n1470), .B(n1471), .Z(n1190) );
  CND2X2 U1696 ( .A(n1472), .B(n1191), .Z(n2124) );
  CIVX2 U1697 ( .A(n1190), .Z(n1191) );
  CND2X1 U1698 ( .A(n1503), .B(n2983), .Z(n1475) );
  COND2X1 U1699 ( .A(n1818), .B(n2073), .C(n2069), .D(n1079), .Z(n1824) );
  CIVXL U1700 ( .A(n3031), .Z(n1193) );
  CNR2X1 U1701 ( .A(n1577), .B(acc[53]), .Z(n1276) );
  CND2IXL U1702 ( .B(n3156), .A(n3033), .Z(n3039) );
  CNR2IX1 U1703 ( .B(n3157), .A(n3156), .Z(n3166) );
  COND1XL U1704 ( .A(n3554), .B(n3350), .C(n3349), .Z(n3351) );
  CND2XL U1705 ( .A(n3574), .B(n3573), .Z(n3576) );
  CND3X1 U1706 ( .A(n1202), .B(n2034), .C(n1971), .Z(n1465) );
  CND3X1 U1707 ( .A(n1202), .B(n2349), .C(n1971), .Z(n1972) );
  CANR2X1 U1708 ( .A(n1464), .B(n2014), .C(n2099), .D(n2117), .Z(n1971) );
  CAN2X2 U1709 ( .A(n1141), .B(n2686), .Z(n1199) );
  CNR2IXL U1710 ( .B(n1113), .A(n3126), .Z(n3133) );
  CND2XL U1711 ( .A(n2169), .B(n2002), .Z(n1919) );
  CND2XL U1712 ( .A(n2002), .B(n2368), .Z(n1261) );
  CMX2XL U1713 ( .A0(h1[1]), .A1(n1192), .S(rst), .Z(n499) );
  CNR2X1 U1714 ( .A(n2378), .B(n2377), .Z(n3574) );
  CND2X1 U1715 ( .A(n2012), .B(n2371), .Z(n1789) );
  CND2X1 U1716 ( .A(n2037), .B(n1194), .Z(n2038) );
  CND2IX1 U1717 ( .B(n3023), .A(n1188), .Z(n2743) );
  CNR2X1 U1718 ( .A(n3022), .B(n3023), .Z(n2711) );
  CIVX3 U1719 ( .A(n1195), .Z(n1503) );
  CAN2X2 U1720 ( .A(n2018), .B(n2146), .Z(n1194) );
  CIVDX2 U1721 ( .A(n3531), .Z0(n3269), .Z1(n3325) );
  CIVDX2 U1722 ( .A(n1544), .Z0(n1195), .Z1(n1196) );
  CIVDX4 U1723 ( .A(h2[4]), .Z0(n2121), .Z1(n2344) );
  CIVDX2 U1724 ( .A(n1521), .Z0(n1596), .Z1(n1198) );
  CND2X4 U1725 ( .A(n1231), .B(h2[2]), .Z(n2172) );
  CNR2X2 U1726 ( .A(n1658), .B(cmd_2[0]), .Z(n1659) );
  CIVDX2 U1727 ( .A(n1330), .Z0(n1223), .Z1(n1893) );
  CIVX2 U1728 ( .A(n2018), .Z(n2129) );
  CAN2X1 U1729 ( .A(n1452), .B(n1451), .Z(n1202) );
  CIVX4 U1730 ( .A(n2121), .Z(n2268) );
  CIVDXL U1731 ( .A(n2452), .Z0(n1203), .Z1(n1204) );
  CIVX2 U1732 ( .A(acc[48]), .Z(n1574) );
  CAN2X1 U1733 ( .A(n2730), .B(n2729), .Z(n1205) );
  CIVX2 U1734 ( .A(acc[41]), .Z(n1432) );
  COR2X1 U1735 ( .A(n3506), .B(n1617), .Z(n1206) );
  CIVX2 U1736 ( .A(acc[43]), .Z(n1434) );
  CAN2XL U1737 ( .A(n2994), .B(n3595), .Z(n1208) );
  CEOX1 U1738 ( .A(n2695), .B(n2694), .Z(n1209) );
  CIVX8 U1739 ( .A(n2087), .Z(n2371) );
  CIVX2 U1740 ( .A(n1501), .Z(n2073) );
  CIVDX1 U1741 ( .A(n1796), .Z0(n1396), .Z1(n2161) );
  CND2X2 U1742 ( .A(n2014), .B(n2121), .Z(n2155) );
  CMX2XL U1743 ( .A0(h1[3]), .A1(h2[3]), .S(rst), .Z(n2539) );
  CND2X2 U1744 ( .A(n2388), .B(n2086), .Z(n2094) );
  CIVXL U1745 ( .A(n1810), .Z(n1813) );
  CIVX8 U1746 ( .A(h2[0]), .Z(n1490) );
  CND2X2 U1747 ( .A(n1490), .B(n1214), .Z(n1317) );
  CNIVX4 U1748 ( .A(n1317), .Z(n1477) );
  CIVX2 U1749 ( .A(n1106), .Z(n1502) );
  CIVX2 U1750 ( .A(n1502), .Z(n1611) );
  CNR2X1 U1751 ( .A(n1611), .B(n1162), .Z(n1212) );
  CNR2X2 U1752 ( .A(n1213), .B(n1212), .Z(n1217) );
  CIVX2 U1753 ( .A(n1084), .Z(n1558) );
  CIVX2 U1754 ( .A(n1558), .Z(n1615) );
  CND2X1 U1755 ( .A(n1615), .B(n1574), .Z(n1216) );
  CNR2X4 U1756 ( .A(n1490), .B(h2[1]), .Z(n1544) );
  CIVX2 U1757 ( .A(n1195), .Z(n1567) );
  CIVX1 U1758 ( .A(acc[47]), .Z(n1350) );
  CND2XL U1759 ( .A(n1567), .B(n1350), .Z(n1215) );
  CND3X2 U1760 ( .A(n1217), .B(n1216), .C(n1215), .Z(n2013) );
  CND2X2 U1761 ( .A(h2[2]), .B(h2[3]), .Z(n2087) );
  CND2X1 U1762 ( .A(n2013), .B(n2371), .Z(n1225) );
  CNR2X1 U1763 ( .A(n1477), .B(n1072), .Z(n1219) );
  CNR2X1 U1764 ( .A(n1555), .B(n858), .Z(n1218) );
  CNR2X2 U1765 ( .A(n1219), .B(n1218), .Z(n1222) );
  CND2XL U1766 ( .A(n1567), .B(n1434), .Z(n1221) );
  CIVX2 U1767 ( .A(n1084), .Z(n1624) );
  CIVX2 U1768 ( .A(n1624), .Z(n1595) );
  CND2X1 U1769 ( .A(n1595), .B(n3632), .Z(n1220) );
  CND3X2 U1770 ( .A(n1222), .B(n1221), .C(n1220), .Z(n2000) );
  CIVX2 U1771 ( .A(h2[3]), .Z(n2089) );
  CNR2X2 U1772 ( .A(n2089), .B(h2[2]), .Z(n1330) );
  CIVX4 U1773 ( .A(n1223), .Z(n2368) );
  CND2X1 U1774 ( .A(n2000), .B(n2368), .Z(n1224) );
  CND2X2 U1775 ( .A(n1225), .B(n1224), .Z(n1950) );
  CNR2X1 U1776 ( .A(h2[3]), .B(h2[2]), .Z(n1796) );
  CND2XL U1777 ( .A(n1648), .B(acc[36]), .Z(n1230) );
  CIVX1 U1778 ( .A(acc[37]), .Z(n3073) );
  CNR2X1 U1779 ( .A(n3073), .B(n1611), .Z(n1227) );
  CND2X2 U1780 ( .A(n1490), .B(n1098), .Z(n1459) );
  CNIVX4 U1781 ( .A(n1459), .Z(n1617) );
  CIVX2 U1782 ( .A(acc[34]), .Z(n2597) );
  CNR2X2 U1783 ( .A(n1227), .B(n1226), .Z(n1229) );
  CND2X1 U1784 ( .A(n1196), .B(acc[35]), .Z(n1228) );
  CIVX2 U1785 ( .A(h2[3]), .Z(n1231) );
  CND2X1 U1786 ( .A(n1649), .B(acc[38]), .Z(n1233) );
  CIVX2 U1787 ( .A(n1341), .Z(n1303) );
  CND2X1 U1788 ( .A(n1395), .B(acc[41]), .Z(n1232) );
  CND2X2 U1789 ( .A(n1233), .B(n1232), .Z(n1906) );
  CND2IX1 U1790 ( .B(n1624), .A(n1166), .Z(n1235) );
  CND2XL U1791 ( .A(n1544), .B(acc[39]), .Z(n1234) );
  COR3X1 U1792 ( .A(n2172), .B(n1906), .C(n1905), .Z(n1236) );
  COND1X1 U1793 ( .A(n1563), .B(n1164), .C(n1236), .Z(n1951) );
  CIVX2 U1794 ( .A(h2[5]), .Z(n1916) );
  CNR2X2 U1795 ( .A(n1916), .B(h2[4]), .Z(n2086) );
  COND1X1 U1796 ( .A(n1950), .B(n1951), .C(n2086), .Z(n1266) );
  CIVX8 U1797 ( .A(h2[6]), .Z(n2337) );
  CND2X4 U1798 ( .A(n2337), .B(h2[5]), .Z(n2018) );
  CND2X1 U1799 ( .A(n2018), .B(n2344), .Z(n2064) );
  CIVX1 U1800 ( .A(acc[30]), .Z(n1364) );
  CIVX2 U1801 ( .A(acc[33]), .Z(n2696) );
  CNR2X1 U1802 ( .A(n2696), .B(n1446), .Z(n1237) );
  CNR2X1 U1803 ( .A(n1238), .B(n1237), .Z(n1241) );
  CND2XL U1804 ( .A(n1648), .B(acc[32]), .Z(n1240) );
  CND2XL U1805 ( .A(n1638), .B(acc[31]), .Z(n1239) );
  CND3X1 U1806 ( .A(n1241), .B(n1239), .C(n1240), .Z(n1995) );
  CIVXL U1807 ( .A(n1995), .Z(n1249) );
  CIVX1 U1808 ( .A(acc[22]), .Z(n1242) );
  CIVXL U1809 ( .A(acc[25]), .Z(n3221) );
  CNR2XL U1810 ( .A(n1577), .B(n3221), .Z(n1243) );
  CNR2XL U1811 ( .A(n1244), .B(n1243), .Z(n1247) );
  CND2XL U1812 ( .A(n1648), .B(acc[24]), .Z(n1246) );
  CND2XL U1813 ( .A(n1638), .B(acc[23]), .Z(n1245) );
  CND3X1 U1814 ( .A(n1247), .B(n1245), .C(n1246), .Z(n2004) );
  CIVX2 U1815 ( .A(n2172), .Z(n2169) );
  CND2X1 U1816 ( .A(n1648), .B(acc[20]), .Z(n1250) );
  CIVX2 U1817 ( .A(n1250), .Z(n1255) );
  CND2X2 U1818 ( .A(n1098), .B(n1490), .Z(n1485) );
  CIVXL U1819 ( .A(n1485), .Z(n1456) );
  CND2X1 U1820 ( .A(n1395), .B(acc[21]), .Z(n1252) );
  CND2XL U1821 ( .A(n1544), .B(acc[19]), .Z(n1251) );
  CNR2X2 U1822 ( .A(n1255), .B(n1254), .Z(n2058) );
  CNR2X2 U1823 ( .A(h2[3]), .B(h2[2]), .Z(n1757) );
  CIVX1 U1824 ( .A(acc[26]), .Z(n3136) );
  CNR2X1 U1825 ( .A(n1617), .B(n3136), .Z(n1257) );
  CIVX2 U1826 ( .A(n1139), .Z(n1447) );
  CNR2X1 U1827 ( .A(n1257), .B(n1256), .Z(n1260) );
  CND2XL U1828 ( .A(n1648), .B(acc[28]), .Z(n1259) );
  CND2XL U1829 ( .A(n1196), .B(acc[27]), .Z(n1258) );
  CND3X1 U1830 ( .A(n1258), .B(n1259), .C(n1260), .Z(n2002) );
  CND2X1 U1831 ( .A(n1261), .B(n1262), .Z(n1263) );
  CNR2X2 U1832 ( .A(n1264), .B(n1263), .Z(n1956) );
  CND2IX2 U1833 ( .B(n2064), .A(n1956), .Z(n1265) );
  CND2X2 U1834 ( .A(n1265), .B(n1266), .Z(n2026) );
  CIVX2 U1835 ( .A(n2026), .Z(n1311) );
  CIVX2 U1836 ( .A(n1485), .Z(n1553) );
  CND2XL U1837 ( .A(n1553), .B(acc[62]), .Z(n1797) );
  CND2IXL U1838 ( .B(n2089), .A(n1797), .Z(n1268) );
  CND2X1 U1839 ( .A(n1567), .B(acc[63]), .Z(n1798) );
  CIVXL U1840 ( .A(n1798), .Z(n1267) );
  CND2XL U1841 ( .A(n1567), .B(n1066), .Z(n1270) );
  CND2X1 U1842 ( .A(n1615), .B(n1181), .Z(n1269) );
  CNR2X2 U1843 ( .A(n1095), .B(h2[2]), .Z(n1272) );
  CIVX2 U1844 ( .A(acc[51]), .Z(n1473) );
  CND2X1 U1845 ( .A(n1503), .B(n1473), .Z(n1274) );
  CND2X1 U1846 ( .A(n1581), .B(n1355), .Z(n1273) );
  CIVX2 U1847 ( .A(n1275), .Z(n1279) );
  CNR2X2 U1848 ( .A(n1277), .B(n1276), .Z(n1278) );
  CND2X2 U1849 ( .A(n1279), .B(n1278), .Z(n2015) );
  CND2X1 U1850 ( .A(n2015), .B(n2176), .Z(n1288) );
  CIVX1 U1851 ( .A(acc[55]), .Z(n1469) );
  CND2XL U1852 ( .A(n1567), .B(n1469), .Z(n1281) );
  CND2X1 U1853 ( .A(n1588), .B(n1109), .Z(n1280) );
  CND2X1 U1854 ( .A(n1281), .B(n1280), .Z(n1282) );
  CIVX2 U1855 ( .A(n1282), .Z(n1286) );
  CNR2X1 U1856 ( .A(acc[57]), .B(n1577), .Z(n1284) );
  CNR2X1 U1857 ( .A(n1477), .B(n1088), .Z(n1283) );
  CNR2X2 U1858 ( .A(n1284), .B(n1283), .Z(n1285) );
  CND2X2 U1859 ( .A(n1286), .B(n1285), .Z(n2012) );
  CND2X1 U1860 ( .A(n2012), .B(n2169), .Z(n1287) );
  CND2X2 U1861 ( .A(n1287), .B(n1288), .Z(n1952) );
  CND2X1 U1862 ( .A(h2[5]), .B(h2[4]), .Z(n1758) );
  CIVX2 U1863 ( .A(n1758), .Z(n2090) );
  CND2X2 U1864 ( .A(n2402), .B(n2090), .Z(n2025) );
  CIVX3 U1865 ( .A(n1553), .Z(n1633) );
  COND2XL U1866 ( .A(n1446), .B(acc[5]), .C(acc[2]), .D(n1633), .Z(n1290) );
  CIVX2 U1867 ( .A(n1312), .Z(n1632) );
  COND2XL U1868 ( .A(n1170), .B(acc[3]), .C(acc[4]), .D(n1101), .Z(n1289) );
  CIVDX2 U1869 ( .A(n1757), .Z0(n1675), .Z1(n2137) );
  CNR2X1 U1870 ( .A(n1675), .B(h2[4]), .Z(n2151) );
  CND2X1 U1871 ( .A(n2151), .B(n2018), .Z(n1680) );
  COND1XL U1872 ( .A(n1290), .B(n1289), .C(n2050), .Z(n1291) );
  CND2X1 U1873 ( .A(n1595), .B(acc[16]), .Z(n1293) );
  CND2XL U1874 ( .A(n1567), .B(acc[15]), .Z(n1292) );
  CND2X1 U1875 ( .A(n1293), .B(n1292), .Z(n1297) );
  CIVDX1 U1876 ( .A(n1303), .Z0(n1577), .Z1(n1508) );
  CIVXL U1877 ( .A(n1459), .Z(n1509) );
  CND2XL U1878 ( .A(n1509), .B(acc[14]), .Z(n1294) );
  CND2X1 U1879 ( .A(n1295), .B(n1294), .Z(n1296) );
  CNR2X2 U1880 ( .A(n1297), .B(n1296), .Z(n2052) );
  CND2XL U1881 ( .A(n2052), .B(n2113), .Z(n1310) );
  CND2XL U1882 ( .A(n1503), .B(acc[11]), .Z(n1301) );
  CND2X1 U1883 ( .A(n1595), .B(acc[12]), .Z(n1300) );
  CND2X1 U1884 ( .A(n1197), .B(acc[13]), .Z(n1299) );
  CIVXL U1885 ( .A(n1485), .Z(n1570) );
  CND2XL U1886 ( .A(n1570), .B(acc[10]), .Z(n1298) );
  CND4X1 U1887 ( .A(n1301), .B(n1300), .C(n1299), .D(n1298), .Z(n2053) );
  CIVXL U1888 ( .A(n2053), .Z(n1302) );
  CNR2X4 U1889 ( .A(n1223), .B(h2[4]), .Z(n2146) );
  CND2X1 U1890 ( .A(n1302), .B(n2146), .Z(n1309) );
  CND2XL U1891 ( .A(n1196), .B(acc[7]), .Z(n1307) );
  CIVDX2 U1892 ( .A(n1395), .Z0(n1446), .Z1(n1455) );
  CND2XL U1893 ( .A(n1455), .B(acc[9]), .Z(n1305) );
  CIVXL U1894 ( .A(n1485), .Z(n1649) );
  CND2XL U1895 ( .A(n1649), .B(acc[6]), .Z(n1304) );
  CAN4X1 U1896 ( .A(n1307), .B(n1306), .C(n1305), .D(n1304), .Z(n2051) );
  CIVX2 U1897 ( .A(n2155), .Z(n2007) );
  CND2X1 U1898 ( .A(n2051), .B(n2007), .Z(n1308) );
  CND3X2 U1899 ( .A(n1311), .B(n2025), .C(n2024), .Z(n2820) );
  CNR2X1 U1900 ( .A(n2018), .B(n2344), .Z(n2582) );
  CIVX2 U1901 ( .A(n1312), .Z(n1414) );
  COND2XL U1902 ( .A(n1632), .B(n858), .C(acc[44]), .D(n1195), .Z(n1855) );
  CIVXL U1903 ( .A(n1855), .Z(n1316) );
  CIVDX1 U1904 ( .A(n1303), .Z0(n1634), .Z1(n1197) );
  CIVX2 U1905 ( .A(acc[46]), .Z(n1535) );
  CND2X2 U1906 ( .A(n1198), .B(n1535), .Z(n1314) );
  CIVXL U1907 ( .A(n1459), .Z(n1401) );
  CND2X1 U1908 ( .A(n1401), .B(n1434), .Z(n1313) );
  CIVX2 U1909 ( .A(n1856), .Z(n1315) );
  CND2X2 U1910 ( .A(n1316), .B(n1315), .Z(n2162) );
  CND2X2 U1911 ( .A(n2162), .B(n2371), .Z(n1334) );
  CIVX2 U1912 ( .A(n1317), .Z(n1575) );
  CIVX3 U1913 ( .A(n1575), .Z(n1547) );
  CNR2X1 U1914 ( .A(acc[31]), .B(n1547), .Z(n1318) );
  CIVX2 U1915 ( .A(n1318), .Z(n1320) );
  COR2X1 U1916 ( .A(acc[34]), .B(n1548), .Z(n1319) );
  CND2X2 U1917 ( .A(n1320), .B(n1319), .Z(n1844) );
  CIVDX2 U1918 ( .A(n1544), .Z0(n1625), .Z1(n1638) );
  CNR2X1 U1919 ( .A(h2[3]), .B(h2[2]), .Z(n1695) );
  COND1X2 U1920 ( .A(n1844), .B(n1323), .C(n2125), .Z(n1333) );
  CND2X2 U1921 ( .A(n1843), .B(n1842), .Z(n2140) );
  CIVX2 U1922 ( .A(n2172), .Z(n2014) );
  CND2X2 U1923 ( .A(n2140), .B(n2014), .Z(n1332) );
  CND2X1 U1924 ( .A(n1508), .B(n1073), .Z(n1325) );
  CIVXL U1925 ( .A(n1459), .Z(n1520) );
  CIVX1 U1926 ( .A(acc[39]), .Z(n1554) );
  CND2X1 U1927 ( .A(n1520), .B(n1554), .Z(n1324) );
  CND2X2 U1928 ( .A(n1325), .B(n1324), .Z(n1861) );
  CIVX2 U1929 ( .A(n1861), .Z(n1329) );
  CND2X1 U1930 ( .A(n1196), .B(n1167), .Z(n1327) );
  CIVX2 U1931 ( .A(n1414), .Z(n1581) );
  CND2X1 U1932 ( .A(n1581), .B(n1432), .Z(n1326) );
  CND2X2 U1933 ( .A(n1327), .B(n1326), .Z(n1862) );
  CIVX2 U1934 ( .A(n1862), .Z(n1328) );
  CND2X2 U1935 ( .A(n1329), .B(n1328), .Z(n2142) );
  CND2X2 U1936 ( .A(n2142), .B(n1893), .Z(n1331) );
  CND4X2 U1937 ( .A(n1334), .B(n1333), .C(n1332), .D(n1331), .Z(n1967) );
  CIVX2 U1938 ( .A(n1967), .Z(n2375) );
  CNR2X1 U1939 ( .A(n1632), .B(n1080), .Z(n1336) );
  CNR2X1 U1940 ( .A(n1180), .B(n1625), .Z(n1335) );
  CNR2X1 U1941 ( .A(n1336), .B(n1335), .Z(n1340) );
  CNR2X1 U1942 ( .A(n1633), .B(n1065), .Z(n1338) );
  CNR2X2 U1943 ( .A(n1338), .B(n1337), .Z(n1339) );
  CND2X2 U1944 ( .A(n1340), .B(n1339), .Z(n2370) );
  CND2X1 U1945 ( .A(n2370), .B(n2371), .Z(n1347) );
  CNR2X1 U1946 ( .A(n1547), .B(acc[55]), .Z(n1343) );
  CIVX2 U1947 ( .A(n1106), .Z(n1521) );
  CNR2X1 U1948 ( .A(acc[58]), .B(n1596), .Z(n1342) );
  CNR2X2 U1949 ( .A(n1343), .B(n1342), .Z(n2164) );
  CNR2X1 U1950 ( .A(n1632), .B(acc[57]), .Z(n1345) );
  CNR2X1 U1951 ( .A(n1345), .B(n1344), .Z(n2163) );
  CND2XL U1952 ( .A(n2164), .B(n2163), .Z(n1847) );
  CND2XL U1953 ( .A(n2369), .B(n2368), .Z(n1346) );
  CND2X1 U1954 ( .A(n1346), .B(n1347), .Z(n1968) );
  CND2X1 U1955 ( .A(n1196), .B(n1574), .Z(n1349) );
  CND2X1 U1956 ( .A(n1595), .B(n1163), .Z(n1348) );
  CND2X2 U1957 ( .A(n1349), .B(n1348), .Z(n1857) );
  CIVX2 U1958 ( .A(n1857), .Z(n1354) );
  CIVX2 U1959 ( .A(n1126), .Z(n2983) );
  CND2X1 U1960 ( .A(n1456), .B(n1350), .Z(n1351) );
  CND2X2 U1961 ( .A(n1352), .B(n1351), .Z(n1858) );
  CIVX2 U1962 ( .A(n1858), .Z(n1353) );
  CND2X2 U1963 ( .A(n1354), .B(n1353), .Z(n2372) );
  CND2X1 U1964 ( .A(n1196), .B(n1355), .Z(n1357) );
  CIVX2 U1965 ( .A(acc[53]), .Z(n2454) );
  CND2X1 U1966 ( .A(n1581), .B(n2454), .Z(n1356) );
  CND2X1 U1967 ( .A(n1359), .B(n1358), .Z(n1696) );
  CIVXL U1968 ( .A(n1696), .Z(n1360) );
  CND2IX1 U1969 ( .B(n1697), .A(n1360), .Z(n2168) );
  CND2X1 U1970 ( .A(n2129), .B(n2344), .Z(n2177) );
  CANR2X1 U1971 ( .A(n2582), .B(n2375), .C(n1363), .D(n1362), .Z(n1411) );
  CND2XL U1972 ( .A(n1638), .B(acc[28]), .Z(n1368) );
  CIVX2 U1973 ( .A(n1624), .Z(n1643) );
  CND2X1 U1974 ( .A(n1643), .B(n1140), .Z(n1367) );
  CIVX1 U1975 ( .A(acc[27]), .Z(n3495) );
  COR2X1 U1976 ( .A(n3495), .B(n1477), .Z(n1366) );
  COR2X1 U1977 ( .A(n1364), .B(n1446), .Z(n1365) );
  CND4X2 U1978 ( .A(n1368), .B(n1367), .C(n1366), .D(n1365), .Z(n2138) );
  CAN2X1 U1979 ( .A(n1961), .B(n2268), .Z(n1385) );
  CIVX2 U1980 ( .A(n1625), .Z(n1517) );
  CND2X1 U1981 ( .A(n1643), .B(acc[17]), .Z(n1372) );
  CNR2X1 U1982 ( .A(n1370), .B(n1369), .Z(n1371) );
  CND3X2 U1983 ( .A(n1373), .B(n1372), .C(n1371), .Z(n2154) );
  CND2X1 U1984 ( .A(n2154), .B(n2176), .Z(n1960) );
  CND2X1 U1985 ( .A(n1196), .B(acc[24]), .Z(n1374) );
  CIVX2 U1986 ( .A(n1374), .Z(n1376) );
  CIVX1 U1987 ( .A(acc[23]), .Z(n1618) );
  CNR2X1 U1988 ( .A(n1618), .B(n1547), .Z(n1375) );
  CNR2X2 U1989 ( .A(n1376), .B(n1375), .Z(n1381) );
  CNR2X1 U1990 ( .A(n3136), .B(n1634), .Z(n1379) );
  CND2X1 U1991 ( .A(n1648), .B(acc[25]), .Z(n1377) );
  CIVX2 U1992 ( .A(n1377), .Z(n1378) );
  CNR2X2 U1993 ( .A(n1379), .B(n1378), .Z(n1380) );
  CND2X1 U1994 ( .A(n1149), .B(n1893), .Z(n1959) );
  CND2X1 U1995 ( .A(n1484), .B(acc[22]), .Z(n1383) );
  CND2XL U1996 ( .A(n1553), .B(acc[19]), .Z(n1382) );
  CIVX1 U1997 ( .A(acc[21]), .Z(n1384) );
  CIVX1 U1998 ( .A(acc[20]), .Z(n1616) );
  CND2IX1 U1999 ( .B(n1838), .A(n1836), .Z(n2145) );
  CIVX2 U2000 ( .A(n2172), .Z(n1922) );
  CND4X1 U2001 ( .A(n1385), .B(n1960), .C(n1959), .D(n1962), .Z(n1409) );
  CIVXL U2002 ( .A(n1485), .Z(n1580) );
  CND2X1 U2003 ( .A(n1580), .B(acc[63]), .Z(n2173) );
  CIVX2 U2004 ( .A(n2173), .Z(n1963) );
  CND2X1 U2005 ( .A(n2121), .B(n1958), .Z(n2336) );
  CIVX2 U2006 ( .A(n2336), .Z(n2349) );
  CND4X1 U2007 ( .A(n1963), .B(n2161), .C(h2[6]), .D(n2349), .Z(n1390) );
  CNR2X1 U2008 ( .A(h2[5]), .B(h2[6]), .Z(n2153) );
  CIVX2 U2009 ( .A(n2153), .Z(n2763) );
  CND2X1 U2010 ( .A(n1390), .B(n2763), .Z(n1408) );
  CND2X1 U2011 ( .A(n1198), .B(acc[6]), .Z(n1389) );
  CND2X1 U2012 ( .A(n1643), .B(acc[5]), .Z(n1388) );
  CND2XL U2013 ( .A(n1638), .B(acc[4]), .Z(n1387) );
  CND4X1 U2014 ( .A(n1389), .B(n1388), .C(n1387), .D(n1386), .Z(n1681) );
  CIVXL U2015 ( .A(acc[7]), .Z(n3473) );
  CIVXL U2016 ( .A(acc[10]), .Z(n1391) );
  CND2X1 U2017 ( .A(n1643), .B(acc[9]), .Z(n1393) );
  CND3X1 U2018 ( .A(n1394), .B(n1393), .C(n1392), .Z(n1839) );
  CND2XL U2019 ( .A(n1395), .B(acc[2]), .Z(n1399) );
  CND2XL U2020 ( .A(n1196), .B(acc[0]), .Z(n1398) );
  CND2X1 U2021 ( .A(n1643), .B(acc[1]), .Z(n1397) );
  CANR11X1 U2022 ( .A(n1399), .B(n1398), .C(n1397), .D(n1396), .Z(n1400) );
  CANR1XL U2023 ( .A(n1893), .B(n1839), .C(n1400), .Z(n1405) );
  CND2X1 U2024 ( .A(n1615), .B(acc[13]), .Z(n1402) );
  CNR2X1 U2025 ( .A(n1841), .B(n1840), .Z(n1685) );
  CIVX2 U2026 ( .A(n1685), .Z(n2152) );
  CND2X1 U2027 ( .A(n2152), .B(n2371), .Z(n1404) );
  CND3XL U2028 ( .A(n1406), .B(n1405), .C(n1404), .Z(n1407) );
  CND3X1 U2029 ( .A(n1409), .B(n1408), .C(n1407), .Z(n1410) );
  CND2X2 U2030 ( .A(n1411), .B(n1410), .Z(n2028) );
  CIVXL U2031 ( .A(n2086), .Z(n1466) );
  CNR2X1 U2032 ( .A(n1477), .B(n3073), .Z(n1413) );
  CNR2X1 U2033 ( .A(n1413), .B(n1412), .Z(n1416) );
  CIVX3 U2034 ( .A(n1414), .Z(n1588) );
  CND2X1 U2035 ( .A(n1588), .B(acc[39]), .Z(n1415) );
  CNR2XL U2036 ( .A(n1477), .B(n2696), .Z(n1419) );
  CIVX1 U2037 ( .A(acc[36]), .Z(n2961) );
  CNR2X1 U2038 ( .A(n2961), .B(n1446), .Z(n1418) );
  CNR2X1 U2039 ( .A(n1419), .B(n1418), .Z(n1422) );
  CND2X1 U2040 ( .A(n1503), .B(acc[34]), .Z(n1421) );
  CND2X1 U2041 ( .A(n1615), .B(acc[35]), .Z(n1420) );
  CND3X2 U2042 ( .A(n1422), .B(n1421), .C(n1420), .Z(n2098) );
  CIVX2 U2043 ( .A(n2098), .Z(n1423) );
  CND2X2 U2044 ( .A(n1423), .B(n2176), .Z(n1424) );
  CNR2X1 U2045 ( .A(n1632), .B(acc[47]), .Z(n1427) );
  CNR2XL U2046 ( .A(n1625), .B(acc[46]), .Z(n1426) );
  CNR2X1 U2047 ( .A(n1427), .B(n1426), .Z(n1431) );
  CNR2X1 U2048 ( .A(acc[48]), .B(n1555), .Z(n1429) );
  CNR2X1 U2049 ( .A(n1477), .B(n858), .Z(n1428) );
  CNR2X2 U2050 ( .A(n1429), .B(n1428), .Z(n1430) );
  CND2X2 U2051 ( .A(n1431), .B(n1430), .Z(n2126) );
  CIVXL U2052 ( .A(n2126), .Z(n1439) );
  CIVDX1 U2053 ( .A(n1521), .Z0(n1548), .Z1(n1484) );
  CNR2X1 U2054 ( .A(acc[44]), .B(n1548), .Z(n1433) );
  CNR2X2 U2055 ( .A(n1135), .B(n1433), .Z(n1437) );
  CND2X1 U2056 ( .A(n1588), .B(n1434), .Z(n1436) );
  CND2X1 U2057 ( .A(n1503), .B(n1073), .Z(n1435) );
  COND1X1 U2058 ( .A(n2087), .B(n1439), .C(n1438), .Z(n1440) );
  CNR2X2 U2059 ( .A(n1441), .B(n1440), .Z(n2392) );
  CNR2X1 U2060 ( .A(n1632), .B(n3495), .Z(n1443) );
  CNR2XL U2061 ( .A(n1625), .B(n3136), .Z(n1442) );
  CNR2X1 U2062 ( .A(n1442), .B(n1443), .Z(n2115) );
  CND2X1 U2063 ( .A(n1455), .B(acc[28]), .Z(n1445) );
  CND2XL U2064 ( .A(n1509), .B(acc[25]), .Z(n1444) );
  CIVX2 U2065 ( .A(n1935), .Z(n2114) );
  CND2X2 U2066 ( .A(n2115), .B(n2114), .Z(n1776) );
  CND2IX1 U2067 ( .B(n1223), .A(n1776), .Z(n1452) );
  CND2X1 U2068 ( .A(n1503), .B(acc[30]), .Z(n1450) );
  CIVX2 U2069 ( .A(acc[32]), .Z(n1546) );
  COR2X1 U2070 ( .A(n1546), .B(n1611), .Z(n1449) );
  CND2X1 U2071 ( .A(n1588), .B(acc[31]), .Z(n1448) );
  CIVX2 U2072 ( .A(n2064), .Z(n2034) );
  CND2X1 U2073 ( .A(n1588), .B(acc[23]), .Z(n1454) );
  CND2X1 U2074 ( .A(n1638), .B(acc[22]), .Z(n1453) );
  CND2X2 U2075 ( .A(n1454), .B(n1453), .Z(n1936) );
  CND2X1 U2076 ( .A(n1455), .B(acc[24]), .Z(n1458) );
  CND2X1 U2077 ( .A(n1458), .B(n1457), .Z(n1937) );
  CIVXL U2078 ( .A(n2110), .Z(n1464) );
  CND2X1 U2079 ( .A(n1198), .B(acc[20]), .Z(n1463) );
  CND2X1 U2080 ( .A(n1595), .B(acc[19]), .Z(n1462) );
  CIVXL U2081 ( .A(n1459), .Z(n1539) );
  CND2X1 U2082 ( .A(n1539), .B(acc[17]), .Z(n1460) );
  CND4X1 U2083 ( .A(n1463), .B(n1462), .C(n1461), .D(n1460), .Z(n2117) );
  COND1X1 U2084 ( .A(n1466), .B(n2392), .C(n1465), .Z(n1532) );
  CNR2X1 U2085 ( .A(n1547), .B(acc[53]), .Z(n1468) );
  CNR2X1 U2086 ( .A(n1108), .B(n1548), .Z(n1467) );
  CNR2X2 U2087 ( .A(n1468), .B(n1467), .Z(n1472) );
  CND2X1 U2088 ( .A(n1559), .B(n1469), .Z(n1471) );
  CND2X1 U2089 ( .A(n1503), .B(n1089), .Z(n1470) );
  CND2XL U2090 ( .A(n2124), .B(n2122), .Z(n1483) );
  CND2X1 U2091 ( .A(n1581), .B(n1473), .Z(n1474) );
  CIVX2 U2092 ( .A(n1476), .Z(n1481) );
  CNR2X1 U2093 ( .A(n1477), .B(n1162), .Z(n1478) );
  CNR2X2 U2094 ( .A(n1478), .B(n1479), .Z(n1480) );
  CND2X1 U2095 ( .A(n2123), .B(n2099), .Z(n1482) );
  CND2X1 U2096 ( .A(n1483), .B(n1482), .Z(n1500) );
  CND2X1 U2097 ( .A(n1588), .B(n1066), .Z(n1489) );
  CIVX1 U2098 ( .A(acc[58]), .Z(n2740) );
  CND2X1 U2099 ( .A(n1503), .B(n2740), .Z(n1488) );
  CND2X1 U2100 ( .A(n1484), .B(n1181), .Z(n1487) );
  CIVXL U2101 ( .A(n1485), .Z(n1639) );
  CIVX1 U2102 ( .A(acc[57]), .Z(n2951) );
  CND2X1 U2103 ( .A(n1639), .B(n2951), .Z(n1486) );
  CND4X1 U2104 ( .A(n1486), .B(n1488), .C(n1487), .D(n1489), .Z(n2127) );
  CND2X1 U2105 ( .A(n2127), .B(n1893), .Z(n1498) );
  CNR2XL U2106 ( .A(n1490), .B(acc[62]), .Z(n1491) );
  CND2IX1 U2107 ( .B(n1491), .A(n1596), .Z(n1492) );
  CIVX2 U2108 ( .A(n1492), .Z(n1496) );
  CND2XL U2109 ( .A(n1575), .B(n1081), .Z(n1495) );
  CNR2XL U2110 ( .A(n1098), .B(acc[63]), .Z(n1493) );
  CIVX1 U2111 ( .A(n1493), .Z(n1494) );
  CND3X2 U2112 ( .A(n1496), .B(n1495), .C(n1494), .Z(n2218) );
  CND2XL U2113 ( .A(n2218), .B(n2371), .Z(n1497) );
  CND2X1 U2114 ( .A(n1498), .B(n1497), .Z(n1499) );
  CNR2X2 U2115 ( .A(n1500), .B(n1499), .Z(n2403) );
  CNR2IX1 U2116 ( .B(n2018), .A(n2155), .Z(n1501) );
  CND2X1 U2117 ( .A(n1395), .B(acc[8]), .Z(n1507) );
  CND2X1 U2118 ( .A(n1643), .B(acc[7]), .Z(n1506) );
  CND2XL U2119 ( .A(n1503), .B(acc[6]), .Z(n1505) );
  CND2X1 U2120 ( .A(n1639), .B(acc[5]), .Z(n1504) );
  CND4X1 U2121 ( .A(n1507), .B(n1506), .C(n1505), .D(n1504), .Z(n2067) );
  CND2X1 U2122 ( .A(n1643), .B(acc[11]), .Z(n1512) );
  CND2XL U2123 ( .A(n1509), .B(acc[9]), .Z(n1510) );
  CND4X1 U2124 ( .A(n1513), .B(n1512), .C(n1511), .D(n1510), .Z(n2072) );
  CIVX2 U2125 ( .A(n1194), .Z(n1820) );
  COND2X1 U2126 ( .A(n2073), .B(n2067), .C(n2072), .D(n1820), .Z(n1529) );
  COND2XL U2127 ( .A(n1555), .B(acc[4]), .C(acc[1]), .D(n1633), .Z(n1515) );
  COND2XL U2128 ( .A(acc[3]), .B(n1632), .C(acc[2]), .D(n1625), .Z(n1514) );
  CNR2X1 U2129 ( .A(n1515), .B(n1514), .Z(n1516) );
  COAN1X1 U2130 ( .A(n1680), .B(n1516), .C(n2337), .Z(n1527) );
  CND2X1 U2131 ( .A(n1517), .B(acc[14]), .Z(n1519) );
  CND2X1 U2132 ( .A(n1520), .B(acc[13]), .Z(n1523) );
  CND2X1 U2133 ( .A(n1484), .B(acc[16]), .Z(n1522) );
  CND2X1 U2134 ( .A(n1523), .B(n1522), .Z(n1524) );
  CNR2X2 U2135 ( .A(n1525), .B(n1524), .Z(n2109) );
  CND2X1 U2136 ( .A(n2113), .B(n2018), .Z(n1647) );
  CND2X1 U2137 ( .A(n2109), .B(n2059), .Z(n1526) );
  CND2X1 U2138 ( .A(n1527), .B(n1526), .Z(n1528) );
  CNR2X1 U2139 ( .A(n1529), .B(n1528), .Z(n1530) );
  COND1X1 U2140 ( .A(n1758), .B(n2403), .C(n1530), .Z(n1531) );
  CNR2X2 U2141 ( .A(n1532), .B(n1531), .Z(n2135) );
  CAN2X1 U2142 ( .A(n1575), .B(n3632), .Z(n1534) );
  CNR2X1 U2143 ( .A(n1596), .B(acc[47]), .Z(n1533) );
  CNR2X2 U2144 ( .A(n1534), .B(n1533), .Z(n1538) );
  CND2X1 U2145 ( .A(n1595), .B(n1535), .Z(n1536) );
  CND3X2 U2146 ( .A(n1538), .B(n1537), .C(n1536), .Z(n1894) );
  CND2X1 U2147 ( .A(n1894), .B(n2371), .Z(n1543) );
  CND2IXL U2148 ( .B(n1434), .A(n1395), .Z(n1541) );
  CND2X1 U2149 ( .A(n1539), .B(n1166), .Z(n1540) );
  CND2X1 U2150 ( .A(n1541), .B(n1540), .Z(n1810) );
  COND2X1 U2151 ( .A(n1625), .B(n1432), .C(n1073), .D(n1558), .Z(n1811) );
  CNR2X1 U2152 ( .A(n1811), .B(n1810), .Z(n1891) );
  CND2X2 U2153 ( .A(n1543), .B(n1542), .Z(n1565) );
  CIVDX1 U2154 ( .A(n1695), .Z0(n1563), .Z1(n2125) );
  CAN2XL U2155 ( .A(n1544), .B(acc[33]), .Z(n1545) );
  CANR1XL U2156 ( .A(acc[34]), .B(n1615), .C(n1545), .Z(n1552) );
  CIVXL U2157 ( .A(acc[35]), .Z(n1549) );
  COR2X1 U2158 ( .A(n1549), .B(n1548), .Z(n1550) );
  CND3X1 U2159 ( .A(n1552), .B(n1551), .C(n1550), .Z(n1895) );
  CND2X1 U2160 ( .A(n1638), .B(acc[37]), .Z(n1752) );
  CAN2XL U2161 ( .A(n1553), .B(acc[36]), .Z(n1557) );
  CNR2X2 U2162 ( .A(n1557), .B(n1556), .Z(n1753) );
  CIVXL U2163 ( .A(acc[38]), .Z(n1560) );
  CIVXL U2164 ( .A(n1414), .Z(n1559) );
  CND2IX1 U2165 ( .B(n1560), .A(n1588), .Z(n1751) );
  COND2X1 U2166 ( .A(n1895), .B(n1563), .C(n1562), .D(n1561), .Z(n1564) );
  CNR2X2 U2167 ( .A(n1565), .B(n1564), .Z(n2365) );
  CNR2IX1 U2168 ( .B(n2086), .A(n2365), .Z(n1566) );
  CIVX2 U2169 ( .A(n1566), .Z(n1594) );
  CND2XL U2170 ( .A(n1567), .B(n1081), .Z(n1569) );
  CND2X1 U2171 ( .A(n1581), .B(n3630), .Z(n1568) );
  CND2X1 U2172 ( .A(n1572), .B(n1571), .Z(n1755) );
  CNR2X2 U2173 ( .A(n1756), .B(n1755), .Z(n2088) );
  CNR2X1 U2174 ( .A(n2088), .B(n2087), .Z(n1573) );
  CIVX2 U2175 ( .A(n1573), .Z(n2407) );
  CND2X1 U2176 ( .A(n1575), .B(n1574), .Z(n1576) );
  COND1X1 U2177 ( .A(acc[51]), .B(n1577), .C(n1576), .Z(n1578) );
  CND2X1 U2178 ( .A(n1892), .B(n2161), .Z(n2406) );
  CND2X1 U2179 ( .A(n1196), .B(n2951), .Z(n1584) );
  CND2IX1 U2180 ( .B(n1108), .A(n1580), .Z(n1583) );
  CND2X1 U2181 ( .A(n1581), .B(n2740), .Z(n1582) );
  CND4X2 U2182 ( .A(n1585), .B(n1584), .C(n1583), .D(n1582), .Z(n1878) );
  CND2X1 U2183 ( .A(n1878), .B(n2368), .Z(n2405) );
  CNR2X1 U2184 ( .A(n1633), .B(acc[52]), .Z(n1587) );
  CNR2X1 U2185 ( .A(acc[55]), .B(n1446), .Z(n1586) );
  CNR2X2 U2186 ( .A(n1587), .B(n1586), .Z(n1591) );
  CND2XL U2187 ( .A(n1196), .B(n2454), .Z(n1590) );
  CND2X1 U2188 ( .A(n1588), .B(n1089), .Z(n1589) );
  CND3X2 U2189 ( .A(n1591), .B(n1590), .C(n1589), .Z(n1877) );
  CND2X1 U2190 ( .A(n1877), .B(n1922), .Z(n2404) );
  CND2XL U2191 ( .A(n1638), .B(acc[25]), .Z(n1602) );
  CND2X1 U2192 ( .A(n709), .B(acc[26]), .Z(n1601) );
  CNR2X1 U2193 ( .A(n3495), .B(n1596), .Z(n1599) );
  CIVX1 U2194 ( .A(acc[24]), .Z(n1597) );
  CNR2X1 U2195 ( .A(n1599), .B(n1598), .Z(n1600) );
  CND3X1 U2196 ( .A(n1601), .B(n1602), .C(n1600), .Z(n1981) );
  CIVX2 U2197 ( .A(acc[31]), .Z(n3054) );
  CNR2X1 U2198 ( .A(n1604), .B(n1603), .Z(n1607) );
  CND2XL U2199 ( .A(n1638), .B(n1140), .Z(n1606) );
  CND2X1 U2200 ( .A(n1615), .B(acc[30]), .Z(n1605) );
  CND2X1 U2201 ( .A(n1899), .B(n2371), .Z(n1608) );
  CND2X1 U2202 ( .A(n1609), .B(n1608), .Z(n1946) );
  CIVX1 U2203 ( .A(acc[16]), .Z(n3506) );
  CND2X1 U2204 ( .A(n1503), .B(acc[17]), .Z(n1610) );
  CND2X2 U2205 ( .A(n1206), .B(n1610), .Z(n1614) );
  CIVX1 U2206 ( .A(acc[19]), .Z(n2734) );
  CND2X1 U2207 ( .A(n1648), .B(acc[18]), .Z(n1612) );
  CIVX2 U2208 ( .A(n1067), .Z(n1819) );
  CND2X1 U2209 ( .A(n1819), .B(n2176), .Z(n1945) );
  CND2XL U2210 ( .A(n1638), .B(acc[21]), .Z(n1623) );
  CND2X1 U2211 ( .A(n1615), .B(acc[22]), .Z(n1622) );
  CNR2X1 U2212 ( .A(n1617), .B(n1616), .Z(n1620) );
  CNR2X1 U2213 ( .A(n1618), .B(n1611), .Z(n1619) );
  CNR2X1 U2214 ( .A(n1620), .B(n1619), .Z(n1621) );
  CND3XL U2215 ( .A(n1945), .B(n1944), .C(n2034), .Z(n1667) );
  CNR2IXL U2216 ( .B(acc[10]), .A(n1558), .Z(n1627) );
  CNR2IX1 U2217 ( .B(acc[9]), .A(n1625), .Z(n1626) );
  CNR2XL U2218 ( .A(n1627), .B(n1626), .Z(n1631) );
  CND2X1 U2219 ( .A(n1395), .B(acc[11]), .Z(n1628) );
  CND2X2 U2220 ( .A(n1631), .B(n1630), .Z(n1821) );
  CIVX2 U2221 ( .A(n1821), .Z(n2036) );
  CND2X1 U2222 ( .A(n2036), .B(n1194), .Z(n1646) );
  COND2XL U2223 ( .A(acc[2]), .B(n1632), .C(acc[1]), .D(n1625), .Z(n1636) );
  CND2IX1 U2224 ( .B(n1636), .A(n1635), .Z(n1637) );
  CANR1X2 U2225 ( .A(n2050), .B(n1637), .C(h2[6]), .Z(n1645) );
  CND2X1 U2226 ( .A(n1638), .B(acc[5]), .Z(n1642) );
  CND2X1 U2227 ( .A(n1639), .B(acc[4]), .Z(n1641) );
  CND2XL U2228 ( .A(n1521), .B(acc[7]), .Z(n1640) );
  CAN3X1 U2229 ( .A(n1642), .B(n1641), .C(n1640), .Z(n2042) );
  CND2X1 U2230 ( .A(n1643), .B(acc[6]), .Z(n2041) );
  CND4X1 U2231 ( .A(n2042), .B(n2007), .C(n2041), .D(n2018), .Z(n1644) );
  CIVDX1 U2232 ( .A(n1647), .Z0(n2059), .Z1(n2069) );
  CND2XL U2233 ( .A(n1567), .B(acc[13]), .Z(n1652) );
  CND2XL U2234 ( .A(n1649), .B(acc[12]), .Z(n1651) );
  CND2X1 U2235 ( .A(n1197), .B(acc[15]), .Z(n1650) );
  CND3X1 U2236 ( .A(n1652), .B(n1651), .C(n1650), .Z(n1653) );
  CIVX2 U2237 ( .A(n2037), .Z(n1818) );
  COND1XL U2238 ( .A(n1946), .B(n1667), .C(n1666), .Z(n1655) );
  CNR2X1 U2239 ( .A(n1669), .B(n1655), .Z(n1656) );
  CND3X1 U2240 ( .A(n1656), .B(n2028), .C(n2135), .Z(n2669) );
  CIVXL U2241 ( .A(push_2), .Z(n1657) );
  CNR2X1 U2242 ( .A(n1657), .B(cmd_2[1]), .Z(n2495) );
  CIVXL U2243 ( .A(n2495), .Z(n1658) );
  CANR2XL U2244 ( .A(n1659), .B(mulout[2]), .C(acc[2]), .D(n3617), .Z(n1663)
         );
  CNR2X1 U2245 ( .A(acc[2]), .B(mulout[2]), .Z(n2222) );
  CND2X1 U2246 ( .A(acc[2]), .B(mulout[2]), .Z(n2225) );
  CND2X1 U2247 ( .A(acc[0]), .B(mulout[0]), .Z(n1674) );
  CNR2X1 U2248 ( .A(acc[1]), .B(mulout[1]), .Z(n1670) );
  CND2X1 U2249 ( .A(acc[1]), .B(mulout[1]), .Z(n1671) );
  COND1X1 U2250 ( .A(n1674), .B(n1670), .C(n1671), .Z(n2228) );
  CIVX1 U2251 ( .A(n2228), .Z(n1703) );
  CEOXL U2252 ( .A(n1660), .B(n1703), .Z(n1661) );
  CAN2X2 U2253 ( .A(n2495), .B(cmd_2[0]), .Z(n3595) );
  CND2XL U2254 ( .A(n1661), .B(n3595), .Z(n1662) );
  COND3X1 U2255 ( .A(n1664), .B(n3325), .C(n1663), .D(n1662), .Z(n1665) );
  CIVX2 U2256 ( .A(n1665), .Z(n3626) );
  COND1X1 U2257 ( .A(n1946), .B(n1667), .C(n1666), .Z(n1668) );
  CNR2X2 U2258 ( .A(n1669), .B(n1668), .Z(n2181) );
  CND2XL U2259 ( .A(n2181), .B(n2028), .Z(n1673) );
  CIVXL U2260 ( .A(push_2), .Z(n3617) );
  CND2X1 U2261 ( .A(n2136), .B(n2371), .Z(n1677) );
  CND2IX1 U2262 ( .B(n1675), .A(n2145), .Z(n1676) );
  CIVX2 U2263 ( .A(n2148), .Z(n1679) );
  COND1X2 U2264 ( .A(n2172), .B(n1679), .C(n1678), .Z(n1885) );
  CNR2XL U2265 ( .A(n1887), .B(n1885), .Z(n1690) );
  CNR2X1 U2266 ( .A(n1839), .B(n2073), .Z(n1683) );
  CIVDX1 U2267 ( .A(n1680), .Z0(n2050), .Z1(n2068) );
  CNR2X1 U2268 ( .A(n2068), .B(n1681), .Z(n1682) );
  CNR2X2 U2269 ( .A(n1683), .B(n1682), .Z(n1688) );
  CIVX2 U2270 ( .A(n2154), .Z(n1684) );
  CANR1X2 U2271 ( .A(n2059), .B(n1684), .C(h2[6]), .Z(n1687) );
  CND2X1 U2272 ( .A(n1685), .B(n1194), .Z(n1686) );
  CND3X2 U2273 ( .A(n1688), .B(n1687), .C(n1686), .Z(n1689) );
  CANR1X2 U2274 ( .A(n2034), .B(n1690), .C(n1689), .Z(n2095) );
  CND2X2 U2275 ( .A(n2142), .B(n2169), .Z(n1692) );
  CND2X2 U2276 ( .A(n2140), .B(n2176), .Z(n1691) );
  CND2X2 U2277 ( .A(n1692), .B(n1691), .Z(n1882) );
  CND2X2 U2278 ( .A(n2372), .B(n2371), .Z(n1693) );
  CND2X2 U2279 ( .A(n1694), .B(n1693), .Z(n1883) );
  COND1X1 U2280 ( .A(n1882), .B(n1883), .C(n2086), .Z(n1702) );
  CIVDX1 U2281 ( .A(n1695), .Z0(n2706), .Z1(n2099) );
  CNR2X1 U2282 ( .A(n1697), .B(n1696), .Z(n1864) );
  CND2X1 U2283 ( .A(n2370), .B(n2368), .Z(n1700) );
  CND2X1 U2284 ( .A(n2164), .B(n2163), .Z(n2369) );
  CND2X2 U2285 ( .A(n1700), .B(n1699), .Z(n1874) );
  COND1XL U2286 ( .A(n1876), .B(n1874), .C(n2090), .Z(n1701) );
  CIVX2 U2287 ( .A(n2669), .Z(n2823) );
  CIVX2 U2288 ( .A(n2820), .Z(n2290) );
  COND1XL U2289 ( .A(n2222), .B(n1703), .C(n2225), .Z(n1705) );
  CNR2X1 U2290 ( .A(acc[3]), .B(mulout[3]), .Z(n2224) );
  CND2X1 U2291 ( .A(acc[3]), .B(mulout[3]), .Z(n2223) );
  CMX2XL U2292 ( .A0(n710), .A1(q[1]), .S(pushin), .Z(n1707) );
  CMX2XL U2293 ( .A0(n1094), .A1(q[3]), .S(n3624), .Z(n1708) );
  CMX2XL U2294 ( .A0(q0[5]), .A1(q[5]), .S(n3624), .Z(n1709) );
  CMX2XL U2295 ( .A0(q0[11]), .A1(q[11]), .S(pushin), .Z(n1710) );
  CMX2XL U2296 ( .A0(q0[17]), .A1(q[17]), .S(n3624), .Z(n1711) );
  CMX2XL U2297 ( .A0(q0[20]), .A1(q[20]), .S(pushin), .Z(n1712) );
  CMX2XL U2298 ( .A0(q0[21]), .A1(q[21]), .S(n3624), .Z(n1713) );
  CMX2XL U2299 ( .A0(q0[22]), .A1(q[22]), .S(pushin), .Z(n1714) );
  CMX2XL U2300 ( .A0(q0[31]), .A1(q[31]), .S(n3624), .Z(n1715) );
  CMX2XL U2301 ( .A0(q0[24]), .A1(q[24]), .S(n3624), .Z(n1716) );
  CMX2XL U2302 ( .A0(n1077), .A1(q[25]), .S(n3624), .Z(n1717) );
  CMX2XL U2303 ( .A0(q0[23]), .A1(q[23]), .S(pushin), .Z(n1718) );
  CMX2XL U2304 ( .A0(q0[30]), .A1(q[30]), .S(n3624), .Z(n1719) );
  CMX2XL U2305 ( .A0(q0[27]), .A1(q[27]), .S(n3624), .Z(n1720) );
  CMX2XL U2306 ( .A0(h0[7]), .A1(h[7]), .S(n3624), .Z(n1721) );
  CMX2XL U2307 ( .A0(h0[8]), .A1(h[8]), .S(n3624), .Z(n1722) );
  CMX2XL U2308 ( .A0(h0[9]), .A1(h[9]), .S(n3624), .Z(n1723) );
  CMX2XL U2309 ( .A0(h0[10]), .A1(h[10]), .S(n3624), .Z(n1724) );
  CMX2XL U2310 ( .A0(h0[11]), .A1(h[11]), .S(n3624), .Z(n1725) );
  CMX2XL U2311 ( .A0(h0[12]), .A1(h[12]), .S(n3624), .Z(n1726) );
  CMX2XL U2312 ( .A0(h0[13]), .A1(h[13]), .S(n3624), .Z(n1727) );
  CMX2XL U2313 ( .A0(h0[14]), .A1(h[14]), .S(n3624), .Z(n1728) );
  CMX2XL U2314 ( .A0(h0[15]), .A1(h[15]), .S(n3624), .Z(n1729) );
  CMX2XL U2315 ( .A0(h0[16]), .A1(h[16]), .S(n3624), .Z(n1730) );
  CMX2XL U2316 ( .A0(h0[17]), .A1(h[17]), .S(n3624), .Z(n1731) );
  CMX2XL U2317 ( .A0(h0[18]), .A1(h[18]), .S(n3624), .Z(n1732) );
  CMX2XL U2318 ( .A0(h0[19]), .A1(h[19]), .S(n3624), .Z(n1733) );
  CMX2XL U2319 ( .A0(h0[20]), .A1(h[20]), .S(n3624), .Z(n1734) );
  CMX2XL U2320 ( .A0(h0[21]), .A1(h[21]), .S(n3624), .Z(n1735) );
  CMX2XL U2321 ( .A0(h0[22]), .A1(h[22]), .S(n3624), .Z(n1736) );
  CMX2XL U2322 ( .A0(h0[23]), .A1(h[23]), .S(n3624), .Z(n1737) );
  CMX2XL U2323 ( .A0(h0[24]), .A1(h[24]), .S(pushin), .Z(n1738) );
  CMX2XL U2324 ( .A0(h0[25]), .A1(h[25]), .S(pushin), .Z(n1739) );
  CMX2XL U2325 ( .A0(h0[26]), .A1(h[26]), .S(pushin), .Z(n1740) );
  CMX2XL U2326 ( .A0(h0[27]), .A1(h[27]), .S(pushin), .Z(n1741) );
  CMX2XL U2327 ( .A0(h0[28]), .A1(h[28]), .S(pushin), .Z(n1742) );
  CMX2XL U2328 ( .A0(h0[29]), .A1(h[29]), .S(pushin), .Z(n1743) );
  CMX2XL U2329 ( .A0(h0[30]), .A1(h[30]), .S(pushin), .Z(n1744) );
  CMX2XL U2330 ( .A0(h0[31]), .A1(h[31]), .S(pushin), .Z(n1745) );
  CMX2XL U2331 ( .A0(q0[28]), .A1(q[28]), .S(n3624), .Z(n1746) );
  CMX2XL U2332 ( .A0(q0[0]), .A1(q[0]), .S(pushin), .Z(n1747) );
  CMX2XL U2333 ( .A0(n708), .A1(q[13]), .S(pushin), .Z(n1748) );
  CMX2XL U2334 ( .A0(q0[19]), .A1(q[19]), .S(n3624), .Z(n1749) );
  CND3XL U2335 ( .A(cmd_2[0]), .B(cmd_2[1]), .C(push_2), .Z(n3435) );
  CMX2XL U2336 ( .A0(q0[15]), .A1(q[15]), .S(n3624), .Z(n1750) );
  CIVX2 U2337 ( .A(n1979), .Z(n1754) );
  CND3X2 U2338 ( .A(n1753), .B(n1752), .C(n1751), .Z(n1889) );
  CND2XL U2339 ( .A(n1889), .B(n2368), .Z(n1980) );
  CND2XL U2340 ( .A(n1895), .B(n2169), .Z(n1977) );
  CND4X1 U2341 ( .A(n1754), .B(n2349), .C(n1980), .D(n1977), .Z(n1768) );
  CND2X4 U2342 ( .A(n1758), .B(n2337), .Z(n2507) );
  CANR1X1 U2343 ( .A(h2[5]), .B(n2312), .C(n2507), .Z(n2351) );
  COND1XL U2344 ( .A(n1916), .B(n2707), .C(n2351), .Z(n1762) );
  CND2XL U2345 ( .A(n1892), .B(n2014), .Z(n1759) );
  CND2X1 U2346 ( .A(n1759), .B(n1760), .Z(n1991) );
  CIVX2 U2347 ( .A(n1763), .Z(n1767) );
  CND2XL U2348 ( .A(n1877), .B(n2368), .Z(n1764) );
  CND2X1 U2349 ( .A(n1765), .B(n1764), .Z(n1992) );
  CND2X1 U2350 ( .A(n1992), .B(n2344), .Z(n1766) );
  CND2XL U2351 ( .A(n2124), .B(n2371), .Z(n1770) );
  CND2X1 U2352 ( .A(n1770), .B(n1769), .Z(n1771) );
  CIVX2 U2353 ( .A(n1771), .Z(n1775) );
  CND2X1 U2354 ( .A(n2126), .B(n2169), .Z(n1773) );
  CND2X2 U2355 ( .A(n1775), .B(n1774), .Z(n2335) );
  CND2X2 U2356 ( .A(n2335), .B(n2086), .Z(n1787) );
  CND2XL U2357 ( .A(n2100), .B(n1922), .Z(n2203) );
  CND2XL U2358 ( .A(n2103), .B(n2371), .Z(n2202) );
  CND3XL U2359 ( .A(n2204), .B(n2202), .C(n2203), .Z(n1777) );
  CIVXL U2360 ( .A(n1777), .Z(n1778) );
  CND2XL U2361 ( .A(n2098), .B(n1893), .Z(n2201) );
  CND3XL U2362 ( .A(n1778), .B(n2034), .C(n2201), .Z(n1786) );
  CIVXL U2363 ( .A(n2127), .Z(n1781) );
  CIVX2 U2364 ( .A(n2218), .Z(n2708) );
  CND2X1 U2365 ( .A(n2708), .B(n2122), .Z(n1779) );
  CIVX1 U2366 ( .A(n1779), .Z(n1780) );
  CANR1X1 U2367 ( .A(n1781), .B(n2125), .C(n1780), .Z(n2339) );
  COND1XL U2368 ( .A(n2072), .B(n2068), .C(n2337), .Z(n1782) );
  CIVXL U2369 ( .A(n2146), .Z(n2003) );
  CIVXL U2370 ( .A(n2109), .Z(n1783) );
  CND4X1 U2371 ( .A(n1787), .B(n1786), .C(n1784), .D(n1785), .Z(n2607) );
  CND2X1 U2372 ( .A(n2013), .B(n2169), .Z(n1791) );
  CND2X1 U2373 ( .A(n2000), .B(n2161), .Z(n1790) );
  CIVX1 U2374 ( .A(n2113), .Z(n2147) );
  CND2XL U2375 ( .A(n2058), .B(n2146), .Z(n1793) );
  CND3X2 U2376 ( .A(n1794), .B(n1793), .C(n1792), .Z(n1795) );
  CANR2X2 U2377 ( .A(n1129), .B(n2086), .C(n2018), .D(n1795), .Z(n1809) );
  CIVDX1 U2378 ( .A(n1796), .Z0(n1800), .Z1(n2373) );
  CND2X2 U2379 ( .A(n1798), .B(n1797), .Z(n2713) );
  CND2X1 U2380 ( .A(n2713), .B(n1922), .Z(n1799) );
  COND1XL U2381 ( .A(n2053), .B(n2068), .C(n2337), .Z(n1801) );
  CANR1X1 U2382 ( .A(n2090), .B(n2332), .C(n1801), .Z(n1808) );
  CNR2X1 U2383 ( .A(n1906), .B(n1905), .Z(n2001) );
  CIVX2 U2384 ( .A(n2002), .Z(n1802) );
  COND2X2 U2385 ( .A(n2087), .B(n2001), .C(n1802), .D(n1563), .Z(n1806) );
  CND2XL U2386 ( .A(n1922), .B(n1995), .Z(n1803) );
  CND2X1 U2387 ( .A(n1804), .B(n1803), .Z(n1805) );
  CND2X1 U2388 ( .A(n2190), .B(n2034), .Z(n1807) );
  CND3X2 U2389 ( .A(n1809), .B(n1808), .C(n1807), .Z(n2608) );
  CNR2X2 U2390 ( .A(n2607), .B(n2608), .Z(n2296) );
  CNR2IXL U2391 ( .B(n2373), .A(n1811), .Z(n1812) );
  CND2X1 U2392 ( .A(n1892), .B(n2368), .Z(n1816) );
  CND2X1 U2393 ( .A(n1894), .B(n2169), .Z(n1815) );
  CND2X1 U2394 ( .A(n1877), .B(n2371), .Z(n1814) );
  CND4X2 U2395 ( .A(n1817), .B(n1816), .C(n1815), .D(n1814), .Z(n2319) );
  CNR3X2 U2396 ( .A(n1824), .B(n1823), .C(n1822), .Z(n1834) );
  CND2XL U2397 ( .A(n1895), .B(n1893), .Z(n1826) );
  CND2X1 U2398 ( .A(n1826), .B(n1825), .Z(n1830) );
  CND2XL U2399 ( .A(n1889), .B(n2371), .Z(n1828) );
  CND2X1 U2400 ( .A(n1828), .B(n1827), .Z(n1829) );
  CNR2X2 U2401 ( .A(n1830), .B(n1829), .Z(n2189) );
  CND2X2 U2402 ( .A(n2189), .B(n2034), .Z(n1833) );
  CIVX1 U2403 ( .A(n1878), .Z(n1831) );
  CND2X1 U2404 ( .A(n2321), .B(n2090), .Z(n1832) );
  CND4X2 U2405 ( .A(n1834), .B(n1835), .C(n1833), .D(n1832), .Z(n2605) );
  CIVXL U2406 ( .A(n1836), .Z(n1837) );
  COND1XL U2407 ( .A(n1838), .B(n1837), .C(n2113), .Z(n1871) );
  CND2X1 U2408 ( .A(n1839), .B(n2151), .Z(n1868) );
  CND3XL U2409 ( .A(n1843), .B(n1842), .C(n2371), .Z(n2196) );
  CND3XL U2410 ( .A(n1865), .B(n2196), .C(n2198), .Z(n1853) );
  CND2X1 U2411 ( .A(n2154), .B(n2146), .Z(n1869) );
  CND2X1 U2412 ( .A(n1847), .B(n2373), .Z(n1850) );
  CND2X1 U2413 ( .A(n2370), .B(n2014), .Z(n1849) );
  CANR1X1 U2414 ( .A(h2[3]), .B(n2173), .C(n2371), .Z(n1848) );
  CND2X1 U2415 ( .A(n2324), .B(n2090), .Z(n1851) );
  COND11X2 U2416 ( .A(n1852), .B(n1854), .C(n1853), .D(n1851), .Z(n2604) );
  CNR2XL U2417 ( .A(n1856), .B(n1855), .Z(n1860) );
  COND1X1 U2418 ( .A(n1858), .B(n1857), .C(n2368), .Z(n1859) );
  CNR2X1 U2419 ( .A(n2129), .B(n2344), .Z(n1867) );
  CIVX2 U2420 ( .A(n1865), .Z(n1866) );
  CNR2IX1 U2421 ( .B(n1867), .A(n1866), .Z(n1870) );
  CND4X1 U2422 ( .A(n1107), .B(n1870), .C(n1869), .D(n1868), .Z(n1872) );
  CNR3X2 U2423 ( .A(n2605), .B(n2604), .C(n2603), .Z(n2297) );
  CND2X2 U2424 ( .A(n2296), .B(n2297), .Z(n2670) );
  CIVX2 U2425 ( .A(n2670), .Z(n2523) );
  CIVX2 U2426 ( .A(n1874), .Z(n1875) );
  CND2IX2 U2427 ( .B(n1876), .A(n1875), .Z(n2380) );
  CND2X1 U2428 ( .A(n1877), .B(n2176), .Z(n1880) );
  CND2X1 U2429 ( .A(n1878), .B(h2[2]), .Z(n1879) );
  CND2X2 U2430 ( .A(n1880), .B(n1879), .Z(n2092) );
  CND2X1 U2431 ( .A(n2508), .B(h2[5]), .Z(n1881) );
  CNR2X2 U2432 ( .A(n1882), .B(n1883), .Z(n2381) );
  CIVXL U2433 ( .A(n2349), .Z(n1884) );
  CND2X2 U2434 ( .A(n1189), .B(n1888), .Z(n2509) );
  CIVX2 U2435 ( .A(n1889), .Z(n1890) );
  CND2X2 U2436 ( .A(n1890), .B(n2137), .Z(n2387) );
  CND2X1 U2437 ( .A(n1891), .B(n2014), .Z(n2386) );
  CND2X1 U2438 ( .A(n1892), .B(n2371), .Z(n2385) );
  CND2X1 U2439 ( .A(n1894), .B(n1893), .Z(n2384) );
  CND3X1 U2440 ( .A(n1898), .B(n1896), .C(n1897), .Z(n2829) );
  CND2X1 U2441 ( .A(n1899), .B(n2368), .Z(n2035) );
  CND2X1 U2442 ( .A(n2035), .B(n2349), .Z(n1900) );
  CNR2X2 U2443 ( .A(n2829), .B(n1900), .Z(n1901) );
  CIVX2 U2444 ( .A(n1901), .Z(n1902) );
  CNR3X2 U2445 ( .A(n1904), .B(n2509), .C(n2506), .Z(n2317) );
  CND2X1 U2446 ( .A(n2000), .B(n1922), .Z(n1911) );
  CIVXL U2447 ( .A(n1905), .Z(n1908) );
  CIVX2 U2448 ( .A(n1906), .Z(n1907) );
  CND3X1 U2449 ( .A(n1908), .B(n2099), .C(n1907), .Z(n1910) );
  CIVX2 U2450 ( .A(n2045), .Z(n2376) );
  COR2X1 U2451 ( .A(n2121), .B(n2376), .Z(n3395) );
  CND2X1 U2452 ( .A(n2127), .B(h2[2]), .Z(n1913) );
  CND2X2 U2453 ( .A(n1914), .B(n1913), .Z(n2080) );
  CND2X1 U2454 ( .A(n2218), .B(h2[3]), .Z(n1915) );
  CND2X1 U2455 ( .A(n1915), .B(n2087), .Z(n2081) );
  CNR2X1 U2456 ( .A(n2081), .B(n2080), .Z(n3571) );
  COR2X1 U2457 ( .A(n1916), .B(n3571), .Z(n1921) );
  CND2XL U2458 ( .A(n1164), .B(n2371), .Z(n1917) );
  CND2XL U2459 ( .A(n2004), .B(n2373), .Z(n1918) );
  CND2X1 U2460 ( .A(n1919), .B(n1918), .Z(n2049) );
  CND2X1 U2461 ( .A(n1153), .B(n1922), .Z(n1925) );
  CND2IX1 U2462 ( .B(n1223), .A(n2126), .Z(n1924) );
  CND4X2 U2463 ( .A(n1926), .B(n1925), .C(n1924), .D(n1923), .Z(n2395) );
  CND2XL U2464 ( .A(n2395), .B(n2344), .Z(n3356) );
  CND2X2 U2465 ( .A(n2012), .B(n2161), .Z(n1927) );
  CND2X2 U2466 ( .A(n1927), .B(n2087), .Z(n2378) );
  CIVX2 U2467 ( .A(n2378), .Z(n1931) );
  CIVX2 U2468 ( .A(n2713), .Z(n2353) );
  CND2X2 U2469 ( .A(n2353), .B(h2[3]), .Z(n1929) );
  CND2X1 U2470 ( .A(n2011), .B(h2[2]), .Z(n1928) );
  CND2X2 U2471 ( .A(n1929), .B(n1928), .Z(n2377) );
  CIVX2 U2472 ( .A(n2377), .Z(n1930) );
  CND2X2 U2473 ( .A(n1931), .B(n1930), .Z(n2044) );
  CND2XL U2474 ( .A(n2044), .B(h2[5]), .Z(n3394) );
  CND2XL U2475 ( .A(n2098), .B(n2371), .Z(n1933) );
  CND2XL U2476 ( .A(n2100), .B(n2368), .Z(n1932) );
  CND2X1 U2477 ( .A(n1933), .B(n1932), .Z(n2066) );
  CIVXL U2478 ( .A(n2066), .Z(n1941) );
  CIVXL U2479 ( .A(n2115), .Z(n1934) );
  CND2X1 U2480 ( .A(n1939), .B(n1938), .Z(n2065) );
  CIVXL U2481 ( .A(n2065), .Z(n1940) );
  CND3X1 U2482 ( .A(n1941), .B(n2349), .C(n1940), .Z(n3354) );
  CND3X1 U2483 ( .A(n3356), .B(n3394), .C(n3354), .Z(n1942) );
  CNR2X2 U2484 ( .A(n1943), .B(n1942), .Z(n2360) );
  CND2X2 U2485 ( .A(n2360), .B(n2317), .Z(n2553) );
  CND2X2 U2486 ( .A(n2523), .B(n2585), .Z(n2033) );
  CND3XL U2487 ( .A(n1945), .B(n1944), .C(n2349), .Z(n1947) );
  CNR2X1 U2488 ( .A(n1947), .B(n1946), .Z(n1949) );
  CNR2X2 U2489 ( .A(n1950), .B(n1951), .Z(n2363) );
  COND1X2 U2490 ( .A(n1953), .B(n1952), .C(h2[5]), .Z(n1954) );
  COND1X1 U2491 ( .A(n2121), .B(n2363), .C(n1954), .Z(n2917) );
  CIVX2 U2492 ( .A(n2507), .Z(n3355) );
  CNR2X2 U2493 ( .A(n2917), .B(n2850), .Z(n1957) );
  CANR1X1 U2494 ( .A(n2349), .B(n1956), .C(n2507), .Z(n2916) );
  CND3X2 U2495 ( .A(n1957), .B(n2852), .C(n2916), .Z(n2421) );
  CIVX2 U2496 ( .A(n2421), .Z(n1976) );
  CIVX2 U2497 ( .A(h2[5]), .Z(n1958) );
  COND2X2 U2498 ( .A(n1958), .B(n2403), .C(n2392), .D(n2121), .Z(n2847) );
  CND2X1 U2499 ( .A(n1960), .B(n1959), .Z(n1966) );
  CND2X1 U2500 ( .A(n1963), .B(n2373), .Z(n2409) );
  CANR1X1 U2501 ( .A(n2090), .B(n2409), .C(h2[6]), .Z(n1964) );
  COND1X1 U2502 ( .A(n1966), .B(n1965), .C(n1964), .Z(n2520) );
  CNR2X2 U2503 ( .A(n2847), .B(n2520), .Z(n1974) );
  COND1X1 U2504 ( .A(n1161), .B(n1968), .C(n2086), .Z(n1969) );
  CND2X1 U2505 ( .A(n1970), .B(n1969), .Z(n2521) );
  CND2X1 U2506 ( .A(n1972), .B(n3355), .Z(n2848) );
  CNR2X2 U2507 ( .A(n2521), .B(n2848), .Z(n1973) );
  CND2X2 U2508 ( .A(n1974), .B(n1973), .Z(n2420) );
  CIVX2 U2509 ( .A(n2420), .Z(n1975) );
  CND2X2 U2510 ( .A(n1976), .B(n1975), .Z(n2554) );
  CIVX3 U2511 ( .A(n2554), .Z(n2586) );
  CND2IXL U2512 ( .B(n2121), .A(n1977), .Z(n1978) );
  CIVXL U2513 ( .A(n1978), .Z(n1990) );
  CIVXL U2514 ( .A(n1981), .Z(n1982) );
  CND2X1 U2515 ( .A(n1983), .B(n2146), .Z(n1986) );
  CND2XL U2516 ( .A(n2037), .B(n2151), .Z(n1984) );
  CND4X1 U2517 ( .A(n1985), .B(n1986), .C(n1987), .D(n1984), .Z(n1988) );
  CNR2X1 U2518 ( .A(n1992), .B(n1991), .Z(n2315) );
  CND2X1 U2519 ( .A(n2315), .B(n2582), .Z(n1994) );
  CND2X1 U2520 ( .A(n2137), .B(n2344), .Z(n2128) );
  CIVX1 U2521 ( .A(n2128), .Z(n2017) );
  CND3XL U2522 ( .A(n2707), .B(n2129), .C(n2017), .Z(n1993) );
  CND2X2 U2523 ( .A(n1994), .B(n1993), .Z(n2299) );
  CIVX2 U2524 ( .A(n1999), .Z(n2346) );
  CND2IX1 U2525 ( .B(n2087), .A(n1119), .Z(n2347) );
  COND1XL U2526 ( .A(n2147), .B(n2002), .C(n2153), .Z(n2006) );
  CNR2XL U2527 ( .A(n2004), .B(n2003), .Z(n2005) );
  CNR2X1 U2528 ( .A(n2006), .B(n2005), .Z(n2009) );
  CANR2X1 U2529 ( .A(n2012), .B(n2368), .C(n2371), .D(n2011), .Z(n2342) );
  CND2X1 U2530 ( .A(n1177), .B(n2582), .Z(n2016) );
  CIVX2 U2531 ( .A(n2016), .Z(n2020) );
  CND2XL U2532 ( .A(n2713), .B(n2017), .Z(n2423) );
  CNR2X1 U2533 ( .A(n2423), .B(n2018), .Z(n2019) );
  CANR1X2 U2534 ( .A(n2342), .B(n2020), .C(n2019), .Z(n2021) );
  CND2X2 U2535 ( .A(n2022), .B(n2021), .Z(n3384) );
  COND1X2 U2536 ( .A(n2298), .B(n2299), .C(n3384), .Z(n2023) );
  CIVX2 U2537 ( .A(n2023), .Z(n2030) );
  CNR2X1 U2538 ( .A(n2027), .B(n2026), .Z(n2029) );
  CIVX2 U2539 ( .A(n2522), .Z(n2031) );
  CND2X2 U2540 ( .A(n2031), .B(n2586), .Z(n2032) );
  CND2X1 U2541 ( .A(n2035), .B(n2034), .Z(n2828) );
  CND2IX1 U2542 ( .B(n2073), .A(n2036), .Z(n2039) );
  CNR2X2 U2543 ( .A(n2826), .B(n2825), .Z(n2043) );
  COND1X1 U2544 ( .A(n2828), .B(n1160), .C(n2043), .Z(n2048) );
  CND2X2 U2545 ( .A(n2044), .B(n2090), .Z(n2047) );
  CND2X2 U2546 ( .A(n1146), .B(n2086), .Z(n2046) );
  CND2X2 U2547 ( .A(n2047), .B(n2046), .Z(n2824) );
  CNR2X2 U2548 ( .A(n2048), .B(n2824), .Z(n2079) );
  CNR3X1 U2549 ( .A(n1120), .B(n2049), .C(n2064), .Z(n2063) );
  CND2X1 U2550 ( .A(n2051), .B(n2050), .Z(n2057) );
  CND2X1 U2551 ( .A(n2052), .B(n1194), .Z(n2056) );
  CNR2X1 U2552 ( .A(n2053), .B(n2073), .Z(n2054) );
  CIVX2 U2553 ( .A(n2054), .Z(n2055) );
  CND3X1 U2554 ( .A(n2057), .B(n2056), .C(n2055), .Z(n2061) );
  CANR1XL U2555 ( .A(n2059), .B(n2058), .C(h2[6]), .Z(n2060) );
  CNR3X1 U2556 ( .A(n2066), .B(n2065), .C(n2064), .Z(n2078) );
  CNR2X1 U2557 ( .A(n2068), .B(n2067), .Z(n2071) );
  COND1X2 U2558 ( .A(n2069), .B(n2117), .C(n2337), .Z(n2070) );
  CNR2X2 U2559 ( .A(n2071), .B(n2070), .Z(n2076) );
  CND2X1 U2560 ( .A(n2109), .B(n1194), .Z(n2074) );
  CND3X1 U2561 ( .A(n2076), .B(n2075), .C(n2074), .Z(n2077) );
  CNR2X2 U2562 ( .A(n2078), .B(n2077), .Z(n2833) );
  CND3X2 U2563 ( .A(n2079), .B(n1115), .C(n2833), .Z(n2445) );
  CIVX2 U2564 ( .A(n2080), .Z(n2083) );
  CIVX2 U2565 ( .A(n2081), .Z(n2082) );
  CND2X2 U2566 ( .A(n2083), .B(n2082), .Z(n2397) );
  CND2X2 U2567 ( .A(n2397), .B(n2090), .Z(n2085) );
  CND2X2 U2568 ( .A(n2395), .B(n2086), .Z(n2084) );
  CND2X2 U2569 ( .A(n2085), .B(n2084), .Z(n2832) );
  COND1XL U2570 ( .A(n2089), .B(n2088), .C(n2087), .Z(n2091) );
  CND2X2 U2571 ( .A(n2094), .B(n2093), .Z(n2830) );
  CNR2X2 U2572 ( .A(n2445), .B(n1118), .Z(n2793) );
  CND2XL U2573 ( .A(n2103), .B(n2368), .Z(n2107) );
  CIVXL U2574 ( .A(n1153), .Z(n2105) );
  CND2IX1 U2575 ( .B(n2087), .A(n2105), .Z(n2106) );
  CND3X2 U2576 ( .A(n2108), .B(n2107), .C(n2106), .Z(n2220) );
  CND2XL U2577 ( .A(n2110), .B(n2146), .Z(n2111) );
  CND3X1 U2578 ( .A(n2112), .B(n2111), .C(n2153), .Z(n2119) );
  CND3XL U2579 ( .A(n2115), .B(n2114), .C(n2113), .Z(n2116) );
  COND1X1 U2580 ( .A(n2121), .B(n2220), .C(n2120), .Z(n2134) );
  CND2XL U2581 ( .A(n2124), .B(n2368), .Z(n2215) );
  CND2XL U2582 ( .A(n2216), .B(n2215), .Z(n2132) );
  CND2XL U2583 ( .A(n2127), .B(n2371), .Z(n2214) );
  CND3XL U2584 ( .A(n2217), .B(n2582), .C(n2214), .Z(n2131) );
  CNR2XL U2585 ( .A(n2218), .B(n2128), .Z(n2428) );
  CND2XL U2586 ( .A(n2428), .B(n2129), .Z(n2130) );
  COAN1X1 U2587 ( .A(n2132), .B(n2131), .C(n2130), .Z(n2133) );
  CND2X2 U2588 ( .A(n2134), .B(n2133), .Z(n2417) );
  CND2X1 U2589 ( .A(n2135), .B(n2417), .Z(n2184) );
  CND2XL U2590 ( .A(n2136), .B(n2169), .Z(n2258) );
  CND2XL U2591 ( .A(n2138), .B(n2137), .Z(n2257) );
  CND3XL U2592 ( .A(n1179), .B(n2257), .C(n2268), .Z(n2139) );
  CIVXL U2593 ( .A(n2139), .Z(n2144) );
  CIVXL U2594 ( .A(n2140), .Z(n2141) );
  CND2X1 U2595 ( .A(n2141), .B(n2368), .Z(n2260) );
  CIVXL U2596 ( .A(n2142), .Z(n2143) );
  CND2X1 U2597 ( .A(n2143), .B(n2371), .Z(n2259) );
  CND3X1 U2598 ( .A(n2144), .B(n2260), .C(n2259), .Z(n2160) );
  CNR2XL U2599 ( .A(n1149), .B(n2147), .Z(n2149) );
  CNR2X1 U2600 ( .A(n2150), .B(n2149), .Z(n2159) );
  COND1XL U2601 ( .A(n2155), .B(n2154), .C(n2153), .Z(n2156) );
  CNR2X1 U2602 ( .A(n2157), .B(n2156), .Z(n2158) );
  CND3X2 U2603 ( .A(n2160), .B(n2159), .C(n2158), .Z(n2295) );
  CND2X1 U2604 ( .A(n2162), .B(n2161), .Z(n2264) );
  CIVXL U2605 ( .A(n2163), .Z(n2166) );
  CIVXL U2606 ( .A(n2164), .Z(n2165) );
  CND2X2 U2607 ( .A(n2264), .B(n2265), .Z(n2437) );
  CIVX1 U2608 ( .A(n2582), .Z(n2167) );
  CNR2X2 U2609 ( .A(n2437), .B(n2167), .Z(n2180) );
  CND2X1 U2610 ( .A(n2168), .B(n2368), .Z(n2433) );
  CIVX2 U2611 ( .A(n2433), .Z(n2171) );
  CIVX2 U2612 ( .A(n2431), .Z(n2170) );
  CNR2X1 U2613 ( .A(n2171), .B(n2170), .Z(n2179) );
  CANR1X1 U2614 ( .A(n2176), .B(n2175), .C(n2174), .Z(n2434) );
  CANR1X1 U2615 ( .A(n2180), .B(n2179), .C(n2178), .Z(n2294) );
  CND2X1 U2616 ( .A(n2295), .B(n2294), .Z(n2182) );
  CND2X2 U2617 ( .A(n2181), .B(n2182), .Z(n2183) );
  CNR2X2 U2618 ( .A(n2184), .B(n2183), .Z(n2504) );
  CND2X2 U2619 ( .A(n2793), .B(n2504), .Z(n3129) );
  CND2X1 U2620 ( .A(n2319), .B(n2268), .Z(n2186) );
  CND2X1 U2621 ( .A(n2186), .B(n2185), .Z(n2282) );
  CND2XL U2622 ( .A(n2332), .B(h2[5]), .Z(n2187) );
  CAN2X2 U2623 ( .A(n1074), .B(n3127), .Z(n2415) );
  CND2X2 U2624 ( .A(n2416), .B(n2415), .Z(n2191) );
  CIVX2 U2625 ( .A(n2191), .Z(n2213) );
  CND2X2 U2626 ( .A(n2335), .B(n2344), .Z(n2193) );
  CND2X2 U2627 ( .A(n2193), .B(n2192), .Z(n3132) );
  CIVX2 U2628 ( .A(n3132), .Z(n2211) );
  CAN2X1 U2629 ( .A(n1152), .B(n2196), .Z(n2279) );
  CND2X1 U2630 ( .A(n2197), .B(n2349), .Z(n2200) );
  CIVX2 U2631 ( .A(n2198), .Z(n2199) );
  CND3XL U2632 ( .A(n2204), .B(n2202), .C(n2203), .Z(n2205) );
  COND1X1 U2633 ( .A(n2206), .B(n2205), .C(n3355), .Z(n3131) );
  CIVX2 U2634 ( .A(n3131), .Z(n2207) );
  CANR1X1 U2635 ( .A(h2[5]), .B(n1169), .C(n2507), .Z(n2280) );
  CND2X2 U2636 ( .A(n2207), .B(n2280), .Z(n2208) );
  CIVX2 U2637 ( .A(n2208), .Z(n2209) );
  CIVX2 U2638 ( .A(n1104), .Z(n2212) );
  CND2X2 U2639 ( .A(n2212), .B(n2213), .Z(n2561) );
  CNR2X1 U2640 ( .A(n2561), .B(n3129), .Z(n2275) );
  CND2X1 U2641 ( .A(n2215), .B(n2214), .Z(n2427) );
  CND2X1 U2642 ( .A(n2217), .B(n2216), .Z(n2426) );
  CND2XL U2643 ( .A(n2218), .B(h2[5]), .Z(n2219) );
  CND2X1 U2644 ( .A(n1178), .B(n2219), .Z(n2556) );
  CIVX2 U2645 ( .A(n2220), .Z(n2221) );
  CNR2X1 U2646 ( .A(n2556), .B(n1182), .Z(n3106) );
  CND2X1 U2647 ( .A(n3106), .B(n3269), .Z(n2270) );
  CNR2X1 U2648 ( .A(n1139), .B(mulout[29]), .Z(n2458) );
  CND2X1 U2649 ( .A(n1139), .B(mulout[29]), .Z(n2457) );
  CNR2X1 U2650 ( .A(acc[16]), .B(mulout[16]), .Z(n2858) );
  CNR2X1 U2651 ( .A(acc[17]), .B(mulout[17]), .Z(n2855) );
  CNR2X1 U2652 ( .A(n2858), .B(n2855), .Z(n2927) );
  CNR2X1 U2653 ( .A(acc[18]), .B(mulout[18]), .Z(n2924) );
  CNR2X1 U2654 ( .A(acc[19]), .B(mulout[19]), .Z(n2732) );
  CNR2X1 U2655 ( .A(n2924), .B(n2732), .Z(n2242) );
  CND2X1 U2656 ( .A(n2927), .B(n2242), .Z(n3363) );
  CNR2X1 U2657 ( .A(acc[20]), .B(mulout[20]), .Z(n3366) );
  CNR2X1 U2658 ( .A(acc[21]), .B(mulout[21]), .Z(n3361) );
  CNR2X1 U2659 ( .A(n3366), .B(n3361), .Z(n3094) );
  CNR2X1 U2660 ( .A(acc[22]), .B(mulout[22]), .Z(n3398) );
  CNR2X1 U2661 ( .A(acc[23]), .B(mulout[23]), .Z(n3089) );
  CNR2X1 U2662 ( .A(n3398), .B(n3089), .Z(n2244) );
  CND2X1 U2663 ( .A(n3094), .B(n2244), .Z(n2246) );
  CNR2X1 U2664 ( .A(n3363), .B(n2246), .Z(n2456) );
  CIVX1 U2665 ( .A(n2456), .Z(n3483) );
  CNR2X1 U2666 ( .A(acc[24]), .B(mulout[24]), .Z(n3215) );
  CNR2X1 U2667 ( .A(acc[25]), .B(mulout[25]), .Z(n3212) );
  CNR2X1 U2668 ( .A(n3215), .B(n3212), .Z(n3482) );
  CNR2X1 U2669 ( .A(acc[26]), .B(mulout[26]), .Z(n3145) );
  CNR2X1 U2670 ( .A(acc[27]), .B(mulout[27]), .Z(n3479) );
  CNR2X1 U2671 ( .A(n3145), .B(n3479), .Z(n2248) );
  CND2X1 U2672 ( .A(n3482), .B(n2248), .Z(n3195) );
  CIVX1 U2673 ( .A(n3195), .Z(n3112) );
  CNR2X1 U2674 ( .A(acc[28]), .B(mulout[28]), .Z(n2455) );
  CIVX1 U2675 ( .A(n2455), .Z(n3193) );
  CND2XL U2676 ( .A(n3112), .B(n3193), .Z(n2251) );
  CNR2XL U2677 ( .A(n3483), .B(n2251), .Z(n2253) );
  CNR2X1 U2678 ( .A(acc[4]), .B(mulout[4]), .Z(n3294) );
  CNR2X1 U2679 ( .A(acc[5]), .B(mulout[5]), .Z(n3292) );
  CNR2X1 U2680 ( .A(n3294), .B(n3292), .Z(n2843) );
  CNR2X1 U2681 ( .A(acc[6]), .B(mulout[6]), .Z(n3467) );
  CNR2X1 U2682 ( .A(acc[7]), .B(mulout[7]), .Z(n3468) );
  CNR2X1 U2683 ( .A(n3467), .B(n3468), .Z(n2230) );
  CND2X1 U2684 ( .A(n2843), .B(n2230), .Z(n2232) );
  CNR2X1 U2685 ( .A(n2222), .B(n2224), .Z(n2227) );
  COND1XL U2686 ( .A(n2225), .B(n2224), .C(n2223), .Z(n2226) );
  CANR1X1 U2687 ( .A(n2228), .B(n2227), .C(n2226), .Z(n2841) );
  CND2X1 U2688 ( .A(acc[4]), .B(mulout[4]), .Z(n3438) );
  CND2X1 U2689 ( .A(acc[5]), .B(mulout[5]), .Z(n3293) );
  COND1XL U2690 ( .A(n3438), .B(n3292), .C(n3293), .Z(n2842) );
  CND2X1 U2691 ( .A(acc[6]), .B(mulout[6]), .Z(n3465) );
  CND2X1 U2692 ( .A(acc[7]), .B(mulout[7]), .Z(n3469) );
  COND1XL U2693 ( .A(n3465), .B(n3468), .C(n3469), .Z(n2229) );
  CANR1XL U2694 ( .A(n2842), .B(n2230), .C(n2229), .Z(n2231) );
  COND1X1 U2695 ( .A(n2232), .B(n2841), .C(n2231), .Z(n2303) );
  CNR2X1 U2696 ( .A(acc[8]), .B(mulout[8]), .Z(n3375) );
  CNR2X1 U2697 ( .A(acc[9]), .B(mulout[9]), .Z(n3282) );
  CNR2X1 U2698 ( .A(n3375), .B(n3282), .Z(n2611) );
  CNR2X1 U2699 ( .A(acc[10]), .B(mulout[10]), .Z(n2615) );
  CNR2X1 U2700 ( .A(acc[11]), .B(mulout[11]), .Z(n2908) );
  CNR2X1 U2701 ( .A(n2615), .B(n2908), .Z(n2234) );
  CND2X1 U2702 ( .A(n2611), .B(n2234), .Z(n3453) );
  CNR2X1 U2703 ( .A(acc[12]), .B(mulout[12]), .Z(n2302) );
  CNR2X1 U2704 ( .A(acc[13]), .B(mulout[13]), .Z(n2304) );
  CNR2X1 U2705 ( .A(n2302), .B(n2304), .Z(n2531) );
  CNR2X1 U2706 ( .A(acc[14]), .B(mulout[14]), .Z(n2527) );
  CNR2X1 U2707 ( .A(acc[15]), .B(mulout[15]), .Z(n2525) );
  CNR2X1 U2708 ( .A(n2527), .B(n2525), .Z(n2236) );
  CND2X1 U2709 ( .A(n2531), .B(n2236), .Z(n2238) );
  CNR2X1 U2710 ( .A(n3453), .B(n2238), .Z(n2240) );
  CND2X1 U2711 ( .A(acc[8]), .B(mulout[8]), .Z(n3376) );
  CND2X1 U2712 ( .A(acc[9]), .B(mulout[9]), .Z(n3283) );
  COND1X1 U2713 ( .A(n3376), .B(n3282), .C(n3283), .Z(n2612) );
  CND2X1 U2714 ( .A(acc[10]), .B(mulout[10]), .Z(n2910) );
  CND2X1 U2715 ( .A(acc[11]), .B(mulout[11]), .Z(n2909) );
  COND1XL U2716 ( .A(n2910), .B(n2908), .C(n2909), .Z(n2233) );
  CANR1X1 U2717 ( .A(n2612), .B(n2234), .C(n2233), .Z(n3451) );
  CND2X1 U2718 ( .A(acc[12]), .B(mulout[12]), .Z(n3454) );
  CND2XL U2719 ( .A(acc[13]), .B(mulout[13]), .Z(n2305) );
  COND1XL U2720 ( .A(n3454), .B(n2304), .C(n2305), .Z(n2529) );
  CND2X1 U2721 ( .A(acc[14]), .B(mulout[14]), .Z(n3379) );
  CND2X1 U2722 ( .A(acc[15]), .B(mulout[15]), .Z(n2526) );
  COND1XL U2723 ( .A(n3379), .B(n2525), .C(n2526), .Z(n2235) );
  CANR1XL U2724 ( .A(n2529), .B(n2236), .C(n2235), .Z(n2237) );
  COND1XL U2725 ( .A(n2238), .B(n3451), .C(n2237), .Z(n2239) );
  CANR1X1 U2726 ( .A(n2303), .B(n2240), .C(n2239), .Z(n2467) );
  CIVX2 U2727 ( .A(n2467), .Z(n3504) );
  CND2X1 U2728 ( .A(acc[16]), .B(mulout[16]), .Z(n3502) );
  CND2X1 U2729 ( .A(acc[17]), .B(mulout[17]), .Z(n2856) );
  COND1X1 U2730 ( .A(n3502), .B(n2855), .C(n2856), .Z(n2926) );
  CND2X1 U2731 ( .A(acc[18]), .B(mulout[18]), .Z(n2925) );
  CND2X1 U2732 ( .A(acc[19]), .B(mulout[19]), .Z(n2733) );
  COND1X1 U2733 ( .A(n2925), .B(n2732), .C(n2733), .Z(n2241) );
  CANR1X1 U2734 ( .A(n2926), .B(n2242), .C(n2241), .Z(n3365) );
  CND2X1 U2735 ( .A(acc[20]), .B(mulout[20]), .Z(n3364) );
  CND2X1 U2736 ( .A(acc[21]), .B(mulout[21]), .Z(n3362) );
  COND1XL U2737 ( .A(n3364), .B(n3361), .C(n3362), .Z(n3092) );
  CND2X1 U2738 ( .A(acc[22]), .B(mulout[22]), .Z(n3399) );
  CND2X1 U2739 ( .A(acc[23]), .B(mulout[23]), .Z(n3090) );
  COND1XL U2740 ( .A(n3399), .B(n3089), .C(n3090), .Z(n2243) );
  CANR1XL U2741 ( .A(n3092), .B(n2244), .C(n2243), .Z(n2245) );
  COND1X1 U2742 ( .A(n2246), .B(n3365), .C(n2245), .Z(n2465) );
  CIVX1 U2743 ( .A(n2465), .Z(n3489) );
  CND2X1 U2744 ( .A(acc[24]), .B(mulout[24]), .Z(n3214) );
  CND2X1 U2745 ( .A(acc[25]), .B(mulout[25]), .Z(n3213) );
  COND1XL U2746 ( .A(n3214), .B(n3212), .C(n3213), .Z(n3486) );
  CND2X1 U2747 ( .A(acc[26]), .B(mulout[26]), .Z(n3484) );
  CND2X1 U2748 ( .A(acc[27]), .B(mulout[27]), .Z(n3480) );
  COND1XL U2749 ( .A(n3484), .B(n3479), .C(n3480), .Z(n2247) );
  CANR1XL U2750 ( .A(n3486), .B(n2248), .C(n2247), .Z(n3194) );
  CIVXL U2751 ( .A(n3194), .Z(n3114) );
  CND2X1 U2752 ( .A(acc[28]), .B(mulout[28]), .Z(n3192) );
  CIVXL U2753 ( .A(n3192), .Z(n2249) );
  CANR1XL U2754 ( .A(n3193), .B(n3114), .C(n2249), .Z(n2250) );
  COND1XL U2755 ( .A(n2251), .B(n3489), .C(n2250), .Z(n2252) );
  CANR1XL U2756 ( .A(n2253), .B(n3504), .C(n2252), .Z(n2254) );
  CEOXL U2757 ( .A(n2255), .B(n2254), .Z(n2256) );
  CND2XL U2758 ( .A(n2256), .B(n3595), .Z(n2272) );
  CND3XL U2759 ( .A(n2258), .B(n2257), .C(n2349), .Z(n2263) );
  CND2X1 U2760 ( .A(n2260), .B(n2259), .Z(n2262) );
  CND2XL U2761 ( .A(n2434), .B(h2[5]), .Z(n2261) );
  COAN1X1 U2762 ( .A(n2263), .B(n2262), .C(n2261), .Z(n2330) );
  CND3X1 U2763 ( .A(n2431), .B(n2265), .C(n3355), .Z(n2266) );
  COND2X2 U2764 ( .A(n2268), .B(n2507), .C(n2267), .D(n2266), .Z(n2329) );
  CND2X1 U2765 ( .A(n2330), .B(n2329), .Z(n3478) );
  CIVXL U2766 ( .A(n3478), .Z(n3205) );
  CANR2XL U2767 ( .A(n1659), .B(mulout[29]), .C(n1140), .D(n3617), .Z(n2269)
         );
  COND1XL U2768 ( .A(n3205), .B(n2270), .C(n2269), .Z(n2271) );
  CNR2IXL U2769 ( .B(n2272), .A(n2271), .Z(n2273) );
  CIVXL U2770 ( .A(n3207), .Z(n2277) );
  CNR2XL U2771 ( .A(n3106), .B(n3478), .Z(n2276) );
  CIVXL U2772 ( .A(n3101), .Z(n3190) );
  CAN2XL U2773 ( .A(n3190), .B(n3269), .Z(n3206) );
  CIVX2 U2774 ( .A(n3129), .Z(n2549) );
  CND2X1 U2775 ( .A(n1155), .B(n2549), .Z(n3099) );
  CANR2XL U2776 ( .A(n1131), .B(n2344), .C(n2279), .D(n2278), .Z(n2281) );
  CND2XL U2777 ( .A(n2280), .B(n2281), .Z(n3128) );
  CNR2XL U2778 ( .A(n3128), .B(n3325), .Z(n3088) );
  CND2XL U2779 ( .A(n3088), .B(n3225), .Z(n2284) );
  COAN1X1 U2780 ( .A(n3099), .B(n2284), .C(n2283), .Z(n2289) );
  CIVXL U2781 ( .A(n3225), .Z(n2287) );
  CND2XL U2782 ( .A(n3128), .B(n3269), .Z(n3100) );
  CANR2XL U2783 ( .A(n1659), .B(mulout[24]), .C(acc[24]), .D(n3617), .Z(n2285)
         );
  COND1XL U2784 ( .A(n3225), .B(n3100), .C(n2285), .Z(n2286) );
  CANR11X1 U2785 ( .A(n3269), .B(n2287), .C(n3099), .D(n2286), .Z(n2288) );
  CND2X1 U2786 ( .A(n2289), .B(n2288), .Z(n545) );
  CMX2XL U2787 ( .A0(h1[6]), .A1(h2[6]), .S(rst), .Z(n504) );
  CND2XL U2788 ( .A(n3387), .B(n3269), .Z(n2301) );
  CIVXL U2789 ( .A(n2669), .Z(n2293) );
  CND2X1 U2790 ( .A(n2793), .B(n2290), .Z(n2291) );
  CIVX2 U2791 ( .A(n2291), .Z(n2292) );
  CND2X2 U2792 ( .A(n2292), .B(n2293), .Z(n3463) );
  CND2X1 U2793 ( .A(n2295), .B(n712), .Z(n2905) );
  CND2X1 U2794 ( .A(n2296), .B(n713), .Z(n3448) );
  CIVXL U2795 ( .A(n3448), .Z(n3444) );
  CNR2X1 U2796 ( .A(n2299), .B(n1175), .Z(n1102) );
  CIVXL U2797 ( .A(n1102), .Z(n3445) );
  CIVXL U2798 ( .A(n3453), .Z(n2528) );
  CIVX1 U2799 ( .A(n2302), .Z(n3455) );
  CIVX2 U2800 ( .A(n2303), .Z(n3452) );
  CIVXL U2801 ( .A(n3451), .Z(n2530) );
  CAOR2XL U2802 ( .A(n1659), .B(mulout[13]), .C(acc[13]), .D(n3617), .Z(n2306)
         );
  CANR1XL U2803 ( .A(n3595), .B(n2307), .C(n2306), .Z(n2310) );
  CIVXL U2804 ( .A(n2707), .Z(n2313) );
  CNR2X1 U2805 ( .A(n2313), .B(n2312), .Z(n2314) );
  CMXI2X1 U2806 ( .A0(n2315), .A1(n2314), .S(n2344), .Z(n2316) );
  CIVX2 U2807 ( .A(n2318), .Z(n2328) );
  CIVXL U2808 ( .A(n2319), .Z(n2320) );
  CNR2IX1 U2809 ( .B(n2337), .A(n2336), .Z(n3573) );
  CND2X1 U2810 ( .A(n2320), .B(n3573), .Z(n2884) );
  CNR2IX2 U2811 ( .B(n2268), .A(n2763), .Z(n2435) );
  CND2X1 U2812 ( .A(n2661), .B(n2435), .Z(n2883) );
  CND2X1 U2813 ( .A(n2884), .B(n2883), .Z(n2326) );
  CIVX2 U2814 ( .A(n2322), .Z(n2323) );
  CNR2IX1 U2815 ( .B(n2337), .A(n2336), .Z(n2979) );
  CND2X1 U2816 ( .A(n2323), .B(n2979), .Z(n2882) );
  CND2X1 U2817 ( .A(n2660), .B(n2435), .Z(n2881) );
  CND2X1 U2818 ( .A(n2882), .B(n2881), .Z(n2325) );
  CND2X1 U2819 ( .A(n2326), .B(n2325), .Z(n2548) );
  CNR2X1 U2820 ( .A(n1102), .B(n2548), .Z(n2327) );
  CND2X2 U2821 ( .A(n2328), .B(n2327), .Z(n2658) );
  CND2X2 U2822 ( .A(n2330), .B(n2329), .Z(n2555) );
  CNR2X2 U2823 ( .A(n2820), .B(n2555), .Z(n2359) );
  CIVXL U2824 ( .A(n1130), .Z(n2331) );
  CND2X1 U2825 ( .A(n2331), .B(n2979), .Z(n2334) );
  CIVX2 U2826 ( .A(n2332), .Z(n2663) );
  CND2X1 U2827 ( .A(n2663), .B(n2435), .Z(n2333) );
  CND2X2 U2828 ( .A(n2334), .B(n2333), .Z(n3528) );
  CIVX2 U2829 ( .A(n2335), .Z(n2338) );
  CNR2IX1 U2830 ( .B(n2337), .A(n2336), .Z(n2671) );
  CND2X2 U2831 ( .A(n2338), .B(n2671), .Z(n2341) );
  CIVXL U2832 ( .A(n2339), .Z(n2662) );
  CND2X1 U2833 ( .A(n2662), .B(n2435), .Z(n2340) );
  CND2X2 U2834 ( .A(n2341), .B(n2340), .Z(n3529) );
  CIVX2 U2835 ( .A(n1091), .Z(n2358) );
  CND2XL U2836 ( .A(n2343), .B(n2342), .Z(n2422) );
  CIVX2 U2837 ( .A(n2348), .Z(n2350) );
  CIVXL U2838 ( .A(n2351), .Z(n2352) );
  CANR1XL U2839 ( .A(h2[5]), .B(n2353), .C(n2352), .Z(n2354) );
  CNR2X2 U2840 ( .A(n1184), .B(n3101), .Z(n2357) );
  CND4X2 U2841 ( .A(n2359), .B(n2360), .C(n2357), .D(n2358), .Z(n2659) );
  CNR2X2 U2842 ( .A(n2658), .B(n2659), .Z(n2362) );
  CNR2X1 U2843 ( .A(n3448), .B(n2669), .Z(n2361) );
  CND2X2 U2844 ( .A(n2362), .B(n2361), .Z(n3554) );
  CIVX3 U2845 ( .A(n3554), .Z(n3551) );
  CIVX2 U2846 ( .A(n2435), .Z(n2396) );
  CND4X1 U2847 ( .A(n2407), .B(n2406), .C(n2405), .D(n2404), .Z(n2364) );
  CND2X1 U2848 ( .A(n2369), .B(n2368), .Z(n2410) );
  CND3XL U2849 ( .A(n2411), .B(n2410), .C(n2435), .Z(n2374) );
  CANR2XL U2850 ( .A(n2373), .B(n2372), .C(n2371), .D(n2370), .Z(n2413) );
  CIVX2 U2851 ( .A(n2380), .Z(n2447) );
  CND2X1 U2852 ( .A(n2447), .B(n2435), .Z(n2383) );
  CND2XL U2853 ( .A(n2671), .B(n1147), .Z(n2382) );
  CND2X1 U2854 ( .A(n2383), .B(n2382), .Z(n2874) );
  CIVXL U2855 ( .A(n2388), .Z(n2389) );
  CND2X1 U2856 ( .A(n2389), .B(n2979), .Z(n2391) );
  CND2X2 U2857 ( .A(n2391), .B(n2390), .Z(n2967) );
  CND2X2 U2858 ( .A(n2874), .B(n2967), .Z(n2401) );
  CND2X1 U2859 ( .A(n2392), .B(n3573), .Z(n2394) );
  CND2X1 U2860 ( .A(n2403), .B(n2435), .Z(n2393) );
  CND2X2 U2861 ( .A(n2394), .B(n2393), .Z(n2580) );
  CIVX2 U2862 ( .A(n2671), .Z(n3248) );
  CNR2X1 U2863 ( .A(n2395), .B(n3248), .Z(n2399) );
  COR2X2 U2864 ( .A(n2398), .B(n2399), .Z(n3060) );
  CND2X2 U2865 ( .A(n2580), .B(n3060), .Z(n2400) );
  CND2X1 U2866 ( .A(n2403), .B(n3573), .Z(n3299) );
  CNR2X2 U2867 ( .A(n2978), .B(n3299), .Z(n2414) );
  CND4XL U2868 ( .A(n2406), .B(n2407), .C(n2405), .D(n2404), .Z(n2408) );
  CNR2X1 U2869 ( .A(n3248), .B(n2408), .Z(n3326) );
  CIVX2 U2870 ( .A(n2409), .Z(n3250) );
  CND3X2 U2871 ( .A(n2414), .B(n3326), .C(n3348), .Z(n2746) );
  CIVXL U2872 ( .A(n2746), .Z(n2419) );
  CND2X1 U2873 ( .A(n3384), .B(n2417), .Z(n2675) );
  CNR3X1 U2874 ( .A(n2676), .B(n2674), .C(n2675), .Z(n2418) );
  CND3X1 U2875 ( .A(n1116), .B(n2419), .C(n2418), .Z(n2446) );
  CNR2X2 U2876 ( .A(n2421), .B(n2420), .Z(n2792) );
  CIVXL U2877 ( .A(n2422), .Z(n2425) );
  CIVX1 U2878 ( .A(n2423), .Z(n2424) );
  CANR1X1 U2879 ( .A(n2121), .B(n2425), .C(n2424), .Z(n2764) );
  CIVX1 U2880 ( .A(n2426), .Z(n2430) );
  CNR2X1 U2881 ( .A(n2427), .B(n2344), .Z(n2429) );
  CANR1X1 U2882 ( .A(n2430), .B(n2429), .C(n2428), .Z(n2569) );
  CNR2X2 U2883 ( .A(n2764), .B(n2569), .Z(n2442) );
  CNR2X1 U2884 ( .A(n2763), .B(n2344), .Z(n2432) );
  CIVX2 U2885 ( .A(n2434), .Z(n2672) );
  CND2X2 U2886 ( .A(n2672), .B(n2435), .Z(n2436) );
  CIVX2 U2887 ( .A(n2440), .Z(n2441) );
  CND3X2 U2888 ( .A(n2905), .B(n2441), .C(n2442), .Z(n2443) );
  CIVX2 U2889 ( .A(n2443), .Z(n2794) );
  CNR2X2 U2890 ( .A(n2444), .B(n2445), .Z(n2505) );
  CND3X2 U2891 ( .A(n2505), .B(n2792), .C(n1093), .Z(n2977) );
  CNR2X2 U2892 ( .A(n2446), .B(n2977), .Z(n3555) );
  CND2X1 U2893 ( .A(n2447), .B(n2979), .Z(n3569) );
  CND2X1 U2894 ( .A(n2448), .B(n2671), .Z(n3271) );
  CNR2X1 U2895 ( .A(n3569), .B(n3271), .Z(n2664) );
  CIVXL U2896 ( .A(n3571), .Z(n3353) );
  CNR2X1 U2897 ( .A(n3353), .B(n3248), .Z(n2451) );
  CIVXL U2898 ( .A(n2451), .Z(n2449) );
  CAN3XL U2899 ( .A(n2664), .B(n3269), .C(n2449), .Z(n2450) );
  CND2IX1 U2900 ( .B(n3276), .A(n2450), .Z(n2503) );
  CIVXL U2901 ( .A(n3271), .Z(n3261) );
  CND2X1 U2902 ( .A(n2451), .B(n3269), .Z(n2452) );
  CND2X1 U2903 ( .A(n1203), .B(n3569), .Z(n2453) );
  COR2X1 U2904 ( .A(mulout[53]), .B(acc[53]), .Z(n2639) );
  CND2X1 U2905 ( .A(mulout[53]), .B(acc[53]), .Z(n2637) );
  CND2XL U2906 ( .A(n2639), .B(n2637), .Z(n2494) );
  CNR2X1 U2907 ( .A(mulout[45]), .B(n858), .Z(n2574) );
  CNR2X1 U2908 ( .A(mulout[44]), .B(acc[44]), .Z(n2576) );
  CNR2X1 U2909 ( .A(n2574), .B(n2576), .Z(n3343) );
  CNR2X1 U2910 ( .A(mulout[46]), .B(acc[46]), .Z(n3346) );
  CNR2X1 U2911 ( .A(mulout[47]), .B(acc[47]), .Z(n3341) );
  CNR2X1 U2912 ( .A(n3346), .B(n3341), .Z(n2486) );
  CND2X1 U2913 ( .A(n3343), .B(n2486), .Z(n3304) );
  CNR2X1 U2914 ( .A(mulout[48]), .B(acc[48]), .Z(n3330) );
  CNR2X1 U2915 ( .A(mulout[49]), .B(n1162), .Z(n3301) );
  CNR2X1 U2916 ( .A(n3330), .B(n3301), .Z(n2989) );
  CNR2X1 U2917 ( .A(mulout[50]), .B(n1127), .Z(n3563) );
  CNR2X1 U2918 ( .A(mulout[51]), .B(acc[51]), .Z(n3558) );
  CNR2X1 U2919 ( .A(n3563), .B(n3558), .Z(n2488) );
  CND2X1 U2920 ( .A(n2989), .B(n2488), .Z(n2490) );
  CNR2X1 U2921 ( .A(n3304), .B(n2490), .Z(n3265) );
  CIVX1 U2922 ( .A(n3265), .Z(n3586) );
  CNR2X1 U2923 ( .A(mulout[52]), .B(acc[52]), .Z(n2636) );
  CNR2X1 U2924 ( .A(n3586), .B(n2636), .Z(n2492) );
  CNR2X1 U2925 ( .A(n2455), .B(n2458), .Z(n3115) );
  CNR2X1 U2926 ( .A(acc[30]), .B(mulout[30]), .Z(n3109) );
  CNR2X1 U2927 ( .A(acc[31]), .B(mulout[31]), .Z(n3041) );
  CNR2X1 U2928 ( .A(n3109), .B(n3041), .Z(n2460) );
  CND2X1 U2929 ( .A(n3115), .B(n2460), .Z(n2462) );
  CNR2X1 U2930 ( .A(n3195), .B(n2462), .Z(n2464) );
  CND2XL U2931 ( .A(n2456), .B(n2464), .Z(n2468) );
  COND1XL U2932 ( .A(n3192), .B(n2458), .C(n2457), .Z(n3113) );
  CND2X1 U2933 ( .A(acc[30]), .B(mulout[30]), .Z(n3110) );
  CND2X1 U2934 ( .A(acc[31]), .B(mulout[31]), .Z(n3042) );
  COND1XL U2935 ( .A(n3110), .B(n3041), .C(n3042), .Z(n2459) );
  CANR1XL U2936 ( .A(n3113), .B(n2460), .C(n2459), .Z(n2461) );
  COND1XL U2937 ( .A(n2462), .B(n3194), .C(n2461), .Z(n2463) );
  CANR1X1 U2938 ( .A(n2465), .B(n2464), .C(n2463), .Z(n2466) );
  COND1X1 U2939 ( .A(n2468), .B(n2467), .C(n2466), .Z(n2540) );
  CNR2X1 U2940 ( .A(mulout[43]), .B(acc[43]), .Z(n2543) );
  CNR2X1 U2941 ( .A(mulout[42]), .B(n1072), .Z(n3542) );
  CNR2X1 U2942 ( .A(n2543), .B(n3542), .Z(n2480) );
  CNR2X1 U2943 ( .A(mulout[41]), .B(acc[41]), .Z(n2891) );
  CNR2X1 U2944 ( .A(mulout[40]), .B(n1166), .Z(n2887) );
  CNR2X1 U2945 ( .A(n2891), .B(n2887), .Z(n3539) );
  CND2X1 U2946 ( .A(n2480), .B(n3539), .Z(n2482) );
  COR2X1 U2947 ( .A(mulout[36]), .B(acc[36]), .Z(n3065) );
  COR2X1 U2948 ( .A(mulout[37]), .B(acc[37]), .Z(n3069) );
  CND2X1 U2949 ( .A(n3065), .B(n3069), .Z(n2871) );
  COR2X1 U2950 ( .A(mulout[38]), .B(acc[38]), .Z(n3613) );
  COR2X1 U2951 ( .A(mulout[39]), .B(acc[39]), .Z(n3616) );
  CND2X1 U2952 ( .A(n3613), .B(n3616), .Z(n2476) );
  CNR2X1 U2953 ( .A(n2871), .B(n2476), .Z(n2478) );
  COR2X1 U2954 ( .A(mulout[34]), .B(acc[34]), .Z(n2782) );
  COR2X1 U2955 ( .A(mulout[35]), .B(acc[35]), .Z(n2784) );
  CND2X1 U2956 ( .A(n2782), .B(n2784), .Z(n2473) );
  COR2X1 U2957 ( .A(mulout[33]), .B(acc[33]), .Z(n2693) );
  CNR2X1 U2958 ( .A(acc[32]), .B(mulout[32]), .Z(n2691) );
  CIVX2 U2959 ( .A(n2691), .Z(n3515) );
  CND2X1 U2960 ( .A(n2693), .B(n3515), .Z(n2777) );
  CNR2X1 U2961 ( .A(n2473), .B(n2777), .Z(n3062) );
  CND2X1 U2962 ( .A(n2478), .B(n3062), .Z(n3004) );
  CNR2X1 U2963 ( .A(n2482), .B(n3004), .Z(n2484) );
  CND2X1 U2964 ( .A(acc[32]), .B(mulout[32]), .Z(n3514) );
  CIVXL U2965 ( .A(n3514), .Z(n2470) );
  CND2X1 U2966 ( .A(mulout[33]), .B(acc[33]), .Z(n2692) );
  CIVX1 U2967 ( .A(n2692), .Z(n2469) );
  CANR1X1 U2968 ( .A(n2470), .B(n2693), .C(n2469), .Z(n2779) );
  CND2X1 U2969 ( .A(mulout[34]), .B(acc[34]), .Z(n2596) );
  CIVXL U2970 ( .A(n2596), .Z(n2780) );
  CND2X1 U2971 ( .A(mulout[35]), .B(acc[35]), .Z(n2783) );
  CIVXL U2972 ( .A(n2783), .Z(n2471) );
  CANR1XL U2973 ( .A(n2780), .B(n2784), .C(n2471), .Z(n2472) );
  CND2X1 U2974 ( .A(mulout[36]), .B(acc[36]), .Z(n2972) );
  CIVXL U2975 ( .A(n2972), .Z(n3063) );
  CND2X1 U2976 ( .A(mulout[37]), .B(acc[37]), .Z(n3068) );
  CND2X1 U2977 ( .A(mulout[38]), .B(acc[38]), .Z(n2872) );
  CIVXL U2978 ( .A(n2872), .Z(n3611) );
  CND2X1 U2979 ( .A(mulout[39]), .B(acc[39]), .Z(n3615) );
  CIVXL U2980 ( .A(n3615), .Z(n2474) );
  CANR1XL U2981 ( .A(n3611), .B(n3616), .C(n2474), .Z(n2475) );
  COND1XL U2982 ( .A(n2476), .B(n2870), .C(n2475), .Z(n2477) );
  CANR1X1 U2983 ( .A(n3064), .B(n2478), .C(n2477), .Z(n3003) );
  CND2X1 U2984 ( .A(mulout[40]), .B(n1166), .Z(n3005) );
  CND2X1 U2985 ( .A(mulout[41]), .B(acc[41]), .Z(n2892) );
  COND1X1 U2986 ( .A(n3005), .B(n2891), .C(n2892), .Z(n3537) );
  CND2X1 U2987 ( .A(mulout[42]), .B(n1072), .Z(n3543) );
  CND2X1 U2988 ( .A(mulout[43]), .B(acc[43]), .Z(n2544) );
  COND1XL U2989 ( .A(n3543), .B(n2543), .C(n2544), .Z(n2479) );
  CANR1XL U2990 ( .A(n3537), .B(n2480), .C(n2479), .Z(n2481) );
  COND1X1 U2991 ( .A(n3003), .B(n2482), .C(n2481), .Z(n2483) );
  CANR1X1 U2992 ( .A(n2540), .B(n2484), .C(n2483), .Z(n2648) );
  CIVX2 U2993 ( .A(n2648), .Z(n3591) );
  CND2X1 U2994 ( .A(mulout[44]), .B(acc[44]), .Z(n2624) );
  CND2X1 U2995 ( .A(mulout[45]), .B(n858), .Z(n2575) );
  COND1X1 U2996 ( .A(n2624), .B(n2574), .C(n2575), .Z(n3344) );
  CND2X1 U2997 ( .A(mulout[46]), .B(acc[46]), .Z(n3345) );
  CND2X1 U2998 ( .A(mulout[47]), .B(acc[47]), .Z(n3342) );
  COND1XL U2999 ( .A(n3345), .B(n3341), .C(n3342), .Z(n2485) );
  CANR1X1 U3000 ( .A(n3344), .B(n2486), .C(n2485), .Z(n3305) );
  CND2X1 U3001 ( .A(mulout[48]), .B(acc[48]), .Z(n3331) );
  CND2X1 U3002 ( .A(mulout[49]), .B(n1162), .Z(n3302) );
  COND1XL U3003 ( .A(n3331), .B(n3301), .C(n3302), .Z(n2988) );
  CND2X1 U3004 ( .A(mulout[50]), .B(n1127), .Z(n3561) );
  CND2XL U3005 ( .A(mulout[51]), .B(acc[51]), .Z(n3559) );
  COND1XL U3006 ( .A(n3561), .B(n3558), .C(n3559), .Z(n2487) );
  CANR1XL U3007 ( .A(n2988), .B(n2488), .C(n2487), .Z(n2489) );
  COND1X1 U3008 ( .A(n2490), .B(n3305), .C(n2489), .Z(n3264) );
  CIVX1 U3009 ( .A(n3264), .Z(n3588) );
  CND2X1 U3010 ( .A(mulout[52]), .B(acc[52]), .Z(n3262) );
  CANR1X1 U3011 ( .A(n2492), .B(n3591), .C(n2491), .Z(n2493) );
  CAN2X1 U3012 ( .A(n2495), .B(cmd_2[0]), .Z(n3620) );
  COR2X1 U3013 ( .A(n2498), .B(n2497), .Z(n2500) );
  CND3X1 U3014 ( .A(n2503), .B(n2502), .C(n2501), .Z(n516) );
  CNR2IX2 U3015 ( .B(n2505), .A(n1132), .Z(n2686) );
  CNR2X2 U3016 ( .A(n711), .B(n2670), .Z(n3525) );
  CND3X1 U3017 ( .A(n2686), .B(n2586), .C(n3525), .Z(n3413) );
  CIVX2 U3018 ( .A(n3413), .Z(n3357) );
  CIVXL U3019 ( .A(n3366), .Z(n2510) );
  CND2XL U3020 ( .A(n2510), .B(n3364), .Z(n2512) );
  CIVXL U3021 ( .A(n3363), .Z(n3091) );
  CIVXL U3022 ( .A(n3365), .Z(n3093) );
  CANR1XL U3023 ( .A(n3091), .B(n3504), .C(n3093), .Z(n2511) );
  CEOXL U3024 ( .A(n2512), .B(n2511), .Z(n2513) );
  CND2IXL U3025 ( .B(n2701), .A(n2513), .Z(n2515) );
  CANR2XL U3026 ( .A(n1659), .B(mulout[20]), .C(acc[20]), .D(n3617), .Z(n2514)
         );
  CND2X1 U3027 ( .A(n2515), .B(n2514), .Z(n2516) );
  CNR2X1 U3028 ( .A(n3359), .B(n3325), .Z(n2518) );
  CND2X2 U3029 ( .A(n2031), .B(n2523), .Z(n2551) );
  CIVX4 U3030 ( .A(n2551), .Z(n2588) );
  CEOX1 U3031 ( .A(n2849), .B(n3002), .Z(n2536) );
  CANR2XL U3032 ( .A(n1659), .B(mulout[15]), .C(acc[15]), .D(n3617), .Z(n2524)
         );
  CIVX1 U3033 ( .A(n2527), .Z(n3380) );
  CND2XL U3034 ( .A(n2528), .B(n2531), .Z(n2533) );
  CANR1XL U3035 ( .A(n2531), .B(n2530), .C(n2529), .Z(n2532) );
  CND2XL U3036 ( .A(n2534), .B(n3620), .Z(n2535) );
  COND3X1 U3037 ( .A(n2536), .B(n3325), .C(n721), .D(n2535), .Z(n554) );
  CNIVXL U3038 ( .A(q0[29]), .Z(n2537) );
  CMX2XL U3039 ( .A0(n2537), .A1(q[29]), .S(n3624), .Z(n599) );
  CNIVXL U3040 ( .A(q0[9]), .Z(n2538) );
  CMX2XL U3041 ( .A0(n2538), .A1(q[9]), .S(n3624), .Z(n579) );
  CIVX4 U3042 ( .A(rst), .Z(n3629) );
  CIVX2 U3043 ( .A(n2540), .Z(n3614) );
  CIVXL U3044 ( .A(n3539), .Z(n2541) );
  CIVXL U3045 ( .A(n3004), .Z(n3536) );
  CIVXL U3046 ( .A(n3003), .Z(n3538) );
  CIVXL U3047 ( .A(n3537), .Z(n2542) );
  CNR2IXL U3048 ( .B(acc[43]), .A(n3580), .Z(n2545) );
  CANR1XL U3049 ( .A(n1659), .B(mulout[43]), .C(n2545), .Z(n2546) );
  CND2XL U3050 ( .A(n2547), .B(n2546), .Z(n2567) );
  CIVX2 U3051 ( .A(n2572), .Z(n2563) );
  CNR2X2 U3052 ( .A(n2554), .B(n2553), .Z(n2593) );
  CNR2X2 U3053 ( .A(n2555), .B(n3101), .Z(n2559) );
  CIVX2 U3054 ( .A(n1184), .Z(n3102) );
  CNR2X2 U3055 ( .A(n2557), .B(n2556), .Z(n2558) );
  CND3X2 U3056 ( .A(n2559), .B(n3102), .C(n2558), .Z(n2560) );
  COND1XL U3057 ( .A(n2572), .B(n2568), .C(n3269), .Z(n2562) );
  CANR1XL U3058 ( .A(n2563), .B(n1105), .C(n2562), .Z(n2564) );
  CND2X1 U3059 ( .A(n2565), .B(n2564), .Z(n2566) );
  CND2IX1 U3060 ( .B(n2567), .A(n2566), .Z(n526) );
  CND2X1 U3061 ( .A(n2631), .B(n2572), .Z(n2766) );
  CIVX2 U3062 ( .A(n3129), .Z(n3526) );
  CND3X1 U3063 ( .A(n3526), .B(n2568), .C(n3525), .Z(n2573) );
  CNR2X1 U3064 ( .A(n2569), .B(n2763), .Z(n2769) );
  CAN2X1 U3065 ( .A(n2769), .B(n3269), .Z(n2570) );
  COND11X2 U3066 ( .A(n2766), .B(n3015), .C(n2573), .D(n2570), .Z(n2571) );
  CIVXL U3067 ( .A(n2769), .Z(n2765) );
  CIVX2 U3068 ( .A(n2573), .Z(n2630) );
  CIVX2 U3069 ( .A(n3015), .Z(n2629) );
  CND2X2 U3070 ( .A(n2630), .B(n2629), .Z(n2774) );
  CIVX1 U3071 ( .A(n2576), .Z(n2625) );
  CND2IX1 U3072 ( .B(n2579), .A(n2578), .Z(n524) );
  CNIVX1 U3073 ( .A(n2580), .Z(n2689) );
  CND2XL U3074 ( .A(n2689), .B(n3269), .Z(n2699) );
  CIVXL U3075 ( .A(n2699), .Z(n2688) );
  CND2X2 U3076 ( .A(n2586), .B(n2585), .Z(n2587) );
  CIVX2 U3077 ( .A(n2587), .Z(n3524) );
  CND2X2 U3078 ( .A(n2588), .B(n3524), .Z(n2687) );
  CIVX2 U3079 ( .A(n2687), .Z(n2589) );
  CND3XL U3080 ( .A(n1110), .B(n1176), .C(n2689), .Z(n2591) );
  CIVX2 U3081 ( .A(n3513), .Z(n3511) );
  CNR2X1 U3082 ( .A(n2591), .B(n3511), .Z(n2592) );
  CND3X1 U3083 ( .A(n1141), .B(n2593), .C(n2592), .Z(n2786) );
  CIVX2 U3084 ( .A(n1105), .Z(n2594) );
  CND2IX2 U3085 ( .B(n2786), .A(n2594), .Z(n3085) );
  CND2XL U3086 ( .A(n2595), .B(n3085), .Z(n2601) );
  CANR1XL U3087 ( .A(n3595), .B(n2599), .C(n2598), .Z(n2600) );
  CND2XL U3088 ( .A(n2601), .B(n2600), .Z(n535) );
  CND2XL U3089 ( .A(n1112), .B(n3269), .Z(n2602) );
  CND2IXL U3090 ( .B(n2602), .A(n3280), .Z(n2606) );
  CIVX2 U3091 ( .A(n3463), .Z(n3443) );
  CNR2X1 U3092 ( .A(n1064), .B(n2603), .Z(n3464) );
  CNIVXL U3093 ( .A(n2605), .Z(n3373) );
  CNR2X2 U3094 ( .A(n3372), .B(n3373), .Z(n3288) );
  CIVDXL U3095 ( .A(n1099), .Z0(n3280), .Z1(n3287) );
  CIVXL U3096 ( .A(n2608), .Z(n2609) );
  CND2XL U3097 ( .A(n2609), .B(n3269), .Z(n2618) );
  CIVXL U3098 ( .A(n2618), .Z(n2610) );
  CIVXL U3099 ( .A(n2611), .Z(n2614) );
  CIVXL U3100 ( .A(n2612), .Z(n2613) );
  COND1XL U3101 ( .A(n2614), .B(n3452), .C(n2613), .Z(n2911) );
  CIVX1 U3102 ( .A(n2615), .Z(n2912) );
  CND2XL U3103 ( .A(n2912), .B(n2910), .Z(n2616) );
  CENX1 U3104 ( .A(n2911), .B(n2616), .Z(n2617) );
  CND2XL U3105 ( .A(n2617), .B(n3620), .Z(n2620) );
  CIVXL U3106 ( .A(n3373), .Z(n3281) );
  CNR2IXL U3107 ( .B(n2620), .A(n2619), .Z(n2621) );
  CNR2XL U3108 ( .A(n3632), .B(n3580), .Z(n2626) );
  CANR1XL U3109 ( .A(n1659), .B(mulout[44]), .C(n2626), .Z(n2627) );
  CND2XL U3110 ( .A(n2628), .B(n2627), .Z(n2634) );
  CND2XL U3111 ( .A(n2631), .B(n3269), .Z(n2632) );
  CND2IXL U3112 ( .B(n2634), .A(n2633), .Z(n525) );
  CNR2X1 U3113 ( .A(mulout[59]), .B(n1065), .Z(n2723) );
  CIVXL U3114 ( .A(n2723), .Z(n2635) );
  CND2X1 U3115 ( .A(mulout[59]), .B(n1065), .Z(n2721) );
  CND2XL U3116 ( .A(n2635), .B(n2721), .Z(n2654) );
  COR2X1 U3117 ( .A(mulout[57]), .B(acc[57]), .Z(n2946) );
  COR2X1 U3118 ( .A(mulout[58]), .B(acc[58]), .Z(n2757) );
  CND2X1 U3119 ( .A(n2946), .B(n2757), .Z(n2720) );
  CIVXL U3120 ( .A(n2720), .Z(n2652) );
  CNR2X1 U3121 ( .A(mulout[55]), .B(acc[55]), .Z(n3417) );
  CNR2X1 U3122 ( .A(mulout[56]), .B(n1108), .Z(n2797) );
  CNR2X1 U3123 ( .A(n3417), .B(n2797), .Z(n2642) );
  CNR2X1 U3124 ( .A(mulout[54]), .B(n1088), .Z(n2800) );
  CIVX2 U3125 ( .A(n2800), .Z(n3585) );
  CND2X1 U3126 ( .A(n2642), .B(n3585), .Z(n2644) );
  CIVX2 U3127 ( .A(n2636), .Z(n3263) );
  CND2X1 U3128 ( .A(n3263), .B(n2639), .Z(n3589) );
  CNR2X1 U3129 ( .A(n2644), .B(n3589), .Z(n2646) );
  CND2XL U3130 ( .A(n3265), .B(n2646), .Z(n2649) );
  CIVXL U3131 ( .A(n3262), .Z(n2640) );
  CIVX1 U3132 ( .A(n2637), .Z(n2638) );
  CANR1X1 U3133 ( .A(n2640), .B(n2639), .C(n2638), .Z(n3587) );
  CND2X1 U3134 ( .A(mulout[54]), .B(n1088), .Z(n3584) );
  CIVXL U3135 ( .A(n3584), .Z(n3421) );
  CND2X1 U3136 ( .A(mulout[55]), .B(acc[55]), .Z(n3418) );
  CND2X1 U3137 ( .A(mulout[56]), .B(n1108), .Z(n2798) );
  COND1XL U3138 ( .A(n3418), .B(n2797), .C(n2798), .Z(n2641) );
  CANR1XL U3139 ( .A(n3421), .B(n2642), .C(n2641), .Z(n2643) );
  COND1XL U3140 ( .A(n3587), .B(n2644), .C(n2643), .Z(n2645) );
  CANR1X1 U3141 ( .A(n2646), .B(n3264), .C(n2645), .Z(n2647) );
  COND1X1 U3142 ( .A(n2649), .B(n2648), .C(n2647), .Z(n3240) );
  CND2X1 U3143 ( .A(mulout[57]), .B(acc[57]), .Z(n2945) );
  CIVX2 U3144 ( .A(n2945), .Z(n2758) );
  CND2X1 U3145 ( .A(mulout[58]), .B(acc[58]), .Z(n2756) );
  CIVXL U3146 ( .A(n2756), .Z(n2650) );
  CANR1X1 U3147 ( .A(n2757), .B(n2758), .C(n2650), .Z(n2722) );
  CIVX1 U3148 ( .A(n2722), .Z(n2651) );
  CANR1X1 U3149 ( .A(n2652), .B(n3240), .C(n2651), .Z(n2653) );
  CEOXL U3150 ( .A(n2654), .B(n2653), .Z(n2655) );
  CAN2XL U3151 ( .A(n2655), .B(n3620), .Z(n2657) );
  CNR2XL U3152 ( .A(n2657), .B(n2656), .Z(n2685) );
  CIVX2 U3153 ( .A(n2658), .Z(n2668) );
  CIVX2 U3154 ( .A(n2659), .Z(n2667) );
  CND2X1 U3155 ( .A(n2660), .B(n3573), .Z(n3431) );
  CND2X1 U3156 ( .A(n2661), .B(n2979), .Z(n2949) );
  CND2X1 U3157 ( .A(n2662), .B(n2671), .Z(n2943) );
  CND2XL U3158 ( .A(n3574), .B(n3571), .Z(n2747) );
  CND2XL U3159 ( .A(n2663), .B(n2979), .Z(n2750) );
  CNR2X1 U3160 ( .A(n2665), .B(n2746), .Z(n2666) );
  CND3X2 U3161 ( .A(n2668), .B(n2667), .C(n2666), .Z(n3025) );
  CND2X1 U3162 ( .A(n2672), .B(n2671), .Z(n3162) );
  CIVX1 U3163 ( .A(n3162), .Z(n3155) );
  CND2XL U3164 ( .A(n3155), .B(n1188), .Z(n2673) );
  CNR2XL U3165 ( .A(n2673), .B(n3025), .Z(n2679) );
  CND3X1 U3166 ( .A(n2793), .B(n2794), .C(n2792), .Z(n3023) );
  CNR3X2 U3167 ( .A(n2676), .B(n2675), .C(n1103), .Z(n2677) );
  CND2X2 U3168 ( .A(n2677), .B(n3521), .Z(n3022) );
  CIVX2 U3169 ( .A(n3022), .Z(n3030) );
  CNR2XL U3170 ( .A(n1154), .B(n2745), .Z(n2678) );
  CND2XL U3171 ( .A(n2679), .B(n2678), .Z(n2683) );
  CIVX2 U3172 ( .A(n2743), .Z(n3031) );
  CND2XL U3173 ( .A(n3031), .B(n1168), .Z(n2680) );
  CANR1XL U3174 ( .A(n3162), .B(n3025), .C(n3325), .Z(n2681) );
  CND3XL U3175 ( .A(n2683), .B(n2682), .C(n2681), .Z(n2684) );
  CND2XL U3176 ( .A(n2684), .B(n2685), .Z(n510) );
  CND2X1 U3177 ( .A(n1176), .B(n3269), .Z(n3520) );
  CNR2XL U3178 ( .A(n3520), .B(n2689), .Z(n2703) );
  CIVX2 U3179 ( .A(n2690), .Z(n3058) );
  CIVXL U3180 ( .A(n3595), .Z(n2701) );
  COND1XL U3181 ( .A(n2691), .B(n3614), .C(n3514), .Z(n2695) );
  CND2X1 U3182 ( .A(n2693), .B(n2692), .Z(n2694) );
  CNR2XL U3183 ( .A(n2696), .B(n3580), .Z(n2697) );
  CANR1XL U3184 ( .A(mulout[33]), .B(n1659), .C(n2697), .Z(n2698) );
  COAN1XL U3185 ( .A(n1176), .B(n2699), .C(n2698), .Z(n2700) );
  COND1XL U3186 ( .A(n2701), .B(n1209), .C(n2700), .Z(n2702) );
  CND2X1 U3187 ( .A(n2705), .B(n2704), .Z(n536) );
  CNR2X1 U3188 ( .A(n3248), .B(n2706), .Z(n2712) );
  CND2XL U3189 ( .A(n2707), .B(n2712), .Z(n3159) );
  CND2X1 U3190 ( .A(n2708), .B(n2712), .Z(n3158) );
  CNR3XL U3191 ( .A(n3162), .B(n3159), .C(n3158), .Z(n2709) );
  CAN2XL U3192 ( .A(n3021), .B(n2709), .Z(n2710) );
  CND2X1 U3193 ( .A(n2710), .B(n2711), .Z(n3246) );
  CIVX1 U3194 ( .A(n3246), .Z(n2715) );
  CND2XL U3195 ( .A(n2713), .B(n2712), .Z(n3245) );
  CND2X1 U3196 ( .A(n2715), .B(n2714), .Z(n2718) );
  CANR1XL U3197 ( .A(n3245), .B(n3025), .C(n3531), .Z(n2717) );
  CND2XL U3198 ( .A(n3246), .B(n3245), .Z(n2716) );
  CND3X1 U3199 ( .A(n2718), .B(n2717), .C(n2716), .Z(n2731) );
  CNR2X1 U3200 ( .A(mulout[62]), .B(acc[62]), .Z(n3238) );
  CIVXL U3201 ( .A(n3238), .Z(n2719) );
  CND2X1 U3202 ( .A(mulout[62]), .B(acc[62]), .Z(n3236) );
  CNR2X1 U3203 ( .A(n2720), .B(n2723), .Z(n3172) );
  CNR2X1 U3204 ( .A(mulout[60]), .B(n1180), .Z(n3176) );
  CNR2X1 U3205 ( .A(mulout[61]), .B(n1080), .Z(n3169) );
  CNR2X1 U3206 ( .A(n3176), .B(n3169), .Z(n2724) );
  CND2XL U3207 ( .A(n3172), .B(n2724), .Z(n3235) );
  CIVX1 U3208 ( .A(n3235), .Z(n2726) );
  COND1X1 U3209 ( .A(n2723), .B(n2722), .C(n2721), .Z(n3173) );
  CND2X1 U3210 ( .A(mulout[60]), .B(n1180), .Z(n3174) );
  CND2X1 U3211 ( .A(mulout[61]), .B(n1080), .Z(n3170) );
  CIVX1 U3212 ( .A(n3237), .Z(n2725) );
  CANR1X1 U3213 ( .A(n2726), .B(n3240), .C(n2725), .Z(n2727) );
  CNR2IX1 U3214 ( .B(acc[62]), .A(n3580), .Z(n2728) );
  CANR1XL U3215 ( .A(n1659), .B(mulout[62]), .C(n2728), .Z(n2729) );
  CND2X1 U3216 ( .A(n2731), .B(n1205), .Z(n507) );
  CENXL U3217 ( .A(n3359), .B(n3413), .Z(n2738) );
  CANR1XL U3218 ( .A(n3620), .B(n2736), .C(n2735), .Z(n2737) );
  CIVXL U3219 ( .A(n3025), .Z(n2742) );
  CND2XL U3220 ( .A(mulout[58]), .B(n1659), .Z(n2739) );
  COND1XL U3221 ( .A(n3580), .B(n2740), .C(n2739), .Z(n2752) );
  CIVXL U3222 ( .A(n2752), .Z(n2741) );
  CNR2XL U3223 ( .A(n3554), .B(n2745), .Z(n2755) );
  CNR2X2 U3224 ( .A(n2746), .B(n3271), .Z(n3572) );
  CND2XL U3225 ( .A(n2748), .B(n3269), .Z(n2749) );
  CNR3XL U3226 ( .A(n2977), .B(n2937), .C(n2749), .Z(n2754) );
  CNR2XL U3227 ( .A(n2750), .B(n3325), .Z(n2751) );
  COR2XL U3228 ( .A(n2752), .B(n2751), .Z(n2753) );
  CANR1XL U3229 ( .A(n2755), .B(n2754), .C(n2753), .Z(n2761) );
  CND2XL U3230 ( .A(n2759), .B(n3595), .Z(n2760) );
  CNR2XL U3231 ( .A(n2764), .B(n2763), .Z(n2767) );
  COR4X1 U3232 ( .A(n2767), .B(n3325), .C(n2766), .D(n2765), .Z(n2775) );
  CND2X1 U3233 ( .A(n2767), .B(n3269), .Z(n2768) );
  CIVXL U3234 ( .A(n3346), .Z(n2770) );
  CNR2IX1 U3235 ( .B(n2771), .A(n1207), .Z(n2772) );
  COND3X1 U3236 ( .A(n2775), .B(n2774), .C(n2773), .D(n2772), .Z(n523) );
  CIVXL U3237 ( .A(n3061), .Z(n2787) );
  CIVXL U3238 ( .A(n2777), .Z(n2778) );
  CIVXL U3239 ( .A(n2779), .Z(n2781) );
  CND2IXL U3240 ( .B(n3061), .A(n3002), .Z(n2788) );
  CND3XL U3241 ( .A(n2790), .B(n2789), .C(n2788), .Z(n534) );
  CIVX2 U3242 ( .A(n2949), .Z(n2939) );
  CNR2XL U3243 ( .A(n2939), .B(n3531), .Z(n2791) );
  CAN3XL U3244 ( .A(n2792), .B(n2505), .C(n2794), .Z(n2795) );
  CND2IX1 U3245 ( .B(n3022), .A(n2795), .Z(n3350) );
  CIVX2 U3246 ( .A(n3350), .Z(n2796) );
  CND2X2 U3247 ( .A(n2796), .B(n3551), .Z(n3577) );
  CIVX2 U3248 ( .A(n3577), .Z(n3575) );
  CIVXL U3249 ( .A(n2797), .Z(n2799) );
  CND2XL U3250 ( .A(n2799), .B(n2798), .Z(n2808) );
  CNR2X1 U3251 ( .A(n2800), .B(n3417), .Z(n2802) );
  CIVX1 U3252 ( .A(n3589), .Z(n3420) );
  CND2X1 U3253 ( .A(n2802), .B(n3420), .Z(n2804) );
  CNR2XL U3254 ( .A(n3586), .B(n2804), .Z(n2806) );
  CIVXL U3255 ( .A(n3587), .Z(n3422) );
  COND1XL U3256 ( .A(n3584), .B(n3417), .C(n3418), .Z(n2801) );
  CANR1XL U3257 ( .A(n3422), .B(n2802), .C(n2801), .Z(n2803) );
  COND1XL U3258 ( .A(n2804), .B(n3588), .C(n2803), .Z(n2805) );
  CANR1XL U3259 ( .A(n2806), .B(n3591), .C(n2805), .Z(n2807) );
  CEOXL U3260 ( .A(n2808), .B(n2807), .Z(n2809) );
  CAN2XL U3261 ( .A(n2809), .B(n3620), .Z(n2814) );
  CND2X1 U3262 ( .A(n2939), .B(n3269), .Z(n2815) );
  CNR2XL U3263 ( .A(n1109), .B(n3580), .Z(n2810) );
  CANR1XL U3264 ( .A(n1659), .B(mulout[56]), .C(n2810), .Z(n2811) );
  COND1XL U3265 ( .A(n2815), .B(n2812), .C(n2811), .Z(n2813) );
  CNR2XL U3266 ( .A(n2814), .B(n2813), .Z(n2818) );
  CIVX2 U3267 ( .A(n2815), .Z(n2816) );
  CND2XL U3268 ( .A(n3577), .B(n2816), .Z(n2817) );
  CND3XL U3269 ( .A(n2817), .B(n2819), .C(n2818), .Z(n513) );
  CNR2XL U3270 ( .A(n1186), .B(n2821), .Z(n2822) );
  CIVXL U3271 ( .A(n2835), .Z(n2839) );
  CNR2XL U3272 ( .A(n2825), .B(n2826), .Z(n2827) );
  CNIVXL U3273 ( .A(n2830), .Z(n2831) );
  CIVX1 U3274 ( .A(n3437), .Z(n2836) );
  CIVXL U3275 ( .A(n2832), .Z(n2834) );
  CND2XL U3276 ( .A(n2834), .B(n2833), .Z(n3297) );
  CANR4CX1 U3277 ( .A(n3297), .B(n2836), .C(n2835), .D(n3325), .Z(n2837) );
  CANR2XL U3278 ( .A(n1659), .B(mulout[6]), .C(acc[6]), .D(n3617), .Z(n2840)
         );
  CIVXL U3279 ( .A(n2841), .Z(n3440) );
  CANR1XL U3280 ( .A(n2843), .B(n3440), .C(n2842), .Z(n3466) );
  CND2XL U3281 ( .A(n2844), .B(n3595), .Z(n2845) );
  CND2IXL U3282 ( .B(n2863), .A(n3269), .Z(n2920) );
  CND3X1 U3283 ( .A(n3526), .B(n3525), .C(n2849), .Z(n3500) );
  CIVXL U3284 ( .A(n3500), .Z(n2854) );
  CIVXL U3285 ( .A(n2850), .Z(n2851) );
  CIVX1 U3286 ( .A(n3501), .Z(n2853) );
  CND2X1 U3287 ( .A(n2854), .B(n2853), .Z(n2929) );
  CIVXL U3288 ( .A(n2855), .Z(n2857) );
  CND2XL U3289 ( .A(n2857), .B(n2856), .Z(n2861) );
  CIVX1 U3290 ( .A(n2858), .Z(n3503) );
  CIVXL U3291 ( .A(n3502), .Z(n2859) );
  CANR1XL U3292 ( .A(n3503), .B(n3504), .C(n2859), .Z(n2860) );
  CEOXL U3293 ( .A(n2861), .B(n2860), .Z(n2862) );
  CND2XL U3294 ( .A(n2862), .B(n3595), .Z(n2866) );
  CAOR2XL U3295 ( .A(acc[17]), .B(n3617), .C(n1659), .D(mulout[17]), .Z(n2864)
         );
  CANR4CXL U3296 ( .A(n3501), .B(n3500), .C(n2930), .D(n2864), .Z(n2865) );
  COND3XL U3297 ( .A(n2920), .B(n2929), .C(n2866), .D(n2865), .Z(n552) );
  CIVXL U3298 ( .A(n2874), .Z(n3076) );
  CNR3XL U3299 ( .A(n3076), .B(n2873), .C(n3325), .Z(n2867) );
  CND3XL U3300 ( .A(n2867), .B(n3083), .C(n2967), .Z(n2869) );
  CIVXL U3301 ( .A(n3085), .Z(n2868) );
  CND2IXL U3302 ( .B(n2869), .A(n2868), .Z(n2880) );
  CIVXL U3303 ( .A(n3062), .Z(n2971) );
  CNR2XL U3304 ( .A(n2971), .B(n2871), .Z(n3610) );
  CIVXL U3305 ( .A(n3064), .Z(n2970) );
  COND1XL U3306 ( .A(n2871), .B(n2970), .C(n2870), .Z(n3612) );
  CND2X1 U3307 ( .A(n2873), .B(n3269), .Z(n2877) );
  CNR2X1 U3308 ( .A(n2876), .B(n2875), .Z(n2879) );
  CND2IXL U3309 ( .B(n2877), .A(n3085), .Z(n2878) );
  CND3XL U3310 ( .A(n2880), .B(n2879), .C(n2878), .Z(n531) );
  CIVX1 U3311 ( .A(n2886), .Z(n2902) );
  CND2X1 U3312 ( .A(n2882), .B(n2881), .Z(n3604) );
  CND2X1 U3313 ( .A(n2884), .B(n2883), .Z(n3530) );
  CANR2X1 U3314 ( .A(mulout[41]), .B(n1659), .C(acc[41]), .D(n3617), .Z(n2885)
         );
  COND4CXL U3315 ( .A(n3604), .B(n3530), .C(n2886), .D(n2885), .Z(n2897) );
  CIVX1 U3316 ( .A(n2887), .Z(n3006) );
  CND2XL U3317 ( .A(n3536), .B(n3006), .Z(n2890) );
  CIVXL U3318 ( .A(n3005), .Z(n2888) );
  CANR1XL U3319 ( .A(n3006), .B(n3538), .C(n2888), .Z(n2889) );
  COND1XL U3320 ( .A(n2890), .B(n3614), .C(n2889), .Z(n2894) );
  CENX1 U3321 ( .A(n2894), .B(n2893), .Z(n2895) );
  CND2XL U3322 ( .A(n2895), .B(n3595), .Z(n2896) );
  CND2IXL U3323 ( .B(n2897), .A(n2896), .Z(n2898) );
  CAN2X1 U3324 ( .A(n3530), .B(n3269), .Z(n3014) );
  CIVXL U3325 ( .A(n3604), .Z(n2899) );
  CNR2XL U3326 ( .A(n2899), .B(n3529), .Z(n2900) );
  CND2XL U3327 ( .A(n3014), .B(n2900), .Z(n2901) );
  CNR2XL U3328 ( .A(n3002), .B(n2901), .Z(n2903) );
  CMXI2XL U3329 ( .A0(n2903), .A1(n2902), .S(n1083), .Z(n2904) );
  CNIVXL U3330 ( .A(n2905), .Z(n3446) );
  CNR2X1 U3331 ( .A(n3463), .B(n3448), .Z(n2906) );
  CENXL U3332 ( .A(n3446), .B(n2906), .Z(n2915) );
  CANR2XL U3333 ( .A(n1659), .B(mulout[11]), .C(acc[11]), .D(n3617), .Z(n2907)
         );
  CND2XL U3334 ( .A(n2913), .B(n3620), .Z(n2914) );
  COND3XL U3335 ( .A(n2915), .B(n3531), .C(n844), .D(n2914), .Z(n558) );
  CNIVXL U3336 ( .A(n1157), .Z(n2918) );
  CAN2XL U3337 ( .A(n2931), .B(n3269), .Z(n2923) );
  CIVXL U3338 ( .A(n2931), .Z(n2921) );
  CANR2XL U3339 ( .A(n1659), .B(mulout[18]), .C(acc[18]), .D(n3617), .Z(n2919)
         );
  COND1XL U3340 ( .A(n2921), .B(n2920), .C(n2919), .Z(n2922) );
  CANR1X1 U3341 ( .A(n2923), .B(n2929), .C(n2922), .Z(n2936) );
  CND2XL U3342 ( .A(n2928), .B(n3620), .Z(n2935) );
  CIVXL U3343 ( .A(n2929), .Z(n2933) );
  CND3X1 U3344 ( .A(n2936), .B(n2934), .C(n2935), .Z(n551) );
  CIVXL U3345 ( .A(n3554), .Z(n2938) );
  CNR3X1 U3346 ( .A(n3022), .B(n2977), .C(n2937), .Z(n3432) );
  CND2XL U3347 ( .A(n3432), .B(n2938), .Z(n2944) );
  CIVXL U3348 ( .A(n2944), .Z(n2942) );
  CND3XL U3349 ( .A(n2939), .B(n3269), .C(n1137), .Z(n2940) );
  CND2XL U3350 ( .A(n2942), .B(n2941), .Z(n2960) );
  CNR2X1 U3351 ( .A(n1137), .B(n3325), .Z(n2953) );
  CND2XL U3352 ( .A(n2944), .B(n2953), .Z(n2959) );
  CND2XL U3353 ( .A(n2946), .B(n2945), .Z(n2947) );
  CENXL U3354 ( .A(n3240), .B(n2947), .Z(n2948) );
  CAN2XL U3355 ( .A(n2948), .B(n3595), .Z(n2957) );
  CND2X1 U3356 ( .A(n2953), .B(n2949), .Z(n2950) );
  COND1XL U3357 ( .A(n3580), .B(n2951), .C(n2950), .Z(n2952) );
  CANR1XL U3358 ( .A(n2953), .B(n3431), .C(n2952), .Z(n2955) );
  CND2XL U3359 ( .A(mulout[57]), .B(n1659), .Z(n2954) );
  CND2XL U3360 ( .A(n2955), .B(n2954), .Z(n2956) );
  CNR2XL U3361 ( .A(n2957), .B(n2956), .Z(n2958) );
  CND3XL U3362 ( .A(n2960), .B(n2959), .C(n2958), .Z(n512) );
  CIVXL U3363 ( .A(n2967), .Z(n3075) );
  CNR2IXL U3364 ( .B(n3269), .A(n3075), .Z(n2966) );
  CND3XL U3365 ( .A(n3076), .B(n3269), .C(n2967), .Z(n2964) );
  CNR2XL U3366 ( .A(n2961), .B(n3580), .Z(n2962) );
  CANR1XL U3367 ( .A(mulout[36]), .B(n1659), .C(n2962), .Z(n2963) );
  CND2X1 U3368 ( .A(n2964), .B(n2963), .Z(n2965) );
  CANR1X1 U3369 ( .A(n2966), .B(n3085), .C(n2965), .Z(n2976) );
  CIVXL U3370 ( .A(n3085), .Z(n2969) );
  CNR3XL U3371 ( .A(n3076), .B(n2967), .C(n3325), .Z(n2968) );
  CND2X1 U3372 ( .A(n2969), .B(n2968), .Z(n2975) );
  CND2XL U3373 ( .A(n2973), .B(n3620), .Z(n2974) );
  CND3X1 U3374 ( .A(n2976), .B(n2975), .C(n2974), .Z(n533) );
  CIVX1 U3375 ( .A(n3348), .Z(n3340) );
  CIVXL U3376 ( .A(n2982), .Z(n2980) );
  CND2XL U3377 ( .A(n3321), .B(n2980), .Z(n3001) );
  CND2XL U3378 ( .A(mulout[50]), .B(n1659), .Z(n2981) );
  COND1XL U3379 ( .A(n3326), .B(n2982), .C(n2981), .Z(n2986) );
  CIVXL U3380 ( .A(n3299), .Z(n3320) );
  CNR3XL U3381 ( .A(n3320), .B(n2996), .C(n3325), .Z(n2985) );
  CNR2XL U3382 ( .A(n1125), .B(n3580), .Z(n2984) );
  CNR3XL U3383 ( .A(n2986), .B(n2985), .C(n2984), .Z(n2995) );
  CIVXL U3384 ( .A(n3563), .Z(n2987) );
  CND2XL U3385 ( .A(n2987), .B(n3561), .Z(n2993) );
  CIVXL U3386 ( .A(n3304), .Z(n3333) );
  CND2XL U3387 ( .A(n3333), .B(n2989), .Z(n3560) );
  CIVX1 U3388 ( .A(n3560), .Z(n2991) );
  CIVXL U3389 ( .A(n3305), .Z(n3332) );
  CANR1XL U3390 ( .A(n2989), .B(n3332), .C(n2988), .Z(n3562) );
  CIVXL U3391 ( .A(n3562), .Z(n2990) );
  CANR1XL U3392 ( .A(n2991), .B(n3591), .C(n2990), .Z(n2992) );
  CEOXL U3393 ( .A(n2993), .B(n2992), .Z(n2994) );
  CNR2IX1 U3394 ( .B(n2995), .A(n1208), .Z(n3000) );
  CNR2X1 U3395 ( .A(n3299), .B(n3325), .Z(n2997) );
  CAN3XL U3396 ( .A(n2997), .B(n3326), .C(n2996), .Z(n2998) );
  CNR2IX2 U3397 ( .B(n3604), .A(n3002), .Z(n3016) );
  CIVX1 U3398 ( .A(n3016), .Z(n3013) );
  COND1XL U3399 ( .A(n3004), .B(n3614), .C(n3003), .Z(n3008) );
  CND2X1 U3400 ( .A(n3006), .B(n3005), .Z(n3007) );
  CENX1 U3401 ( .A(n3008), .B(n3007), .Z(n3009) );
  CND2XL U3402 ( .A(n3009), .B(n3595), .Z(n3011) );
  CANR2XL U3403 ( .A(mulout[40]), .B(n1659), .C(n1166), .D(n3617), .Z(n3010)
         );
  CND2X1 U3404 ( .A(n3011), .B(n3010), .Z(n3012) );
  CANR1X1 U3405 ( .A(n3014), .B(n3013), .C(n3012), .Z(n3020) );
  CND2XL U3406 ( .A(n1083), .B(n3014), .Z(n3019) );
  CND2XL U3407 ( .A(n3016), .B(n3017), .Z(n3018) );
  CNR2X1 U3408 ( .A(n3159), .B(n3325), .Z(n3029) );
  CIVXL U3409 ( .A(n3021), .Z(n3024) );
  CND2XL U3410 ( .A(n3162), .B(n3029), .Z(n3026) );
  COND1XL U3411 ( .A(n3580), .B(n1181), .C(n3026), .Z(n3027) );
  CAOR1XL U3412 ( .A(n1659), .B(mulout[60]), .C(n3027), .Z(n3028) );
  CND3X2 U3413 ( .A(n3031), .B(n3255), .C(n1168), .Z(n3156) );
  CIVXL U3414 ( .A(n3159), .Z(n3154) );
  CNR2IXL U3415 ( .B(n3269), .A(n3154), .Z(n3032) );
  CAN2XL U3416 ( .A(n3155), .B(n3032), .Z(n3033) );
  CIVXL U3417 ( .A(n3176), .Z(n3034) );
  CND2XL U3418 ( .A(n3034), .B(n3174), .Z(n3036) );
  CANR1XL U3419 ( .A(n3172), .B(n3240), .C(n3173), .Z(n3035) );
  CEOXL U3420 ( .A(n3036), .B(n3035), .Z(n3037) );
  CND2XL U3421 ( .A(n3037), .B(n3620), .Z(n3038) );
  CND2XL U3422 ( .A(n3040), .B(n3269), .Z(n3059) );
  CIVXL U3423 ( .A(n3041), .Z(n3043) );
  CND2XL U3424 ( .A(n3043), .B(n3042), .Z(n3053) );
  CIVXL U3425 ( .A(n3115), .Z(n3044) );
  CNR2XL U3426 ( .A(n3044), .B(n3109), .Z(n3047) );
  CND2XL U3427 ( .A(n3047), .B(n3112), .Z(n3049) );
  CNR2XL U3428 ( .A(n3483), .B(n3049), .Z(n3051) );
  CIVXL U3429 ( .A(n3113), .Z(n3045) );
  COND1XL U3430 ( .A(n3109), .B(n3045), .C(n3110), .Z(n3046) );
  CANR1XL U3431 ( .A(n3114), .B(n3047), .C(n3046), .Z(n3048) );
  COND1XL U3432 ( .A(n3049), .B(n3489), .C(n3048), .Z(n3050) );
  CANR1XL U3433 ( .A(n3051), .B(n3504), .C(n3050), .Z(n3052) );
  CEOXL U3434 ( .A(n3053), .B(n3052), .Z(n3056) );
  CMX2XL U3435 ( .A0(h1[0]), .A1(n1185), .S(rst), .Z(n498) );
  COR3XL U3436 ( .A(n3061), .B(n3075), .C(n3083), .Z(n3082) );
  CND2XL U3437 ( .A(n3062), .B(n3065), .Z(n3067) );
  CANR1XL U3438 ( .A(n3065), .B(n3064), .C(n3063), .Z(n3066) );
  COND1XL U3439 ( .A(n3067), .B(n3614), .C(n3066), .Z(n3071) );
  CND2X1 U3440 ( .A(n3069), .B(n3068), .Z(n3070) );
  CENX1 U3441 ( .A(n3071), .B(n3070), .Z(n3072) );
  CND2XL U3442 ( .A(n3072), .B(n3595), .Z(n3080) );
  CNR2XL U3443 ( .A(n3073), .B(n3580), .Z(n3074) );
  CANR1XL U3444 ( .A(mulout[37]), .B(n1659), .C(n3074), .Z(n3078) );
  CNR2IX1 U3445 ( .B(n3078), .A(n3077), .Z(n3079) );
  CAN2XL U3446 ( .A(n3080), .B(n3079), .Z(n3081) );
  COAN1X1 U3447 ( .A(n3082), .B(n3085), .C(n3081), .Z(n3087) );
  CAN2XL U3448 ( .A(n3083), .B(n3269), .Z(n3084) );
  CND2XL U3449 ( .A(n3085), .B(n3084), .Z(n3086) );
  CND2X1 U3450 ( .A(n3087), .B(n3086), .Z(n532) );
  CND2XL U3451 ( .A(n3099), .B(n3088), .Z(n3098) );
  CND2XL U3452 ( .A(n3091), .B(n3094), .Z(n3400) );
  CANR1XL U3453 ( .A(n3094), .B(n3093), .C(n3092), .Z(n3401) );
  CAOR2XL U3454 ( .A(n1659), .B(mulout[23]), .C(acc[23]), .D(n3617), .Z(n3095)
         );
  CANR1XL U3455 ( .A(n3620), .B(n3096), .C(n3095), .Z(n3097) );
  COND3XL U3456 ( .A(n3100), .B(n3099), .C(n3098), .D(n3097), .Z(n546) );
  CNR2XL U3457 ( .A(n3478), .B(n3101), .Z(n3105) );
  CND4XL U3458 ( .A(n3105), .B(n3269), .C(n3106), .D(n1117), .Z(n3125) );
  CIVXL U3459 ( .A(n3104), .Z(n3108) );
  CANR2XL U3460 ( .A(n1659), .B(mulout[30]), .C(acc[30]), .D(n3617), .Z(n3103)
         );
  COND4CXL U3461 ( .A(n3106), .B(n3105), .C(n3104), .D(n3103), .Z(n3107) );
  CANR1XL U3462 ( .A(n3108), .B(n3207), .C(n3107), .Z(n3124) );
  CIVX1 U3463 ( .A(n3109), .Z(n3111) );
  CND2X1 U3464 ( .A(n3111), .B(n3110), .Z(n3121) );
  CND2XL U3465 ( .A(n3112), .B(n3115), .Z(n3117) );
  CNR2XL U3466 ( .A(n3483), .B(n3117), .Z(n3119) );
  CANR1XL U3467 ( .A(n3115), .B(n3114), .C(n3113), .Z(n3116) );
  COND1XL U3468 ( .A(n3117), .B(n3489), .C(n3116), .Z(n3118) );
  CANR1XL U3469 ( .A(n3119), .B(n3504), .C(n3118), .Z(n3120) );
  CEOXL U3470 ( .A(n3121), .B(n3120), .Z(n3122) );
  CND2XL U3471 ( .A(n3122), .B(n3595), .Z(n3123) );
  COND3XL U3472 ( .A(n1145), .B(n3125), .C(n3123), .D(n3124), .Z(n539) );
  CND2X1 U3473 ( .A(n3133), .B(n3269), .Z(n3139) );
  CIVX1 U3474 ( .A(n3139), .Z(n3144) );
  CNR2XL U3475 ( .A(n3129), .B(n3128), .Z(n3130) );
  CND2X1 U3476 ( .A(n3130), .B(n1155), .Z(n3229) );
  CNR2XL U3477 ( .A(n3225), .B(n3325), .Z(n3135) );
  CNR2XL U3478 ( .A(n3132), .B(n1134), .Z(n3230) );
  CIVXL U3479 ( .A(n3133), .Z(n3134) );
  CND3XL U3480 ( .A(n3135), .B(n3230), .C(n3134), .Z(n3142) );
  CNR2XL U3481 ( .A(n3136), .B(n3580), .Z(n3137) );
  CANR1XL U3482 ( .A(mulout[26]), .B(n1659), .C(n3137), .Z(n3138) );
  COND1XL U3483 ( .A(n3230), .B(n3139), .C(n3138), .Z(n3140) );
  CANR1XL U3484 ( .A(n3144), .B(n3225), .C(n3140), .Z(n3141) );
  COND1XL U3485 ( .A(n3142), .B(n3229), .C(n3141), .Z(n3143) );
  CIVX1 U3486 ( .A(n3145), .Z(n3487) );
  CND2X1 U3487 ( .A(n3487), .B(n3484), .Z(n3151) );
  CIVXL U3488 ( .A(n3482), .Z(n3147) );
  CNR2XL U3489 ( .A(n3483), .B(n3147), .Z(n3149) );
  CIVXL U3490 ( .A(n3486), .Z(n3146) );
  COND1XL U3491 ( .A(n3147), .B(n3489), .C(n3146), .Z(n3148) );
  CANR1XL U3492 ( .A(n3149), .B(n3504), .C(n3148), .Z(n3150) );
  CEOXL U3493 ( .A(n3151), .B(n3150), .Z(n3152) );
  CND2XL U3494 ( .A(n3152), .B(n3620), .Z(n3153) );
  CAN4X1 U3495 ( .A(n3155), .B(n3154), .C(n3269), .D(n3158), .Z(n3157) );
  CNR2X1 U3496 ( .A(n3158), .B(n3531), .Z(n3167) );
  CND2XL U3497 ( .A(n3167), .B(n3159), .Z(n3160) );
  COND1XL U3498 ( .A(n3580), .B(n1081), .C(n3160), .Z(n3161) );
  CANR1XL U3499 ( .A(n3167), .B(n3162), .C(n3161), .Z(n3164) );
  CND2XL U3500 ( .A(mulout[61]), .B(n1659), .Z(n3163) );
  CND2XL U3501 ( .A(n3164), .B(n3163), .Z(n3165) );
  CNR2X1 U3502 ( .A(n3166), .B(n3165), .Z(n3184) );
  CND2XL U3503 ( .A(n3168), .B(n3167), .Z(n3183) );
  CIVX1 U3504 ( .A(n3169), .Z(n3171) );
  CND2X1 U3505 ( .A(n3171), .B(n3170), .Z(n3180) );
  CIVXL U3506 ( .A(n3173), .Z(n3175) );
  COND1XL U3507 ( .A(n3176), .B(n3175), .C(n3174), .Z(n3177) );
  CANR1XL U3508 ( .A(n3178), .B(n3240), .C(n3177), .Z(n3179) );
  CEOXL U3509 ( .A(n3180), .B(n3179), .Z(n3181) );
  CND2XL U3510 ( .A(n3181), .B(n3595), .Z(n3182) );
  CND3X1 U3511 ( .A(n3184), .B(n3183), .C(n3182), .Z(n508) );
  CNIVX1 U3512 ( .A(n3629), .Z(n3633) );
  CNIVXL U3513 ( .A(n839), .Z(n3185) );
  CMX2XL U3514 ( .A0(n3185), .A1(h[3]), .S(n3624), .Z(n605) );
  CNIVXL U3515 ( .A(n817), .Z(n3186) );
  CMX2XL U3516 ( .A0(n3186), .A1(h[2]), .S(n3624), .Z(n604) );
  CNIVXL U3517 ( .A(n820), .Z(n3187) );
  CMX2XL U3518 ( .A0(n3187), .A1(h[1]), .S(n3624), .Z(n603) );
  CNIVXL U3519 ( .A(n836), .Z(n3188) );
  CMX2XL U3520 ( .A0(n3188), .A1(h[4]), .S(n3624), .Z(n606) );
  CMX2XL U3521 ( .A0(n841), .A1(h[6]), .S(n3624), .Z(n608) );
  CMX2XL U3522 ( .A0(n828), .A1(h[5]), .S(n3624), .Z(n607) );
  CMX2X1 U3523 ( .A0(h1[4]), .A1(n2344), .S(rst), .Z(n502) );
  CIVDX1 U3524 ( .A(n3435), .Z0(n3628), .Z1(n3189) );
  CMX2XL U3525 ( .A0(acc[11]), .A1(z[11]), .S(n3189), .Z(n655) );
  CMX2XL U3526 ( .A0(acc[4]), .A1(z[4]), .S(n3189), .Z(n662) );
  CMX2XL U3527 ( .A0(acc[2]), .A1(z[2]), .S(n3189), .Z(n664) );
  CMX2XL U3528 ( .A0(acc[24]), .A1(z[24]), .S(n3189), .Z(n642) );
  CMX2XL U3529 ( .A0(acc[20]), .A1(z[20]), .S(n3189), .Z(n646) );
  CMX2XL U3530 ( .A0(acc[25]), .A1(z[25]), .S(n3189), .Z(n641) );
  CMX2XL U3531 ( .A0(acc[27]), .A1(z[27]), .S(n3189), .Z(n639) );
  CMX2XL U3532 ( .A0(acc[17]), .A1(z[17]), .S(n3189), .Z(n649) );
  CMX2XL U3533 ( .A0(acc[7]), .A1(z[7]), .S(n3189), .Z(n659) );
  CMX2XL U3534 ( .A0(acc[13]), .A1(z[13]), .S(n3189), .Z(n653) );
  CMX2XL U3535 ( .A0(acc[8]), .A1(z[8]), .S(n3189), .Z(n658) );
  CMX2XL U3536 ( .A0(acc[18]), .A1(z[18]), .S(n3189), .Z(n648) );
  CMX2XL U3537 ( .A0(acc[5]), .A1(z[5]), .S(n3189), .Z(n661) );
  CMX2XL U3538 ( .A0(acc[14]), .A1(z[14]), .S(n3189), .Z(n652) );
  CMX2XL U3539 ( .A0(acc[6]), .A1(z[6]), .S(n3189), .Z(n660) );
  CMX2XL U3540 ( .A0(acc[3]), .A1(z[3]), .S(n3189), .Z(n663) );
  CMX2XL U3541 ( .A0(acc[26]), .A1(z[26]), .S(n3189), .Z(n640) );
  CMX2XL U3542 ( .A0(acc[15]), .A1(z[15]), .S(n3189), .Z(n651) );
  CMX2XL U3543 ( .A0(acc[21]), .A1(z[21]), .S(n3189), .Z(n645) );
  CMX2XL U3544 ( .A0(acc[22]), .A1(z[22]), .S(n3189), .Z(n644) );
  CMX2XL U3545 ( .A0(acc[23]), .A1(z[23]), .S(n3189), .Z(n643) );
  CMX2XL U3546 ( .A0(acc[16]), .A1(z[16]), .S(n3189), .Z(n650) );
  CMX2XL U3547 ( .A0(acc[12]), .A1(z[12]), .S(n3189), .Z(n654) );
  CMX2XL U3548 ( .A0(acc[10]), .A1(z[10]), .S(n3189), .Z(n656) );
  CMX2XL U3549 ( .A0(acc[19]), .A1(z[19]), .S(n3189), .Z(n647) );
  CMX2XL U3550 ( .A0(acc[9]), .A1(z[9]), .S(n3189), .Z(n657) );
  CNR3XL U3551 ( .A(n3190), .B(n3478), .C(n3325), .Z(n3191) );
  CNR2IXL U3552 ( .B(n3191), .A(n3207), .Z(n3204) );
  CND2X1 U3553 ( .A(n3193), .B(n3192), .Z(n3199) );
  CNR2XL U3554 ( .A(n3483), .B(n3195), .Z(n3197) );
  COND1XL U3555 ( .A(n3195), .B(n3489), .C(n3194), .Z(n3196) );
  CANR1XL U3556 ( .A(n3197), .B(n3504), .C(n3196), .Z(n3198) );
  CEOXL U3557 ( .A(n3199), .B(n3198), .Z(n3200) );
  CND2XL U3558 ( .A(n3200), .B(n3595), .Z(n3202) );
  CANR2XL U3559 ( .A(n1659), .B(mulout[28]), .C(acc[28]), .D(n3617), .Z(n3201)
         );
  CND2X1 U3560 ( .A(n3202), .B(n3201), .Z(n3203) );
  CNR2X1 U3561 ( .A(n3204), .B(n3203), .Z(n3209) );
  COND1XL U3562 ( .A(n3478), .B(n3207), .C(n3206), .Z(n3208) );
  CND2X1 U3563 ( .A(n3209), .B(n3208), .Z(n541) );
  CIVXL U3564 ( .A(n3229), .Z(n3211) );
  CNR3XL U3565 ( .A(n3230), .B(n3225), .C(n3325), .Z(n3210) );
  CND2X1 U3566 ( .A(n3211), .B(n3210), .Z(n3232) );
  CNR2XL U3567 ( .A(n3483), .B(n3215), .Z(n3217) );
  COND1XL U3568 ( .A(n3215), .B(n3489), .C(n3214), .Z(n3216) );
  CANR1XL U3569 ( .A(n3217), .B(n3504), .C(n3216), .Z(n3218) );
  CEOXL U3570 ( .A(n3219), .B(n3218), .Z(n3220) );
  CND2XL U3571 ( .A(n3220), .B(n3595), .Z(n3224) );
  CNR2XL U3572 ( .A(n3221), .B(n3580), .Z(n3222) );
  CANR1XL U3573 ( .A(mulout[25]), .B(n1659), .C(n3222), .Z(n3223) );
  CND2XL U3574 ( .A(n3224), .B(n3223), .Z(n3227) );
  CND3XL U3575 ( .A(n3225), .B(n3230), .C(n3269), .Z(n3226) );
  CND2IXL U3576 ( .B(n3227), .A(n3226), .Z(n3228) );
  CANR11XL U3577 ( .A(n3230), .B(n3269), .C(n3229), .D(n3228), .Z(n3231) );
  COR2XL U3578 ( .A(mulout[63]), .B(acc[63]), .Z(n3234) );
  CND2XL U3579 ( .A(mulout[63]), .B(acc[63]), .Z(n3233) );
  CND2XL U3580 ( .A(n3234), .B(n3233), .Z(n3243) );
  CNR2XL U3581 ( .A(n3235), .B(n3238), .Z(n3241) );
  COND1XL U3582 ( .A(n3238), .B(n3237), .C(n3236), .Z(n3239) );
  CANR1XL U3583 ( .A(n3241), .B(n3240), .C(n3239), .Z(n3242) );
  CEOXL U3584 ( .A(n3243), .B(n3242), .Z(n3244) );
  CND2XL U3585 ( .A(n3244), .B(n3595), .Z(n3258) );
  CNR2XL U3586 ( .A(n3245), .B(n3247), .Z(n3256) );
  CIVXL U3587 ( .A(n3246), .Z(n3254) );
  CNR2XL U3588 ( .A(n3248), .B(n3247), .Z(n3249) );
  CANR2XL U3589 ( .A(n3250), .B(n3249), .C(acc[63]), .D(n3617), .Z(n3252) );
  CND2XL U3590 ( .A(mulout[63]), .B(n1659), .Z(n3251) );
  CND2X1 U3591 ( .A(n3252), .B(n3251), .Z(n3253) );
  CANR11X1 U3592 ( .A(n3256), .B(n3255), .C(n3254), .D(n3253), .Z(n3257) );
  CND2X1 U3593 ( .A(n3258), .B(n3257), .Z(n506) );
  CIVXL U3594 ( .A(n3276), .Z(n3260) );
  CNR3XL U3595 ( .A(n3261), .B(n3569), .C(n3325), .Z(n3259) );
  CND2X1 U3596 ( .A(n3260), .B(n3259), .Z(n3279) );
  CAN2XL U3597 ( .A(n3261), .B(n3269), .Z(n3277) );
  CND2X1 U3598 ( .A(n3263), .B(n3262), .Z(n3267) );
  CANR1XL U3599 ( .A(n3265), .B(n3591), .C(n3264), .Z(n3266) );
  CEOXL U3600 ( .A(n3267), .B(n3266), .Z(n3268) );
  CND2XL U3601 ( .A(n3268), .B(n3595), .Z(n3274) );
  CND2X1 U3602 ( .A(n3569), .B(n3269), .Z(n3553) );
  CND2XL U3603 ( .A(n3617), .B(acc[52]), .Z(n3270) );
  COND1XL U3604 ( .A(n3271), .B(n3553), .C(n3270), .Z(n3272) );
  CANR1XL U3605 ( .A(n1659), .B(mulout[52]), .C(n3272), .Z(n3273) );
  CND2X1 U3606 ( .A(n3274), .B(n3273), .Z(n3275) );
  CANR1X1 U3607 ( .A(n3277), .B(n3276), .C(n3275), .Z(n3278) );
  CND2X1 U3608 ( .A(n3279), .B(n3278), .Z(n517) );
  CAN2XL U3609 ( .A(n3280), .B(n3269), .Z(n3286) );
  CANR1X1 U3610 ( .A(n3286), .B(n3285), .C(n3284), .Z(n3291) );
  CND2XL U3611 ( .A(n3287), .B(n3269), .Z(n3289) );
  CND2IX1 U3612 ( .B(n3289), .A(n3288), .Z(n3290) );
  CND2X1 U3613 ( .A(n3291), .B(n3290), .Z(n560) );
  CIVX1 U3614 ( .A(n3294), .Z(n3439) );
  CANR2X1 U3615 ( .A(n1659), .B(mulout[5]), .C(acc[5]), .D(n3617), .Z(n3296)
         );
  CIVXL U3616 ( .A(n3326), .Z(n3311) );
  CNR2X1 U3617 ( .A(n3311), .B(n3325), .Z(n3327) );
  CND2X1 U3618 ( .A(n3327), .B(n3299), .Z(n3300) );
  CNR2X1 U3619 ( .A(n3321), .B(n3300), .Z(n3319) );
  CIVXL U3620 ( .A(n3301), .Z(n3303) );
  CND2XL U3621 ( .A(n3303), .B(n3302), .Z(n3309) );
  CNR2XL U3622 ( .A(n3304), .B(n3330), .Z(n3307) );
  COND1XL U3623 ( .A(n3330), .B(n3305), .C(n3331), .Z(n3306) );
  CANR1XL U3624 ( .A(n3307), .B(n3591), .C(n3306), .Z(n3308) );
  CEOXL U3625 ( .A(n3309), .B(n3308), .Z(n3310) );
  CND2XL U3626 ( .A(n3310), .B(n3595), .Z(n3317) );
  CAN2X1 U3627 ( .A(n1659), .B(mulout[49]), .Z(n3315) );
  COR2XL U3628 ( .A(n3580), .B(n1163), .Z(n3313) );
  CND3XL U3629 ( .A(n3311), .B(n3320), .C(n3269), .Z(n3312) );
  CND2XL U3630 ( .A(n3313), .B(n3312), .Z(n3314) );
  CNR2XL U3631 ( .A(n3315), .B(n3314), .Z(n3316) );
  CND2XL U3632 ( .A(n3317), .B(n3316), .Z(n3318) );
  CND2XL U3633 ( .A(n3320), .B(n3269), .Z(n3322) );
  CND2IXL U3634 ( .B(n3322), .A(n3321), .Z(n3323) );
  CIVX1 U3635 ( .A(n3327), .Z(n3335) );
  CANR2XL U3636 ( .A(mulout[48]), .B(n1659), .C(acc[48]), .D(n3617), .Z(n3328)
         );
  COAN1XL U3637 ( .A(n3335), .B(n3329), .C(n3328), .Z(n3338) );
  CND2XL U3638 ( .A(n3595), .B(n3334), .Z(n3337) );
  CND4X1 U3639 ( .A(n3339), .B(n3338), .C(n3337), .D(n3336), .Z(n521) );
  CAN2XL U3640 ( .A(n3348), .B(n3269), .Z(n3349) );
  CNR2X1 U3641 ( .A(n3359), .B(n3360), .Z(n3405) );
  CND4XL U3642 ( .A(n3357), .B(n3269), .C(n3405), .D(n3402), .Z(n3371) );
  CNR2X1 U3643 ( .A(n3402), .B(n3325), .Z(n3397) );
  CAOR2XL U3644 ( .A(acc[21]), .B(n3617), .C(n1659), .D(mulout[21]), .Z(n3358)
         );
  CANR4CX1 U3645 ( .A(n3360), .B(n3359), .C(n3397), .D(n3358), .Z(n3370) );
  CND2XL U3646 ( .A(n3367), .B(n3620), .Z(n3369) );
  CND4X1 U3647 ( .A(n3371), .B(n3370), .C(n3369), .D(n3368), .Z(n548) );
  CANR2XL U3648 ( .A(n1659), .B(mulout[8]), .C(acc[8]), .D(n3617), .Z(n3374)
         );
  CND2XL U3649 ( .A(n3377), .B(n3595), .Z(n3378) );
  CANR1XL U3650 ( .A(n3383), .B(n3385), .C(n3382), .Z(n3392) );
  CND2XL U3651 ( .A(n1151), .B(n3269), .Z(n3388) );
  CIVXL U3652 ( .A(acc[14]), .Z(n3386) );
  CIVXL U3653 ( .A(n3403), .Z(n3396) );
  CND3XL U3654 ( .A(n3405), .B(n3397), .C(n3396), .Z(n3414) );
  CIVXL U3655 ( .A(n3402), .Z(n3406) );
  CND2X1 U3656 ( .A(n3403), .B(n3269), .Z(n3409) );
  CANR2XL U3657 ( .A(n1659), .B(mulout[22]), .C(acc[22]), .D(n3617), .Z(n3404)
         );
  COND4CX1 U3658 ( .A(n3406), .B(n3405), .C(n3409), .D(n3404), .Z(n3407) );
  CNR2IX1 U3659 ( .B(n3408), .A(n3407), .Z(n3412) );
  CIVX1 U3660 ( .A(n3409), .Z(n3410) );
  CIVXL U3661 ( .A(n3430), .Z(n3416) );
  CANR2XL U3662 ( .A(mulout[55]), .B(n1659), .C(acc[55]), .D(n3617), .Z(n3415)
         );
  CIVXL U3663 ( .A(n3417), .Z(n3419) );
  CND2X1 U3664 ( .A(n3419), .B(n3418), .Z(n3428) );
  CND2XL U3665 ( .A(n3420), .B(n3585), .Z(n3424) );
  CNR2XL U3666 ( .A(n3586), .B(n3424), .Z(n3426) );
  CANR1XL U3667 ( .A(n3585), .B(n3422), .C(n3421), .Z(n3423) );
  COND1XL U3668 ( .A(n3424), .B(n3588), .C(n3423), .Z(n3425) );
  CANR1XL U3669 ( .A(n3426), .B(n3591), .C(n3425), .Z(n3427) );
  CEOXL U3670 ( .A(n3428), .B(n3427), .Z(n3429) );
  CMX2XL U3671 ( .A0(q0[4]), .A1(q[4]), .S(pushin), .Z(n574) );
  CMX2XL U3672 ( .A0(q0[18]), .A1(q[18]), .S(pushin), .Z(n588) );
  CMX2XL U3673 ( .A0(q0[10]), .A1(q[10]), .S(pushin), .Z(n580) );
  CMX2XL U3674 ( .A0(q0[12]), .A1(q[12]), .S(pushin), .Z(n582) );
  CMX2XL U3675 ( .A0(q0[8]), .A1(q[8]), .S(pushin), .Z(n578) );
  CMX2XL U3676 ( .A0(q0[14]), .A1(q[14]), .S(pushin), .Z(n584) );
  CMX2XL U3677 ( .A0(q0[16]), .A1(q[16]), .S(pushin), .Z(n586) );
  CMX2XL U3678 ( .A0(q0[6]), .A1(q[6]), .S(pushin), .Z(n576) );
  CMX2XL U3679 ( .A0(q0[2]), .A1(q[2]), .S(pushin), .Z(n572) );
  CMX2XL U3680 ( .A0(acc[30]), .A1(z[30]), .S(n3435), .Z(n636) );
  CMX2XL U3681 ( .A0(acc[28]), .A1(z[28]), .S(n3435), .Z(n638) );
  CMX2XL U3682 ( .A0(acc[31]), .A1(z[31]), .S(n3435), .Z(n634) );
  CMX2XL U3683 ( .A0(acc[1]), .A1(z[1]), .S(n3435), .Z(n665) );
  CMX2XL U3684 ( .A0(q0[26]), .A1(q[26]), .S(n3624), .Z(n596) );
  CNIVXL U3685 ( .A(h0[0]), .Z(n3436) );
  CMX2XL U3686 ( .A0(n3436), .A1(h[0]), .S(n3624), .Z(n602) );
  CIVXL U3687 ( .A(acc[4]), .Z(n3442) );
  CND2XL U3688 ( .A(n1659), .B(mulout[4]), .Z(n3441) );
  CNR2XL U3689 ( .A(n3443), .B(n3445), .Z(n3462) );
  CND3XL U3690 ( .A(n3444), .B(n3446), .C(n3445), .Z(n3450) );
  COND1XL U3691 ( .A(n3446), .B(n3445), .C(n3269), .Z(n3447) );
  CANR1XL U3692 ( .A(n1102), .B(n3448), .C(n3447), .Z(n3449) );
  COND1XL U3693 ( .A(n3450), .B(n1114), .C(n3449), .Z(n3461) );
  CIVXL U3694 ( .A(acc[12]), .Z(n3457) );
  CND2XL U3695 ( .A(n1659), .B(mulout[12]), .Z(n3456) );
  COND1XL U3696 ( .A(n3580), .B(n3457), .C(n3456), .Z(n3458) );
  CANR1XL U3697 ( .A(n3620), .B(n3459), .C(n3458), .Z(n3460) );
  COND1XL U3698 ( .A(n3462), .B(n3461), .C(n3460), .Z(n557) );
  CEOXL U3699 ( .A(n3464), .B(n3463), .Z(n3477) );
  COND1XL U3700 ( .A(n3467), .B(n3466), .C(n3465), .Z(n3471) );
  CENX1 U3701 ( .A(n3471), .B(n3470), .Z(n3475) );
  CND2XL U3702 ( .A(n1659), .B(mulout[7]), .Z(n3472) );
  COND1XL U3703 ( .A(n3580), .B(n3473), .C(n3472), .Z(n3474) );
  CANR1XL U3704 ( .A(n3620), .B(n3475), .C(n3474), .Z(n3476) );
  COND1XL U3705 ( .A(n3325), .B(n3477), .C(n3476), .Z(n562) );
  CENXL U3706 ( .A(n3478), .B(n3207), .Z(n3499) );
  CIVXL U3707 ( .A(n3479), .Z(n3481) );
  CND2XL U3708 ( .A(n3481), .B(n3480), .Z(n3494) );
  CND2XL U3709 ( .A(n3482), .B(n3487), .Z(n3490) );
  CNR2XL U3710 ( .A(n3483), .B(n3490), .Z(n3492) );
  CIVXL U3711 ( .A(n3484), .Z(n3485) );
  CANR1XL U3712 ( .A(n3487), .B(n3486), .C(n3485), .Z(n3488) );
  COND1XL U3713 ( .A(n3490), .B(n3489), .C(n3488), .Z(n3491) );
  CANR1XL U3714 ( .A(n3492), .B(n3504), .C(n3491), .Z(n3493) );
  CEOXL U3715 ( .A(n3494), .B(n3493), .Z(n3497) );
  CANR1XL U3716 ( .A(n3595), .B(n3497), .C(n3496), .Z(n3498) );
  CENXL U3717 ( .A(n3501), .B(n1159), .Z(n3510) );
  CND2XL U3718 ( .A(n1659), .B(mulout[16]), .Z(n3505) );
  COND1XL U3719 ( .A(n3580), .B(n3506), .C(n3505), .Z(n3507) );
  CANR1XL U3720 ( .A(n3595), .B(n3508), .C(n3507), .Z(n3509) );
  CNR2XL U3721 ( .A(n1176), .B(n3325), .Z(n3512) );
  CNR2IX1 U3722 ( .B(n3512), .A(n3511), .Z(n3517) );
  CANR1X1 U3723 ( .A(n3517), .B(n3519), .C(n3516), .Z(n3518) );
  COND1XL U3724 ( .A(n3520), .B(n3519), .C(n3518), .Z(n537) );
  CND2XL U3725 ( .A(n3528), .B(n3269), .Z(n3527) );
  CAN2XL U3726 ( .A(n1141), .B(n1116), .Z(n3523) );
  CND2X1 U3727 ( .A(n3523), .B(n3524), .Z(n3605) );
  CND2XL U3728 ( .A(n1068), .B(n3525), .Z(n3602) );
  CIVX1 U3729 ( .A(n3602), .Z(n3608) );
  CIVXL U3730 ( .A(n3605), .Z(n3534) );
  CND2XL U3731 ( .A(mulout[42]), .B(n1659), .Z(n3532) );
  COND1XL U3732 ( .A(n3580), .B(n1073), .C(n3532), .Z(n3533) );
  CND2XL U3733 ( .A(n3539), .B(n3536), .Z(n3541) );
  CANR1XL U3734 ( .A(n3539), .B(n3538), .C(n3537), .Z(n3540) );
  COND1XL U3735 ( .A(n3541), .B(n3614), .C(n3540), .Z(n3546) );
  CIVXL U3736 ( .A(n3542), .Z(n3544) );
  CND2X1 U3737 ( .A(n3544), .B(n3543), .Z(n3545) );
  CENX1 U3738 ( .A(n3546), .B(n3545), .Z(n3547) );
  CND2XL U3739 ( .A(n3547), .B(n3620), .Z(n3548) );
  CNR2X1 U3740 ( .A(n3569), .B(n3325), .Z(n3557) );
  CIVXL U3741 ( .A(n3557), .Z(n3552) );
  COR2XL U3742 ( .A(n3552), .B(n3551), .Z(n3568) );
  CNR2XL U3743 ( .A(n3554), .B(n3553), .Z(n3556) );
  CMXI2X1 U3744 ( .A0(n3557), .A1(n3556), .S(n3555), .Z(n3567) );
  CAOR2XL U3745 ( .A(mulout[51]), .B(n1659), .C(acc[51]), .D(n3617), .Z(n3564)
         );
  CANR1XL U3746 ( .A(n3595), .B(n3565), .C(n3564), .Z(n3566) );
  CIVXL U3747 ( .A(n3569), .Z(n3570) );
  CAN3X1 U3748 ( .A(n3572), .B(n1111), .C(n3570), .Z(n3578) );
  CNR2XL U3749 ( .A(n3576), .B(n3325), .Z(n3583) );
  CND2XL U3750 ( .A(n3577), .B(n3583), .Z(n3600) );
  CIVXL U3751 ( .A(n3578), .Z(n3582) );
  CND2XL U3752 ( .A(mulout[54]), .B(n1659), .Z(n3579) );
  COND1XL U3753 ( .A(n3580), .B(n1089), .C(n3579), .Z(n3581) );
  CANR1XL U3754 ( .A(n3583), .B(n3582), .C(n3581), .Z(n3598) );
  CND2X1 U3755 ( .A(n3585), .B(n3584), .Z(n3594) );
  CNR2XL U3756 ( .A(n3586), .B(n3589), .Z(n3592) );
  COND1XL U3757 ( .A(n3589), .B(n3588), .C(n3587), .Z(n3590) );
  CANR1XL U3758 ( .A(n3592), .B(n3591), .C(n3590), .Z(n3593) );
  CEOXL U3759 ( .A(n3594), .B(n3593), .Z(n3596) );
  CND2XL U3760 ( .A(n3596), .B(n3595), .Z(n3597) );
  CAN2XL U3761 ( .A(n3598), .B(n3597), .Z(n3599) );
  CND3XL U3762 ( .A(n3600), .B(n3601), .C(n3599), .Z(n515) );
  CNR2XL U3763 ( .A(n3604), .B(n3325), .Z(n3603) );
  CNR2IXL U3764 ( .B(n3603), .A(n3602), .Z(n3607) );
  CND2XL U3765 ( .A(n3604), .B(n3269), .Z(n3609) );
  CIVX1 U3766 ( .A(n3609), .Z(n3606) );
  CMXI2XL U3767 ( .A0(n3607), .A1(n3606), .S(n3605), .Z(n3623) );
  COR2X1 U3768 ( .A(n3609), .B(n3608), .Z(n3622) );
  CAOR2XL U3769 ( .A(n1659), .B(mulout[39]), .C(acc[39]), .D(n3617), .Z(n3618)
         );
  CANR1XL U3770 ( .A(n3620), .B(n3619), .C(n3618), .Z(n3621) );
  CND3XL U3771 ( .A(n3621), .B(n3622), .C(n3623), .Z(n530) );
  CDLY1XL U3772 ( .A(q0[7]), .Z(n3625) );
  CMX2XL U3773 ( .A0(n3625), .A1(q[7]), .S(n3624), .Z(n577) );
endmodule

