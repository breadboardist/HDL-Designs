
module sqrt64_DW01_add_5 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n13, n27, n28, n29, n30, n31, n32, n33, n34, n35, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n49, n50, n51, n52, n53,
         n54, n55, n56, n61, n62, n63, n64, n65, n68, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n92, n93, n94, n95, n96, n97, n98, n99, n101, n104, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n143, n144, n146, n147, n148,
         n151, n152, n153, n154, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n174, n175, n176,
         n177, n178, n179, n180, n183, n185, n186, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n204,
         n205, n206, n207, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n225, n226, n228, n229, n230, n233, n234,
         n235, n236, n237, n238, n241, n244, n245, n246, n247, n248, n249,
         n258, n262, n263, n264, n265, n266, n270, n273, n274, n279, n280,
         n281, n282, n283, n284, n285, n289, n290, n293, n295, n296, n298,
         n299, n300, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n321, n325, n326, n327, n330, n333, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n347, n348, n351, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n373, n375, n376, n377, n380, n381, n382, n384, n385, n390,
         n392, n393, n394, n395, n396, n399, n400, n401, n402, n403, n404,
         n405, n409, n410, n411, n412, n413, n416, n417, n420, n421, n422,
         n423, n426, n427, n428, n429, n430, n431, n432, n435, n436, n437,
         n440, n442, n443, n445, n446, n447, n448, n457, n458, n459, n460,
         n461, n462, n465, n466, n467, n468, n469, n475, n477, n478, n479,
         n480, n481, n482, n483, n485, n486, n487, n488, n489, n491, n492,
         n493, n498, n501, n502, n505, n508, n509, n510, n512, n513, n514,
         n515, n524, n525, n526, n527, n528, n535, n536, n537, n538, n541,
         n543, n544, n545, n546, n549, n552, n553, n554, n561, n562, n563,
         n567, n574, n576, n581, n583, n584, n585, n586, n587, n588, n590,
         n591, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n607, n608, n609, net13590, net13593, net13619,
         net13644, net13692, net13691, net14013, net14079, net14212, net14374,
         net14373, net14586, net14643, net14657, net14687, net14700, n324,
         n323, n322, n449, net17164, net23257, net26826, n408, n391, n389,
         n388, n383, n372, n352, n346, n308, n306, n304, n242, n332, n309,
         n307, n305, n303, n302, n276, n275, n261, n257, n256, n255, n254,
         n253, n252, n243, n2, n560, n559, n558, n557, net14704, n580, n575,
         n573, n571, net26819, net14691, net14666, n519, n507, n506, n500,
         n470, n455, n453, n451, n569, n565, net14006, net26810, net14198,
         n566, n564, n556, n534, n533, n532, n531, n530, n529, n518, n499,
         n456, n452, n450, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n877, n878, n879;
  assign n68 = A[59];
  assign n111 = A[55];
  assign n131 = A[53];
  assign n193 = A[47];
  assign n213 = A[45];
  assign n299 = A[35];
  assign n340 = A[31];
  assign n360 = A[29];
  assign n446 = A[19];
  assign n485 = A[15];
  assign n567 = A[3];
  assign n576 = A[1];

  COND1X1 U54 ( .A(n117), .B(n77), .C(n78), .Z(n76) );
  CNR2X2 U57 ( .A(n81), .B(n92), .Z(n79) );
  CNR2X2 U61 ( .A(B[58]), .B(A[58]), .Z(n81) );
  CEOX2 U63 ( .A(n92), .B(n93), .Z(SUM[57]) );
  CANR1X1 U75 ( .A(n94), .B(net13691), .C(n95), .Z(n93) );
  CANR1X1 U79 ( .A(n98), .B(n119), .C(n99), .Z(n97) );
  CNR2X2 U84 ( .A(n104), .B(n112), .Z(n98) );
  CNR2X2 U88 ( .A(B[56]), .B(A[56]), .Z(n104) );
  CEOX2 U90 ( .A(n112), .B(n113), .Z(SUM[55]) );
  CND2X2 U106 ( .A(n138), .B(n122), .Z(n116) );
  CANR1X1 U107 ( .A(n143), .B(n122), .C(n123), .Z(n117) );
  CNR2X2 U108 ( .A(n124), .B(n132), .Z(n122) );
  CNR2X2 U112 ( .A(B[54]), .B(A[54]), .Z(n124) );
  CEOX2 U138 ( .A(n151), .B(n152), .Z(SUM[51]) );
  CANR1X1 U139 ( .A(n147), .B(net13692), .C(n148), .Z(n146) );
  CANR1X1 U146 ( .A(n153), .B(net13692), .C(n154), .Z(n152) );
  CNR2X2 U159 ( .A(B[50]), .B(A[50]), .Z(n163) );
  CANR1X1 U173 ( .A(n176), .B(net13691), .C(n177), .Z(n175) );
  CNR2X2 U186 ( .A(B[48]), .B(A[48]), .Z(n186) );
  CND2X2 U187 ( .A(B[48]), .B(A[48]), .Z(n183) );
  CEOX2 U188 ( .A(n194), .B(n195), .Z(SUM[47]) );
  CANR1X1 U197 ( .A(n196), .B(net13692), .C(n197), .Z(n195) );
  CND2X2 U204 ( .A(n220), .B(n204), .Z(n198) );
  CNR2X2 U206 ( .A(n206), .B(n214), .Z(n204) );
  CNR2X2 U210 ( .A(B[46]), .B(A[46]), .Z(n206) );
  CND2X2 U211 ( .A(B[46]), .B(A[46]), .Z(n207) );
  CEOX2 U212 ( .A(n214), .B(n215), .Z(SUM[45]) );
  CANR1X1 U221 ( .A(n216), .B(net13692), .C(n217), .Z(n215) );
  CNR2X2 U234 ( .A(B[44]), .B(A[44]), .Z(n226) );
  CND2X2 U235 ( .A(B[44]), .B(A[44]), .Z(n219) );
  CEOX2 U236 ( .A(n233), .B(n234), .Z(SUM[43]) );
  CANR1X1 U237 ( .A(n229), .B(net13691), .C(n230), .Z(n228) );
  CNR2X2 U249 ( .A(n273), .B(n241), .Z(n235) );
  CNR2X2 U274 ( .A(n262), .B(n825), .Z(n258) );
  CND2X2 U295 ( .A(n290), .B(n279), .Z(n273) );
  CNR2X2 U297 ( .A(n281), .B(n821), .Z(n279) );
  CNR2X2 U301 ( .A(B[38]), .B(A[38]), .Z(n281) );
  CNR2X2 U316 ( .A(n296), .B(n300), .Z(n290) );
  CENX2 U322 ( .A(n300), .B(net13691), .Z(SUM[35]) );
  CNR2X2 U365 ( .A(B[32]), .B(A[32]), .Z(n333) );
  CND2X2 U383 ( .A(n351), .B(n843), .Z(n345) );
  CNR2X2 U389 ( .A(B[30]), .B(A[30]), .Z(n353) );
  CANR1X1 U392 ( .A(n356), .B(n448), .C(n357), .Z(n355) );
  CNR2X2 U413 ( .A(B[28]), .B(A[28]), .Z(n373) );
  CANR1X1 U446 ( .A(n401), .B(n448), .C(n402), .Z(n400) );
  CNR2X2 U457 ( .A(B[24]), .B(A[24]), .Z(n409) );
  CEOX2 U459 ( .A(n416), .B(n417), .Z(SUM[23]) );
  CANR1X1 U460 ( .A(n412), .B(n448), .C(n413), .Z(n411) );
  CANR1X1 U467 ( .A(n422), .B(net17164), .C(n423), .Z(n417) );
  CND2X2 U474 ( .A(n426), .B(n437), .Z(n420) );
  CNR2X2 U476 ( .A(n428), .B(n435), .Z(n426) );
  CNR2X2 U480 ( .A(B[22]), .B(A[22]), .Z(n428) );
  CEOX2 U482 ( .A(n435), .B(n436), .Z(SUM[21]) );
  CANR1X1 U490 ( .A(n437), .B(net17164), .C(n442), .Z(n436) );
  CNR2X2 U495 ( .A(n443), .B(n447), .Z(n437) );
  COND1X1 U519 ( .A(net26826), .B(n459), .C(n460), .Z(n458) );
  COND1X1 U528 ( .A(n467), .B(n528), .C(n468), .Z(n466) );
  COND1X1 U544 ( .A(n480), .B(net26826), .C(n481), .Z(n479) );
  CND2X2 U565 ( .A(B[14]), .B(A[14]), .Z(n493) );
  COND1X1 U578 ( .A(n509), .B(n528), .C(n510), .Z(n508) );
  CNR2X2 U585 ( .A(B[12]), .B(A[12]), .Z(n513) );
  COND1X1 U588 ( .A(n824), .B(net26826), .C(n872), .Z(n515) );
  CNR2X2 U629 ( .A(n554), .B(n549), .Z(n544) );
  CNR2X2 U637 ( .A(B[6]), .B(A[6]), .Z(n553) );
  CND2X2 U638 ( .A(B[6]), .B(A[6]), .Z(n554) );
  CND2X2 U650 ( .A(B[4]), .B(A[4]), .Z(n562) );
  CNR2X2 U330 ( .A(n306), .B(n345), .Z(n304) );
  CANR1X1 U423 ( .A(n382), .B(net17164), .C(n383), .Z(n381) );
  CNR2X2 U643 ( .A(n562), .B(n559), .Z(n558) );
  CND2X2 U668 ( .A(net14704), .B(n576), .Z(n575) );
  CND2X2 U655 ( .A(n571), .B(n567), .Z(n566) );
  CNR2X2 U516 ( .A(B[18]), .B(A[18]), .Z(n456) );
  COR2X1 U680 ( .A(B[60]), .B(A[60]), .Z(n811) );
  CNIVXL U681 ( .A(n562), .Z(n812) );
  CIVDXL U682 ( .A(n561), .Z0(n813), .Z1(n814) );
  COAN1XL U683 ( .A(n493), .B(n475), .C(n478), .Z(n815) );
  CNR2X4 U684 ( .A(n373), .B(n380), .Z(n843) );
  CNR2X2 U685 ( .A(n513), .B(n507), .Z(n505) );
  CIVXL U686 ( .A(n392), .Z(n599) );
  COND1X2 U687 ( .A(n346), .B(n306), .C(n307), .Z(n305) );
  CAOR1X1 U688 ( .A(n557), .B(net14586), .C(n558), .Z(net14079) );
  CANR1X1 U689 ( .A(n99), .B(n79), .C(n80), .Z(n78) );
  CIVX1 U690 ( .A(n82), .Z(n80) );
  CEOX2 U691 ( .A(n68), .B(n873), .Z(SUM[59]) );
  CAOR1X1 U692 ( .A(n71), .B(net14374), .C(n72), .Z(n873) );
  COR2X1 U693 ( .A(B[12]), .B(A[12]), .Z(n816) );
  CANR1X2 U694 ( .A(n284), .B(net13691), .C(n285), .Z(n283) );
  CNR2X4 U695 ( .A(n475), .B(n492), .Z(n469) );
  CNR2IX1 U696 ( .B(n469), .A(n465), .Z(n461) );
  CIVX1 U697 ( .A(n818), .Z(n845) );
  CNR2X4 U698 ( .A(n333), .B(n341), .Z(n327) );
  CND2X2 U699 ( .A(n327), .B(n308), .Z(n306) );
  CIVXL U700 ( .A(n333), .Z(n596) );
  CND2XL U701 ( .A(n532), .B(n543), .Z(n817) );
  CANR1X2 U702 ( .A(n265), .B(net13692), .C(n266), .Z(n264) );
  CIVXL U703 ( .A(n608), .Z(net13590) );
  CANR1X1 U704 ( .A(n290), .B(net13692), .C(n295), .Z(n818) );
  CANR1X1 U705 ( .A(n290), .B(net13692), .C(n295), .Z(n289) );
  COND1X1 U706 ( .A(n814), .B(n563), .C(n812), .Z(n560) );
  CIVXL U707 ( .A(n502), .Z(n819) );
  CNR2XL U708 ( .A(n492), .B(n486), .Z(n482) );
  CND2X2 U709 ( .A(n304), .B(n382), .Z(n302) );
  CIVXL U710 ( .A(n353), .Z(n597) );
  CIVXL U711 ( .A(n75), .Z(n73) );
  CNR2X1 U712 ( .A(n77), .B(n116), .Z(n75) );
  CNR2X2 U713 ( .A(B[16]), .B(A[16]), .Z(n477) );
  COND1X2 U714 ( .A(n575), .B(n565), .C(n566), .Z(n564) );
  CANR1X1 U715 ( .A(n544), .B(n532), .C(n533), .Z(n820) );
  CANR1XL U716 ( .A(n544), .B(n532), .C(n533), .Z(n531) );
  CNR2X1 U717 ( .A(n163), .B(n174), .Z(n161) );
  CANR1X2 U718 ( .A(n185), .B(n161), .C(n162), .Z(n160) );
  COND1X1 U719 ( .A(n199), .B(n159), .C(n160), .Z(n158) );
  CENX1 U720 ( .A(n865), .B(n126), .Z(SUM[54]) );
  CANR1X1 U721 ( .A(n127), .B(net13692), .C(n128), .Z(n126) );
  CND2IX2 U722 ( .B(n321), .A(net14700), .Z(n837) );
  CANR1X1 U723 ( .A(n605), .B(n502), .C(n491), .Z(n489) );
  CENX1 U724 ( .A(n340), .B(n342), .Z(SUM[31]) );
  COND1XL U725 ( .A(net13590), .B(n546), .C(n823), .Z(n537) );
  CENXL U726 ( .A(n869), .B(n165), .Z(SUM[50]) );
  COND1X1 U727 ( .A(n365), .B(n385), .C(n366), .Z(n364) );
  CND2X2 U728 ( .A(net14006), .B(n567), .Z(n565) );
  COR2X2 U729 ( .A(A[2]), .B(B[2]), .Z(net14006) );
  CIVX2 U730 ( .A(n449), .Z(net17164) );
  CNIVXL U731 ( .A(n541), .Z(n823) );
  CIVX2 U732 ( .A(n449), .Z(n448) );
  CENX1 U733 ( .A(n525), .B(n524), .Z(SUM[11]) );
  CANR1X2 U734 ( .A(n383), .B(n304), .C(n305), .Z(n303) );
  CAN2X2 U735 ( .A(n529), .B(n450), .Z(net14198) );
  COND1X2 U736 ( .A(n302), .B(net14666), .C(n303), .Z(n2) );
  CNR2X2 U737 ( .A(n561), .B(n559), .Z(n557) );
  CNR2X2 U738 ( .A(B[4]), .B(A[4]), .Z(n561) );
  CND2X1 U739 ( .A(n811), .B(n68), .Z(n55) );
  CND2X1 U740 ( .A(n879), .B(n180), .Z(n159) );
  CNR2X2 U741 ( .A(n159), .B(n198), .Z(n157) );
  CND2X1 U742 ( .A(B[36]), .B(A[36]), .Z(n293) );
  CND2X1 U743 ( .A(B[32]), .B(A[32]), .Z(n330) );
  CND2X1 U744 ( .A(B[50]), .B(A[50]), .Z(n164) );
  CND2X2 U745 ( .A(n518), .B(n505), .Z(n499) );
  CND2XL U746 ( .A(net23257), .B(A[0]), .Z(net13593) );
  CIVDX1 U747 ( .A(A[37]), .Z0(n821), .Z1(n822) );
  COR2XL U748 ( .A(n526), .B(n524), .Z(n824) );
  CIVX1 U749 ( .A(net14373), .Z(net14374) );
  CIVDX1 U750 ( .A(A[39]), .Z0(n825), .Z1(n826) );
  CIVX1 U751 ( .A(A[33]), .Z(n321) );
  COR2XL U752 ( .A(net23257), .B(A[0]), .Z(n827) );
  CIVX1 U753 ( .A(n500), .Z(n502) );
  CIVXL U754 ( .A(n309), .Z(n828) );
  CND2XL U755 ( .A(n878), .B(n207), .Z(n13) );
  CIVX1 U756 ( .A(n492), .Z(n605) );
  CNR2XL U757 ( .A(n384), .B(n345), .Z(n343) );
  CNR2X4 U758 ( .A(n353), .B(n361), .Z(n351) );
  CIVX2 U759 ( .A(n499), .Z(n501) );
  CIVX2 U760 ( .A(n580), .Z(net14704) );
  CND2X4 U761 ( .A(n846), .B(n847), .Z(SUM[37]) );
  CND2X1 U762 ( .A(n532), .B(n543), .Z(n530) );
  COND1XL U763 ( .A(n500), .B(n829), .C(n815), .Z(n830) );
  CIVXL U764 ( .A(n469), .Z(n829) );
  CIVXL U765 ( .A(n830), .Z(n468) );
  CNR2IX2 U766 ( .B(A[9]), .A(n538), .Z(n532) );
  CNR2X2 U767 ( .A(net14198), .B(n451), .Z(n449) );
  CNR2X1 U768 ( .A(net26819), .B(net14198), .Z(net14666) );
  CNR2X2 U769 ( .A(n452), .B(n499), .Z(n450) );
  CND2X2 U770 ( .A(n469), .B(n831), .Z(n452) );
  CNR2X2 U771 ( .A(n456), .B(n465), .Z(n831) );
  CIVX2 U772 ( .A(A[17]), .Z(n465) );
  COND1X1 U773 ( .A(n530), .B(n556), .C(n820), .Z(n529) );
  CANR1X1 U774 ( .A(n564), .B(n557), .C(n558), .Z(n556) );
  COND1X1 U775 ( .A(n499), .B(n528), .C(n819), .Z(n498) );
  CNR2X2 U776 ( .A(n526), .B(n524), .Z(n518) );
  CIVX2 U777 ( .A(A[11]), .Z(n524) );
  CIVXL U778 ( .A(n456), .Z(n603) );
  COND1X1 U779 ( .A(n817), .B(net26810), .C(n531), .Z(net14687) );
  CNR2X2 U780 ( .A(n541), .B(n534), .Z(n533) );
  CIVX2 U781 ( .A(A[9]), .Z(n534) );
  CEOX1 U782 ( .A(n534), .B(n535), .Z(SUM[9]) );
  CANR1XL U783 ( .A(n564), .B(n557), .C(n558), .Z(net26810) );
  CIVX2 U784 ( .A(n573), .Z(n571) );
  CIVXL U785 ( .A(n571), .Z(net14657) );
  CND2XL U786 ( .A(net14006), .B(net14657), .Z(n35) );
  CANR1XL U787 ( .A(n574), .B(net14006), .C(n571), .Z(n569) );
  CND2X1 U788 ( .A(B[2]), .B(A[2]), .Z(n573) );
  COND1X1 U789 ( .A(n565), .B(net14643), .C(n832), .Z(net14586) );
  CND2XL U790 ( .A(n571), .B(n567), .Z(n832) );
  CENXL U791 ( .A(n567), .B(n569), .Z(SUM[3]) );
  COND1XL U792 ( .A(n500), .B(net14691), .C(n453), .Z(net26819) );
  CANR1X2 U793 ( .A(n519), .B(n505), .C(n506), .Z(n500) );
  COND1X1 U794 ( .A(n500), .B(net14691), .C(n453), .Z(n451) );
  CNR2X1 U795 ( .A(n514), .B(n507), .Z(n506) );
  CIVX2 U796 ( .A(A[13]), .Z(n507) );
  CENX1 U797 ( .A(n508), .B(n507), .Z(SUM[13]) );
  CNR2X2 U798 ( .A(n527), .B(n524), .Z(n519) );
  CND2XL U799 ( .A(n831), .B(n469), .Z(net14691) );
  CANR1X1 U800 ( .A(n470), .B(n831), .C(n455), .Z(n453) );
  CIVX2 U801 ( .A(n457), .Z(n455) );
  COND1XL U802 ( .A(n493), .B(n475), .C(n478), .Z(n470) );
  CND2XL U803 ( .A(net14704), .B(n576), .Z(net14643) );
  CENX1 U804 ( .A(net13593), .B(n576), .Z(SUM[1]) );
  CND2X1 U805 ( .A(B[0]), .B(A[0]), .Z(n580) );
  CDLY1XL U806 ( .A(B[0]), .Z(net23257) );
  CIVX2 U807 ( .A(A[5]), .Z(n559) );
  CENXL U808 ( .A(n560), .B(n559), .Z(SUM[5]) );
  CIVXL U809 ( .A(n543), .Z(n545) );
  CIVXL U810 ( .A(n544), .Z(n546) );
  CND2XL U811 ( .A(n813), .B(n562), .Z(n34) );
  CENX2 U812 ( .A(A[41]), .B(n253), .Z(SUM[41]) );
  CANR1X2 U813 ( .A(n254), .B(net13692), .C(n255), .Z(n253) );
  CIVX2 U814 ( .A(n257), .Z(n255) );
  CNIVX4 U815 ( .A(n2), .Z(net13692) );
  CIVX2 U816 ( .A(n256), .Z(n254) );
  CIVX2 U817 ( .A(A[41]), .Z(n252) );
  CNR2X2 U818 ( .A(n245), .B(n252), .Z(n243) );
  CNR2X1 U819 ( .A(n256), .B(n252), .Z(n248) );
  CNR2X1 U820 ( .A(n257), .B(n252), .Z(n249) );
  CANR1XL U821 ( .A(n258), .B(n276), .C(n261), .Z(n257) );
  CIVX2 U822 ( .A(n263), .Z(n261) );
  CANR1X2 U823 ( .A(n261), .B(n243), .C(n244), .Z(n242) );
  CIVX1 U824 ( .A(n274), .Z(n276) );
  CANR1X2 U825 ( .A(n275), .B(net13692), .C(n276), .Z(n270) );
  CNIVX4 U826 ( .A(n2), .Z(net13691) );
  CANR1X2 U827 ( .A(n332), .B(n308), .C(n309), .Z(n307) );
  CIVX1 U828 ( .A(n311), .Z(n309) );
  CIVX2 U829 ( .A(n330), .Z(n332) );
  CANR1XL U830 ( .A(n327), .B(n348), .C(n332), .Z(n326) );
  CND2XL U831 ( .A(n275), .B(n258), .Z(n256) );
  CIVX2 U832 ( .A(n273), .Z(n275) );
  CND2X2 U833 ( .A(n258), .B(n243), .Z(n241) );
  CAN2XL U834 ( .A(net13619), .B(n263), .Z(net14013) );
  COND1X2 U835 ( .A(n241), .B(n274), .C(n242), .Z(n236) );
  CNR2XL U836 ( .A(n274), .B(n825), .Z(n266) );
  CIVX2 U837 ( .A(n383), .Z(n385) );
  COND1X2 U838 ( .A(n388), .B(n421), .C(n389), .Z(n383) );
  CANR1X2 U839 ( .A(n408), .B(n390), .C(n391), .Z(n389) );
  CIVX2 U840 ( .A(n393), .Z(n391) );
  CIVX1 U841 ( .A(n410), .Z(n408) );
  CANR1X1 U842 ( .A(n405), .B(n423), .C(n408), .Z(n404) );
  CND2X1 U843 ( .A(n405), .B(n390), .Z(n388) );
  CANR1X4 U844 ( .A(n372), .B(n351), .C(n352), .Z(n346) );
  COND1X1 U845 ( .A(n345), .B(n385), .C(n346), .Z(n344) );
  CIVX2 U846 ( .A(n346), .Z(n348) );
  CIVX2 U847 ( .A(n354), .Z(n352) );
  CIVX2 U848 ( .A(n366), .Z(n372) );
  CND2XL U849 ( .A(n372), .B(n360), .Z(n359) );
  CNR2X2 U850 ( .A(n310), .B(n321), .Z(n308) );
  CIVXL U851 ( .A(net14687), .Z(net26826) );
  CIVX1 U852 ( .A(net14687), .Z(n528) );
  CNR2X2 U853 ( .A(B[10]), .B(A[10]), .Z(n526) );
  COND1X1 U854 ( .A(n96), .B(n3), .C(n97), .Z(n95) );
  CND2IX2 U855 ( .B(n822), .A(n845), .Z(n846) );
  CIVXL U856 ( .A(n373), .Z(n598) );
  CAN2XL U857 ( .A(n598), .B(n366), .Z(n867) );
  CIVX1 U858 ( .A(n236), .Z(n238) );
  CAN2X1 U859 ( .A(net17164), .B(n323), .Z(n838) );
  CIVDXL U860 ( .A(n199), .Z0(n201) );
  CND2XL U861 ( .A(n603), .B(n457), .Z(n27) );
  CND2XL U862 ( .A(n604), .B(n478), .Z(n28) );
  CNR2IXL U863 ( .B(n327), .A(n321), .Z(n317) );
  CENX1 U864 ( .A(n131), .B(n133), .Z(SUM[53]) );
  CNR2X1 U865 ( .A(n384), .B(n325), .Z(n323) );
  CEOXL U866 ( .A(n31), .B(n528), .Z(SUM[10]) );
  CNR2XL U867 ( .A(n330), .B(n321), .Z(n318) );
  CIVXL U868 ( .A(net14586), .Z(n563) );
  CENXL U869 ( .A(n549), .B(n833), .Z(SUM[7]) );
  CAOR1XL U870 ( .A(n609), .B(net14079), .C(n552), .Z(n833) );
  CAN2XL U871 ( .A(net17164), .B(n323), .Z(n834) );
  CNR2X1 U872 ( .A(n834), .B(n324), .Z(net14700) );
  CND2X2 U873 ( .A(n836), .B(n837), .Z(SUM[33]) );
  CND2IX2 U874 ( .B(A[33]), .A(n835), .Z(n836) );
  CIVX2 U875 ( .A(n322), .Z(n835) );
  CNR2X2 U876 ( .A(n838), .B(n324), .Z(n322) );
  COND1X1 U877 ( .A(n325), .B(n385), .C(n326), .Z(n324) );
  CND2X2 U878 ( .A(n174), .B(n840), .Z(n841) );
  CND2X1 U879 ( .A(n839), .B(n175), .Z(n842) );
  CND2X2 U880 ( .A(n841), .B(n842), .Z(SUM[49]) );
  CIVX2 U881 ( .A(n174), .Z(n839) );
  CIVX1 U882 ( .A(n175), .Z(n840) );
  COND1XL U883 ( .A(n136), .B(n3), .C(n137), .Z(n135) );
  CENXL U884 ( .A(n860), .B(n430), .Z(SUM[22]) );
  CANR1X1 U885 ( .A(n343), .B(n448), .C(n344), .Z(n342) );
  COND1X1 U886 ( .A(n358), .B(n385), .C(n359), .Z(n357) );
  CANR1X1 U887 ( .A(n336), .B(n448), .C(n337), .Z(n335) );
  CND2X1 U888 ( .A(n347), .B(n327), .Z(n325) );
  CEOX2 U889 ( .A(n380), .B(n381), .Z(SUM[27]) );
  CNR2X4 U890 ( .A(n392), .B(n399), .Z(n390) );
  CND2X2 U891 ( .A(n604), .B(n485), .Z(n475) );
  CIVXL U892 ( .A(n552), .Z(n844) );
  CND2XL U893 ( .A(B[16]), .B(A[16]), .Z(n478) );
  CND2X2 U894 ( .A(net13691), .B(n299), .Z(n298) );
  CNR2X2 U895 ( .A(n553), .B(n549), .Z(n543) );
  CANR1X1 U896 ( .A(n536), .B(net14079), .C(n537), .Z(n535) );
  CIVXL U897 ( .A(n554), .Z(n552) );
  CANR1XL U898 ( .A(n166), .B(net13691), .C(n167), .Z(n165) );
  CENXL U899 ( .A(n871), .B(n312), .Z(SUM[34]) );
  CIVX1 U900 ( .A(n310), .Z(n595) );
  CND2X2 U901 ( .A(n849), .B(n850), .Z(SUM[29]) );
  CANR1XL U902 ( .A(n313), .B(net17164), .C(n314), .Z(n312) );
  CANR1X1 U903 ( .A(n395), .B(n448), .C(n396), .Z(n394) );
  CND2XL U904 ( .A(B[24]), .B(A[24]), .Z(n410) );
  CIVXL U905 ( .A(net13691), .Z(net14373) );
  CENX2 U906 ( .A(n826), .B(n270), .Z(SUM[39]) );
  CANR1X1 U907 ( .A(n248), .B(net13691), .C(n249), .Z(n247) );
  CANR1XL U908 ( .A(n431), .B(net17164), .C(n432), .Z(n430) );
  CENXL U909 ( .A(n448), .B(n447), .Z(SUM[19]) );
  CENXL U910 ( .A(n35), .B(n574), .Z(SUM[2]) );
  CENXL U911 ( .A(net14079), .B(n33), .Z(SUM[6]) );
  CANR1XL U912 ( .A(n543), .B(net14079), .C(n544), .Z(n856) );
  CEOX2 U913 ( .A(n855), .B(n247), .Z(SUM[42]) );
  CANR1X1 U914 ( .A(n189), .B(net13691), .C(n190), .Z(n188) );
  CEOX2 U915 ( .A(n399), .B(n400), .Z(SUM[25]) );
  CANR1X1 U916 ( .A(n107), .B(net13692), .C(n108), .Z(n106) );
  CND2X2 U917 ( .A(n289), .B(n822), .Z(n847) );
  CANR1X1 U918 ( .A(n134), .B(net13692), .C(n135), .Z(n133) );
  CND2X1 U919 ( .A(B[10]), .B(A[10]), .Z(n527) );
  CENX2 U920 ( .A(n874), .B(n298), .Z(SUM[36]) );
  CEOX2 U921 ( .A(n13), .B(n857), .Z(SUM[46]) );
  CANR1X1 U922 ( .A(n209), .B(net13691), .C(n210), .Z(n857) );
  COND1XL U923 ( .A(n178), .B(n238), .C(n179), .Z(n177) );
  CNR2X1 U924 ( .A(n237), .B(n178), .Z(n176) );
  CIVX1 U925 ( .A(n362), .Z(n848) );
  COND1XL U926 ( .A(n116), .B(n3), .C(n117), .Z(n115) );
  CND2X1 U927 ( .A(n361), .B(n848), .Z(n849) );
  CANR1X1 U928 ( .A(n114), .B(net13691), .C(n115), .Z(n113) );
  CND2X1 U929 ( .A(net14212), .B(n362), .Z(n850) );
  CIVXL U930 ( .A(n361), .Z(net14212) );
  CENX1 U931 ( .A(n866), .B(n411), .Z(SUM[24]) );
  CND2X1 U932 ( .A(B[40]), .B(A[40]), .Z(n263) );
  CND2X1 U933 ( .A(n98), .B(n79), .Z(n77) );
  CND2XL U934 ( .A(n118), .B(n98), .Z(n96) );
  CENXL U935 ( .A(n854), .B(n83), .Z(SUM[58]) );
  CND2X2 U936 ( .A(B[28]), .B(A[28]), .Z(n366) );
  CND2X2 U937 ( .A(n235), .B(n157), .Z(n4) );
  CND2XL U938 ( .A(n200), .B(n180), .Z(n178) );
  CEOX2 U939 ( .A(n852), .B(n146), .Z(SUM[52]) );
  COND1X1 U940 ( .A(net13644), .B(n528), .C(n527), .Z(n525) );
  CEOX2 U941 ( .A(n851), .B(n228), .Z(SUM[44]) );
  CEOXL U942 ( .A(n32), .B(n856), .Z(SUM[8]) );
  CENXL U943 ( .A(n859), .B(n40), .Z(SUM[62]) );
  CAN2XL U944 ( .A(n583), .B(n82), .Z(n854) );
  CANR1XL U945 ( .A(n53), .B(n76), .C(n54), .Z(n52) );
  CNR2XL U946 ( .A(n237), .B(n233), .Z(n229) );
  CNR2X2 U947 ( .A(B[14]), .B(A[14]), .Z(n492) );
  CIVX2 U948 ( .A(n477), .Z(n604) );
  CNR2XL U949 ( .A(n237), .B(n168), .Z(n166) );
  CIVX2 U950 ( .A(n382), .Z(n384) );
  CND2XL U951 ( .A(n88), .B(n118), .Z(n86) );
  CND2XL U952 ( .A(n590), .B(n219), .Z(n851) );
  CND2XL U953 ( .A(n586), .B(n137), .Z(n852) );
  CAN2XL U954 ( .A(n584), .B(n101), .Z(n863) );
  CAN2XL U955 ( .A(n585), .B(n125), .Z(n865) );
  CNR2XL U956 ( .A(n237), .B(n218), .Z(n216) );
  CENX1 U957 ( .A(n853), .B(n61), .Z(SUM[60]) );
  CAN2XL U958 ( .A(n811), .B(n56), .Z(n853) );
  CNR2X2 U959 ( .A(n144), .B(n151), .Z(n138) );
  CAN2XL U960 ( .A(n600), .B(n410), .Z(n866) );
  CND2XL U961 ( .A(n591), .B(n246), .Z(n855) );
  CNR2XL U962 ( .A(n56), .B(n47), .Z(n46) );
  CAN2XL U963 ( .A(n597), .B(n354), .Z(n868) );
  CAN2XL U964 ( .A(n601), .B(n429), .Z(n860) );
  CENXL U965 ( .A(n47), .B(n858), .Z(SUM[61]) );
  CNR2XL U966 ( .A(n101), .B(n92), .Z(n89) );
  CNR2IXL U967 ( .B(n98), .A(n92), .Z(n88) );
  CNR2XL U968 ( .A(n293), .B(n821), .Z(n285) );
  CNR2XL U969 ( .A(n404), .B(n399), .Z(n396) );
  CNR2XL U970 ( .A(n384), .B(n380), .Z(n376) );
  COR2XL U971 ( .A(n527), .B(n524), .Z(n872) );
  CIVX1 U972 ( .A(n111), .Z(n112) );
  CAN2XL U973 ( .A(n594), .B(n293), .Z(n874) );
  CND2XL U974 ( .A(n200), .B(n193), .Z(n191) );
  CND2XL U975 ( .A(n347), .B(n340), .Z(n338) );
  CNR2XL U976 ( .A(n315), .B(n384), .Z(n313) );
  CANR1XL U977 ( .A(n41), .B(net14374), .C(n42), .Z(n40) );
  CND2XL U978 ( .A(n75), .B(n45), .Z(n43) );
  CND2XL U979 ( .A(n816), .B(n514), .Z(n30) );
  CANR1XL U980 ( .A(n180), .B(n201), .C(n185), .Z(n179) );
  CND2XL U981 ( .A(n170), .B(n200), .Z(n168) );
  CND2XL U982 ( .A(n317), .B(n347), .Z(n315) );
  CND2XL U983 ( .A(n461), .B(n501), .Z(n459) );
  CND2XL U984 ( .A(n75), .B(n53), .Z(n51) );
  CAOR1XL U985 ( .A(n49), .B(net14374), .C(n50), .Z(n858) );
  CND2XL U986 ( .A(n501), .B(n482), .Z(n480) );
  CND2XL U987 ( .A(n501), .B(n605), .Z(n488) );
  CENX1 U988 ( .A(n458), .B(n27), .Z(SUM[18]) );
  CND2XL U989 ( .A(n844), .B(n609), .Z(n33) );
  CAN2X1 U990 ( .A(n581), .B(n39), .Z(n859) );
  CENX1 U991 ( .A(n861), .B(n188), .Z(SUM[48]) );
  CAN2XL U992 ( .A(n588), .B(n183), .Z(n861) );
  CENX1 U993 ( .A(n862), .B(n335), .Z(SUM[32]) );
  CAN2XL U994 ( .A(n596), .B(n330), .Z(n862) );
  CENX1 U995 ( .A(n863), .B(n106), .Z(SUM[56]) );
  CENX1 U996 ( .A(n864), .B(n394), .Z(SUM[26]) );
  CAN2XL U997 ( .A(n599), .B(n393), .Z(n864) );
  CENX1 U998 ( .A(n867), .B(n375), .Z(SUM[28]) );
  CENX1 U999 ( .A(n868), .B(n355), .Z(SUM[30]) );
  CEOXL U1000 ( .A(n34), .B(n563), .Z(SUM[4]) );
  CAN2XL U1001 ( .A(n587), .B(n164), .Z(n869) );
  COND1XL U1002 ( .A(n218), .B(n238), .C(n219), .Z(n217) );
  CENX1 U1003 ( .A(n283), .B(n870), .Z(SUM[38]) );
  CAN2XL U1004 ( .A(n593), .B(n282), .Z(n870) );
  CNR2XL U1005 ( .A(n237), .B(n198), .Z(n196) );
  CAN2XL U1006 ( .A(n595), .B(n828), .Z(n871) );
  CNR2X1 U1007 ( .A(n4), .B(n136), .Z(n134) );
  CANR1XL U1008 ( .A(n502), .B(n461), .C(n462), .Z(n460) );
  CNR2XL U1009 ( .A(n815), .B(n465), .Z(n462) );
  CANR1XL U1010 ( .A(n119), .B(n88), .C(n89), .Z(n87) );
  CNR2XL U1011 ( .A(n55), .B(n47), .Z(n45) );
  CANR1XL U1012 ( .A(n45), .B(n76), .C(n46), .Z(n44) );
  COND1XL U1013 ( .A(n168), .B(n238), .C(n169), .Z(n167) );
  CANR1XL U1014 ( .A(n201), .B(n170), .C(n171), .Z(n169) );
  CNR2XL U1015 ( .A(n183), .B(n174), .Z(n171) );
  COND1XL U1016 ( .A(n385), .B(n315), .C(n316), .Z(n314) );
  CANR1XL U1017 ( .A(n348), .B(n317), .C(n318), .Z(n316) );
  CNR2IXL U1018 ( .B(n180), .A(n174), .Z(n170) );
  CNR2XL U1019 ( .A(n440), .B(n435), .Z(n432) );
  CNR2XL U1020 ( .A(n237), .B(n211), .Z(n209) );
  CNR2IXL U1021 ( .B(n437), .A(n435), .Z(n431) );
  CNR2XL U1022 ( .A(n238), .B(n233), .Z(n230) );
  CNR2XL U1023 ( .A(n385), .B(n380), .Z(n377) );
  CNR2XL U1024 ( .A(n237), .B(n191), .Z(n189) );
  CNR2XL U1025 ( .A(n384), .B(n338), .Z(n336) );
  CNR2XL U1026 ( .A(n273), .B(n825), .Z(n265) );
  CNR2X1 U1027 ( .A(n403), .B(n399), .Z(n395) );
  CNR2XL U1028 ( .A(n420), .B(n416), .Z(n412) );
  CNR2XL U1029 ( .A(n384), .B(n358), .Z(n356) );
  CNR2IXL U1030 ( .B(n290), .A(n821), .Z(n284) );
  CENX1 U1031 ( .A(n264), .B(net14013), .Z(SUM[40]) );
  CND2XL U1032 ( .A(n119), .B(n111), .Z(n110) );
  CND2XL U1033 ( .A(n143), .B(n131), .Z(n130) );
  CEOX1 U1034 ( .A(A[63]), .B(n37), .Z(SUM[63]) );
  COND1XL U1035 ( .A(n38), .B(n40), .C(n39), .Z(n37) );
  COND1XL U1036 ( .A(n211), .B(n238), .C(n212), .Z(n210) );
  CENX1 U1037 ( .A(n875), .B(n445), .Z(SUM[20]) );
  CAN2XL U1038 ( .A(n602), .B(n440), .Z(n875) );
  CNR2X1 U1039 ( .A(B[52]), .B(A[52]), .Z(n144) );
  CND2XL U1040 ( .A(n76), .B(n68), .Z(n65) );
  COND1XL U1041 ( .A(n191), .B(n238), .C(n192), .Z(n190) );
  COND1XL U1042 ( .A(n338), .B(n385), .C(n339), .Z(n337) );
  CNR2X1 U1043 ( .A(B[62]), .B(A[62]), .Z(n38) );
  CND2X1 U1044 ( .A(B[60]), .B(A[60]), .Z(n56) );
  CND2X1 U1045 ( .A(B[56]), .B(A[56]), .Z(n101) );
  CND2X1 U1046 ( .A(B[52]), .B(A[52]), .Z(n137) );
  CND2X1 U1047 ( .A(B[22]), .B(A[22]), .Z(n429) );
  CND2X1 U1048 ( .A(B[58]), .B(A[58]), .Z(n82) );
  CND2X1 U1049 ( .A(B[54]), .B(A[54]), .Z(n125) );
  CND2X1 U1050 ( .A(B[30]), .B(A[30]), .Z(n354) );
  CND2X1 U1051 ( .A(B[18]), .B(A[18]), .Z(n457) );
  CND2X1 U1052 ( .A(B[62]), .B(A[62]), .Z(n39) );
  CND2XL U1053 ( .A(n220), .B(n213), .Z(n211) );
  CAN2XL U1054 ( .A(n827), .B(net13593), .Z(SUM[0]) );
  CND2XL U1055 ( .A(n75), .B(n68), .Z(n64) );
  CND2XL U1056 ( .A(n118), .B(n111), .Z(n109) );
  CND2XL U1057 ( .A(n138), .B(n131), .Z(n129) );
  CANR1X1 U1058 ( .A(n376), .B(n448), .C(n377), .Z(n375) );
  CANR1X1 U1059 ( .A(n363), .B(net17164), .C(n364), .Z(n362) );
  CNR2XL U1060 ( .A(n4), .B(n43), .Z(n41) );
  CNR2XL U1061 ( .A(n4), .B(n51), .Z(n49) );
  CNR2XL U1062 ( .A(n4), .B(n73), .Z(n71) );
  CNR2XL U1063 ( .A(n4), .B(n64), .Z(n62) );
  CNR2XL U1064 ( .A(n4), .B(n86), .Z(n84) );
  CNR2XL U1065 ( .A(n4), .B(n109), .Z(n107) );
  CNR2X1 U1066 ( .A(n4), .B(n116), .Z(n114) );
  CNR2XL U1067 ( .A(n4), .B(n129), .Z(n127) );
  CNR2XL U1068 ( .A(n4), .B(n96), .Z(n94) );
  CNR2X1 U1069 ( .A(n4), .B(n151), .Z(n147) );
  CIVXL U1070 ( .A(n4), .Z(n153) );
  CANR1XL U1071 ( .A(n62), .B(net14374), .C(n63), .Z(n61) );
  CANR1XL U1072 ( .A(n84), .B(net14374), .C(n85), .Z(n83) );
  COND1XL U1073 ( .A(n129), .B(n3), .C(n130), .Z(n128) );
  CANR1X1 U1074 ( .A(n235), .B(net13691), .C(n236), .Z(n234) );
  CNR2X1 U1075 ( .A(B[36]), .B(A[36]), .Z(n296) );
  CND2X1 U1076 ( .A(B[38]), .B(A[38]), .Z(n282) );
  CNR2X1 U1077 ( .A(B[40]), .B(A[40]), .Z(n262) );
  CND2X1 U1078 ( .A(B[42]), .B(A[42]), .Z(n246) );
  CNR2X1 U1079 ( .A(B[42]), .B(A[42]), .Z(n245) );
  CND2X1 U1080 ( .A(n225), .B(n213), .Z(n212) );
  CND2X1 U1081 ( .A(n201), .B(n193), .Z(n192) );
  CIVXL U1082 ( .A(n3), .Z(n154) );
  CIVXL U1083 ( .A(net14643), .Z(n574) );
  CNR2X2 U1084 ( .A(B[26]), .B(A[26]), .Z(n392) );
  CND2X2 U1085 ( .A(n405), .B(n390), .Z(n877) );
  CND2XL U1086 ( .A(n607), .B(n527), .Z(n31) );
  CANR1XL U1087 ( .A(n816), .B(n519), .C(n512), .Z(n510) );
  CND2XL U1088 ( .A(n518), .B(n816), .Z(n509) );
  CIVXL U1089 ( .A(n607), .Z(net13644) );
  CIVXL U1090 ( .A(n526), .Z(n607) );
  CNR2X4 U1091 ( .A(n226), .B(n233), .Z(n220) );
  CNR2X1 U1092 ( .A(n545), .B(net13590), .Z(n536) );
  CANR1XL U1093 ( .A(n482), .B(n502), .C(n483), .Z(n481) );
  COR2XL U1094 ( .A(A[46]), .B(B[46]), .Z(n878) );
  CNR2X1 U1095 ( .A(n163), .B(n174), .Z(n879) );
  CND2X1 U1096 ( .A(n422), .B(n405), .Z(n403) );
  COR2XL U1097 ( .A(B[40]), .B(A[40]), .Z(net13619) );
  CIVX1 U1098 ( .A(n421), .Z(n423) );
  CNR2XL U1099 ( .A(n421), .B(n416), .Z(n413) );
  CIVXL U1100 ( .A(n186), .Z(n588) );
  CENX1 U1101 ( .A(n498), .B(n29), .Z(SUM[14]) );
  CENX1 U1102 ( .A(n487), .B(n486), .Z(SUM[15]) );
  CND2X1 U1103 ( .A(B[26]), .B(A[26]), .Z(n393) );
  CND2X1 U1104 ( .A(n843), .B(n360), .Z(n358) );
  CND2X1 U1105 ( .A(n348), .B(n340), .Z(n339) );
  CND2X1 U1106 ( .A(B[34]), .B(A[34]), .Z(n311) );
  CIVXL U1107 ( .A(n245), .Z(n591) );
  CIVXL U1108 ( .A(n514), .Z(n512) );
  CND2X1 U1109 ( .A(B[12]), .B(A[12]), .Z(n514) );
  CIVXL U1110 ( .A(n553), .Z(n609) );
  CNR2X2 U1111 ( .A(B[34]), .B(A[34]), .Z(n310) );
  CIVXL U1112 ( .A(n538), .Z(n608) );
  CNR2X2 U1113 ( .A(B[8]), .B(A[8]), .Z(n538) );
  CND2X1 U1114 ( .A(B[20]), .B(A[20]), .Z(n440) );
  CNR2X1 U1115 ( .A(B[20]), .B(A[20]), .Z(n443) );
  CND2XL U1116 ( .A(n823), .B(n608), .Z(n32) );
  COND1X1 U1117 ( .A(n488), .B(n528), .C(n489), .Z(n487) );
  CNR2X4 U1118 ( .A(n409), .B(n416), .Z(n405) );
  CNR2X4 U1119 ( .A(n420), .B(n877), .Z(n382) );
  CNR2X4 U1120 ( .A(n186), .B(n194), .Z(n180) );
  COND1XL U1121 ( .A(n198), .B(n238), .C(n199), .Z(n197) );
  CND2XL U1122 ( .A(n501), .B(n469), .Z(n467) );
  CENX1 U1123 ( .A(n466), .B(n465), .Z(SUM[17]) );
  CND2X2 U1124 ( .A(B[8]), .B(A[8]), .Z(n541) );
  CND2XL U1125 ( .A(n605), .B(n493), .Z(n29) );
  CNR2XL U1126 ( .A(n493), .B(n486), .Z(n483) );
  CNR2X1 U1127 ( .A(n384), .B(n365), .Z(n363) );
  CANR1X2 U1128 ( .A(n442), .B(n426), .C(n427), .Z(n421) );
  CANR1X2 U1129 ( .A(n236), .B(n157), .C(n158), .Z(n3) );
  CANR1X2 U1130 ( .A(n225), .B(n204), .C(n205), .Z(n199) );
  CND2X1 U1131 ( .A(n448), .B(n446), .Z(n445) );
  COND1XL U1132 ( .A(n43), .B(n3), .C(n44), .Z(n42) );
  COND1XL U1133 ( .A(n64), .B(n3), .C(n65), .Z(n63) );
  COND1XL U1134 ( .A(n51), .B(n3), .C(n52), .Z(n50) );
  COND1XL U1135 ( .A(n86), .B(n3), .C(n87), .Z(n85) );
  COND1XL U1136 ( .A(n73), .B(n3), .C(n74), .Z(n72) );
  CNR2XL U1137 ( .A(n3), .B(n151), .Z(n148) );
  COND1XL U1138 ( .A(n109), .B(n3), .C(n110), .Z(n108) );
  CENX1 U1139 ( .A(n479), .B(n28), .Z(SUM[16]) );
  CANR1X2 U1140 ( .A(n295), .B(n279), .C(n280), .Z(n274) );
  CENX1 U1141 ( .A(n515), .B(n30), .Z(SUM[12]) );
  CIVX2 U1142 ( .A(A[57]), .Z(n92) );
  CIVX2 U1143 ( .A(n76), .Z(n74) );
  CIVX2 U1144 ( .A(n443), .Z(n602) );
  CIVX2 U1145 ( .A(n428), .Z(n601) );
  CIVX2 U1146 ( .A(n409), .Z(n600) );
  CIVX2 U1147 ( .A(n296), .Z(n594) );
  CIVX2 U1148 ( .A(n281), .Z(n593) );
  CIVX2 U1149 ( .A(n226), .Z(n590) );
  CIVX2 U1150 ( .A(n163), .Z(n587) );
  CIVX2 U1151 ( .A(n144), .Z(n586) );
  CIVX2 U1152 ( .A(n124), .Z(n585) );
  CIVX2 U1153 ( .A(n104), .Z(n584) );
  CIVX2 U1154 ( .A(n81), .Z(n583) );
  CIVX2 U1155 ( .A(n38), .Z(n581) );
  CIVX2 U1156 ( .A(A[7]), .Z(n549) );
  CIVX2 U1157 ( .A(n56), .Z(n54) );
  CIVX2 U1158 ( .A(n55), .Z(n53) );
  CIVX2 U1159 ( .A(n493), .Z(n491) );
  CIVX2 U1160 ( .A(n485), .Z(n486) );
  CIVX2 U1161 ( .A(A[61]), .Z(n47) );
  CIVX2 U1162 ( .A(n446), .Z(n447) );
  CIVX2 U1163 ( .A(n440), .Z(n442) );
  CIVX2 U1164 ( .A(A[21]), .Z(n435) );
  CIVX2 U1165 ( .A(n429), .Z(n427) );
  CIVX2 U1166 ( .A(n420), .Z(n422) );
  CIVX2 U1167 ( .A(A[23]), .Z(n416) );
  CIVX2 U1168 ( .A(n404), .Z(n402) );
  CIVX2 U1169 ( .A(n403), .Z(n401) );
  CIVX2 U1170 ( .A(A[25]), .Z(n399) );
  CIVX2 U1171 ( .A(A[27]), .Z(n380) );
  CIVX2 U1172 ( .A(n843), .Z(n365) );
  CIVX2 U1173 ( .A(n360), .Z(n361) );
  CIVX2 U1174 ( .A(n345), .Z(n347) );
  CIVX2 U1175 ( .A(n340), .Z(n341) );
  CIVX2 U1176 ( .A(n299), .Z(n300) );
  CIVX2 U1177 ( .A(n293), .Z(n295) );
  CIVX2 U1178 ( .A(n282), .Z(n280) );
  CIVX2 U1179 ( .A(n246), .Z(n244) );
  CIVX2 U1180 ( .A(n235), .Z(n237) );
  CIVX2 U1181 ( .A(A[43]), .Z(n233) );
  CIVX2 U1182 ( .A(n219), .Z(n225) );
  CIVX2 U1183 ( .A(n220), .Z(n218) );
  CIVX2 U1184 ( .A(n213), .Z(n214) );
  CIVX2 U1185 ( .A(n207), .Z(n205) );
  CIVX2 U1186 ( .A(n198), .Z(n200) );
  CIVX2 U1187 ( .A(n193), .Z(n194) );
  CIVX2 U1188 ( .A(n183), .Z(n185) );
  CIVX2 U1189 ( .A(A[49]), .Z(n174) );
  CIVX2 U1190 ( .A(n164), .Z(n162) );
  CIVX2 U1191 ( .A(A[51]), .Z(n151) );
  CIVX2 U1192 ( .A(n137), .Z(n143) );
  CIVX2 U1193 ( .A(n138), .Z(n136) );
  CIVX2 U1194 ( .A(n131), .Z(n132) );
  CIVX2 U1195 ( .A(n125), .Z(n123) );
  CIVX2 U1196 ( .A(n117), .Z(n119) );
  CIVX2 U1197 ( .A(n116), .Z(n118) );
  CIVX2 U1198 ( .A(n101), .Z(n99) );
endmodule


module sqrt64_DW01_add_10 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n8, n9, n12, n13, n16, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47,
         n48, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n67, n74, n76, n78, n79, n84, n85, n86, n87, n88, n105,
         n106, n110, n116, n120, n121, n122, n123, n124, n125, n126, n144,
         n145, n146, n147, n148, n149, n150, n152, n153, n154, n155, n156,
         n157, n158, n164, n166, n167, n168, n169, n170, n171, n172, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n188, n189, n190,
         n191, n192, n193, n196, n197, n198, n200, n201, n204, n206, n208,
         n209, n210, n211, n212, n213, n216, n217, n218, n219, n220, n221,
         n222, n225, n226, n227, n228, n229, n230, n231, n234, n235, n238,
         n239, n240, n241, n244, n245, n246, n247, n248, n249, n250, n251,
         n254, n255, n256, n257, n259, n262, n263, n264, n266, n267, n268,
         n269, n279, n280, n281, n282, n283, n288, n289, n290, n297, n298,
         n299, n300, n301, n303, n304, n305, n306, n309, n310, n314, n315,
         n316, n317, n318, n319, n321, n322, n323, n324, n325, n326, n327,
         n337, n338, n339, n340, n341, n347, n348, n349, n351, n352, n359,
         n360, n366, n372, n377, n378, n379, n380, n381, n382, n388, n389,
         n390, n391, n392, n393, n400, n401, n402, n403, n404, n405, n406,
         n411, n412, n415, n418, n419, n421, n423, n424, n425, n426, n427,
         n428, n430, n433, n434, n435, n436, n437, n443, n445, n446, n448,
         n450, n451, n452, n453, n454, n455, n456, n458, n460, n461, n462,
         n463, n467, n468, n469, n470, n471, n472, n473, n474, n478, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n505, n507, n508, n509, n510, n511, n512, n513, n514, n516, n519,
         n520, n521, n522, n523, n526, n527, n529, n530, n531, n532, n533,
         n534, n535, n536, n538, n541, n542, n543, n544, n545, n551, n552,
         n553, n554, n556, n558, n559, n560, n561, n562, n563, n564, n566,
         n568, n569, n570, n571, n575, n576, n577, n578, n579, n580, n581,
         n582, n586, n588, n589, n590, n591, n593, n596, n597, n598, n599,
         n601, n603, n604, n606, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n623, n625, n626, n627,
         n628, n630, n636, n640, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n653, n654, n655, n659, n660, n661, n665, n668,
         n669, n671, n675, n677, n678, n679, n680, n681, n682, n683, n684,
         n687, n689, n692, n693, n695, \B[0] , net13575, net13631, net14046,
         net14085, net14087, net14090, net14094, net14098, net14130, net14129,
         net14384, net14588, net14587, net14622, net14626, net14628, net14690,
         net14721, net14742, n350, n664, n357, n132, n129, n118, n10, net14584,
         net14710, net14569, n183, n165, n161, n160, n159, n141, n139, n138,
         n137, n136, n135, n134, n133, n128, n127, net14743, n657, net19919,
         net19921, net26798, net26801, net26821, net26823, net14110, net14104,
         n92, n89, n637, n97, n96, n95, n94, n93, n108, n103, n662, n345, n336,
         n334, n333, n328, n313, n395, n370, n307, n658, n294, n292, n284,
         n275, net14379, n287, n278, n277, n207, n205, n2, n199, n119, n117,
         n115, n114, n113, net14638, net14585, net14362, net14204, n413, n386,
         n375, n373, n371, n369, n368, n367, n308, n276, n274, n272, n271,
         n112, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n962, n963, n964, n965, n966;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  CNR2X2 U107 ( .A(B[55]), .B(A[55]), .Z(n144) );
  CND2X2 U129 ( .A(n164), .B(n182), .Z(n158) );
  CNR2X2 U135 ( .A(B[53]), .B(A[53]), .Z(n166) );
  CANR1X1 U150 ( .A(n178), .B(n269), .C(n179), .Z(n177) );
  COND1X1 U152 ( .A(n180), .B(n201), .C(n181), .Z(n179) );
  CNR2X2 U159 ( .A(n193), .B(n188), .Z(n182) );
  CANR1X1 U166 ( .A(n191), .B(net14129), .C(n192), .Z(n190) );
  CND2X2 U183 ( .A(n222), .B(n206), .Z(n204) );
  CNR2X2 U185 ( .A(n208), .B(n213), .Z(n206) );
  CNR2X2 U189 ( .A(B[49]), .B(A[49]), .Z(n208) );
  CANR1X1 U192 ( .A(n211), .B(net14129), .C(n212), .Z(n210) );
  CANR1X1 U202 ( .A(n218), .B(n269), .C(n219), .Z(n217) );
  CANR1X1 U206 ( .A(n222), .B(n241), .C(n225), .Z(n221) );
  CNR2X2 U209 ( .A(n231), .B(n226), .Z(n222) );
  CNR2X2 U213 ( .A(B[47]), .B(A[47]), .Z(n226) );
  CANR1X1 U216 ( .A(n229), .B(net26801), .C(n230), .Z(n228) );
  CANR1X1 U226 ( .A(n240), .B(net26801), .C(n241), .Z(n235) );
  CNR2X2 U235 ( .A(n251), .B(n246), .Z(n244) );
  CNR2X2 U239 ( .A(B[45]), .B(A[45]), .Z(n246) );
  CANR1X1 U252 ( .A(n256), .B(n269), .C(n257), .Z(n255) );
  CNR2X2 U261 ( .A(B[43]), .B(A[43]), .Z(n262) );
  CANR1X1 U264 ( .A(n655), .B(n269), .C(n266), .Z(n264) );
  CNR2X2 U342 ( .A(B[36]), .B(A[36]), .Z(n322) );
  CND2X2 U343 ( .A(A[36]), .B(B[36]), .Z(n323) );
  COND1X1 U345 ( .A(n325), .B(net26798), .C(n326), .Z(n324) );
  CNR2X2 U352 ( .A(n915), .B(n349), .Z(n327) );
  CANR1X1 U484 ( .A(n434), .B(n451), .C(n435), .Z(n433) );
  COND1X1 U511 ( .A(n455), .B(n472), .C(n456), .Z(n454) );
  CND2X2 U512 ( .A(n675), .B(n902), .Z(n455) );
  CANR1X1 U513 ( .A(n467), .B(n902), .C(n458), .Z(n456) );
  CNR2X2 U571 ( .A(B[18]), .B(A[18]), .Z(n497) );
  CND2X2 U607 ( .A(n683), .B(n682), .Z(n526) );
  COND1X1 U655 ( .A(n580), .B(n563), .C(n564), .Z(n562) );
  CNR2X2 U308 ( .A(B[39]), .B(A[39]), .Z(n297) );
  CND2X2 U71 ( .A(n138), .B(n118), .Z(n116) );
  CNR2X2 U103 ( .A(n153), .B(n144), .Z(n138) );
  CANR1X1 U94 ( .A(n134), .B(n269), .C(n135), .Z(n133) );
  CNR2X2 U328 ( .A(net14690), .B(n322), .Z(n313) );
  CNR2X2 U69 ( .A(n158), .B(n116), .Z(n114) );
  CANR1X1 U176 ( .A(n198), .B(net14129), .C(n199), .Z(n197) );
  CND2X2 U326 ( .A(n313), .B(n327), .Z(n307) );
  COND1X1 U279 ( .A(n287), .B(n277), .C(n278), .Z(n276) );
  CANR1X1 U277 ( .A(n292), .B(n275), .C(n276), .Z(n274) );
  COND1X1 U275 ( .A(net14362), .B(n308), .C(n274), .Z(n272) );
  COR2X1 U763 ( .A(B[21]), .B(A[21]), .Z(n894) );
  CND2X1 U764 ( .A(n275), .B(net14742), .Z(net14362) );
  COR2XL U765 ( .A(n436), .B(n418), .Z(n895) );
  CIVX2 U766 ( .A(n552), .Z(n684) );
  CANR1X2 U767 ( .A(n108), .B(net14046), .C(n103), .Z(n97) );
  CIVXL U768 ( .A(net13631), .Z(n896) );
  COR2X1 U769 ( .A(A[11]), .B(B[11]), .Z(n897) );
  COR2XL U770 ( .A(A[11]), .B(B[11]), .Z(n966) );
  CIVXL U771 ( .A(n226), .Z(n650) );
  CNR2X2 U772 ( .A(B[35]), .B(A[35]), .Z(n900) );
  CNR2XL U773 ( .A(A[35]), .B(B[35]), .Z(n337) );
  COR2X1 U774 ( .A(B[34]), .B(A[34]), .Z(net14085) );
  CNIVXL U775 ( .A(n664), .Z(n898) );
  CANR1XL U776 ( .A(n390), .B(n451), .C(n391), .Z(n389) );
  CND2XL U777 ( .A(n677), .B(n487), .Z(n46) );
  CENXL U778 ( .A(n488), .B(n46), .Z(SUM[20]) );
  CANR1XL U779 ( .A(n901), .B(n898), .C(n896), .Z(n899) );
  COND1X2 U780 ( .A(n1), .B(n620), .C(n621), .Z(n619) );
  CNR2X2 U781 ( .A(n471), .B(n455), .Z(n453) );
  CND2X1 U782 ( .A(B[19]), .B(A[19]), .Z(n490) );
  CND2X1 U783 ( .A(n897), .B(n687), .Z(n563) );
  CIVXL U784 ( .A(n437), .Z(n435) );
  CENXL U785 ( .A(n339), .B(n31), .Z(SUM[35]) );
  CND2X2 U786 ( .A(B[35]), .B(A[35]), .Z(n338) );
  CANR1X2 U787 ( .A(n894), .B(n485), .C(n478), .Z(n472) );
  CNR2X2 U788 ( .A(B[15]), .B(A[15]), .Z(n530) );
  CIVXL U789 ( .A(n545), .Z(n543) );
  COR2X2 U790 ( .A(B[12]), .B(A[12]), .Z(n951) );
  CND2X1 U791 ( .A(B[11]), .B(A[11]), .Z(n568) );
  CNR2XL U792 ( .A(B[8]), .B(A[8]), .Z(n590) );
  COND1X1 U793 ( .A(n196), .B(n188), .C(n189), .Z(n183) );
  COND1X1 U794 ( .A(n176), .B(n166), .C(n167), .Z(n165) );
  CND2X1 U795 ( .A(net14094), .B(net14046), .Z(n96) );
  CIVXL U796 ( .A(n183), .Z(n181) );
  CNR2X1 U797 ( .A(B[48]), .B(A[48]), .Z(n213) );
  CND2X1 U798 ( .A(B[63]), .B(A[63]), .Z(n67) );
  CAN2X1 U799 ( .A(B[32]), .B(A[32]), .Z(n901) );
  COR2X1 U800 ( .A(A[23]), .B(B[23]), .Z(n902) );
  CAOR1XL U801 ( .A(n956), .B(n79), .C(n74), .Z(n903) );
  COAN1XL U802 ( .A(n92), .B(n84), .C(n85), .Z(n904) );
  COR2XL U803 ( .A(A[1]), .B(B[1]), .Z(n905) );
  CIVX1 U804 ( .A(n158), .Z(n160) );
  CND2X2 U805 ( .A(n256), .B(n244), .Z(n238) );
  CND2X2 U806 ( .A(net14204), .B(n907), .Z(n908) );
  CND2X2 U807 ( .A(n908), .B(n113), .Z(n2) );
  CIVX2 U808 ( .A(n112), .Z(n907) );
  CIVX1 U809 ( .A(net14585), .Z(net14204) );
  CND2XL U810 ( .A(net14204), .B(n907), .Z(net14130) );
  CANR1X1 U811 ( .A(net14638), .B(n367), .C(n272), .Z(net14585) );
  CNR2X1 U812 ( .A(net14362), .B(n307), .Z(net14638) );
  CND2X2 U813 ( .A(n198), .B(n114), .Z(n112) );
  COND1X2 U814 ( .A(n368), .B(n452), .C(n369), .Z(n367) );
  CIVXL U815 ( .A(n367), .Z(net26798) );
  CIVX2 U816 ( .A(n367), .Z(n366) );
  CANR1X1 U817 ( .A(n271), .B(n367), .C(n272), .Z(net14584) );
  CANR1X2 U818 ( .A(n413), .B(n370), .C(n371), .Z(n369) );
  COND1X1 U819 ( .A(n372), .B(n393), .C(n373), .Z(n371) );
  CANR1X1 U820 ( .A(n386), .B(net14090), .C(n375), .Z(n373) );
  CIVX2 U821 ( .A(n377), .Z(n375) );
  CIVXL U822 ( .A(n388), .Z(n386) );
  CANR1XL U823 ( .A(net14098), .B(n395), .C(n386), .Z(n382) );
  COND1X1 U824 ( .A(n418), .B(n437), .C(n419), .Z(n413) );
  CND2X1 U825 ( .A(n906), .B(n370), .Z(n368) );
  CNR2X1 U826 ( .A(n436), .B(n418), .Z(n906) );
  CANR1X1 U827 ( .A(n313), .B(n328), .C(n314), .Z(n308) );
  CNR2X1 U828 ( .A(net14362), .B(n307), .Z(n271) );
  CANR1X1 U829 ( .A(net14094), .B(n2), .C(n108), .Z(n106) );
  CANR1X2 U830 ( .A(n94), .B(n2), .C(n95), .Z(n93) );
  CANR1X1 U831 ( .A(n199), .B(n114), .C(n115), .Z(n113) );
  COND1X2 U832 ( .A(n204), .B(n239), .C(n205), .Z(n199) );
  CIVX2 U833 ( .A(n199), .Z(n201) );
  CANR1XL U834 ( .A(n199), .B(n114), .C(n115), .Z(net14626) );
  CANR1X2 U835 ( .A(n225), .B(n206), .C(n207), .Z(n205) );
  COND1X2 U836 ( .A(n216), .B(n208), .C(n209), .Z(n207) );
  COND1X1 U837 ( .A(n116), .B(net14384), .C(n117), .Z(n115) );
  CANR1X1 U838 ( .A(n139), .B(n118), .C(n119), .Z(n117) );
  COND1XL U839 ( .A(n132), .B(n120), .C(n121), .Z(n119) );
  CNR2X2 U840 ( .A(B[41]), .B(A[41]), .Z(n277) );
  CNR2X1 U841 ( .A(n284), .B(n277), .Z(n275) );
  COR2XL U842 ( .A(A[41]), .B(B[41]), .Z(net14379) );
  CND2X1 U843 ( .A(B[41]), .B(A[41]), .Z(n278) );
  CND2X1 U844 ( .A(B[40]), .B(A[40]), .Z(n287) );
  CND2XL U845 ( .A(n287), .B(n657), .Z(n26) );
  COND1XL U846 ( .A(net19919), .B(n294), .C(n287), .Z(n283) );
  CND2XL U847 ( .A(net14379), .B(n278), .Z(n25) );
  CNR2X1 U848 ( .A(B[40]), .B(A[40]), .Z(n284) );
  COND1X1 U849 ( .A(n305), .B(n297), .C(n298), .Z(n292) );
  CANR1XL U850 ( .A(net14743), .B(n310), .C(n292), .Z(n290) );
  CIVXL U851 ( .A(n292), .Z(n294) );
  CIVXL U852 ( .A(n305), .Z(n303) );
  CND2XL U853 ( .A(n659), .B(n305), .Z(n28) );
  CNR2X1 U854 ( .A(n304), .B(n297), .Z(net14742) );
  CNR2XL U855 ( .A(n304), .B(n297), .Z(net14743) );
  CIVXL U856 ( .A(n297), .Z(n658) );
  CND2XL U857 ( .A(n658), .B(n298), .Z(n27) );
  CIVXL U858 ( .A(n284), .Z(n657) );
  COND1XL U859 ( .A(n307), .B(n366), .C(net26821), .Z(n306) );
  CIVX2 U860 ( .A(n307), .Z(n309) );
  CIVX1 U861 ( .A(n452), .Z(n451) );
  CNR2X2 U862 ( .A(n392), .B(n372), .Z(n370) );
  COND1XL U863 ( .A(n392), .B(n415), .C(n393), .Z(n391) );
  CIVX2 U864 ( .A(n393), .Z(n395) );
  CANR1X1 U865 ( .A(n313), .B(n328), .C(n314), .Z(net14587) );
  COND1X2 U866 ( .A(n350), .B(n333), .C(n334), .Z(n328) );
  CIVXL U867 ( .A(n328), .Z(n326) );
  CANR1X2 U868 ( .A(n345), .B(n662), .C(n336), .Z(n334) );
  CIVX2 U869 ( .A(n338), .Z(n336) );
  CIVX2 U870 ( .A(n900), .Z(n662) );
  CND2XL U871 ( .A(n662), .B(n338), .Z(n31) );
  CIVX2 U872 ( .A(n347), .Z(n345) );
  CANR1XL U873 ( .A(net14085), .B(n352), .C(n345), .Z(n341) );
  CND2IX1 U874 ( .B(n900), .A(net14085), .Z(n333) );
  CENX2 U875 ( .A(net14110), .B(n93), .Z(SUM[60]) );
  CIVX2 U876 ( .A(n97), .Z(n95) );
  CIVX2 U877 ( .A(n96), .Z(n94) );
  COND1XL U878 ( .A(n97), .B(net14104), .C(n904), .Z(n79) );
  COND1XL U879 ( .A(n89), .B(n97), .C(n92), .Z(n88) );
  CIVX2 U880 ( .A(n105), .Z(n103) );
  CIVX2 U881 ( .A(n110), .Z(n108) );
  CNR2XL U882 ( .A(net14104), .B(n96), .Z(n78) );
  CNR2XL U883 ( .A(n96), .B(n89), .Z(n87) );
  CAN2X1 U884 ( .A(n637), .B(n92), .Z(net14110) );
  CIVX2 U885 ( .A(n89), .Z(n637) );
  CND2X1 U886 ( .A(B[60]), .B(A[60]), .Z(n92) );
  CNR2X1 U887 ( .A(B[60]), .B(A[60]), .Z(n89) );
  COR2XL U888 ( .A(n89), .B(n84), .Z(net14104) );
  CIVXL U889 ( .A(n267), .Z(n655) );
  CND2XL U890 ( .A(B[55]), .B(A[55]), .Z(n145) );
  CIVXL U891 ( .A(n651), .Z(n909) );
  CIVXL U892 ( .A(n231), .Z(n651) );
  CNR2X1 U893 ( .A(B[17]), .B(A[17]), .Z(n508) );
  CND2X1 U894 ( .A(A[17]), .B(B[17]), .Z(n509) );
  COND1X1 U895 ( .A(n418), .B(n437), .C(n419), .Z(net26823) );
  CIVXL U896 ( .A(net19921), .Z(net26821) );
  CIVXL U897 ( .A(n647), .Z(n910) );
  CIVX1 U898 ( .A(net14584), .Z(net26801) );
  CIVX1 U899 ( .A(net14584), .Z(n269) );
  CNR2X1 U900 ( .A(B[10]), .B(A[10]), .Z(n576) );
  CIVX1 U901 ( .A(n577), .Z(n575) );
  CND2X1 U902 ( .A(B[57]), .B(A[57]), .Z(n121) );
  CND2X1 U903 ( .A(n351), .B(net14085), .Z(n340) );
  CNR2X4 U904 ( .A(n544), .B(n526), .Z(n520) );
  CIVX1 U905 ( .A(net26823), .Z(n415) );
  CANR1XL U906 ( .A(n412), .B(n451), .C(net26823), .Z(n411) );
  CANR1XL U907 ( .A(n249), .B(net26801), .C(n250), .Z(n248) );
  COND1X1 U908 ( .A(n323), .B(n315), .C(n316), .Z(n314) );
  CENX1 U909 ( .A(n911), .B(n177), .Z(SUM[52]) );
  CAN2XL U910 ( .A(n645), .B(n176), .Z(n911) );
  CENXL U911 ( .A(n912), .B(net26801), .Z(SUM[42]) );
  CND2XL U912 ( .A(n655), .B(n268), .Z(n912) );
  CENXL U913 ( .A(n913), .B(n248), .Z(SUM[45]) );
  CAN2XL U914 ( .A(n920), .B(n247), .Z(n913) );
  CANR1XL U915 ( .A(n78), .B(n964), .C(n79), .Z(n940) );
  CIVXL U916 ( .A(net14587), .Z(net19921) );
  CIVXL U917 ( .A(net14587), .Z(n310) );
  CIVXL U918 ( .A(n657), .Z(net19919) );
  CENX1 U919 ( .A(n914), .B(n255), .Z(SUM[44]) );
  CAN2XL U920 ( .A(n653), .B(n254), .Z(n914) );
  COND1X2 U921 ( .A(n234), .B(n226), .C(n227), .Z(n225) );
  CNR2IXL U922 ( .B(net14743), .A(net19919), .Z(n282) );
  CEOX1 U923 ( .A(n133), .B(n10), .Z(SUM[56]) );
  COND1X1 U924 ( .A(n136), .B(n201), .C(n137), .Z(n135) );
  CANR1X1 U925 ( .A(n138), .B(n161), .C(net14569), .Z(n137) );
  CIVXL U926 ( .A(n141), .Z(net14569) );
  CIVXL U927 ( .A(n139), .Z(n141) );
  COND1XL U928 ( .A(n129), .B(n141), .C(n132), .Z(n128) );
  CIVX1 U929 ( .A(n159), .Z(n161) );
  CANR1XL U930 ( .A(n161), .B(n127), .C(n128), .Z(n126) );
  CANR1XL U931 ( .A(n643), .B(n161), .C(n152), .Z(n150) );
  CANR1X1 U932 ( .A(n183), .B(net14710), .C(n165), .Z(n159) );
  CNR2X1 U933 ( .A(n200), .B(n136), .Z(n134) );
  CIVX2 U934 ( .A(n198), .Z(n200) );
  CND2X1 U935 ( .A(n160), .B(n138), .Z(n136) );
  CND2XL U936 ( .A(n127), .B(n160), .Z(n125) );
  CND2XL U937 ( .A(n160), .B(n643), .Z(n149) );
  CNR2IX1 U938 ( .B(n138), .A(n129), .Z(n127) );
  COND1X1 U939 ( .A(n154), .B(n144), .C(n145), .Z(n139) );
  CANR1XL U940 ( .A(n645), .B(n183), .C(n174), .Z(n172) );
  CANR1X1 U941 ( .A(n183), .B(net14710), .C(n165), .Z(net14384) );
  CNR2XL U942 ( .A(n175), .B(n166), .Z(net14710) );
  CIVXL U943 ( .A(net14584), .Z(net14129) );
  CND2IXL U944 ( .B(n129), .A(n132), .Z(n10) );
  CNR2X1 U945 ( .A(B[56]), .B(A[56]), .Z(n129) );
  CNR2X1 U946 ( .A(n129), .B(n120), .Z(n118) );
  CND2X1 U947 ( .A(B[56]), .B(A[56]), .Z(n132) );
  CNR2X1 U948 ( .A(B[44]), .B(A[44]), .Z(n251) );
  CIVXL U949 ( .A(n268), .Z(n266) );
  CND2X1 U950 ( .A(B[44]), .B(A[44]), .Z(n254) );
  CNR2X2 U951 ( .A(B[51]), .B(A[51]), .Z(n188) );
  CND2X1 U952 ( .A(B[51]), .B(A[51]), .Z(n189) );
  CIVX1 U953 ( .A(n357), .Z(n664) );
  CNR2X1 U954 ( .A(B[33]), .B(A[33]), .Z(n357) );
  CND2X1 U955 ( .A(n664), .B(n665), .Z(n349) );
  CANR1X2 U956 ( .A(n901), .B(n664), .C(net14087), .Z(n350) );
  CND2XL U957 ( .A(n898), .B(net13631), .Z(n33) );
  CAN2X1 U958 ( .A(B[33]), .B(A[33]), .Z(net14087) );
  CIVXL U959 ( .A(n899), .Z(n352) );
  CNR2X1 U960 ( .A(B[38]), .B(A[38]), .Z(n304) );
  CND2IX1 U961 ( .B(n337), .A(net14085), .Z(n915) );
  CND2XL U962 ( .A(n288), .B(n26), .Z(n917) );
  CND2X1 U963 ( .A(n916), .B(net14721), .Z(n918) );
  CND2X1 U964 ( .A(n918), .B(n917), .Z(SUM[40]) );
  CIVXL U965 ( .A(n288), .Z(n916) );
  CIVX2 U966 ( .A(n26), .Z(net14721) );
  COND1X1 U967 ( .A(n289), .B(n366), .C(n290), .Z(n288) );
  CIVX1 U968 ( .A(n610), .Z(n609) );
  CND2X1 U969 ( .A(net14098), .B(net14090), .Z(n372) );
  CND2X2 U970 ( .A(n669), .B(n668), .Z(n392) );
  CIVX1 U971 ( .A(n360), .Z(n665) );
  CNR2X2 U972 ( .A(B[37]), .B(A[37]), .Z(net14690) );
  CNR2X2 U973 ( .A(B[37]), .B(A[37]), .Z(n315) );
  CIVXL U974 ( .A(n492), .Z(n491) );
  CND2XL U975 ( .A(n962), .B(n625), .Z(n63) );
  CANR1X2 U976 ( .A(n593), .B(n955), .C(n586), .Z(n580) );
  CENX1 U977 ( .A(n919), .B(n235), .Z(SUM[46]) );
  CAN2XL U978 ( .A(n651), .B(n234), .Z(n919) );
  CIVXL U979 ( .A(n144), .Z(n642) );
  COND1X2 U980 ( .A(n497), .B(n505), .C(n498), .Z(n496) );
  CIVXL U981 ( .A(n182), .Z(n180) );
  CIVX1 U982 ( .A(n489), .Z(n678) );
  CIVXL U983 ( .A(n484), .Z(n482) );
  CIVXL U984 ( .A(n326), .Z(net14628) );
  CIVXL U985 ( .A(n153), .Z(n643) );
  CANR1X1 U986 ( .A(n606), .B(n959), .C(n601), .Z(n599) );
  CIVXL U987 ( .A(n321), .Z(net14622) );
  CND2X2 U988 ( .A(n689), .B(n955), .Z(n579) );
  CNR2X1 U989 ( .A(B[46]), .B(A[46]), .Z(n231) );
  COND1X1 U990 ( .A(n149), .B(n201), .C(n150), .Z(n148) );
  CIVXL U991 ( .A(n327), .Z(n325) );
  CIVXL U992 ( .A(n120), .Z(n640) );
  CND2XL U993 ( .A(B[30]), .B(A[30]), .Z(n388) );
  CIVXL U994 ( .A(n352), .Z(net14588) );
  CNR2X2 U995 ( .A(B[29]), .B(A[29]), .Z(n400) );
  CND2X1 U996 ( .A(n958), .B(n953), .Z(n436) );
  CENXL U997 ( .A(n348), .B(n32), .Z(SUM[34]) );
  CND2X1 U998 ( .A(B[46]), .B(A[46]), .Z(n234) );
  CND2X1 U999 ( .A(B[47]), .B(A[47]), .Z(n227) );
  CIVX1 U1000 ( .A(n322), .Z(n661) );
  CIVXL U1001 ( .A(n568), .Z(n566) );
  CND2XL U1002 ( .A(n661), .B(net14622), .Z(n30) );
  CANR1X2 U1003 ( .A(n448), .B(n953), .C(n443), .Z(n437) );
  CND2X1 U1004 ( .A(B[52]), .B(A[52]), .Z(n176) );
  CENXL U1005 ( .A(n299), .B(n27), .Z(SUM[39]) );
  CENX1 U1006 ( .A(n921), .B(n106), .Z(SUM[59]) );
  CNR2XL U1007 ( .A(B[2]), .B(A[2]), .Z(n627) );
  CEOX1 U1008 ( .A(n939), .B(n146), .Z(SUM[55]) );
  CIVXL U1009 ( .A(n166), .Z(n644) );
  COR2XL U1010 ( .A(B[45]), .B(A[45]), .Z(n920) );
  CND2X2 U1011 ( .A(B[42]), .B(A[42]), .Z(n268) );
  COND1X2 U1012 ( .A(n254), .B(n246), .C(n247), .Z(n245) );
  COND1X2 U1013 ( .A(n268), .B(n262), .C(n263), .Z(n257) );
  CIVXL U1014 ( .A(n208), .Z(n648) );
  COND1X2 U1015 ( .A(n598), .B(n610), .C(n599), .Z(n597) );
  CENXL U1016 ( .A(n306), .B(n28), .Z(SUM[38]) );
  CANR1X2 U1017 ( .A(n556), .B(n684), .C(n551), .Z(n545) );
  CND2X1 U1018 ( .A(B[50]), .B(A[50]), .Z(n196) );
  CIVXL U1019 ( .A(n323), .Z(n321) );
  CNR2X2 U1020 ( .A(B[52]), .B(A[52]), .Z(n175) );
  CAN2XL U1021 ( .A(net14046), .B(n105), .Z(n921) );
  CNR2XL U1022 ( .A(n220), .B(n213), .Z(n211) );
  CND2X2 U1023 ( .A(B[37]), .B(A[37]), .Z(n316) );
  CND2X2 U1024 ( .A(n13), .B(n923), .Z(n924) );
  CND2XL U1025 ( .A(n168), .B(n922), .Z(n925) );
  CND2X2 U1026 ( .A(n924), .B(n925), .Z(SUM[53]) );
  CIVX2 U1027 ( .A(n13), .Z(n922) );
  CIVX1 U1028 ( .A(n168), .Z(n923) );
  CANR1X1 U1029 ( .A(n169), .B(net26801), .C(n170), .Z(n168) );
  CND2X2 U1030 ( .A(n927), .B(n9), .Z(n928) );
  CND2XL U1031 ( .A(n122), .B(n926), .Z(n929) );
  CND2X2 U1032 ( .A(n929), .B(n928), .Z(SUM[57]) );
  CIVX2 U1033 ( .A(n9), .Z(n926) );
  CIVX1 U1034 ( .A(n122), .Z(n927) );
  CND2XL U1035 ( .A(n640), .B(n121), .Z(n9) );
  CND2X2 U1036 ( .A(n12), .B(n931), .Z(n932) );
  CND2XL U1037 ( .A(n155), .B(n930), .Z(n933) );
  CND2X2 U1038 ( .A(n932), .B(n933), .Z(SUM[54]) );
  CIVX2 U1039 ( .A(n12), .Z(n930) );
  CIVX1 U1040 ( .A(n155), .Z(n931) );
  CANR1X1 U1041 ( .A(n156), .B(net26801), .C(n157), .Z(n155) );
  CANR1XL U1042 ( .A(n661), .B(net14628), .C(n321), .Z(n319) );
  CIVXL U1043 ( .A(n257), .Z(n259) );
  CIVXL U1044 ( .A(n304), .Z(n659) );
  CIVXL U1045 ( .A(n436), .Z(n434) );
  COND1XL U1046 ( .A(n349), .B(n366), .C(net14588), .Z(n348) );
  CANR1X1 U1047 ( .A(n147), .B(n269), .C(n148), .Z(n146) );
  CND2X2 U1048 ( .A(n681), .B(n680), .Z(n502) );
  CANR1X2 U1049 ( .A(n516), .B(n680), .C(n507), .Z(n505) );
  CIVX2 U1050 ( .A(n514), .Z(n516) );
  CND2X1 U1051 ( .A(B[29]), .B(A[29]), .Z(n401) );
  CND2X1 U1052 ( .A(n964), .B(n8), .Z(n936) );
  CIVX1 U1053 ( .A(n964), .Z(n934) );
  CND2XL U1054 ( .A(n962), .B(n695), .Z(n620) );
  CANR1X2 U1055 ( .A(n630), .B(n962), .C(n623), .Z(n621) );
  CND2X1 U1056 ( .A(net14130), .B(net14626), .Z(n964) );
  CIVXL U1057 ( .A(n8), .Z(n935) );
  CNR2XL U1058 ( .A(n436), .B(n418), .Z(n412) );
  CND2X1 U1059 ( .A(n934), .B(n935), .Z(n937) );
  CND2X2 U1060 ( .A(n936), .B(n937), .Z(SUM[58]) );
  CAN2XL U1061 ( .A(n636), .B(n85), .Z(n938) );
  CENXL U1062 ( .A(n938), .B(n86), .Z(SUM[61]) );
  CND2XL U1063 ( .A(net14094), .B(n110), .Z(n8) );
  CNR2X1 U1064 ( .A(n175), .B(n166), .Z(n164) );
  CNR2XL U1065 ( .A(n895), .B(n381), .Z(n379) );
  CANR1X1 U1066 ( .A(n430), .B(n954), .C(n421), .Z(n419) );
  CENX1 U1067 ( .A(n947), .B(n940), .Z(SUM[62]) );
  CANR1XL U1068 ( .A(n542), .B(n559), .C(n543), .Z(n541) );
  COND1XL U1069 ( .A(n300), .B(n366), .C(n301), .Z(n299) );
  COND1XL U1070 ( .A(n340), .B(n366), .C(n341), .Z(n339) );
  CANR1X1 U1071 ( .A(n575), .B(n966), .C(n566), .Z(n564) );
  COR2X1 U1072 ( .A(B[58]), .B(A[58]), .Z(net14094) );
  CEOX2 U1073 ( .A(n944), .B(n228), .Z(SUM[47]) );
  CND2XL U1074 ( .A(B[18]), .B(A[18]), .Z(n498) );
  CNR2X1 U1075 ( .A(B[22]), .B(A[22]), .Z(n468) );
  CND2X1 U1076 ( .A(n484), .B(n894), .Z(n471) );
  CANR1XL U1077 ( .A(n952), .B(n964), .C(n903), .Z(n945) );
  CENXL U1078 ( .A(n960), .B(n945), .Z(SUM[63]) );
  CND2X1 U1079 ( .A(B[20]), .B(A[20]), .Z(n487) );
  CNR2X1 U1080 ( .A(n946), .B(n489), .Z(n484) );
  CNR2XL U1081 ( .A(B[20]), .B(A[20]), .Z(n946) );
  CNR2X1 U1082 ( .A(n522), .B(n502), .Z(n500) );
  CANR1X1 U1083 ( .A(n123), .B(net26801), .C(n124), .Z(n122) );
  CND2XL U1084 ( .A(n644), .B(n167), .Z(n13) );
  CAN2XL U1085 ( .A(n646), .B(n189), .Z(n949) );
  CND2XL U1086 ( .A(n642), .B(n145), .Z(n939) );
  CIVXL U1087 ( .A(n176), .Z(n174) );
  CIVX1 U1088 ( .A(n588), .Z(n586) );
  CND2XL U1089 ( .A(n693), .B(n617), .Z(n62) );
  CND2XL U1090 ( .A(n689), .B(n591), .Z(n58) );
  CND2XL U1091 ( .A(n678), .B(n490), .Z(n47) );
  CENXL U1092 ( .A(n941), .B(n519), .Z(SUM[16]) );
  CAN2XL U1093 ( .A(n681), .B(n514), .Z(n941) );
  CEOXL U1094 ( .A(n59), .B(n604), .Z(SUM[7]) );
  CND2XL U1095 ( .A(n959), .B(n603), .Z(n59) );
  CEOXL U1096 ( .A(n35), .B(n378), .Z(SUM[31]) );
  CND2XL U1097 ( .A(net14090), .B(n377), .Z(n35) );
  CNR2XL U1098 ( .A(n613), .B(n616), .Z(n611) );
  CEOXL U1099 ( .A(n41), .B(n446), .Z(SUM[25]) );
  CND2XL U1100 ( .A(n953), .B(n445), .Z(n41) );
  CEOXL U1101 ( .A(n39), .B(n424), .Z(SUM[27]) );
  CND2XL U1102 ( .A(n954), .B(n423), .Z(n39) );
  CNR2XL U1103 ( .A(n436), .B(n427), .Z(n425) );
  CEOXL U1104 ( .A(n37), .B(n402), .Z(SUM[29]) );
  CEOXL U1105 ( .A(n53), .B(n554), .Z(SUM[13]) );
  CEOXL U1106 ( .A(n48), .B(n499), .Z(SUM[18]) );
  CND2XL U1107 ( .A(n581), .B(n687), .Z(n570) );
  CND2XL U1108 ( .A(n955), .B(n588), .Z(n57) );
  CEOXL U1109 ( .A(n451), .B(n942), .Z(SUM[24]) );
  CAN2XL U1110 ( .A(n958), .B(n450), .Z(n942) );
  CND2XL U1111 ( .A(n687), .B(n577), .Z(n56) );
  CND2XL U1112 ( .A(n957), .B(n608), .Z(n60) );
  CND2XL U1113 ( .A(n647), .B(n196), .Z(n16) );
  CND2XL U1114 ( .A(n671), .B(n428), .Z(n40) );
  CND2XL U1115 ( .A(net14098), .B(n388), .Z(n36) );
  CEOX1 U1116 ( .A(n943), .B(n264), .Z(SUM[43]) );
  CND2XL U1117 ( .A(n654), .B(n263), .Z(n943) );
  CND2IXL U1118 ( .B(n392), .A(net14098), .Z(n381) );
  CIVX1 U1119 ( .A(n76), .Z(n74) );
  CNR2XL U1120 ( .A(B[19]), .B(A[19]), .Z(n489) );
  CEOXL U1121 ( .A(n64), .B(n1), .Z(SUM[2]) );
  CND2XL U1122 ( .A(n650), .B(n227), .Z(n944) );
  CNR2XL U1123 ( .A(B[32]), .B(A[32]), .Z(n360) );
  CND2XL U1124 ( .A(B[61]), .B(A[61]), .Z(n85) );
  CND2XL U1125 ( .A(B[5]), .B(A[5]), .Z(n614) );
  COR2XL U1126 ( .A(B[24]), .B(A[24]), .Z(n958) );
  COR2XL U1127 ( .A(B[63]), .B(A[63]), .Z(n963) );
  CNR2XL U1128 ( .A(n200), .B(n125), .Z(n123) );
  CNR2XL U1129 ( .A(n200), .B(n171), .Z(n169) );
  CNR2XL U1130 ( .A(n200), .B(n149), .Z(n147) );
  CENX1 U1131 ( .A(n559), .B(n54), .Z(SUM[12]) );
  CEOXL U1132 ( .A(n34), .B(net26798), .Z(SUM[32]) );
  CND2XL U1133 ( .A(n665), .B(net13575), .Z(n34) );
  COND1XL U1134 ( .A(n158), .B(n201), .C(net14384), .Z(n157) );
  CNR2X2 U1135 ( .A(n238), .B(n204), .Z(n198) );
  COND1XL U1136 ( .A(n570), .B(n596), .C(n571), .Z(n569) );
  CENX1 U1137 ( .A(n279), .B(n25), .Z(SUM[41]) );
  COND1XL U1138 ( .A(n280), .B(n366), .C(n281), .Z(n279) );
  CENX1 U1139 ( .A(n317), .B(n29), .Z(SUM[37]) );
  COND1XL U1140 ( .A(n318), .B(n366), .C(n319), .Z(n317) );
  CENX1 U1141 ( .A(n470), .B(n44), .Z(SUM[22]) );
  CND2XL U1142 ( .A(n675), .B(n469), .Z(n44) );
  COND1XL U1143 ( .A(n471), .B(n491), .C(n472), .Z(n470) );
  CENX1 U1144 ( .A(n461), .B(n43), .Z(SUM[23]) );
  COND1XL U1145 ( .A(n462), .B(n491), .C(n463), .Z(n461) );
  CND2XL U1146 ( .A(n473), .B(n675), .Z(n462) );
  CENX1 U1147 ( .A(n578), .B(n56), .Z(SUM[10]) );
  COND1XL U1148 ( .A(n579), .B(n596), .C(n580), .Z(n578) );
  CENX1 U1149 ( .A(n609), .B(n60), .Z(SUM[6]) );
  CENX1 U1150 ( .A(n589), .B(n57), .Z(SUM[9]) );
  COND1XL U1151 ( .A(n590), .B(n596), .C(n591), .Z(n589) );
  CENX1 U1152 ( .A(n615), .B(n61), .Z(SUM[5]) );
  CND2X1 U1153 ( .A(n692), .B(n614), .Z(n61) );
  COND1XL U1154 ( .A(n616), .B(n618), .C(n617), .Z(n615) );
  CNR2X1 U1155 ( .A(n200), .B(n180), .Z(n178) );
  CAN2X1 U1156 ( .A(n956), .B(n76), .Z(n947) );
  CANR1XL U1157 ( .A(n87), .B(n964), .C(n88), .Z(n86) );
  CEOX1 U1158 ( .A(n16), .B(n197), .Z(SUM[50]) );
  CENX1 U1159 ( .A(n948), .B(n210), .Z(SUM[49]) );
  CAN2X1 U1160 ( .A(n648), .B(n209), .Z(n948) );
  CENX1 U1161 ( .A(n949), .B(n190), .Z(SUM[51]) );
  CEOX1 U1162 ( .A(n40), .B(n433), .Z(SUM[26]) );
  CANR1XL U1163 ( .A(n958), .B(n451), .C(n448), .Z(n446) );
  CEOX1 U1164 ( .A(n38), .B(n411), .Z(SUM[28]) );
  CND2XL U1165 ( .A(n669), .B(n406), .Z(n38) );
  CEOX1 U1166 ( .A(n36), .B(n389), .Z(SUM[30]) );
  CANR1XL U1167 ( .A(n425), .B(n451), .C(n426), .Z(n424) );
  CANR1XL U1168 ( .A(n379), .B(n451), .C(n380), .Z(n378) );
  CANR1XL U1169 ( .A(n403), .B(n451), .C(n404), .Z(n402) );
  CNR2XL U1170 ( .A(n895), .B(n405), .Z(n403) );
  CND2X1 U1171 ( .A(n679), .B(n498), .Z(n48) );
  CANR1XL U1172 ( .A(n500), .B(n559), .C(n501), .Z(n499) );
  CEOX1 U1173 ( .A(n51), .B(n532), .Z(SUM[15]) );
  CND2XL U1174 ( .A(n682), .B(n531), .Z(n51) );
  CANR1XL U1175 ( .A(n533), .B(n559), .C(n534), .Z(n532) );
  CEOX1 U1176 ( .A(n52), .B(n541), .Z(SUM[14]) );
  CND2XL U1177 ( .A(n683), .B(n536), .Z(n52) );
  CEOX1 U1178 ( .A(n49), .B(n510), .Z(SUM[17]) );
  CND2XL U1179 ( .A(n509), .B(n680), .Z(n49) );
  CANR1XL U1180 ( .A(n511), .B(n559), .C(n512), .Z(n510) );
  CND2XL U1181 ( .A(n684), .B(n553), .Z(n53) );
  CANR1XL U1182 ( .A(n951), .B(n559), .C(n556), .Z(n554) );
  CEOXL U1183 ( .A(n47), .B(n491), .Z(SUM[19]) );
  CEOXL U1184 ( .A(n62), .B(n618), .Z(SUM[4]) );
  CEOXL U1185 ( .A(n58), .B(n596), .Z(SUM[8]) );
  CANR1XL U1186 ( .A(n957), .B(n609), .C(n606), .Z(n604) );
  CANR1X1 U1187 ( .A(n611), .B(n619), .C(n612), .Z(n610) );
  COND1XL U1188 ( .A(n617), .B(n613), .C(n614), .Z(n612) );
  CND2XL U1189 ( .A(n643), .B(n154), .Z(n12) );
  CNR2XL U1190 ( .A(n200), .B(n158), .Z(n156) );
  COAN1X1 U1191 ( .A(n406), .B(n400), .C(n401), .Z(n393) );
  CNR2IXL U1192 ( .B(n256), .A(n251), .Z(n249) );
  CNR2X1 U1193 ( .A(n579), .B(n563), .Z(n561) );
  CND2X1 U1194 ( .A(n959), .B(n957), .Z(n598) );
  COND1XL U1195 ( .A(n360), .B(n366), .C(net13575), .Z(n359) );
  CENX1 U1196 ( .A(n950), .B(n217), .Z(SUM[48]) );
  CAN2X1 U1197 ( .A(n649), .B(n216), .Z(n950) );
  CANR1XL U1198 ( .A(n659), .B(net19921), .C(n303), .Z(n301) );
  CANR1XL U1199 ( .A(n675), .B(n474), .C(n467), .Z(n463) );
  CANR1XL U1200 ( .A(n687), .B(n582), .C(n575), .Z(n571) );
  COND1XL U1201 ( .A(n125), .B(n201), .C(n126), .Z(n124) );
  COND1XL U1202 ( .A(n171), .B(n201), .C(n172), .Z(n170) );
  COND1XL U1203 ( .A(n381), .B(n415), .C(n382), .Z(n380) );
  COND1XL U1204 ( .A(n405), .B(n415), .C(n406), .Z(n404) );
  CNR2X2 U1205 ( .A(n502), .B(n497), .Z(n495) );
  CND2X1 U1206 ( .A(n671), .B(n954), .Z(n418) );
  CIVX2 U1207 ( .A(n513), .Z(n681) );
  CND2XL U1208 ( .A(n282), .B(n309), .Z(n280) );
  CAN2XL U1209 ( .A(n78), .B(n956), .Z(n952) );
  COND1XL U1210 ( .A(n482), .B(n491), .C(n483), .Z(n481) );
  COND1XL U1211 ( .A(n489), .B(n491), .C(n490), .Z(n488) );
  CENX1 U1212 ( .A(n626), .B(n63), .Z(SUM[3]) );
  COND1XL U1213 ( .A(n627), .B(n1), .C(n628), .Z(n626) );
  CND2XL U1214 ( .A(n695), .B(n628), .Z(n64) );
  CNR2X1 U1215 ( .A(B[28]), .B(A[28]), .Z(n405) );
  CNR2X1 U1216 ( .A(B[4]), .B(A[4]), .Z(n616) );
  CNR2X1 U1217 ( .A(B[61]), .B(A[61]), .Z(n84) );
  CNR2X1 U1218 ( .A(B[5]), .B(A[5]), .Z(n613) );
  CNR2X1 U1219 ( .A(B[26]), .B(A[26]), .Z(n427) );
  CNR2X1 U1220 ( .A(B[42]), .B(A[42]), .Z(n267) );
  CNR2X1 U1221 ( .A(B[54]), .B(A[54]), .Z(n153) );
  CNR2X1 U1222 ( .A(B[16]), .B(A[16]), .Z(n513) );
  CNR2X2 U1223 ( .A(B[57]), .B(A[57]), .Z(n120) );
  COR2X1 U1224 ( .A(B[30]), .B(A[30]), .Z(net14098) );
  CNR2X1 U1225 ( .A(B[14]), .B(A[14]), .Z(n535) );
  COR2X1 U1226 ( .A(B[25]), .B(A[25]), .Z(n953) );
  COR2X1 U1227 ( .A(B[27]), .B(A[27]), .Z(n954) );
  COR2X1 U1228 ( .A(B[9]), .B(A[9]), .Z(n955) );
  CND2X1 U1229 ( .A(B[54]), .B(A[54]), .Z(n154) );
  COR2X1 U1230 ( .A(B[62]), .B(A[62]), .Z(n956) );
  COR2X1 U1231 ( .A(B[6]), .B(A[6]), .Z(n957) );
  COR2X1 U1232 ( .A(A[31]), .B(B[31]), .Z(net14090) );
  CND2X1 U1233 ( .A(B[28]), .B(A[28]), .Z(n406) );
  CND2X1 U1234 ( .A(B[8]), .B(A[8]), .Z(n591) );
  CND2X1 U1235 ( .A(B[2]), .B(A[2]), .Z(n628) );
  COR2X1 U1236 ( .A(B[7]), .B(A[7]), .Z(n959) );
  CND2X1 U1237 ( .A(B[48]), .B(A[48]), .Z(n216) );
  CND2X1 U1238 ( .A(B[26]), .B(A[26]), .Z(n428) );
  CND2X1 U1239 ( .A(B[16]), .B(A[16]), .Z(n514) );
  CND2X1 U1240 ( .A(B[14]), .B(A[14]), .Z(n536) );
  CND2X1 U1241 ( .A(B[4]), .B(A[4]), .Z(n617) );
  CND2X1 U1242 ( .A(B[58]), .B(A[58]), .Z(n110) );
  CND2X1 U1243 ( .A(B[62]), .B(A[62]), .Z(n76) );
  CND2X1 U1244 ( .A(B[22]), .B(A[22]), .Z(n469) );
  CND2X1 U1245 ( .A(B[24]), .B(A[24]), .Z(n450) );
  CND2X1 U1246 ( .A(B[25]), .B(A[25]), .Z(n445) );
  CND2X1 U1247 ( .A(B[27]), .B(A[27]), .Z(n423) );
  CND2X1 U1248 ( .A(B[31]), .B(A[31]), .Z(n377) );
  CND2X1 U1249 ( .A(B[9]), .B(A[9]), .Z(n588) );
  CND2X1 U1250 ( .A(B[10]), .B(A[10]), .Z(n577) );
  CND2X1 U1251 ( .A(B[7]), .B(A[7]), .Z(n603) );
  CND2X1 U1252 ( .A(B[6]), .B(A[6]), .Z(n608) );
  CNR2XL U1253 ( .A(n238), .B(n909), .Z(n229) );
  CND2X1 U1254 ( .A(B[23]), .B(A[23]), .Z(n460) );
  CAN2X1 U1255 ( .A(n963), .B(n67), .Z(n960) );
  CND2X1 U1256 ( .A(A[1]), .B(B[1]), .Z(n1) );
  CAN2XL U1257 ( .A(n905), .B(n1), .Z(SUM[1]) );
  COR2X1 U1258 ( .A(B[59]), .B(A[59]), .Z(net14046) );
  COR2X1 U1259 ( .A(B[3]), .B(A[3]), .Z(n962) );
  CND2X1 U1260 ( .A(B[59]), .B(A[59]), .Z(n105) );
  CND2X1 U1261 ( .A(B[3]), .B(A[3]), .Z(n625) );
  CND2X1 U1262 ( .A(n240), .B(n222), .Z(n220) );
  COND1XL U1263 ( .A(n427), .B(n437), .C(n428), .Z(n426) );
  CANR1X2 U1264 ( .A(n538), .B(n682), .C(n529), .Z(n527) );
  CND2XL U1265 ( .A(n902), .B(n460), .Z(n43) );
  CND2X2 U1266 ( .A(n951), .B(n684), .Z(n544) );
  COND1XL U1267 ( .A(n213), .B(n221), .C(n216), .Z(n212) );
  CIVXL U1268 ( .A(n213), .Z(n649) );
  CANR1XL U1269 ( .A(n282), .B(net19921), .C(n283), .Z(n281) );
  CIVXL U1270 ( .A(n485), .Z(n483) );
  COND1X1 U1271 ( .A(n490), .B(n486), .C(n487), .Z(n485) );
  CND2X2 U1272 ( .A(n520), .B(n495), .Z(n493) );
  CIVXL U1273 ( .A(n251), .Z(n653) );
  COND1XL U1274 ( .A(n251), .B(n259), .C(n254), .Z(n250) );
  COND1X2 U1275 ( .A(n526), .B(n545), .C(n527), .Z(n521) );
  CANR1X2 U1276 ( .A(n495), .B(n521), .C(n496), .Z(n494) );
  CND2X1 U1277 ( .A(B[43]), .B(A[43]), .Z(n263) );
  CNR2X2 U1278 ( .A(n267), .B(n262), .Z(n256) );
  CIVXL U1279 ( .A(n521), .Z(n523) );
  CND2X1 U1280 ( .A(n182), .B(n645), .Z(n171) );
  CIVXL U1281 ( .A(n262), .Z(n654) );
  CND2X1 U1282 ( .A(B[39]), .B(A[39]), .Z(n298) );
  CIVXL U1283 ( .A(n239), .Z(n241) );
  COND1X2 U1284 ( .A(n493), .B(n560), .C(n494), .Z(n492) );
  CIVXL U1285 ( .A(n472), .Z(n474) );
  CND2X1 U1286 ( .A(B[15]), .B(A[15]), .Z(n531) );
  CANR1X2 U1287 ( .A(n597), .B(n561), .C(n562), .Z(n560) );
  COND1XL U1288 ( .A(n535), .B(n545), .C(n536), .Z(n534) );
  COND1XL U1289 ( .A(n910), .B(n201), .C(n196), .Z(n192) );
  CNR2XL U1290 ( .A(n200), .B(n910), .Z(n191) );
  CIVXL U1291 ( .A(n193), .Z(n647) );
  CNR2X1 U1292 ( .A(B[50]), .B(A[50]), .Z(n193) );
  CND2XL U1293 ( .A(n894), .B(n480), .Z(n45) );
  CND2X1 U1294 ( .A(B[21]), .B(A[21]), .Z(n480) );
  CENX1 U1295 ( .A(n481), .B(n45), .Z(SUM[21]) );
  CNR2XL U1296 ( .A(B[20]), .B(A[20]), .Z(n965) );
  CNR2X1 U1297 ( .A(B[20]), .B(A[20]), .Z(n486) );
  CNR2X1 U1298 ( .A(n895), .B(n392), .Z(n390) );
  CIVX2 U1299 ( .A(n400), .Z(n668) );
  CIVXL U1300 ( .A(net14087), .Z(net13631) );
  CND2XL U1301 ( .A(n668), .B(n401), .Z(n37) );
  CND2XL U1302 ( .A(n897), .B(n568), .Z(n55) );
  CENX1 U1303 ( .A(n569), .B(n55), .Z(SUM[11]) );
  CENX1 U1304 ( .A(n324), .B(n30), .Z(SUM[36]) );
  CND2XL U1305 ( .A(n327), .B(n661), .Z(n318) );
  CND2XL U1306 ( .A(n309), .B(net14742), .Z(n289) );
  CND2X1 U1307 ( .A(n309), .B(n659), .Z(n300) );
  CND2X1 U1308 ( .A(B[38]), .B(A[38]), .Z(n305) );
  CENX1 U1309 ( .A(n359), .B(n33), .Z(SUM[33]) );
  CNR2X1 U1310 ( .A(B[13]), .B(A[13]), .Z(n552) );
  CND2X1 U1311 ( .A(B[13]), .B(A[13]), .Z(n553) );
  CND2XL U1312 ( .A(n660), .B(n316), .Z(n29) );
  CIVXL U1313 ( .A(n544), .Z(n542) );
  CNR2XL U1314 ( .A(n544), .B(n535), .Z(n533) );
  CND2XL U1315 ( .A(net14085), .B(n347), .Z(n32) );
  CND2X1 U1316 ( .A(B[34]), .B(A[34]), .Z(n347) );
  CND2X1 U1317 ( .A(B[53]), .B(A[53]), .Z(n167) );
  COND1XL U1318 ( .A(n502), .B(n523), .C(n505), .Z(n501) );
  CIVX1 U1319 ( .A(n901), .Z(net13575) );
  CND2X1 U1320 ( .A(B[49]), .B(A[49]), .Z(n209) );
  CIVXL U1321 ( .A(n188), .Z(n646) );
  COND1XL U1322 ( .A(n909), .B(n239), .C(n234), .Z(n230) );
  CND2X1 U1323 ( .A(B[45]), .B(A[45]), .Z(n247) );
  CIVXL U1324 ( .A(net14690), .Z(n660) );
  CANR1XL U1325 ( .A(n520), .B(n559), .C(n521), .Z(n519) );
  CND2X1 U1326 ( .A(B[12]), .B(A[12]), .Z(n558) );
  CNR2XL U1327 ( .A(n522), .B(n513), .Z(n511) );
  COND1XL U1328 ( .A(n513), .B(n523), .C(n514), .Z(n512) );
  CIVX1 U1329 ( .A(n560), .Z(n559) );
  CANR1X2 U1330 ( .A(n257), .B(n244), .C(n245), .Z(n239) );
  CND2X1 U1331 ( .A(n951), .B(n558), .Z(n54) );
  CANR1X2 U1332 ( .A(n453), .B(n492), .C(n454), .Z(n452) );
  CIVX2 U1333 ( .A(n616), .Z(n693) );
  CIVX2 U1334 ( .A(n613), .Z(n692) );
  CIVX2 U1335 ( .A(n497), .Z(n679) );
  CIVX2 U1336 ( .A(n965), .Z(n677) );
  CIVX2 U1337 ( .A(n84), .Z(n636) );
  CIVX2 U1338 ( .A(n628), .Z(n630) );
  CIVX2 U1339 ( .A(n627), .Z(n695) );
  CIVX2 U1340 ( .A(n625), .Z(n623) );
  CIVX2 U1341 ( .A(n619), .Z(n618) );
  CIVX2 U1342 ( .A(n608), .Z(n606) );
  CIVX2 U1343 ( .A(n603), .Z(n601) );
  CIVX2 U1344 ( .A(n597), .Z(n596) );
  CIVX2 U1345 ( .A(n591), .Z(n593) );
  CIVX2 U1346 ( .A(n590), .Z(n689) );
  CIVX2 U1347 ( .A(n580), .Z(n582) );
  CIVX2 U1348 ( .A(n579), .Z(n581) );
  CIVX2 U1349 ( .A(n576), .Z(n687) );
  CIVX2 U1350 ( .A(n558), .Z(n556) );
  CIVX2 U1351 ( .A(n553), .Z(n551) );
  CIVX2 U1352 ( .A(n536), .Z(n538) );
  CIVX2 U1353 ( .A(n535), .Z(n683) );
  CIVX2 U1354 ( .A(n531), .Z(n529) );
  CIVX2 U1355 ( .A(n530), .Z(n682) );
  CIVX2 U1356 ( .A(n520), .Z(n522) );
  CIVX2 U1357 ( .A(n509), .Z(n507) );
  CIVX2 U1358 ( .A(n508), .Z(n680) );
  CIVX2 U1359 ( .A(n480), .Z(n478) );
  CIVX2 U1360 ( .A(n471), .Z(n473) );
  CIVX2 U1361 ( .A(n469), .Z(n467) );
  CIVX2 U1362 ( .A(n468), .Z(n675) );
  CIVX2 U1363 ( .A(n460), .Z(n458) );
  CIVX2 U1364 ( .A(n450), .Z(n448) );
  CIVX2 U1365 ( .A(n445), .Z(n443) );
  CIVX2 U1366 ( .A(n428), .Z(n430) );
  CIVX2 U1367 ( .A(n427), .Z(n671) );
  CIVX2 U1368 ( .A(n423), .Z(n421) );
  CIVX2 U1369 ( .A(n405), .Z(n669) );
  CIVX2 U1370 ( .A(n349), .Z(n351) );
  CIVX2 U1371 ( .A(n238), .Z(n240) );
  CIVX2 U1372 ( .A(n221), .Z(n219) );
  CIVX2 U1373 ( .A(n220), .Z(n218) );
  CIVX2 U1374 ( .A(n175), .Z(n645) );
  CIVX2 U1375 ( .A(n154), .Z(n152) );
endmodule


module sqrt64_DW_cmp_4 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [63:0] A;
  input [63:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n34, n56, n58, n60, n62, n70, n87, n89, n91, n93, n107, n109, n117,
         n129, n154, n156, n158, n160, n164, n172, n176, n199, n207, n222,
         n312, n316, n320, n322, n325, n326, n327, n328, n329, n330, n331,
         n333, n334, n335, n336, n340, n342, n346, n348, n350, net14039,
         net14042, n99, n98, n97, n96, n95, n94, n92, n90, n88, n86, n85, n84,
         n83, n82, n81, n80, n79, n78, n77, n76, n75, n74, n73, n72, n71, n69,
         n68, n67, n66, n65, n63, n61, n59, n57, n55, n54, n53, n52, n51, n50,
         n5, n49, n48, n351, n349, n347, n345, n344, n343, n341, n339, n338,
         n337, n332, n324, n323, n321, n319, n318, n317, n315, n314, n313,
         n311, n310, n309, n308, n307, n306, n305, n304, n303, n302, n301,
         n300, n3, n299, n298, n297, n296, n294, n293, n290, n289, n288, n286,
         n285, n282, n280, n273, n272, n271, n270, n269, n268, n267, n266,
         n265, n264, n262, n255, n254, n253, n244, n243, n238, n236, n234,
         n233, n232, n231, n230, n229, n228, n227, n226, n225, n224, n223,
         n221, n220, n219, n218, n217, n216, n215, n214, n213, n212, n211,
         n210, n209, n208, n206, n205, n204, n203, n202, n201, n192, n191,
         n190, n189, n188, n18, n179, n178, n170, n169, n168, n167, n166, n16,
         n157, n147, n146, n145, n144, n143, n142, n141, n132, n131, n122,
         n121, n120, n119, n110, n100, n1, n46, n44, n42, n352, net19772, n6,
         n4, n362, n361, n360, n2, n15, n17, net23082, net14590, n32, n30, n28,
         n26, n20, n47, n45, n43, n358, n357, n356, n353, n35, n33, n31, n29,
         n27, n23, n21, n19, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767;

  CNR2X2 U57 ( .A(A[51]), .B(n350), .Z(n56) );
  CNR2X2 U59 ( .A(n62), .B(n60), .Z(n58) );
  CNR2X2 U71 ( .A(A[47]), .B(n346), .Z(n70) );
  CNR2X2 U161 ( .A(A[30]), .B(n329), .Z(n160) );
  COND1X1 U54 ( .A(n57), .B(n54), .C(n55), .Z(n53) );
  CNR2X2 U53 ( .A(n56), .B(n54), .Z(n52) );
  CNR2X2 U61 ( .A(A[50]), .B(n349), .Z(n60) );
  COND1X1 U60 ( .A(n63), .B(n60), .C(n61), .Z(n59) );
  CANR1X1 U52 ( .A(n59), .B(n52), .C(n53), .Z(n51) );
  CNR2X2 U69 ( .A(A[48]), .B(n347), .Z(n68) );
  COND1X1 U68 ( .A(n71), .B(n68), .C(n69), .Z(n67) );
  COND1X1 U74 ( .A(n77), .B(n74), .C(n75), .Z(n73) );
  CANR1X1 U66 ( .A(n73), .B(n66), .C(n67), .Z(n65) );
  CNR2X2 U86 ( .A(A[44]), .B(n343), .Z(n85) );
  COND1X1 U85 ( .A(n88), .B(n85), .C(n86), .Z(n84) );
  CANR1X1 U83 ( .A(n90), .B(n83), .C(n84), .Z(n82) );
  CANR1X1 U111 ( .A(n2755), .B(net14039), .C(n2723), .Z(n110) );
  COND1X1 U99 ( .A(n99), .B(n110), .C(n100), .Z(n98) );
  CANR1X1 U123 ( .A(n2764), .B(n2712), .C(n2722), .Z(n122) );
  CANR1X1 U133 ( .A(n2746), .B(n2716), .C(n2748), .Z(n132) );
  CANR1X1 U97 ( .A(n120), .B(n97), .C(n98), .Z(n96) );
  CANR1X1 U148 ( .A(n2725), .B(n2715), .C(n2761), .Z(n147) );
  CANR1X1 U158 ( .A(n2757), .B(n158), .C(n2713), .Z(n157) );
  CANR1X1 U170 ( .A(n2762), .B(n170), .C(n2721), .Z(n169) );
  CNR2X2 U145 ( .A(n146), .B(n156), .Z(n144) );
  CANR1X1 U193 ( .A(n2763), .B(n2753), .C(n2720), .Z(n192) );
  CANR1X1 U235 ( .A(n2760), .B(n2750), .C(n236), .Z(n234) );
  CANR1X1 U245 ( .A(n2756), .B(n2749), .C(n2719), .Z(n244) );
  CANR1X1 U256 ( .A(n2759), .B(n2752), .C(n2718), .Z(n255) );
  CANR1X1 U274 ( .A(n2758), .B(n2751), .C(n2717), .Z(n273) );
  CANR1X1 U231 ( .A(n253), .B(n231), .C(n232), .Z(n230) );
  CANR1X1 U79 ( .A(n79), .B(n141), .C(n80), .Z(n78) );
  CND2X2 U51 ( .A(n58), .B(n52), .Z(n50) );
  CANR1X1 U7 ( .A(n2742), .B(n2711), .C(n2727), .Z(n6) );
  COND1X1 U3 ( .A(n3), .B(n6), .C(n4), .Z(n2) );
  COND1X1 U16 ( .A(n16), .B(n78), .C(n17), .Z(n15) );
  COND1X1 U44 ( .A(n47), .B(n44), .C(n45), .Z(n43) );
  CNR2X2 U31 ( .A(A[58]), .B(n357), .Z(n30) );
  CANR1X1 U18 ( .A(n18), .B(n49), .C(n19), .Z(n17) );
  COND1X1 U20 ( .A(n20), .B(n35), .C(n21), .Z(n19) );
  COR2X1 U1562 ( .A(A[62]), .B(n361), .Z(n2711) );
  CNR2X2 U1563 ( .A(n2743), .B(n2744), .Z(net19772) );
  CNR2IX1 U1564 ( .B(B[55]), .A(A[55]), .Z(n2744) );
  CND2X1 U1565 ( .A(n2732), .B(n28), .Z(n20) );
  CND2IX1 U1566 ( .B(n107), .A(net14042), .Z(n99) );
  COR2X1 U1567 ( .A(A[36]), .B(n335), .Z(n2712) );
  CAN2X1 U1568 ( .A(A[30]), .B(n329), .Z(n2713) );
  COR2X1 U1569 ( .A(A[26]), .B(n325), .Z(n2714) );
  COR2X1 U1570 ( .A(A[38]), .B(n337), .Z(net14039) );
  CNR2X1 U1571 ( .A(A[28]), .B(n327), .Z(n172) );
  COND1XL U1572 ( .A(n254), .B(n264), .C(n255), .Z(n253) );
  CND2IXL U1573 ( .B(n129), .A(n2712), .Z(n121) );
  CNR2X1 U1574 ( .A(A[63]), .B(n362), .Z(n3) );
  COND1XL U1575 ( .A(n214), .B(n211), .C(n212), .Z(n210) );
  COND1XL U1576 ( .A(n216), .B(n230), .C(n217), .Z(n215) );
  CANR1XL U1577 ( .A(n225), .B(n218), .C(n219), .Z(n217) );
  CNR2X1 U1578 ( .A(n178), .B(n168), .Z(n166) );
  CNR2X1 U1579 ( .A(A[49]), .B(n348), .Z(n62) );
  COND1XL U1580 ( .A(n94), .B(n91), .C(n92), .Z(n90) );
  CNR2XL U1581 ( .A(n131), .B(n121), .Z(n119) );
  COR2X1 U1582 ( .A(A[32]), .B(n331), .Z(n2715) );
  COR2X1 U1583 ( .A(A[34]), .B(n333), .Z(n2716) );
  CAN2X1 U1584 ( .A(A[6]), .B(n305), .Z(n2717) );
  CAN2X1 U1585 ( .A(A[10]), .B(n309), .Z(n2718) );
  CAN2X1 U1586 ( .A(A[12]), .B(n311), .Z(n2719) );
  CAN2XL U1587 ( .A(A[24]), .B(n323), .Z(n2720) );
  CAN2X1 U1588 ( .A(A[28]), .B(n327), .Z(n2721) );
  CAN2X1 U1589 ( .A(A[36]), .B(n335), .Z(n2722) );
  CAN2XL U1590 ( .A(A[38]), .B(n337), .Z(n2723) );
  CAN2X1 U1591 ( .A(A[39]), .B(n338), .Z(n2724) );
  CAN2XL U1592 ( .A(A[31]), .B(n330), .Z(n2725) );
  COR2XL U1593 ( .A(A[13]), .B(n312), .Z(n2726) );
  CAN2X1 U1594 ( .A(A[62]), .B(n361), .Z(n2727) );
  COR2XL U1595 ( .A(A[61]), .B(n360), .Z(n2728) );
  COR2XL U1596 ( .A(A[25]), .B(n324), .Z(n2729) );
  COR2XL U1597 ( .A(A[11]), .B(n310), .Z(n2730) );
  COR2XL U1598 ( .A(A[33]), .B(n332), .Z(n2731) );
  CNR2XL U1599 ( .A(n26), .B(net23082), .Z(n2732) );
  CANR1XL U1600 ( .A(n2739), .B(n2740), .C(n2741), .Z(n2736) );
  CNR2IX2 U1601 ( .B(B[60]), .A(A[60]), .Z(n2734) );
  CANR1X1 U1602 ( .A(n2733), .B(n27), .C(n2734), .Z(n23) );
  CNR2IX1 U1603 ( .B(B[60]), .A(A[60]), .Z(net23082) );
  CIVX2 U1604 ( .A(B[60]), .Z(n2735) );
  CND2X1 U1605 ( .A(A[60]), .B(n2735), .Z(n2733) );
  CANR1X2 U1606 ( .A(net14590), .B(n29), .C(n23), .Z(n21) );
  CND2X1 U1607 ( .A(A[59]), .B(n358), .Z(n27) );
  CIVX2 U1608 ( .A(B[59]), .Z(n358) );
  CNR2X1 U1609 ( .A(A[59]), .B(n358), .Z(n26) );
  COND1X1 U1610 ( .A(n33), .B(n30), .C(n31), .Z(n29) );
  CND2X1 U1611 ( .A(A[58]), .B(n357), .Z(n31) );
  CIVX2 U1612 ( .A(B[58]), .Z(n357) );
  CND2X2 U1613 ( .A(A[57]), .B(n356), .Z(n33) );
  CIVX2 U1614 ( .A(B[57]), .Z(n356) );
  CNR2X2 U1615 ( .A(A[57]), .B(n356), .Z(n32) );
  CANR1X1 U1616 ( .A(net19772), .B(n43), .C(n2736), .Z(n35) );
  CNR2IX1 U1617 ( .B(B[56]), .A(A[56]), .Z(n2741) );
  CND2XL U1618 ( .A(A[55]), .B(n2738), .Z(n2740) );
  CIVX2 U1619 ( .A(B[55]), .Z(n2738) );
  CND2XL U1620 ( .A(A[56]), .B(n2737), .Z(n2739) );
  CIVX2 U1621 ( .A(B[56]), .Z(n2737) );
  CND2X1 U1622 ( .A(A[54]), .B(n353), .Z(n45) );
  CIVX2 U1623 ( .A(B[54]), .Z(n353) );
  CNR2X2 U1624 ( .A(A[54]), .B(n353), .Z(n44) );
  CND2X1 U1625 ( .A(A[53]), .B(n352), .Z(n47) );
  CIVX2 U1626 ( .A(B[53]), .Z(n352) );
  CNR2X1 U1627 ( .A(n26), .B(net23082), .Z(net14590) );
  CNR2X1 U1628 ( .A(n30), .B(n32), .Z(n28) );
  CANR1X2 U1629 ( .A(n1), .B(n15), .C(n2), .Z(GE_LT_GT_LE) );
  CND2XL U1630 ( .A(A[63]), .B(n362), .Z(n4) );
  CIVX2 U1631 ( .A(B[63]), .Z(n362) );
  CIVX2 U1632 ( .A(B[62]), .Z(n361) );
  CND2X1 U1633 ( .A(n2728), .B(n2711), .Z(n5) );
  CAN2X1 U1634 ( .A(A[61]), .B(n360), .Z(n2742) );
  CIVX2 U1635 ( .A(B[61]), .Z(n360) );
  CNR2IX2 U1636 ( .B(n2766), .A(n50), .Z(n48) );
  CAN2X1 U1637 ( .A(n72), .B(n66), .Z(n2766) );
  CNR2XL U1638 ( .A(n46), .B(n44), .Z(n42) );
  CNR2IX1 U1639 ( .B(B[56]), .A(A[56]), .Z(n2743) );
  CNR2X1 U1640 ( .A(A[53]), .B(n352), .Z(n46) );
  CND2X1 U1641 ( .A(n42), .B(net19772), .Z(n34) );
  CNR2X1 U1642 ( .A(n5), .B(n3), .Z(n1) );
  CND2X1 U1643 ( .A(n48), .B(n18), .Z(n16) );
  CNR2X1 U1644 ( .A(n20), .B(n34), .Z(n18) );
  CNR2X1 U1645 ( .A(n76), .B(n74), .Z(n72) );
  CNR2XL U1646 ( .A(A[45]), .B(n344), .Z(n76) );
  CIVX2 U1647 ( .A(B[45]), .Z(n344) );
  CNR2X1 U1648 ( .A(A[46]), .B(n345), .Z(n74) );
  CNR2X2 U1649 ( .A(n70), .B(n68), .Z(n66) );
  CNR2XL U1650 ( .A(n81), .B(n95), .Z(n79) );
  CND2XL U1651 ( .A(n83), .B(n89), .Z(n81) );
  CND2XL U1652 ( .A(n119), .B(n97), .Z(n95) );
  CND2XL U1653 ( .A(n2731), .B(n2716), .Z(n131) );
  CIVX2 U1654 ( .A(B[33]), .Z(n332) );
  CNR2X1 U1655 ( .A(n109), .B(n99), .Z(n97) );
  COND1XL U1656 ( .A(n188), .B(n142), .C(n143), .Z(n141) );
  CANR1XL U1657 ( .A(n189), .B(n215), .C(n190), .Z(n188) );
  CNR2X1 U1658 ( .A(n201), .B(n191), .Z(n189) );
  CND2XL U1659 ( .A(n209), .B(n203), .Z(n201) );
  CNR2XL U1660 ( .A(n213), .B(n211), .Z(n209) );
  CNR2XL U1661 ( .A(A[19]), .B(n318), .Z(n213) );
  CIVX2 U1662 ( .A(B[19]), .Z(n318) );
  CNR2X1 U1663 ( .A(A[20]), .B(n319), .Z(n211) );
  CNR2XL U1664 ( .A(n207), .B(n205), .Z(n203) );
  CND2IX1 U1665 ( .B(n199), .A(n2753), .Z(n191) );
  CND2XL U1666 ( .A(n218), .B(n224), .Z(n216) );
  CNR2XL U1667 ( .A(n222), .B(n220), .Z(n218) );
  CNR2XL U1668 ( .A(n226), .B(n228), .Z(n224) );
  CNR2X1 U1669 ( .A(A[16]), .B(n315), .Z(n226) );
  CNR2XL U1670 ( .A(A[15]), .B(n314), .Z(n228) );
  CIVX2 U1671 ( .A(B[15]), .Z(n314) );
  CND2IXL U1672 ( .B(n262), .A(n2752), .Z(n254) );
  CNR2XL U1673 ( .A(A[9]), .B(n308), .Z(n262) );
  CIVX2 U1674 ( .A(B[9]), .Z(n308) );
  COR2X1 U1675 ( .A(A[10]), .B(n309), .Z(n2752) );
  CANR1XL U1676 ( .A(n271), .B(n265), .C(n266), .Z(n264) );
  COND1XL U1677 ( .A(n282), .B(n272), .C(n273), .Z(n271) );
  COAN1XL U1678 ( .A(n2765), .B(n285), .C(n286), .Z(n282) );
  COAN1X1 U1679 ( .A(n288), .B(n290), .C(n289), .Z(n2765) );
  CNR2X1 U1680 ( .A(A[3]), .B(n302), .Z(n288) );
  CIVX2 U1681 ( .A(B[3]), .Z(n302) );
  COAN1X1 U1682 ( .A(n293), .B(n2754), .C(n294), .Z(n290) );
  CNR2XL U1683 ( .A(A[2]), .B(n301), .Z(n293) );
  CIVX1 U1684 ( .A(B[2]), .Z(n301) );
  COAN1X1 U1685 ( .A(n298), .B(n296), .C(n297), .Z(n2754) );
  CND2X1 U1686 ( .A(A[0]), .B(n299), .Z(n298) );
  CIVX2 U1687 ( .A(B[0]), .Z(n299) );
  CNR2X1 U1688 ( .A(A[1]), .B(n300), .Z(n296) );
  CIVX1 U1689 ( .A(B[1]), .Z(n300) );
  CND2XL U1690 ( .A(A[1]), .B(n300), .Z(n297) );
  CND2XL U1691 ( .A(A[2]), .B(n301), .Z(n294) );
  CND2XL U1692 ( .A(A[3]), .B(n302), .Z(n289) );
  CNR2XL U1693 ( .A(A[4]), .B(n303), .Z(n285) );
  CIVX2 U1694 ( .A(B[4]), .Z(n303) );
  CND2XL U1695 ( .A(A[4]), .B(n303), .Z(n286) );
  CND2IXL U1696 ( .B(n280), .A(n2751), .Z(n272) );
  CNR2XL U1697 ( .A(A[5]), .B(n304), .Z(n280) );
  CIVX2 U1698 ( .A(B[5]), .Z(n304) );
  COR2X1 U1699 ( .A(A[6]), .B(n305), .Z(n2751) );
  CAN2X1 U1700 ( .A(A[5]), .B(n304), .Z(n2758) );
  CIVX2 U1701 ( .A(B[6]), .Z(n305) );
  CNR2X1 U1702 ( .A(n269), .B(n267), .Z(n265) );
  CNR2X1 U1703 ( .A(A[7]), .B(n306), .Z(n269) );
  CIVX2 U1704 ( .A(B[7]), .Z(n306) );
  CNR2XL U1705 ( .A(A[8]), .B(n307), .Z(n267) );
  COND1XL U1706 ( .A(n270), .B(n267), .C(n268), .Z(n266) );
  CND2XL U1707 ( .A(A[7]), .B(n306), .Z(n270) );
  CND2XL U1708 ( .A(A[8]), .B(n307), .Z(n268) );
  CIVX2 U1709 ( .A(B[8]), .Z(n307) );
  CAN2X1 U1710 ( .A(A[9]), .B(n308), .Z(n2759) );
  CIVX2 U1711 ( .A(B[10]), .Z(n309) );
  CNR2XL U1712 ( .A(n233), .B(n243), .Z(n231) );
  CND2X1 U1713 ( .A(n2750), .B(n2726), .Z(n233) );
  CND2XL U1714 ( .A(n2749), .B(n2730), .Z(n243) );
  COR2X1 U1715 ( .A(A[12]), .B(n311), .Z(n2749) );
  CIVX2 U1716 ( .A(B[11]), .Z(n310) );
  COND1X1 U1717 ( .A(n244), .B(n233), .C(n234), .Z(n232) );
  CAN2X1 U1718 ( .A(A[11]), .B(n310), .Z(n2756) );
  CIVX2 U1719 ( .A(B[12]), .Z(n311) );
  CAN2XL U1720 ( .A(A[13]), .B(n312), .Z(n2760) );
  CIVX2 U1721 ( .A(B[13]), .Z(n312) );
  COR2X1 U1722 ( .A(A[14]), .B(n313), .Z(n2750) );
  CIVXL U1723 ( .A(n238), .Z(n236) );
  CND2XL U1724 ( .A(A[14]), .B(n313), .Z(n238) );
  CIVX2 U1725 ( .A(B[14]), .Z(n313) );
  COND1XL U1726 ( .A(n229), .B(n226), .C(n227), .Z(n225) );
  CND2XL U1727 ( .A(A[15]), .B(n314), .Z(n229) );
  CND2XL U1728 ( .A(A[16]), .B(n315), .Z(n227) );
  CIVX2 U1729 ( .A(B[16]), .Z(n315) );
  COND1XL U1730 ( .A(n223), .B(n220), .C(n221), .Z(n219) );
  CND2XL U1731 ( .A(A[17]), .B(n316), .Z(n223) );
  CIVX2 U1732 ( .A(B[17]), .Z(n316) );
  CNR2X1 U1733 ( .A(A[18]), .B(n317), .Z(n220) );
  CND2XL U1734 ( .A(A[18]), .B(n317), .Z(n221) );
  CIVX2 U1735 ( .A(B[18]), .Z(n317) );
  COND1XL U1736 ( .A(n191), .B(n202), .C(n192), .Z(n190) );
  CANR1XL U1737 ( .A(n210), .B(n203), .C(n204), .Z(n202) );
  CND2XL U1738 ( .A(A[19]), .B(n318), .Z(n214) );
  CND2XL U1739 ( .A(A[20]), .B(n319), .Z(n212) );
  CIVX2 U1740 ( .A(B[20]), .Z(n319) );
  COND1XL U1741 ( .A(n208), .B(n205), .C(n206), .Z(n204) );
  CND2X1 U1742 ( .A(A[21]), .B(n320), .Z(n208) );
  CIVX2 U1743 ( .A(B[21]), .Z(n320) );
  CNR2X1 U1744 ( .A(A[22]), .B(n321), .Z(n205) );
  CND2XL U1745 ( .A(A[22]), .B(n321), .Z(n206) );
  CIVX2 U1746 ( .A(B[22]), .Z(n321) );
  CAN2X1 U1747 ( .A(A[23]), .B(n322), .Z(n2763) );
  CIVX2 U1748 ( .A(B[23]), .Z(n322) );
  COR2X1 U1749 ( .A(A[24]), .B(n323), .Z(n2753) );
  CIVX2 U1750 ( .A(B[24]), .Z(n323) );
  CND2X1 U1751 ( .A(n144), .B(n166), .Z(n142) );
  CND2X1 U1752 ( .A(n2729), .B(n2714), .Z(n178) );
  CIVX2 U1753 ( .A(B[25]), .Z(n324) );
  CND2IX1 U1754 ( .B(n176), .A(n170), .Z(n168) );
  CANR1XL U1755 ( .A(n167), .B(n144), .C(n145), .Z(n143) );
  COND1XL U1756 ( .A(n168), .B(n179), .C(n169), .Z(n167) );
  CANR1XL U1757 ( .A(n2745), .B(n2714), .C(n2747), .Z(n179) );
  CAN2XL U1758 ( .A(A[25]), .B(n324), .Z(n2745) );
  CAN2X1 U1759 ( .A(A[26]), .B(n325), .Z(n2747) );
  CIVX2 U1760 ( .A(B[26]), .Z(n325) );
  CAN2XL U1761 ( .A(A[27]), .B(n326), .Z(n2762) );
  CIVX2 U1762 ( .A(B[27]), .Z(n326) );
  CIVX2 U1763 ( .A(n172), .Z(n170) );
  CIVX2 U1764 ( .A(B[28]), .Z(n327) );
  COND1XL U1765 ( .A(n157), .B(n146), .C(n147), .Z(n145) );
  CAN2X1 U1766 ( .A(A[29]), .B(n328), .Z(n2757) );
  CIVX2 U1767 ( .A(B[29]), .Z(n328) );
  CIVX2 U1768 ( .A(n160), .Z(n158) );
  CIVX2 U1769 ( .A(B[30]), .Z(n329) );
  CND2IX1 U1770 ( .B(n154), .A(n2715), .Z(n146) );
  CIVX2 U1771 ( .A(B[31]), .Z(n330) );
  CAN2X1 U1772 ( .A(A[32]), .B(n331), .Z(n2761) );
  CIVX2 U1773 ( .A(B[32]), .Z(n331) );
  COND1X1 U1774 ( .A(n81), .B(n96), .C(n82), .Z(n80) );
  COND1XL U1775 ( .A(n121), .B(n132), .C(n122), .Z(n120) );
  CAN2X1 U1776 ( .A(A[33]), .B(n332), .Z(n2746) );
  CAN2X1 U1777 ( .A(A[34]), .B(n333), .Z(n2748) );
  CIVX2 U1778 ( .A(B[34]), .Z(n333) );
  CAN2XL U1779 ( .A(A[35]), .B(n334), .Z(n2764) );
  CIVX2 U1780 ( .A(B[35]), .Z(n334) );
  CIVX2 U1781 ( .A(B[36]), .Z(n335) );
  CNR2X1 U1782 ( .A(A[39]), .B(n338), .Z(n107) );
  CND2IX1 U1783 ( .B(A[40]), .A(B[40]), .Z(net14042) );
  CAN2X1 U1784 ( .A(A[37]), .B(n336), .Z(n2755) );
  CIVX2 U1785 ( .A(B[37]), .Z(n336) );
  CIVX2 U1786 ( .A(B[38]), .Z(n337) );
  CANR1X2 U1787 ( .A(n2724), .B(net14042), .C(n2767), .Z(n100) );
  CIVX2 U1788 ( .A(B[39]), .Z(n338) );
  CAN2X1 U1789 ( .A(A[40]), .B(n339), .Z(n2767) );
  CIVX2 U1790 ( .A(B[40]), .Z(n339) );
  CND2X1 U1791 ( .A(A[41]), .B(n340), .Z(n94) );
  CIVX2 U1792 ( .A(B[41]), .Z(n340) );
  CNR2X1 U1793 ( .A(A[42]), .B(n341), .Z(n91) );
  CND2XL U1794 ( .A(A[42]), .B(n341), .Z(n92) );
  CIVX2 U1795 ( .A(B[42]), .Z(n341) );
  CNR2X1 U1796 ( .A(n87), .B(n85), .Z(n83) );
  CND2X1 U1797 ( .A(A[43]), .B(n342), .Z(n88) );
  CIVX2 U1798 ( .A(B[43]), .Z(n342) );
  CND2X1 U1799 ( .A(A[44]), .B(n343), .Z(n86) );
  CIVX2 U1800 ( .A(B[44]), .Z(n343) );
  COND1XL U1801 ( .A(n50), .B(n65), .C(n51), .Z(n49) );
  CND2XL U1802 ( .A(A[45]), .B(n344), .Z(n77) );
  CND2XL U1803 ( .A(A[46]), .B(n345), .Z(n75) );
  CIVX2 U1804 ( .A(B[46]), .Z(n345) );
  CND2X1 U1805 ( .A(A[47]), .B(n346), .Z(n71) );
  CIVX2 U1806 ( .A(B[47]), .Z(n346) );
  CND2XL U1807 ( .A(A[48]), .B(n347), .Z(n69) );
  CIVX2 U1808 ( .A(B[48]), .Z(n347) );
  CND2X1 U1809 ( .A(A[49]), .B(n348), .Z(n63) );
  CIVX2 U1810 ( .A(B[49]), .Z(n348) );
  CND2XL U1811 ( .A(A[50]), .B(n349), .Z(n61) );
  CIVX2 U1812 ( .A(B[50]), .Z(n349) );
  CND2X1 U1813 ( .A(A[51]), .B(n350), .Z(n57) );
  CIVX2 U1814 ( .A(B[51]), .Z(n350) );
  CNR2X2 U1815 ( .A(A[52]), .B(n351), .Z(n54) );
  CND2XL U1816 ( .A(A[52]), .B(n351), .Z(n55) );
  CIVX2 U1817 ( .A(B[52]), .Z(n351) );
  CND2IX1 U1818 ( .B(n164), .A(n158), .Z(n156) );
  CNR2XL U1819 ( .A(A[17]), .B(n316), .Z(n222) );
  CNR2XL U1820 ( .A(A[21]), .B(n320), .Z(n207) );
  CND2IXL U1821 ( .B(n117), .A(net14039), .Z(n109) );
  CNR2XL U1822 ( .A(A[29]), .B(n328), .Z(n164) );
  CNR2XL U1823 ( .A(n91), .B(n93), .Z(n89) );
  CNR2XL U1824 ( .A(A[41]), .B(n340), .Z(n93) );
  CNR2XL U1825 ( .A(A[37]), .B(n336), .Z(n117) );
  CNR2X1 U1826 ( .A(A[43]), .B(n342), .Z(n87) );
  CNR2X1 U1827 ( .A(A[35]), .B(n334), .Z(n129) );
  CNR2X1 U1828 ( .A(A[27]), .B(n326), .Z(n176) );
  CNR2X1 U1829 ( .A(A[23]), .B(n322), .Z(n199) );
  CNR2X1 U1830 ( .A(A[31]), .B(n330), .Z(n154) );
endmodule


module sqrt64 ( clk, rdy, reset, x, acc );
  input [63:0] x;
  output [31:0] acc;
  input clk, reset;
  output rdy;
  wire   N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91,
         N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126,
         N128, N130, N131, N132, N133, N134, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n98, N9, N8, N7, N63, N62, N61, N60, N6, N59, N58, N57,
         N56, N55, N54, N53, N52, N51, N50, N5, N49, N48, N47, N46, N45, N44,
         N43, N42, N41, N40, N4, N39, N38, N37, N36, N35, N34, N33, N32, N31,
         N30, N3, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N2, N19,
         N18, N17, N16, N15, N14, N13, N12, N11, N10, N1, N0, net3640,
         net10635, net10636, net10639, net10644, net10816, net11095, net11163,
         net11166, net13656, net13668, net13671, net13702, net13725, net13724,
         net14219, net14218, net14242, net14241, net14250, net14249, net14327,
         net14518, net14502, net14488, net14486, net14483, net14606, net14615,
         net14652, net14651, net14734, net17171, net17179, net23250, net23249,
         net26377, net26430, net26435, net26437, net26606, net26601, net26813,
         net26812, net31721, net31723, net31747, net13672, net26633, net26596,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601;
  wire   [4:0] bitl;
  wire   [63:0] bit2;
  wire   [63:0] acc2;
  wire   [63:0] guess2;

  CFD4QX4 \bitl_reg[0]  ( .D(n118), .CP(clk), .SD(n230), .Q(bitl[0]) );
  CFD4QX4 \bitl_reg[1]  ( .D(N130), .CP(clk), .SD(n230), .Q(net17179) );
  CFD4QX4 \bitl_reg[2]  ( .D(N131), .CP(clk), .SD(n230), .Q(bitl[2]) );
  CFD4QX4 \bitl_reg[3]  ( .D(N132), .CP(clk), .SD(n230), .Q(bitl[3]) );
  CFD4QX4 \bitl_reg[4]  ( .D(N133), .CP(clk), .SD(n230), .Q(bitl[4]) );
  sqrt64_DW01_add_5 add_1_root_add_0_root_add_39_2 ( .A({n161, n162, n145, 
        n144, acc2[59:56], n172, n164, n175, n166, n174, n171, n193, n169, 
        n179, acc2[46], n178, n170, net14488, n190, net14502, acc2[40], n152, 
        n181, n151, n185, n187, n184, n142, n158, n180, n155, n189, net14518, 
        n149, n183, net14483, n156, n143, n157, n146, n192, n150, n159, n154, 
        n188, n176, n163, n153, n182, n148, n186, n194, n165, net14486, n167, 
        n147, n168, n173, n191, n160, n177}), .B({1'b0, n200, 1'b0, bit2[60], 
        1'b0, bit2[58], 1'b0, bit2[56], 1'b0, bit2[54], 1'b0, bit2[52], 1'b0, 
        bit2[50], 1'b0, bit2[48], 1'b0, bit2[46], 1'b0, bit2[44], 1'b0, 
        bit2[42], 1'b0, bit2[40], 1'b0, bit2[38], 1'b0, bit2[36], 1'b0, 
        bit2[34], 1'b0, bit2[32], 1'b0, n113, 1'b0, bit2[28], 1'b0, bit2[26], 
        1'b0, bit2[24], 1'b0, bit2[22], 1'b0, bit2[20], 1'b0, bit2[18], 1'b0, 
        bit2[16], 1'b0, bit2[14], 1'b0, bit2[12], 1'b0, bit2[10], 1'b0, 
        bit2[8], 1'b0, bit2[6], 1'b0, bit2[4], 1'b0, bit2[2], 1'b0, bit2[0]}), 
        .CI(1'b0), .SUM({N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, 
        N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  sqrt64_DW01_add_10 add_0_root_add_0_root_add_39_2 ( .A({N126, N125, N124, 
        N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, 
        N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, 
        N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, 
        N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, 
        N71, N70, N69, N68, N67, N66, N65, N64, 1'b0}), .B({N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, 
        N1, N0}), .CI(1'b0), .SUM(guess2) );
  sqrt64_DW_cmp_4 lte_55 ( .A(guess2), .B(x), .TC(1'b0), .GE_LT(1'b0), 
        .GE_GT_EQ(1'b0), .GE_LT_GT_LE(N128) );
  CFD2XL \acc2_reg[9]  ( .D(n43), .CP(clk), .CD(n225), .Q(n194) );
  CFD2XL \acc2_reg[49]  ( .D(n83), .CP(clk), .CD(n228), .Q(n193) );
  CFD2XL \acc2_reg[20]  ( .D(n54), .CP(clk), .CD(n226), .Q(n192) );
  CFD2XL \acc2_reg[2]  ( .D(n36), .CP(clk), .CD(n225), .Q(n191) );
  CFD2XL \acc2_reg[42]  ( .D(n76), .CP(clk), .CD(n228), .Q(n190) );
  CFD2XL \acc2_reg[29]  ( .D(n63), .CP(clk), .CD(n227), .Q(n189) );
  CFD2XL \acc2_reg[16]  ( .D(n50), .CP(clk), .CD(n226), .Q(n188) );
  CFD2XL \acc2_reg[35]  ( .D(n69), .CP(clk), .CD(n227), .Q(n187) );
  CFD2XL \acc2_reg[10]  ( .D(n44), .CP(clk), .CD(n225), .Q(n186) );
  CFD2XL \acc2_reg[36]  ( .D(n70), .CP(clk), .CD(n227), .Q(n185) );
  CFD2XL \acc2_reg[34]  ( .D(n68), .CP(clk), .CD(n227), .Q(n184) );
  CFD2XL \acc2_reg[26]  ( .D(n60), .CP(clk), .CD(n227), .Q(n183) );
  CFD2XL \acc2_reg[12]  ( .D(n46), .CP(clk), .CD(n226), .Q(n182) );
  CFD2XL \acc2_reg[38]  ( .D(n72), .CP(clk), .CD(n228), .Q(n181) );
  CFD2XL \acc2_reg[31]  ( .D(n65), .CP(clk), .CD(n227), .Q(n180) );
  CFD2XL \acc2_reg[47]  ( .D(n81), .CP(clk), .CD(n228), .Q(n179) );
  CFD2XL \acc2_reg[45]  ( .D(n79), .CP(clk), .CD(n228), .Q(n178) );
  CFD2XL \acc2_reg[0]  ( .D(n34), .CP(clk), .CD(n225), .Q(n177) );
  CFD2XL \acc2_reg[15]  ( .D(n49), .CP(clk), .CD(n226), .Q(n176) );
  CFD2XL \acc2_reg[53]  ( .D(n87), .CP(clk), .CD(n229), .Q(n175) );
  CFD2XL \acc2_reg[51]  ( .D(n85), .CP(clk), .CD(n229), .Q(n174) );
  CFD2XL \acc2_reg[3]  ( .D(n37), .CP(clk), .CD(n225), .Q(n173) );
  CFD2XL \acc2_reg[55]  ( .D(n89), .CP(clk), .CD(n229), .Q(n172) );
  CFD2XL \acc2_reg[50]  ( .D(n84), .CP(clk), .CD(n228), .Q(n171) );
  CFD2XL \acc2_reg[44]  ( .D(n78), .CP(clk), .CD(n228), .Q(n170) );
  CFD2XL \acc2_reg[48]  ( .D(n82), .CP(clk), .CD(n228), .Q(n169) );
  CFD2XL \acc2_reg[4]  ( .D(n38), .CP(clk), .CD(n225), .Q(n168) );
  CFD2XL \acc2_reg[6]  ( .D(n40), .CP(clk), .CD(n225), .Q(n167) );
  CFD2XL \acc2_reg[52]  ( .D(n86), .CP(clk), .CD(n229), .Q(n166) );
  CFD2XL \acc2_reg[8]  ( .D(n42), .CP(clk), .CD(n225), .Q(n165) );
  CFD2XL \acc2_reg[54]  ( .D(n88), .CP(clk), .CD(n229), .Q(n164) );
  CFD2XL \acc2_reg[14]  ( .D(n48), .CP(clk), .CD(n226), .Q(n163) );
  CFD2XL \acc2_reg[62]  ( .D(n96), .CP(clk), .CD(n229), .Q(n162) );
  CFD2XL \acc2_reg[63]  ( .D(n98), .CP(clk), .CD(n229), .Q(n161) );
  CFD2XL \acc2_reg[1]  ( .D(n35), .CP(clk), .CD(n225), .Q(n160) );
  CFD2XL \acc2_reg[18]  ( .D(n52), .CP(clk), .CD(n226), .Q(n159) );
  CFD2XL \acc2_reg[32]  ( .D(n66), .CP(clk), .CD(n227), .Q(n158) );
  CFD2XL \acc2_reg[22]  ( .D(n56), .CP(clk), .CD(n226), .Q(n157) );
  CFD2XL \acc2_reg[28]  ( .D(n62), .CP(clk), .CD(n227), .Q(net14518) );
  CFD2XL \acc2_reg[24]  ( .D(n58), .CP(clk), .CD(n226), .Q(n156) );
  CFD2XL \acc2_reg[30]  ( .D(n64), .CP(clk), .CD(n227), .Q(n155) );
  CFD2XL \acc2_reg[13]  ( .D(n47), .CP(clk), .CD(n226), .Q(n153) );
  CFD2XL \acc2_reg[39]  ( .D(n73), .CP(clk), .CD(n228), .Q(n152) );
  CFD2XL \acc2_reg[19]  ( .D(n53), .CP(clk), .CD(n226), .Q(n150) );
  CFD2XL \acc2_reg[27]  ( .D(n61), .CP(clk), .CD(n227), .Q(n149) );
  CFD2XL \acc2_reg[11]  ( .D(n45), .CP(clk), .CD(n225), .Q(n148) );
  CFD2XL \acc2_reg[5]  ( .D(n39), .CP(clk), .CD(n225), .Q(n147) );
  CFD2XL \acc2_reg[43]  ( .D(n77), .CP(clk), .CD(n228), .Q(net14488) );
  CFD2XL \acc2_reg[21]  ( .D(n55), .CP(clk), .CD(n226), .Q(n146) );
  CFD2XL \acc2_reg[61]  ( .D(n95), .CP(clk), .CD(n229), .Q(n145) );
  CFD2XL \acc2_reg[60]  ( .D(n94), .CP(clk), .CD(n229), .Q(n144) );
  CFD2XL \acc2_reg[23]  ( .D(n57), .CP(clk), .CD(n226), .Q(n143) );
  CFD2XL \acc2_reg[33]  ( .D(n67), .CP(clk), .CD(n227), .Q(n142) );
  CFD2XL \acc2_reg[17]  ( .D(n51), .CP(clk), .CD(n226), .Q(n154) );
  CFD2XL \acc2_reg[37]  ( .D(n71), .CP(clk), .CD(n227), .Q(n151) );
  CFD2XL \acc2_reg[25]  ( .D(n59), .CP(clk), .CD(n227), .Q(net14483) );
  CFD2XL \acc2_reg[59]  ( .D(n93), .CP(clk), .CD(n229), .Q(acc2[59]), .QN(n578) );
  CFD2XL \acc2_reg[58]  ( .D(n92), .CP(clk), .CD(n229), .Q(acc2[58]), .QN(n580) );
  CFD2XL \acc2_reg[56]  ( .D(n90), .CP(clk), .CD(n229), .Q(acc2[56]), .QN(n583) );
  CFD2XL \acc2_reg[46]  ( .D(n80), .CP(clk), .CD(n228), .Q(acc2[46]), .QN(n585) );
  CFD2XL \acc2_reg[40]  ( .D(n74), .CP(clk), .CD(n228), .Q(acc2[40]), .QN(n587) );
  CFD2XL \acc2_reg[7]  ( .D(n41), .CP(clk), .CD(n225), .Q(net14486) );
  CFD2XL \bitl_reg[5]  ( .D(N134), .CP(clk), .CD(n601), .Q(rdy), .QN(n572) );
  CFD2XL \acc_reg[23]  ( .D(n10), .CP(clk), .CD(n601), .Q(acc[23]), .QN(n312)
         );
  CFD2XL \acc_reg[20]  ( .D(n13), .CP(clk), .CD(n601), .Q(acc[20]), .QN(n313)
         );
  CFD2XL \acc_reg[19]  ( .D(n14), .CP(clk), .CD(n601), .Q(acc[19]), .QN(n324)
         );
  CFD2XL \acc_reg[16]  ( .D(n17), .CP(clk), .CD(n601), .Q(acc[16]), .QN(n325)
         );
  CFD2XL \acc_reg[22]  ( .D(n11), .CP(clk), .CD(n601), .Q(acc[22]), .QN(n311)
         );
  CFD2XL \acc_reg[21]  ( .D(n12), .CP(clk), .CD(n601), .Q(acc[21]), .QN(n314)
         );
  CFD2XL \acc_reg[18]  ( .D(n15), .CP(clk), .CD(n601), .Q(acc[18]), .QN(n323)
         );
  CFD2XL \acc_reg[17]  ( .D(n16), .CP(clk), .CD(n601), .Q(acc[17]), .QN(n326)
         );
  CFD2XL \acc2_reg[57]  ( .D(n91), .CP(clk), .CD(n601), .Q(acc2[57]), .QN(n582) );
  CFD2XL \acc_reg[7]  ( .D(n26), .CP(clk), .CD(n601), .Q(acc[7]), .QN(n348) );
  CFD2XL \acc_reg[6]  ( .D(n27), .CP(clk), .CD(n601), .Q(acc[6]), .QN(n347) );
  CFD2XL \acc_reg[5]  ( .D(n28), .CP(clk), .CD(n601), .Q(acc[5]), .QN(n350) );
  CFD2XL \acc_reg[4]  ( .D(n29), .CP(clk), .CD(n601), .Q(acc[4]), .QN(n349) );
  CFD2XL \acc_reg[3]  ( .D(n30), .CP(clk), .CD(n601), .Q(acc[3]), .QN(n337) );
  CFD2XL \acc_reg[2]  ( .D(n31), .CP(clk), .CD(n601), .Q(acc[2]), .QN(n336) );
  CFD2XL \acc_reg[31]  ( .D(n2), .CP(clk), .CD(n601), .Q(acc[31]), .QN(n356)
         );
  CFD2XL \acc_reg[30]  ( .D(n3), .CP(clk), .CD(n601), .Q(acc[30]), .QN(n331)
         );
  CFD2XL \acc_reg[29]  ( .D(n4), .CP(clk), .CD(n601), .Q(acc[29]), .QN(n333)
         );
  CFD2XL \acc_reg[28]  ( .D(n5), .CP(clk), .CD(n601), .Q(acc[28]), .QN(n332)
         );
  CFD2XL \acc_reg[27]  ( .D(n6), .CP(clk), .CD(n601), .Q(acc[27]), .QN(n306)
         );
  CFD2XL \acc_reg[26]  ( .D(n7), .CP(clk), .CD(n601), .Q(acc[26]), .QN(n305)
         );
  CFD2XL \acc_reg[25]  ( .D(n8), .CP(clk), .CD(n601), .Q(acc[25]), .QN(n308)
         );
  CFD2XL \acc_reg[24]  ( .D(n9), .CP(clk), .CD(n601), .Q(acc[24]), .QN(n307)
         );
  CFD2XL \acc_reg[15]  ( .D(n18), .CP(clk), .CD(n601), .Q(acc[15]), .QN(n318)
         );
  CFD2XL \acc_reg[14]  ( .D(n19), .CP(clk), .CD(n601), .Q(acc[14]), .QN(n317)
         );
  CFD2XL \acc_reg[13]  ( .D(n20), .CP(clk), .CD(n601), .Q(acc[13]), .QN(n320)
         );
  CFD2XL \acc_reg[12]  ( .D(n21), .CP(clk), .CD(n601), .Q(acc[12]), .QN(n319)
         );
  CFD2XL \acc_reg[11]  ( .D(n22), .CP(clk), .CD(n601), .Q(acc[11]), .QN(n342)
         );
  CFD2XL \acc_reg[8]  ( .D(n25), .CP(clk), .CD(n601), .Q(acc[8]), .QN(n343) );
  CFD2XL \acc_reg[10]  ( .D(n23), .CP(clk), .CD(n601), .Q(acc[10]), .QN(n341)
         );
  CFD2XL \acc_reg[9]  ( .D(n24), .CP(clk), .CD(n601), .Q(acc[9]), .QN(n344) );
  CFD2X2 \acc_reg[1]  ( .D(n32), .CP(clk), .CD(n601), .Q(acc[1]), .QN(n338) );
  CFD2X1 \acc_reg[0]  ( .D(n33), .CP(clk), .CD(n601), .Q(acc[0]), .QN(n598) );
  CFD2X2 \acc2_reg[41]  ( .D(n75), .CP(clk), .CD(n228), .Q(net14502) );
  CIVX1 U102 ( .A(n591), .Z(n592) );
  CNR2X1 U103 ( .A(n591), .B(n137), .Z(bit2[16]) );
  CIVXL U104 ( .A(net14502), .Z(n126) );
  CND2X1 U105 ( .A(net31721), .B(n571), .Z(n600) );
  CNIVX1 U106 ( .A(n333), .Z(n100) );
  CNIVX1 U107 ( .A(n331), .Z(n101) );
  CAN2X1 U108 ( .A(n483), .B(n107), .Z(n102) );
  CIVX2 U109 ( .A(bitl[4]), .Z(net26435) );
  CIVXL U110 ( .A(n594), .Z(n103) );
  CAN2X2 U111 ( .A(n595), .B(net14651), .Z(bit2[12]) );
  CNIVX4 U112 ( .A(n198), .Z(n140) );
  CAN2X1 U113 ( .A(n196), .B(n564), .Z(N74) );
  CND2X2 U114 ( .A(net26633), .B(n125), .Z(net26596) );
  CIVX1 U115 ( .A(bitl[0]), .Z(net26606) );
  CANR2X1 U116 ( .A(net14241), .B(n336), .C(n338), .D(net26377), .Z(n254) );
  CANR2XL U117 ( .A(n109), .B(n336), .C(n596), .D(n338), .Z(n296) );
  CAN2X2 U118 ( .A(n210), .B(n596), .Z(n113) );
  CAN2X2 U119 ( .A(n593), .B(bitl[3]), .Z(n210) );
  CAN2X1 U120 ( .A(n210), .B(net13725), .Z(bit2[26]) );
  CDLY1XL U121 ( .A(guess2[50]), .Z(n104) );
  COND1X2 U122 ( .A(n550), .B(n224), .C(n518), .Z(N98) );
  CIVX1 U123 ( .A(n522), .Z(n558) );
  CAN2X2 U124 ( .A(n590), .B(net10636), .Z(bit2[34]) );
  CIVX1 U125 ( .A(n379), .Z(n469) );
  CIVXL U126 ( .A(n377), .Z(n470) );
  COND2XL U127 ( .A(n197), .B(n537), .C(n536), .D(n112), .Z(N89) );
  CAN2XL U128 ( .A(n102), .B(net10636), .Z(bit2[58]) );
  CANR2XL U129 ( .A(net14218), .B(n312), .C(net10636), .D(n311), .Z(n316) );
  CANR2XL U130 ( .A(net14242), .B(n313), .C(net10636), .D(n324), .Z(n290) );
  CANR2XL U131 ( .A(net14242), .B(n318), .C(net10636), .D(n317), .Z(n322) );
  CANR2XL U132 ( .A(net14242), .B(n333), .C(net10636), .D(n332), .Z(n262) );
  CANR2XL U133 ( .A(net14242), .B(n349), .C(net10636), .D(n337), .Z(n297) );
  CANR2XL U134 ( .A(net14242), .B(n337), .C(net10636), .D(n336), .Z(n340) );
  CANR2XL U135 ( .A(net14242), .B(n331), .C(net10636), .D(n333), .Z(n241) );
  CDLY1XL U136 ( .A(guess2[38]), .Z(n105) );
  CIVX2 U137 ( .A(n487), .Z(n593) );
  CIVXL U138 ( .A(net14606), .Z(n106) );
  CIVXL U139 ( .A(n106), .Z(n107) );
  CAN2X2 U140 ( .A(n209), .B(net14606), .Z(n211) );
  CIVX1 U141 ( .A(bitl[2]), .Z(net14249) );
  CNIVX1 U142 ( .A(net14652), .Z(n108) );
  CNIVX4 U143 ( .A(net14652), .Z(n109) );
  CNIVX4 U144 ( .A(net14652), .Z(n110) );
  CAN2X2 U145 ( .A(net17179), .B(net13672), .Z(net14652) );
  CNR2X2 U146 ( .A(bitl[4]), .B(bitl[2]), .Z(n125) );
  CIVX3 U147 ( .A(n294), .Z(n136) );
  CND2X2 U148 ( .A(net26435), .B(bitl[2]), .Z(n487) );
  CND3X1 U149 ( .A(net23249), .B(bitl[3]), .C(net10644), .Z(n591) );
  COND1XL U150 ( .A(n218), .B(n549), .C(n353), .Z(n563) );
  CIVX2 U151 ( .A(n489), .Z(n524) );
  CND2X1 U152 ( .A(net13671), .B(net13668), .Z(n137) );
  COND1XL U153 ( .A(n539), .B(n489), .C(n382), .Z(N120) );
  CIVX2 U154 ( .A(bitl[0]), .Z(net13672) );
  COND1XL U155 ( .A(n422), .B(n224), .C(n421), .Z(N117) );
  CIVX2 U156 ( .A(n396), .Z(n483) );
  COND1XL U157 ( .A(n205), .B(n224), .C(n492), .Z(N109) );
  COND1XL U158 ( .A(n203), .B(n224), .C(n495), .Z(N107) );
  COND1XL U159 ( .A(n460), .B(n224), .C(n459), .Z(N113) );
  CAN2X1 U160 ( .A(n565), .B(n196), .Z(N73) );
  CIVX12 U161 ( .A(net31747), .Z(net14327) );
  CND2XL U162 ( .A(net14327), .B(net11163), .Z(n130) );
  CND2XL U163 ( .A(net31721), .B(net11163), .Z(n129) );
  CND2XL U164 ( .A(net14327), .B(net11163), .Z(n128) );
  CIVDX1 U165 ( .A(n555), .Z0(n111), .Z1(n112) );
  CIVXL U166 ( .A(net26377), .Z(net13656) );
  CAN2X1 U167 ( .A(bitl[2]), .B(n114), .Z(n209) );
  CMXI2XL U168 ( .A0(n115), .A1(n581), .S(net31721), .Z(n91) );
  CMXI2XL U169 ( .A0(n119), .A1(n584), .S(net31723), .Z(n80) );
  CMXI2XL U170 ( .A0(n122), .A1(n579), .S(net31723), .Z(n92) );
  CMXI2XL U171 ( .A0(n117), .A1(n577), .S(net31723), .Z(n93) );
  CMXI2XL U172 ( .A0(n120), .A1(n586), .S(net31721), .Z(n74) );
  CMXI2XL U173 ( .A0(n126), .A1(n127), .S(net31721), .Z(n75) );
  CMXI2XL U174 ( .A0(n123), .A1(n223), .S(net31723), .Z(n90) );
  CAOR1XL U175 ( .A(n398), .B(n217), .C(n397), .Z(n503) );
  CANR2XL U176 ( .A(n483), .B(n386), .C(n217), .D(n385), .Z(n387) );
  CANR2XL U177 ( .A(n483), .B(n417), .C(n217), .D(n416), .Z(n418) );
  CANR2XL U178 ( .A(n483), .B(n416), .C(n217), .D(n414), .Z(n365) );
  CANR2XL U179 ( .A(n477), .B(n483), .C(n484), .D(n217), .Z(n329) );
  CANR2XL U180 ( .A(n440), .B(n483), .C(n441), .D(n217), .Z(n360) );
  CANR2XL U181 ( .A(n484), .B(n483), .C(n482), .D(n217), .Z(n485) );
  CANR2XL U182 ( .A(n483), .B(n404), .C(n217), .D(n403), .Z(n405) );
  CANR2XL U183 ( .A(n468), .B(n483), .C(n463), .D(n217), .Z(n291) );
  CANR2XL U184 ( .A(n441), .B(n483), .C(n438), .D(n217), .Z(n248) );
  CANR2XL U185 ( .A(n469), .B(n483), .C(n467), .D(n217), .Z(n425) );
  CANR2XL U186 ( .A(n454), .B(n483), .C(n450), .D(n217), .Z(n269) );
  CANR2XL U187 ( .A(n483), .B(n374), .C(n217), .D(n373), .Z(n375) );
  CANR2XL U188 ( .A(n450), .B(n483), .C(n449), .D(n217), .Z(n451) );
  CIVX2 U189 ( .A(bitl[3]), .Z(n114) );
  CIVX2 U190 ( .A(bitl[3]), .Z(net10639) );
  CNIVX1 U191 ( .A(net10639), .Z(net26430) );
  CNIVX1 U192 ( .A(n582), .Z(n115) );
  CNIVX1 U193 ( .A(n356), .Z(n116) );
  CNIVX1 U194 ( .A(n578), .Z(n117) );
  CNIVX1 U195 ( .A(net13656), .Z(n118) );
  CNIVX1 U196 ( .A(n585), .Z(n119) );
  CNIVX1 U197 ( .A(n587), .Z(n120) );
  CNIVX1 U198 ( .A(net23249), .Z(n121) );
  CNIVX1 U199 ( .A(n580), .Z(n122) );
  CNIVX1 U200 ( .A(n583), .Z(n123) );
  CND2X1 U201 ( .A(n131), .B(n596), .Z(n124) );
  CIVX2 U202 ( .A(n124), .Z(bit2[14]) );
  CNR2IX1 U203 ( .B(bitl[0]), .A(net26596), .Z(bit2[2]) );
  CMX2XL U204 ( .A0(net14488), .A1(guess2[43]), .S(net14327), .Z(n77) );
  CIVX4 U205 ( .A(N128), .Z(net31747) );
  CMX2XL U206 ( .A0(net14518), .A1(guess2[28]), .S(net14327), .Z(n62) );
  CMX2XL U207 ( .A0(net14483), .A1(guess2[25]), .S(net14327), .Z(n59) );
  CMX2XL U208 ( .A0(net14486), .A1(guess2[7]), .S(net14327), .Z(n41) );
  CNR2IX1 U209 ( .B(net26606), .A(net26596), .Z(bit2[0]) );
  CNR2X2 U210 ( .A(bitl[3]), .B(net17179), .Z(net26633) );
  CIVXL U211 ( .A(bitl[4]), .Z(net26437) );
  CIVX1 U212 ( .A(bitl[4]), .Z(net10644) );
  CAN2XL U213 ( .A(net17179), .B(net13672), .Z(net14651) );
  CIVX2 U214 ( .A(guess2[41]), .Z(n127) );
  CIVX1 U215 ( .A(net31747), .Z(net31721) );
  CIVXL U216 ( .A(net31747), .Z(net31723) );
  CIVXL U217 ( .A(n110), .Z(net26812) );
  CIVX2 U218 ( .A(net26812), .Z(net26813) );
  CIVX2 U219 ( .A(n294), .Z(n596) );
  CIVDX2 U220 ( .A(n557), .Z0(n196), .Z1(n197) );
  COND2XL U221 ( .A(n528), .B(n489), .C(rdy), .D(n488), .Z(n490) );
  COND2XL U222 ( .A(n526), .B(n489), .C(n208), .D(n112), .Z(N111) );
  COND2XL U223 ( .A(n547), .B(n489), .C(n546), .D(n427), .Z(n428) );
  CIVX2 U224 ( .A(bitl[2]), .Z(net23249) );
  CIVXL U225 ( .A(n594), .Z(n131) );
  CIVX1 U226 ( .A(bitl[0]), .Z(net3640) );
  COND2XL U227 ( .A(n197), .B(n539), .C(n538), .D(n112), .Z(N88) );
  CIVXL U228 ( .A(bitl[2]), .Z(net14250) );
  CANR2XL U229 ( .A(n442), .B(n140), .C(n443), .D(n199), .Z(n359) );
  CAN2XL U230 ( .A(n196), .B(n562), .Z(N76) );
  COND1X1 U231 ( .A(n546), .B(net26430), .C(n303), .Z(n562) );
  CAN2X2 U232 ( .A(n210), .B(n108), .Z(bit2[28]) );
  CNIVX3 U233 ( .A(n209), .Z(n199) );
  CND2X2 U234 ( .A(net26601), .B(net3640), .Z(net11095) );
  CND2X2 U235 ( .A(bitl[0]), .B(net26601), .Z(net11166) );
  CIVX2 U236 ( .A(net17179), .Z(net26601) );
  CIVXL U237 ( .A(net26606), .Z(net26377) );
  CDLY1XL U238 ( .A(guess2[45]), .Z(n132) );
  CND2X2 U239 ( .A(n217), .B(net14606), .Z(n588) );
  CIVX1 U240 ( .A(net26437), .Z(net14606) );
  CIVXL U241 ( .A(net23249), .Z(net23250) );
  CDLY1XL U242 ( .A(guess2[57]), .Z(n133) );
  CDLY1XL U243 ( .A(guess2[52]), .Z(n134) );
  CDLY1XL U244 ( .A(guess2[59]), .Z(n135) );
  CNR2IX1 U245 ( .B(net17179), .A(n271), .Z(n491) );
  CIVXL U246 ( .A(net14249), .Z(net17171) );
  CIVXL U247 ( .A(n121), .Z(net14734) );
  COND3XL U248 ( .A(n233), .B(n599), .C(n232), .D(n272), .Z(N134) );
  CAN2X2 U249 ( .A(n590), .B(net14242), .Z(bit2[32]) );
  CDLY1XL U250 ( .A(guess2[60]), .Z(n138) );
  CAN2XL U251 ( .A(n196), .B(n563), .Z(N75) );
  CIVXL U252 ( .A(n563), .Z(n532) );
  CANR2XL U253 ( .A(n201), .B(n202), .C(n524), .D(n563), .Z(n495) );
  CAN2X1 U254 ( .A(n211), .B(net14241), .Z(bit2[40]) );
  CIVXL U255 ( .A(n219), .Z(n139) );
  CAN2X2 U256 ( .A(n592), .B(net13724), .Z(bit2[18]) );
  CIVX1 U257 ( .A(net11095), .Z(net10635) );
  CND2X1 U258 ( .A(n141), .B(n359), .Z(n564) );
  CNIVXL U259 ( .A(net11095), .Z(net14219) );
  CAN2X2 U260 ( .A(n592), .B(n596), .Z(bit2[22]) );
  CDLY1XL U261 ( .A(bitl[3]), .Z(net14615) );
  CIVX4 U262 ( .A(net11166), .Z(net13725) );
  CAN2X2 U263 ( .A(n103), .B(net13725), .Z(bit2[10]) );
  CIVX2 U264 ( .A(bitl[0]), .Z(net13671) );
  CIVX2 U265 ( .A(n570), .Z(n546) );
  COND2X2 U266 ( .A(n598), .B(n298), .C(net17171), .D(n377), .Z(n570) );
  CND2X2 U267 ( .A(n297), .B(n296), .Z(n377) );
  CND2XL U268 ( .A(n473), .B(net26430), .Z(n427) );
  CND2XL U269 ( .A(n524), .B(net26430), .Z(n508) );
  CND2XL U270 ( .A(n111), .B(net26430), .Z(net10816) );
  CND2XL U271 ( .A(n390), .B(net26430), .Z(n540) );
  COR2XL U272 ( .A(n218), .B(n551), .Z(n141) );
  COND3X1 U273 ( .A(acc[0]), .B(net13668), .C(n219), .D(n254), .Z(n551) );
  CND2XL U274 ( .A(n590), .B(n572), .Z(n553) );
  CAN2XL U275 ( .A(n590), .B(n108), .Z(bit2[36]) );
  CND2X2 U276 ( .A(bitl[3]), .B(net14250), .Z(n431) );
  CIVX2 U277 ( .A(n432), .Z(n590) );
  CND2X2 U278 ( .A(n593), .B(net10639), .Z(n594) );
  CANR2XL U279 ( .A(net14241), .B(n324), .C(net13725), .D(n323), .Z(n328) );
  CANR2XL U280 ( .A(net14241), .B(n323), .C(net13724), .D(n326), .Z(n245) );
  CANR2XL U281 ( .A(net14241), .B(n320), .C(net10636), .D(n319), .Z(n274) );
  CANR2XL U282 ( .A(net14241), .B(n332), .C(net10636), .D(n306), .Z(n284) );
  CANR2XL U283 ( .A(net14241), .B(n342), .C(net13724), .D(n341), .Z(n346) );
  CANR2XL U284 ( .A(net14241), .B(n305), .C(net10636), .D(n308), .Z(n243) );
  CANR2XL U285 ( .A(net14241), .B(n317), .C(net13725), .D(n320), .Z(n251) );
  CANR2XL U286 ( .A(net14241), .B(n344), .C(net13724), .D(n343), .Z(n276) );
  CANR2XL U287 ( .A(net14241), .B(n348), .C(net10636), .D(n347), .Z(n352) );
  CANR2XL U288 ( .A(net14241), .B(n347), .C(net10636), .D(n350), .Z(n256) );
  CANR2XL U289 ( .A(net14241), .B(n343), .C(net10636), .D(n348), .Z(n302) );
  CAN2X2 U290 ( .A(n589), .B(net14241), .Z(bit2[48]) );
  CAN2X1 U291 ( .A(n210), .B(net14241), .Z(bit2[24]) );
  CAN2X2 U292 ( .A(n595), .B(net10635), .Z(bit2[8]) );
  CND3X1 U293 ( .A(net14249), .B(net10644), .C(net10639), .Z(n513) );
  CAN2X2 U294 ( .A(n597), .B(net14651), .Z(bit2[4]) );
  CND2X2 U295 ( .A(net14606), .B(n198), .Z(n432) );
  CDLY1XL U296 ( .A(guess2[56]), .Z(n195) );
  CIVX2 U297 ( .A(net17179), .Z(net13668) );
  CIVXL U298 ( .A(n133), .Z(n581) );
  CND2XL U299 ( .A(net26437), .B(n572), .Z(n557) );
  CIVXL U300 ( .A(guess2[46]), .Z(n584) );
  CIVXL U301 ( .A(n135), .Z(n577) );
  CAN2X2 U302 ( .A(net23249), .B(n114), .Z(n198) );
  CIVX2 U303 ( .A(net14219), .Z(net14218) );
  CIVX2 U304 ( .A(net11095), .Z(net14241) );
  CIVX2 U305 ( .A(net11095), .Z(net14242) );
  CANR2XL U306 ( .A(n476), .B(n140), .C(n478), .D(n199), .Z(n353) );
  CANR2XL U307 ( .A(n575), .B(n483), .C(n456), .D(n217), .Z(n280) );
  CANR2XL U308 ( .A(n470), .B(n483), .C(n469), .D(n217), .Z(n471) );
  CANR2XL U309 ( .A(n463), .B(n483), .C(n462), .D(n217), .Z(n464) );
  CANR2XL U310 ( .A(n453), .B(n140), .C(n455), .D(n199), .Z(n281) );
  CANR2XL U311 ( .A(n493), .B(n140), .C(n461), .D(n199), .Z(n465) );
  CANR2XL U312 ( .A(n468), .B(n140), .C(n467), .D(n199), .Z(n472) );
  CIVXL U313 ( .A(guess2[58]), .Z(n579) );
  COND1XL U314 ( .A(n112), .B(n545), .C(n506), .Z(N101) );
  CIVXL U315 ( .A(n545), .Z(n420) );
  CAN2X1 U316 ( .A(n589), .B(net10636), .Z(bit2[50]) );
  CANR2XL U317 ( .A(n481), .B(n140), .C(n482), .D(n199), .Z(n330) );
  CAN2X1 U318 ( .A(n211), .B(n109), .Z(bit2[44]) );
  CMXI2XL U319 ( .A0(n598), .A1(n338), .S(net13671), .Z(n277) );
  CANR2XL U320 ( .A(n110), .B(n333), .C(n136), .D(n332), .Z(n334) );
  CIVX1 U321 ( .A(n363), .Z(n391) );
  COR2XL U322 ( .A(net14218), .B(n139), .Z(N130) );
  CMX2XL U323 ( .A0(n172), .A1(guess2[55]), .S(net14327), .Z(n89) );
  CMX2XL U324 ( .A0(n164), .A1(guess2[54]), .S(net14327), .Z(n88) );
  CMX2XL U325 ( .A0(n175), .A1(guess2[53]), .S(net14327), .Z(n87) );
  CMX2XL U326 ( .A0(n166), .A1(n134), .S(net14327), .Z(n86) );
  CMX2XL U327 ( .A0(n174), .A1(guess2[51]), .S(net14327), .Z(n85) );
  CMX2XL U328 ( .A0(n171), .A1(n104), .S(net14327), .Z(n84) );
  CMX2XL U329 ( .A0(n193), .A1(guess2[49]), .S(net14327), .Z(n83) );
  CMX2XL U330 ( .A0(n169), .A1(guess2[48]), .S(net14327), .Z(n82) );
  CMX2XL U331 ( .A0(n185), .A1(guess2[36]), .S(net14327), .Z(n70) );
  CMX2XL U332 ( .A0(n151), .A1(guess2[37]), .S(net14327), .Z(n71) );
  CMX2XL U333 ( .A0(n181), .A1(n105), .S(net14327), .Z(n72) );
  CMX2XL U334 ( .A0(n152), .A1(guess2[39]), .S(net14327), .Z(n73) );
  CMX2XL U335 ( .A0(n190), .A1(guess2[42]), .S(net14327), .Z(n76) );
  CMX2XL U336 ( .A0(n170), .A1(guess2[44]), .S(net14327), .Z(n78) );
  CMX2XL U337 ( .A0(n178), .A1(n132), .S(net14327), .Z(n79) );
  CMX2XL U338 ( .A0(n179), .A1(guess2[47]), .S(net14327), .Z(n81) );
  CMX2XL U339 ( .A0(n160), .A1(guess2[1]), .S(net14327), .Z(n35) );
  CMX2XL U340 ( .A0(n153), .A1(guess2[13]), .S(net14327), .Z(n47) );
  CMX2XL U341 ( .A0(n163), .A1(guess2[14]), .S(net14327), .Z(n48) );
  CMX2XL U342 ( .A0(n176), .A1(guess2[15]), .S(net14327), .Z(n49) );
  CMX2XL U343 ( .A0(n188), .A1(guess2[16]), .S(net14327), .Z(n50) );
  CMX2XL U344 ( .A0(n154), .A1(guess2[17]), .S(net14327), .Z(n51) );
  CMX2XL U345 ( .A0(n159), .A1(guess2[18]), .S(net14327), .Z(n52) );
  CMX2XL U346 ( .A0(n150), .A1(guess2[19]), .S(net14327), .Z(n53) );
  CMX2XL U347 ( .A0(n192), .A1(guess2[20]), .S(net14327), .Z(n54) );
  CMX2XL U348 ( .A0(n146), .A1(guess2[21]), .S(net14327), .Z(n55) );
  CMX2XL U349 ( .A0(n157), .A1(guess2[22]), .S(net14327), .Z(n56) );
  CMX2XL U350 ( .A0(n143), .A1(guess2[23]), .S(net14327), .Z(n57) );
  CMX2XL U351 ( .A0(n156), .A1(guess2[24]), .S(net14327), .Z(n58) );
  CMX2XL U352 ( .A0(n182), .A1(guess2[12]), .S(net14327), .Z(n46) );
  CMX2XL U353 ( .A0(n148), .A1(guess2[11]), .S(net14327), .Z(n45) );
  CMX2XL U354 ( .A0(n186), .A1(guess2[10]), .S(net14327), .Z(n44) );
  CMX2XL U355 ( .A0(n194), .A1(guess2[9]), .S(net14327), .Z(n43) );
  CMX2XL U356 ( .A0(n165), .A1(guess2[8]), .S(net14327), .Z(n42) );
  CMX2XL U357 ( .A0(n167), .A1(guess2[6]), .S(net14327), .Z(n40) );
  CMX2XL U358 ( .A0(n147), .A1(guess2[5]), .S(net14327), .Z(n39) );
  CMX2XL U359 ( .A0(n168), .A1(guess2[4]), .S(net14327), .Z(n38) );
  CMX2XL U360 ( .A0(n173), .A1(guess2[3]), .S(net14327), .Z(n37) );
  CMX2XL U361 ( .A0(n191), .A1(guess2[2]), .S(net14327), .Z(n36) );
  CMX2XL U362 ( .A0(n183), .A1(guess2[26]), .S(net14327), .Z(n60) );
  CMX2XL U363 ( .A0(n149), .A1(guess2[27]), .S(net14327), .Z(n61) );
  CMX2XL U364 ( .A0(n189), .A1(guess2[29]), .S(net14327), .Z(n63) );
  CMX2XL U365 ( .A0(n155), .A1(guess2[30]), .S(net14327), .Z(n64) );
  CMX2XL U366 ( .A0(n180), .A1(guess2[31]), .S(net14327), .Z(n65) );
  CMX2XL U367 ( .A0(n158), .A1(guess2[32]), .S(net14327), .Z(n66) );
  CMX2XL U368 ( .A0(n142), .A1(guess2[33]), .S(net14327), .Z(n67) );
  CMX2XL U369 ( .A0(n177), .A1(guess2[0]), .S(net14327), .Z(n34) );
  CMX2XL U370 ( .A0(n184), .A1(guess2[34]), .S(net14327), .Z(n68) );
  CMX2XL U371 ( .A0(n187), .A1(guess2[35]), .S(net14327), .Z(n69) );
  CMX2XL U372 ( .A0(n144), .A1(n138), .S(net14327), .Z(n94) );
  CMX2XL U373 ( .A0(n145), .A1(guess2[61]), .S(net14327), .Z(n95) );
  CMX2XL U374 ( .A0(n162), .A1(guess2[62]), .S(net14327), .Z(n96) );
  CMX2XL U375 ( .A0(n161), .A1(guess2[63]), .S(net14327), .Z(n98) );
  CND2IXL U376 ( .B(n393), .A(acc[31]), .Z(n394) );
  CMXI2XL U377 ( .A0(acc[30]), .A1(acc[31]), .S(net13671), .Z(n271) );
  CMX2XL U378 ( .A0(n493), .A1(n461), .S(net14734), .Z(n215) );
  CMX2XL U379 ( .A0(n491), .A1(n448), .S(net14734), .Z(n214) );
  CMX2XL U380 ( .A0(n202), .A1(n481), .S(net14734), .Z(n216) );
  COND1XL U381 ( .A(n558), .B(n224), .C(n525), .Z(N96) );
  COND1XL U382 ( .A(n112), .B(n537), .C(n499), .Z(N105) );
  COND1XL U383 ( .A(n541), .B(n489), .C(n392), .Z(N119) );
  COND1XL U384 ( .A(n112), .B(n541), .C(n502), .Z(N103) );
  COND1XL U385 ( .A(n203), .B(n489), .C(n354), .Z(N123) );
  COND1XL U386 ( .A(n537), .B(n489), .C(n370), .Z(N121) );
  COND1XL U387 ( .A(n498), .B(n363), .C(n362), .Z(N122) );
  COND1XL U388 ( .A(n205), .B(n489), .C(n282), .Z(N125) );
  COND1XL U389 ( .A(n204), .B(n489), .C(n304), .Z(N124) );
  COND1XL U390 ( .A(n552), .B(n224), .C(n521), .Z(N97) );
  COND1XL U391 ( .A(n498), .B(n497), .C(n496), .Z(N106) );
  CIVX2 U392 ( .A(n272), .Z(n473) );
  COND1XL U393 ( .A(n393), .B(n234), .C(n116), .Z(n2) );
  COND1XL U394 ( .A(n238), .B(n234), .C(n101), .Z(n3) );
  COND1XL U395 ( .A(n239), .B(n234), .C(n100), .Z(n4) );
  COND1XL U396 ( .A(n298), .B(n234), .C(n332), .Z(n5) );
  COND1XL U397 ( .A(n357), .B(n234), .C(n306), .Z(n6) );
  COND1XL U398 ( .A(n235), .B(n234), .C(n305), .Z(n7) );
  COND1XL U399 ( .A(n236), .B(n234), .C(n308), .Z(n8) );
  COND1XL U400 ( .A(n599), .B(n234), .C(n307), .Z(n9) );
  COND1XL U401 ( .A(n393), .B(n600), .C(n348), .Z(n26) );
  COND1XL U402 ( .A(n238), .B(n221), .C(n347), .Z(n27) );
  COND1XL U403 ( .A(n239), .B(n221), .C(n350), .Z(n28) );
  COND1XL U404 ( .A(n298), .B(n600), .C(n349), .Z(n29) );
  COND1XL U405 ( .A(n357), .B(n222), .C(n337), .Z(n30) );
  COND1XL U406 ( .A(n235), .B(n221), .C(n336), .Z(n31) );
  COND1XL U407 ( .A(n236), .B(n222), .C(n338), .Z(n32) );
  COND1XL U408 ( .A(n599), .B(n600), .C(n598), .Z(n33) );
  COND1XL U409 ( .A(n128), .B(n238), .C(n311), .Z(n11) );
  COND1XL U410 ( .A(n239), .B(n129), .C(n314), .Z(n12) );
  COND1XL U411 ( .A(n130), .B(n235), .C(n323), .Z(n15) );
  COND1XL U412 ( .A(n236), .B(n129), .C(n326), .Z(n16) );
  COND1XL U413 ( .A(n393), .B(n237), .C(n318), .Z(n18) );
  COND1XL U414 ( .A(n599), .B(n237), .C(n343), .Z(n25) );
  COND1XL U415 ( .A(n393), .B(n130), .C(n312), .Z(n10) );
  COND1XL U416 ( .A(n298), .B(n128), .C(n313), .Z(n13) );
  COND1XL U417 ( .A(n357), .B(n128), .C(n324), .Z(n14) );
  COND1XL U418 ( .A(n599), .B(n130), .C(n325), .Z(n17) );
  CAN2XL U419 ( .A(n102), .B(n139), .Z(n200) );
  CAN2XL U420 ( .A(n210), .B(n572), .Z(n201) );
  CAN2X1 U421 ( .A(n335), .B(n334), .Z(n202) );
  CAN2X1 U422 ( .A(n330), .B(n329), .Z(n203) );
  CAN2X1 U423 ( .A(n292), .B(n291), .Z(n204) );
  CAN2X1 U424 ( .A(n270), .B(n269), .Z(n205) );
  CAN2XL U425 ( .A(n597), .B(n572), .Z(n206) );
  CAN2XL U426 ( .A(n102), .B(n572), .Z(n207) );
  CAN2X1 U427 ( .A(n486), .B(n485), .Z(n208) );
  COND1XL U428 ( .A(n378), .B(net26430), .C(n231), .Z(N132) );
  CNIVX1 U429 ( .A(n601), .Z(n226) );
  CNIVX1 U430 ( .A(n601), .Z(n227) );
  CNIVX1 U431 ( .A(n601), .Z(n225) );
  CNIVX1 U432 ( .A(n601), .Z(n228) );
  CNIVX1 U433 ( .A(n601), .Z(n229) );
  CNIVX1 U434 ( .A(n601), .Z(n230) );
  CND4XL U435 ( .A(n369), .B(n368), .C(n367), .D(n396), .Z(n536) );
  CND2XL U436 ( .A(n140), .B(n417), .Z(n369) );
  CAN2XL U437 ( .A(rdy), .B(n597), .Z(n212) );
  CAN2XL U438 ( .A(rdy), .B(n590), .Z(n213) );
  CIVDX4 U439 ( .A(n431), .Z0(n217), .Z1(n218) );
  CIVXL U440 ( .A(n358), .Z(n498) );
  CANR2XL U441 ( .A(n438), .B(n483), .C(n437), .D(n217), .Z(n439) );
  CIVX2 U442 ( .A(net11166), .Z(net13724) );
  CIVX2 U443 ( .A(net11166), .Z(net10636) );
  CIVXL U444 ( .A(n136), .Z(n219) );
  CIVXL U445 ( .A(n136), .Z(n220) );
  CIVXL U446 ( .A(n564), .Z(n534) );
  CANR2XL U447 ( .A(n524), .B(n564), .C(n111), .D(n533), .Z(n496) );
  CANR2XL U448 ( .A(n473), .B(n564), .C(n524), .D(n533), .Z(n362) );
  CIVXL U449 ( .A(net14241), .Z(net13702) );
  CIVXL U450 ( .A(n562), .Z(n531) );
  CANR2XL U451 ( .A(n201), .B(n493), .C(n524), .D(n562), .Z(n494) );
  CANR2XL U452 ( .A(n207), .B(n493), .C(n473), .D(n562), .Z(n304) );
  CIVXL U453 ( .A(guess2[40]), .Z(n586) );
  CND2XL U454 ( .A(n277), .B(net13668), .Z(n554) );
  CAN2X2 U455 ( .A(n211), .B(n136), .Z(bit2[46]) );
  COND1XL U456 ( .A(n235), .B(n237), .C(n341), .Z(n23) );
  COND1XL U457 ( .A(n236), .B(n237), .C(n344), .Z(n24) );
  COND1XL U458 ( .A(n238), .B(n237), .C(n317), .Z(n19) );
  COND1XL U459 ( .A(n239), .B(n237), .C(n320), .Z(n20) );
  COND1XL U460 ( .A(n298), .B(n237), .C(n319), .Z(n21) );
  COND1XL U461 ( .A(n357), .B(n237), .C(n342), .Z(n22) );
  CND2XL U462 ( .A(net31721), .B(n571), .Z(n221) );
  CND2IX1 U463 ( .B(n363), .A(net31721), .Z(n234) );
  CND2IX1 U464 ( .B(n497), .A(net31721), .Z(n237) );
  CAN2XL U465 ( .A(n571), .B(n570), .Z(N68) );
  CAN2X2 U466 ( .A(n596), .B(n597), .Z(bit2[6]) );
  CAN2XL U467 ( .A(n592), .B(net14651), .Z(bit2[20]) );
  CND2XL U468 ( .A(rdy), .B(net10644), .Z(n489) );
  CANR2XL U469 ( .A(n467), .B(n140), .C(n469), .D(n199), .Z(n303) );
  CANR2XL U470 ( .A(net13668), .B(n356), .C(net13656), .D(n331), .Z(n293) );
  CANR2XL U471 ( .A(n448), .B(n140), .C(n449), .D(n199), .Z(n270) );
  CANR2XL U472 ( .A(n398), .B(n140), .C(n437), .D(n199), .Z(n249) );
  CANR2XL U473 ( .A(n202), .B(n140), .C(n481), .D(n199), .Z(n486) );
  CANR2XL U474 ( .A(n140), .B(n384), .C(n199), .D(n383), .Z(n388) );
  CANR2XL U475 ( .A(n140), .B(n372), .C(n199), .D(n371), .Z(n376) );
  CANR2XL U476 ( .A(n140), .B(n364), .C(n199), .D(n415), .Z(n366) );
  CANR2XL U477 ( .A(n437), .B(n140), .C(n438), .D(n199), .Z(n361) );
  CANR2XL U478 ( .A(n491), .B(n199), .C(n449), .D(n483), .Z(n410) );
  CANR2XL U479 ( .A(n140), .B(n402), .C(n199), .D(n401), .Z(n406) );
  CANR2XL U480 ( .A(n202), .B(n199), .C(n482), .D(n483), .Z(n429) );
  CANR2XL U481 ( .A(n463), .B(n140), .C(n468), .D(n199), .Z(n426) );
  CANR2XL U482 ( .A(n140), .B(n415), .C(n199), .D(n414), .Z(n419) );
  CANR2XL U483 ( .A(n461), .B(n140), .C(n462), .D(n199), .Z(n292) );
  CANR2XL U484 ( .A(n493), .B(n199), .C(n462), .D(n483), .Z(n423) );
  CANR2XL U485 ( .A(n484), .B(n140), .C(n477), .D(n199), .Z(n434) );
  CANR2XL U486 ( .A(n454), .B(n140), .C(n453), .D(n199), .Z(n458) );
  CANR2XL U487 ( .A(n477), .B(n140), .C(n476), .D(n199), .Z(n480) );
  CANR2XL U488 ( .A(n441), .B(n140), .C(n440), .D(n199), .Z(n445) );
  CANR2XL U489 ( .A(n440), .B(n140), .C(n442), .D(n199), .Z(n258) );
  CANR2XL U490 ( .A(n491), .B(n140), .C(n448), .D(n199), .Z(n452) );
  CEOXL U491 ( .A(n107), .B(n466), .Z(N133) );
  CND2XL U492 ( .A(rdy), .B(n107), .Z(n272) );
  CND2XL U493 ( .A(n107), .B(n572), .Z(n555) );
  CND2XL U494 ( .A(net14327), .B(n571), .Z(n222) );
  CND2XL U495 ( .A(net13724), .B(n121), .Z(n236) );
  CND2XL U496 ( .A(net26813), .B(n121), .Z(n235) );
  COND1XL U497 ( .A(n470), .B(net23249), .C(n381), .Z(n538) );
  COND2XL U498 ( .A(n357), .B(n356), .C(net23249), .D(n355), .Z(n358) );
  CND2XL U499 ( .A(n136), .B(n121), .Z(n357) );
  CND2XL U500 ( .A(net14615), .B(n196), .Z(n497) );
  CND2XL U501 ( .A(n111), .B(net14615), .Z(n363) );
  COND1XL U502 ( .A(net14615), .B(n498), .C(n439), .Z(n517) );
  COND2XL U503 ( .A(n396), .B(n395), .C(net14615), .D(n394), .Z(n397) );
  CND2XL U504 ( .A(net14615), .B(n554), .Z(n368) );
  CANR2XL U505 ( .A(net14615), .B(n380), .C(n140), .D(n379), .Z(n381) );
  CIVXL U506 ( .A(n195), .Z(n223) );
  COND1XL U507 ( .A(net14218), .B(n121), .C(n599), .Z(N131) );
  COND3XL U508 ( .A(acc[29]), .B(n220), .C(net13702), .D(n293), .Z(n295) );
  CND2XL U509 ( .A(net17171), .B(n412), .Z(n367) );
  CMXI2XL U510 ( .A0(n399), .A1(n551), .S(net17171), .Z(n400) );
  CMXI2XL U511 ( .A0(n389), .A1(n549), .S(net17171), .Z(n390) );
  CMXI2XL U512 ( .A0(n412), .A1(n554), .S(net17171), .Z(n413) );
  CND2XL U513 ( .A(net23250), .B(net14242), .Z(n298) );
  CND2XL U514 ( .A(net13724), .B(net14734), .Z(n239) );
  CND2XL U515 ( .A(net14734), .B(net26813), .Z(n238) );
  CND2XL U516 ( .A(net17171), .B(n136), .Z(n393) );
  CND2XL U517 ( .A(bitl[3]), .B(net23250), .Z(n396) );
  COND1XL U518 ( .A(n218), .B(n411), .C(n410), .Z(n505) );
  COND1XL U519 ( .A(n218), .B(n430), .C(n429), .Z(n514) );
  COND1XL U520 ( .A(n218), .B(n424), .C(n423), .Z(n507) );
  CIVX2 U521 ( .A(n111), .Z(n224) );
  CIVX2 U522 ( .A(reset), .Z(n601) );
  CND2X1 U523 ( .A(bitl[0]), .B(net17179), .Z(n294) );
  CND2X1 U524 ( .A(net14242), .B(n121), .Z(n599) );
  CIVX2 U525 ( .A(n599), .Z(n378) );
  CND2X1 U526 ( .A(n378), .B(net26430), .Z(n231) );
  CIVX2 U527 ( .A(n231), .Z(n466) );
  CND2X1 U528 ( .A(n196), .B(net26430), .Z(n233) );
  CND2X1 U529 ( .A(rdy), .B(n231), .Z(n232) );
  CIVX2 U530 ( .A(n497), .Z(n501) );
  CIVX2 U531 ( .A(n233), .Z(n571) );
  CIVX2 U532 ( .A(net10816), .Z(net11163) );
  CANR2X1 U533 ( .A(n110), .B(n332), .C(n136), .D(n306), .Z(n240) );
  CND2X1 U534 ( .A(n241), .B(n240), .Z(n355) );
  CIVX2 U535 ( .A(n355), .Z(n398) );
  CANR2X1 U536 ( .A(n110), .B(n307), .C(n136), .D(n312), .Z(n242) );
  CND2X1 U537 ( .A(n243), .B(n242), .Z(n395) );
  CIVX2 U538 ( .A(n395), .Z(n437) );
  CANR2X1 U539 ( .A(n110), .B(n325), .C(n136), .D(n318), .Z(n244) );
  CND2X1 U540 ( .A(n245), .B(n244), .Z(n401) );
  CIVX2 U541 ( .A(n401), .Z(n441) );
  CANR2X1 U542 ( .A(net14242), .B(n311), .C(net13725), .D(n314), .Z(n247) );
  CANR2X1 U543 ( .A(n109), .B(n313), .C(n136), .D(n324), .Z(n246) );
  CND2X1 U544 ( .A(n247), .B(n246), .Z(n402) );
  CIVX2 U545 ( .A(n402), .Z(n438) );
  CND2X1 U546 ( .A(n249), .B(n248), .Z(n527) );
  CANR2X1 U547 ( .A(n109), .B(n319), .C(n136), .D(n342), .Z(n250) );
  CND2X1 U548 ( .A(n251), .B(n250), .Z(n403) );
  CIVX2 U549 ( .A(n403), .Z(n440) );
  CANR2X1 U550 ( .A(net14242), .B(n341), .C(net13724), .D(n344), .Z(n253) );
  CANR2X1 U551 ( .A(n110), .B(n343), .C(n136), .D(n348), .Z(n252) );
  CND2X1 U552 ( .A(n253), .B(n252), .Z(n404) );
  CIVX2 U553 ( .A(n404), .Z(n442) );
  CIVX2 U554 ( .A(n551), .Z(n574) );
  CANR2X1 U555 ( .A(n110), .B(n349), .C(n136), .D(n337), .Z(n255) );
  CND2X1 U556 ( .A(n256), .B(n255), .Z(n399) );
  CIVX2 U557 ( .A(n399), .Z(n443) );
  CANR2X1 U558 ( .A(n574), .B(n483), .C(n443), .D(n217), .Z(n257) );
  CND2X1 U559 ( .A(n258), .B(n257), .Z(n560) );
  CIVX2 U560 ( .A(n560), .Z(n528) );
  CND2X1 U561 ( .A(n200), .B(acc[31]), .Z(n259) );
  COND2X1 U562 ( .A(n528), .B(n272), .C(rdy), .D(n259), .Z(n260) );
  CAOR1X1 U563 ( .A(n524), .B(n527), .C(n260), .Z(N126) );
  CANR2X1 U564 ( .A(n110), .B(n306), .C(n136), .D(n305), .Z(n261) );
  CND2X1 U565 ( .A(n262), .B(n261), .Z(n411) );
  CIVX2 U566 ( .A(n411), .Z(n448) );
  CANR2X1 U567 ( .A(net14218), .B(n308), .C(net13725), .D(n307), .Z(n264) );
  CANR2X1 U568 ( .A(n110), .B(n312), .C(n136), .D(n311), .Z(n263) );
  CND2X1 U569 ( .A(n264), .B(n263), .Z(n364) );
  CIVX2 U570 ( .A(n364), .Z(n449) );
  CANR2X1 U571 ( .A(net14218), .B(n326), .C(net13724), .D(n325), .Z(n266) );
  CANR2X1 U572 ( .A(n110), .B(n318), .C(n136), .D(n317), .Z(n265) );
  CND2X1 U573 ( .A(n266), .B(n265), .Z(n414) );
  CIVX2 U574 ( .A(n414), .Z(n454) );
  CANR2X1 U575 ( .A(net14218), .B(n314), .C(net13725), .D(n313), .Z(n268) );
  CANR2X1 U576 ( .A(n109), .B(n324), .C(n136), .D(n323), .Z(n267) );
  CND2X1 U577 ( .A(n268), .B(n267), .Z(n415) );
  CIVX2 U578 ( .A(n415), .Z(n450) );
  CANR2X1 U579 ( .A(n109), .B(n342), .C(n136), .D(n341), .Z(n273) );
  CND2X1 U580 ( .A(n274), .B(n273), .Z(n416) );
  CIVX2 U581 ( .A(n416), .Z(n453) );
  CANR2X1 U582 ( .A(n109), .B(n348), .C(n136), .D(n347), .Z(n275) );
  CND2X1 U583 ( .A(n276), .B(n275), .Z(n417) );
  CIVX2 U584 ( .A(n417), .Z(n455) );
  CIVX2 U585 ( .A(n554), .Z(n575) );
  CANR2X1 U586 ( .A(net14242), .B(n350), .C(net13725), .D(n349), .Z(n279) );
  CANR2X1 U587 ( .A(n110), .B(n337), .C(n136), .D(n336), .Z(n278) );
  CND2X1 U588 ( .A(n279), .B(n278), .Z(n412) );
  CIVX2 U589 ( .A(n412), .Z(n456) );
  CND2X1 U590 ( .A(n281), .B(n280), .Z(n561) );
  CANR2X1 U591 ( .A(n207), .B(n491), .C(n473), .D(n561), .Z(n282) );
  CANR2X1 U592 ( .A(n110), .B(n305), .C(n136), .D(n308), .Z(n283) );
  CND2X1 U593 ( .A(n284), .B(n283), .Z(n424) );
  CIVX2 U594 ( .A(n424), .Z(n461) );
  CANR2X1 U595 ( .A(net14242), .B(n307), .C(net13724), .D(n312), .Z(n286) );
  CANR2X1 U596 ( .A(n109), .B(n311), .C(n136), .D(n314), .Z(n285) );
  CND2X1 U597 ( .A(n286), .B(n285), .Z(n372) );
  CIVX2 U598 ( .A(n372), .Z(n462) );
  CANR2X1 U599 ( .A(net14242), .B(n325), .C(net13725), .D(n318), .Z(n288) );
  CANR2X1 U600 ( .A(n109), .B(n317), .C(n136), .D(n320), .Z(n287) );
  CND2X1 U601 ( .A(n288), .B(n287), .Z(n373) );
  CIVX2 U602 ( .A(n373), .Z(n468) );
  CANR2X1 U603 ( .A(n110), .B(n323), .C(n136), .D(n326), .Z(n289) );
  CND2X1 U604 ( .A(n290), .B(n289), .Z(n371) );
  CIVX2 U605 ( .A(n371), .Z(n463) );
  CIVX2 U606 ( .A(n295), .Z(n493) );
  CANR2X1 U607 ( .A(net14242), .B(n319), .C(net13725), .D(n342), .Z(n300) );
  CANR2X1 U608 ( .A(n109), .B(n341), .C(n136), .D(n344), .Z(n299) );
  CND2X1 U609 ( .A(n300), .B(n299), .Z(n374) );
  CIVX2 U610 ( .A(n374), .Z(n467) );
  CANR2X1 U611 ( .A(n109), .B(n347), .C(n136), .D(n350), .Z(n301) );
  CND2X1 U612 ( .A(n302), .B(n301), .Z(n379) );
  CANR2X1 U613 ( .A(net14218), .B(n306), .C(net13725), .D(n305), .Z(n310) );
  CANR2X1 U614 ( .A(n109), .B(n308), .C(n136), .D(n307), .Z(n309) );
  CND2X1 U615 ( .A(n310), .B(n309), .Z(n430) );
  CIVX2 U616 ( .A(n430), .Z(n481) );
  CANR2X1 U617 ( .A(n110), .B(n314), .C(n136), .D(n313), .Z(n315) );
  CND2X1 U618 ( .A(n316), .B(n315), .Z(n384) );
  CIVX2 U619 ( .A(n384), .Z(n482) );
  CANR2X1 U620 ( .A(n109), .B(n320), .C(n136), .D(n319), .Z(n321) );
  CND2X1 U621 ( .A(n322), .B(n321), .Z(n385) );
  CIVX2 U622 ( .A(n385), .Z(n477) );
  CANR2X1 U623 ( .A(n109), .B(n326), .C(n136), .D(n325), .Z(n327) );
  CND2X1 U624 ( .A(n328), .B(n327), .Z(n383) );
  CIVX2 U625 ( .A(n383), .Z(n484) );
  CANR2X1 U626 ( .A(net14218), .B(n356), .C(net13724), .D(n331), .Z(n335) );
  CANR2X1 U627 ( .A(n110), .B(n338), .C(n136), .D(n598), .Z(n339) );
  CND2X1 U628 ( .A(n340), .B(n339), .Z(n549) );
  CANR2X1 U629 ( .A(n110), .B(n344), .C(n136), .D(n343), .Z(n345) );
  CND2X1 U630 ( .A(n346), .B(n345), .Z(n386) );
  CIVX2 U631 ( .A(n386), .Z(n476) );
  CANR2X1 U632 ( .A(n109), .B(n350), .C(n136), .D(n349), .Z(n351) );
  CND2X1 U633 ( .A(n352), .B(n351), .Z(n389) );
  CIVX2 U634 ( .A(n389), .Z(n478) );
  CANR2X1 U635 ( .A(n207), .B(n202), .C(n473), .D(n563), .Z(n354) );
  CND2X1 U636 ( .A(n361), .B(n360), .Z(n533) );
  CND2X1 U637 ( .A(n366), .B(n365), .Z(n537) );
  CIVX2 U638 ( .A(n536), .Z(n565) );
  CANR2X1 U639 ( .A(n391), .B(n214), .C(n473), .D(n565), .Z(n370) );
  CND2X1 U640 ( .A(n376), .B(n375), .Z(n539) );
  CND2X1 U641 ( .A(acc[0]), .B(n378), .Z(n380) );
  CIVX2 U642 ( .A(n538), .Z(n566) );
  CANR2X1 U643 ( .A(n391), .B(n215), .C(n473), .D(n566), .Z(n382) );
  CND2X1 U644 ( .A(n388), .B(n387), .Z(n541) );
  CIVX2 U645 ( .A(n540), .Z(n567) );
  CANR2X1 U646 ( .A(n391), .B(n216), .C(n473), .D(n567), .Z(n392) );
  CIVX2 U647 ( .A(n503), .Z(n409) );
  CND2X1 U648 ( .A(n400), .B(net26430), .Z(n542) );
  CIVX2 U649 ( .A(n542), .Z(n568) );
  CND2X1 U650 ( .A(n406), .B(n405), .Z(n543) );
  CIVX2 U651 ( .A(n543), .Z(n407) );
  CANR2X1 U652 ( .A(n473), .B(n568), .C(n524), .D(n407), .Z(n408) );
  COND1X1 U653 ( .A(n409), .B(n224), .C(n408), .Z(N118) );
  CIVX2 U654 ( .A(n505), .Z(n422) );
  CND2X1 U655 ( .A(n413), .B(net26430), .Z(n544) );
  CIVX2 U656 ( .A(n544), .Z(n569) );
  CND2X1 U657 ( .A(n419), .B(n418), .Z(n545) );
  CANR2X1 U658 ( .A(n473), .B(n569), .C(n524), .D(n420), .Z(n421) );
  CND2X1 U659 ( .A(n426), .B(n425), .Z(n511) );
  CIVX2 U660 ( .A(n511), .Z(n547) );
  CAOR1X1 U661 ( .A(n111), .B(n507), .C(n428), .Z(N116) );
  CIVX2 U662 ( .A(n514), .Z(n436) );
  CIVX2 U663 ( .A(n549), .Z(n573) );
  CANR2X1 U664 ( .A(n478), .B(n483), .C(n476), .D(n217), .Z(n433) );
  CND2X1 U665 ( .A(n434), .B(n433), .Z(n512) );
  CANR2X1 U666 ( .A(n213), .B(n573), .C(n524), .D(n512), .Z(n435) );
  COND1X1 U667 ( .A(n436), .B(n224), .C(n435), .Z(N115) );
  CIVX2 U668 ( .A(n517), .Z(n447) );
  CANR2X1 U669 ( .A(n443), .B(n483), .C(n442), .D(n217), .Z(n444) );
  CND2X1 U670 ( .A(n445), .B(n444), .Z(n516) );
  CANR2X1 U671 ( .A(n213), .B(n574), .C(n524), .D(n516), .Z(n446) );
  COND1X1 U672 ( .A(n447), .B(n224), .C(n446), .Z(N114) );
  CND2X1 U673 ( .A(n452), .B(n451), .Z(n520) );
  CIVX2 U674 ( .A(n520), .Z(n460) );
  CANR2X1 U675 ( .A(n456), .B(n483), .C(n455), .D(n217), .Z(n457) );
  CND2X1 U676 ( .A(n458), .B(n457), .Z(n519) );
  CANR2X1 U677 ( .A(n213), .B(n575), .C(n524), .D(n519), .Z(n459) );
  CND2X1 U678 ( .A(n465), .B(n464), .Z(n523) );
  CIVX2 U679 ( .A(n523), .Z(n475) );
  CND2X1 U680 ( .A(n466), .B(acc[0]), .Z(n556) );
  CIVX2 U681 ( .A(n556), .Z(n576) );
  CND2X1 U682 ( .A(n472), .B(n471), .Z(n522) );
  CANR2X1 U683 ( .A(n473), .B(n576), .C(n524), .D(n522), .Z(n474) );
  COND1X1 U684 ( .A(n475), .B(n224), .C(n474), .Z(N112) );
  CANR2X1 U685 ( .A(n573), .B(n483), .C(n478), .D(n217), .Z(n479) );
  CND2X1 U686 ( .A(n480), .B(n479), .Z(n559) );
  CIVX2 U687 ( .A(n559), .Z(n526) );
  CND2X1 U688 ( .A(n113), .B(acc[31]), .Z(n488) );
  CAOR1X1 U689 ( .A(n111), .B(n527), .C(n490), .Z(N110) );
  CANR2X1 U690 ( .A(n201), .B(n491), .C(n524), .D(n561), .Z(n492) );
  COND1X1 U691 ( .A(n204), .B(n224), .C(n494), .Z(N108) );
  CANR2X1 U692 ( .A(n501), .B(n214), .C(n524), .D(n565), .Z(n499) );
  CANR2X1 U693 ( .A(n501), .B(n215), .C(n524), .D(n566), .Z(n500) );
  COND1X1 U694 ( .A(n112), .B(n539), .C(n500), .Z(N104) );
  CANR2X1 U695 ( .A(n501), .B(n216), .C(n524), .D(n567), .Z(n502) );
  CANR2X1 U696 ( .A(n524), .B(n568), .C(n196), .D(n503), .Z(n504) );
  COND1X1 U697 ( .A(n112), .B(n543), .C(n504), .Z(N102) );
  CANR2X1 U698 ( .A(n524), .B(n569), .C(n196), .D(n505), .Z(n506) );
  CIVX2 U699 ( .A(n507), .Z(n509) );
  COND2X1 U700 ( .A(n509), .B(n197), .C(n546), .D(n508), .Z(n510) );
  CAOR1X1 U701 ( .A(n111), .B(n511), .C(n510), .Z(N100) );
  CIVX2 U702 ( .A(n512), .Z(n548) );
  CIVX2 U703 ( .A(n513), .Z(n597) );
  CANR2X1 U704 ( .A(n212), .B(n573), .C(n196), .D(n514), .Z(n515) );
  COND1X1 U705 ( .A(n548), .B(n224), .C(n515), .Z(N99) );
  CIVX2 U706 ( .A(n516), .Z(n550) );
  CANR2X1 U707 ( .A(n212), .B(n574), .C(n196), .D(n517), .Z(n518) );
  CIVX2 U708 ( .A(n519), .Z(n552) );
  CANR2X1 U709 ( .A(n212), .B(n575), .C(n196), .D(n520), .Z(n521) );
  CANR2X1 U710 ( .A(n524), .B(n576), .C(n196), .D(n523), .Z(n525) );
  COND2X1 U711 ( .A(n208), .B(n197), .C(n526), .D(n224), .Z(N95) );
  CIVX2 U712 ( .A(n527), .Z(n529) );
  COND2X1 U713 ( .A(n529), .B(n197), .C(n528), .D(n224), .Z(N94) );
  CIVX2 U714 ( .A(n561), .Z(n530) );
  COND2X1 U715 ( .A(n205), .B(n197), .C(n530), .D(n224), .Z(N93) );
  COND2X1 U716 ( .A(n204), .B(n197), .C(n531), .D(n224), .Z(N92) );
  COND2X1 U717 ( .A(n203), .B(n197), .C(n532), .D(n224), .Z(N91) );
  CIVX2 U718 ( .A(n533), .Z(n535) );
  COND2X1 U719 ( .A(n535), .B(n197), .C(n534), .D(n112), .Z(N90) );
  COND2X1 U720 ( .A(n197), .B(n541), .C(n540), .D(n112), .Z(N87) );
  COND2X1 U721 ( .A(n197), .B(n543), .C(n542), .D(n112), .Z(N86) );
  COND2X1 U722 ( .A(n197), .B(n545), .C(n544), .D(n112), .Z(N85) );
  COND2X1 U723 ( .A(n547), .B(n197), .C(n546), .D(net10816), .Z(N84) );
  COND2X1 U724 ( .A(n549), .B(n553), .C(n548), .D(n197), .Z(N83) );
  COND2X1 U725 ( .A(n551), .B(n553), .C(n550), .D(n197), .Z(N82) );
  COND2X1 U726 ( .A(n554), .B(n553), .C(n552), .D(n197), .Z(N81) );
  COND2X1 U727 ( .A(n558), .B(n197), .C(n556), .D(n112), .Z(N80) );
  CAN2X1 U728 ( .A(n196), .B(n559), .Z(N79) );
  CAN2X1 U729 ( .A(n196), .B(n560), .Z(N78) );
  CAN2X1 U730 ( .A(n196), .B(n561), .Z(N77) );
  CAN2X1 U731 ( .A(n566), .B(n196), .Z(N72) );
  CAN2X1 U732 ( .A(n567), .B(n196), .Z(N71) );
  CAN2X1 U733 ( .A(n568), .B(n196), .Z(N70) );
  CAN2X1 U734 ( .A(n569), .B(n196), .Z(N69) );
  CAN2X1 U735 ( .A(n573), .B(n206), .Z(N67) );
  CAN2X1 U736 ( .A(n574), .B(n206), .Z(N66) );
  CAN2X1 U737 ( .A(n206), .B(n575), .Z(N65) );
  CAN2X1 U738 ( .A(n576), .B(n196), .Z(N64) );
  CAN2X1 U739 ( .A(n102), .B(net26813), .Z(bit2[60]) );
  CAN2X1 U740 ( .A(n102), .B(net14218), .Z(bit2[56]) );
  CIVX2 U741 ( .A(n588), .Z(n589) );
  CAN2X1 U742 ( .A(n589), .B(n136), .Z(bit2[54]) );
  CAN2X1 U743 ( .A(n589), .B(n109), .Z(bit2[52]) );
  CAN2X1 U744 ( .A(n211), .B(net13725), .Z(bit2[42]) );
  CAN2X1 U745 ( .A(n590), .B(n596), .Z(bit2[38]) );
  CIVX2 U746 ( .A(n594), .Z(n595) );
endmodule

