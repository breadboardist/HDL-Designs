
module sfilt_DW01_add_2 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n6, n8, n9, n10, n11, n12, n13, n14, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n88, n89, n90, n91, n92, n93, n95, n96, n97, n98, n99,
         n100, n103, n104, n105, n106, n107, n108, n109, n110, n113, n114,
         n115, n116, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n135, n136, n137, n138,
         n139, n141, n142, n143, n144, n145, n146, n148, n149, n150, n151,
         n152, n153, n155, n156, n157, n158, n159, n160, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n193, n194, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n207, n208, n209, n211, n212, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n232, n233, n234, n235, n236, n238, n239,
         n240, n241, n242, n243, n245, n246, n247, n248, n249, n250, n252,
         n253, n254, n255, n256, n257, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n290, n291, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n304, n305, n306, n308, n309, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n327,
         n328, n329, n330, n332, n333, n334, n335, n336, n338, n339, n340,
         n341, n342, n344, n345, n346, n347, n348, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n370, n374, n375, n376, n377, n378, n379, n383,
         n384, n385, n585, n586, n587, n588, n589;
  assign n22 = A[61];
  assign n28 = A[60];
  assign n55 = A[56];
  assign n69 = A[54];
  assign n89 = A[51];
  assign n95 = A[50];
  assign n113 = A[47];
  assign n121 = A[46];
  assign n127 = A[45];
  assign n135 = A[44];
  assign n141 = A[43];
  assign n149 = A[42];
  assign n155 = A[41];
  assign n163 = A[40];
  assign n167 = A[39];
  assign n175 = A[38];
  assign n179 = A[37];
  assign n185 = A[36];
  assign n189 = A[35];
  assign n197 = A[34];
  assign n201 = A[33];
  assign n207 = A[32];
  assign n211 = A[31];
  assign n218 = A[30];
  assign n224 = A[29];
  assign n232 = A[28];
  assign n238 = A[27];
  assign n246 = A[26];
  assign n252 = A[25];
  assign n260 = A[24];
  assign n264 = A[23];
  assign n272 = A[22];
  assign n276 = A[21];
  assign n282 = A[20];
  assign n286 = A[19];
  assign n294 = A[18];
  assign n298 = A[17];
  assign n304 = A[16];
  assign n308 = A[15];
  assign n315 = A[14];
  assign n320 = A[13];
  assign n327 = A[12];
  assign n332 = A[11];
  assign n339 = A[10];
  assign n344 = A[9];
  assign n351 = A[8];
  assign n354 = A[7];
  assign n360 = A[6];
  assign n364 = A[5];
  assign n370 = A[4];
  assign n374 = A[3];
  assign n379 = A[2];
  assign n383 = A[1];

  CNR2X2 U359 ( .A(n312), .B(n357), .Z(n311) );
  CENX1 U454 ( .A(n105), .B(n104), .Z(SUM[49]) );
  CNR2XL U455 ( .A(n588), .B(n106), .Z(n105) );
  COR2XL U456 ( .A(n21), .B(n17), .Z(n585) );
  CNR2XL U457 ( .A(n588), .B(n19), .Z(n18) );
  CNR2XL U458 ( .A(n588), .B(n25), .Z(n24) );
  CNR2XL U459 ( .A(n588), .B(n44), .Z(n43) );
  CNR2XL U460 ( .A(n588), .B(n92), .Z(n91) );
  CNR2XL U461 ( .A(n588), .B(n13), .Z(n12) );
  CNR2XL U462 ( .A(n588), .B(n31), .Z(n30) );
  CNR2XL U463 ( .A(n588), .B(n98), .Z(n97) );
  CNR2X1 U464 ( .A(n3), .B(n221), .Z(n220) );
  CNR2X1 U465 ( .A(n3), .B(n263), .Z(n262) );
  CNR2X1 U466 ( .A(n3), .B(n285), .Z(n284) );
  CNR2X1 U467 ( .A(n3), .B(n297), .Z(n296) );
  CIVXL U468 ( .A(n311), .Z(n3) );
  CNR2XL U469 ( .A(n588), .B(n52), .Z(n51) );
  CNR2XL U470 ( .A(n588), .B(n72), .Z(n71) );
  CNR2XL U471 ( .A(n3), .B(n309), .Z(n306) );
  CND2XL U472 ( .A(n589), .B(n32), .Z(n31) );
  CND2XL U473 ( .A(n589), .B(n99), .Z(n98) );
  CNR2XL U474 ( .A(n588), .B(n110), .Z(n109) );
  CNR2XL U475 ( .A(n588), .B(n116), .Z(n115) );
  CND2XL U476 ( .A(n230), .B(n224), .Z(n223) );
  CND2XL U477 ( .A(n302), .B(n298), .Z(n297) );
  CND2XL U478 ( .A(n61), .B(n47), .Z(n46) );
  CND2XL U479 ( .A(n171), .B(n139), .Z(n138) );
  CNR2XL U480 ( .A(n146), .B(n142), .Z(n139) );
  CND2XL U481 ( .A(n171), .B(n159), .Z(n158) );
  CND2XL U482 ( .A(n171), .B(n167), .Z(n166) );
  CNIVX2 U483 ( .A(n8), .Z(n589) );
  CND2XL U484 ( .A(n171), .B(n125), .Z(n124) );
  CNR2XL U485 ( .A(n146), .B(n126), .Z(n125) );
  CNR2X1 U486 ( .A(n301), .B(n293), .Z(n290) );
  CND2XL U487 ( .A(n61), .B(n55), .Z(n54) );
  CEOXL U488 ( .A(n333), .B(n334), .Z(SUM[11]) );
  CNR2X2 U489 ( .A(n160), .B(n148), .Z(n145) );
  CNR2XL U490 ( .A(n194), .B(n184), .Z(n183) );
  CNR2XL U491 ( .A(n588), .B(n130), .Z(n129) );
  CNR2XL U492 ( .A(n146), .B(n132), .Z(n131) );
  CNR2XL U493 ( .A(n588), .B(n138), .Z(n137) );
  CNR2XL U494 ( .A(n588), .B(n144), .Z(n143) );
  CNR2XL U495 ( .A(n588), .B(n152), .Z(n151) );
  CNR2XL U496 ( .A(n160), .B(n156), .Z(n153) );
  CNR2XL U497 ( .A(n588), .B(n158), .Z(n157) );
  CNR2XL U498 ( .A(n588), .B(n166), .Z(n165) );
  CNR2XL U499 ( .A(n588), .B(n170), .Z(n169) );
  CNR2XL U500 ( .A(n588), .B(n182), .Z(n181) );
  CNR2XL U501 ( .A(n588), .B(n188), .Z(n187) );
  CNR2XL U502 ( .A(n588), .B(n194), .Z(n191) );
  CND2XL U503 ( .A(n205), .B(n201), .Z(n200) );
  CNR2XL U504 ( .A(n588), .B(n200), .Z(n199) );
  CNR2XL U505 ( .A(n588), .B(n204), .Z(n203) );
  CNR2XL U506 ( .A(n588), .B(n212), .Z(n209) );
  CND2XL U507 ( .A(n268), .B(n228), .Z(n227) );
  CNR2XL U508 ( .A(n243), .B(n229), .Z(n228) );
  CNR2XL U509 ( .A(n243), .B(n239), .Z(n236) );
  CND2XL U510 ( .A(n589), .B(n20), .Z(n19) );
  CND2XL U511 ( .A(n589), .B(n26), .Z(n25) );
  CND2XL U512 ( .A(n589), .B(n45), .Z(n44) );
  CND2XL U513 ( .A(n589), .B(n93), .Z(n92) );
  CND2XL U514 ( .A(n589), .B(n14), .Z(n13) );
  CNR2XL U515 ( .A(n588), .B(n38), .Z(n37) );
  CND2XL U516 ( .A(n589), .B(n39), .Z(n38) );
  CNR2XL U517 ( .A(n86), .B(n40), .Z(n39) );
  CND2XL U518 ( .A(n41), .B(n61), .Z(n40) );
  CNR2XL U519 ( .A(n588), .B(n58), .Z(n57) );
  CND2XL U520 ( .A(n589), .B(n59), .Z(n58) );
  CIVXL U521 ( .A(n28), .Z(n29) );
  CND2XL U522 ( .A(n290), .B(n286), .Z(n285) );
  CNR2X2 U523 ( .A(n100), .B(n88), .Z(n85) );
  CNR2X2 U524 ( .A(n257), .B(n245), .Z(n242) );
  CNR2XL U525 ( .A(n291), .B(n281), .Z(n280) );
  CNR2XL U526 ( .A(n114), .B(n108), .Z(n107) );
  CNR2XL U527 ( .A(n336), .B(n324), .Z(n323) );
  CNR2XL U528 ( .A(n348), .B(n345), .Z(n342) );
  CNR2XL U529 ( .A(n588), .B(n124), .Z(n123) );
  CND2XL U530 ( .A(n133), .B(n127), .Z(n126) );
  CNR2XL U531 ( .A(n588), .B(n178), .Z(n177) );
  CND2XL U532 ( .A(n183), .B(n179), .Z(n178) );
  CNR2XL U533 ( .A(n376), .B(n367), .Z(n366) );
  CEOXL U534 ( .A(n375), .B(n376), .Z(SUM[3]) );
  CNR2IXL U535 ( .B(n47), .A(n42), .Z(n41) );
  CND2XL U536 ( .A(n356), .B(n335), .Z(n334) );
  CIVX1 U537 ( .A(A[62]), .Z(n17) );
  CIVXL U538 ( .A(n22), .Z(n23) );
  CND2XL U539 ( .A(n280), .B(n276), .Z(n275) );
  CNR2X2 U540 ( .A(n348), .B(n338), .Z(n335) );
  CND2XL U541 ( .A(n368), .B(n364), .Z(n363) );
  CEOXL U542 ( .A(n1), .B(n384), .Z(SUM[1]) );
  CEOXL U543 ( .A(n586), .B(n379), .Z(SUM[2]) );
  CNR2XL U544 ( .A(n1), .B(n384), .Z(n586) );
  CEOXL U545 ( .A(n587), .B(n370), .Z(SUM[4]) );
  CNR2XL U546 ( .A(n376), .B(n375), .Z(n587) );
  CND2IXL U547 ( .B(n385), .A(n1), .Z(n10) );
  CENXL U548 ( .A(n151), .B(n150), .Z(SUM[42]) );
  CEOXL U549 ( .A(n316), .B(n317), .Z(SUM[14]) );
  CEOXL U550 ( .A(n321), .B(n322), .Z(SUM[13]) );
  CEOXL U551 ( .A(n328), .B(n329), .Z(SUM[12]) );
  CEOXL U552 ( .A(n340), .B(n341), .Z(SUM[10]) );
  CEOXL U553 ( .A(n345), .B(n346), .Z(SUM[9]) );
  CEOXL U554 ( .A(n352), .B(n353), .Z(SUM[8]) );
  CND2X1 U555 ( .A(n155), .B(n149), .Z(n148) );
  CNR2X1 U556 ( .A(n204), .B(n196), .Z(n193) );
  CND2X1 U557 ( .A(n201), .B(n197), .Z(n196) );
  CNR2X1 U558 ( .A(n588), .B(n84), .Z(n83) );
  CND2X1 U559 ( .A(n589), .B(n85), .Z(n84) );
  CNR2X1 U560 ( .A(n9), .B(n21), .Z(n20) );
  CNR2X1 U561 ( .A(n9), .B(n29), .Z(n26) );
  CNR2XL U562 ( .A(n86), .B(n46), .Z(n45) );
  CNR2XL U563 ( .A(n86), .B(n60), .Z(n59) );
  CNR2X1 U564 ( .A(n100), .B(n96), .Z(n93) );
  CNR2X1 U565 ( .A(n9), .B(n585), .Z(n14) );
  CND2X1 U566 ( .A(n589), .B(n113), .Z(n110) );
  CND2X1 U567 ( .A(n171), .B(n131), .Z(n130) );
  CND2XL U568 ( .A(n171), .B(n145), .Z(n144) );
  CND2XL U569 ( .A(n171), .B(n153), .Z(n152) );
  CND2XL U570 ( .A(n193), .B(n189), .Z(n188) );
  CNR2X1 U571 ( .A(n3), .B(n227), .Z(n226) );
  CNR2X1 U572 ( .A(n3), .B(n235), .Z(n234) );
  CND2XL U573 ( .A(n268), .B(n236), .Z(n235) );
  CNR2X1 U574 ( .A(n3), .B(n241), .Z(n240) );
  CND2XL U575 ( .A(n268), .B(n242), .Z(n241) );
  CNR2X1 U576 ( .A(n3), .B(n249), .Z(n248) );
  CND2XL U577 ( .A(n268), .B(n250), .Z(n249) );
  CNR2X1 U578 ( .A(n257), .B(n253), .Z(n250) );
  CNR2X1 U579 ( .A(n3), .B(n255), .Z(n254) );
  CND2XL U580 ( .A(n268), .B(n256), .Z(n255) );
  CNR2X1 U581 ( .A(n3), .B(n279), .Z(n278) );
  CNR2X1 U582 ( .A(n3), .B(n291), .Z(n288) );
  CND2X1 U583 ( .A(n141), .B(n135), .Z(n132) );
  CND2X1 U584 ( .A(n163), .B(n167), .Z(n160) );
  CNR2X1 U585 ( .A(n170), .B(n118), .Z(n8) );
  CND2X1 U586 ( .A(n145), .B(n119), .Z(n118) );
  CNR2X1 U587 ( .A(n132), .B(n120), .Z(n119) );
  CND2X1 U588 ( .A(n89), .B(n95), .Z(n88) );
  CND2X1 U589 ( .A(n252), .B(n246), .Z(n245) );
  CNR2X1 U590 ( .A(n56), .B(n50), .Z(n47) );
  CND2X1 U591 ( .A(n298), .B(n294), .Z(n293) );
  CND2XL U592 ( .A(n589), .B(n107), .Z(n106) );
  CND2XL U593 ( .A(n589), .B(n53), .Z(n52) );
  CNR2XL U594 ( .A(n86), .B(n54), .Z(n53) );
  CND2XL U595 ( .A(n589), .B(n73), .Z(n72) );
  CNR2XL U596 ( .A(n86), .B(n74), .Z(n73) );
  CND2XL U597 ( .A(n268), .B(n222), .Z(n221) );
  CNR2X1 U598 ( .A(n243), .B(n223), .Z(n222) );
  CND2XL U599 ( .A(n268), .B(n264), .Z(n263) );
  CNR2XL U600 ( .A(n3), .B(n267), .Z(n266) );
  CNR2XL U601 ( .A(n3), .B(n301), .Z(n300) );
  CND2X1 U602 ( .A(n173), .B(n193), .Z(n170) );
  CNR2X1 U603 ( .A(n184), .B(n174), .Z(n173) );
  CND2X1 U604 ( .A(n179), .B(n175), .Z(n174) );
  CND2X1 U605 ( .A(n33), .B(n85), .Z(n9) );
  CNR2X1 U606 ( .A(n60), .B(n34), .Z(n33) );
  CND2X1 U607 ( .A(n47), .B(n35), .Z(n34) );
  CNR2X1 U608 ( .A(n36), .B(n42), .Z(n35) );
  CNR2X1 U609 ( .A(n229), .B(n217), .Z(n216) );
  CND2X1 U610 ( .A(n224), .B(n218), .Z(n217) );
  CND2X1 U611 ( .A(n238), .B(n232), .Z(n229) );
  CND2X1 U612 ( .A(n207), .B(n211), .Z(n204) );
  CND2X1 U613 ( .A(n75), .B(n63), .Z(n60) );
  CNR2X1 U614 ( .A(n70), .B(n64), .Z(n63) );
  CND2X1 U615 ( .A(n260), .B(n264), .Z(n257) );
  CND2X1 U616 ( .A(n103), .B(n113), .Z(n100) );
  CNR2X1 U617 ( .A(n108), .B(n104), .Z(n103) );
  CND2X1 U618 ( .A(n189), .B(n185), .Z(n184) );
  CND2X1 U619 ( .A(n28), .B(n22), .Z(n21) );
  CNIVX4 U620 ( .A(n6), .Z(n588) );
  CND2X1 U621 ( .A(n311), .B(n214), .Z(n6) );
  CNR2X1 U622 ( .A(n267), .B(n215), .Z(n214) );
  CND2X1 U623 ( .A(n242), .B(n216), .Z(n215) );
  CND2XL U624 ( .A(n356), .B(n342), .Z(n341) );
  CND2XL U625 ( .A(n356), .B(n347), .Z(n346) );
  CND2XL U626 ( .A(n323), .B(n356), .Z(n322) );
  CND2XL U627 ( .A(n330), .B(n356), .Z(n329) );
  CNR2XL U628 ( .A(n336), .B(n333), .Z(n330) );
  CND2X1 U629 ( .A(n127), .B(n121), .Z(n120) );
  CND2X1 U630 ( .A(n335), .B(n313), .Z(n312) );
  CNR2X1 U631 ( .A(n324), .B(n314), .Z(n313) );
  CND2X1 U632 ( .A(n320), .B(n315), .Z(n314) );
  CND2X1 U633 ( .A(n344), .B(n339), .Z(n338) );
  CNR2X1 U634 ( .A(n82), .B(n78), .Z(n75) );
  CNR2XL U635 ( .A(n588), .B(n66), .Z(n65) );
  CND2XL U636 ( .A(n589), .B(n67), .Z(n66) );
  CNR2XL U637 ( .A(n86), .B(n68), .Z(n67) );
  CND2XL U638 ( .A(n75), .B(n69), .Z(n68) );
  CNR2XL U639 ( .A(n588), .B(n80), .Z(n79) );
  CND2XL U640 ( .A(n589), .B(n81), .Z(n80) );
  CNR2XL U641 ( .A(n86), .B(n82), .Z(n81) );
  CNR2XL U642 ( .A(n3), .B(n275), .Z(n274) );
  CNR2X1 U643 ( .A(n363), .B(n376), .Z(n362) );
  CNR2X1 U644 ( .A(n378), .B(n1), .Z(n377) );
  CND2X1 U645 ( .A(n383), .B(n379), .Z(n378) );
  CND2X1 U646 ( .A(n290), .B(n270), .Z(n267) );
  CNR2X1 U647 ( .A(n281), .B(n271), .Z(n270) );
  CND2X1 U648 ( .A(n276), .B(n272), .Z(n271) );
  CND2X1 U649 ( .A(n332), .B(n327), .Z(n324) );
  CND2X1 U650 ( .A(n308), .B(n304), .Z(n301) );
  CND2X1 U651 ( .A(n374), .B(n370), .Z(n367) );
  CND2X1 U652 ( .A(n354), .B(n351), .Z(n348) );
  CND2X1 U653 ( .A(n286), .B(n282), .Z(n281) );
  CND2X1 U654 ( .A(n358), .B(n377), .Z(n357) );
  CNR2X1 U655 ( .A(n367), .B(n359), .Z(n358) );
  CND2X1 U656 ( .A(n364), .B(n360), .Z(n359) );
  CND2XL U657 ( .A(n356), .B(n354), .Z(n353) );
  CND2XL U658 ( .A(n318), .B(n356), .Z(n317) );
  CNR2XL U659 ( .A(n336), .B(n319), .Z(n318) );
  CND2XL U660 ( .A(n325), .B(n320), .Z(n319) );
  CND2X1 U661 ( .A(B[0]), .B(A[0]), .Z(n1) );
  CNR2XL U662 ( .A(B[0]), .B(A[0]), .Z(n385) );
  CENX1 U663 ( .A(n115), .B(n114), .Z(SUM[47]) );
  CENX1 U664 ( .A(n165), .B(n164), .Z(SUM[40]) );
  CENX1 U665 ( .A(n177), .B(n176), .Z(SUM[38]) );
  CENX1 U666 ( .A(n169), .B(n168), .Z(SUM[39]) );
  CENX1 U667 ( .A(n181), .B(n180), .Z(SUM[37]) );
  CENX1 U668 ( .A(n191), .B(n190), .Z(SUM[35]) );
  CENX1 U669 ( .A(n199), .B(n198), .Z(SUM[34]) );
  CENX1 U670 ( .A(n203), .B(n202), .Z(SUM[33]) );
  CENX1 U671 ( .A(n209), .B(n208), .Z(SUM[32]) );
  CEOXL U672 ( .A(n212), .B(n588), .Z(SUM[31]) );
  CENX1 U673 ( .A(n220), .B(n219), .Z(SUM[30]) );
  CENX1 U674 ( .A(n226), .B(n225), .Z(SUM[29]) );
  CENX1 U675 ( .A(n234), .B(n233), .Z(SUM[28]) );
  CENX1 U676 ( .A(n240), .B(n239), .Z(SUM[27]) );
  CENX1 U677 ( .A(n248), .B(n247), .Z(SUM[26]) );
  CENX1 U678 ( .A(n12), .B(n11), .Z(SUM[63]) );
  CENXL U679 ( .A(n37), .B(n36), .Z(SUM[59]) );
  CENXL U680 ( .A(n57), .B(n56), .Z(SUM[56]) );
  CENX1 U681 ( .A(n18), .B(n17), .Z(SUM[62]) );
  CENX1 U682 ( .A(n24), .B(n23), .Z(SUM[61]) );
  CENX1 U683 ( .A(n30), .B(n29), .Z(SUM[60]) );
  CENX1 U684 ( .A(n43), .B(n42), .Z(SUM[58]) );
  CENX1 U685 ( .A(n51), .B(n50), .Z(SUM[57]) );
  CENX1 U686 ( .A(n65), .B(n64), .Z(SUM[55]) );
  CENX1 U687 ( .A(n71), .B(n70), .Z(SUM[54]) );
  CENX1 U688 ( .A(n79), .B(n78), .Z(SUM[53]) );
  CENX1 U689 ( .A(n83), .B(n82), .Z(SUM[52]) );
  CENX1 U690 ( .A(n91), .B(n90), .Z(SUM[51]) );
  CENX1 U691 ( .A(n97), .B(n96), .Z(SUM[50]) );
  CENX1 U692 ( .A(n143), .B(n142), .Z(SUM[43]) );
  CENX1 U693 ( .A(n157), .B(n156), .Z(SUM[41]) );
  CENX1 U694 ( .A(n123), .B(n122), .Z(SUM[46]) );
  CENX1 U695 ( .A(n129), .B(n128), .Z(SUM[45]) );
  CENX1 U696 ( .A(n137), .B(n136), .Z(SUM[44]) );
  CENX1 U697 ( .A(n187), .B(n186), .Z(SUM[36]) );
  CENX1 U698 ( .A(n109), .B(n108), .Z(SUM[48]) );
  CENX1 U699 ( .A(n254), .B(n253), .Z(SUM[25]) );
  CENX1 U700 ( .A(n262), .B(n261), .Z(SUM[24]) );
  CENX1 U701 ( .A(n266), .B(n265), .Z(SUM[23]) );
  CENX1 U702 ( .A(n274), .B(n273), .Z(SUM[22]) );
  CENX1 U703 ( .A(n278), .B(n277), .Z(SUM[21]) );
  CENX1 U704 ( .A(n284), .B(n283), .Z(SUM[20]) );
  CENX1 U705 ( .A(n288), .B(n287), .Z(SUM[19]) );
  CENX1 U706 ( .A(n296), .B(n295), .Z(SUM[18]) );
  CENX1 U707 ( .A(n300), .B(n299), .Z(SUM[17]) );
  CENX1 U708 ( .A(n306), .B(n305), .Z(SUM[16]) );
  CEOXL U709 ( .A(n309), .B(n3), .Z(SUM[15]) );
  CENX1 U710 ( .A(n356), .B(n355), .Z(SUM[7]) );
  CENX1 U711 ( .A(n362), .B(n361), .Z(SUM[6]) );
  CENX1 U712 ( .A(n366), .B(n365), .Z(SUM[5]) );
  CIVX2 U713 ( .A(n100), .Z(n99) );
  CIVX2 U714 ( .A(n95), .Z(n96) );
  CIVX2 U715 ( .A(n89), .Z(n90) );
  CIVX2 U716 ( .A(n85), .Z(n86) );
  CIVX2 U717 ( .A(A[52]), .Z(n82) );
  CIVX2 U718 ( .A(A[53]), .Z(n78) );
  CIVX2 U719 ( .A(n75), .Z(n74) );
  CIVX2 U720 ( .A(n69), .Z(n70) );
  CIVX2 U721 ( .A(A[55]), .Z(n64) );
  CIVX2 U722 ( .A(n60), .Z(n61) );
  CIVX2 U723 ( .A(n55), .Z(n56) );
  CIVX2 U724 ( .A(A[57]), .Z(n50) );
  CIVX2 U725 ( .A(A[58]), .Z(n42) );
  CIVX2 U726 ( .A(n383), .Z(n384) );
  CIVX2 U727 ( .A(n377), .Z(n376) );
  CIVX2 U728 ( .A(n374), .Z(n375) );
  CIVX2 U729 ( .A(n367), .Z(n368) );
  CIVX2 U730 ( .A(n364), .Z(n365) );
  CIVX2 U731 ( .A(n360), .Z(n361) );
  CIVX2 U732 ( .A(A[59]), .Z(n36) );
  CIVX2 U733 ( .A(n357), .Z(n356) );
  CIVX2 U734 ( .A(n354), .Z(n355) );
  CIVX2 U735 ( .A(n351), .Z(n352) );
  CIVX2 U736 ( .A(n348), .Z(n347) );
  CIVX2 U737 ( .A(n344), .Z(n345) );
  CIVX2 U738 ( .A(n339), .Z(n340) );
  CIVX2 U739 ( .A(n335), .Z(n336) );
  CIVX2 U740 ( .A(n332), .Z(n333) );
  CIVX2 U741 ( .A(n327), .Z(n328) );
  CIVX2 U742 ( .A(n324), .Z(n325) );
  CIVX2 U743 ( .A(n320), .Z(n321) );
  CIVX2 U744 ( .A(n9), .Z(n32) );
  CIVX2 U745 ( .A(n315), .Z(n316) );
  CIVX2 U746 ( .A(n308), .Z(n309) );
  CIVX2 U747 ( .A(n304), .Z(n305) );
  CIVX2 U748 ( .A(n301), .Z(n302) );
  CIVX2 U749 ( .A(n298), .Z(n299) );
  CIVX2 U750 ( .A(n294), .Z(n295) );
  CIVX2 U751 ( .A(n290), .Z(n291) );
  CIVX2 U752 ( .A(n286), .Z(n287) );
  CIVX2 U753 ( .A(n282), .Z(n283) );
  CIVX2 U754 ( .A(n280), .Z(n279) );
  CIVX2 U755 ( .A(n276), .Z(n277) );
  CIVX2 U756 ( .A(n272), .Z(n273) );
  CIVX2 U757 ( .A(n267), .Z(n268) );
  CIVX2 U758 ( .A(n264), .Z(n265) );
  CIVX2 U759 ( .A(n260), .Z(n261) );
  CIVX2 U760 ( .A(n257), .Z(n256) );
  CIVX2 U761 ( .A(n252), .Z(n253) );
  CIVX2 U762 ( .A(n246), .Z(n247) );
  CIVX2 U763 ( .A(n242), .Z(n243) );
  CIVX2 U764 ( .A(n238), .Z(n239) );
  CIVX2 U765 ( .A(n232), .Z(n233) );
  CIVX2 U766 ( .A(n229), .Z(n230) );
  CIVX2 U767 ( .A(n224), .Z(n225) );
  CIVX2 U768 ( .A(n218), .Z(n219) );
  CIVX2 U769 ( .A(n211), .Z(n212) );
  CIVX2 U770 ( .A(n207), .Z(n208) );
  CIVX2 U771 ( .A(n204), .Z(n205) );
  CIVX2 U772 ( .A(n201), .Z(n202) );
  CIVX2 U773 ( .A(n197), .Z(n198) );
  CIVX2 U774 ( .A(n193), .Z(n194) );
  CIVX2 U775 ( .A(n189), .Z(n190) );
  CIVX2 U776 ( .A(n185), .Z(n186) );
  CIVX2 U777 ( .A(n183), .Z(n182) );
  CIVX2 U778 ( .A(n179), .Z(n180) );
  CIVX2 U779 ( .A(n175), .Z(n176) );
  CIVX2 U780 ( .A(n170), .Z(n171) );
  CIVX2 U781 ( .A(n167), .Z(n168) );
  CIVX2 U782 ( .A(n163), .Z(n164) );
  CIVX2 U783 ( .A(n160), .Z(n159) );
  CIVX2 U784 ( .A(n155), .Z(n156) );
  CIVX2 U785 ( .A(n149), .Z(n150) );
  CIVX2 U786 ( .A(n145), .Z(n146) );
  CIVX2 U787 ( .A(n141), .Z(n142) );
  CIVX2 U788 ( .A(n135), .Z(n136) );
  CIVX2 U789 ( .A(n132), .Z(n133) );
  CIVX2 U790 ( .A(n127), .Z(n128) );
  CIVX2 U791 ( .A(n121), .Z(n122) );
  CIVX2 U792 ( .A(n589), .Z(n116) );
  CIVX2 U793 ( .A(n113), .Z(n114) );
  CIVX2 U794 ( .A(A[63]), .Z(n11) );
  CIVX2 U795 ( .A(A[48]), .Z(n108) );
  CIVX2 U796 ( .A(A[49]), .Z(n104) );
  CIVX2 U797 ( .A(n10), .Z(SUM[0]) );
endmodule


module sfilt_DW01_add_6 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n6, n7, n9, n11, n12, n13, n14, n15, n16, n17, n19, n21,
         n22, n23, n24, n25, n26, n28, n29, n30, n36, n37, n38, n39, n40, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n80, n95, n96, n97, n98, n99, n100, n102,
         n115, n116, n117, n118, n122, n124, n125, n126, n127, n128, n129,
         n130, n131, n134, n135, n136, n137, n138, n139, n141, n144, n145,
         n146, n147, n148, n150, n151, n152, n153, n154, n155, n160, n162,
         n163, n164, n165, n166, n167, n168, n169, n172, n173, n174, n175,
         n176, n177, n179, n191, n209, n210, n211, n218, n219, n220, n221,
         n222, n232, n233, n234, n235, n236, n237, n241, n242, n243, n244,
         n247, n251, n252, n253, n254, n256, n257, n258, n259, n260, n262,
         n263, n270, n271, n272, n277, n278, n279, n280, n286, n287, n288,
         n289, n290, n291, n297, n298, n299, n300, n301, n302, n305, n306,
         n307, n308, n313, n314, n316, n318, n319, n320, n321, n322, n323,
         n325, n328, n329, n330, n331, n332, n338, n339, n340, n341, n343,
         n345, n346, n347, n348, n349, n350, n351, n353, n354, n355, n356,
         n357, n358, n362, n364, n365, n366, n367, n368, n369, n373, n374,
         n375, n376, n377, n378, n380, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n397, n398, n399, n400, n402,
         n405, n406, n407, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n422, n424, n425, n426, n427, n429, n432,
         n433, n434, n435, n437, n439, n440, n441, n442, n443, n444, n445,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n460, n462, n463, n464, n465, n467, n470, n471, n472, n473,
         n475, n477, n478, n480, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n497, n499, n500, n502,
         n504, n505, n506, n508, n510, n511, n512, n513, n515, n517, n518,
         n520, n522, n523, n524, n526, n528, n529, n530, n531, n532, n534,
         n536, n537, n538, n539, n542, n543, n544, n546, n548, n549, n550,
         n551, n552, n558, n559, n560, n561, n570, n571, n572, n573, n574,
         n576, n578, n580, n581, n583, n585, n586, n587, n588, n589, n590,
         n591, n593, n595, n596, n597, n599, n602, n603, n610, net16249,
         net17506, net17505, net18014, net18013, net18589, net18840, net18843,
         net18964, n93, n94, n91, n90, n89, n88, n87, n86, n85, n84, n83, n82,
         n81, n8, n79, n553, n103, n101, net17940, n577, n310, n296, n295,
         n294, n293, n292, n224, net18512, n569, n250, n245, n240, n231, n229,
         n228, n227, n226, n225, net18513, n281, n276, n275, n274, n269, n267,
         n266, n261, n566, n565, n213, n212, n208, n207, n206, n204, n203,
         n202, n201, n200, n20, n198, n268, n158, n556, n555, n5, n161, n159,
         n123, n114, n111, n110, n109, n108, n107, n106, n105, n104, n10, n564,
         n199, n195, n194, n193, n192, n190, n189, n188, n186, n185, n184,
         n183, n182, n18, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883;

  CND2X2 U8 ( .A(n552), .B(n72), .Z(n7) );
  CNR2X2 U10 ( .A(A[63]), .B(B[63]), .Z(n71) );
  COND1X1 U41 ( .A(n96), .B(net18014), .C(n97), .Z(n95) );
  CANR1X1 U43 ( .A(n819), .B(n850), .C(n99), .Z(n97) );
  CND2X2 U72 ( .A(n122), .B(n138), .Z(n6) );
  CNR2X2 U78 ( .A(A[58]), .B(B[58]), .Z(n124) );
  COND1X1 U81 ( .A(n127), .B(n852), .C(n128), .Z(n126) );
  CANR1X1 U83 ( .A(n129), .B(n850), .C(n130), .Z(n128) );
  COND1X1 U93 ( .A(n136), .B(n852), .C(n137), .Z(n135) );
  CNR2X2 U100 ( .A(n151), .B(n144), .Z(n138) );
  COND1X1 U117 ( .A(n154), .B(n852), .C(n155), .Z(n153) );
  CNR2X2 U128 ( .A(A[54]), .B(B[54]), .Z(n162) );
  CNR2X2 U202 ( .A(A[48]), .B(B[48]), .Z(n218) );
  CND2X2 U209 ( .A(A[47]), .B(B[47]), .Z(n222) );
  CNR2X2 U294 ( .A(A[40]), .B(B[40]), .Z(n286) );
  CNR2X2 U311 ( .A(A[38]), .B(B[38]), .Z(n297) );
  CND2X2 U331 ( .A(n580), .B(n848), .Z(n313) );
  CND2X2 U359 ( .A(n824), .B(n581), .Z(n331) );
  CANR1X1 U428 ( .A(n400), .B(n387), .C(n388), .Z(n386) );
  CNR2X2 U443 ( .A(A[27]), .B(B[27]), .Z(n394) );
  CNR2X2 U38 ( .A(A[61]), .B(B[61]), .Z(n93) );
  CANR1X1 U19 ( .A(n103), .B(n80), .C(n81), .Z(n79) );
  CNR2X2 U24 ( .A(A[62]), .B(B[62]), .Z(n82) );
  COND1X1 U21 ( .A(n94), .B(n82), .C(n83), .Z(n81) );
  CANR1X1 U33 ( .A(n91), .B(n103), .C(n821), .Z(n90) );
  CANR1X1 U29 ( .A(n820), .B(n850), .C(n88), .Z(n86) );
  COND1X1 U27 ( .A(n85), .B(net18013), .C(n86), .Z(n84) );
  CNR2X2 U212 ( .A(net17940), .B(n260), .Z(n224) );
  COND1X1 U308 ( .A(n305), .B(n297), .C(n298), .Z(n296) );
  CNR2X2 U242 ( .A(n257), .B(net18589), .Z(n244) );
  CNR2X2 U216 ( .A(n237), .B(n857), .Z(n228) );
  CNR2X2 U290 ( .A(n286), .B(n289), .Z(n280) );
  CNR2X2 U266 ( .A(n275), .B(net18513), .Z(n266) );
  CNR2X2 U198 ( .A(n221), .B(n218), .Z(n212) );
  COND1X1 U181 ( .A(n203), .B(net18013), .C(n204), .Z(n202) );
  CND2X2 U122 ( .A(n160), .B(n176), .Z(n158) );
  CNR2X2 U64 ( .A(A[59]), .B(B[59]), .Z(n111) );
  CNR2X2 U52 ( .A(A[60]), .B(B[60]), .Z(n104) );
  CND2X2 U172 ( .A(n198), .B(n212), .Z(n192) );
  CNR2X2 U150 ( .A(n189), .B(n182), .Z(n176) );
  CNR2X2 U154 ( .A(A[52]), .B(B[52]), .Z(n182) );
  CND2XL U683 ( .A(n553), .B(n83), .Z(n8) );
  CND2X1 U684 ( .A(A[62]), .B(B[62]), .Z(n83) );
  COND1X2 U685 ( .A(n190), .B(n182), .C(n183), .Z(n177) );
  CND2X2 U686 ( .A(A[51]), .B(B[51]), .Z(n190) );
  CIVX2 U687 ( .A(n384), .Z(n383) );
  CIVXL U688 ( .A(n443), .Z(n595) );
  CNR2XL U689 ( .A(A[20]), .B(B[20]), .Z(n443) );
  CND2XL U690 ( .A(n595), .B(n444), .Z(n50) );
  CIVXL U691 ( .A(n499), .Z(n497) );
  CIVX1 U692 ( .A(n506), .Z(n505) );
  CIVX1 U693 ( .A(n464), .Z(n599) );
  CNR2X2 U694 ( .A(A[12]), .B(B[12]), .Z(n490) );
  CENXL U695 ( .A(n412), .B(n45), .Z(SUM[25]) );
  CNR2X1 U696 ( .A(n419), .B(n416), .Z(n414) );
  CIVXL U697 ( .A(n416), .Z(n591) );
  CANR1XL U698 ( .A(n307), .B(n346), .C(n834), .Z(n306) );
  CANR1X1 U699 ( .A(n329), .B(n346), .C(n330), .Z(n328) );
  CANR1X1 U700 ( .A(n320), .B(n346), .C(n321), .Z(n319) );
  CNIVX1 U701 ( .A(n305), .Z(n814) );
  COND1X1 U702 ( .A(n411), .B(n405), .C(n406), .Z(n400) );
  CND2XL U703 ( .A(n591), .B(n417), .Z(n46) );
  CIVX1 U704 ( .A(n484), .Z(n861) );
  CIVXL U705 ( .A(n380), .Z(n815) );
  CIVXL U706 ( .A(n380), .Z(n816) );
  COND1XL U707 ( .A(n278), .B(n291), .C(n279), .Z(n277) );
  CIVX1 U708 ( .A(n347), .Z(n346) );
  CIVXL U709 ( .A(n332), .Z(n330) );
  CIVX1 U710 ( .A(n818), .Z(n263) );
  COND1XL U711 ( .A(n313), .B(n332), .C(n314), .Z(n817) );
  CANR1X1 U712 ( .A(n281), .B(n266), .C(n267), .Z(n818) );
  CANR1X1 U713 ( .A(n281), .B(n266), .C(n267), .Z(n261) );
  CNR2XL U714 ( .A(n100), .B(n6), .Z(n819) );
  CNR2XL U715 ( .A(n100), .B(n6), .Z(n98) );
  CIVX1 U716 ( .A(n141), .Z(n837) );
  COND1X1 U717 ( .A(n131), .B(n141), .C(n134), .Z(n130) );
  COND1X2 U718 ( .A(n114), .B(n104), .C(n105), .Z(n103) );
  CIVX2 U719 ( .A(n290), .Z(n854) );
  CNR2IX1 U720 ( .B(n176), .A(n169), .Z(n167) );
  CNR2X2 U721 ( .A(A[53]), .B(B[53]), .Z(n169) );
  CND2X1 U722 ( .A(n102), .B(n80), .Z(n78) );
  CNR2XL U723 ( .A(n6), .B(n89), .Z(n820) );
  CNR2XL U724 ( .A(n6), .B(n89), .Z(n87) );
  CIVX1 U725 ( .A(n839), .Z(n141) );
  CIVX1 U726 ( .A(n93), .Z(n91) );
  CNR2X1 U727 ( .A(n93), .B(n82), .Z(n80) );
  CIVXL U728 ( .A(n413), .Z(n412) );
  CIVDXL U729 ( .A(n200), .Z0(n565) );
  CIVX1 U730 ( .A(n212), .Z(n210) );
  CIVXL U731 ( .A(n82), .Z(n553) );
  CND2X2 U732 ( .A(A[39]), .B(B[39]), .Z(n290) );
  CAN2XL U733 ( .A(A[61]), .B(B[61]), .Z(n821) );
  CIVXL U734 ( .A(n104), .Z(n555) );
  CIVX1 U735 ( .A(n318), .Z(n316) );
  COND1X2 U736 ( .A(n208), .B(n200), .C(n201), .Z(n199) );
  CIVX1 U737 ( .A(n4), .Z(n154) );
  CND2X1 U738 ( .A(A[52]), .B(B[52]), .Z(n183) );
  CND2X2 U739 ( .A(A[46]), .B(B[46]), .Z(n231) );
  CENXL U740 ( .A(n95), .B(n9), .Z(SUM[61]) );
  CIVX1 U741 ( .A(n245), .Z(n247) );
  COND1X2 U742 ( .A(n258), .B(n250), .C(n251), .Z(n245) );
  CND2X2 U743 ( .A(A[45]), .B(B[45]), .Z(n240) );
  CANR1XL U744 ( .A(n195), .B(n167), .C(n168), .Z(n166) );
  COND1X1 U745 ( .A(n313), .B(n332), .C(n314), .Z(n308) );
  CND2X1 U746 ( .A(A[49]), .B(B[49]), .Z(n208) );
  COND1XL U747 ( .A(n169), .B(n179), .C(n172), .Z(n168) );
  CND2X1 U748 ( .A(A[59]), .B(B[59]), .Z(n114) );
  CND2X1 U749 ( .A(n102), .B(n91), .Z(n89) );
  CANR1X1 U750 ( .A(n485), .B(n493), .C(n486), .Z(n484) );
  CANR1X1 U751 ( .A(n870), .B(n442), .C(n437), .Z(n435) );
  COND1X1 U752 ( .A(n454), .B(n458), .C(n455), .Z(n453) );
  CND2X1 U753 ( .A(A[36]), .B(B[36]), .Z(n318) );
  CIVXL U754 ( .A(B[36]), .Z(n849) );
  CANR1XL U755 ( .A(n572), .B(n263), .C(n256), .Z(n254) );
  CND2XL U756 ( .A(n555), .B(n105), .Z(n10) );
  CND2X1 U757 ( .A(n565), .B(n201), .Z(n20) );
  COND1XL U758 ( .A(n165), .B(net18014), .C(n166), .Z(n164) );
  CND2XL U759 ( .A(n558), .B(n134), .Z(n13) );
  CNIVX1 U760 ( .A(n221), .Z(n822) );
  COR2X1 U761 ( .A(A[31]), .B(B[31]), .Z(n823) );
  COR2X1 U762 ( .A(A[33]), .B(B[33]), .Z(n824) );
  CENXL U763 ( .A(n418), .B(n46), .Z(SUM[24]) );
  CENXL U764 ( .A(n383), .B(n825), .Z(SUM[29]) );
  CAN2XL U765 ( .A(n586), .B(n816), .Z(n825) );
  CENXL U766 ( .A(n826), .B(n391), .Z(SUM[28]) );
  CAN2XL U767 ( .A(n587), .B(n390), .Z(n826) );
  CENXL U768 ( .A(n827), .B(n407), .Z(SUM[26]) );
  CAN2XL U769 ( .A(n589), .B(n406), .Z(n827) );
  CENXL U770 ( .A(n828), .B(n398), .Z(SUM[27]) );
  CAN2XL U771 ( .A(n588), .B(n397), .Z(n828) );
  CANR1X1 U772 ( .A(n520), .B(n875), .C(n515), .Z(n513) );
  CND2X1 U773 ( .A(n593), .B(n871), .Z(n419) );
  CIVXL U774 ( .A(n484), .Z(n483) );
  CANR1X1 U775 ( .A(n480), .B(n873), .C(n475), .Z(n473) );
  CIVXL U776 ( .A(n477), .Z(n475) );
  CIVXL U777 ( .A(n482), .Z(n480) );
  CIVXL U778 ( .A(n493), .Z(n492) );
  CENXL U779 ( .A(n376), .B(n40), .Z(SUM[30]) );
  CENXL U780 ( .A(n356), .B(n38), .Z(SUM[32]) );
  CENXL U781 ( .A(n365), .B(n39), .Z(SUM[31]) );
  CANR1XL U782 ( .A(n300), .B(n346), .C(n301), .Z(n299) );
  CENXL U783 ( .A(n291), .B(n829), .Z(SUM[39]) );
  CAN2XL U784 ( .A(n576), .B(n290), .Z(n829) );
  CIVX1 U785 ( .A(n375), .Z(n373) );
  CNR2XL U786 ( .A(A[19]), .B(B[19]), .Z(n448) );
  CIVXL U787 ( .A(n405), .Z(n589) );
  CIVX1 U788 ( .A(n374), .Z(n585) );
  CENXL U789 ( .A(n830), .B(n328), .Z(SUM[35]) );
  CAN2XL U790 ( .A(n580), .B(n323), .Z(n830) );
  CENXL U791 ( .A(n831), .B(n319), .Z(SUM[36]) );
  CAN2XL U792 ( .A(n848), .B(n318), .Z(n831) );
  CENXL U793 ( .A(n832), .B(n306), .Z(SUM[37]) );
  CAN2XL U794 ( .A(n578), .B(n814), .Z(n832) );
  CENXL U795 ( .A(n277), .B(n29), .Z(SUM[41]) );
  CENXL U796 ( .A(n252), .B(n26), .Z(SUM[44]) );
  COND1XL U797 ( .A(n253), .B(n291), .C(n254), .Z(n252) );
  CENXL U798 ( .A(n833), .B(n299), .Z(SUM[38]) );
  CAN2XL U799 ( .A(n577), .B(n298), .Z(n833) );
  CNR2X1 U800 ( .A(A[34]), .B(B[34]), .Z(n339) );
  CIVX1 U801 ( .A(n297), .Z(n577) );
  CENXL U802 ( .A(n164), .B(n16), .Z(SUM[54]) );
  CIVXL U803 ( .A(n310), .Z(n834) );
  CENXL U804 ( .A(n153), .B(n15), .Z(SUM[55]) );
  COND1XL U805 ( .A(n260), .B(n291), .C(net18840), .Z(n259) );
  CANR1XL U806 ( .A(n109), .B(n3), .C(n110), .Z(n108) );
  COND1XL U807 ( .A(n107), .B(net18013), .C(n108), .Z(n106) );
  CIVXL U808 ( .A(n389), .Z(n587) );
  CNR2X1 U809 ( .A(n389), .B(n394), .Z(n387) );
  CNIVXL U810 ( .A(n176), .Z(n835) );
  CNR2X1 U811 ( .A(n6), .B(n78), .Z(n76) );
  CIVXL U812 ( .A(n6), .Z(n118) );
  COR2XL U813 ( .A(B[58]), .B(A[58]), .Z(n836) );
  CND2XL U814 ( .A(n883), .B(n882), .Z(SUM[49]) );
  CIVX1 U815 ( .A(n189), .Z(n564) );
  COND1X1 U816 ( .A(n134), .B(n124), .C(n125), .Z(n858) );
  CANR1X1 U817 ( .A(n564), .B(n195), .C(n188), .Z(n186) );
  COND1X1 U818 ( .A(n152), .B(n144), .C(n145), .Z(n139) );
  CIVXL U819 ( .A(n195), .Z(n838) );
  CIVXL U820 ( .A(n257), .Z(n572) );
  COND1X1 U821 ( .A(n134), .B(n124), .C(n125), .Z(n123) );
  COND1X1 U822 ( .A(n152), .B(n144), .C(n145), .Z(n839) );
  CND2XL U823 ( .A(n4), .B(n98), .Z(n96) );
  CNR2XL U824 ( .A(n131), .B(n124), .Z(n840) );
  CANR1XL U825 ( .A(n560), .B(n3), .C(n150), .Z(n148) );
  CIVX1 U826 ( .A(n275), .Z(n574) );
  COND1XL U827 ( .A(n293), .B(n846), .C(n294), .Z(n841) );
  COND1X1 U828 ( .A(n347), .B(n293), .C(n294), .Z(n842) );
  COND1XL U829 ( .A(n347), .B(n293), .C(n294), .Z(n845) );
  CDLY1XL U830 ( .A(net18512), .Z(n843) );
  COND1XL U831 ( .A(n293), .B(n846), .C(n294), .Z(n292) );
  COND1X1 U832 ( .A(n347), .B(n293), .C(n294), .Z(n844) );
  CND2X2 U833 ( .A(A[55]), .B(B[55]), .Z(n152) );
  COND1X1 U834 ( .A(n416), .B(n420), .C(n417), .Z(n415) );
  CANR1XL U835 ( .A(n348), .B(n384), .C(n349), .Z(n846) );
  CND2X2 U836 ( .A(n864), .B(n863), .Z(SUM[48]) );
  CENXL U837 ( .A(n106), .B(n10), .Z(SUM[60]) );
  CND2XL U838 ( .A(n881), .B(net16249), .Z(n883) );
  COND1XL U839 ( .A(n366), .B(n383), .C(n367), .Z(n365) );
  CNR2X1 U840 ( .A(A[35]), .B(B[35]), .Z(n322) );
  CANR1XL U841 ( .A(n118), .B(n3), .C(n859), .Z(n117) );
  CNR2X4 U842 ( .A(A[50]), .B(B[50]), .Z(n200) );
  CND2X2 U843 ( .A(A[50]), .B(B[50]), .Z(n201) );
  CND2X1 U844 ( .A(A[37]), .B(B[37]), .Z(n305) );
  CND2X1 U845 ( .A(A[35]), .B(B[35]), .Z(n323) );
  CENXL U846 ( .A(n259), .B(n847), .Z(SUM[43]) );
  CND2XL U847 ( .A(n572), .B(n258), .Z(n847) );
  CND2X2 U848 ( .A(n307), .B(n295), .Z(n293) );
  CND2IX2 U849 ( .B(A[36]), .A(n849), .Z(n848) );
  CNR2X2 U850 ( .A(n366), .B(n350), .Z(n348) );
  COND1X2 U851 ( .A(n158), .B(n193), .C(n159), .Z(n850) );
  COND1X1 U852 ( .A(n158), .B(n193), .C(n159), .Z(n3) );
  CIVX1 U853 ( .A(n193), .Z(n195) );
  CENXL U854 ( .A(n84), .B(n8), .Z(SUM[62]) );
  COND1X2 U855 ( .A(n172), .B(n162), .C(n163), .Z(n161) );
  COND1XL U856 ( .A(n210), .B(n2), .C(n211), .Z(n209) );
  COND1X1 U857 ( .A(n89), .B(n5), .C(n90), .Z(n88) );
  CANR1X1 U858 ( .A(n839), .B(n840), .C(n858), .Z(n853) );
  CND2X2 U859 ( .A(n228), .B(n244), .Z(n226) );
  COND1XL U860 ( .A(n100), .B(n5), .C(n101), .Z(n99) );
  CIVX1 U861 ( .A(n260), .Z(n262) );
  CIVXL U862 ( .A(n433), .Z(n432) );
  CND2X1 U863 ( .A(n228), .B(n244), .Z(net17940) );
  COND1X2 U864 ( .A(n226), .B(n261), .C(n227), .Z(n851) );
  COND1XL U865 ( .A(n818), .B(n226), .C(n227), .Z(n225) );
  CIVXL U866 ( .A(n209), .Z(n881) );
  COND1X2 U867 ( .A(n350), .B(n367), .C(n351), .Z(n349) );
  CND2X2 U868 ( .A(n583), .B(n823), .Z(n350) );
  CND2X1 U869 ( .A(n561), .B(n163), .Z(n16) );
  CANR1X1 U870 ( .A(n224), .B(n292), .C(n225), .Z(n852) );
  CANR1X1 U871 ( .A(n224), .B(n841), .C(n851), .Z(net18014) );
  CIVXL U872 ( .A(n162), .Z(n561) );
  CAN2XL U873 ( .A(n138), .B(n558), .Z(n129) );
  CIVX2 U874 ( .A(n367), .Z(n369) );
  CNR2X1 U875 ( .A(n131), .B(n124), .Z(n122) );
  CND2X2 U876 ( .A(A[41]), .B(B[41]), .Z(n276) );
  CENX1 U877 ( .A(n184), .B(n18), .Z(SUM[52]) );
  CND2IXL U878 ( .B(n182), .A(n183), .Z(n18) );
  COND1X1 U879 ( .A(n185), .B(net18013), .C(n186), .Z(n184) );
  CIVX2 U880 ( .A(n190), .Z(n188) );
  CANR1XL U881 ( .A(n835), .B(n195), .C(n177), .Z(n175) );
  CND2XL U882 ( .A(n194), .B(n564), .Z(n185) );
  CND2XL U883 ( .A(n564), .B(n190), .Z(n19) );
  CIVX2 U884 ( .A(n192), .Z(n194) );
  CND2XL U885 ( .A(n167), .B(n194), .Z(n165) );
  CND2XL U886 ( .A(n194), .B(n835), .Z(n174) );
  CANR1X2 U887 ( .A(n844), .B(n224), .C(n851), .Z(net18013) );
  CANR1X2 U888 ( .A(n213), .B(n198), .C(n199), .Z(n193) );
  COND1XL U889 ( .A(n192), .B(net18014), .C(n838), .Z(n191) );
  CNR2X1 U890 ( .A(A[51]), .B(B[51]), .Z(n189) );
  CNR2X4 U891 ( .A(n192), .B(n158), .Z(n4) );
  CANR1X1 U892 ( .A(n845), .B(n224), .C(n851), .Z(n2) );
  CIVX2 U893 ( .A(n842), .Z(n291) );
  CANR1XL U894 ( .A(n566), .B(n213), .C(n206), .Z(n204) );
  CIVX2 U895 ( .A(n213), .Z(n211) );
  CND2XL U896 ( .A(n566), .B(n208), .Z(n21) );
  COND1XL U897 ( .A(n111), .B(n853), .C(n114), .Z(n110) );
  CND2XL U898 ( .A(n109), .B(n4), .Z(n107) );
  CND2X1 U899 ( .A(A[60]), .B(B[60]), .Z(n105) );
  CNR2X2 U900 ( .A(n111), .B(n104), .Z(n102) );
  CNR2X1 U901 ( .A(n6), .B(n111), .Z(n109) );
  CANR1X2 U902 ( .A(n177), .B(n160), .C(n161), .Z(n159) );
  CIVX2 U903 ( .A(n111), .Z(n556) );
  CANR1X1 U904 ( .A(n139), .B(n122), .C(n123), .Z(n5) );
  COND1XL U905 ( .A(n78), .B(n853), .C(n79), .Z(n77) );
  CND2XL U906 ( .A(n556), .B(n114), .Z(n11) );
  CIVXL U907 ( .A(n177), .Z(n179) );
  CNR2X1 U908 ( .A(A[42]), .B(B[42]), .Z(n268) );
  COND1X1 U909 ( .A(n276), .B(n268), .C(n269), .Z(n267) );
  CND2X1 U910 ( .A(A[42]), .B(B[42]), .Z(n269) );
  CNR2X1 U911 ( .A(A[42]), .B(B[42]), .Z(net18513) );
  CENX1 U912 ( .A(n202), .B(n20), .Z(SUM[50]) );
  CIVX2 U913 ( .A(n208), .Z(n206) );
  CIVX2 U914 ( .A(n207), .Z(n566) );
  CND2XL U915 ( .A(n212), .B(n566), .Z(n203) );
  CNR2X2 U916 ( .A(n207), .B(n200), .Z(n198) );
  COND1X2 U917 ( .A(n222), .B(n218), .C(n219), .Z(n213) );
  CNR2X1 U918 ( .A(A[49]), .B(B[49]), .Z(n207) );
  CND2IXL U919 ( .B(n822), .A(n222), .Z(n23) );
  COND1X1 U920 ( .A(n822), .B(n2), .C(n222), .Z(n220) );
  CND2IXL U921 ( .B(n218), .A(n219), .Z(n22) );
  CND2X2 U922 ( .A(n856), .B(n287), .Z(n281) );
  CIVXL U923 ( .A(n281), .Z(n279) );
  CANR1XL U924 ( .A(n574), .B(n281), .C(n274), .Z(n272) );
  CND2X2 U925 ( .A(n854), .B(n855), .Z(n856) );
  CIVX2 U926 ( .A(n286), .Z(n855) );
  CND2X2 U927 ( .A(n266), .B(n280), .Z(n260) );
  CIVX1 U928 ( .A(n276), .Z(n274) );
  CND2X1 U929 ( .A(n574), .B(n276), .Z(n29) );
  CND2XL U930 ( .A(n573), .B(n269), .Z(n28) );
  CND2XL U931 ( .A(n855), .B(n287), .Z(n30) );
  COND1XL U932 ( .A(n289), .B(n291), .C(n290), .Z(n288) );
  CNR2X1 U933 ( .A(A[41]), .B(B[41]), .Z(n275) );
  CANR1X2 U934 ( .A(n245), .B(n228), .C(n229), .Z(n227) );
  COND1X1 U935 ( .A(n240), .B(net18512), .C(n231), .Z(n229) );
  CNR2X1 U936 ( .A(A[44]), .B(B[44]), .Z(n250) );
  CNR2X1 U937 ( .A(A[46]), .B(B[46]), .Z(n857) );
  CNR2X2 U938 ( .A(A[46]), .B(B[46]), .Z(net18512) );
  CIVXL U939 ( .A(n843), .Z(n569) );
  CND2XL U940 ( .A(n231), .B(n569), .Z(n24) );
  CNR2X2 U941 ( .A(A[45]), .B(B[45]), .Z(n237) );
  CND2XL U942 ( .A(A[45]), .B(B[45]), .Z(net18964) );
  CANR1X2 U943 ( .A(n295), .B(n308), .C(n296), .Z(n294) );
  CIVXL U944 ( .A(n817), .Z(n310) );
  COND1XL U945 ( .A(n302), .B(n310), .C(n814), .Z(n301) );
  CNR2X2 U946 ( .A(n302), .B(n297), .Z(n295) );
  CNR2IXL U947 ( .B(n307), .A(n302), .Z(n300) );
  CND2XL U948 ( .A(n91), .B(n94), .Z(n9) );
  CND2XL U949 ( .A(n4), .B(n87), .Z(n85) );
  CIVXL U950 ( .A(n103), .Z(n101) );
  CND2X1 U951 ( .A(A[61]), .B(B[61]), .Z(n94) );
  CNR2XL U952 ( .A(n487), .B(n490), .Z(n485) );
  CND2XL U953 ( .A(n559), .B(n145), .Z(n14) );
  CNR2XL U954 ( .A(A[16]), .B(B[16]), .Z(n464) );
  CND2XL U955 ( .A(n836), .B(n125), .Z(n12) );
  CIVXL U956 ( .A(n247), .Z(net18843) );
  CIVXL U957 ( .A(n263), .Z(net18840) );
  CAOR1XL U958 ( .A(n839), .B(n840), .C(n858), .Z(n859) );
  CND2X1 U959 ( .A(A[53]), .B(B[53]), .Z(n172) );
  CNR2X4 U960 ( .A(A[56]), .B(B[56]), .Z(n144) );
  CANR1X2 U961 ( .A(n348), .B(n384), .C(n349), .Z(n347) );
  COR2X1 U962 ( .A(B[17]), .B(A[17]), .Z(n872) );
  CIVX1 U963 ( .A(n465), .Z(n467) );
  CND2X1 U964 ( .A(n599), .B(n872), .Z(n457) );
  COND1X1 U965 ( .A(n506), .B(n494), .C(n495), .Z(n493) );
  CNR2X1 U966 ( .A(A[30]), .B(B[30]), .Z(n374) );
  CNR2X1 U967 ( .A(B[44]), .B(A[44]), .Z(net18589) );
  CND2X2 U968 ( .A(net17505), .B(net17506), .Z(n864) );
  CND2XL U969 ( .A(n209), .B(n21), .Z(n882) );
  CANR1XL U970 ( .A(n76), .B(n3), .C(n77), .Z(n75) );
  CANR1X2 U971 ( .A(n362), .B(n583), .C(n353), .Z(n351) );
  CANR1X1 U972 ( .A(n429), .B(n871), .C(n422), .Z(n420) );
  CIVXL U973 ( .A(n427), .Z(n429) );
  COND1X1 U974 ( .A(n491), .B(n487), .C(n488), .Z(n486) );
  CANR1X1 U975 ( .A(n502), .B(n876), .C(n497), .Z(n495) );
  CND2X2 U976 ( .A(A[57]), .B(B[57]), .Z(n134) );
  CIVX1 U977 ( .A(n323), .Z(n325) );
  CNR2XL U978 ( .A(n448), .B(n443), .Z(n441) );
  COND1X1 U979 ( .A(n449), .B(n443), .C(n444), .Z(n442) );
  CANR1X2 U980 ( .A(n325), .B(n848), .C(n316), .Z(n314) );
  CNR2X1 U981 ( .A(A[37]), .B(B[37]), .Z(n302) );
  COND1X2 U982 ( .A(n385), .B(n413), .C(n386), .Z(n384) );
  CNR2X2 U983 ( .A(A[57]), .B(B[57]), .Z(n131) );
  CENXL U984 ( .A(n37), .B(n346), .Z(SUM[33]) );
  CANR1X2 U985 ( .A(n380), .B(n585), .C(n373), .Z(n367) );
  CNR2X1 U986 ( .A(A[55]), .B(B[55]), .Z(n151) );
  CANR1X1 U987 ( .A(n138), .B(n850), .C(n837), .Z(n137) );
  CANR1X1 U988 ( .A(n467), .B(n872), .C(n460), .Z(n458) );
  CIVX1 U989 ( .A(n462), .Z(n460) );
  CIVXL U990 ( .A(n258), .Z(n256) );
  CNR2X1 U991 ( .A(A[43]), .B(B[43]), .Z(n257) );
  CANR1X2 U992 ( .A(n343), .B(n581), .C(n338), .Z(n332) );
  CND2X1 U993 ( .A(A[44]), .B(B[44]), .Z(n251) );
  CNR2X2 U994 ( .A(n331), .B(n313), .Z(n307) );
  CENXL U995 ( .A(n288), .B(n30), .Z(SUM[40]) );
  CND2X1 U996 ( .A(A[56]), .B(B[56]), .Z(n145) );
  CENXL U997 ( .A(n241), .B(n25), .Z(SUM[45]) );
  CND2X2 U998 ( .A(n860), .B(n861), .Z(n862) );
  CND2X2 U999 ( .A(n862), .B(n473), .Z(n471) );
  CIVX2 U1000 ( .A(n472), .Z(n860) );
  CND2XL U1001 ( .A(n874), .B(n873), .Z(n472) );
  CND2X1 U1002 ( .A(n220), .B(n22), .Z(n863) );
  CIVX1 U1003 ( .A(n220), .Z(net17505) );
  CIVX2 U1004 ( .A(n22), .Z(net17506) );
  CND2X2 U1005 ( .A(A[29]), .B(B[29]), .Z(n378) );
  CNR2X1 U1006 ( .A(A[29]), .B(B[29]), .Z(n377) );
  CND2XL U1007 ( .A(A[40]), .B(B[40]), .Z(n287) );
  CIVX1 U1008 ( .A(n377), .Z(n586) );
  CENXL U1009 ( .A(n270), .B(n28), .Z(SUM[42]) );
  CENXL U1010 ( .A(n232), .B(n24), .Z(SUM[46]) );
  CNR2X1 U1011 ( .A(A[32]), .B(B[32]), .Z(n354) );
  CND2X1 U1012 ( .A(A[28]), .B(B[28]), .Z(n390) );
  CENXL U1013 ( .A(n191), .B(n19), .Z(SUM[51]) );
  CENXL U1014 ( .A(n173), .B(n17), .Z(SUM[53]) );
  CENXL U1015 ( .A(n115), .B(n11), .Z(SUM[59]) );
  CENXL U1016 ( .A(n146), .B(n14), .Z(SUM[56]) );
  CENXL U1017 ( .A(n73), .B(n7), .Z(SUM[63]) );
  CNR2X2 U1018 ( .A(A[28]), .B(B[28]), .Z(n389) );
  CND2XL U1019 ( .A(A[38]), .B(B[38]), .Z(n298) );
  CANR1X1 U1020 ( .A(n471), .B(n452), .C(n453), .Z(n451) );
  CANR1XL U1021 ( .A(n471), .B(n452), .C(n453), .Z(n865) );
  CND2X1 U1022 ( .A(n875), .B(n869), .Z(n512) );
  CND2X1 U1023 ( .A(A[5]), .B(B[5]), .Z(n531) );
  CNR2X1 U1024 ( .A(n457), .B(n454), .Z(n452) );
  COND1XL U1025 ( .A(n174), .B(net18013), .C(n175), .Z(n173) );
  CANR1XL U1026 ( .A(n537), .B(n880), .C(n534), .Z(n532) );
  CND2X1 U1027 ( .A(A[54]), .B(B[54]), .Z(n163) );
  CND2X1 U1028 ( .A(A[25]), .B(B[25]), .Z(n411) );
  CND2X1 U1029 ( .A(A[43]), .B(B[43]), .Z(n258) );
  CND2XL U1030 ( .A(n4), .B(n129), .Z(n127) );
  CND2XL U1031 ( .A(n4), .B(n138), .Z(n136) );
  CND2XL U1032 ( .A(n262), .B(n572), .Z(n253) );
  CND2XL U1033 ( .A(n235), .B(n262), .Z(n233) );
  COND1X1 U1034 ( .A(n451), .B(n434), .C(n435), .Z(n433) );
  CND2XL U1035 ( .A(n441), .B(n870), .Z(n434) );
  CANR1X1 U1036 ( .A(n877), .B(n511), .C(n508), .Z(n506) );
  CANR1X1 U1037 ( .A(n878), .B(n529), .C(n526), .Z(n524) );
  COND1X1 U1038 ( .A(n532), .B(n530), .C(n531), .Z(n529) );
  CNR2X2 U1039 ( .A(n162), .B(n169), .Z(n160) );
  COND1X1 U1040 ( .A(n397), .B(n389), .C(n390), .Z(n388) );
  COND1X1 U1041 ( .A(n524), .B(n512), .C(n513), .Z(n511) );
  CIVXL U1042 ( .A(n850), .Z(n155) );
  CND2IXL U1043 ( .B(n169), .A(n172), .Z(n17) );
  CANR1X1 U1044 ( .A(n549), .B(n879), .C(n546), .Z(n544) );
  CIVXL U1045 ( .A(n424), .Z(n422) );
  CND2XL U1046 ( .A(n870), .B(n439), .Z(n49) );
  CND2XL U1047 ( .A(n873), .B(n477), .Z(n55) );
  CND2XL U1048 ( .A(n596), .B(n449), .Z(n51) );
  CND2XL U1049 ( .A(n874), .B(n482), .Z(n56) );
  CND2XL U1050 ( .A(n603), .B(n491), .Z(n58) );
  CND2XL U1051 ( .A(n875), .B(n517), .Z(n62) );
  CND2XL U1052 ( .A(n876), .B(n499), .Z(n59) );
  CND2XL U1053 ( .A(n868), .B(n504), .Z(n60) );
  CND2XL U1054 ( .A(n869), .B(n522), .Z(n63) );
  CND2XL U1055 ( .A(n880), .B(n536), .Z(n66) );
  CND2XL U1056 ( .A(n879), .B(n548), .Z(n69) );
  CND2IXL U1057 ( .B(n542), .A(n543), .Z(n68) );
  CNR2XL U1058 ( .A(A[22]), .B(B[22]), .Z(n426) );
  CNR2XL U1059 ( .A(A[3]), .B(B[3]), .Z(n538) );
  COND1XL U1060 ( .A(n74), .B(net18013), .C(n75), .Z(n73) );
  CND2XL U1061 ( .A(A[14]), .B(B[14]), .Z(n482) );
  CND2XL U1062 ( .A(B[26]), .B(A[26]), .Z(n406) );
  CND2XL U1063 ( .A(B[24]), .B(A[24]), .Z(n417) );
  CND2XL U1064 ( .A(A[13]), .B(B[13]), .Z(n488) );
  CND2XL U1065 ( .A(A[18]), .B(B[18]), .Z(n455) );
  CND2XL U1066 ( .A(A[20]), .B(B[20]), .Z(n444) );
  CND2XL U1067 ( .A(A[3]), .B(B[3]), .Z(n539) );
  COR2XL U1068 ( .A(A[7]), .B(B[7]), .Z(n869) );
  CENXL U1069 ( .A(n66), .B(n537), .Z(SUM[4]) );
  CND2IXL U1070 ( .B(n550), .A(n551), .Z(n70) );
  CIVXL U1071 ( .A(n402), .Z(n866) );
  CIVXL U1072 ( .A(n400), .Z(n402) );
  CND2XL U1073 ( .A(n4), .B(n118), .Z(n116) );
  CND2XL U1074 ( .A(n4), .B(n76), .Z(n74) );
  CANR1XL U1075 ( .A(n244), .B(n263), .C(net18843), .Z(n243) );
  CND2XL U1076 ( .A(n4), .B(n560), .Z(n147) );
  CND2XL U1077 ( .A(n280), .B(n574), .Z(n271) );
  CND2XL U1078 ( .A(n262), .B(n244), .Z(n242) );
  CNR2IXL U1079 ( .B(n244), .A(n237), .Z(n235) );
  COND1XL U1080 ( .A(n867), .B(n538), .C(n539), .Z(n537) );
  CND2X1 U1081 ( .A(n876), .B(n868), .Z(n494) );
  CND2X1 U1082 ( .A(n399), .B(n387), .Z(n385) );
  COND1XL U1083 ( .A(n116), .B(net18014), .C(n117), .Z(n115) );
  COND1XL U1084 ( .A(n147), .B(net18013), .C(n148), .Z(n146) );
  CANR1X1 U1085 ( .A(n414), .B(n433), .C(n415), .Z(n413) );
  CNR2X1 U1086 ( .A(n405), .B(n410), .Z(n399) );
  CANR1XL U1087 ( .A(n823), .B(n369), .C(n362), .Z(n358) );
  CND2XL U1088 ( .A(n570), .B(net18964), .Z(n25) );
  CND2XL U1089 ( .A(n571), .B(n251), .Z(n26) );
  CND2XL U1090 ( .A(n824), .B(n345), .Z(n37) );
  CND2XL U1091 ( .A(n583), .B(n355), .Z(n38) );
  COND1XL U1092 ( .A(n357), .B(n383), .C(n358), .Z(n356) );
  CND2XL U1093 ( .A(n368), .B(n823), .Z(n357) );
  CND2XL U1094 ( .A(n823), .B(n364), .Z(n39) );
  CND2XL U1095 ( .A(n585), .B(n375), .Z(n40) );
  COND1XL U1096 ( .A(n377), .B(n383), .C(n815), .Z(n376) );
  CANR1XL U1097 ( .A(n263), .B(n235), .C(n236), .Z(n234) );
  CND2XL U1098 ( .A(n560), .B(n152), .Z(n15) );
  COND1XL U1099 ( .A(n271), .B(n291), .C(n272), .Z(n270) );
  CEOXL U1100 ( .A(n341), .B(n36), .Z(SUM[34]) );
  CND2XL U1101 ( .A(n581), .B(n340), .Z(n36) );
  CANR1XL U1102 ( .A(n824), .B(n346), .C(n343), .Z(n341) );
  CANR1XL U1103 ( .A(n392), .B(n412), .C(n393), .Z(n391) );
  CANR1XL U1104 ( .A(n399), .B(n412), .C(n866), .Z(n398) );
  CANR1XL U1105 ( .A(n590), .B(n412), .C(n409), .Z(n407) );
  CNR2XL U1106 ( .A(n331), .B(n322), .Z(n320) );
  COAN1X1 U1107 ( .A(n542), .B(n544), .C(n543), .Z(n867) );
  CND2X1 U1108 ( .A(n585), .B(n586), .Z(n366) );
  CND2XL U1109 ( .A(n590), .B(n411), .Z(n45) );
  COND1XL U1110 ( .A(n419), .B(n432), .C(n420), .Z(n418) );
  CENX1 U1111 ( .A(n425), .B(n47), .Z(SUM[23]) );
  CND2X1 U1112 ( .A(n871), .B(n424), .Z(n47) );
  COND1XL U1113 ( .A(n426), .B(n432), .C(n427), .Z(n425) );
  CENX1 U1114 ( .A(n450), .B(n51), .Z(SUM[19]) );
  CENX1 U1115 ( .A(n456), .B(n52), .Z(SUM[18]) );
  CND2X1 U1116 ( .A(n597), .B(n455), .Z(n52) );
  COND1XL U1117 ( .A(n457), .B(n470), .C(n458), .Z(n456) );
  CENX1 U1118 ( .A(n463), .B(n53), .Z(SUM[17]) );
  CND2X1 U1119 ( .A(n872), .B(n462), .Z(n53) );
  COND1XL U1120 ( .A(n464), .B(n470), .C(n465), .Z(n463) );
  CENX1 U1121 ( .A(n483), .B(n56), .Z(SUM[14]) );
  CENX1 U1122 ( .A(n489), .B(n57), .Z(SUM[13]) );
  CND2X1 U1123 ( .A(n602), .B(n488), .Z(n57) );
  COND1XL U1124 ( .A(n490), .B(n492), .C(n491), .Z(n489) );
  COND1XL U1125 ( .A(n394), .B(n402), .C(n397), .Z(n393) );
  CEOXL U1126 ( .A(n48), .B(n432), .Z(SUM[22]) );
  CND2XL U1127 ( .A(n593), .B(n427), .Z(n48) );
  CEOXL U1128 ( .A(n49), .B(n440), .Z(SUM[21]) );
  CANR1XL U1129 ( .A(n441), .B(n450), .C(n442), .Z(n440) );
  CEOXL U1130 ( .A(n50), .B(n445), .Z(SUM[20]) );
  CANR1XL U1131 ( .A(n596), .B(n450), .C(n447), .Z(n445) );
  CEOXL U1132 ( .A(n54), .B(n470), .Z(SUM[16]) );
  CND2XL U1133 ( .A(n599), .B(n465), .Z(n54) );
  CEOXL U1134 ( .A(n55), .B(n478), .Z(SUM[15]) );
  CANR1XL U1135 ( .A(n874), .B(n483), .C(n480), .Z(n478) );
  CNR2IXL U1136 ( .B(n399), .A(n394), .Z(n392) );
  CENX1 U1137 ( .A(n60), .B(n505), .Z(SUM[10]) );
  CENX1 U1138 ( .A(n61), .B(n511), .Z(SUM[9]) );
  CND2X1 U1139 ( .A(n877), .B(n510), .Z(n61) );
  CENX1 U1140 ( .A(n63), .B(n523), .Z(SUM[7]) );
  CENX1 U1141 ( .A(n64), .B(n529), .Z(SUM[6]) );
  CND2X1 U1142 ( .A(n878), .B(n528), .Z(n64) );
  CEOXL U1143 ( .A(n58), .B(n492), .Z(SUM[12]) );
  CEOXL U1144 ( .A(n59), .B(n500), .Z(SUM[11]) );
  CANR1XL U1145 ( .A(n868), .B(n505), .C(n502), .Z(n500) );
  CEOXL U1146 ( .A(n518), .B(n62), .Z(SUM[8]) );
  CANR1XL U1147 ( .A(n869), .B(n523), .C(n520), .Z(n518) );
  CEOXL U1148 ( .A(n532), .B(n65), .Z(SUM[5]) );
  CND2X1 U1149 ( .A(n610), .B(n531), .Z(n65) );
  CND2IX1 U1150 ( .B(n538), .A(n539), .Z(n67) );
  CNR2X1 U1151 ( .A(A[39]), .B(B[39]), .Z(n289) );
  CNR2X1 U1152 ( .A(A[24]), .B(B[24]), .Z(n416) );
  CNR2X1 U1153 ( .A(A[18]), .B(B[18]), .Z(n454) );
  CNR2X1 U1154 ( .A(A[26]), .B(B[26]), .Z(n405) );
  CNR2X1 U1155 ( .A(A[47]), .B(B[47]), .Z(n221) );
  CNR2X1 U1156 ( .A(A[13]), .B(B[13]), .Z(n487) );
  CNR2X1 U1157 ( .A(A[25]), .B(B[25]), .Z(n410) );
  CND2X1 U1158 ( .A(A[63]), .B(B[63]), .Z(n72) );
  CNR2X1 U1159 ( .A(A[5]), .B(B[5]), .Z(n530) );
  COR2X1 U1160 ( .A(A[10]), .B(B[10]), .Z(n868) );
  COR2X1 U1161 ( .A(A[21]), .B(B[21]), .Z(n870) );
  COR2X1 U1162 ( .A(A[23]), .B(B[23]), .Z(n871) );
  COR2X1 U1163 ( .A(A[15]), .B(B[15]), .Z(n873) );
  CND2X1 U1164 ( .A(A[22]), .B(B[22]), .Z(n427) );
  CND2X1 U1165 ( .A(A[16]), .B(B[16]), .Z(n465) );
  COR2X1 U1166 ( .A(A[14]), .B(B[14]), .Z(n874) );
  COR2X1 U1167 ( .A(A[8]), .B(B[8]), .Z(n875) );
  COR2X1 U1168 ( .A(B[11]), .B(A[11]), .Z(n876) );
  CND2X1 U1169 ( .A(A[19]), .B(B[19]), .Z(n449) );
  CND2X1 U1170 ( .A(A[27]), .B(B[27]), .Z(n397) );
  CND2X1 U1171 ( .A(A[12]), .B(B[12]), .Z(n491) );
  CND2X1 U1172 ( .A(A[33]), .B(B[33]), .Z(n345) );
  CND2X1 U1173 ( .A(A[34]), .B(B[34]), .Z(n340) );
  CND2X1 U1174 ( .A(A[31]), .B(B[31]), .Z(n364) );
  CND2X1 U1175 ( .A(A[30]), .B(B[30]), .Z(n375) );
  CND2X1 U1176 ( .A(A[32]), .B(B[32]), .Z(n355) );
  CND2X1 U1177 ( .A(A[10]), .B(B[10]), .Z(n504) );
  CND2X1 U1178 ( .A(A[7]), .B(B[7]), .Z(n522) );
  CND2X1 U1179 ( .A(A[23]), .B(B[23]), .Z(n424) );
  CND2X1 U1180 ( .A(A[17]), .B(B[17]), .Z(n462) );
  CND2X1 U1181 ( .A(A[21]), .B(B[21]), .Z(n439) );
  CND2X1 U1182 ( .A(A[8]), .B(B[8]), .Z(n517) );
  CND2X1 U1183 ( .A(A[15]), .B(B[15]), .Z(n477) );
  CND2X1 U1184 ( .A(A[11]), .B(B[11]), .Z(n499) );
  CND2X1 U1185 ( .A(A[9]), .B(B[9]), .Z(n510) );
  CND2X1 U1186 ( .A(A[1]), .B(B[1]), .Z(n548) );
  CND2X1 U1187 ( .A(A[4]), .B(B[4]), .Z(n536) );
  CND2X1 U1188 ( .A(A[6]), .B(B[6]), .Z(n528) );
  CND2X1 U1189 ( .A(A[58]), .B(B[58]), .Z(n125) );
  COR2X1 U1190 ( .A(A[9]), .B(B[9]), .Z(n877) );
  COR2X1 U1191 ( .A(A[6]), .B(B[6]), .Z(n878) );
  COR2X1 U1192 ( .A(A[1]), .B(B[1]), .Z(n879) );
  COR2X1 U1193 ( .A(A[4]), .B(B[4]), .Z(n880) );
  CNR2X1 U1194 ( .A(A[2]), .B(B[2]), .Z(n542) );
  CND2X1 U1195 ( .A(A[0]), .B(B[0]), .Z(n551) );
  CND2X1 U1196 ( .A(A[2]), .B(B[2]), .Z(n543) );
  CEOXL U1197 ( .A(n867), .B(n67), .Z(SUM[3]) );
  CEOXL U1198 ( .A(n544), .B(n68), .Z(SUM[2]) );
  CENX1 U1199 ( .A(n69), .B(n549), .Z(SUM[1]) );
  CNR2XL U1200 ( .A(A[0]), .B(B[0]), .Z(n550) );
  CND2X1 U1201 ( .A(A[48]), .B(B[48]), .Z(n219) );
  CIVXL U1202 ( .A(n237), .Z(n570) );
  COND1XL U1203 ( .A(n237), .B(n247), .C(net18964), .Z(n236) );
  CIVXL U1204 ( .A(net18589), .Z(n571) );
  COND1XL U1205 ( .A(n242), .B(n291), .C(n243), .Z(n241) );
  COND1XL U1206 ( .A(n291), .B(n233), .C(n234), .Z(n232) );
  CIVXL U1207 ( .A(net18513), .Z(n573) );
  CEOXL U1208 ( .A(n23), .B(net18013), .Z(SUM[47]) );
  COND1XL U1209 ( .A(n322), .B(n332), .C(n323), .Z(n321) );
  CIVX2 U1210 ( .A(n21), .Z(net16249) );
  CENX1 U1211 ( .A(n135), .B(n13), .Z(SUM[57]) );
  CENX1 U1212 ( .A(n126), .B(n12), .Z(SUM[58]) );
  CIVX2 U1213 ( .A(n530), .Z(n610) );
  CIVX2 U1214 ( .A(n490), .Z(n603) );
  CIVX2 U1215 ( .A(n487), .Z(n602) );
  CIVX2 U1216 ( .A(n454), .Z(n597) );
  CIVX2 U1217 ( .A(n394), .Z(n588) );
  CIVX2 U1218 ( .A(n302), .Z(n578) );
  CIVX2 U1219 ( .A(n289), .Z(n576) );
  CIVX2 U1220 ( .A(n144), .Z(n559) );
  CIVX2 U1221 ( .A(n131), .Z(n558) );
  CIVX2 U1222 ( .A(n71), .Z(n552) );
  CIVX2 U1223 ( .A(n551), .Z(n549) );
  CIVX2 U1224 ( .A(n548), .Z(n546) );
  CIVX2 U1225 ( .A(n536), .Z(n534) );
  CIVX2 U1226 ( .A(n528), .Z(n526) );
  CIVX2 U1227 ( .A(n524), .Z(n523) );
  CIVX2 U1228 ( .A(n522), .Z(n520) );
  CIVX2 U1229 ( .A(n517), .Z(n515) );
  CIVX2 U1230 ( .A(n510), .Z(n508) );
  CIVX2 U1231 ( .A(n504), .Z(n502) );
  CIVX2 U1232 ( .A(n471), .Z(n470) );
  CIVX2 U1233 ( .A(n865), .Z(n450) );
  CIVX2 U1234 ( .A(n449), .Z(n447) );
  CIVX2 U1235 ( .A(n448), .Z(n596) );
  CIVX2 U1236 ( .A(n439), .Z(n437) );
  CIVX2 U1237 ( .A(n426), .Z(n593) );
  CIVX2 U1238 ( .A(n411), .Z(n409) );
  CIVX2 U1239 ( .A(n410), .Z(n590) );
  CIVX2 U1240 ( .A(n378), .Z(n380) );
  CIVX2 U1241 ( .A(n366), .Z(n368) );
  CIVX2 U1242 ( .A(n364), .Z(n362) );
  CIVX2 U1243 ( .A(n355), .Z(n353) );
  CIVX2 U1244 ( .A(n354), .Z(n583) );
  CIVX2 U1245 ( .A(n345), .Z(n343) );
  CIVX2 U1246 ( .A(n340), .Z(n338) );
  CIVX2 U1247 ( .A(n339), .Z(n581) );
  CIVX2 U1248 ( .A(n331), .Z(n329) );
  CIVX2 U1249 ( .A(n322), .Z(n580) );
  CIVX2 U1250 ( .A(n280), .Z(n278) );
  CIVX2 U1251 ( .A(n152), .Z(n150) );
  CIVX2 U1252 ( .A(n151), .Z(n560) );
  CIVX2 U1253 ( .A(n102), .Z(n100) );
  CIVX2 U1254 ( .A(n70), .Z(SUM[0]) );
endmodule


module sfilt_DW_mult_tc_4 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n9, n12, n15, n18, n21, n24, n27, n30, n39, n45, n48, n54,
         n57, n63, n66, n75, n78, n81, n84, n87, n90, n93, n96, n99, n102,
         n105, n111, n117, n120, n123, n129, n135, n136, n144, n145, n150,
         n151, n152, n153, n154, n155, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n171, n175, n176, n177,
         n178, n179, n182, n183, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n198, n200, n201, n202, n204, n205,
         n206, n207, n208, n209, n210, n212, n213, n214, n216, n218, n219,
         n220, n221, n222, n223, n224, n225, n227, n229, n230, n231, n232,
         n233, n236, n241, n242, n244, n246, n247, n248, n249, n253, n255,
         n256, n257, n258, n259, n260, n261, n262, n264, n265, n266, n267,
         n268, n269, n272, n273, n274, n275, n277, n279, n280, n281, n282,
         n283, n286, n291, n292, n293, n294, n295, n296, n298, n299, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n314, n316,
         n317, n318, n319, n320, n323, n324, n327, n328, n329, n330, n331,
         n332, n333, n334, n340, n341, n342, n343, n344, n345, n349, n351,
         n352, n353, n354, n355, n356, n359, n360, n361, n362, n363, n364,
         n365, n366, n369, n370, n371, n372, n373, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n392, n393,
         n394, n395, n396, n397, n399, n402, n403, n404, n405, n406, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n426, n427, n428, n432, n433, n434, n435, n439, n441, n445, n448,
         n449, n450, n451, n452, n456, n469, n470, n471, n472, n487, n488,
         n489, n490, n495, n496, n497, n498, n506, n507, n508, n510, n511,
         n513, n514, n516, n517, n520, n522, n523, n524, n525, n526, n528,
         n529, n530, n531, n532, n533, n534, n540, n541, n542, n543, n544,
         n545, n551, n552, n553, n554, n555, n556, n560, n561, n562, n564,
         n567, n568, n569, n571, n572, n573, n574, n575, n576, n577, n579,
         n582, n583, n584, n585, n586, n590, n591, n592, n593, n594, n595,
         n596, n603, n604, n605, n606, n611, n612, n613, n614, n616, n618,
         n619, n620, n621, n622, n623, n624, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n639, n641, n642, n643,
         n644, n646, n651, n652, n654, n656, n657, n658, n659, n660, n661,
         n662, n664, n665, n666, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n681, n683, n684, n686, n688, n689,
         n690, n691, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n704, n706, n707, n708, n709, n710, n712, n714, n718, n720,
         n721, n722, n723, n724, n726, n728, n729, n731, n736, n738, n739,
         n741, n742, n744, n745, n746, n747, n748, n750, n751, n758, n760,
         n761, n762, n765, n766, n767, n768, n770, n772, n773, n774, n776,
         n778, n779, n780, n781, n784, n785, n786, n788, n791, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1110, n1111, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1135, n1137, n1139, n1145, n1146, n1147, n1148, n1149,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1161, n1162,
         n1163, n1164, n1165, n1167, n1171, n1173, n1180, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1203, n1204, n1205, n1206, n1207, n1210, n1211,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2812, n2813, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2825, n2826,
         n2827, net15916, net15914, net15912, net15910, net15974, net15988,
         net16102, net16104, net16270, net16274, net16301, net16309, net16413,
         net16416, net16420, net16419, net16426, net16433, net16439, net16438,
         net16437, net16451, net16465, net16472, net16471, net16490, net16497,
         net16496, net16512, net16511, net16510, net16541, net16959, net17136,
         net17154, net17211, net17279, net17278, net17297, net17411, net17410,
         net17419, net17425, net17439, net17438, net17451, net17512, net17728,
         net17727, net17738, net17759, net17758, net17756, net17755, net17791,
         net17930, net17986, net18061, net18180, net18200, net18199, net18211,
         net18209, net18218, net18310, net18400, net18496, net18534, net18532,
         net18548, net18561, net18574, net18593, net18592, net18610, net18614,
         net18627, net18628, net18689, net18718, net18772, net18817, net18824,
         net18828, net18827, net18832, net18863, net18897, net18896, net18914,
         net18913, net19006, net19057, net19060, net18507, net18505, n2650,
         n462, n458, n444, n170, net18204, n549, net17942, n535, n515, n754,
         n753, n559, n550, n548, n547, n546, n479, n478, n474, n468, n467,
         n461, n459, n149, net18527, n494, n491, n485, n484, n483, n482, n481,
         n1184, net18519, n512, n505, n504, n499, net16974, net16962, n1134,
         n1107, n1106, n1083, net17985, net17984, n1973, n1212, n1185, n1175,
         n1174, n1172, n1166, n1141, n1140, net18422, net18420, net18419,
         net15980, n2095, n1880, n2004, n1911, n1856, n1825, n1794, n1763,
         n1202, n1179, n1178, n1177, n1176, n1169, n1168, n114, net18261,
         net17725, net17724, net17723, n2126, n2005, n1942, n1881, n1826,
         n1209, n1208, n1183, n1182, n1181, n1170, net19067, net19066,
         net17989, net17987, n1824, n1793, n1151, n1150, n1144, n1143, n1142,
         n1138, n1136, n1113, n1112, n1109, n1108, net17483, net17482, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n57 = a[13];
  assign n66 = a[15];
  assign n75 = a[17];
  assign n84 = a[19];
  assign n93 = a[21];
  assign n102 = a[23];
  assign n111 = a[25];
  assign n120 = a[27];
  assign n129 = a[29];
  assign n136 = a[31];
  assign n145 = b[0];
  assign n2780 = b[31];
  assign n2781 = b[30];
  assign n2782 = b[29];
  assign n2783 = b[28];
  assign n2784 = b[27];
  assign n2785 = b[26];
  assign n2786 = b[25];
  assign n2787 = b[24];
  assign n2788 = b[23];
  assign n2789 = b[22];
  assign n2790 = b[21];
  assign n2791 = b[20];
  assign n2792 = b[19];
  assign n2793 = b[18];
  assign n2794 = b[17];
  assign n2795 = b[16];
  assign n2796 = b[15];
  assign n2797 = b[14];
  assign n2798 = b[13];
  assign n2799 = b[12];
  assign n2800 = b[11];
  assign n2801 = b[10];
  assign n2802 = b[9];
  assign n2803 = b[8];
  assign n2804 = b[7];
  assign n2805 = b[6];
  assign n2806 = b[5];
  assign n2807 = b[4];
  assign n2808 = b[3];
  assign n2809 = b[2];
  assign n2810 = b[1];

  CNR2X2 U181 ( .A(n274), .B(n4483), .Z(n233) );
  CANR1X1 U188 ( .A(n4497), .B(n253), .C(n244), .Z(n242) );
  CANR1X1 U214 ( .A(n736), .B(n273), .C(n264), .Z(n262) );
  CND2X2 U229 ( .A(n283), .B(n4490), .Z(n274) );
  CANR1X1 U230 ( .A(n4490), .B(n286), .C(n277), .Z(n275) );
  COND1X1 U244 ( .A(n4482), .B(n334), .C(n4477), .Z(n286) );
  CNR2X2 U255 ( .A(n813), .B(n818), .Z(n295) );
  CANR1X1 U260 ( .A(n739), .B(n308), .C(n301), .Z(n299) );
  CNR2X2 U265 ( .A(n826), .B(n819), .Z(n302) );
  CND2X2 U266 ( .A(n826), .B(n819), .Z(n303) );
  COND1X1 U272 ( .A(n309), .B(n3732), .C(n310), .Z(n308) );
  COND1X1 U284 ( .A(n318), .B(net16472), .C(n319), .Z(n317) );
  CANR1X1 U286 ( .A(n320), .B(n356), .C(n323), .Z(n319) );
  CNR2X2 U295 ( .A(n835), .B(n844), .Z(n324) );
  COND1X1 U298 ( .A(n329), .B(net16472), .C(n330), .Z(n328) );
  CANR1X1 U308 ( .A(n349), .B(n742), .C(n340), .Z(n334) );
  CNR2X2 U313 ( .A(n845), .B(n854), .Z(n341) );
  COND1X1 U316 ( .A(n344), .B(net16472), .C(n345), .Z(n343) );
  CANR1X1 U318 ( .A(n4479), .B(n356), .C(n349), .Z(n345) );
  COND1X1 U328 ( .A(n353), .B(net16472), .C(n4074), .Z(n352) );
  CNR2X2 U335 ( .A(n361), .B(n416), .Z(n359) );
  COND1X1 U336 ( .A(n417), .B(n361), .C(n362), .Z(n360) );
  CNR2X2 U339 ( .A(n365), .B(n389), .Z(n363) );
  CNR2X2 U347 ( .A(n878), .B(n867), .Z(n369) );
  COND1X1 U350 ( .A(n372), .B(net16472), .C(n373), .Z(n371) );
  CANR1X1 U352 ( .A(n745), .B(n384), .C(n377), .Z(n373) );
  CNR2X2 U359 ( .A(n879), .B(n892), .Z(n378) );
  CND2X2 U360 ( .A(n3567), .B(n892), .Z(n379) );
  COND1X1 U362 ( .A(n381), .B(net16472), .C(n382), .Z(n380) );
  COND1X1 U366 ( .A(n385), .B(n441), .C(n386), .Z(n384) );
  CNR2X2 U375 ( .A(n893), .B(n906), .Z(n389) );
  COND1X1 U378 ( .A(n394), .B(net16472), .C(n395), .Z(n393) );
  CNR2X2 U389 ( .A(n907), .B(n922), .Z(n402) );
  COND1X1 U392 ( .A(n405), .B(net16472), .C(n406), .Z(n404) );
  CNR2X2 U405 ( .A(n3196), .B(n416), .Z(n414) );
  COND1X1 U406 ( .A(n416), .B(n441), .C(n417), .Z(n415) );
  COND1X1 U420 ( .A(n427), .B(net16471), .C(n428), .Z(n426) );
  COND1X1 U450 ( .A(n451), .B(net16471), .C(n452), .Z(n450) );
  COND1X1 U548 ( .A(n525), .B(n545), .C(n526), .Z(n524) );
  COND1X1 U572 ( .A(n4073), .B(n545), .C(n544), .Z(n542) );
  CND2X2 U576 ( .A(n1245), .B(n1274), .Z(n544) );
  CNR2X2 U608 ( .A(n1333), .B(n1360), .Z(n567) );
  CNR2X2 U629 ( .A(n1387), .B(n1412), .Z(n582) );
  COND1X1 U632 ( .A(n585), .B(n611), .C(n586), .Z(n584) );
  CNR2X2 U641 ( .A(n1436), .B(n1413), .Z(n591) );
  COND1X1 U760 ( .A(n674), .B(n676), .C(n675), .Z(n673) );
  CFA1X1 U858 ( .A(n800), .B(n1769), .CI(n1741), .CO(n796), .S(n797) );
  CFA1X1 U859 ( .A(n1770), .B(n804), .CI(n801), .CO(n798), .S(n799) );
  CFA1X1 U861 ( .A(n1742), .B(n805), .CI(n808), .CO(n802), .S(n803) );
  CFA1X1 U862 ( .A(n810), .B(n1802), .CI(n1771), .CO(n804), .S(n805) );
  CFA1X1 U863 ( .A(n816), .B(n814), .CI(n809), .CO(n806), .S(n807) );
  CFA1X1 U864 ( .A(n1803), .B(n811), .CI(n1772), .CO(n808), .S(n809) );
  CFA1X1 U866 ( .A(n817), .B(n815), .CI(n820), .CO(n812), .S(n813) );
  CFA1X1 U867 ( .A(n1743), .B(n822), .CI(n1804), .CO(n814), .S(n815) );
  CFA1X1 U868 ( .A(n824), .B(n1835), .CI(n1773), .CO(n816), .S(n817) );
  CFA1X1 U869 ( .A(n823), .B(n828), .CI(n821), .CO(n818), .S(n819) );
  CFA1X1 U870 ( .A(n825), .B(n830), .CI(n832), .CO(n820), .S(n821) );
  CFA1X1 U871 ( .A(n1774), .B(n1836), .CI(n1805), .CO(n822), .S(n823) );
  CFA1X1 U873 ( .A(n838), .B(n836), .CI(n829), .CO(n826), .S(n827) );
  CFA1X1 U874 ( .A(n840), .B(n831), .CI(n833), .CO(n828), .S(n829) );
  CFA1X1 U875 ( .A(n1744), .B(n1806), .CI(n1775), .CO(n830), .S(n831) );
  CFA1X1 U877 ( .A(n839), .B(n837), .CI(n846), .CO(n834), .S(n835) );
  CFA1X1 U878 ( .A(n850), .B(n848), .CI(n841), .CO(n836), .S(n837) );
  CFA1X1 U879 ( .A(n1807), .B(n852), .CI(n843), .CO(n838), .S(n839) );
  CFA1X1 U880 ( .A(n1745), .B(n1776), .CI(n1838), .CO(n840), .S(n841) );
  CFA1X1 U882 ( .A(n849), .B(n847), .CI(n856), .CO(n844), .S(n845) );
  CFA1X1 U883 ( .A(n851), .B(n858), .CI(n853), .CO(n846), .S(n847) );
  CFA1X1 U884 ( .A(n1894), .B(n860), .CI(n862), .CO(n848), .S(n849) );
  CFA1X1 U885 ( .A(n1869), .B(n1839), .CI(n1746), .CO(n850), .S(n851) );
  CFA1X1 U887 ( .A(n859), .B(n857), .CI(n868), .CO(n854), .S(n855) );
  CFA1X1 U888 ( .A(n861), .B(n870), .CI(n872), .CO(n856), .S(n857) );
  CFA1X1 U889 ( .A(n876), .B(n863), .CI(n874), .CO(n858), .S(n859) );
  CFA1X1 U890 ( .A(n1809), .B(n865), .CI(n1778), .CO(n860), .S(n861) );
  CFA1X1 U891 ( .A(n1747), .B(n1840), .CI(n1895), .CO(n862), .S(n863) );
  CFA1X1 U894 ( .A(n884), .B(n882), .CI(n873), .CO(n868), .S(n869) );
  CFA1X1 U895 ( .A(n886), .B(n877), .CI(n875), .CO(n870), .S(n871) );
  CFA1X1 U896 ( .A(n1748), .B(n888), .CI(n1927), .CO(n872), .S(n873) );
  CFA1X1 U898 ( .A(n890), .B(n1810), .CI(n1841), .CO(n876), .S(n877) );
  CFA1X1 U899 ( .A(n883), .B(n881), .CI(n894), .CO(n878), .S(n879) );
  CFA1X1 U901 ( .A(n900), .B(n887), .CI(n889), .CO(n882), .S(n883) );
  CFA1X1 U902 ( .A(n891), .B(n902), .CI(n904), .CO(n884), .S(n885) );
  CFA1X1 U903 ( .A(n1842), .B(n1811), .CI(n1780), .CO(n886), .S(n887) );
  CFA1X1 U904 ( .A(n1749), .B(n1897), .CI(n1928), .CO(n888), .S(n889) );
  CFA1X1 U906 ( .A(n897), .B(n895), .CI(n908), .CO(n892), .S(n893) );
  CFA1X1 U908 ( .A(n905), .B(n914), .CI(n901), .CO(n896), .S(n897) );
  CFA1X1 U909 ( .A(n918), .B(n903), .CI(n916), .CO(n898), .S(n899) );
  CFA1X1 U910 ( .A(n1750), .B(n1960), .CI(n1898), .CO(n900), .S(n901) );
  CFA1X1 U912 ( .A(n920), .B(n1781), .CI(n1929), .CO(n904), .S(n905) );
  CFA1X1 U913 ( .A(n911), .B(n909), .CI(n924), .CO(n906), .S(n907) );
  CFA1X1 U916 ( .A(n934), .B(n919), .CI(n932), .CO(n912), .S(n913) );
  CFA1X1 U917 ( .A(n1844), .B(n936), .CI(n921), .CO(n914), .S(n915) );
  CFA1X1 U918 ( .A(n1899), .B(n1813), .CI(n1782), .CO(n916), .S(n917) );
  CFA1X1 U922 ( .A(n944), .B(n942), .CI(n929), .CO(n924), .S(n925) );
  CFA1X1 U924 ( .A(n948), .B(n935), .CI(n937), .CO(n928), .S(n929) );
  CFA1X1 U925 ( .A(n1814), .B(n950), .CI(n952), .CO(n930), .S(n931) );
  CFA1X1 U926 ( .A(n1752), .B(n1993), .CI(n1783), .CO(n932), .S(n933) );
  CFA1X1 U928 ( .A(n954), .B(n1845), .CI(n1962), .CO(n936), .S(n937) );
  CFA1X1 U929 ( .A(n943), .B(n941), .CI(n958), .CO(n938), .S(n939) );
  CFA1X1 U931 ( .A(n966), .B(n947), .CI(n964), .CO(n942), .S(n943) );
  CFA1X1 U932 ( .A(n953), .B(n949), .CI(n951), .CO(n944), .S(n945) );
  CFA1X1 U933 ( .A(n972), .B(n968), .CI(n970), .CO(n946), .S(n947) );
  CFA1X1 U934 ( .A(n1963), .B(n955), .CI(n1932), .CO(n948), .S(n949) );
  CFA1X1 U935 ( .A(n1815), .B(n1846), .CI(n1901), .CO(n950), .S(n951) );
  CFA1X1 U938 ( .A(n961), .B(n959), .CI(n976), .CO(n956), .S(n957) );
  CFA1X1 U939 ( .A(n980), .B(n978), .CI(n963), .CO(n958), .S(n959) );
  CFA1X1 U940 ( .A(n982), .B(n965), .CI(n967), .CO(n960), .S(n961) );
  CFA1X1 U941 ( .A(n973), .B(n984), .CI(n969), .CO(n962), .S(n963) );
  CFA1X1 U943 ( .A(n1964), .B(n990), .CI(n1933), .CO(n966), .S(n967) );
  CFA1X1 U944 ( .A(n1754), .B(n1816), .CI(n1785), .CO(n968), .S(n969) );
  CFA1X1 U945 ( .A(n1847), .B(n1902), .CI(n1873), .CO(n970), .S(n971) );
  CFA1X1 U948 ( .A(n1000), .B(n998), .CI(n981), .CO(n976), .S(n977) );
  CFA1X1 U950 ( .A(n989), .B(n1004), .CI(n987), .CO(n980), .S(n981) );
  CFA1X1 U952 ( .A(n993), .B(n1010), .CI(n1012), .CO(n984), .S(n985) );
  CFA1X1 U953 ( .A(n1903), .B(n1848), .CI(n1817), .CO(n986), .S(n987) );
  CFA1X1 U954 ( .A(n1755), .B(n1786), .CI(n1934), .CO(n988), .S(n989) );
  CFA1X1 U955 ( .A(n1874), .B(n1996), .CI(n1965), .CO(n990), .S(n991) );
  CFA1X1 U959 ( .A(n1005), .B(n1003), .CI(n1022), .CO(n998), .S(n999) );
  CFA1X1 U960 ( .A(n1011), .B(n1024), .CI(n1026), .CO(n1000), .S(n1001) );
  CFA1X1 U962 ( .A(n1032), .B(n1028), .CI(n1030), .CO(n1004), .S(n1005) );
  CFA1X1 U963 ( .A(n1756), .B(n2057), .CI(n1997), .CO(n1006), .S(n1007) );
  CFA1X1 U965 ( .A(n2027), .B(n1935), .CI(n1904), .CO(n1010), .S(n1011) );
  CFA1X1 U966 ( .A(n1818), .B(n1034), .CI(n1966), .CO(n1012), .S(n1013) );
  CFA1X1 U973 ( .A(n1850), .B(n1056), .CI(n1035), .CO(n1026), .S(n1027) );
  CFA1X1 U974 ( .A(n1788), .B(n1819), .CI(n1967), .CO(n1028), .S(n1029) );
  CFA1X1 U976 ( .A(n1936), .B(n1905), .CI(n2028), .CO(n1032), .S(n1033) );
  CFA1X1 U979 ( .A(n1064), .B(n1062), .CI(n1043), .CO(n1038), .S(n1039) );
  CFA1X1 U981 ( .A(n1070), .B(n1068), .CI(n1049), .CO(n1042), .S(n1043) );
  CFA1X1 U983 ( .A(n1074), .B(n1055), .CI(n1072), .CO(n1046), .S(n1047) );
  CFA1X1 U984 ( .A(n1968), .B(n1076), .CI(n1078), .CO(n1048), .S(n1049) );
  CFA1X1 U985 ( .A(n1758), .B(n2090), .CI(n1906), .CO(n1050), .S(n1051) );
  CFA1X1 U986 ( .A(n1876), .B(n1851), .CI(n2059), .CO(n1052), .S(n1053) );
  CFA1X1 U988 ( .A(n1789), .B(n1999), .CI(n3584), .CO(n1056), .S(n1057) );
  CFA1X1 U991 ( .A(n1069), .B(n1067), .CI(n1090), .CO(n1062), .S(n1063) );
  CFA1X1 U992 ( .A(n1094), .B(n1092), .CI(n1071), .CO(n1064), .S(n1065) );
  CFA1X1 U995 ( .A(n1104), .B(n1098), .CI(n1100), .CO(n1070), .S(n1071) );
  CFA1X1 U996 ( .A(n1938), .B(n1081), .CI(n1907), .CO(n1072), .S(n1073) );
  CFA1X1 U997 ( .A(n1969), .B(n1852), .CI(n1821), .CO(n1074), .S(n1075) );
  CFA1X1 U998 ( .A(n1790), .B(n2000), .CI(n1759), .CO(n1076), .S(n1077) );
  CFA1X1 U999 ( .A(n1877), .B(n2060), .CI(n2091), .CO(n1078), .S(n1079) );
  CFA1X1 U1006 ( .A(n1103), .B(n1105), .CI(n1099), .CO(n1092), .S(n1093) );
  CFA1X1 U1009 ( .A(n1760), .B(n2123), .CI(n1853), .CO(n1098), .S(n1099) );
  CFA1X1 U1010 ( .A(n1878), .B(n2001), .CI(n1822), .CO(n1100), .S(n1101) );
  CFA1X1 U1011 ( .A(n1791), .B(n2030), .CI(n1970), .CO(n1102), .S(n1103) );
  CFA1X1 U1020 ( .A(n1131), .B(n1154), .CI(n1156), .CO(n1120), .S(n1121) );
  CFA1X1 U1024 ( .A(n1940), .B(n2031), .CI(n2124), .CO(n1128), .S(n1129) );
  CFA1X1 U1034 ( .A(n2094), .B(n1972), .CI(n1855), .CO(n1148), .S(n1149) );
  CFA1X1 U1037 ( .A(n1910), .B(n1941), .CI(n2032), .CO(n1154), .S(n1155) );
  CFA1X1 U1060 ( .A(n1234), .B(n1232), .CI(n1238), .CO(n1200), .S(n1201) );
  CFA1X1 U1062 ( .A(n1795), .B(n1974), .CI(n1764), .CO(n1204), .S(n1205) );
  CFA1X1 U1074 ( .A(n1266), .B(n1262), .CI(n1264), .CO(n1228), .S(n1229) );
  CFA1X1 U1079 ( .A(n2097), .B(n2066), .CI(n1882), .CO(n1238), .S(n1239) );
  CFA1X1 U1089 ( .A(n1296), .B(n1292), .CI(n1294), .CO(n1258), .S(n1259) );
  CFA1X1 U1090 ( .A(n1273), .B(n1298), .CI(n1300), .CO(n1260), .S(n1261) );
  CFA1X1 U1095 ( .A(n2159), .B(n2007), .CI(n1976), .CO(n1270), .S(n1271) );
  COR2X1 U1097 ( .A(n2189), .B(n1883), .Z(n1272) );
  CFA1X1 U1102 ( .A(n1318), .B(n1316), .CI(n1291), .CO(n1282), .S(n1283) );
  CFA1X1 U1105 ( .A(n1322), .B(n1326), .CI(n1324), .CO(n1288), .S(n1289) );
  CFA1X1 U1107 ( .A(n1724), .B(n1977), .CI(n1798), .CO(n1292), .S(n1293) );
  CFA1X1 U1108 ( .A(n1767), .B(n1829), .CI(n1915), .CO(n1294), .S(n1295) );
  CFA1X1 U1109 ( .A(n2068), .B(n2008), .CI(n2037), .CO(n1296), .S(n1297) );
  CFA1X1 U1110 ( .A(n2130), .B(n2190), .CI(n2099), .CO(n1298), .S(n1299) );
  CFA1X1 U1111 ( .A(n2160), .B(n1860), .CI(n1946), .CO(n1300), .S(n1301) );
  CHA1X1 U1112 ( .A(n2221), .B(n1884), .CO(n1302), .S(n1303) );
  CFA1X1 U1121 ( .A(n2100), .B(n1356), .CI(n3255), .CO(n1320), .S(n1321) );
  CFA1X1 U1122 ( .A(n2131), .B(n2009), .CI(n2069), .CO(n1322), .S(n1323) );
  CFA1X1 U1123 ( .A(n1916), .B(n1978), .CI(n1947), .CO(n1324), .S(n1325) );
  CFA1X1 U1125 ( .A(n1799), .B(n2191), .CI(n2222), .CO(n1328), .S(n1329) );
  CFA1X1 U1126 ( .A(n1768), .B(n2161), .CI(n2038), .CO(n1330), .S(n1331) );
  CFA1X1 U1128 ( .A(n1339), .B(n1364), .CI(n1341), .CO(n1334), .S(n1335) );
  CFA1X1 U1135 ( .A(n2101), .B(n1359), .CI(n2070), .CO(n1348), .S(n1349) );
  CFA1X1 U1136 ( .A(n2132), .B(n2010), .CI(n1979), .CO(n1350), .S(n1351) );
  CFA1X1 U1138 ( .A(n1831), .B(n1862), .CI(n2039), .CO(n1354), .S(n1355) );
  CFA1X1 U1139 ( .A(n2223), .B(n1948), .CI(n1886), .CO(n1356), .S(n1357) );
  CFA1X1 U1143 ( .A(n1371), .B(n1369), .CI(n1394), .CO(n1364), .S(n1365) );
  CFA1X1 U1149 ( .A(n2102), .B(n2011), .CI(n2071), .CO(n1376), .S(n1377) );
  CFA1X1 U1150 ( .A(n2133), .B(n1980), .CI(n1949), .CO(n1378), .S(n1379) );
  CFA1X1 U1152 ( .A(n2224), .B(n1832), .CI(n2193), .CO(n1382), .S(n1383) );
  CFA1X1 U1156 ( .A(n1420), .B(n1418), .CI(n1397), .CO(n1390), .S(n1391) );
  CFA1X1 U1163 ( .A(n1888), .B(n1919), .CI(n2103), .CO(n1404), .S(n1405) );
  CFA1X1 U1165 ( .A(n2164), .B(n1833), .CI(n2225), .CO(n1408), .S(n1409) );
  CHA1X1 U1166 ( .A(n2041), .B(n1726), .CO(n1410), .S(n1411) );
  CFA1X1 U1171 ( .A(n1431), .B(n1427), .CI(n1429), .CO(n1420), .S(n1421) );
  CFA1X1 U1174 ( .A(n2135), .B(n1458), .CI(n2104), .CO(n1426), .S(n1427) );
  CFA1X1 U1178 ( .A(n1834), .B(n2165), .CI(n1889), .CO(n1434), .S(n1435) );
  CFA1X1 U1187 ( .A(n2196), .B(n2014), .CI(n1952), .CO(n1452), .S(n1453) );
  CFA1X1 U1188 ( .A(n2043), .B(n1866), .CI(n1921), .CO(n1454), .S(n1455) );
  CFA1X1 U1194 ( .A(n1494), .B(n1473), .CI(n1492), .CO(n1466), .S(n1467) );
  CFA1X1 U1197 ( .A(n2106), .B(n1500), .CI(n3758), .CO(n1472), .S(n1473) );
  CFA1X1 U1198 ( .A(n2137), .B(n2015), .CI(n2075), .CO(n1474), .S(n1475) );
  CFA1X1 U1201 ( .A(n1867), .B(n1891), .CI(n2167), .CO(n1480), .S(n1481) );
  CFA1X1 U1205 ( .A(n1514), .B(n1495), .CI(n1501), .CO(n1488), .S(n1489) );
  CFA1X1 U1208 ( .A(n1892), .B(n1503), .CI(n1985), .CO(n1494), .S(n1495) );
  CFA1X1 U1209 ( .A(n1954), .B(n2198), .CI(n1923), .CO(n1496), .S(n1497) );
  CFA1X1 U1210 ( .A(n2168), .B(n2016), .CI(n2229), .CO(n1498), .S(n1499) );
  CFA1X1 U1215 ( .A(n1532), .B(n1530), .CI(n1515), .CO(n1508), .S(n1509) );
  CFA1X1 U1219 ( .A(n2139), .B(n2108), .CI(n2077), .CO(n1516), .S(n1517) );
  CFA1X1 U1220 ( .A(n2230), .B(n2017), .CI(n1986), .CO(n1518), .S(n1519) );
  CFA1X1 U1222 ( .A(n1893), .B(n2199), .CI(n2169), .CO(n1522), .S(n1523) );
  CFA1X1 U1225 ( .A(n1552), .B(n1550), .CI(n1535), .CO(n1528), .S(n1529) );
  CFA1X1 U1236 ( .A(n1561), .B(n1557), .CI(n1559), .CO(n1550), .S(n1551) );
  CFA1X1 U1239 ( .A(n2232), .B(n2079), .CI(n2019), .CO(n1556), .S(n1557) );
  CFA1X1 U1246 ( .A(n1594), .B(n1592), .CI(n1579), .CO(n1570), .S(n1571) );
  CFA1X1 U1247 ( .A(n2142), .B(n2080), .CI(n2111), .CO(n1572), .S(n1573) );
  CFA1X1 U1249 ( .A(n1958), .B(n1989), .CI(n2202), .CO(n1576), .S(n1577) );
  CFA1X1 U1253 ( .A(n1591), .B(n1602), .CI(n1604), .CO(n1584), .S(n1585) );
  CFA1X1 U1255 ( .A(n2143), .B(n1608), .CI(n1610), .CO(n1588), .S(n1589) );
  CFA1X1 U1256 ( .A(n2234), .B(n2112), .CI(n2081), .CO(n1590), .S(n1591) );
  CFA1X1 U1258 ( .A(n1959), .B(n2203), .CI(n2173), .CO(n1594), .S(n1595) );
  CFA1X1 U1261 ( .A(n1609), .B(n1618), .CI(n1607), .CO(n1600), .S(n1601) );
  CFA1X1 U1263 ( .A(n3292), .B(n1611), .CI(n2022), .CO(n1604), .S(n1605) );
  CFA1X1 U1264 ( .A(n2113), .B(n1991), .CI(n2051), .CO(n1606), .S(n1607) );
  CFA1X1 U1265 ( .A(n2204), .B(n4503), .CI(n2235), .CO(n1608), .S(n1609) );
  CFA1X1 U1268 ( .A(n1632), .B(n1630), .CI(n1619), .CO(n1614), .S(n1615) );
  CFA1X1 U1271 ( .A(n2236), .B(n2145), .CI(n2114), .CO(n1620), .S(n1621) );
  CFA1X1 U1272 ( .A(n2175), .B(n2023), .CI(n2083), .CO(n1622), .S(n1623) );
  CFA1X1 U1276 ( .A(n1648), .B(n1635), .CI(n1646), .CO(n1630), .S(n1631) );
  CFA1X1 U1277 ( .A(n2115), .B(n1650), .CI(n1639), .CO(n1632), .S(n1633) );
  CFA1X1 U1281 ( .A(n1645), .B(n1643), .CI(n1654), .CO(n1640), .S(n1641) );
  CFA1X1 U1282 ( .A(n1649), .B(n1656), .CI(n1647), .CO(n1642), .S(n1643) );
  CFA1X1 U1283 ( .A(n1660), .B(n1651), .CI(n1658), .CO(n1644), .S(n1645) );
  CFA1X1 U1285 ( .A(n2207), .B(n2116), .CI(n2085), .CO(n1648), .S(n1649) );
  CFA1X1 U1286 ( .A(n2025), .B(n2054), .CI(n2177), .CO(n1650), .S(n1651) );
  CFA1X1 U1287 ( .A(n1657), .B(n1655), .CI(n1666), .CO(n1652), .S(n1653) );
  CFA1X1 U1288 ( .A(n1661), .B(n1668), .CI(n1659), .CO(n1654), .S(n1655) );
  CFA1X1 U1290 ( .A(n2178), .B(n2086), .CI(n2055), .CO(n1658), .S(n1659) );
  CFA1X1 U1291 ( .A(n2208), .B(n2117), .CI(n2239), .CO(n1660), .S(n1661) );
  CHA1X1 U1292 ( .A(n1733), .B(n2148), .CO(n1662), .S(n1663) );
  CFA1X1 U1293 ( .A(n1676), .B(n1667), .CI(n1669), .CO(n1664), .S(n1665) );
  CFA1X1 U1295 ( .A(n2149), .B(n1680), .CI(n1682), .CO(n1668), .S(n1669) );
  CFA1X1 U1296 ( .A(n2240), .B(n2118), .CI(n2087), .CO(n1670), .S(n1671) );
  CFA1X1 U1298 ( .A(n1679), .B(n1677), .CI(n1686), .CO(n1674), .S(n1675) );
  CFA1X1 U1299 ( .A(n1690), .B(n1681), .CI(n1688), .CO(n1676), .S(n1677) );
  CFA1X1 U1301 ( .A(n2241), .B(n2180), .CI(n2088), .CO(n1680), .S(n1681) );
  CFA1X1 U1305 ( .A(n2242), .B(n2151), .CI(n2120), .CO(n1688), .S(n1689) );
  CFA1X1 U1306 ( .A(n2089), .B(n2181), .CI(n2211), .CO(n1690), .S(n1691) );
  CFA1X1 U1307 ( .A(n1702), .B(n1695), .CI(n1697), .CO(n1692), .S(n1693) );
  CFA1X1 U1308 ( .A(n2243), .B(n1704), .CI(n1699), .CO(n1694), .S(n1695) );
  CFA1X1 U1309 ( .A(n2182), .B(n2152), .CI(n2121), .CO(n1696), .S(n1697) );
  CFA1X1 U1311 ( .A(n1708), .B(n1703), .CI(n1705), .CO(n1700), .S(n1701) );
  CFA1X1 U1312 ( .A(n2244), .B(n1710), .CI(n2153), .CO(n1702), .S(n1703) );
  CFA1X1 U1313 ( .A(n2122), .B(n2213), .CI(n2183), .CO(n1704), .S(n1705) );
  CFA1X1 U1314 ( .A(n1711), .B(n1709), .CI(n1714), .CO(n1706), .S(n1707) );
  CHA1X1 U1316 ( .A(n2214), .B(n1736), .CO(n1710), .S(n1711) );
  CFA1X1 U1317 ( .A(n2246), .B(n1715), .CI(n1718), .CO(n1712), .S(n1713) );
  CFA1X1 U1318 ( .A(n2155), .B(n4459), .CI(n2215), .CO(n1714), .S(n1715) );
  CFA1X1 U1319 ( .A(n2216), .B(n1719), .CI(n2186), .CO(n1716), .S(n1717) );
  CHA1X1 U1320 ( .A(n1737), .B(n2247), .CO(n1718), .S(n1719) );
  CFA1X1 U1321 ( .A(n3745), .B(n2217), .CI(n2248), .CO(n1720), .S(n1721) );
  COND2X1 U1323 ( .A(n144), .B(n4604), .C(n2284), .D(n3277), .Z(n1724) );
  COND2X1 U1332 ( .A(n4511), .B(n2260), .C(n2259), .D(n3277), .Z(n1744) );
  COND2X1 U1333 ( .A(n4511), .B(n2261), .C(n2260), .D(n3277), .Z(n1745) );
  COND2X1 U1335 ( .A(n4511), .B(n2263), .C(n2262), .D(n3277), .Z(n1747) );
  COND2X1 U1336 ( .A(n4511), .B(n2264), .C(n2263), .D(n3277), .Z(n1748) );
  COND2X1 U1337 ( .A(n4511), .B(n2265), .C(n2264), .D(n3277), .Z(n1749) );
  COND2X1 U1338 ( .A(n4511), .B(n2266), .C(n2265), .D(n3277), .Z(n1750) );
  COND2X1 U1339 ( .A(n4511), .B(n2267), .C(n2266), .D(n3277), .Z(n1751) );
  COND2X1 U1340 ( .A(n4511), .B(n2268), .C(n2267), .D(n3277), .Z(n1752) );
  COND2X1 U1341 ( .A(n4511), .B(n2269), .C(n2268), .D(n3277), .Z(n1753) );
  COND2X1 U1342 ( .A(n4511), .B(n2270), .C(n2269), .D(n3277), .Z(n1754) );
  COND2X1 U1343 ( .A(n4511), .B(n2271), .C(n2270), .D(n3277), .Z(n1755) );
  COND2X1 U1344 ( .A(n4511), .B(n2272), .C(n2271), .D(n3277), .Z(n1756) );
  COND2X1 U1345 ( .A(n4511), .B(n2273), .C(n2272), .D(n3277), .Z(n1757) );
  COND2X1 U1346 ( .A(n144), .B(n2274), .C(n2273), .D(n3277), .Z(n1758) );
  COND2X1 U1347 ( .A(n4511), .B(n2275), .C(n2274), .D(n3277), .Z(n1759) );
  COND2X1 U1348 ( .A(n4511), .B(n2276), .C(n2275), .D(n3277), .Z(n1760) );
  COND2X1 U1349 ( .A(n4511), .B(n2277), .C(n2276), .D(n3277), .Z(n1761) );
  COND2X1 U1350 ( .A(n144), .B(n2278), .C(n2277), .D(n3277), .Z(n1762) );
  COND2X1 U1352 ( .A(n144), .B(n2280), .C(n3277), .D(n2279), .Z(n1764) );
  COND2X1 U1354 ( .A(n144), .B(n2282), .C(n2281), .D(net16497), .Z(n1766) );
  COND2X1 U1396 ( .A(net18310), .B(n2290), .C(net16438), .D(n2289), .Z(n1774)
         );
  COND2X1 U1401 ( .A(net18310), .B(n2295), .C(net16438), .D(n2294), .Z(n1779)
         );
  COND2X1 U1402 ( .A(net18310), .B(n2296), .C(net16438), .D(n2295), .Z(n1780)
         );
  COND2X1 U1404 ( .A(net18310), .B(n2298), .C(net16438), .D(n2297), .Z(n1782)
         );
  COND2X1 U1406 ( .A(net18310), .B(n2300), .C(net16438), .D(n2299), .Z(n1784)
         );
  COND2X1 U1407 ( .A(net18310), .B(n2301), .C(net16439), .D(n2300), .Z(n1785)
         );
  COND2X1 U1409 ( .A(net18310), .B(n2303), .C(net16438), .D(n2302), .Z(n1787)
         );
  COND2X1 U1410 ( .A(net18310), .B(n2304), .C(net16439), .D(n2303), .Z(n1788)
         );
  COND2X1 U1411 ( .A(net18310), .B(n2305), .C(net16438), .D(n2304), .Z(n1789)
         );
  COND2X1 U1412 ( .A(net18310), .B(n2306), .C(net16439), .D(n2305), .Z(n1790)
         );
  COND2X1 U1413 ( .A(net18310), .B(n2307), .C(net16438), .D(n2306), .Z(n1791)
         );
  COND2X1 U1414 ( .A(net18310), .B(n2308), .C(net16438), .D(n2307), .Z(n1792)
         );
  COND2X1 U1417 ( .A(net18310), .B(n2311), .C(net16438), .D(n2310), .Z(n1795)
         );
  COND2X1 U1419 ( .A(n135), .B(n2313), .C(net16439), .D(n2312), .Z(n1797) );
  COND2X1 U1420 ( .A(net18310), .B(n2314), .C(net16438), .D(n2313), .Z(n1798)
         );
  COND2X1 U1462 ( .A(net17738), .B(n2322), .C(n123), .D(n2321), .Z(n1806) );
  COND2X1 U1465 ( .A(net17738), .B(n2325), .C(n123), .D(n2324), .Z(n1809) );
  COND2X1 U1466 ( .A(net17738), .B(n2326), .C(n123), .D(n2325), .Z(n1810) );
  COND2X1 U1467 ( .A(net17738), .B(n2327), .C(n123), .D(n2326), .Z(n1811) );
  COND2X1 U1468 ( .A(net17738), .B(n2328), .C(n123), .D(n2327), .Z(n1812) );
  COND2X1 U1469 ( .A(net17738), .B(n2329), .C(n123), .D(n2328), .Z(n1813) );
  COND2X1 U1471 ( .A(net17738), .B(n2331), .C(n123), .D(n2330), .Z(n1815) );
  COND2X1 U1472 ( .A(net17738), .B(n2332), .C(n123), .D(n2331), .Z(n1816) );
  COND2X1 U1473 ( .A(net17738), .B(n2333), .C(n123), .D(n2332), .Z(n1817) );
  COND2X1 U1474 ( .A(net17738), .B(n2334), .C(n123), .D(n2333), .Z(n1818) );
  COND2X1 U1475 ( .A(net17738), .B(n2335), .C(n123), .D(n2334), .Z(n1819) );
  COND2X1 U1476 ( .A(net17738), .B(n2336), .C(n123), .D(n2335), .Z(n1820) );
  COND2X1 U1477 ( .A(net17738), .B(n2337), .C(n123), .D(n2336), .Z(n1821) );
  COND2X1 U1478 ( .A(net17738), .B(n2338), .C(n123), .D(n2337), .Z(n1822) );
  COND2X1 U1479 ( .A(net17738), .B(n2339), .C(n123), .D(n2338), .Z(n1823) );
  COND2X1 U1483 ( .A(net17738), .B(n2343), .C(n123), .D(n2342), .Z(n1827) );
  COND2X1 U1484 ( .A(net17738), .B(n2344), .C(n123), .D(n2343), .Z(n1828) );
  COND2X1 U1485 ( .A(net17738), .B(n2345), .C(n123), .D(n2344), .Z(n1829) );
  COND2X1 U1486 ( .A(net17738), .B(n2346), .C(n123), .D(n2345), .Z(n1830) );
  COND2X1 U1487 ( .A(net17738), .B(n2347), .C(n123), .D(n2346), .Z(n1831) );
  COND2X1 U1489 ( .A(net17738), .B(n2349), .C(n123), .D(n2348), .Z(n1833) );
  COND2X1 U1524 ( .A(net18628), .B(n4281), .C(n2383), .D(net16433), .Z(n1727)
         );
  COND2X1 U1526 ( .A(net18628), .B(n2352), .C(n3667), .D(n2351), .Z(n1836) );
  COND2X1 U1527 ( .A(n117), .B(n2353), .C(n3667), .D(n2352), .Z(n1837) );
  COND2X1 U1530 ( .A(net18628), .B(n2356), .C(n3667), .D(n2355), .Z(n1840) );
  COND2X1 U1531 ( .A(net18628), .B(n2357), .C(n3667), .D(n2356), .Z(n1841) );
  COND2X1 U1532 ( .A(n117), .B(n2358), .C(net16433), .D(n2357), .Z(n1842) );
  COND2X1 U1533 ( .A(net18628), .B(n2359), .C(net16433), .D(n2358), .Z(n1843)
         );
  COND2X1 U1534 ( .A(n117), .B(n2360), .C(n3667), .D(n2359), .Z(n1844) );
  COND2X1 U1535 ( .A(net18628), .B(n2361), .C(net16433), .D(n2360), .Z(n1845)
         );
  COND2X1 U1536 ( .A(net18628), .B(n2362), .C(net16433), .D(n2361), .Z(n1846)
         );
  COND2X1 U1537 ( .A(net18628), .B(n2363), .C(net16433), .D(n2362), .Z(n1847)
         );
  COND2X1 U1538 ( .A(n117), .B(n2364), .C(net16433), .D(n2363), .Z(n1848) );
  COND2X1 U1539 ( .A(n117), .B(n2365), .C(net16433), .D(n2364), .Z(n1849) );
  COND2X1 U1540 ( .A(net18628), .B(n2366), .C(n3667), .D(n2365), .Z(n1850) );
  COND2X1 U1541 ( .A(n117), .B(n2367), .C(net16433), .D(n2366), .Z(n1851) );
  COND2X1 U1542 ( .A(n117), .B(n2368), .C(net16433), .D(n2367), .Z(n1852) );
  COND2X1 U1543 ( .A(net18628), .B(n2369), .C(net16433), .D(n2368), .Z(n1853)
         );
  COND2X1 U1544 ( .A(n117), .B(n2370), .C(net16433), .D(n2369), .Z(n1854) );
  COND2X1 U1547 ( .A(net18628), .B(n2373), .C(net16433), .D(n2372), .Z(n1857)
         );
  COND2X1 U1548 ( .A(n117), .B(n2374), .C(net16433), .D(n2373), .Z(n1858) );
  COND2X1 U1549 ( .A(n117), .B(n2375), .C(net16433), .D(n2374), .Z(n1859) );
  COND2X1 U1550 ( .A(n117), .B(n2376), .C(net16433), .D(n2375), .Z(n1860) );
  COND2X1 U1552 ( .A(net18628), .B(n2378), .C(net16433), .D(n2377), .Z(n1862)
         );
  COND2X1 U1553 ( .A(n117), .B(n2379), .C(net16433), .D(n2378), .Z(n1863) );
  COND2X1 U1554 ( .A(n117), .B(n2380), .C(net16433), .D(n2379), .Z(n1864) );
  COND2X1 U1556 ( .A(net18628), .B(n2382), .C(net16433), .D(n2381), .Z(n1866)
         );
  COND2X1 U1599 ( .A(n3301), .B(n2391), .C(net17425), .D(n2390), .Z(n920) );
  COND2X1 U1601 ( .A(net17727), .B(n2393), .C(n2392), .D(net17425), .Z(n954)
         );
  COND2X1 U1602 ( .A(n4013), .B(n2394), .C(n2393), .D(net17425), .Z(n1873) );
  COND2X1 U1603 ( .A(n4013), .B(n2395), .C(n2394), .D(net16426), .Z(n1874) );
  COND2X1 U1604 ( .A(n4012), .B(n2396), .C(n2395), .D(net16426), .Z(n1875) );
  COND2X1 U1605 ( .A(n3302), .B(n2397), .C(n2396), .D(net16426), .Z(n1034) );
  COND2X1 U1606 ( .A(n3301), .B(n2398), .C(n2397), .D(net16426), .Z(n1876) );
  COND2X1 U1608 ( .A(n4012), .B(n2400), .C(n2399), .D(net16426), .Z(n1878) );
  COND2X1 U1619 ( .A(n2411), .B(net17727), .C(n2410), .D(net16426), .Z(n1888)
         );
  COND2X1 U1620 ( .A(n3301), .B(n2412), .C(net16426), .D(n2411), .Z(n1889) );
  COND2X1 U1660 ( .A(net18627), .B(n2418), .C(n4508), .D(n2417), .Z(n1895) );
  COND2X1 U1661 ( .A(net18627), .B(n2419), .C(n3891), .D(n2418), .Z(n1896) );
  COND2X1 U1662 ( .A(net18627), .B(n2420), .C(n3891), .D(n2419), .Z(n1897) );
  COND2X1 U1663 ( .A(net18627), .B(n2421), .C(n4508), .D(n2420), .Z(n1898) );
  COND2X1 U1664 ( .A(net18627), .B(n2422), .C(n3891), .D(n2421), .Z(n1899) );
  COND2X1 U1665 ( .A(net18627), .B(n2423), .C(n3891), .D(n2422), .Z(n1900) );
  COND2X1 U1666 ( .A(net18627), .B(n2424), .C(n4508), .D(n2423), .Z(n1901) );
  COND2X1 U1667 ( .A(net18627), .B(n2425), .C(n3891), .D(n2424), .Z(n1902) );
  COND2X1 U1668 ( .A(net18627), .B(n2426), .C(n4508), .D(n2425), .Z(n1903) );
  COND2X1 U1669 ( .A(net18627), .B(n2427), .C(n3891), .D(n2426), .Z(n1904) );
  COND2X1 U1670 ( .A(net18627), .B(n2428), .C(n3891), .D(n2427), .Z(n1905) );
  COND2X1 U1671 ( .A(net18627), .B(n2429), .C(n4508), .D(n2428), .Z(n1906) );
  COND2X1 U1672 ( .A(net18627), .B(n2430), .C(n3891), .D(n2429), .Z(n1907) );
  COND2X1 U1673 ( .A(n99), .B(n2431), .C(n3891), .D(n2430), .Z(n1908) );
  COND2X1 U1674 ( .A(n99), .B(n2432), .C(n3771), .D(n2431), .Z(n1909) );
  COND2X1 U1675 ( .A(n99), .B(n2433), .C(net16416), .D(n2432), .Z(n1910) );
  COND2X1 U1678 ( .A(net18627), .B(n2436), .C(n3771), .D(n2435), .Z(n1913) );
  COND2X1 U1679 ( .A(net18627), .B(n2437), .C(n4508), .D(n2436), .Z(n1914) );
  COND2X1 U1680 ( .A(n99), .B(n2438), .C(n2437), .D(net16416), .Z(n1915) );
  COND2X1 U1681 ( .A(n99), .B(n2439), .C(n4508), .D(n2438), .Z(n1916) );
  COND2X1 U1682 ( .A(net18627), .B(n2440), .C(n3891), .D(n2439), .Z(n1917) );
  COND2X1 U1683 ( .A(net18627), .B(n2441), .C(n3891), .D(n2440), .Z(n1918) );
  COND2X1 U1684 ( .A(net18627), .B(n2442), .C(n4508), .D(n2441), .Z(n1919) );
  COND2X1 U1685 ( .A(net18627), .B(n2443), .C(n4508), .D(n2442), .Z(n1920) );
  COND2X1 U1686 ( .A(net18627), .B(n2444), .C(n3891), .D(n2443), .Z(n1921) );
  COND2X1 U1687 ( .A(n99), .B(n2445), .C(n2444), .D(n4508), .Z(n1922) );
  COND2X1 U1688 ( .A(n99), .B(n2446), .C(n3891), .D(n2445), .Z(n1923) );
  COND2X1 U1689 ( .A(net18627), .B(n2447), .C(n3771), .D(n2446), .Z(n1924) );
  COND2X1 U1690 ( .A(n99), .B(n2448), .C(n3771), .D(n2447), .Z(n1925) );
  COND2X1 U1727 ( .A(n3991), .B(n2451), .C(net16511), .D(n2450), .Z(n1928) );
  COND2X1 U1728 ( .A(n3991), .B(n2452), .C(net16512), .D(n2451), .Z(n1929) );
  COND2X1 U1731 ( .A(n90), .B(n2455), .C(net16511), .D(n2454), .Z(n1932) );
  COND2X1 U1733 ( .A(n3991), .B(n2457), .C(net16512), .D(n2456), .Z(n1934) );
  COND2X1 U1735 ( .A(n3991), .B(n2459), .C(net16511), .D(n2458), .Z(n1936) );
  COND2X1 U1737 ( .A(n3991), .B(n2461), .C(net16511), .D(n2460), .Z(n1938) );
  COND2X1 U1740 ( .A(n90), .B(n2464), .C(net16512), .D(n2463), .Z(n1941) );
  COND2X1 U1742 ( .A(n90), .B(n2466), .C(net16511), .D(n2465), .Z(n1943) );
  COND2X1 U1743 ( .A(n3991), .B(n2467), .C(net16512), .D(n2466), .Z(n1944) );
  COND2X1 U1745 ( .A(n2469), .B(n90), .C(net16511), .D(n2468), .Z(n1946) );
  COND2X1 U1746 ( .A(n3991), .B(n2470), .C(net16512), .D(n2469), .Z(n1947) );
  COND2X1 U1747 ( .A(n90), .B(n2471), .C(net16512), .D(n2470), .Z(n1948) );
  COND2X1 U1748 ( .A(n3991), .B(n2472), .C(net16512), .D(n2471), .Z(n1949) );
  COND2X1 U1749 ( .A(n90), .B(n2473), .C(net16511), .D(n2472), .Z(n1950) );
  COND2X1 U1750 ( .A(n3991), .B(n2474), .C(net16511), .D(n2473), .Z(n1951) );
  COND2X1 U1751 ( .A(n90), .B(n2475), .C(net16511), .D(n2474), .Z(n1952) );
  COND2X1 U1752 ( .A(n3991), .B(n2476), .C(net16512), .D(n2475), .Z(n1953) );
  COND2X1 U1753 ( .A(n3991), .B(n2477), .C(net16511), .D(n2476), .Z(n1954) );
  COND2X1 U1755 ( .A(n3991), .B(n2479), .C(net16511), .D(n2478), .Z(n1956) );
  COND2X1 U1757 ( .A(n3991), .B(n2481), .C(net16511), .D(n2480), .Z(n1958) );
  COND2X1 U1794 ( .A(n4120), .B(n2484), .C(net16413), .D(n2483), .Z(n1961) );
  COND2X1 U1795 ( .A(n4120), .B(n2485), .C(n4217), .D(n2484), .Z(n1962) );
  COND2X1 U1798 ( .A(n81), .B(n2488), .C(n4217), .D(n2487), .Z(n1965) );
  COND2X1 U1799 ( .A(n81), .B(n2489), .C(n4217), .D(n2488), .Z(n1966) );
  COND2X1 U1800 ( .A(n81), .B(n2490), .C(n4217), .D(n2489), .Z(n1967) );
  COND2X1 U1802 ( .A(n4120), .B(n2492), .C(net16413), .D(n2491), .Z(n1969) );
  COND2X1 U1803 ( .A(n4120), .B(n2493), .C(net16413), .D(n2492), .Z(n1970) );
  COND2X1 U1804 ( .A(n4120), .B(n2494), .C(net16413), .D(n2493), .Z(n1971) );
  COND2X1 U1805 ( .A(n81), .B(n2495), .C(n4217), .D(n2494), .Z(n1972) );
  COND2X1 U1807 ( .A(n81), .B(n2497), .C(n4217), .D(n2496), .Z(n1974) );
  COND2X1 U1808 ( .A(n4120), .B(n2498), .C(n2497), .D(n78), .Z(n1975) );
  COND2X1 U1809 ( .A(n81), .B(n2499), .C(net16413), .D(n2498), .Z(n1976) );
  COND2X1 U1810 ( .A(n81), .B(n2500), .C(net16413), .D(n2499), .Z(n1977) );
  COND2X1 U1811 ( .A(n4120), .B(n2501), .C(net16413), .D(n2500), .Z(n1978) );
  COND2X1 U1812 ( .A(n4120), .B(n2502), .C(net16413), .D(n2501), .Z(n1979) );
  COND2X1 U1813 ( .A(n4120), .B(n2503), .C(net16413), .D(n2502), .Z(n1980) );
  COND2X1 U1814 ( .A(n81), .B(n2504), .C(net16413), .D(n2503), .Z(n1981) );
  COND2X1 U1815 ( .A(n4120), .B(n2505), .C(net16413), .D(n2504), .Z(n1982) );
  COND2X1 U1816 ( .A(n4120), .B(n2506), .C(net16413), .D(n2505), .Z(n1983) );
  COND2X1 U1818 ( .A(n4120), .B(n2508), .C(n4217), .D(n2507), .Z(n1985) );
  COND2X1 U1819 ( .A(n81), .B(n2509), .C(net16413), .D(n2508), .Z(n1986) );
  COND2X1 U1820 ( .A(n81), .B(n2510), .C(n4217), .D(n2509), .Z(n1987) );
  COND2X1 U1822 ( .A(n4120), .B(n2512), .C(n4217), .D(n2511), .Z(n1989) );
  COND2X1 U1824 ( .A(n81), .B(n2514), .C(n4217), .D(n2513), .Z(n1991) );
  COND2X1 U1862 ( .A(n2518), .B(net17279), .C(n3122), .D(n2517), .Z(n1995) );
  COND2X1 U1863 ( .A(n2519), .B(n3117), .C(n3121), .D(n2518), .Z(n1996) );
  COND2X1 U1864 ( .A(net17279), .B(n2520), .C(n3122), .D(n2519), .Z(n1997) );
  COND2X1 U1865 ( .A(n3117), .B(n2521), .C(n3121), .D(n2520), .Z(n1998) );
  COND2X1 U1866 ( .A(n2522), .B(n3113), .C(n3122), .D(n2521), .Z(n1999) );
  COND2X1 U1867 ( .A(n3117), .B(n2523), .C(n3121), .D(n2522), .Z(n2000) );
  COND2X1 U1868 ( .A(net17279), .B(n2524), .C(n3122), .D(n2523), .Z(n2001) );
  COND2X1 U1869 ( .A(net16301), .B(n2525), .C(net16465), .D(n2524), .Z(n2002)
         );
  COND2X1 U1873 ( .A(net17278), .B(n2529), .C(net16465), .D(n2528), .Z(n2006)
         );
  COND2X1 U1874 ( .A(n3117), .B(n2530), .C(n3121), .D(n2529), .Z(n2007) );
  COND2X1 U1875 ( .A(n3142), .B(n2531), .C(n3121), .D(n2530), .Z(n2008) );
  COND2X1 U1876 ( .A(net16301), .B(n2532), .C(net16465), .D(n2531), .Z(n2009)
         );
  COND2X1 U1877 ( .A(n3133), .B(n2533), .C(n3122), .D(n2532), .Z(n2010) );
  COND2X1 U1878 ( .A(n2534), .B(net17278), .C(net16465), .D(n2533), .Z(n2011)
         );
  COND2X1 U1880 ( .A(net17278), .B(n2536), .C(n3121), .D(n2535), .Z(n2013) );
  COND2X1 U1881 ( .A(net17278), .B(n2537), .C(net16465), .D(n2536), .Z(n2014)
         );
  COND2X1 U1882 ( .A(n3117), .B(n2538), .C(n3122), .D(n2537), .Z(n2015) );
  COND2X1 U1883 ( .A(n3117), .B(n2539), .C(n3122), .D(n2538), .Z(n2016) );
  COND2X1 U1884 ( .A(n3117), .B(n2540), .C(n3122), .D(n2539), .Z(n2017) );
  COND2X1 U1886 ( .A(net16301), .B(n2542), .C(net16465), .D(n2541), .Z(n2019)
         );
  COND2X1 U1887 ( .A(n3117), .B(n2543), .C(n3121), .D(n2542), .Z(n2020) );
  COND2X1 U1888 ( .A(net17279), .B(n2544), .C(n3122), .D(n2543), .Z(n2021) );
  COND2X1 U1890 ( .A(net17279), .B(n2546), .C(n3121), .D(n2545), .Z(n2023) );
  COND2X1 U1928 ( .A(n63), .B(n2550), .C(n2549), .D(n4505), .Z(n992) );
  COND2X1 U1929 ( .A(n63), .B(n2551), .C(n2550), .D(n4505), .Z(n2027) );
  COND2X1 U1930 ( .A(n63), .B(n2552), .C(n2551), .D(n4505), .Z(n2028) );
  COND2X1 U1931 ( .A(n63), .B(n2553), .C(n4505), .D(n2552), .Z(n2029) );
  COND2X1 U1933 ( .A(n63), .B(n2555), .C(n2554), .D(n4505), .Z(n2030) );
  COND2X1 U1934 ( .A(n63), .B(n3269), .C(n2555), .D(n4505), .Z(n2031) );
  COND2X1 U1936 ( .A(n63), .B(n2558), .C(n2557), .D(n4505), .Z(n2033) );
  COND2X1 U1937 ( .A(n63), .B(n2559), .C(n2558), .D(n4505), .Z(n2034) );
  COND2X1 U1938 ( .A(n63), .B(n2560), .C(n2559), .D(n4505), .Z(n2035) );
  COND2X1 U1940 ( .A(n63), .B(n2562), .C(n2561), .D(n4505), .Z(n2037) );
  COND2X1 U1942 ( .A(n4316), .B(n2564), .C(n2563), .D(n4505), .Z(n2039) );
  COND2X1 U1945 ( .A(n63), .B(n2567), .C(n2566), .D(n4505), .Z(n2042) );
  COND2X1 U1946 ( .A(n63), .B(n2568), .C(n2567), .D(n4505), .Z(n2043) );
  COND2X1 U1947 ( .A(n4316), .B(n2569), .C(n2568), .D(n4505), .Z(n2044) );
  COND2X1 U1948 ( .A(n63), .B(n2570), .C(n2569), .D(n4505), .Z(n2045) );
  COND2X1 U1949 ( .A(n63), .B(n2571), .C(n2570), .D(n4505), .Z(n2046) );
  COND2X1 U1951 ( .A(n4316), .B(n2573), .C(n2572), .D(n4505), .Z(n2048) );
  COND2X1 U1953 ( .A(n63), .B(n2575), .C(n2574), .D(n4505), .Z(n2050) );
  COND2X1 U1954 ( .A(n63), .B(n2576), .C(n2575), .D(n4505), .Z(n2051) );
  COND2X1 U1956 ( .A(n4316), .B(n2578), .C(n2577), .D(n4505), .Z(n2053) );
  COND2X1 U1958 ( .A(n63), .B(n2580), .C(n2579), .D(n4505), .Z(n2055) );
  CAOR1X1 U1994 ( .A(n4507), .B(n54), .C(n2582), .Z(n2057) );
  COND2X1 U1996 ( .A(n54), .B(n2584), .C(n4507), .D(n2583), .Z(n2059) );
  COND2X1 U1997 ( .A(n54), .B(n2585), .C(n4506), .D(n2584), .Z(n2060) );
  COND2X1 U1998 ( .A(n4184), .B(n2586), .C(n4506), .D(n2585), .Z(n2061) );
  COND2X1 U2000 ( .A(n54), .B(n2588), .C(n4506), .D(n2587), .Z(n2063) );
  COND2X1 U2002 ( .A(n4184), .B(n2590), .C(n4507), .D(n2589), .Z(n2065) );
  COND2X1 U2004 ( .A(n54), .B(n2592), .C(n4507), .D(n2591), .Z(n2067) );
  COND2X1 U2005 ( .A(n54), .B(n2593), .C(n4506), .D(n2592), .Z(n2068) );
  COND2X1 U2006 ( .A(n54), .B(n2594), .C(n4506), .D(n2593), .Z(n2069) );
  COND2X1 U2008 ( .A(n54), .B(n2596), .C(n4507), .D(n2595), .Z(n2071) );
  COND2X1 U2009 ( .A(n54), .B(n2597), .C(n4506), .D(n2596), .Z(n2072) );
  COND2X1 U2011 ( .A(n54), .B(n2599), .C(n4507), .D(n2598), .Z(n2074) );
  COND2X1 U2012 ( .A(n54), .B(n2600), .C(n4507), .D(n2599), .Z(n2075) );
  COND2X1 U2014 ( .A(n54), .B(n2602), .C(n4506), .D(n2601), .Z(n2077) );
  COND2X1 U2015 ( .A(n4184), .B(n2603), .C(n4507), .D(n2602), .Z(n2078) );
  COND2X1 U2016 ( .A(n54), .B(n2604), .C(n4507), .D(n2603), .Z(n2079) );
  COND2X1 U2017 ( .A(n4184), .B(n2605), .C(n4506), .D(n2604), .Z(n2080) );
  COND2X1 U2018 ( .A(n4184), .B(n2606), .C(n4507), .D(n2605), .Z(n2081) );
  COND2X1 U2020 ( .A(n54), .B(n2608), .C(n4507), .D(n2607), .Z(n2083) );
  COND2X1 U2021 ( .A(n54), .B(n2609), .C(n4507), .D(n2608), .Z(n2084) );
  COND2X1 U2022 ( .A(n54), .B(n2610), .C(n4506), .D(n2609), .Z(n2085) );
  COND2X1 U2025 ( .A(n54), .B(n2613), .C(n4506), .D(n2612), .Z(n2088) );
  COND2X1 U2062 ( .A(n45), .B(n2616), .C(net16420), .D(n2615), .Z(n2091) );
  COND2X1 U2065 ( .A(n45), .B(n2619), .C(net16420), .D(n2618), .Z(n2094) );
  COND2X1 U2070 ( .A(n4064), .B(n2624), .C(net16420), .D(n2623), .Z(n2099) );
  COND2X1 U2071 ( .A(n4064), .B(n2625), .C(net18914), .D(n2624), .Z(n2100) );
  COND2X1 U2072 ( .A(n4064), .B(n2626), .C(net18914), .D(n2625), .Z(n2101) );
  COND2X1 U2073 ( .A(n4064), .B(n2627), .C(net16420), .D(n2626), .Z(n2102) );
  COND2X1 U2074 ( .A(n4064), .B(n2628), .C(net16420), .D(n2627), .Z(n2103) );
  COND2X1 U2075 ( .A(n4063), .B(n2629), .C(net16420), .D(n2628), .Z(n2104) );
  COND2X1 U2076 ( .A(n4063), .B(n2630), .C(net18914), .D(n2629), .Z(n2105) );
  COND2X1 U2077 ( .A(n4064), .B(n2631), .C(net18914), .D(n2630), .Z(n2106) );
  COND2X1 U2078 ( .A(n4064), .B(n2632), .C(net16420), .D(n2631), .Z(n2107) );
  COND2X1 U2079 ( .A(n4063), .B(n2633), .C(net16420), .D(n2632), .Z(n2108) );
  COND2X1 U2080 ( .A(n45), .B(n2634), .C(net16420), .D(n2633), .Z(n2109) );
  COND2X1 U2081 ( .A(n4063), .B(n2635), .C(net16420), .D(n2634), .Z(n2110) );
  COND2X1 U2082 ( .A(n4064), .B(n2636), .C(net18914), .D(n2635), .Z(n2111) );
  COND2X1 U2083 ( .A(n4063), .B(n2637), .C(net18914), .D(n2636), .Z(n2112) );
  COND2X1 U2084 ( .A(n4063), .B(n2638), .C(net16420), .D(n2637), .Z(n2113) );
  COND2X1 U2085 ( .A(n45), .B(n2639), .C(net16420), .D(n2638), .Z(n2114) );
  COND2X1 U2087 ( .A(n4064), .B(n2641), .C(net18914), .D(n2640), .Z(n2116) );
  COND2X1 U2088 ( .A(n4064), .B(n2642), .C(net18914), .D(n2641), .Z(n2117) );
  COND2X1 U2089 ( .A(n4064), .B(n2643), .C(net16420), .D(n2642), .Z(n2118) );
  COND2X1 U2091 ( .A(n4064), .B(n2645), .C(net18914), .D(n2644), .Z(n2120) );
  COND2X1 U2092 ( .A(n4064), .B(n2646), .C(net16420), .D(n2645), .Z(n2121) );
  COND2X1 U2129 ( .A(net18896), .B(n2649), .C(net16490), .D(n2648), .Z(n2124)
         );
  COND2X1 U2132 ( .A(net18896), .B(n2652), .C(n3644), .D(n2651), .Z(n2127) );
  COND2X1 U2133 ( .A(net18896), .B(n2653), .C(n3644), .D(n4059), .Z(n2128) );
  COND2X1 U2134 ( .A(net16309), .B(n2654), .C(n3644), .D(n2653), .Z(n2129) );
  COND2X1 U2135 ( .A(net18896), .B(n2655), .C(n3644), .D(n2654), .Z(n2130) );
  COND2X1 U2136 ( .A(net18896), .B(n2656), .C(n2655), .D(n3644), .Z(n2131) );
  COND2X1 U2137 ( .A(net18896), .B(n2657), .C(n3644), .D(n2656), .Z(n2132) );
  COND2X1 U2138 ( .A(net18896), .B(n2658), .C(n3644), .D(n2657), .Z(n2133) );
  COND2X1 U2140 ( .A(net18610), .B(n2660), .C(n3644), .D(n2659), .Z(n2135) );
  COND2X1 U2141 ( .A(net16309), .B(n2661), .C(n3644), .D(n2660), .Z(n2136) );
  COND2X1 U2142 ( .A(net16309), .B(n2662), .C(n3644), .D(n2661), .Z(n2137) );
  COND2X1 U2145 ( .A(net18897), .B(n2665), .C(n3644), .D(n2664), .Z(n2140) );
  COND2X1 U2151 ( .A(net18896), .B(n2671), .C(net16490), .D(n2670), .Z(n2146)
         );
  COND2X1 U2201 ( .A(net18772), .B(n2687), .C(net17297), .D(n2686), .Z(n2161)
         );
  COND2X1 U2202 ( .A(net18772), .B(n2688), .C(net17297), .D(n2687), .Z(n2162)
         );
  COND2X1 U2203 ( .A(net18772), .B(n2689), .C(net16451), .D(n2688), .Z(n2163)
         );
  COND2X1 U2204 ( .A(net18772), .B(n2690), .C(net17297), .D(n2689), .Z(n2164)
         );
  COND2X1 U2206 ( .A(net18772), .B(n2692), .C(net16451), .D(n2691), .Z(n2166)
         );
  COND2X1 U2207 ( .A(net18772), .B(n2693), .C(net16451), .D(n2692), .Z(n2167)
         );
  COND2X1 U2208 ( .A(net18772), .B(n2694), .C(net16451), .D(n2693), .Z(n2168)
         );
  COND2X1 U2210 ( .A(n27), .B(n2696), .C(net17297), .D(n2695), .Z(n2170) );
  COND2X1 U2213 ( .A(net18772), .B(n2699), .C(net17297), .D(n2698), .Z(n2173)
         );
  COND2X1 U2215 ( .A(n27), .B(n2701), .C(net16451), .D(n2700), .Z(n2175) );
  COND2X1 U2216 ( .A(net18772), .B(n2702), .C(net16451), .D(n2701), .Z(n2176)
         );
  COND2X1 U2217 ( .A(net18772), .B(n2703), .C(net16451), .D(n2702), .Z(n2177)
         );
  COND2X1 U2218 ( .A(net18772), .B(n2704), .C(net16451), .D(n2703), .Z(n2178)
         );
  COND2X1 U2219 ( .A(net18772), .B(n2705), .C(net16451), .D(n2704), .Z(n2179)
         );
  COND2X1 U2220 ( .A(net18772), .B(n2706), .C(net16451), .D(n2705), .Z(n2180)
         );
  COND2X1 U2221 ( .A(net18772), .B(n2707), .C(net16451), .D(n2706), .Z(n2181)
         );
  COND2X1 U2226 ( .A(net18772), .B(n2712), .C(net16451), .D(n2711), .Z(n2186)
         );
  CAOR1X1 U2262 ( .A(n4510), .B(n4461), .C(n2714), .Z(n2188) );
  COND2X1 U2264 ( .A(n4461), .B(n2716), .C(n2715), .D(n4510), .Z(n2189) );
  COND2X1 U2265 ( .A(n4461), .B(n2717), .C(n2716), .D(n4510), .Z(n2190) );
  COND2X1 U2268 ( .A(n4461), .B(n2720), .C(n2719), .D(n4510), .Z(n2193) );
  COND2X1 U2269 ( .A(n4461), .B(n2721), .C(n2720), .D(n4510), .Z(n2194) );
  COND2X1 U2272 ( .A(n4461), .B(n2724), .C(n2723), .D(n4510), .Z(n2197) );
  COND2X1 U2273 ( .A(n4461), .B(n2725), .C(n2724), .D(n4510), .Z(n2198) );
  COND2X1 U2274 ( .A(n4461), .B(n2726), .C(n2725), .D(n4510), .Z(n2199) );
  COND2X1 U2275 ( .A(n4461), .B(n2727), .C(n2726), .D(n4510), .Z(n2200) );
  COND2X1 U2276 ( .A(n4460), .B(n2728), .C(n2727), .D(n4510), .Z(n2201) );
  COND2X1 U2277 ( .A(n4461), .B(n2729), .C(n2728), .D(n4510), .Z(n2202) );
  COND2X1 U2278 ( .A(n4461), .B(n2730), .C(n2729), .D(n4510), .Z(n2203) );
  COND2X1 U2279 ( .A(n4461), .B(n2731), .C(n2730), .D(n4510), .Z(n2204) );
  COND2X1 U2282 ( .A(n4461), .B(n2734), .C(n2733), .D(n4510), .Z(n2207) );
  COND2X1 U2283 ( .A(n4461), .B(n2735), .C(n2734), .D(n4510), .Z(n2208) );
  COND2X1 U2284 ( .A(n4461), .B(n2736), .C(n2735), .D(n4510), .Z(n2209) );
  COND2X1 U2290 ( .A(n4461), .B(n2742), .C(n4510), .D(n2741), .Z(n2215) );
  COND2X1 U2292 ( .A(n4461), .B(n2744), .C(n2743), .D(n4510), .Z(n2217) );
  CAOR1X1 U2329 ( .A(n6), .B(n3211), .C(n2747), .Z(n2220) );
  COND2X1 U2330 ( .A(n9), .B(n2748), .C(n6), .D(n2747), .Z(n2221) );
  COND2X1 U2331 ( .A(n3210), .B(n2749), .C(n6), .D(n2748), .Z(n2222) );
  COND2X1 U2332 ( .A(n9), .B(n2750), .C(n6), .D(n2749), .Z(n2223) );
  COND2X1 U2333 ( .A(n3211), .B(n2751), .C(n6), .D(n2750), .Z(n2224) );
  COND2X1 U2334 ( .A(n9), .B(n2752), .C(n6), .D(n2751), .Z(n2225) );
  COND2X1 U2335 ( .A(n3210), .B(n4270), .C(n6), .D(n2752), .Z(n2226) );
  COND2X1 U2336 ( .A(n9), .B(n2754), .C(n6), .D(n2753), .Z(n2227) );
  COND2X1 U2338 ( .A(n3210), .B(n2756), .C(n6), .D(n2755), .Z(n2229) );
  COND2X1 U2339 ( .A(n9), .B(n2757), .C(n6), .D(n2756), .Z(n2230) );
  COND2X1 U2341 ( .A(n3210), .B(n2759), .C(n6), .D(n2758), .Z(n2232) );
  COND2X1 U2343 ( .A(n3210), .B(n2761), .C(n6), .D(n2760), .Z(n2234) );
  COND2X1 U2344 ( .A(n9), .B(n2762), .C(n6), .D(n2761), .Z(n2235) );
  COND2X1 U2345 ( .A(n3211), .B(n2763), .C(n6), .D(n2762), .Z(n2236) );
  COND2X1 U2346 ( .A(n3211), .B(n2764), .C(n6), .D(n2763), .Z(n2237) );
  COND2X1 U2347 ( .A(n3210), .B(n2765), .C(n6), .D(n2764), .Z(n2238) );
  COND2X1 U2348 ( .A(n3211), .B(n2766), .C(n6), .D(n2765), .Z(n2239) );
  COND2X1 U2350 ( .A(n3211), .B(n2768), .C(n6), .D(n2767), .Z(n2241) );
  COND2X1 U2351 ( .A(n3211), .B(n2769), .C(n6), .D(n2768), .Z(n2242) );
  COND2X1 U2352 ( .A(n3210), .B(n2770), .C(n6), .D(n2769), .Z(n2243) );
  COND2X1 U2353 ( .A(n3211), .B(n2771), .C(n6), .D(n2770), .Z(n2244) );
  COND2X1 U2354 ( .A(n3210), .B(n2772), .C(n6), .D(n2771), .Z(n2245) );
  COND2X1 U2355 ( .A(n3210), .B(n2773), .C(n6), .D(n2772), .Z(n2246) );
  COND2X1 U2356 ( .A(n3211), .B(n2774), .C(n6), .D(n2773), .Z(n2247) );
  COND2X1 U2357 ( .A(n3211), .B(n2775), .C(n6), .D(n2774), .Z(n2248) );
  COND2X1 U2358 ( .A(n3211), .B(n2776), .C(n6), .D(n2775), .Z(n2249) );
  COND2X1 U2359 ( .A(n3211), .B(n2777), .C(n6), .D(n2776), .Z(n2250) );
  COND2X1 U2360 ( .A(n3210), .B(n2778), .C(n6), .D(n2777), .Z(n2251) );
  CND2IX1 U2394 ( .B(n3244), .A(n4571), .Z(n2779) );
  CND2X2 U441 ( .A(n3937), .B(n751), .Z(n444) );
  CNR2X2 U473 ( .A(n1036), .B(n1015), .Z(n468) );
  COND2X1 U2196 ( .A(n2682), .B(net18772), .C(net17297), .D(n2681), .Z(n1184)
         );
  CNR2X2 U521 ( .A(n1107), .B(n1132), .Z(n504) );
  COND2X1 U2066 ( .A(n45), .B(n2620), .C(net16420), .D(n2619), .Z(n2095) );
  COND2X1 U1351 ( .A(n144), .B(n2279), .C(n2278), .D(n3277), .Z(n1763) );
  COND2X1 U1481 ( .A(net17738), .B(n2341), .C(n123), .D(n2340), .Z(n1825) );
  COND2X1 U1416 ( .A(net18310), .B(n2310), .C(net16438), .D(n2309), .Z(n1794)
         );
  CFA1X1 U1049 ( .A(n1763), .B(n1825), .CI(n1794), .CO(n1178), .S(n1179) );
  COND2X1 U1871 ( .A(net16301), .B(n2527), .C(n3122), .D(n2526), .Z(n2004) );
  COND2X1 U1676 ( .A(net18627), .B(n2434), .C(n4508), .D(n2433), .Z(n1911) );
  COND2X1 U1546 ( .A(net18628), .B(n2372), .C(net16433), .D(n2371), .Z(n1856)
         );
  CFA1X1 U1048 ( .A(n2004), .B(n1911), .CI(n1856), .CO(n1176), .S(n1177) );
  COND2X1 U2131 ( .A(n3920), .B(net18897), .C(net16490), .D(n2650), .Z(n2126)
         );
  CFA1X1 U1033 ( .A(n1182), .B(n1176), .CI(n1178), .CO(n1146), .S(n1147) );
  CFA1X1 U1051 ( .A(n1880), .B(n2095), .CI(n2126), .CO(n1182), .S(n1183) );
  COND2X1 U1872 ( .A(n3142), .B(n2528), .C(n3122), .D(n2527), .Z(n2005) );
  COND2X1 U1612 ( .A(n3301), .B(n2404), .C(n2403), .D(net17425), .Z(n1881) );
  CFA1X1 U1058 ( .A(n1211), .B(n1230), .CI(n1209), .CO(n1196), .S(n1197) );
  COND2X1 U1741 ( .A(n3991), .B(n2465), .C(net16512), .D(n2464), .Z(n1942) );
  CFA1X1 U1030 ( .A(n1172), .B(n1170), .CI(n1174), .CO(n1140), .S(n1141) );
  COND2X1 U1480 ( .A(net17738), .B(n2340), .C(n123), .D(n2339), .Z(n1824) );
  COND2X1 U1415 ( .A(n135), .B(n2309), .C(net16438), .D(n2308), .Z(n1793) );
  CFA1X1 U1035 ( .A(n1762), .B(n1824), .CI(n1793), .CO(n1150), .S(n1151) );
  CFA1X1 U1001 ( .A(n1087), .B(n1085), .CI(n1108), .CO(n1082), .S(n1083) );
  CND2X1 U2507 ( .A(n3427), .B(n2237), .Z(n4362) );
  CND2X1 U2508 ( .A(n2076), .B(n2107), .Z(n3702) );
  CND2X1 U2509 ( .A(n3992), .B(n3753), .Z(n3995) );
  CENX1 U2510 ( .A(n1542), .B(n1540), .Z(n3842) );
  CENX2 U2511 ( .A(net17419), .B(n4553), .Z(n2399) );
  CIVX2 U2512 ( .A(n3772), .Z(n3534) );
  COND2X2 U2513 ( .A(n4316), .B(n2566), .C(n2565), .D(n4505), .Z(n2041) );
  CEOX2 U2514 ( .A(n1576), .B(n1574), .Z(n3022) );
  CEOX2 U2515 ( .A(n3022), .B(n1572), .Z(n1553) );
  CND2XL U2516 ( .A(n1572), .B(n1574), .Z(n3023) );
  CND2XL U2517 ( .A(n1572), .B(n1576), .Z(n3024) );
  CND2XL U2518 ( .A(n1574), .B(n1576), .Z(n3025) );
  CND3X1 U2519 ( .A(n3023), .B(n3024), .C(n3025), .Z(n1552) );
  CND3X2 U2520 ( .A(n4258), .B(n4259), .C(n4260), .Z(n1574) );
  CIVX3 U2521 ( .A(n3777), .Z(net16301) );
  CNIVX4 U2522 ( .A(n4588), .Z(n3026) );
  CNIVX1 U2523 ( .A(n4588), .Z(n4086) );
  CAN2X1 U2524 ( .A(n4373), .B(n3762), .Z(n3027) );
  CNR2X1 U2525 ( .A(n671), .B(n674), .Z(n669) );
  CNR2X2 U2526 ( .A(n1641), .B(n1652), .Z(n671) );
  CIVX4 U2527 ( .A(net18913), .Z(net18914) );
  CIVXL U2528 ( .A(n4598), .Z(n3028) );
  CND2XL U2529 ( .A(n1139), .B(n1164), .Z(n3936) );
  CND2XL U2530 ( .A(n1155), .B(n1180), .Z(net19067) );
  CND2X1 U2531 ( .A(n4594), .B(a[22]), .Z(n3031) );
  CND2X2 U2532 ( .A(n3029), .B(n3030), .Z(n3032) );
  CND2X4 U2533 ( .A(n3031), .B(n3032), .Z(n3890) );
  CIVX2 U2534 ( .A(n4594), .Z(n3029) );
  CIVX2 U2535 ( .A(a[22]), .Z(n3030) );
  CIVX4 U2536 ( .A(n3890), .Z(net16426) );
  CND2X1 U2537 ( .A(n3657), .B(n1307), .Z(n3035) );
  CND2X2 U2538 ( .A(n3033), .B(n3034), .Z(n3036) );
  CND2X2 U2539 ( .A(n3035), .B(n3036), .Z(n1305) );
  CIVX1 U2540 ( .A(n3657), .Z(n3033) );
  CIVXL U2541 ( .A(n1307), .Z(n3034) );
  COND2XL U2542 ( .A(net18897), .B(n2669), .C(net16490), .D(n2668), .Z(n2144)
         );
  CND2XL U2543 ( .A(n773), .B(n628), .Z(n191) );
  CND2XL U2544 ( .A(n1485), .B(n1506), .Z(n3793) );
  CND2X1 U2545 ( .A(n1506), .B(n1487), .Z(n3795) );
  CFA1X1 U2546 ( .A(n1765), .B(n1858), .CI(n1796), .CO(n1234), .S(n1235) );
  COND2X1 U2547 ( .A(net18310), .B(n2312), .C(net16438), .D(n2311), .Z(n1796)
         );
  CNIVXL U2548 ( .A(n1181), .Z(net18689) );
  COND1XL U2549 ( .A(n544), .B(n540), .C(n541), .Z(n3037) );
  CND2XL U2550 ( .A(n1289), .B(n1287), .Z(n3040) );
  CND2X2 U2551 ( .A(n3038), .B(n3039), .Z(n3041) );
  CND2X2 U2552 ( .A(n3040), .B(n3041), .Z(n4487) );
  CIVXL U2553 ( .A(n1289), .Z(n3038) );
  CIVX1 U2554 ( .A(n1287), .Z(n3039) );
  CENX2 U2555 ( .A(n1414), .B(n1391), .Z(n4154) );
  CND3X2 U2556 ( .A(n4079), .B(n4080), .C(n4081), .Z(n1414) );
  COND2X2 U2557 ( .A(n4460), .B(n2723), .C(n2722), .D(n4510), .Z(n2196) );
  CND2X1 U2558 ( .A(n4333), .B(n4334), .Z(n2479) );
  CNIVX1 U2559 ( .A(n1117), .Z(n3143) );
  CANR1X1 U2560 ( .A(n562), .B(n549), .C(n550), .Z(n3042) );
  CND2X1 U2561 ( .A(n1323), .B(n1331), .Z(n3045) );
  CND2X2 U2562 ( .A(n3043), .B(n3044), .Z(n3046) );
  CND2X2 U2563 ( .A(n3045), .B(n3046), .Z(n4014) );
  CIVX2 U2564 ( .A(n1323), .Z(n3043) );
  CIVX2 U2565 ( .A(n1331), .Z(n3044) );
  CANR1X1 U2566 ( .A(n562), .B(n549), .C(n550), .Z(n548) );
  CIVX1 U2567 ( .A(n3874), .Z(net18897) );
  CND3X2 U2568 ( .A(n4318), .B(net17759), .C(net17758), .Z(n1084) );
  CND2IX1 U2569 ( .B(net18199), .A(n1110), .Z(n4318) );
  CIVX3 U2570 ( .A(net18824), .Z(net16438) );
  CENX1 U2571 ( .A(net16541), .B(n4560), .Z(n2689) );
  CENXL U2572 ( .A(n3047), .B(n1599), .Z(n1597) );
  CENX2 U2573 ( .A(n1601), .B(n1614), .Z(n3047) );
  COND2XL U2574 ( .A(n4063), .B(n2640), .C(net18914), .D(n2639), .Z(n2115) );
  CNR2XL U2575 ( .A(n4063), .B(n2621), .Z(n4257) );
  CENXL U2576 ( .A(n4582), .B(n2785), .Z(n2521) );
  CENXL U2577 ( .A(n4582), .B(n4554), .Z(n2530) );
  CEOX2 U2578 ( .A(n1313), .B(n1311), .Z(n3048) );
  CEOX2 U2579 ( .A(n1336), .B(n3048), .Z(n1307) );
  CND2X1 U2580 ( .A(n1336), .B(n1311), .Z(n3049) );
  CND2X1 U2581 ( .A(n1336), .B(n1313), .Z(n3050) );
  CND2XL U2582 ( .A(n1311), .B(n1313), .Z(n3051) );
  CND3X2 U2583 ( .A(n3049), .B(n3050), .C(n3051), .Z(n1306) );
  CND3X2 U2584 ( .A(n3391), .B(n3393), .C(n3392), .Z(n1336) );
  CIVX1 U2585 ( .A(n1306), .Z(n3581) );
  CND2X1 U2586 ( .A(n1328), .B(n1330), .Z(n3105) );
  CND2XL U2587 ( .A(n1330), .B(n1303), .Z(n3107) );
  CIVXL U2588 ( .A(net16426), .Z(n3899) );
  CEOX2 U2589 ( .A(net18209), .B(n4546), .Z(n2406) );
  CENX1 U2590 ( .A(n4597), .B(n4542), .Z(n2344) );
  CIVX2 U2591 ( .A(n4462), .Z(n3248) );
  CNIVX1 U2592 ( .A(n1136), .Z(n3219) );
  CND2X1 U2593 ( .A(n1302), .B(n2067), .Z(n3547) );
  CND2IX1 U2594 ( .B(n1226), .A(n3604), .Z(n3605) );
  CND2XL U2595 ( .A(n4121), .B(n4555), .Z(n3054) );
  CND2X1 U2596 ( .A(n3052), .B(n3053), .Z(n3055) );
  CND2X1 U2597 ( .A(n3054), .B(n3055), .Z(n2562) );
  CIVXL U2598 ( .A(n4121), .Z(n3052) );
  CIVXL U2599 ( .A(n4555), .Z(n3053) );
  CENX2 U2600 ( .A(n3056), .B(n1355), .Z(n1345) );
  CENX2 U2601 ( .A(n1382), .B(n3366), .Z(n3056) );
  CENX2 U2602 ( .A(n2065), .B(n1240), .Z(n3775) );
  CEOX2 U2603 ( .A(n1491), .B(n1508), .Z(n3057) );
  CEOX2 U2604 ( .A(n3057), .B(n1489), .Z(n1485) );
  CND2X1 U2605 ( .A(n1489), .B(n1508), .Z(n3058) );
  CND2X1 U2606 ( .A(n1489), .B(n1491), .Z(n3059) );
  CND2XL U2607 ( .A(n1508), .B(n1491), .Z(n3060) );
  CND3X2 U2608 ( .A(n3058), .B(n3059), .C(n3060), .Z(n1484) );
  CENX2 U2609 ( .A(n1465), .B(n1484), .Z(n4478) );
  CENX1 U2610 ( .A(n3061), .B(n1363), .Z(n1361) );
  CENX1 U2611 ( .A(n1388), .B(n1365), .Z(n3061) );
  CNIVX4 U2612 ( .A(n1190), .Z(n3488) );
  CND3XL U2613 ( .A(n4261), .B(n4262), .C(n4263), .Z(n3062) );
  CND3XL U2614 ( .A(n4261), .B(n4262), .C(n4263), .Z(n3063) );
  CND3XL U2615 ( .A(n4261), .B(n4262), .C(n4263), .Z(n1568) );
  CND2X1 U2616 ( .A(n1424), .B(n1405), .Z(n3375) );
  CND2X1 U2617 ( .A(n1424), .B(n1407), .Z(n3374) );
  CEO3X1 U2618 ( .A(n1913), .B(n2006), .C(n1243), .Z(n1233) );
  CND2XL U2619 ( .A(n1913), .B(n1243), .Z(n3064) );
  CND2XL U2620 ( .A(n1913), .B(n2006), .Z(n3065) );
  CND2X1 U2621 ( .A(n1243), .B(n2006), .Z(n3066) );
  CND3X1 U2622 ( .A(n3064), .B(n3065), .C(n3066), .Z(n1232) );
  CIVX1 U2623 ( .A(n1242), .Z(n1243) );
  CNIVX1 U2624 ( .A(n2134), .Z(n3755) );
  CND2X1 U2625 ( .A(n355), .B(n320), .Z(n318) );
  CENX1 U2626 ( .A(n4585), .B(n4562), .Z(n2489) );
  CENX1 U2627 ( .A(n3097), .B(n3067), .Z(n1247) );
  CENX1 U2628 ( .A(n1251), .B(n1253), .Z(n3067) );
  CND2X1 U2629 ( .A(n4478), .B(n1463), .Z(n3070) );
  CND2X2 U2630 ( .A(n3068), .B(n3069), .Z(n3071) );
  CND2X2 U2631 ( .A(n3070), .B(n3071), .Z(n1461) );
  CIVX2 U2632 ( .A(n4478), .Z(n3068) );
  CIVXL U2633 ( .A(n1463), .Z(n3069) );
  CND2X1 U2634 ( .A(n3633), .B(n3073), .Z(n3074) );
  CND2XL U2635 ( .A(n3072), .B(n3098), .Z(n3075) );
  CND2X1 U2636 ( .A(n3074), .B(n3075), .Z(n1465) );
  CIVX2 U2637 ( .A(n3633), .Z(n3072) );
  CIVXL U2638 ( .A(n3098), .Z(n3073) );
  CEO3X1 U2639 ( .A(n1479), .B(n1475), .C(n1477), .Z(n3098) );
  CIVXL U2640 ( .A(n1329), .Z(n3076) );
  CIVX1 U2641 ( .A(n3076), .Z(n3077) );
  CIVX2 U2642 ( .A(n3719), .Z(n3078) );
  CIVX2 U2643 ( .A(n3719), .Z(n4593) );
  CENX1 U2644 ( .A(n3079), .B(n2018), .Z(n1537) );
  CENX1 U2645 ( .A(n1956), .B(n2109), .Z(n3079) );
  CND2XL U2646 ( .A(n3645), .B(n4542), .Z(n3082) );
  CND2X1 U2647 ( .A(n3080), .B(n3081), .Z(n3083) );
  CND2X1 U2648 ( .A(n3082), .B(n3083), .Z(n2542) );
  CIVXL U2649 ( .A(n3645), .Z(n3080) );
  CIVXL U2650 ( .A(n4542), .Z(n3081) );
  CNR2IX2 U2651 ( .B(n2820), .A(net16959), .Z(net17154) );
  CND2X2 U2652 ( .A(n3834), .B(n3835), .Z(n3084) );
  CENX2 U2653 ( .A(n4601), .B(a[30]), .Z(n3085) );
  CENXL U2654 ( .A(n4601), .B(a[30]), .Z(n3086) );
  CENX2 U2655 ( .A(n4601), .B(a[30]), .Z(net18548) );
  CNIVX2 U2656 ( .A(n3669), .Z(n4501) );
  CND2X1 U2657 ( .A(n3268), .B(n896), .Z(n3089) );
  CND2X2 U2658 ( .A(n3087), .B(n3088), .Z(n3090) );
  CND2X2 U2659 ( .A(n3089), .B(n3090), .Z(n881) );
  CIVX2 U2660 ( .A(n3268), .Z(n3087) );
  CIVXL U2661 ( .A(n896), .Z(n3088) );
  CND2X1 U2662 ( .A(n885), .B(n898), .Z(n3093) );
  CND2X2 U2663 ( .A(n3091), .B(n3092), .Z(n3094) );
  CND2X2 U2664 ( .A(n3093), .B(n3094), .Z(n3268) );
  CIVX1 U2665 ( .A(n885), .Z(n3091) );
  CIVXL U2666 ( .A(n898), .Z(n3092) );
  CND2X2 U2667 ( .A(n4199), .B(n4200), .Z(n3095) );
  CND2X2 U2668 ( .A(n4199), .B(n4200), .Z(n4310) );
  CIVX1 U2669 ( .A(n628), .Z(n626) );
  CENX1 U2670 ( .A(n1337), .B(n1362), .Z(n3779) );
  CND2XL U2671 ( .A(n1362), .B(n1337), .Z(n4172) );
  CIVX1 U2672 ( .A(n3874), .Z(net16309) );
  CIVX2 U2673 ( .A(n3144), .Z(n3669) );
  CEOX2 U2674 ( .A(n3621), .B(n4554), .Z(n2563) );
  CIVX2 U2675 ( .A(n4121), .Z(n3621) );
  CIVX1 U2676 ( .A(n1278), .Z(n3096) );
  CIVX2 U2677 ( .A(n3096), .Z(n3097) );
  CENX1 U2678 ( .A(n1219), .B(n1246), .Z(n3823) );
  CND2X1 U2679 ( .A(n2813), .B(net16437), .Z(n135) );
  CIVX8 U2680 ( .A(n3579), .Z(n4505) );
  CIVX2 U2681 ( .A(n4397), .Z(n3099) );
  CIVX2 U2682 ( .A(a[18]), .Z(n4397) );
  CIVXL U2683 ( .A(n1861), .Z(n3100) );
  CIVX1 U2684 ( .A(n3100), .Z(n3101) );
  CND2X2 U2685 ( .A(n4411), .B(n4412), .Z(n2413) );
  CND2X1 U2686 ( .A(n2809), .B(net17419), .Z(n4411) );
  CND2X1 U2687 ( .A(n1472), .B(n1449), .Z(n4192) );
  CNR2X2 U2688 ( .A(n1361), .B(n1386), .Z(n572) );
  CIVXL U2689 ( .A(net18419), .Z(n3102) );
  CENX2 U2690 ( .A(n3103), .B(n960), .Z(n941) );
  CENX2 U2691 ( .A(n962), .B(n945), .Z(n3103) );
  CEOX2 U2692 ( .A(n1303), .B(n1330), .Z(n3104) );
  CEOX2 U2693 ( .A(n3104), .B(n1328), .Z(n1291) );
  CND2X2 U2694 ( .A(n1328), .B(n1303), .Z(n3106) );
  CND3X2 U2695 ( .A(n3105), .B(n3106), .C(n3107), .Z(n1290) );
  CND2XL U2696 ( .A(n1269), .B(n1290), .Z(n4125) );
  CND2X1 U2697 ( .A(n4233), .B(n1257), .Z(n3110) );
  CND2X2 U2698 ( .A(n3108), .B(n3109), .Z(n3111) );
  CND2X2 U2699 ( .A(n3110), .B(n3111), .Z(n1251) );
  CIVX2 U2700 ( .A(n4233), .Z(n3108) );
  CIVXL U2701 ( .A(n1257), .Z(n3109) );
  CENX1 U2702 ( .A(n1286), .B(n1284), .Z(n4233) );
  CIVX3 U2703 ( .A(n4094), .Z(n4575) );
  CND2X2 U2704 ( .A(n1505), .B(n1524), .Z(n623) );
  CENX1 U2705 ( .A(n3112), .B(n1039), .Z(n4041) );
  CENX1 U2706 ( .A(n1060), .B(n1041), .Z(n3112) );
  CIVXL U2707 ( .A(n3777), .Z(n3113) );
  CIVX8 U2708 ( .A(a[8]), .Z(net18420) );
  CNIVXL U2709 ( .A(n3454), .Z(n3114) );
  CND2X1 U2710 ( .A(n1548), .B(n1533), .Z(n3805) );
  CIVXL U2711 ( .A(n1548), .Z(n3611) );
  CND2X2 U2712 ( .A(n4441), .B(n4442), .Z(n3115) );
  CIVX1 U2713 ( .A(net17930), .Z(n3116) );
  COND2X1 U2714 ( .A(n90), .B(n2463), .C(net16511), .D(n2462), .Z(n1940) );
  CENX2 U2715 ( .A(net17411), .B(n4556), .Z(n2396) );
  CIVX3 U2716 ( .A(net18824), .Z(net16439) );
  CIVX3 U2717 ( .A(net17154), .Z(n3117) );
  CIVX2 U2718 ( .A(net17154), .Z(net17278) );
  CND2X1 U2719 ( .A(n1464), .B(n1443), .Z(n4197) );
  CIVX1 U2720 ( .A(a[20]), .Z(n4440) );
  CIVXL U2721 ( .A(a[20]), .Z(n3876) );
  CENX2 U2722 ( .A(n3118), .B(n1196), .Z(n1165) );
  CENX2 U2723 ( .A(n1198), .B(n1171), .Z(n3118) );
  CND2X2 U2724 ( .A(n4441), .B(n4442), .Z(n96) );
  CIVXL U2725 ( .A(n1304), .Z(n3119) );
  CIVXL U2726 ( .A(n3119), .Z(n3120) );
  CND3XL U2727 ( .A(n4030), .B(n4031), .C(n4032), .Z(n3894) );
  CIVX3 U2728 ( .A(n3380), .Z(n3121) );
  CIVX3 U2729 ( .A(n3380), .Z(n3122) );
  CIVX2 U2730 ( .A(n3380), .Z(net16465) );
  CIVX3 U2731 ( .A(net18218), .Z(n3328) );
  CND2X1 U2732 ( .A(n1442), .B(n1419), .Z(n4079) );
  COND2X1 U2733 ( .A(n3991), .B(n2458), .C(net16512), .D(n2457), .Z(n1935) );
  CND2X4 U2734 ( .A(n3222), .B(n3223), .Z(n1171) );
  CND2XL U2735 ( .A(n383), .B(n745), .Z(n372) );
  CIVXL U2736 ( .A(n3977), .Z(n3519) );
  CND2XL U2737 ( .A(n1157), .B(n1180), .Z(n3919) );
  CND2XL U2738 ( .A(n1155), .B(n1157), .Z(net19066) );
  CND2X1 U2739 ( .A(n1490), .B(n3124), .Z(n3125) );
  CND2X2 U2740 ( .A(n3123), .B(n1471), .Z(n3126) );
  CND2X2 U2741 ( .A(n3125), .B(n3126), .Z(n3633) );
  CIVX2 U2742 ( .A(n1490), .Z(n3123) );
  CIVX1 U2743 ( .A(n1471), .Z(n3124) );
  CFA1X1 U2744 ( .A(n1520), .B(n1499), .CI(n1497), .CO(n1490), .S(n1491) );
  CND2XL U2745 ( .A(n3828), .B(n2785), .Z(n3129) );
  CND2X1 U2746 ( .A(n3127), .B(n3128), .Z(n3130) );
  CND2X1 U2747 ( .A(n3129), .B(n3130), .Z(n2389) );
  CIVXL U2748 ( .A(n3828), .Z(n3127) );
  CIVXL U2749 ( .A(n2785), .Z(n3128) );
  CND2XL U2750 ( .A(n1327), .B(n1325), .Z(n4535) );
  CEOX1 U2751 ( .A(n1885), .B(n1830), .Z(n3513) );
  CENXL U2752 ( .A(n1389), .B(n4154), .Z(n3131) );
  CENX1 U2753 ( .A(n1389), .B(n4154), .Z(n1387) );
  CNR2X2 U2754 ( .A(n1545), .B(n1562), .Z(n633) );
  CND2X2 U2755 ( .A(n1545), .B(n1562), .Z(n634) );
  CEOX2 U2756 ( .A(n1549), .B(n1564), .Z(n4387) );
  CENX2 U2757 ( .A(n1529), .B(n1546), .Z(n3772) );
  CND2X1 U2758 ( .A(n1467), .B(n1488), .Z(n3698) );
  CIVX4 U2759 ( .A(n3248), .Z(n4507) );
  CIVX1 U2760 ( .A(n605), .Z(n770) );
  CIVX1 U2761 ( .A(n1417), .Z(n3962) );
  CENX2 U2762 ( .A(n3132), .B(n3164), .Z(n1231) );
  CENX2 U2763 ( .A(n1272), .B(n1268), .Z(n3132) );
  CIVXL U2764 ( .A(n3777), .Z(n3133) );
  CENXL U2765 ( .A(n4579), .B(n2785), .Z(n2587) );
  CENXL U2766 ( .A(n4579), .B(n4563), .Z(n2586) );
  CENXL U2767 ( .A(n4579), .B(n4561), .Z(n2589) );
  CND2XL U2768 ( .A(n1135), .B(n1137), .Z(n4385) );
  CFA1XL U2769 ( .A(n1751), .B(n1930), .CI(n1961), .CO(n918), .S(n919) );
  CENX2 U2770 ( .A(n1124), .B(n1122), .Z(n3881) );
  CND3X2 U2771 ( .A(n3151), .B(n3152), .C(n3153), .Z(n1122) );
  CND2XL U2772 ( .A(net15912), .B(n4545), .Z(n3136) );
  CND2X1 U2773 ( .A(n3134), .B(n3135), .Z(n3137) );
  CND2X1 U2774 ( .A(n3136), .B(n3137), .Z(n2407) );
  CIVXL U2775 ( .A(net15912), .Z(n3134) );
  CIVXL U2776 ( .A(n4545), .Z(n3135) );
  CIVX3 U2777 ( .A(net17410), .Z(net17411) );
  CND2XL U2778 ( .A(n4572), .B(n2785), .Z(n3140) );
  CND2X1 U2779 ( .A(n3138), .B(n3139), .Z(n3141) );
  CND2X1 U2780 ( .A(n3140), .B(n3141), .Z(n2719) );
  CIVXL U2781 ( .A(n4572), .Z(n3138) );
  CIVXL U2782 ( .A(n2785), .Z(n3139) );
  CIVXL U2783 ( .A(n3777), .Z(n3142) );
  CIVXL U2784 ( .A(n84), .Z(n3144) );
  CNIVXL U2785 ( .A(n2107), .Z(n3145) );
  CND2IX2 U2786 ( .B(n471), .A(n3194), .Z(n3196) );
  CNR2X2 U2787 ( .A(n1037), .B(n1058), .Z(n471) );
  CENX1 U2788 ( .A(n4512), .B(n4556), .Z(n2726) );
  CND3X1 U2789 ( .A(n3916), .B(n3917), .C(n3918), .Z(n1138) );
  CFA1X2 U2790 ( .A(n2158), .B(n1944), .CI(n2128), .CO(n1240), .S(n1241) );
  CEOX2 U2791 ( .A(n3471), .B(n991), .Z(n983) );
  CEOX2 U2792 ( .A(n871), .B(n880), .Z(n3146) );
  CEOX2 U2793 ( .A(n3146), .B(n869), .Z(n867) );
  CND2XL U2794 ( .A(n869), .B(n880), .Z(n3147) );
  CND2X1 U2795 ( .A(n869), .B(n871), .Z(n3148) );
  CND2XL U2796 ( .A(n880), .B(n871), .Z(n3149) );
  CND3XL U2797 ( .A(n3147), .B(n3148), .C(n3149), .Z(n866) );
  CND3X2 U2798 ( .A(n3298), .B(n3299), .C(n3300), .Z(n880) );
  COR2X2 U2799 ( .A(n855), .B(n866), .Z(n4479) );
  CND2X1 U2800 ( .A(n855), .B(n866), .Z(n351) );
  CND2IX2 U2801 ( .B(n1063), .A(n3231), .Z(n3233) );
  CEO3X2 U2802 ( .A(n2074), .B(n2105), .C(n2136), .Z(n1451) );
  CND3X2 U2803 ( .A(n3862), .B(n3863), .C(n3864), .Z(n1492) );
  CND2X1 U2804 ( .A(n1522), .B(n1516), .Z(n3862) );
  CEOX2 U2805 ( .A(n3761), .B(n4553), .Z(n2498) );
  CENX1 U2806 ( .A(n1220), .B(n1193), .Z(n3585) );
  CENXL U2807 ( .A(n4579), .B(net16102), .Z(n2584) );
  COND2XL U2808 ( .A(n2589), .B(n54), .C(n4506), .D(n2588), .Z(n2064) );
  CND2IX1 U2809 ( .B(n3244), .A(n3078), .Z(n2449) );
  CIVXL U2810 ( .A(n643), .Z(n776) );
  CND2X1 U2811 ( .A(n1581), .B(n1596), .Z(n644) );
  CND2XL U2812 ( .A(n1247), .B(n1276), .Z(n4097) );
  CEOX1 U2813 ( .A(n2002), .B(n1971), .Z(n3150) );
  CEOX1 U2814 ( .A(n3150), .B(n1909), .Z(n1123) );
  CND2XL U2815 ( .A(n1909), .B(n1971), .Z(n3151) );
  CND2X1 U2816 ( .A(n2002), .B(n1909), .Z(n3152) );
  CND2X1 U2817 ( .A(n1971), .B(n2002), .Z(n3153) );
  CND2X1 U2818 ( .A(n2062), .B(n1823), .Z(n3399) );
  CND2X1 U2819 ( .A(n1246), .B(n1219), .Z(n4380) );
  CND2X2 U2820 ( .A(n3521), .B(n3522), .Z(n1219) );
  CND2XL U2821 ( .A(n4319), .B(n4320), .Z(n3154) );
  CND2X1 U2822 ( .A(n1367), .B(n1392), .Z(n3544) );
  CND2X2 U2823 ( .A(n1395), .B(n3156), .Z(n3157) );
  CND2X1 U2824 ( .A(n1393), .B(n3155), .Z(n3158) );
  CND2X2 U2825 ( .A(n3157), .B(n3158), .Z(n3626) );
  CIVXL U2826 ( .A(n1395), .Z(n3155) );
  CIVX2 U2827 ( .A(n1393), .Z(n3156) );
  CEOX2 U2828 ( .A(n3373), .B(n1424), .Z(n1395) );
  CND2X1 U2829 ( .A(n3462), .B(n3776), .Z(n3161) );
  CND2X2 U2830 ( .A(n3159), .B(n3160), .Z(n3162) );
  CND2X2 U2831 ( .A(n3161), .B(n3162), .Z(n1311) );
  CIVXL U2832 ( .A(n3462), .Z(n3159) );
  CIVX2 U2833 ( .A(n3776), .Z(n3160) );
  CIVX1 U2834 ( .A(n1270), .Z(n3163) );
  CIVX2 U2835 ( .A(n3163), .Z(n3164) );
  CIVXL U2836 ( .A(n3190), .Z(n3165) );
  CND3X1 U2837 ( .A(n3692), .B(n3693), .C(n3694), .Z(n1230) );
  CIVX2 U2838 ( .A(n1258), .Z(n3186) );
  CANR1XL U2839 ( .A(n646), .B(n3490), .C(n639), .Z(n4226) );
  CEO3X1 U2840 ( .A(n1144), .B(n1142), .C(n1119), .Z(n1113) );
  CND2XL U2841 ( .A(n1144), .B(n1119), .Z(n3166) );
  CND2X1 U2842 ( .A(n3170), .B(n1142), .Z(n3167) );
  CND2X1 U2843 ( .A(n1119), .B(n1142), .Z(n3168) );
  CND3X2 U2844 ( .A(n3166), .B(n3167), .C(n3168), .Z(n1112) );
  CIVXL U2845 ( .A(n1144), .Z(n3169) );
  CIVXL U2846 ( .A(n3169), .Z(n3170) );
  CND3X2 U2847 ( .A(n3738), .B(n3739), .C(n3740), .Z(n1142) );
  CENX1 U2848 ( .A(n1152), .B(net18574), .Z(n1119) );
  CND2X1 U2849 ( .A(n3332), .B(n1112), .Z(net17758) );
  CND3X1 U2850 ( .A(net19066), .B(net19067), .C(n3919), .Z(n1144) );
  CIVX3 U2851 ( .A(n3753), .Z(n3993) );
  COND2XL U2852 ( .A(n4120), .B(n2487), .C(net16413), .D(n2486), .Z(n1964) );
  CND2XL U2853 ( .A(n1461), .B(n1482), .Z(n3171) );
  CND2XL U2854 ( .A(n1461), .B(n1482), .Z(n3172) );
  CND2X1 U2855 ( .A(n1482), .B(n1461), .Z(n606) );
  COND2X1 U2856 ( .A(n54), .B(n2591), .C(n4507), .D(n2590), .Z(n2066) );
  CNR2X1 U2857 ( .A(n636), .B(n633), .Z(n631) );
  CIVX1 U2858 ( .A(n641), .Z(n639) );
  CND2X1 U2859 ( .A(n1218), .B(n1193), .Z(n4043) );
  CND2X1 U2860 ( .A(n1218), .B(n1220), .Z(n4044) );
  CND2X2 U2861 ( .A(n1252), .B(n1225), .Z(n4032) );
  CND2IX1 U2862 ( .B(n1438), .A(n1417), .Z(n3963) );
  CND3XL U2863 ( .A(n4195), .B(n4197), .C(n4196), .Z(n3173) );
  CND3XL U2864 ( .A(n4195), .B(n4197), .C(n4196), .Z(n3174) );
  CND3XL U2865 ( .A(n4195), .B(n4197), .C(n4196), .Z(n1438) );
  CIVX1 U2866 ( .A(n3289), .Z(n3290) );
  CND2IX2 U2867 ( .B(n4464), .A(n3175), .Z(n1242) );
  COR2X1 U2868 ( .A(n2714), .B(n15), .Z(n3175) );
  CND2X1 U2869 ( .A(n1136), .B(n1113), .Z(n3417) );
  CND3X1 U2870 ( .A(n4027), .B(n4028), .C(n4029), .Z(n1318) );
  CEO3X1 U2871 ( .A(n1127), .B(n1146), .C(n1121), .Z(n1115) );
  CNIVXL U2872 ( .A(n1459), .Z(n3176) );
  CND3X2 U2873 ( .A(net17989), .B(net17987), .C(n3915), .Z(n1136) );
  CND3X1 U2874 ( .A(n3998), .B(n4000), .C(n3999), .Z(n3517) );
  CIVX4 U2875 ( .A(n3085), .Z(net16496) );
  CIVX1 U2876 ( .A(n3580), .Z(n3249) );
  CIVX2 U2877 ( .A(net15910), .Z(net17410) );
  CNR2XL U2878 ( .A(n594), .B(n4155), .Z(n3177) );
  CEO3X2 U2879 ( .A(n1519), .B(n1517), .C(n1534), .Z(n1511) );
  CND2XL U2880 ( .A(n1519), .B(n1534), .Z(n3178) );
  CND2XL U2881 ( .A(n1519), .B(n1517), .Z(n3179) );
  CND2XL U2882 ( .A(n1534), .B(n1517), .Z(n3180) );
  CND3X2 U2883 ( .A(n3178), .B(n3179), .C(n3180), .Z(n1510) );
  CNR2IX1 U2884 ( .B(n3751), .A(net16433), .Z(n1867) );
  CND2X1 U2885 ( .A(n878), .B(n867), .Z(n370) );
  CND2X1 U2886 ( .A(n744), .B(n370), .Z(n162) );
  CFA1X1 U2887 ( .A(n1975), .B(n1827), .CI(n2035), .CO(n1236), .S(n1237) );
  CND2XL U2888 ( .A(n1366), .B(n1368), .Z(n3393) );
  CND2XL U2889 ( .A(n1343), .B(n1366), .Z(n3391) );
  CEOX1 U2890 ( .A(n1343), .B(n1366), .Z(n3390) );
  CNIVXL U2891 ( .A(n4113), .Z(n3181) );
  CEOX1 U2892 ( .A(n1041), .B(n1060), .Z(n3182) );
  CEOX1 U2893 ( .A(n3182), .B(n1039), .Z(n1037) );
  CND2XL U2894 ( .A(n1039), .B(n1060), .Z(n3183) );
  CND2XL U2895 ( .A(n1039), .B(n1041), .Z(n3184) );
  CND2XL U2896 ( .A(n1060), .B(n1041), .Z(n3185) );
  CND3X1 U2897 ( .A(n3183), .B(n3184), .C(n3185), .Z(n1036) );
  CNIVX1 U2898 ( .A(n2040), .Z(n4530) );
  CND2X1 U2899 ( .A(n1258), .B(n1231), .Z(n3188) );
  CND2X2 U2900 ( .A(n3186), .B(n3187), .Z(n3189) );
  CND2X2 U2901 ( .A(n3189), .B(n3188), .Z(n4203) );
  CIVX2 U2902 ( .A(n1231), .Z(n3187) );
  CND2X1 U2903 ( .A(n4583), .B(a[16]), .Z(n3192) );
  CND2X2 U2904 ( .A(n3190), .B(n3191), .Z(n3193) );
  CND2X2 U2905 ( .A(n3192), .B(n3193), .Z(n78) );
  CIVX2 U2906 ( .A(n4583), .Z(n3190) );
  CIVX1 U2907 ( .A(a[16]), .Z(n3191) );
  CIVX3 U2908 ( .A(n4121), .Z(n4467) );
  CAN2X1 U2909 ( .A(n753), .B(n3195), .Z(n3194) );
  CIVX2 U2910 ( .A(n444), .Z(n3195) );
  CENX2 U2911 ( .A(n1381), .B(n3437), .Z(n1371) );
  CIVXL U2912 ( .A(n1167), .Z(n3197) );
  CIVX2 U2913 ( .A(n3197), .Z(n3198) );
  CEO3X1 U2914 ( .A(n1200), .B(n1175), .C(n1173), .Z(n1167) );
  CEOX2 U2915 ( .A(n1378), .B(n1384), .Z(n3199) );
  CEOX2 U2916 ( .A(n3199), .B(n1376), .Z(n1347) );
  CND2X1 U2917 ( .A(n1376), .B(n1384), .Z(n3200) );
  CND2X1 U2918 ( .A(n1376), .B(n1378), .Z(n3201) );
  CND2XL U2919 ( .A(n1384), .B(n1378), .Z(n3202) );
  CND3X1 U2920 ( .A(n3200), .B(n3201), .C(n3202), .Z(n1346) );
  CIVX1 U2921 ( .A(n3893), .Z(n3273) );
  CIVX1 U2922 ( .A(n1390), .Z(n3203) );
  CIVX2 U2923 ( .A(n3203), .Z(n3204) );
  CEOX1 U2924 ( .A(n3653), .B(n983), .Z(n979) );
  COND2XL U2925 ( .A(n90), .B(n2456), .C(net16512), .D(n2455), .Z(n1933) );
  COND2XL U2926 ( .A(n90), .B(n2453), .C(net16512), .D(n2452), .Z(n1930) );
  CENX1 U2927 ( .A(n4597), .B(n4541), .Z(n2346) );
  CENX1 U2928 ( .A(n1373), .B(n1396), .Z(n3594) );
  CND2X1 U2929 ( .A(n896), .B(n885), .Z(n3299) );
  CIVXL U2930 ( .A(n498), .Z(n3205) );
  CIVXL U2931 ( .A(n3205), .Z(n3206) );
  CEO3X1 U2932 ( .A(n2220), .B(n1766), .C(n1859), .Z(n1267) );
  CND2XL U2933 ( .A(n2220), .B(n1859), .Z(n3207) );
  CND2XL U2934 ( .A(n2220), .B(n1766), .Z(n3208) );
  CND2X1 U2935 ( .A(n1859), .B(n1766), .Z(n3209) );
  CND3X1 U2936 ( .A(n3207), .B(n3208), .C(n3209), .Z(n1266) );
  CND2X2 U2937 ( .A(n2827), .B(n6), .Z(n3210) );
  CND2X2 U2938 ( .A(n2827), .B(n6), .Z(n3211) );
  CND2X2 U2939 ( .A(n2827), .B(n6), .Z(n9) );
  CND3X1 U2940 ( .A(n3417), .B(n3418), .C(n3419), .Z(n1108) );
  CNIVX1 U2941 ( .A(n4121), .Z(n3790) );
  CIVX1 U2942 ( .A(n1247), .Z(n3680) );
  CIVX2 U2943 ( .A(n444), .Z(n3212) );
  CNR2IX2 U2944 ( .B(n754), .A(n3213), .Z(n3420) );
  CND2X2 U2945 ( .A(n753), .B(n3212), .Z(n3213) );
  CIVXL U2946 ( .A(n528), .Z(n3214) );
  CND2X2 U2947 ( .A(n1250), .B(n3216), .Z(n3217) );
  CND2X1 U2948 ( .A(n1221), .B(n3215), .Z(n3218) );
  CND2X2 U2949 ( .A(n3217), .B(n3218), .Z(n3704) );
  CIVX1 U2950 ( .A(n1250), .Z(n3215) );
  CIVX2 U2951 ( .A(n1221), .Z(n3216) );
  CND2X1 U2952 ( .A(n3905), .B(n1282), .Z(n3998) );
  CENXL U2953 ( .A(n4603), .B(n4565), .Z(n2252) );
  CENXL U2954 ( .A(n4603), .B(net16104), .Z(n2255) );
  CENXL U2955 ( .A(n4603), .B(net16102), .Z(n2254) );
  CENXL U2956 ( .A(n4603), .B(n4563), .Z(n2256) );
  CENXL U2957 ( .A(n4603), .B(n4560), .Z(n2260) );
  CENXL U2958 ( .A(n4603), .B(n4561), .Z(n2259) );
  CND2IXL U2959 ( .B(n3244), .A(n4603), .Z(n2284) );
  CENXL U2960 ( .A(n4569), .B(n4603), .Z(n2279) );
  CIVXL U2961 ( .A(n1080), .Z(n1081) );
  CND2X1 U2962 ( .A(n3527), .B(net18689), .Z(n3222) );
  CND2X2 U2963 ( .A(n3220), .B(n3221), .Z(n3223) );
  CIVX2 U2964 ( .A(n3527), .Z(n3220) );
  CIVX1 U2965 ( .A(net18689), .Z(n3221) );
  CND2X1 U2966 ( .A(n1171), .B(n1198), .Z(n3434) );
  CND2X1 U2967 ( .A(n1196), .B(n1171), .Z(n3432) );
  CEO3X2 U2968 ( .A(n1020), .B(n1018), .C(n1001), .Z(n997) );
  CEOX2 U2969 ( .A(n999), .B(n1016), .Z(n3224) );
  CEOX2 U2970 ( .A(n3224), .B(n997), .Z(n995) );
  CND2X1 U2971 ( .A(n1020), .B(n1018), .Z(n3225) );
  CND2X1 U2972 ( .A(n1020), .B(n1001), .Z(n3226) );
  CND2X2 U2973 ( .A(n1018), .B(n1001), .Z(n3227) );
  CND3X2 U2974 ( .A(n3225), .B(n3226), .C(n3227), .Z(n996) );
  CND2XL U2975 ( .A(n999), .B(n1016), .Z(n3228) );
  CND2XL U2976 ( .A(n999), .B(n997), .Z(n3229) );
  CND2XL U2977 ( .A(n1016), .B(n997), .Z(n3230) );
  CND3X1 U2978 ( .A(n3228), .B(n3229), .C(n3230), .Z(n994) );
  CEO3XL U2979 ( .A(n1605), .B(n1616), .C(n1603), .Z(n1599) );
  CND2X1 U2980 ( .A(n1063), .B(n1084), .Z(n3232) );
  CND2X2 U2981 ( .A(n3232), .B(n3233), .Z(n4042) );
  CIVX1 U2982 ( .A(n1084), .Z(n3231) );
  CENX2 U2983 ( .A(n4042), .B(n1061), .Z(n1059) );
  CIVX2 U2984 ( .A(n469), .Z(n467) );
  CENXL U2985 ( .A(n3078), .B(n4553), .Z(n2432) );
  CIVX3 U2986 ( .A(n4593), .Z(n3877) );
  CIVX1 U2987 ( .A(n1110), .Z(net18561) );
  COND1XL U2988 ( .A(n530), .B(n522), .C(n523), .Z(n3234) );
  CND2X1 U2989 ( .A(n1254), .B(n3949), .Z(n3237) );
  CND2X2 U2990 ( .A(n3235), .B(n3236), .Z(n3238) );
  CND2X2 U2991 ( .A(n3237), .B(n3238), .Z(n1221) );
  CIVX2 U2992 ( .A(n3949), .Z(n3235) );
  CIVXL U2993 ( .A(n1254), .Z(n3236) );
  CIVX3 U2994 ( .A(n4599), .Z(n4597) );
  CIVXL U2995 ( .A(n3520), .Z(n3239) );
  CIVX12 U2996 ( .A(n4604), .Z(n4603) );
  CEOX2 U2997 ( .A(n1179), .B(n1177), .Z(n3240) );
  CEOX2 U2998 ( .A(n3240), .B(n1202), .Z(n1169) );
  CND2XL U2999 ( .A(n1202), .B(n1177), .Z(n3241) );
  CND2X1 U3000 ( .A(n1202), .B(n1179), .Z(n3242) );
  CND2XL U3001 ( .A(n1177), .B(n1179), .Z(n3243) );
  CND3X1 U3002 ( .A(n3241), .B(n3242), .C(n3243), .Z(n1168) );
  CND3X1 U3003 ( .A(n3922), .B(n3923), .C(n3924), .Z(n1202) );
  CIVX4 U3004 ( .A(net18548), .Z(n3277) );
  CANR1X1 U3005 ( .A(n646), .B(n4481), .C(n639), .Z(n637) );
  CIVX4 U3006 ( .A(n4500), .Z(n4506) );
  CND3X1 U3007 ( .A(n4176), .B(n4177), .C(n4178), .Z(n1592) );
  CIVX3 U3008 ( .A(n3659), .Z(n4573) );
  CIVX2 U3009 ( .A(n12), .Z(n3658) );
  CENX1 U3010 ( .A(n593), .B(n186), .Z(product[26]) );
  COND1X1 U3011 ( .A(n594), .B(n611), .C(n3773), .Z(n593) );
  CIVX2 U3012 ( .A(n3896), .Z(n611) );
  CIVX4 U3013 ( .A(n3749), .Z(n3244) );
  CIVX2 U3014 ( .A(n3749), .Z(n3751) );
  CAOR1X1 U3015 ( .A(n3996), .B(n669), .C(n670), .Z(n4465) );
  CANR1XL U3016 ( .A(n4492), .B(n707), .C(n704), .Z(n3245) );
  CANR1XL U3017 ( .A(n4492), .B(n707), .C(n704), .Z(n3246) );
  CANR1X1 U3018 ( .A(n4492), .B(n707), .C(n704), .Z(n702) );
  COND2X1 U3019 ( .A(net18772), .B(n2685), .C(net17297), .D(n2684), .Z(n2159)
         );
  CND2X1 U3020 ( .A(n1466), .B(n1443), .Z(n4196) );
  COND2XL U3021 ( .A(n90), .B(n4208), .C(n2482), .D(net16511), .Z(n1730) );
  CENXL U3022 ( .A(n3760), .B(n4552), .Z(n2499) );
  CIVX2 U3023 ( .A(n1279), .Z(n3580) );
  CND2IXL U3024 ( .B(n1728), .A(n2138), .Z(n3976) );
  COR2X1 U3025 ( .A(n1580), .B(n1563), .Z(n3490) );
  CIVXL U3026 ( .A(n4086), .Z(n4332) );
  CIVX2 U3027 ( .A(n120), .Z(n4599) );
  COR2X1 U3028 ( .A(n81), .B(n2507), .Z(n4303) );
  CENX1 U3029 ( .A(n4122), .B(n3247), .Z(product[38]) );
  CAN2XL U3030 ( .A(n494), .B(n3756), .Z(n3247) );
  CND3X1 U3031 ( .A(n3630), .B(n3631), .C(n3632), .Z(n1478) );
  CANR1X2 U3032 ( .A(n658), .B(n4465), .C(n3989), .Z(n657) );
  CIVX3 U3033 ( .A(n4462), .Z(n4500) );
  CND2XL U3034 ( .A(n2045), .B(n2107), .Z(n3701) );
  COND1X1 U3035 ( .A(n3556), .B(n545), .C(net16270), .Z(n3250) );
  COND1XL U3036 ( .A(n3556), .B(n545), .C(net16270), .Z(n513) );
  CND3X2 U3037 ( .A(n4170), .B(n4171), .C(n4172), .Z(n1332) );
  CEOX2 U3038 ( .A(n4299), .B(n1468), .Z(n1441) );
  CEOX2 U3039 ( .A(n1445), .B(n1447), .Z(n4299) );
  CENX1 U3040 ( .A(net18614), .B(n3251), .Z(product[28]) );
  CND2X1 U3041 ( .A(n766), .B(n573), .Z(n3251) );
  CND2XL U3042 ( .A(n2200), .B(n2140), .Z(n3799) );
  CND2XL U3043 ( .A(n1925), .B(n2140), .Z(n3798) );
  CENX2 U3044 ( .A(n170), .B(n459), .Z(product[42]) );
  CENX2 U3045 ( .A(n3533), .B(n3760), .Z(n3252) );
  CENX2 U3046 ( .A(n3533), .B(n3760), .Z(n2819) );
  CENX1 U3047 ( .A(n3253), .B(n1320), .Z(n1285) );
  CENX1 U3048 ( .A(n1301), .B(n1297), .Z(n3253) );
  CND2X1 U3049 ( .A(n754), .B(n753), .Z(n3254) );
  CIVX2 U3050 ( .A(n471), .Z(n754) );
  CEOX1 U3051 ( .A(n4465), .B(n4472), .Z(product[15]) );
  CAN2XL U3052 ( .A(n2192), .B(n1725), .Z(n3255) );
  CNIVX2 U3053 ( .A(n1111), .Z(n3256) );
  CND3X2 U3054 ( .A(n4134), .B(n4135), .C(n4136), .Z(n3487) );
  COR2X1 U3055 ( .A(n939), .B(n956), .Z(n3257) );
  CEO3X2 U3056 ( .A(n3154), .B(n1941), .C(n1910), .Z(n3906) );
  CEO3X1 U3057 ( .A(n1571), .B(n1584), .C(n1569), .Z(n1565) );
  CND2XL U3058 ( .A(n1571), .B(n1569), .Z(n3258) );
  CND2X1 U3059 ( .A(n1571), .B(n1584), .Z(n3259) );
  CND2X1 U3060 ( .A(n1569), .B(n1584), .Z(n3260) );
  CND3X2 U3061 ( .A(n3258), .B(n3259), .C(n3260), .Z(n1564) );
  CND2X1 U3062 ( .A(n1549), .B(n1564), .Z(n4391) );
  CND2X1 U3063 ( .A(n4599), .B(a[28]), .Z(n3263) );
  CND2X2 U3064 ( .A(n3261), .B(n3262), .Z(n3264) );
  CND2X4 U3065 ( .A(n3263), .B(n3264), .Z(net18824) );
  CIVX2 U3066 ( .A(n4599), .Z(n3261) );
  CIVX1 U3067 ( .A(a[28]), .Z(n3262) );
  CND2XL U3068 ( .A(n4085), .B(n2809), .Z(n4333) );
  CENXL U3069 ( .A(n4086), .B(n4545), .Z(n2473) );
  COR2X1 U3070 ( .A(n4461), .B(n2718), .Z(n4246) );
  CND2XL U3071 ( .A(n4582), .B(n4559), .Z(n3266) );
  CND2XL U3072 ( .A(n3646), .B(n3265), .Z(n3267) );
  CND2X1 U3073 ( .A(n3266), .B(n3267), .Z(n2525) );
  CIVXL U3074 ( .A(n4559), .Z(n3265) );
  CIVX1 U3075 ( .A(n416), .Z(n418) );
  CIVX1 U3076 ( .A(net18718), .Z(net15910) );
  CND3X2 U3077 ( .A(n3356), .B(n3358), .C(n3357), .Z(n1018) );
  CND3X4 U3078 ( .A(n4293), .B(n4295), .C(n4294), .Z(n1086) );
  CND2IX1 U3079 ( .B(n3728), .A(n3993), .Z(n3994) );
  CIVX1 U3080 ( .A(a[10]), .Z(n3728) );
  CND2XL U3081 ( .A(n4359), .B(n4360), .Z(n3269) );
  CND2X1 U3082 ( .A(n4357), .B(n4358), .Z(n4360) );
  CND2XL U3083 ( .A(n1268), .B(n1272), .Z(n3694) );
  CND2IX1 U3084 ( .B(n1112), .A(net18199), .Z(n4201) );
  CAN2XL U3085 ( .A(n754), .B(n472), .Z(net19060) );
  CEO3X1 U3086 ( .A(n1622), .B(n1624), .C(n1620), .Z(n1603) );
  CND2XL U3087 ( .A(n1622), .B(n1620), .Z(n3270) );
  CND2XL U3088 ( .A(n1622), .B(n1624), .Z(n3271) );
  CND2X1 U3089 ( .A(n1620), .B(n1624), .Z(n3272) );
  CND3X1 U3090 ( .A(n3270), .B(n3271), .C(n3272), .Z(n1602) );
  CND2XL U3091 ( .A(n3893), .B(n4542), .Z(n3275) );
  CND2X2 U3092 ( .A(n3273), .B(n3274), .Z(n3276) );
  CND2X2 U3093 ( .A(n3275), .B(n3276), .Z(n2608) );
  CIVXL U3094 ( .A(n4542), .Z(n3274) );
  CND2X4 U3095 ( .A(net16510), .B(n2818), .Z(n3991) );
  COND2XL U3096 ( .A(n4064), .B(n2644), .C(net18914), .D(n2643), .Z(n2119) );
  CIVX1 U3097 ( .A(n39), .Z(n4094) );
  CENX1 U3098 ( .A(n4567), .B(n3893), .Z(n2611) );
  CENX1 U3099 ( .A(n4597), .B(n2809), .Z(n2347) );
  CND2X1 U3100 ( .A(n1009), .B(n1007), .Z(n3687) );
  COND2XL U3101 ( .A(net18772), .B(n2710), .C(net17297), .D(n2709), .Z(n2184)
         );
  COND2XL U3102 ( .A(net18772), .B(n2708), .C(net16451), .D(n2707), .Z(n2182)
         );
  CAOR1XL U3103 ( .A(net17297), .B(n27), .C(n2681), .Z(n2156) );
  CND2X1 U3104 ( .A(n1288), .B(n1261), .Z(n3407) );
  CND2X2 U3105 ( .A(n3651), .B(n3652), .Z(n2685) );
  CND2X1 U3106 ( .A(n1112), .B(n1110), .Z(net17759) );
  CENX1 U3107 ( .A(n3747), .B(n3893), .Z(n2613) );
  CEO3X1 U3108 ( .A(n1488), .B(n1467), .C(n1486), .Z(n1463) );
  CND2X1 U3109 ( .A(n1270), .B(n1272), .Z(n3693) );
  CND2X1 U3110 ( .A(n1270), .B(n1268), .Z(n3692) );
  CEOX1 U3111 ( .A(n1797), .B(n2036), .Z(n3278) );
  CEOX1 U3112 ( .A(n3278), .B(n1828), .Z(n1269) );
  CND2X1 U3113 ( .A(n1828), .B(n2036), .Z(n3279) );
  CND2X1 U3114 ( .A(n1828), .B(n1797), .Z(n3280) );
  CND2X1 U3115 ( .A(n2036), .B(n1797), .Z(n3281) );
  CND3X2 U3116 ( .A(n3279), .B(n3280), .C(n3281), .Z(n1268) );
  CENX1 U3117 ( .A(net15974), .B(n2785), .Z(n2653) );
  CEO3X2 U3118 ( .A(n933), .B(n931), .C(n946), .Z(n927) );
  CND2X1 U3119 ( .A(n933), .B(n931), .Z(n3282) );
  CND2XL U3120 ( .A(n933), .B(n946), .Z(n3283) );
  CND2X1 U3121 ( .A(n931), .B(n946), .Z(n3284) );
  CND3X2 U3122 ( .A(n3282), .B(n3283), .C(n3284), .Z(n926) );
  CEOX2 U3123 ( .A(n928), .B(n913), .Z(n3285) );
  CEOX2 U3124 ( .A(n3285), .B(n926), .Z(n909) );
  CND2XL U3125 ( .A(n928), .B(n913), .Z(n3286) );
  CND2XL U3126 ( .A(n928), .B(n926), .Z(n3287) );
  CND2XL U3127 ( .A(n913), .B(n926), .Z(n3288) );
  CND3X1 U3128 ( .A(n3286), .B(n3287), .C(n3288), .Z(n908) );
  CENX1 U3129 ( .A(n1075), .B(n1073), .Z(n3333) );
  CENX1 U3130 ( .A(net16541), .B(n4554), .Z(n2695) );
  CENX1 U3131 ( .A(n4592), .B(n4548), .Z(n2437) );
  CIVX3 U3132 ( .A(n3718), .Z(n4592) );
  CENX1 U3133 ( .A(n4592), .B(n4547), .Z(n2438) );
  CIVX1 U3134 ( .A(n4238), .Z(n4075) );
  CNR2X1 U3135 ( .A(n594), .B(n4155), .Z(n576) );
  CIVXL U3136 ( .A(n1415), .Z(n3289) );
  CEO3X1 U3137 ( .A(n1442), .B(n1419), .C(n1440), .Z(n1415) );
  COND1X2 U3138 ( .A(n628), .B(n622), .C(n623), .Z(n621) );
  CNR2X2 U3139 ( .A(n1483), .B(n1504), .Z(n4269) );
  CIVX3 U3140 ( .A(n4183), .Z(n4184) );
  CND2X1 U3141 ( .A(n4091), .B(n4092), .Z(n2003) );
  CENX1 U3142 ( .A(n1096), .B(n3333), .Z(n1067) );
  CIVX1 U3143 ( .A(n2082), .Z(n3291) );
  CIVX2 U3144 ( .A(n3291), .Z(n3292) );
  CIVXL U3145 ( .A(n1425), .Z(n3293) );
  CIVX1 U3146 ( .A(n3293), .Z(n3294) );
  CEO3X1 U3147 ( .A(n1452), .B(n1450), .C(n1456), .Z(n1425) );
  CIVXL U3148 ( .A(n3086), .Z(net16497) );
  CIVXL U3149 ( .A(n4601), .Z(n4463) );
  CIVXL U3150 ( .A(n4600), .Z(n4342) );
  CENX2 U3151 ( .A(n3295), .B(n3219), .Z(n1109) );
  CENX1 U3152 ( .A(n1138), .B(n1113), .Z(n3295) );
  CIVX3 U3153 ( .A(n3807), .Z(net18896) );
  CENX1 U3154 ( .A(n3908), .B(n4559), .Z(n2657) );
  CND2X1 U3155 ( .A(n1277), .B(n3249), .Z(n4382) );
  CENX1 U3156 ( .A(n4085), .B(n4546), .Z(n2472) );
  CND2X1 U3157 ( .A(n1522), .B(n1518), .Z(n3863) );
  CENX1 U3158 ( .A(net17419), .B(n4554), .Z(n2398) );
  COND1XL U3159 ( .A(n700), .B(n3246), .C(n701), .Z(n3296) );
  CANR1XL U3160 ( .A(n4485), .B(n4493), .C(n712), .Z(n3297) );
  COND1X1 U3161 ( .A(n700), .B(n702), .C(n701), .Z(n699) );
  CANR1X1 U3162 ( .A(n4485), .B(n4493), .C(n712), .Z(n710) );
  COR2XL U3163 ( .A(net17279), .B(n2541), .Z(n3983) );
  COND2XL U3164 ( .A(n3133), .B(n2547), .C(n3121), .D(n2546), .Z(n2024) );
  CND2X2 U3165 ( .A(n1093), .B(n1114), .Z(n4294) );
  CENX1 U3166 ( .A(n4580), .B(n4560), .Z(n2557) );
  CIVX8 U3167 ( .A(n111), .Z(n4596) );
  CND2X1 U3168 ( .A(n896), .B(n898), .Z(n3298) );
  CND2XL U3169 ( .A(n898), .B(n885), .Z(n3300) );
  CND2X2 U3170 ( .A(n3095), .B(n3084), .Z(n3301) );
  CND2X2 U3171 ( .A(n4310), .B(n105), .Z(n3302) );
  CND2X1 U3172 ( .A(n3095), .B(n3084), .Z(net17727) );
  CAN2X1 U3173 ( .A(n4373), .B(n3762), .Z(n690) );
  CND2X4 U3174 ( .A(n24), .B(n2825), .Z(n27) );
  CND2X1 U3175 ( .A(n1590), .B(n1577), .Z(n3305) );
  CND2X2 U3176 ( .A(n3303), .B(n3304), .Z(n3306) );
  CND2X2 U3177 ( .A(n3305), .B(n3306), .Z(n3912) );
  CIVX1 U3178 ( .A(n1590), .Z(n3303) );
  CIVX1 U3179 ( .A(n1577), .Z(n3304) );
  COND2X1 U3180 ( .A(net18772), .B(n2700), .C(net16451), .D(n2699), .Z(n2174)
         );
  CENX1 U3181 ( .A(n3893), .B(n4543), .Z(n2607) );
  CIVX2 U3182 ( .A(net18218), .Z(net16419) );
  CIVXL U3183 ( .A(n1239), .Z(n3307) );
  CIVXL U3184 ( .A(n3307), .Z(n3308) );
  CENX2 U3185 ( .A(net18420), .B(n4577), .Z(n3309) );
  CENX1 U3186 ( .A(net18420), .B(n4577), .Z(n3310) );
  CENX2 U3187 ( .A(net18420), .B(n4577), .Z(n2823) );
  CND2X1 U3188 ( .A(n1280), .B(n1255), .Z(n4000) );
  CIVX3 U3189 ( .A(n4311), .Z(n4598) );
  CND2X1 U3190 ( .A(n4575), .B(n4561), .Z(n3313) );
  CND2X1 U3191 ( .A(n3311), .B(n3312), .Z(n3314) );
  CND2X2 U3192 ( .A(n3313), .B(n3314), .Z(n2622) );
  CIVX1 U3193 ( .A(n4575), .Z(n3311) );
  CIVXL U3194 ( .A(n4561), .Z(n3312) );
  CND2XL U3195 ( .A(n1134), .B(n1109), .Z(n3710) );
  CND2X1 U3196 ( .A(n1164), .B(n1162), .Z(n3935) );
  CND2XL U3197 ( .A(n1242), .B(n2188), .Z(n3928) );
  CND2XL U3198 ( .A(n1242), .B(n2096), .Z(n3929) );
  CND2XL U3199 ( .A(n4580), .B(n2785), .Z(n3317) );
  CND2X1 U3200 ( .A(n3315), .B(n3316), .Z(n3318) );
  CND2X2 U3201 ( .A(n3317), .B(n3318), .Z(n2554) );
  CIVXL U3202 ( .A(n4580), .Z(n3315) );
  CIVXL U3203 ( .A(n2785), .Z(n3316) );
  CIVXL U3204 ( .A(n1462), .Z(n3319) );
  CIVXL U3205 ( .A(n3319), .Z(n3320) );
  CEO3X1 U3206 ( .A(n1536), .B(n1521), .C(n1523), .Z(n1513) );
  CND2XL U3207 ( .A(n1536), .B(n1521), .Z(n3321) );
  CND2XL U3208 ( .A(n1536), .B(n1523), .Z(n3322) );
  CND2X1 U3209 ( .A(n1521), .B(n1523), .Z(n3323) );
  CND3X1 U3210 ( .A(n3321), .B(n3322), .C(n3323), .Z(n1512) );
  CEOX2 U3211 ( .A(n1510), .B(n1493), .Z(n3324) );
  CEOX2 U3212 ( .A(n3324), .B(n1512), .Z(n1487) );
  CND2X1 U3213 ( .A(n1510), .B(n1493), .Z(n3325) );
  CND2X1 U3214 ( .A(n1510), .B(n1512), .Z(n3326) );
  CND2X2 U3215 ( .A(n1493), .B(n1512), .Z(n3327) );
  CND3X2 U3216 ( .A(n3325), .B(n3326), .C(n3327), .Z(n1486) );
  CENX2 U3217 ( .A(n1137), .B(n3487), .Z(n4242) );
  CENX1 U3218 ( .A(n4595), .B(n4544), .Z(n2375) );
  CIVX1 U3219 ( .A(net18218), .Z(n3329) );
  CNR2XL U3220 ( .A(n1083), .B(n1106), .Z(n3330) );
  CNR2XL U3221 ( .A(n1083), .B(n1106), .Z(n3331) );
  CIVXL U3222 ( .A(net18199), .Z(n3332) );
  CNR2XL U3223 ( .A(n1083), .B(n1106), .Z(n491) );
  CENX1 U3224 ( .A(net16541), .B(net16102), .Z(n2683) );
  CND2X1 U3225 ( .A(n2197), .B(n2228), .Z(n4119) );
  CENX1 U3226 ( .A(n4582), .B(n4556), .Z(n2528) );
  CENX1 U3227 ( .A(n1309), .B(n1334), .Z(n3657) );
  CENX2 U3228 ( .A(n1315), .B(n1338), .Z(n3401) );
  COND2X1 U3229 ( .A(n63), .B(n2565), .C(n2564), .D(n4505), .Z(n2040) );
  CENX2 U3230 ( .A(n3334), .B(n1312), .Z(n1279) );
  CENX2 U3231 ( .A(n1285), .B(n1310), .Z(n3334) );
  CIVXL U3232 ( .A(n708), .Z(n788) );
  CEO3XL U3233 ( .A(n1702), .B(n1695), .C(n1697), .Z(n3335) );
  CND2X1 U3234 ( .A(n3841), .B(n1422), .Z(n3338) );
  CND2X2 U3235 ( .A(n3336), .B(n3337), .Z(n3339) );
  CND2X2 U3236 ( .A(n3338), .B(n3339), .Z(n1393) );
  CIVX2 U3237 ( .A(n3841), .Z(n3336) );
  CIVXL U3238 ( .A(n1422), .Z(n3337) );
  CIVXL U3239 ( .A(n3727), .Z(n3340) );
  CEO3X1 U3240 ( .A(n2029), .B(n1820), .C(n1937), .Z(n1055) );
  CND2XL U3241 ( .A(n2029), .B(n1820), .Z(n3341) );
  CND2XL U3242 ( .A(n2029), .B(n1937), .Z(n3342) );
  CND2XL U3243 ( .A(n1820), .B(n1937), .Z(n3343) );
  CND3X1 U3244 ( .A(n3341), .B(n3342), .C(n3343), .Z(n1054) );
  CEOX2 U3245 ( .A(n1050), .B(n1052), .Z(n3344) );
  CEOX2 U3246 ( .A(n3344), .B(n1054), .Z(n1025) );
  CND2X1 U3247 ( .A(n1050), .B(n1052), .Z(n3345) );
  CND2X1 U3248 ( .A(n1050), .B(n1054), .Z(n3346) );
  CND2X1 U3249 ( .A(n1052), .B(n1054), .Z(n3347) );
  CND3X2 U3250 ( .A(n3345), .B(n3346), .C(n3347), .Z(n1024) );
  COR2XL U3251 ( .A(n2460), .B(n3991), .Z(n3348) );
  COR2XL U3252 ( .A(net16512), .B(n2459), .Z(n3349) );
  CND2X1 U3253 ( .A(n3348), .B(n3349), .Z(n1937) );
  CNIVX1 U3254 ( .A(n4566), .Z(n3746) );
  CENX1 U3255 ( .A(n4568), .B(net17419), .Z(n2411) );
  CENX1 U3256 ( .A(n3908), .B(n4552), .Z(n2664) );
  CND2X2 U3257 ( .A(n3679), .B(n3680), .Z(n3682) );
  CENX2 U3258 ( .A(n3350), .B(n3906), .Z(n1145) );
  CENX2 U3259 ( .A(n1180), .B(n1157), .Z(n3350) );
  CENXL U3260 ( .A(n4598), .B(n4558), .Z(n2328) );
  CENXL U3261 ( .A(n4598), .B(n4544), .Z(n2342) );
  CENXL U3262 ( .A(n4598), .B(n4553), .Z(n2333) );
  CENXL U3263 ( .A(n4598), .B(n4552), .Z(n2334) );
  CENXL U3264 ( .A(n4569), .B(n4598), .Z(n2345) );
  CND3X2 U3265 ( .A(n3793), .B(n3794), .C(n3795), .Z(n1482) );
  CENXL U3266 ( .A(net15910), .B(n4557), .Z(n2395) );
  CENXL U3267 ( .A(net15910), .B(n4558), .Z(n2394) );
  CENXL U3268 ( .A(net15910), .B(n4544), .Z(n2408) );
  CND2XL U3269 ( .A(net15910), .B(n4559), .Z(n3838) );
  CENXL U3270 ( .A(net15910), .B(n4560), .Z(n2392) );
  CND2X1 U3271 ( .A(n3595), .B(n498), .Z(n3397) );
  CENX1 U3272 ( .A(net16541), .B(n4562), .Z(n2687) );
  CIVX4 U3273 ( .A(net15912), .Z(net18211) );
  CIVXL U3274 ( .A(n1260), .Z(n3351) );
  CIVX1 U3275 ( .A(n3351), .Z(n3352) );
  CND2X1 U3276 ( .A(n1226), .B(n1224), .Z(n4113) );
  CIVX4 U3277 ( .A(a[16]), .Z(n3533) );
  CIVXL U3278 ( .A(n3254), .Z(n3353) );
  CIVX1 U3279 ( .A(n3353), .Z(n3354) );
  CIVX1 U3280 ( .A(net16541), .Z(n3649) );
  CEO3X2 U3281 ( .A(n1222), .B(n1195), .C(n1197), .Z(n1191) );
  CENX1 U3282 ( .A(net16541), .B(n4544), .Z(n2705) );
  CIVX1 U3283 ( .A(net15914), .Z(net18209) );
  CEOX2 U3284 ( .A(n1025), .B(n1044), .Z(n3355) );
  CEOX2 U3285 ( .A(n3355), .B(n1023), .Z(n1019) );
  CND2X1 U3286 ( .A(n1023), .B(n1044), .Z(n3356) );
  CND2X1 U3287 ( .A(n1023), .B(n1025), .Z(n3357) );
  CND2XL U3288 ( .A(n1044), .B(n1025), .Z(n3358) );
  CND2X1 U3289 ( .A(n1471), .B(n1490), .Z(n3636) );
  CAOR1XL U3290 ( .A(n3667), .B(n117), .C(n2351), .Z(n1835) );
  COND2XL U3291 ( .A(n117), .B(n2355), .C(n3667), .D(n2354), .Z(n1839) );
  COND2XL U3292 ( .A(n117), .B(n2354), .C(n3667), .D(n2353), .Z(n1838) );
  CND3X2 U3293 ( .A(n4286), .B(n4287), .C(n4288), .Z(n1530) );
  CENX1 U3294 ( .A(n4585), .B(n4564), .Z(n2484) );
  CIVXL U3295 ( .A(n1479), .Z(n3359) );
  CIVXL U3296 ( .A(n3359), .Z(n3360) );
  COAN1X1 U3297 ( .A(n487), .B(n545), .C(n488), .Z(n4474) );
  CANR1X1 U3298 ( .A(n489), .B(n517), .C(n490), .Z(n488) );
  CEOX2 U3299 ( .A(n1051), .B(n1057), .Z(n3361) );
  CEOX2 U3300 ( .A(n3361), .B(n1053), .Z(n1045) );
  CND2X1 U3301 ( .A(n1053), .B(n1057), .Z(n3362) );
  CND2XL U3302 ( .A(n1053), .B(n1051), .Z(n3363) );
  CND2XL U3303 ( .A(n1057), .B(n1051), .Z(n3364) );
  CND3X1 U3304 ( .A(n3362), .B(n3363), .C(n3364), .Z(n1044) );
  CND3X1 U3305 ( .A(n4524), .B(n4525), .C(n4526), .Z(n3366) );
  CND3X2 U3306 ( .A(n3686), .B(n3687), .C(n3688), .Z(n1002) );
  CANR1X1 U3307 ( .A(n419), .B(n387), .C(n388), .Z(n386) );
  COND2XL U3308 ( .A(n54), .B(n3993), .C(n2614), .D(n4507), .Z(n1734) );
  CND3XL U3309 ( .A(n4537), .B(n4538), .C(n4539), .Z(n3365) );
  CENX2 U3310 ( .A(n1342), .B(n1319), .Z(n3776) );
  CND2X1 U3311 ( .A(n1240), .B(n2065), .Z(n3924) );
  CEO3X2 U3312 ( .A(n1472), .B(n1449), .C(n1470), .Z(n1443) );
  CEO3X1 U3313 ( .A(n1194), .B(n1169), .C(n3198), .Z(n1163) );
  CND2X1 U3314 ( .A(n307), .B(n739), .Z(n298) );
  CND2XL U3315 ( .A(n4512), .B(n4558), .Z(n3369) );
  CND2X1 U3316 ( .A(n3367), .B(n3368), .Z(n3370) );
  CND2X1 U3317 ( .A(n3369), .B(n3370), .Z(n2724) );
  CIVXL U3318 ( .A(n4512), .Z(n3367) );
  CIVXL U3319 ( .A(n4558), .Z(n3368) );
  CND3XL U3320 ( .A(n4000), .B(n3998), .C(n3999), .Z(n3371) );
  CIVXL U3321 ( .A(n639), .Z(n3372) );
  CEOX2 U3322 ( .A(n1405), .B(n1407), .Z(n3373) );
  CND2XL U3323 ( .A(n1407), .B(n1405), .Z(n3376) );
  CND3X1 U3324 ( .A(n3374), .B(n3375), .C(n3376), .Z(n1394) );
  CND2XL U3325 ( .A(n2074), .B(n2136), .Z(n3377) );
  CND2X1 U3326 ( .A(n2074), .B(n2105), .Z(n3378) );
  CND2X1 U3327 ( .A(n2136), .B(n2105), .Z(n3379) );
  CND3X2 U3328 ( .A(n3377), .B(n3378), .C(n3379), .Z(n1450) );
  CFA1X1 U3329 ( .A(n1864), .B(n3755), .CI(n2194), .CO(n1406), .S(n1407) );
  CEOX2 U3330 ( .A(n3640), .B(n1662), .Z(n1647) );
  CIVXL U3331 ( .A(n3296), .Z(n698) );
  CENXL U3332 ( .A(n4085), .B(n4542), .Z(n2476) );
  CND2X4 U3333 ( .A(n3831), .B(n3832), .Z(n3380) );
  CND2X2 U3334 ( .A(n3831), .B(n3832), .Z(net16959) );
  CEO3X2 U3335 ( .A(n1555), .B(n3063), .C(n1570), .Z(n1549) );
  CND2X1 U3336 ( .A(n3062), .B(n1570), .Z(n3381) );
  CND2X1 U3337 ( .A(n1568), .B(n1555), .Z(n3382) );
  CND2X2 U3338 ( .A(n1570), .B(n1555), .Z(n3383) );
  CND3X2 U3339 ( .A(n3381), .B(n3382), .C(n3383), .Z(n1548) );
  COR2X1 U3340 ( .A(n3117), .B(n2526), .Z(n4091) );
  CEO3X2 U3341 ( .A(n1411), .B(n3778), .C(n1434), .Z(n1401) );
  CND2XL U3342 ( .A(n1411), .B(n1434), .Z(n3384) );
  CND2XL U3343 ( .A(n1411), .B(n3778), .Z(n3385) );
  CND2X1 U3344 ( .A(n1434), .B(n3778), .Z(n3386) );
  CND3X1 U3345 ( .A(n3384), .B(n3385), .C(n3386), .Z(n1400) );
  CEO3X1 U3346 ( .A(n1383), .B(n1398), .C(n1400), .Z(n1369) );
  CND2XL U3347 ( .A(n1383), .B(n1398), .Z(n3387) );
  CND2X1 U3348 ( .A(n1383), .B(n1400), .Z(n3388) );
  CND2XL U3349 ( .A(n1398), .B(n1400), .Z(n3389) );
  CND3X1 U3350 ( .A(n3387), .B(n3388), .C(n3389), .Z(n1368) );
  CEOX2 U3351 ( .A(n3390), .B(n1368), .Z(n1337) );
  CND2X1 U3352 ( .A(n1343), .B(n1368), .Z(n3392) );
  CNR2X2 U3353 ( .A(n3116), .B(n4321), .Z(n3394) );
  CNR2XL U3354 ( .A(n2350), .B(n123), .Z(n3395) );
  COR2X1 U3355 ( .A(n3394), .B(n3395), .Z(n1726) );
  CENX2 U3356 ( .A(a[26]), .B(n4596), .Z(n3396) );
  CNIVX1 U3357 ( .A(n2012), .Z(n3778) );
  CND2IXL U3358 ( .B(n3244), .A(n4598), .Z(n2350) );
  CIVX4 U3359 ( .A(n3396), .Z(n123) );
  CENX2 U3360 ( .A(a[26]), .B(n4596), .Z(n3907) );
  CND2X1 U3361 ( .A(n1469), .B(n1490), .Z(n3635) );
  CNR2X1 U3362 ( .A(n409), .B(n402), .Z(n396) );
  CEO3X1 U3363 ( .A(n2062), .B(n1823), .C(n1854), .Z(n1125) );
  CND2XL U3364 ( .A(n2062), .B(n1854), .Z(n3398) );
  CND2X1 U3365 ( .A(n1854), .B(n1823), .Z(n3400) );
  CND3X2 U3366 ( .A(n3398), .B(n3399), .C(n3400), .Z(n1124) );
  COND2X1 U3367 ( .A(n54), .B(n2587), .C(n4506), .D(n2586), .Z(n2062) );
  CNR2X2 U3368 ( .A(n3335), .B(n1700), .Z(n696) );
  CEO3X1 U3369 ( .A(n1509), .B(n1526), .C(n4038), .Z(n4266) );
  CENX2 U3370 ( .A(n3401), .B(n1340), .Z(n1309) );
  CEOX2 U3371 ( .A(n1617), .B(n1628), .Z(n3402) );
  CEOX2 U3372 ( .A(n3402), .B(n1615), .Z(n1613) );
  CND2XL U3373 ( .A(n1615), .B(n1628), .Z(n3403) );
  CND2XL U3374 ( .A(n1615), .B(n1617), .Z(n3404) );
  CND2XL U3375 ( .A(n1628), .B(n1617), .Z(n3405) );
  CND3X1 U3376 ( .A(n3403), .B(n3404), .C(n3405), .Z(n1612) );
  COR2X1 U3377 ( .A(n1597), .B(n1612), .Z(n4169) );
  CND2XL U3378 ( .A(n1247), .B(n1249), .Z(n4098) );
  CAOR1XL U3379 ( .A(net16438), .B(net18310), .C(n2285), .Z(n1769) );
  COND2XL U3380 ( .A(net18310), .B(n2287), .C(net16438), .D(n2286), .Z(n1771)
         );
  COND2XL U3381 ( .A(net18310), .B(n2289), .C(net16438), .D(n2288), .Z(n1773)
         );
  COND2XL U3382 ( .A(net18310), .B(n2293), .C(net16438), .D(n2292), .Z(n1777)
         );
  CNR2X1 U3383 ( .A(net18310), .B(n2316), .Z(n4277) );
  CEO3X2 U3384 ( .A(n1288), .B(n1261), .C(n1259), .Z(n1253) );
  CND2X1 U3385 ( .A(n1288), .B(n1259), .Z(n3406) );
  CND2X2 U3386 ( .A(n1259), .B(n1261), .Z(n3408) );
  CND3X2 U3387 ( .A(n3406), .B(n3407), .C(n3408), .Z(n1252) );
  COND1X1 U3388 ( .A(n530), .B(n522), .C(n523), .Z(n3409) );
  CND2X2 U3389 ( .A(n1223), .B(n1252), .Z(n4030) );
  CND2X1 U3390 ( .A(n1285), .B(n1312), .Z(n4339) );
  CEO3X2 U3391 ( .A(n2056), .B(n2179), .C(n2209), .Z(n1673) );
  CND2XL U3392 ( .A(n2056), .B(n2179), .Z(n3410) );
  CND2XL U3393 ( .A(n2056), .B(n2209), .Z(n3411) );
  CND2XL U3394 ( .A(n2179), .B(n2209), .Z(n3412) );
  CND3X1 U3395 ( .A(n3410), .B(n3411), .C(n3412), .Z(n1672) );
  CEOXL U3396 ( .A(n1663), .B(n1670), .Z(n3413) );
  CEOX1 U3397 ( .A(n3413), .B(n1672), .Z(n1657) );
  CND2X1 U3398 ( .A(n1663), .B(n1670), .Z(n3414) );
  CND2X1 U3399 ( .A(n1663), .B(n1672), .Z(n3415) );
  CND2X1 U3400 ( .A(n1670), .B(n1672), .Z(n3416) );
  CND3X1 U3401 ( .A(n3414), .B(n3415), .C(n3416), .Z(n1656) );
  CND2X1 U3402 ( .A(n1136), .B(n1138), .Z(n3418) );
  CND2XL U3403 ( .A(n1113), .B(n1138), .Z(n3419) );
  CNR2X2 U3404 ( .A(net16974), .B(net16962), .Z(n3874) );
  CENX1 U3405 ( .A(n3748), .B(n3774), .Z(n2481) );
  CIVX3 U3406 ( .A(n39), .Z(n4093) );
  CIVXL U3407 ( .A(n3196), .Z(n3421) );
  CIVX1 U3408 ( .A(n3421), .Z(n3422) );
  CND2XL U3409 ( .A(n4582), .B(n4561), .Z(n3425) );
  CND2X1 U3410 ( .A(n3423), .B(n3424), .Z(n3426) );
  CND2X1 U3411 ( .A(n3425), .B(n3426), .Z(n2523) );
  CIVXL U3412 ( .A(n4582), .Z(n3423) );
  CIVXL U3413 ( .A(n4561), .Z(n3424) );
  CAOR1XL U3414 ( .A(n4508), .B(net18627), .C(n2417), .Z(n1894) );
  COND2XL U3415 ( .A(n63), .B(n2578), .C(n2577), .D(n4505), .Z(n3427) );
  CND2X1 U3416 ( .A(n267), .B(n154), .Z(n3430) );
  CND2X2 U3417 ( .A(n3428), .B(n3429), .Z(n3431) );
  CND2X2 U3418 ( .A(n3430), .B(n3431), .Z(product[58]) );
  CIVX2 U3419 ( .A(n267), .Z(n3428) );
  CIVX2 U3420 ( .A(n154), .Z(n3429) );
  CND2XL U3421 ( .A(n975), .B(n994), .Z(n449) );
  CIVX1 U3422 ( .A(n448), .Z(n751) );
  CIVXL U3423 ( .A(n458), .Z(n456) );
  CND2X1 U3424 ( .A(n1196), .B(n1198), .Z(n3433) );
  CND3X2 U3425 ( .A(n3432), .B(n3433), .C(n3434), .Z(n1164) );
  CEOX1 U3426 ( .A(n2005), .B(n1881), .Z(n3435) );
  CEOX1 U3427 ( .A(n3435), .B(n1826), .Z(n1209) );
  CND3X1 U3428 ( .A(n4110), .B(n4111), .C(n4112), .Z(n1198) );
  CNIVX4 U3429 ( .A(n4566), .Z(n3747) );
  CENX1 U3430 ( .A(n3622), .B(n4551), .Z(n2566) );
  CNIVX2 U3431 ( .A(n1453), .Z(n3436) );
  CENXL U3432 ( .A(n4570), .B(n4541), .Z(n2775) );
  COND1XL U3433 ( .A(n633), .B(n637), .C(n634), .Z(n3788) );
  CND2X1 U3434 ( .A(n1553), .B(n1566), .Z(n4388) );
  CENX2 U3435 ( .A(n1379), .B(n1377), .Z(n3437) );
  CENX2 U3436 ( .A(n3438), .B(n1017), .Z(n1015) );
  CENX2 U3437 ( .A(n1019), .B(n1038), .Z(n3438) );
  CNR2X2 U3438 ( .A(n1059), .B(n1082), .Z(n484) );
  CND3X1 U3439 ( .A(n3524), .B(n3525), .C(n3526), .Z(n1398) );
  CND2XL U3440 ( .A(n1432), .B(n1430), .Z(n3524) );
  CIVX2 U3441 ( .A(n1224), .Z(n3604) );
  CEOX2 U3442 ( .A(n1573), .B(n1588), .Z(n3439) );
  CEOX1 U3443 ( .A(n3439), .B(n1586), .Z(n1567) );
  CND2X1 U3444 ( .A(n1586), .B(n1588), .Z(n3440) );
  CND2X1 U3445 ( .A(n1586), .B(n1573), .Z(n3441) );
  CND2XL U3446 ( .A(n1588), .B(n1573), .Z(n3442) );
  CND3X2 U3447 ( .A(n3440), .B(n3441), .C(n3442), .Z(n1566) );
  CND2X1 U3448 ( .A(n1278), .B(n1253), .Z(n3443) );
  CND2X1 U3449 ( .A(n1278), .B(n1251), .Z(n3444) );
  CND2X1 U3450 ( .A(n1253), .B(n1251), .Z(n3445) );
  CND3X2 U3451 ( .A(n3443), .B(n3444), .C(n3445), .Z(n1246) );
  CND2X2 U3452 ( .A(n1338), .B(n1340), .Z(n4161) );
  CIVX1 U3453 ( .A(n3921), .Z(n3667) );
  CND2X1 U3454 ( .A(n1221), .B(n1250), .Z(n3707) );
  CEO3X1 U3455 ( .A(n2034), .B(n1857), .C(n2127), .Z(n1207) );
  COR2XL U3456 ( .A(n995), .B(n1014), .Z(n3572) );
  CENX2 U3457 ( .A(n4234), .B(n1634), .Z(n1619) );
  CND2X1 U3458 ( .A(n393), .B(n164), .Z(n3448) );
  CND2X2 U3459 ( .A(n3446), .B(n3447), .Z(n3449) );
  CND2X2 U3460 ( .A(n3448), .B(n3449), .Z(product[48]) );
  CIVX1 U3461 ( .A(n393), .Z(n3446) );
  CIVX2 U3462 ( .A(n164), .Z(n3447) );
  CEO3X1 U3463 ( .A(n1088), .B(n1086), .C(n1065), .Z(n1061) );
  CEOX1 U3464 ( .A(n2226), .B(n2073), .Z(n3450) );
  CEOX1 U3465 ( .A(n3450), .B(n2013), .Z(n1429) );
  CND2XL U3466 ( .A(n2073), .B(n2013), .Z(n3451) );
  CND2X1 U3467 ( .A(n2013), .B(n2226), .Z(n3452) );
  CND2XL U3468 ( .A(n2073), .B(n2226), .Z(n3453) );
  CND3X1 U3469 ( .A(n3451), .B(n3452), .C(n3453), .Z(n1428) );
  CEO3X2 U3470 ( .A(n1194), .B(n1169), .C(n3198), .Z(n3454) );
  CND2IX1 U3471 ( .B(n1279), .A(n3581), .Z(n3583) );
  CND2XL U3472 ( .A(n1282), .B(n1255), .Z(n3999) );
  CENX1 U3473 ( .A(n4512), .B(n4548), .Z(n2734) );
  CIVX1 U3474 ( .A(n3749), .Z(n3750) );
  CIVX4 U3475 ( .A(n4566), .Z(n3749) );
  CAN2X1 U3476 ( .A(n1728), .B(n2138), .Z(n3758) );
  CENX2 U3477 ( .A(n1370), .B(n1347), .Z(n3463) );
  CEOX2 U3478 ( .A(n1924), .B(n2046), .Z(n3455) );
  CEOX2 U3479 ( .A(n3455), .B(n1955), .Z(n1521) );
  CND2XL U3480 ( .A(n1955), .B(n2046), .Z(n3456) );
  CND2XL U3481 ( .A(n1955), .B(n1924), .Z(n3457) );
  CND2XL U3482 ( .A(n2046), .B(n1924), .Z(n3458) );
  CND3XL U3483 ( .A(n3456), .B(n3457), .C(n3458), .Z(n1520) );
  COR2X1 U3484 ( .A(n3991), .B(n2478), .Z(n3459) );
  COR2XL U3485 ( .A(net16512), .B(n2477), .Z(n3460) );
  CND2X2 U3486 ( .A(n3459), .B(n3460), .Z(n1955) );
  CNIVX4 U3487 ( .A(n87), .Z(net16512) );
  CENX1 U3488 ( .A(n4582), .B(n4557), .Z(n2527) );
  CIVXL U3489 ( .A(n4573), .Z(n3461) );
  COND1X1 U3490 ( .A(n651), .B(n668), .C(n652), .Z(n3511) );
  CHA1X1 U3491 ( .A(n2212), .B(n1735), .CO(n1698), .S(n1699) );
  CND2X1 U3492 ( .A(n1994), .B(n1753), .Z(n3574) );
  CND2IX1 U3493 ( .B(n3580), .A(n1306), .Z(n3582) );
  CENX2 U3494 ( .A(n3912), .B(n4143), .Z(n1569) );
  CENXL U3495 ( .A(net16541), .B(n4564), .Z(n2682) );
  CENXL U3496 ( .A(net16541), .B(n4553), .Z(n2696) );
  CENXL U3497 ( .A(net16541), .B(n4551), .Z(n2698) );
  CENX1 U3498 ( .A(net16541), .B(n2785), .Z(n2686) );
  CENXL U3499 ( .A(n3077), .B(n4014), .Z(n3462) );
  CENX1 U3500 ( .A(n3077), .B(n4014), .Z(n1317) );
  CENX2 U3501 ( .A(n3463), .B(n1345), .Z(n1339) );
  CENX1 U3502 ( .A(n3886), .B(n1277), .Z(n1275) );
  CNR2X2 U3503 ( .A(n4351), .B(n616), .Z(n614) );
  CENX1 U3504 ( .A(n4512), .B(n4555), .Z(n2727) );
  CIVX4 U3505 ( .A(n3658), .Z(n4572) );
  CNR2X1 U3506 ( .A(n1215), .B(n1244), .Z(n3518) );
  COND1X1 U3507 ( .A(n547), .B(n575), .C(n3042), .Z(n3464) );
  COND1X1 U3508 ( .A(n547), .B(n575), .C(n548), .Z(n546) );
  CND2XL U3509 ( .A(n1951), .B(n1982), .Z(n4175) );
  CENX1 U3510 ( .A(n3893), .B(n4548), .Z(n2602) );
  CND2XL U3511 ( .A(n75), .B(a[18]), .Z(n3951) );
  COND1X1 U3512 ( .A(n675), .B(n671), .C(n672), .Z(n670) );
  COND2X1 U3513 ( .A(n81), .B(n2491), .C(n4217), .D(n2490), .Z(n1968) );
  COND2X1 U3514 ( .A(net17738), .B(n2348), .C(n123), .D(n2347), .Z(n1832) );
  CND2X2 U3515 ( .A(n3596), .B(n3597), .Z(n3599) );
  CIVXL U3516 ( .A(n3475), .Z(n3465) );
  CND2XL U3517 ( .A(n3645), .B(n4555), .Z(n3468) );
  CND2X1 U3518 ( .A(n3466), .B(n3467), .Z(n3469) );
  CND2X1 U3519 ( .A(n3468), .B(n3469), .Z(n2529) );
  CIVXL U3520 ( .A(n3645), .Z(n3466) );
  CIVXL U3521 ( .A(n4555), .Z(n3467) );
  CENX1 U3522 ( .A(n3470), .B(n1908), .Z(n1105) );
  CENXL U3523 ( .A(n2092), .B(n1130), .Z(n3470) );
  CEOX1 U3524 ( .A(n1006), .B(n1008), .Z(n3471) );
  CND2XL U3525 ( .A(n991), .B(n1008), .Z(n3472) );
  CND2XL U3526 ( .A(n991), .B(n1006), .Z(n3473) );
  CND2XL U3527 ( .A(n1008), .B(n1006), .Z(n3474) );
  CND3X1 U3528 ( .A(n3472), .B(n3473), .C(n3474), .Z(n982) );
  CND2XL U3529 ( .A(n4582), .B(net16104), .Z(n3477) );
  CND2X1 U3530 ( .A(n3475), .B(n3476), .Z(n3478) );
  CND2X1 U3531 ( .A(n3477), .B(n3478), .Z(n2519) );
  CIVXL U3532 ( .A(n4582), .Z(n3475) );
  CIVXL U3533 ( .A(net16104), .Z(n3476) );
  CND2XL U3534 ( .A(net16541), .B(n4559), .Z(n3481) );
  CND2X1 U3535 ( .A(n3479), .B(n3480), .Z(n3482) );
  CND2X1 U3536 ( .A(n3481), .B(n3482), .Z(n2690) );
  CIVXL U3537 ( .A(net16541), .Z(n3479) );
  CIVXL U3538 ( .A(n4559), .Z(n3480) );
  CND2X2 U3539 ( .A(n3329), .B(n3310), .Z(n45) );
  CIVX2 U3540 ( .A(n3830), .Z(n3815) );
  CND2XL U3541 ( .A(n4343), .B(net18209), .Z(n4412) );
  CND2XL U3542 ( .A(net18209), .B(n3837), .Z(n3839) );
  CEOX2 U3543 ( .A(n1945), .B(n2129), .Z(n3483) );
  CEOX2 U3544 ( .A(n3483), .B(n1914), .Z(n1265) );
  CND2XL U3545 ( .A(n1914), .B(n2129), .Z(n3484) );
  CND2XL U3546 ( .A(n1914), .B(n1945), .Z(n3485) );
  CND2XL U3547 ( .A(n2129), .B(n1945), .Z(n3486) );
  CND3X1 U3548 ( .A(n3484), .B(n3485), .C(n3486), .Z(n1264) );
  CENX2 U3549 ( .A(n1109), .B(n3489), .Z(n1107) );
  CENX2 U3550 ( .A(n3256), .B(n1134), .Z(n3489) );
  CEO3X2 U3551 ( .A(n1172), .B(n3791), .C(n1174), .Z(n3904) );
  CEOX2 U3552 ( .A(net17986), .B(net18863), .Z(n1137) );
  CENX2 U3553 ( .A(n4487), .B(n1314), .Z(n1281) );
  CND2IX1 U3554 ( .B(n643), .A(n3490), .Z(n636) );
  COND1X1 U3555 ( .A(n544), .B(n540), .C(n541), .Z(n535) );
  CENX2 U3556 ( .A(n1031), .B(n3491), .Z(n1023) );
  CENX2 U3557 ( .A(n1033), .B(n1029), .Z(n3491) );
  CEOX2 U3558 ( .A(n1102), .B(n1077), .Z(n3492) );
  CEOX2 U3559 ( .A(n3492), .B(n1079), .Z(n1069) );
  CND2XL U3560 ( .A(n1077), .B(n1079), .Z(n3493) );
  CND2X1 U3561 ( .A(n1079), .B(n1102), .Z(n3494) );
  CND2XL U3562 ( .A(n1077), .B(n1102), .Z(n3495) );
  CND3X1 U3563 ( .A(n3493), .B(n3495), .C(n3494), .Z(n1068) );
  CIVX3 U3564 ( .A(n3659), .Z(n4512) );
  CND2XL U3565 ( .A(n1127), .B(n1146), .Z(n4291) );
  CEOX2 U3566 ( .A(n3786), .B(n3668), .Z(n1459) );
  CND2IXL U3567 ( .B(a[12]), .A(n4466), .Z(n4469) );
  CIVX1 U3568 ( .A(n414), .Z(n412) );
  CEO3X2 U3569 ( .A(n917), .B(n915), .C(n930), .Z(n911) );
  CND2X2 U3570 ( .A(n917), .B(n915), .Z(n3496) );
  CND2X1 U3571 ( .A(n917), .B(n930), .Z(n3497) );
  CND2X2 U3572 ( .A(n915), .B(n930), .Z(n3498) );
  CND3X4 U3573 ( .A(n3496), .B(n3497), .C(n3498), .Z(n910) );
  CEOX2 U3574 ( .A(n912), .B(n899), .Z(n3499) );
  CEOX2 U3575 ( .A(n3499), .B(n910), .Z(n895) );
  CND2XL U3576 ( .A(n912), .B(n899), .Z(n3500) );
  CND2X1 U3577 ( .A(n912), .B(n910), .Z(n3501) );
  CND2X1 U3578 ( .A(n899), .B(n910), .Z(n3502) );
  CND3X2 U3579 ( .A(n3500), .B(n3501), .C(n3502), .Z(n894) );
  CIVX1 U3580 ( .A(n1135), .Z(n4005) );
  CND2X2 U3581 ( .A(n4040), .B(n4039), .Z(n24) );
  CIVXL U3582 ( .A(n399), .Z(n3503) );
  CEO3X1 U3583 ( .A(n992), .B(n2026), .C(n1995), .Z(n973) );
  CND2XL U3584 ( .A(n1995), .B(n992), .Z(n3504) );
  CND2X1 U3585 ( .A(n1995), .B(n2026), .Z(n3505) );
  CND2X1 U3586 ( .A(n992), .B(n2026), .Z(n3506) );
  CND3X1 U3587 ( .A(n3504), .B(n3505), .C(n3506), .Z(n972) );
  CEOX2 U3588 ( .A(n927), .B(n940), .Z(n3507) );
  CEOX2 U3589 ( .A(n3507), .B(n925), .Z(n923) );
  CND2XL U3590 ( .A(n925), .B(n940), .Z(n3508) );
  CND2X1 U3591 ( .A(n925), .B(n927), .Z(n3509) );
  CND2XL U3592 ( .A(n940), .B(n927), .Z(n3510) );
  CND3X1 U3593 ( .A(n3508), .B(n3509), .C(n3510), .Z(n922) );
  COND1X1 U3594 ( .A(n410), .B(n402), .C(n403), .Z(n397) );
  CND3X2 U3595 ( .A(n3607), .B(n3608), .C(n3609), .Z(n940) );
  CIVX8 U3596 ( .A(n4499), .Z(n4504) );
  COND1XL U3597 ( .A(n668), .B(n651), .C(n652), .Z(n3512) );
  CND2X1 U3598 ( .A(n1994), .B(n1784), .Z(n3575) );
  CIVXL U3599 ( .A(n307), .Z(n305) );
  CND2XL U3600 ( .A(n1486), .B(n1488), .Z(n3699) );
  CEOX1 U3601 ( .A(n3513), .B(n3101), .Z(n1327) );
  CND2XL U3602 ( .A(n1861), .B(n1830), .Z(n3514) );
  CND2XL U3603 ( .A(n1861), .B(n1885), .Z(n3515) );
  CND2XL U3604 ( .A(n1830), .B(n1885), .Z(n3516) );
  CND3X1 U3605 ( .A(n3514), .B(n3515), .C(n3516), .Z(n1326) );
  CNR2X1 U3606 ( .A(n1215), .B(n1244), .Z(n540) );
  COND2XL U3607 ( .A(n4184), .B(n2607), .C(n4506), .D(n2606), .Z(n2082) );
  CND2XL U3608 ( .A(n3239), .B(n3977), .Z(n3521) );
  CND2X1 U3609 ( .A(n3519), .B(n3520), .Z(n3522) );
  CIVXL U3610 ( .A(n1223), .Z(n3520) );
  CANR1X1 U3611 ( .A(n397), .B(n363), .C(n364), .Z(n362) );
  CEOX2 U3612 ( .A(n1428), .B(n1430), .Z(n3523) );
  CEOX2 U3613 ( .A(n3523), .B(n1432), .Z(n1399) );
  CND2X1 U3614 ( .A(n1432), .B(n1428), .Z(n3525) );
  CND2X1 U3615 ( .A(n1430), .B(n1428), .Z(n3526) );
  CENX1 U3616 ( .A(n1208), .B(n1183), .Z(n3527) );
  CND2IX1 U3617 ( .B(n3099), .A(n4589), .Z(n4400) );
  COND2X1 U3618 ( .A(n135), .B(n4601), .C(n2317), .D(net16439), .Z(n1725) );
  CIVX3 U3619 ( .A(n4583), .Z(n4374) );
  CENX1 U3620 ( .A(n1443), .B(n4151), .Z(n3787) );
  CND2IX1 U3621 ( .B(a[4]), .A(net19006), .Z(n3961) );
  CND2X2 U3622 ( .A(n4398), .B(n4440), .Z(n4441) );
  CND2X1 U3623 ( .A(n1421), .B(n1423), .Z(n3625) );
  COND2X1 U3624 ( .A(n3302), .B(n2413), .C(n2412), .D(net16426), .Z(n1890) );
  CND3X1 U3625 ( .A(n4415), .B(n4414), .C(n4416), .Z(n3528) );
  CND3X1 U3626 ( .A(n4414), .B(n4415), .C(n4416), .Z(n1158) );
  CEOX2 U3627 ( .A(n1241), .B(n1237), .Z(n3529) );
  CEOX2 U3628 ( .A(n3529), .B(n3352), .Z(n1225) );
  CND2X1 U3629 ( .A(n1260), .B(n1237), .Z(n3530) );
  CND2X1 U3630 ( .A(n1260), .B(n1241), .Z(n3531) );
  CND2X1 U3631 ( .A(n1237), .B(n1241), .Z(n3532) );
  CND3X2 U3632 ( .A(n3530), .B(n3531), .C(n3532), .Z(n1224) );
  CIVX2 U3633 ( .A(n3777), .Z(net17279) );
  CENX1 U3634 ( .A(a[22]), .B(net15916), .Z(n2816) );
  CND2X1 U3635 ( .A(n3772), .B(n1527), .Z(n3536) );
  CND2X2 U3636 ( .A(n3534), .B(n3535), .Z(n3537) );
  CND2X2 U3637 ( .A(n3536), .B(n3537), .Z(n1525) );
  CIVX1 U3638 ( .A(n1527), .Z(n3535) );
  CENX1 U3639 ( .A(net15974), .B(n4560), .Z(n2656) );
  CND2XL U3640 ( .A(n1363), .B(n1365), .Z(n3538) );
  CND2XL U3641 ( .A(n1363), .B(n1388), .Z(n3539) );
  CND2XL U3642 ( .A(n1365), .B(n1388), .Z(n3540) );
  CND3X1 U3643 ( .A(n3538), .B(n3539), .C(n3540), .Z(n1360) );
  CEOX2 U3644 ( .A(n1392), .B(n1367), .Z(n3541) );
  CEOX2 U3645 ( .A(n3541), .B(n3204), .Z(n1363) );
  CND2X1 U3646 ( .A(n1390), .B(n1367), .Z(n3542) );
  CND2X1 U3647 ( .A(n1390), .B(n1392), .Z(n3543) );
  CND3X2 U3648 ( .A(n3542), .B(n3543), .C(n3544), .Z(n1362) );
  CND2X1 U3649 ( .A(n1335), .B(n1362), .Z(n4170) );
  CEOX2 U3650 ( .A(n2067), .B(n2098), .Z(n3545) );
  CEOX1 U3651 ( .A(n3545), .B(n1302), .Z(n1263) );
  CND2XL U3652 ( .A(n1302), .B(n2098), .Z(n3546) );
  CND2XL U3653 ( .A(n2098), .B(n2067), .Z(n3548) );
  CND3X1 U3654 ( .A(n3546), .B(n3547), .C(n3548), .Z(n1262) );
  CIVX4 U3655 ( .A(net18261), .Z(net16490) );
  CEO3X2 U3656 ( .A(n2061), .B(n1128), .C(n1939), .Z(n1097) );
  CND2XL U3657 ( .A(n2061), .B(n1128), .Z(n3549) );
  CND2XL U3658 ( .A(n2061), .B(n1939), .Z(n3550) );
  CND2XL U3659 ( .A(n1128), .B(n1939), .Z(n3551) );
  CND3X2 U3660 ( .A(n3549), .B(n3550), .C(n3551), .Z(n1096) );
  CND2XL U3661 ( .A(n1075), .B(n1073), .Z(n3552) );
  CND2XL U3662 ( .A(n1075), .B(n1096), .Z(n3553) );
  CND2XL U3663 ( .A(n1073), .B(n1096), .Z(n3554) );
  CND3X1 U3664 ( .A(n3552), .B(n3553), .C(n3554), .Z(n1066) );
  CIVXL U3665 ( .A(n514), .Z(n3555) );
  CIVXL U3666 ( .A(n3555), .Z(n3556) );
  CND2XL U3667 ( .A(n1017), .B(n1038), .Z(n3557) );
  CND2XL U3668 ( .A(n1017), .B(n1019), .Z(n3558) );
  CND2XL U3669 ( .A(n1038), .B(n1019), .Z(n3559) );
  CND3XL U3670 ( .A(n3557), .B(n3558), .C(n3559), .Z(n1014) );
  CND2X1 U3671 ( .A(n1021), .B(n4036), .Z(n3562) );
  CND2X2 U3672 ( .A(n3560), .B(n3561), .Z(n3563) );
  CND2X2 U3673 ( .A(n3562), .B(n3563), .Z(n1017) );
  CIVXL U3674 ( .A(n1021), .Z(n3560) );
  CIVX2 U3675 ( .A(n4036), .Z(n3561) );
  CEO3X1 U3676 ( .A(n1048), .B(n1027), .C(n1046), .Z(n1021) );
  CENX1 U3677 ( .A(n1042), .B(n1040), .Z(n4036) );
  CNIVX2 U3678 ( .A(n3517), .Z(n3708) );
  CENX1 U3679 ( .A(n4582), .B(n4553), .Z(n2531) );
  CEOX2 U3680 ( .A(n1168), .B(n3904), .Z(net17986) );
  CND2XL U3681 ( .A(n1355), .B(n1382), .Z(n3564) );
  CND2XL U3682 ( .A(n1355), .B(n3366), .Z(n3565) );
  CND2XL U3683 ( .A(n1382), .B(n3366), .Z(n3566) );
  CND3X1 U3684 ( .A(n3564), .B(n3565), .C(n3566), .Z(n1344) );
  CEO3X2 U3685 ( .A(n1346), .B(n1321), .C(n1344), .Z(n1313) );
  CENX1 U3686 ( .A(n4579), .B(n4551), .Z(n2599) );
  CENX2 U3687 ( .A(n1147), .B(n1145), .Z(n3895) );
  CND2X2 U3688 ( .A(n4017), .B(n4018), .Z(product[56]) );
  CEO3XL U3689 ( .A(n883), .B(n881), .C(n894), .Z(n3567) );
  CEOX2 U3690 ( .A(n1474), .B(n1476), .Z(n3568) );
  CEOX2 U3691 ( .A(n3568), .B(n3436), .Z(n1447) );
  CND2X1 U3692 ( .A(n1453), .B(n1476), .Z(n3569) );
  CND2X1 U3693 ( .A(n1453), .B(n1474), .Z(n3570) );
  CND2X1 U3694 ( .A(n1476), .B(n1474), .Z(n3571) );
  CND3X2 U3695 ( .A(n3569), .B(n3570), .C(n3571), .Z(n1446) );
  CND3X2 U3696 ( .A(n4117), .B(n4118), .C(n4119), .Z(n1476) );
  CENXL U3697 ( .A(n4597), .B(net16104), .Z(n2321) );
  CENXL U3698 ( .A(n4597), .B(net16102), .Z(n2320) );
  CENXL U3699 ( .A(n4597), .B(n4559), .Z(n2327) );
  CENXL U3700 ( .A(n4597), .B(n4557), .Z(n2329) );
  CEOX1 U3701 ( .A(n1784), .B(n1753), .Z(n3573) );
  CEOX1 U3702 ( .A(n3573), .B(n1994), .Z(n953) );
  CND2XL U3703 ( .A(n1753), .B(n1784), .Z(n3576) );
  CND3X1 U3704 ( .A(n3574), .B(n3575), .C(n3576), .Z(n952) );
  COR2X1 U3705 ( .A(net17279), .B(n2517), .Z(n3577) );
  COR2XL U3706 ( .A(n3121), .B(n2516), .Z(n3578) );
  CND2X2 U3707 ( .A(n3577), .B(n3578), .Z(n1994) );
  CND2X1 U3708 ( .A(n1419), .B(n1440), .Z(n4081) );
  CENX1 U3709 ( .A(n4576), .B(n4555), .Z(n2628) );
  CND2X4 U3710 ( .A(n4371), .B(n4372), .Z(n3579) );
  CND2X2 U3711 ( .A(n3582), .B(n3583), .Z(n3886) );
  COND1X2 U3712 ( .A(net16472), .B(n220), .C(n221), .Z(n219) );
  COND2X1 U3713 ( .A(n63), .B(n2554), .C(n2553), .D(n4505), .Z(n3584) );
  COND2XL U3714 ( .A(n63), .B(n2554), .C(n2553), .D(n4505), .Z(n1080) );
  CIVXL U3715 ( .A(n992), .Z(n993) );
  CENX2 U3716 ( .A(n1229), .B(n1227), .Z(n3949) );
  CEO3X2 U3717 ( .A(n1239), .B(n1235), .C(n1233), .Z(n1227) );
  CENX2 U3718 ( .A(n3585), .B(n3894), .Z(n1189) );
  CENX1 U3719 ( .A(n4582), .B(n4551), .Z(n2533) );
  CEO3X2 U3720 ( .A(n1637), .B(n1633), .C(n1644), .Z(n1629) );
  CEOX2 U3721 ( .A(n1631), .B(n1642), .Z(n3586) );
  CEOX1 U3722 ( .A(n3586), .B(n1629), .Z(n1627) );
  CND2X1 U3723 ( .A(n1637), .B(n1633), .Z(n3587) );
  CND2X1 U3724 ( .A(n1637), .B(n1644), .Z(n3588) );
  CND2X1 U3725 ( .A(n1633), .B(n1644), .Z(n3589) );
  CND3X2 U3726 ( .A(n3587), .B(n3588), .C(n3589), .Z(n1628) );
  CND2XL U3727 ( .A(n1631), .B(n1642), .Z(n3590) );
  CND2X1 U3728 ( .A(n1631), .B(n1629), .Z(n3591) );
  CND2X1 U3729 ( .A(n1642), .B(n1629), .Z(n3592) );
  CND3X2 U3730 ( .A(n3590), .B(n3591), .C(n3592), .Z(n1626) );
  CEOX2 U3731 ( .A(n2176), .B(n1732), .Z(n1639) );
  CIVX2 U3732 ( .A(n3593), .Z(n1638) );
  CND2X1 U3733 ( .A(n2176), .B(n1732), .Z(n3593) );
  CND2IX2 U3734 ( .B(n4325), .A(n3767), .Z(n1732) );
  CND2X1 U3735 ( .A(n1638), .B(n1634), .Z(n4365) );
  CENX1 U3736 ( .A(n1375), .B(n3594), .Z(n1367) );
  CEO3X2 U3737 ( .A(n1242), .B(n2096), .C(n2188), .Z(n1213) );
  CNR2XL U3738 ( .A(n491), .B(n484), .Z(n3595) );
  CND2X1 U3739 ( .A(n3881), .B(n1126), .Z(n3598) );
  CND2X2 U3740 ( .A(n3598), .B(n3599), .Z(n1095) );
  CIVX2 U3741 ( .A(n3881), .Z(n3596) );
  CIVXL U3742 ( .A(n1126), .Z(n3597) );
  CNR2XL U3743 ( .A(n484), .B(n3330), .Z(n482) );
  COND2XL U3744 ( .A(n63), .B(n2577), .C(n4505), .D(n2576), .Z(n2052) );
  CND2X2 U3745 ( .A(n3078), .B(a[22]), .Z(n3835) );
  CIVX1 U3746 ( .A(n3719), .Z(n3833) );
  CENX2 U3747 ( .A(n1191), .B(n1216), .Z(n4476) );
  CNR2X2 U3748 ( .A(n2548), .B(n3121), .Z(n4325) );
  CENX1 U3749 ( .A(n4579), .B(net16104), .Z(n2585) );
  CEO3X2 U3750 ( .A(n1457), .B(n1455), .C(n1451), .Z(n1445) );
  CND2XL U3751 ( .A(n1457), .B(n1451), .Z(n3600) );
  CND2XL U3752 ( .A(n1457), .B(n1455), .Z(n3601) );
  CND2X1 U3753 ( .A(n1451), .B(n1455), .Z(n3602) );
  CND3XL U3754 ( .A(n3600), .B(n3601), .C(n3602), .Z(n1444) );
  CEO3X1 U3755 ( .A(n2227), .B(n1983), .C(n2166), .Z(n1457) );
  CIVX8 U3756 ( .A(n3765), .Z(net16541) );
  CND2X2 U3757 ( .A(n1195), .B(n1197), .Z(n4131) );
  CENX1 U3758 ( .A(n4572), .B(n4560), .Z(n2722) );
  CND2X2 U3759 ( .A(n3753), .B(n4370), .Z(n4371) );
  CND2XL U3760 ( .A(n414), .B(n396), .Z(n394) );
  CND2XL U3761 ( .A(n414), .B(n748), .Z(n405) );
  CIVXL U3762 ( .A(n4312), .Z(n3603) );
  CND2X2 U3763 ( .A(n4113), .B(n3605), .Z(n3880) );
  CND2X1 U3764 ( .A(n1305), .B(n1332), .Z(n559) );
  COAN1X1 U3765 ( .A(n651), .B(n668), .C(n652), .Z(n3606) );
  COND1XL U3766 ( .A(n633), .B(n4226), .C(n634), .Z(n3990) );
  CND3X1 U3767 ( .A(n4367), .B(n4368), .C(n4369), .Z(n1624) );
  COND2X2 U3768 ( .A(n27), .B(n2686), .C(net16451), .D(n2685), .Z(n2160) );
  CND2X1 U3769 ( .A(n960), .B(n945), .Z(n3607) );
  CND2XL U3770 ( .A(n960), .B(n962), .Z(n3608) );
  CND2XL U3771 ( .A(n945), .B(n962), .Z(n3609) );
  COND2X2 U3772 ( .A(n4063), .B(n2623), .C(net18914), .D(n2622), .Z(n2098) );
  CNR2XL U3773 ( .A(n4351), .B(n616), .Z(n3610) );
  CIVX1 U3774 ( .A(n3611), .Z(n3612) );
  COND2XL U3775 ( .A(n63), .B(n2574), .C(n2573), .D(n4505), .Z(n3613) );
  COND2XL U3776 ( .A(n4316), .B(n2574), .C(n2573), .D(n4505), .Z(n2049) );
  CANR1X1 U3777 ( .A(n779), .B(n4465), .C(n664), .Z(n662) );
  CEOX1 U3778 ( .A(n662), .B(n196), .Z(product[16]) );
  CEO3X1 U3779 ( .A(n1589), .B(n1600), .C(n1587), .Z(n1583) );
  CEOX2 U3780 ( .A(n1585), .B(n1598), .Z(n3614) );
  CEOX1 U3781 ( .A(n3614), .B(n1583), .Z(n1581) );
  CND2XL U3782 ( .A(n1589), .B(n1600), .Z(n3615) );
  CND2XL U3783 ( .A(n1589), .B(n1587), .Z(n3616) );
  CND2XL U3784 ( .A(n1600), .B(n1587), .Z(n3617) );
  CND3X1 U3785 ( .A(n3615), .B(n3616), .C(n3617), .Z(n1582) );
  CND2XL U3786 ( .A(n1585), .B(n1598), .Z(n3618) );
  CND2XL U3787 ( .A(n1585), .B(n1583), .Z(n3619) );
  CND2XL U3788 ( .A(n1583), .B(n1598), .Z(n3620) );
  CND3X1 U3789 ( .A(n3619), .B(n3618), .C(n3620), .Z(n1580) );
  CEOX2 U3790 ( .A(n1957), .B(n2048), .Z(n4305) );
  CND2X1 U3791 ( .A(n2048), .B(n1957), .Z(n4308) );
  CND2X1 U3792 ( .A(n4309), .B(n2048), .Z(n4306) );
  CEOX2 U3793 ( .A(n4305), .B(n4309), .Z(n1559) );
  CEOX2 U3794 ( .A(n1498), .B(n1496), .Z(n4346) );
  CND2IX2 U3795 ( .B(n4198), .A(net18211), .Z(n4199) );
  CAN2XL U3796 ( .A(n552), .B(n3822), .Z(net17211) );
  CIVX1 U3797 ( .A(n534), .Z(n532) );
  CIVX1 U3798 ( .A(n2144), .Z(n4502) );
  CIVX8 U3799 ( .A(n129), .Z(n4601) );
  CND2X1 U3800 ( .A(n2816), .B(n3084), .Z(net17728) );
  CND2XL U3801 ( .A(n1216), .B(n1191), .Z(n4523) );
  CND3XL U3802 ( .A(n4537), .B(n4538), .C(n4539), .Z(n1280) );
  CEOX1 U3803 ( .A(net18211), .B(n4551), .Z(n2401) );
  CEO3XL U3804 ( .A(n2024), .B(n2146), .C(n2206), .Z(n1637) );
  CIVX2 U3805 ( .A(n3621), .Z(n3622) );
  CNIVX4 U3806 ( .A(n57), .Z(n4121) );
  CEO3X1 U3807 ( .A(n1444), .B(n1421), .C(n1423), .Z(n1417) );
  CND2XL U3808 ( .A(n1444), .B(n1421), .Z(n3623) );
  CND2X1 U3809 ( .A(n1444), .B(n1423), .Z(n3624) );
  CND3X2 U3810 ( .A(n3623), .B(n3624), .C(n3625), .Z(n1416) );
  CEOX2 U3811 ( .A(n1416), .B(n3626), .Z(n1389) );
  CND2XL U3812 ( .A(n1395), .B(n1393), .Z(n3627) );
  CND2X1 U3813 ( .A(n1395), .B(n1416), .Z(n3628) );
  CND2X1 U3814 ( .A(n1393), .B(n1416), .Z(n3629) );
  CND3X2 U3815 ( .A(n3627), .B(n3628), .C(n3629), .Z(n1388) );
  CEO3X1 U3816 ( .A(n2044), .B(n1922), .C(n1953), .Z(n1479) );
  CND2XL U3817 ( .A(n1922), .B(n1953), .Z(n3630) );
  CND2XL U3818 ( .A(n1922), .B(n2044), .Z(n3631) );
  CND2X1 U3819 ( .A(n1953), .B(n2044), .Z(n3632) );
  CND2X1 U3820 ( .A(n3098), .B(n1471), .Z(n3634) );
  CND3X2 U3821 ( .A(n3634), .B(n3635), .C(n3636), .Z(n1464) );
  CEO3X2 U3822 ( .A(n1479), .B(n1475), .C(n1477), .Z(n1469) );
  CEO3X1 U3823 ( .A(n1271), .B(n1265), .C(n1267), .Z(n1257) );
  CND2XL U3824 ( .A(n1271), .B(n1267), .Z(n3637) );
  CND2X1 U3825 ( .A(n1271), .B(n1265), .Z(n3638) );
  CND2X1 U3826 ( .A(n1267), .B(n1265), .Z(n3639) );
  CND3X2 U3827 ( .A(n3637), .B(n3638), .C(n3639), .Z(n1256) );
  CEOX2 U3828 ( .A(n4219), .B(n4224), .Z(n1433) );
  CIVDX2 U3829 ( .A(a[14]), .Z0(n3986), .Z1(n3985) );
  CEOX2 U3830 ( .A(n2238), .B(n3780), .Z(n3640) );
  CND2X1 U3831 ( .A(n1662), .B(n3780), .Z(n3641) );
  CND2X1 U3832 ( .A(n1662), .B(n2238), .Z(n3642) );
  CND2XL U3833 ( .A(n3780), .B(n2238), .Z(n3643) );
  CND3X2 U3834 ( .A(n3641), .B(n3642), .C(n3643), .Z(n1646) );
  CIVX4 U3835 ( .A(net18261), .Z(n3644) );
  COND2X1 U3836 ( .A(n3302), .B(n2414), .C(n2413), .D(net16426), .Z(n1891) );
  CIVXL U3837 ( .A(n4251), .Z(n3645) );
  CIVXL U3838 ( .A(n4583), .Z(n3646) );
  CENX2 U3839 ( .A(n3647), .B(n1541), .Z(n1531) );
  CENX2 U3840 ( .A(n1539), .B(n1537), .Z(n3647) );
  CND2X2 U3841 ( .A(n3648), .B(a[6]), .Z(n3914) );
  COND2X1 U3842 ( .A(net18896), .B(n2667), .C(n3644), .D(n2666), .Z(n2142) );
  CFA1XL U3843 ( .A(n2184), .B(n2245), .CI(n2154), .CO(n1708), .S(n1709) );
  CIVXL U3844 ( .A(n21), .Z(n3648) );
  CND2XL U3845 ( .A(net16541), .B(n4563), .Z(n3651) );
  CND2X1 U3846 ( .A(n3649), .B(n3650), .Z(n3652) );
  CIVXL U3847 ( .A(n4563), .Z(n3650) );
  CEOX2 U3848 ( .A(n1002), .B(n985), .Z(n3653) );
  CND2X1 U3849 ( .A(n983), .B(n985), .Z(n3654) );
  CND2X1 U3850 ( .A(n983), .B(n1002), .Z(n3655) );
  CND2X1 U3851 ( .A(n985), .B(n1002), .Z(n3656) );
  CND3X2 U3852 ( .A(n3654), .B(n3655), .C(n3656), .Z(n978) );
  CIVX2 U3853 ( .A(n1189), .Z(n4213) );
  CENX1 U3854 ( .A(n3908), .B(n4562), .Z(n2654) );
  CIVX2 U3855 ( .A(n12), .Z(n3659) );
  CIVX2 U3856 ( .A(n12), .Z(n4574) );
  COND2X1 U3857 ( .A(n4316), .B(n2561), .C(n2560), .D(n4505), .Z(n2036) );
  CEO3X2 U3858 ( .A(n1998), .B(n1757), .C(n3666), .Z(n1031) );
  CND2XL U3859 ( .A(n1998), .B(n1757), .Z(n3660) );
  CND2XL U3860 ( .A(n1998), .B(n2058), .Z(n3661) );
  CND2XL U3861 ( .A(n1757), .B(n2058), .Z(n3662) );
  CND3X1 U3862 ( .A(n3660), .B(n3661), .C(n3662), .Z(n1030) );
  CND2XL U3863 ( .A(n1033), .B(n1029), .Z(n3663) );
  CND2XL U3864 ( .A(n1033), .B(n1031), .Z(n3664) );
  CND2XL U3865 ( .A(n1029), .B(n1031), .Z(n3665) );
  CND3X1 U3866 ( .A(n3663), .B(n3664), .C(n3665), .Z(n1022) );
  COAN1X1 U3867 ( .A(n458), .B(n448), .C(n449), .Z(n445) );
  CNIVX1 U3868 ( .A(n2058), .Z(n3666) );
  COND2XL U3869 ( .A(n54), .B(n2583), .C(n4506), .D(n2582), .Z(n2058) );
  COND2X1 U3870 ( .A(n117), .B(n4281), .C(n2383), .D(net16433), .Z(n3668) );
  COAN1X1 U3871 ( .A(n369), .B(n379), .C(n370), .Z(n366) );
  CEO3X2 U3872 ( .A(n1950), .B(n2072), .C(n1981), .Z(n1403) );
  CND2XL U3873 ( .A(n1950), .B(n1981), .Z(n3670) );
  CND2XL U3874 ( .A(n1950), .B(n2072), .Z(n3671) );
  CND2X1 U3875 ( .A(n1981), .B(n2072), .Z(n3672) );
  CND3X1 U3876 ( .A(n3671), .B(n3670), .C(n3672), .Z(n1402) );
  CND2X1 U3877 ( .A(n1403), .B(n3674), .Z(n3675) );
  CND2X1 U3878 ( .A(n3673), .B(n1426), .Z(n3676) );
  CND2X2 U3879 ( .A(n3675), .B(n3676), .Z(n4404) );
  CIVXL U3880 ( .A(n1403), .Z(n3673) );
  CIVXL U3881 ( .A(n1426), .Z(n3674) );
  CENX1 U3882 ( .A(n1404), .B(n1402), .Z(n3978) );
  CND2X4 U3883 ( .A(n3754), .B(n3783), .Z(n4372) );
  CEOX2 U3884 ( .A(n1487), .B(n1506), .Z(n3792) );
  CIVX2 U3885 ( .A(n3), .Z(n3677) );
  CIVX2 U3886 ( .A(n3), .Z(n3678) );
  CIVX2 U3887 ( .A(n3), .Z(n4421) );
  CND2X1 U3888 ( .A(n3733), .B(n1247), .Z(n3681) );
  CND2X2 U3889 ( .A(n3681), .B(n3682), .Z(n1245) );
  CIVX2 U3890 ( .A(n3733), .Z(n3679) );
  CND2X4 U3891 ( .A(n2818), .B(net16510), .Z(n90) );
  CANR1X1 U3892 ( .A(n753), .B(n474), .C(n467), .Z(n3683) );
  CANR1XL U3893 ( .A(n753), .B(n474), .C(n467), .Z(n3684) );
  CANR1X1 U3894 ( .A(n753), .B(n474), .C(n467), .Z(n461) );
  CND2XL U3895 ( .A(n4309), .B(n1957), .Z(n4307) );
  CND3X1 U3896 ( .A(n3710), .B(n3711), .C(n3712), .Z(n1106) );
  CND3X2 U3897 ( .A(n4235), .B(n4236), .C(n4237), .Z(n1506) );
  CND2X1 U3898 ( .A(n1528), .B(n1511), .Z(n4235) );
  CNR2IX1 U3899 ( .B(n3244), .A(n3771), .Z(n1926) );
  CENX2 U3900 ( .A(n1116), .B(n3685), .Z(n1089) );
  CENX2 U3901 ( .A(n1097), .B(n1095), .Z(n3685) );
  CANR1X2 U3902 ( .A(n4480), .B(n659), .C(n654), .Z(n652) );
  CIVXL U3903 ( .A(n3254), .Z(n462) );
  CEO3X1 U3904 ( .A(n1009), .B(n1007), .C(n1013), .Z(n1003) );
  CND2XL U3905 ( .A(n1009), .B(n1013), .Z(n3686) );
  CND2X1 U3906 ( .A(n1013), .B(n1007), .Z(n3688) );
  CEO3X1 U3907 ( .A(n1875), .B(n1787), .C(n1849), .Z(n1009) );
  CND2XL U3908 ( .A(n1875), .B(n1849), .Z(n3689) );
  CND2XL U3909 ( .A(n1875), .B(n1787), .Z(n3690) );
  CND2X1 U3910 ( .A(n1849), .B(n1787), .Z(n3691) );
  CND3XL U3911 ( .A(n3689), .B(n3690), .C(n3691), .Z(n1008) );
  CIVXL U3912 ( .A(n308), .Z(n306) );
  CNR2IX1 U3913 ( .B(n3244), .A(net16512), .Z(n1959) );
  CIVX4 U3914 ( .A(net16420), .Z(net18913) );
  CIVXL U3915 ( .A(n533), .Z(n3695) );
  COND2XL U3916 ( .A(net18628), .B(n2377), .C(net16433), .D(n2376), .Z(n1861)
         );
  CEOX1 U3917 ( .A(n979), .B(n996), .Z(n4165) );
  CND2XL U3918 ( .A(n977), .B(n979), .Z(n4167) );
  CIVX4 U3919 ( .A(n3993), .Z(n3893) );
  CENX1 U3920 ( .A(net15912), .B(n4541), .Z(n2412) );
  CND2X1 U3921 ( .A(n1162), .B(n1139), .Z(n3934) );
  CNIVX4 U3922 ( .A(n3703), .Z(net17297) );
  CENXL U3923 ( .A(n4572), .B(n4565), .Z(n2714) );
  CAOR1X1 U3924 ( .A(n4505), .B(n63), .C(n2549), .Z(n2026) );
  CENX2 U3925 ( .A(n3488), .B(n3696), .Z(n1161) );
  CENX1 U3926 ( .A(n1192), .B(n1165), .Z(n3696) );
  CIVX1 U3927 ( .A(n223), .Z(n221) );
  COND2X1 U3928 ( .A(n4461), .B(n2740), .C(n2739), .D(n4510), .Z(n2213) );
  CENX1 U3929 ( .A(net15974), .B(n4561), .Z(n2655) );
  CND2X1 U3930 ( .A(n1236), .B(n1240), .Z(n3922) );
  CND2XL U3931 ( .A(n1467), .B(n1486), .Z(n3697) );
  CND3X1 U3932 ( .A(n3697), .B(n3699), .C(n3698), .Z(n1462) );
  CEO3XL U3933 ( .A(n2045), .B(n3145), .C(n2076), .Z(n1501) );
  CND2XL U3934 ( .A(n2045), .B(n2076), .Z(n3700) );
  CND3X1 U3935 ( .A(n3700), .B(n3701), .C(n3702), .Z(n1500) );
  COND2X1 U3936 ( .A(n54), .B(n2601), .C(n4507), .D(n2600), .Z(n2076) );
  COR2X2 U3937 ( .A(n4316), .B(n2557), .Z(n4319) );
  CND2X2 U3938 ( .A(n4040), .B(n4039), .Z(n3703) );
  CEOX2 U3939 ( .A(n3708), .B(n3704), .Z(n1217) );
  CND2X1 U3940 ( .A(n3371), .B(n1221), .Z(n3705) );
  CND2X1 U3941 ( .A(n3517), .B(n1250), .Z(n3706) );
  CND3X2 U3942 ( .A(n3705), .B(n3706), .C(n3707), .Z(n1216) );
  CND2XL U3943 ( .A(n3), .B(a[2]), .Z(n3709) );
  CND3X1 U3944 ( .A(n4248), .B(n4249), .C(n4250), .Z(n1250) );
  CIVX1 U3945 ( .A(n317), .Z(n3741) );
  COND2X2 U3946 ( .A(n4012), .B(n2399), .C(n2398), .D(net17425), .Z(n1877) );
  CND2X1 U3947 ( .A(n3256), .B(n1109), .Z(n3711) );
  CND2XL U3948 ( .A(n3256), .B(n1134), .Z(n3712) );
  CEO3XL U3949 ( .A(n1117), .B(n1140), .C(n1115), .Z(n1111) );
  CND3X2 U3950 ( .A(n3934), .B(n3935), .C(n3936), .Z(n1134) );
  CND2X2 U3951 ( .A(n549), .B(n561), .Z(n547) );
  CENX1 U3952 ( .A(n1114), .B(n3713), .Z(n1087) );
  CENX1 U3953 ( .A(n1093), .B(n1091), .Z(n3713) );
  CEOX1 U3954 ( .A(n3858), .B(n1560), .Z(n1535) );
  CND2XL U3955 ( .A(n2201), .B(n2171), .Z(n3857) );
  CND3X2 U3956 ( .A(n4031), .B(n4030), .C(n4032), .Z(n1218) );
  CEOX2 U3957 ( .A(n1973), .B(n1185), .Z(n3714) );
  CEOX1 U3958 ( .A(n3714), .B(n1212), .Z(n1175) );
  CND2XL U3959 ( .A(n1212), .B(n1185), .Z(n3715) );
  CND2X1 U3960 ( .A(n1212), .B(n1973), .Z(n3716) );
  CND2XL U3961 ( .A(n1185), .B(n1973), .Z(n3717) );
  CND3X2 U3962 ( .A(n3715), .B(n3716), .C(n3717), .Z(n1174) );
  CND3X1 U3963 ( .A(n3928), .B(n3929), .C(n3930), .Z(n1212) );
  CIVX1 U3964 ( .A(n1184), .Z(n1185) );
  CND2XL U3965 ( .A(n1256), .B(n1258), .Z(n4426) );
  COND2X2 U3966 ( .A(n2283), .B(n144), .C(n2282), .D(n3277), .Z(n1767) );
  CIVX2 U3967 ( .A(n93), .Z(n3718) );
  CIVX2 U3968 ( .A(n93), .Z(n3719) );
  CND2X1 U3969 ( .A(n1194), .B(n1167), .Z(n3720) );
  CND2XL U3970 ( .A(n1194), .B(n1169), .Z(n3721) );
  CND2X1 U3971 ( .A(n1167), .B(n1169), .Z(n3722) );
  CND3X2 U3972 ( .A(n3720), .B(n3721), .C(n3722), .Z(n1162) );
  CIVX2 U3973 ( .A(n93), .Z(n4594) );
  CEOX2 U3974 ( .A(n1162), .B(n4279), .Z(n1135) );
  CAOR1XL U3975 ( .A(net16451), .B(n27), .C(n2681), .Z(n3723) );
  CIVX2 U3976 ( .A(n1148), .Z(n3865) );
  CND3X2 U3977 ( .A(n4185), .B(n4187), .C(n4186), .Z(n1418) );
  CND2X1 U3978 ( .A(n1446), .B(n1448), .Z(n4186) );
  CND2XL U3979 ( .A(n3308), .B(n1233), .Z(n3724) );
  CND2XL U3980 ( .A(n3308), .B(n1235), .Z(n3725) );
  CND2X1 U3981 ( .A(n1233), .B(n1235), .Z(n3726) );
  CND3X1 U3982 ( .A(n3724), .B(n3725), .C(n3726), .Z(n1226) );
  CND2X1 U3983 ( .A(n1226), .B(n1199), .Z(n4114) );
  CND2X1 U3984 ( .A(n4578), .B(n3728), .Z(n3729) );
  CND2X2 U3985 ( .A(n3727), .B(a[10]), .Z(n3730) );
  CND2X2 U3986 ( .A(n3729), .B(n3730), .Z(n4095) );
  CIVX1 U3987 ( .A(n4578), .Z(n3727) );
  COND2XL U3988 ( .A(n4461), .B(n2737), .C(n2736), .D(n4510), .Z(n2210) );
  COND2XL U3989 ( .A(n4461), .B(n2741), .C(n2740), .D(n4510), .Z(n2214) );
  CANR1X1 U3990 ( .A(n686), .B(n4488), .C(n681), .Z(n679) );
  CENX1 U3991 ( .A(n3893), .B(n4540), .Z(n2612) );
  CND2X2 U3992 ( .A(n4075), .B(net18561), .Z(n4077) );
  CAOR1XL U3993 ( .A(n753), .B(n474), .C(n467), .Z(n3731) );
  CANR1X1 U3994 ( .A(n359), .B(n439), .C(n360), .Z(n3732) );
  CANR1X1 U3995 ( .A(n359), .B(n439), .C(n360), .Z(n354) );
  CIVXL U3996 ( .A(n511), .Z(n758) );
  CENX2 U3997 ( .A(n1249), .B(n1276), .Z(n3733) );
  COND2XL U3998 ( .A(n4012), .B(n2402), .C(n2401), .D(net17425), .Z(n1879) );
  CND2X1 U3999 ( .A(n4078), .B(n3735), .Z(n3736) );
  CND2X2 U4000 ( .A(n3734), .B(n3290), .Z(n3737) );
  CND2X2 U4001 ( .A(n3736), .B(n3737), .Z(n1413) );
  CIVX2 U4002 ( .A(n4078), .Z(n3734) );
  CIVXL U4003 ( .A(n1415), .Z(n3735) );
  CND2X2 U4004 ( .A(n1223), .B(n1225), .Z(n4031) );
  CND2X2 U4005 ( .A(n3658), .B(n3959), .Z(n4040) );
  CNIVX4 U4006 ( .A(n145), .Z(n4566) );
  CIVX1 U4007 ( .A(n4267), .Z(n4015) );
  CNIVX3 U4008 ( .A(n4566), .Z(n3748) );
  CIVX8 U4009 ( .A(n3925), .Z(net16420) );
  CND2X4 U4010 ( .A(n3926), .B(net18422), .Z(n3925) );
  CND2X1 U4011 ( .A(net18200), .B(n4201), .Z(n4238) );
  CEO3X2 U4012 ( .A(n1153), .B(n1151), .C(n1149), .Z(n1143) );
  CND2XL U4013 ( .A(n1153), .B(n1149), .Z(n3738) );
  CND2XL U4014 ( .A(n1153), .B(n1151), .Z(n3739) );
  CND2X1 U4015 ( .A(n1149), .B(n1151), .Z(n3740) );
  CEO3X1 U4016 ( .A(n1879), .B(n2063), .C(n2003), .Z(n1153) );
  COND1X1 U4017 ( .A(n573), .B(n567), .C(n568), .Z(n562) );
  CENX2 U4018 ( .A(n150), .B(n219), .Z(product[62]) );
  CND2X1 U4019 ( .A(n317), .B(n158), .Z(n3743) );
  CND2X2 U4020 ( .A(n3741), .B(n3742), .Z(n3744) );
  CND2X2 U4021 ( .A(n3743), .B(n3744), .Z(product[54]) );
  CIVX2 U4022 ( .A(n158), .Z(n3742) );
  CIVXL U4023 ( .A(n3037), .Z(n533) );
  CENXL U4024 ( .A(n3909), .B(n4565), .Z(n2648) );
  CIVX3 U4025 ( .A(net15980), .Z(n3909) );
  CNIVX2 U4026 ( .A(n2187), .Z(n3745) );
  CND2XL U4027 ( .A(n1207), .B(n1205), .Z(n4110) );
  CIVX3 U4028 ( .A(n4182), .Z(n4582) );
  CND2X2 U4029 ( .A(n4041), .B(n1058), .Z(n472) );
  CIVX1 U4030 ( .A(a[6]), .Z(net17482) );
  CIVX2 U4031 ( .A(net15980), .Z(n3908) );
  CNR2IX4 U4032 ( .B(n2820), .A(n3380), .Z(n3777) );
  CIVX1 U4033 ( .A(n582), .Z(n767) );
  CND2X2 U4034 ( .A(n4417), .B(n4418), .Z(n4420) );
  CIVX1 U4035 ( .A(n3746), .Z(n4417) );
  CENX1 U4036 ( .A(n3790), .B(n4552), .Z(n2565) );
  COND1X1 U4037 ( .A(n678), .B(n690), .C(n679), .Z(n677) );
  CND2X1 U4038 ( .A(n3909), .B(net16102), .Z(n3938) );
  CIVX2 U4039 ( .A(net15980), .Z(net15974) );
  CND2X2 U4040 ( .A(n4419), .B(n4420), .Z(n2283) );
  CIVX1 U4041 ( .A(n75), .Z(n3950) );
  CIVX3 U4042 ( .A(n75), .Z(n4586) );
  CND2X1 U4043 ( .A(n3747), .B(n4603), .Z(n4419) );
  CENX1 U4044 ( .A(n4582), .B(n4552), .Z(n2532) );
  CND2IX1 U4045 ( .B(n3244), .A(n3790), .Z(n2581) );
  CND2IX1 U4046 ( .B(n3244), .A(n4595), .Z(n2383) );
  COND2X1 U4047 ( .A(net18772), .B(net18827), .C(n2713), .D(net16451), .Z(
        n1737) );
  CNIVX4 U4048 ( .A(n2804), .Z(n4544) );
  CNIVX4 U4049 ( .A(n2787), .Z(n4561) );
  COND2X1 U4050 ( .A(n9), .B(n2758), .C(n6), .D(n2757), .Z(n2231) );
  CND2X1 U4051 ( .A(n4330), .B(n4331), .Z(n2738) );
  CIVX3 U4052 ( .A(n4519), .Z(n4520) );
  CND2X1 U4053 ( .A(n1027), .B(n1046), .Z(n4146) );
  CIVXL U4054 ( .A(net17728), .Z(n3902) );
  CENX1 U4055 ( .A(n4573), .B(n4559), .Z(n2723) );
  CENX1 U4056 ( .A(n4579), .B(n4562), .Z(n2588) );
  CENX1 U4057 ( .A(n4463), .B(n4544), .Z(n2309) );
  CENX1 U4058 ( .A(n4602), .B(n2809), .Z(n2281) );
  CND2X1 U4059 ( .A(n4332), .B(n4343), .Z(n4334) );
  CENX1 U4060 ( .A(n3893), .B(n4549), .Z(n2601) );
  CND2X1 U4061 ( .A(n3838), .B(n3839), .Z(n2393) );
  CND2X1 U4062 ( .A(n1449), .B(n1470), .Z(n4194) );
  CND2X2 U4063 ( .A(n3878), .B(n3879), .Z(n3903) );
  COND2X1 U4064 ( .A(n3301), .B(n2409), .C(n2408), .D(net16426), .Z(n1886) );
  CND3X1 U4065 ( .A(n4283), .B(n4284), .C(n4285), .Z(n1540) );
  CND3X2 U4066 ( .A(n4107), .B(n4108), .C(n4109), .Z(n1554) );
  CND2X1 U4067 ( .A(n1578), .B(n2141), .Z(n4107) );
  COR2XL U4068 ( .A(n3211), .B(n2760), .Z(n4264) );
  CNR2IX1 U4069 ( .B(n3244), .A(net16413), .Z(n1992) );
  CND2X1 U4070 ( .A(n320), .B(n4486), .Z(n309) );
  CIVX8 U4071 ( .A(n4509), .Z(n4510) );
  CND3X1 U4072 ( .A(n3181), .B(n4114), .C(n4115), .Z(n1192) );
  CENX1 U4073 ( .A(n3910), .B(n1204), .Z(n1173) );
  CND2X1 U4074 ( .A(n1281), .B(n1283), .Z(n4163) );
  CND2X1 U4075 ( .A(n1048), .B(n1046), .Z(n4145) );
  CND2X1 U4076 ( .A(n620), .B(n4475), .Z(n613) );
  CND2X1 U4077 ( .A(n845), .B(n854), .Z(n342) );
  CND2X1 U4078 ( .A(n233), .B(n4498), .Z(n224) );
  CND2X1 U4079 ( .A(n827), .B(n834), .Z(n316) );
  CND3X1 U4080 ( .A(n3845), .B(n3846), .C(n3847), .Z(n1686) );
  CFA1X1 U4081 ( .A(n1047), .B(n1045), .CI(n1066), .CO(n1040), .S(n1041) );
  CND2X1 U4082 ( .A(n3869), .B(n1386), .Z(n573) );
  CND2X1 U4083 ( .A(n799), .B(n802), .Z(n255) );
  CND2XL U4084 ( .A(n741), .B(n327), .Z(n159) );
  CENX1 U4085 ( .A(n205), .B(n3769), .Z(product[7]) );
  CNIVXL U4086 ( .A(n3028), .Z(n4321) );
  CAN2X1 U4087 ( .A(n3882), .B(n956), .Z(n3752) );
  CIVDX2 U4088 ( .A(n3892), .Z0(n3753), .Z1(n3754) );
  CIVX2 U4089 ( .A(n3464), .Z(n545) );
  CIVX1 U4090 ( .A(n3807), .Z(net18610) );
  COND2XL U4091 ( .A(net18896), .B(n2659), .C(net16490), .D(n2658), .Z(n2134)
         );
  CIVX2 U4092 ( .A(a[4]), .Z(n3959) );
  CIVDXL U4093 ( .A(n3331), .Z0(n3756), .Z1(n3757) );
  COR2X1 U4094 ( .A(n799), .B(n802), .Z(n3759) );
  CENX1 U4095 ( .A(n4580), .B(n4556), .Z(n2561) );
  CIVDX4 U4096 ( .A(n4586), .Z0(n3760), .Z1(n3761) );
  CIVX1 U4097 ( .A(n2809), .Z(n4343) );
  COAN1X1 U4098 ( .A(n693), .B(n697), .C(n694), .Z(n3762) );
  COAN1XL U4099 ( .A(n266), .B(n241), .C(n242), .Z(n3763) );
  COR2XL U4100 ( .A(n2251), .B(n1739), .Z(n3764) );
  CNIVX4 U4101 ( .A(net15988), .Z(n3765) );
  CIVXL U4102 ( .A(n21), .Z(n3766) );
  COND1X1 U4103 ( .A(n666), .B(n660), .C(n661), .Z(n659) );
  CIVXL U4104 ( .A(n660), .Z(n778) );
  CND2XL U4105 ( .A(net17154), .B(n3465), .Z(n3767) );
  CIVX2 U4106 ( .A(n4123), .Z(n629) );
  CNR2X1 U4107 ( .A(n693), .B(n696), .Z(n691) );
  CIVXL U4108 ( .A(n696), .Z(n785) );
  COND1XL U4109 ( .A(n696), .B(n698), .C(n697), .Z(n695) );
  CIVX1 U4110 ( .A(n720), .Z(n718) );
  CIVXL U4111 ( .A(n707), .Z(n3768) );
  CIVXL U4112 ( .A(n3768), .Z(n3769) );
  CIVXL U4113 ( .A(n2185), .Z(n4458) );
  CND2XL U4114 ( .A(n780), .B(n672), .Z(n198) );
  CIVXL U4115 ( .A(n671), .Z(n780) );
  CEOX2 U4116 ( .A(n195), .B(n657), .Z(product[17]) );
  CHA1XL U4117 ( .A(n1738), .B(n2218), .CO(n1722), .S(n1723) );
  CIVX1 U4118 ( .A(n3996), .Z(n676) );
  CENXL U4119 ( .A(n193), .B(n642), .Z(product[19]) );
  COND1XL U4120 ( .A(n3172), .B(n4282), .C(n603), .Z(n3770) );
  CENX2 U4121 ( .A(n3669), .B(n3785), .Z(n3771) );
  CENX1 U4122 ( .A(n3669), .B(n3785), .Z(net16416) );
  CND2X1 U4123 ( .A(n1409), .B(n1426), .Z(n4405) );
  CIVXL U4124 ( .A(n3770), .Z(n3773) );
  CNIVXL U4125 ( .A(n4589), .Z(n3774) );
  CENX1 U4126 ( .A(n3775), .B(n1236), .Z(n1203) );
  CENX1 U4127 ( .A(n3779), .B(n1335), .Z(n1333) );
  CNIVX2 U4128 ( .A(n2147), .Z(n3780) );
  CIVXL U4129 ( .A(n514), .Z(n516) );
  CND3X2 U4130 ( .A(n4128), .B(n4129), .C(n4130), .Z(n1220) );
  CENX1 U4131 ( .A(n3781), .B(n1353), .Z(n1343) );
  CENX1 U4132 ( .A(n1351), .B(n1357), .Z(n3781) );
  CIVX2 U4133 ( .A(n4584), .Z(n3782) );
  CIVX3 U4134 ( .A(n4584), .Z(n4583) );
  COND2X1 U4135 ( .A(n2598), .B(n54), .C(n4506), .D(n2597), .Z(n2073) );
  CND2XL U4136 ( .A(n2125), .B(n3723), .Z(n4072) );
  CIVX3 U4137 ( .A(n4370), .Z(n3783) );
  CFA1XL U4138 ( .A(n1870), .B(n1779), .CI(n1896), .CO(n874), .S(n875) );
  CEOX2 U4139 ( .A(n182), .B(n560), .Z(product[30]) );
  CIVX4 U4140 ( .A(a[20]), .Z(n3784) );
  CIVX8 U4141 ( .A(n3784), .Z(n3785) );
  COND2X1 U4142 ( .A(n3302), .B(n2413), .C(n2412), .D(net16426), .Z(n3786) );
  CENX2 U4143 ( .A(n4596), .B(a[24]), .Z(n2815) );
  CEOX2 U4144 ( .A(a[26]), .B(n4311), .Z(n4280) );
  CIVX8 U4145 ( .A(net17930), .Z(net17738) );
  CENXL U4146 ( .A(n1443), .B(n4151), .Z(n1439) );
  CENX2 U4147 ( .A(a[16]), .B(n4583), .Z(n3789) );
  CENX1 U4148 ( .A(n3026), .B(n4540), .Z(n2480) );
  CND2X1 U4149 ( .A(n1984), .B(n2228), .Z(n4118) );
  CAOR1XL U4150 ( .A(n123), .B(net17738), .C(n2318), .Z(n1802) );
  COND2XL U4151 ( .A(net17738), .B(n2319), .C(n123), .D(n2318), .Z(n1803) );
  COND2XL U4152 ( .A(net17738), .B(n2323), .C(n123), .D(n2322), .Z(n1807) );
  COND2XL U4153 ( .A(net17738), .B(n2320), .C(n123), .D(n2319), .Z(n1804) );
  COND2XL U4154 ( .A(net17738), .B(n2324), .C(n123), .D(n2323), .Z(n1808) );
  COND2XL U4155 ( .A(net17738), .B(n2321), .C(n123), .D(n2320), .Z(n1805) );
  CND2X1 U4156 ( .A(n3), .B(a[2]), .Z(n4423) );
  CAOR1XL U4157 ( .A(n3644), .B(net18896), .C(n2648), .Z(n2123) );
  CIVX3 U4158 ( .A(net18824), .Z(net16437) );
  CNIVX1 U4159 ( .A(n1170), .Z(n3791) );
  CND2X4 U4160 ( .A(n2812), .B(net16496), .Z(n144) );
  CENXL U4161 ( .A(n4572), .B(n4543), .Z(n2739) );
  CENXL U4162 ( .A(n4572), .B(n4546), .Z(n2736) );
  CENXL U4163 ( .A(n4572), .B(n4554), .Z(n2728) );
  CENXL U4164 ( .A(n4572), .B(n4553), .Z(n2729) );
  CENXL U4165 ( .A(n4572), .B(n4550), .Z(n2732) );
  CENXL U4166 ( .A(n4572), .B(net16102), .Z(n2716) );
  CENXL U4167 ( .A(n4573), .B(n4552), .Z(n2730) );
  CENXL U4168 ( .A(n4512), .B(n4541), .Z(n2742) );
  CENXL U4169 ( .A(n4512), .B(n4540), .Z(n2744) );
  CENXL U4170 ( .A(n4512), .B(n4545), .Z(n2737) );
  CENX1 U4171 ( .A(n4512), .B(n4564), .Z(n2715) );
  CENXL U4172 ( .A(n4573), .B(n4542), .Z(n2740) );
  CENXL U4173 ( .A(n4573), .B(n4547), .Z(n2735) );
  CENXL U4174 ( .A(n4573), .B(n4551), .Z(n2731) );
  CENXL U4175 ( .A(n4573), .B(n4549), .Z(n2733) );
  CNIVX4 U4176 ( .A(n3703), .Z(net16451) );
  CIVX4 U4177 ( .A(n136), .Z(n4604) );
  CENX2 U4178 ( .A(net18420), .B(n3836), .Z(net18218) );
  CIVX4 U4179 ( .A(n4093), .Z(n4577) );
  CEOX2 U4180 ( .A(n3792), .B(n1485), .Z(n1483) );
  CND2X1 U4181 ( .A(n1485), .B(n1487), .Z(n3794) );
  CEOX2 U4182 ( .A(n2140), .B(n2200), .Z(n3796) );
  CEOX2 U4183 ( .A(n3796), .B(n1925), .Z(n1539) );
  CND2XL U4184 ( .A(n1925), .B(n2200), .Z(n3797) );
  CND3X1 U4185 ( .A(n3797), .B(n3798), .C(n3799), .Z(n1538) );
  CENX1 U4186 ( .A(n3842), .B(n1538), .Z(n1515) );
  CEO3X1 U4187 ( .A(n1526), .B(n1509), .C(n1507), .Z(n1505) );
  CND2XL U4188 ( .A(n1526), .B(n1507), .Z(n3800) );
  CND2XL U4189 ( .A(n1526), .B(n1509), .Z(n3801) );
  CND2XL U4190 ( .A(n1507), .B(n1509), .Z(n3802) );
  CND3XL U4191 ( .A(n3800), .B(n3801), .C(n3802), .Z(n1504) );
  CEOX2 U4192 ( .A(n1533), .B(n1531), .Z(n3803) );
  CEOX2 U4193 ( .A(n3803), .B(n3612), .Z(n1527) );
  CND2X1 U4194 ( .A(n1548), .B(n1531), .Z(n3804) );
  CND2X1 U4195 ( .A(n1531), .B(n1533), .Z(n3806) );
  CND3X2 U4196 ( .A(n3804), .B(n3806), .C(n3805), .Z(n1526) );
  CND2X1 U4197 ( .A(n3972), .B(n3973), .Z(n1507) );
  CNR2X2 U4198 ( .A(net16974), .B(net16962), .Z(n3807) );
  CENXL U4199 ( .A(n4576), .B(n4567), .Z(n2644) );
  CENXL U4200 ( .A(n4576), .B(n4540), .Z(n2645) );
  CENXL U4201 ( .A(n4576), .B(n4547), .Z(n2636) );
  CENXL U4202 ( .A(n4576), .B(n4548), .Z(n2635) );
  CENXL U4203 ( .A(n4576), .B(n4543), .Z(n2640) );
  CENXL U4204 ( .A(n4576), .B(n4542), .Z(n2641) );
  CENXL U4205 ( .A(n4576), .B(n4541), .Z(n2643) );
  CENXL U4206 ( .A(n4576), .B(n4545), .Z(n2638) );
  CENXL U4207 ( .A(n4576), .B(n4549), .Z(n2634) );
  CANR1X1 U4208 ( .A(n669), .B(n677), .C(n670), .Z(n668) );
  CEO3X2 U4209 ( .A(n2150), .B(n1683), .C(n2119), .Z(n1679) );
  CND2X1 U4210 ( .A(n2150), .B(n1683), .Z(n3808) );
  CND2XL U4211 ( .A(n2150), .B(n2119), .Z(n3809) );
  CND2X1 U4212 ( .A(n1683), .B(n2119), .Z(n3810) );
  CND3X2 U4213 ( .A(n3808), .B(n3809), .C(n3810), .Z(n1678) );
  CEOX2 U4214 ( .A(n1673), .B(n1671), .Z(n3811) );
  CEOX2 U4215 ( .A(n3811), .B(n1678), .Z(n1667) );
  CND2XL U4216 ( .A(n1673), .B(n1671), .Z(n3812) );
  CND2XL U4217 ( .A(n1673), .B(n1678), .Z(n3813) );
  CND2XL U4218 ( .A(n1671), .B(n1678), .Z(n3814) );
  CND3X1 U4219 ( .A(n3812), .B(n3813), .C(n3814), .Z(n1666) );
  COND2X1 U4220 ( .A(n99), .B(n3877), .C(n2449), .D(n3771), .Z(n1729) );
  CND2XL U4221 ( .A(n1305), .B(n1332), .Z(net17791) );
  CND3X2 U4222 ( .A(n4527), .B(n4528), .C(n4529), .Z(n1370) );
  CENX1 U4223 ( .A(n3026), .B(n4543), .Z(n2475) );
  COND2XL U4224 ( .A(n4012), .B(n2402), .C(n2401), .D(net17425), .Z(n3816) );
  CAOR1XL U4225 ( .A(net16511), .B(n3991), .C(n2450), .Z(n1927) );
  COND2XL U4226 ( .A(n3991), .B(n2462), .C(net16511), .D(n2461), .Z(n1939) );
  COND2XL U4227 ( .A(n3991), .B(n2454), .C(net16511), .D(n2453), .Z(n1931) );
  CND2XL U4228 ( .A(n1826), .B(n2005), .Z(n3817) );
  CND2XL U4229 ( .A(n1826), .B(n1881), .Z(n3818) );
  CND2X1 U4230 ( .A(n2005), .B(n1881), .Z(n3819) );
  CND3X1 U4231 ( .A(n3817), .B(n3818), .C(n3819), .Z(n1208) );
  COR2X1 U4232 ( .A(net17738), .B(n2342), .Z(n3820) );
  COR2XL U4233 ( .A(n123), .B(n2341), .Z(n3821) );
  CND2X2 U4234 ( .A(n3820), .B(n3821), .Z(n1826) );
  CND2X1 U4235 ( .A(n1236), .B(n2065), .Z(n3923) );
  CIVX1 U4236 ( .A(n415), .Z(n413) );
  COR2XL U4237 ( .A(n3120), .B(n1275), .Z(n3822) );
  CENX1 U4238 ( .A(n3823), .B(n1217), .Z(n1215) );
  CIVX2 U4239 ( .A(n371), .Z(n4452) );
  CND2X1 U4240 ( .A(n1338), .B(n1315), .Z(n4159) );
  CEOX2 U4241 ( .A(n986), .B(n988), .Z(n3824) );
  CEOX2 U4242 ( .A(n3824), .B(n971), .Z(n965) );
  CND2X1 U4243 ( .A(n971), .B(n988), .Z(n3825) );
  CND2X1 U4244 ( .A(n971), .B(n986), .Z(n3826) );
  CND2XL U4245 ( .A(n988), .B(n986), .Z(n3827) );
  CND3X2 U4246 ( .A(n3825), .B(n3826), .C(n3827), .Z(n964) );
  CIVXL U4247 ( .A(net15916), .Z(n3828) );
  CND3XL U4248 ( .A(n4083), .B(n4082), .C(n4084), .Z(n3829) );
  CND2X2 U4249 ( .A(n4121), .B(n3986), .Z(n3831) );
  CND2X2 U4250 ( .A(n3830), .B(n3985), .Z(n3832) );
  CIVX2 U4251 ( .A(n4466), .Z(n3830) );
  CENX1 U4252 ( .A(n4595), .B(n4556), .Z(n2363) );
  CND3X1 U4253 ( .A(n4394), .B(n4395), .C(n4396), .Z(n1386) );
  CND2X1 U4254 ( .A(n4594), .B(n4198), .Z(n3834) );
  CND2X2 U4255 ( .A(n3834), .B(n3835), .Z(n105) );
  CENX1 U4256 ( .A(n3815), .B(n4563), .Z(n2553) );
  CNIVX4 U4257 ( .A(n30), .Z(n3836) );
  CIVX1 U4258 ( .A(n30), .Z(net15980) );
  CND3X2 U4259 ( .A(n4162), .B(n4163), .C(n4164), .Z(n1276) );
  CIVXL U4260 ( .A(n4559), .Z(n3837) );
  CNIVX4 U4261 ( .A(n2789), .Z(n4559) );
  CND3X2 U4262 ( .A(n4274), .B(n4275), .C(n4276), .Z(n1342) );
  COND1X1 U4263 ( .A(n633), .B(n637), .C(n634), .Z(n632) );
  CNIVX1 U4264 ( .A(n1987), .Z(n3979) );
  COR2XL U4265 ( .A(n1186), .B(n1159), .Z(n3840) );
  CENXL U4266 ( .A(n3833), .B(n4551), .Z(n2434) );
  CANR1XL U4267 ( .A(n748), .B(n415), .C(n408), .Z(n406) );
  CENX2 U4268 ( .A(n1401), .B(n1399), .Z(n3841) );
  CENX1 U4269 ( .A(n604), .B(n187), .Z(product[25]) );
  COND1X1 U4270 ( .A(n605), .B(n611), .C(n3171), .Z(n604) );
  CANR1XL U4271 ( .A(n3511), .B(n631), .C(n3788), .Z(n3843) );
  CIVX3 U4272 ( .A(a[22]), .Z(n4198) );
  CIVXL U4273 ( .A(n954), .Z(n955) );
  CIVX2 U4274 ( .A(n3718), .Z(n4591) );
  CANR1X1 U4275 ( .A(n631), .B(n3511), .C(n632), .Z(n630) );
  CEO3X2 U4276 ( .A(n1698), .B(n1691), .C(n1696), .Z(n1687) );
  CEOX2 U4277 ( .A(n1689), .B(n1694), .Z(n3844) );
  CEOX2 U4278 ( .A(n3844), .B(n1687), .Z(n1685) );
  CND2X1 U4279 ( .A(n1698), .B(n1691), .Z(n3845) );
  CND2X1 U4280 ( .A(n1698), .B(n1696), .Z(n3846) );
  CND2X1 U4281 ( .A(n1691), .B(n1696), .Z(n3847) );
  CND2XL U4282 ( .A(n1689), .B(n1694), .Z(n3848) );
  CND2XL U4283 ( .A(n1689), .B(n1687), .Z(n3849) );
  CND2XL U4284 ( .A(n1694), .B(n1687), .Z(n3850) );
  CND3X1 U4285 ( .A(n3848), .B(n3849), .C(n3850), .Z(n1684) );
  CIVXL U4286 ( .A(n260), .Z(n258) );
  CENX2 U4287 ( .A(n1606), .B(n1595), .Z(n4153) );
  CND2XL U4288 ( .A(n230), .B(n151), .Z(n3853) );
  CND2X1 U4289 ( .A(n3851), .B(n3852), .Z(n3854) );
  CND2X2 U4290 ( .A(n3853), .B(n3854), .Z(product[61]) );
  CIVXL U4291 ( .A(n230), .Z(n3851) );
  CIVX2 U4292 ( .A(n151), .Z(n3852) );
  CND2XL U4293 ( .A(n4498), .B(n229), .Z(n151) );
  CIVXL U4294 ( .A(n1034), .Z(n1035) );
  CEO3X2 U4295 ( .A(n1926), .B(n2201), .C(n2171), .Z(n1561) );
  CND2XL U4296 ( .A(n1926), .B(n2201), .Z(n3855) );
  CND2XL U4297 ( .A(n1926), .B(n2171), .Z(n3856) );
  CND3X1 U4298 ( .A(n3855), .B(n3856), .C(n3857), .Z(n1560) );
  CEOX1 U4299 ( .A(n2078), .B(n1543), .Z(n3858) );
  CND2X1 U4300 ( .A(n2078), .B(n1543), .Z(n3859) );
  CND2X1 U4301 ( .A(n2078), .B(n1560), .Z(n3860) );
  CND2X1 U4302 ( .A(n1543), .B(n1560), .Z(n3861) );
  CND3X2 U4303 ( .A(n3859), .B(n3860), .C(n3861), .Z(n1534) );
  CENX1 U4304 ( .A(n4591), .B(n4560), .Z(n2425) );
  CEO3X1 U4305 ( .A(n1522), .B(n1518), .C(n1516), .Z(n1493) );
  CND2X1 U4306 ( .A(n1516), .B(n1518), .Z(n3864) );
  CIVX1 U4307 ( .A(n275), .Z(n273) );
  CND2X1 U4308 ( .A(n1190), .B(n1192), .Z(n4135) );
  COND2X1 U4309 ( .A(n90), .B(n2468), .C(net16511), .D(n2467), .Z(n1945) );
  CIVX1 U4310 ( .A(n434), .Z(n432) );
  COND2XL U4311 ( .A(n45), .B(n2617), .C(net16420), .D(n2616), .Z(n2092) );
  CND2X1 U4312 ( .A(n1148), .B(n1150), .Z(n3867) );
  CND2X2 U4313 ( .A(n3865), .B(n3866), .Z(n3868) );
  CND2X2 U4314 ( .A(n3867), .B(n3868), .Z(net18574) );
  CIVX2 U4315 ( .A(n1150), .Z(n3866) );
  CND2X1 U4316 ( .A(n1281), .B(n1308), .Z(n4162) );
  COND2XL U4317 ( .A(net18310), .B(n2286), .C(net16439), .D(n2285), .Z(n1770)
         );
  COND2XL U4318 ( .A(net18310), .B(n2288), .C(net16439), .D(n2287), .Z(n1772)
         );
  COND2XL U4319 ( .A(net18310), .B(n2292), .C(net16439), .D(n2291), .Z(n1776)
         );
  COND2XL U4320 ( .A(net18310), .B(n2294), .C(net16439), .D(n2293), .Z(n1778)
         );
  COND2XL U4321 ( .A(net18310), .B(n2291), .C(net16439), .D(n2290), .Z(n1775)
         );
  COND2XL U4322 ( .A(net18310), .B(n2299), .C(net16439), .D(n2298), .Z(n1783)
         );
  COND2XL U4323 ( .A(n135), .B(n2297), .C(net16439), .D(n2296), .Z(n1781) );
  COND2XL U4324 ( .A(net18310), .B(n2302), .C(net16439), .D(n2301), .Z(n1786)
         );
  CNR2IXL U4325 ( .B(n3751), .A(net16439), .Z(n1801) );
  COND1X2 U4326 ( .A(n559), .B(n551), .C(n552), .Z(n550) );
  CEO3XL U4327 ( .A(n1365), .B(n1388), .C(n1363), .Z(n3869) );
  COND2XL U4328 ( .A(n4063), .B(n2618), .C(net16420), .D(n2617), .Z(n2093) );
  CAOR1XL U4329 ( .A(net16420), .B(n4063), .C(n2615), .Z(n2090) );
  CND2XL U4330 ( .A(n1792), .B(n2093), .Z(n3955) );
  CND2X1 U4331 ( .A(n1578), .B(n2110), .Z(n4108) );
  COND1XL U4332 ( .A(n643), .B(n3606), .C(n4218), .Z(n642) );
  CND2X1 U4333 ( .A(n1206), .B(n1210), .Z(n3872) );
  CND2X2 U4334 ( .A(n3870), .B(n3871), .Z(n3873) );
  CND2X2 U4335 ( .A(n3872), .B(n3873), .Z(n3910) );
  CIVXL U4336 ( .A(n1206), .Z(n3870) );
  CIVX2 U4337 ( .A(n1210), .Z(n3871) );
  CANR1XL U4338 ( .A(n396), .B(n415), .C(n3503), .Z(n395) );
  COND2XL U4339 ( .A(net16301), .B(n2545), .C(n3122), .D(n2544), .Z(n2022) );
  CND2XL U4340 ( .A(n746), .B(n392), .Z(n164) );
  CENXL U4341 ( .A(n4121), .B(n4541), .Z(n2577) );
  CENXL U4342 ( .A(n4121), .B(n4548), .Z(n2569) );
  COR2XL U4343 ( .A(net16420), .B(n2620), .Z(n4216) );
  CND2X1 U4344 ( .A(n1320), .B(n1301), .Z(n4101) );
  CND2X1 U4345 ( .A(n1320), .B(n1297), .Z(n4100) );
  CIVX2 U4346 ( .A(n4581), .Z(n4580) );
  CND2X2 U4347 ( .A(n4252), .B(n4253), .Z(n2820) );
  CND2X2 U4348 ( .A(n1193), .B(n1220), .Z(n4045) );
  CND2X1 U4349 ( .A(n272), .B(n736), .Z(n261) );
  CND2XL U4350 ( .A(n2127), .B(n1857), .Z(n4024) );
  CND2XL U4351 ( .A(n2034), .B(n1857), .Z(n4023) );
  CIVX4 U4352 ( .A(n3890), .Z(net17425) );
  CND2XL U4353 ( .A(n784), .B(n694), .Z(n202) );
  CENX1 U4354 ( .A(n4580), .B(n4544), .Z(n2573) );
  COND1XL U4355 ( .A(n4155), .B(n595), .C(n579), .Z(n3875) );
  CND2X2 U4356 ( .A(n3785), .B(n3877), .Z(n3878) );
  CND2X1 U4357 ( .A(n3876), .B(n3833), .Z(n3879) );
  CND2X2 U4358 ( .A(n4467), .B(n3783), .Z(n4468) );
  CENX2 U4359 ( .A(n1199), .B(n3880), .Z(n1193) );
  CEO3XL U4360 ( .A(n943), .B(n941), .C(n958), .Z(n3882) );
  CENX1 U4361 ( .A(n4580), .B(n4562), .Z(n2555) );
  CND2X1 U4362 ( .A(n1308), .B(n1283), .Z(n4164) );
  CENX2 U4363 ( .A(a[6]), .B(n3836), .Z(net16974) );
  COND2XL U4364 ( .A(net17738), .B(n2330), .C(n123), .D(n2329), .Z(n1814) );
  CND2X1 U4365 ( .A(n1538), .B(n1540), .Z(n3883) );
  CND2X1 U4366 ( .A(n1538), .B(n1542), .Z(n3884) );
  CND2X1 U4367 ( .A(n1540), .B(n1542), .Z(n3885) );
  CND3X2 U4368 ( .A(n3883), .B(n3884), .C(n3885), .Z(n1514) );
  CIVX1 U4369 ( .A(n920), .Z(n921) );
  CND2X2 U4370 ( .A(n3887), .B(n3888), .Z(n1855) );
  CND2X1 U4371 ( .A(n2815), .B(n3889), .Z(n3888) );
  CNR2XL U4372 ( .A(n2371), .B(n3921), .Z(n3889) );
  COR2X1 U4373 ( .A(n2370), .B(net16433), .Z(n3887) );
  CENX2 U4374 ( .A(n4595), .B(n4548), .Z(n2371) );
  CENX1 U4375 ( .A(n4595), .B(n4549), .Z(n2370) );
  CIVX2 U4376 ( .A(a[12]), .Z(n4370) );
  CENX4 U4377 ( .A(n3026), .B(n3785), .Z(n3891) );
  COND2X1 U4378 ( .A(n27), .B(n2697), .C(net16451), .D(n2696), .Z(n2171) );
  CND2X1 U4379 ( .A(n748), .B(n410), .Z(n166) );
  CIVX2 U4380 ( .A(n410), .Z(n408) );
  CND2X2 U4381 ( .A(n923), .B(n938), .Z(n410) );
  CENX2 U4382 ( .A(a[28]), .B(n4601), .Z(n2813) );
  CIVX8 U4383 ( .A(n4601), .Z(n4600) );
  CND2XL U4384 ( .A(n1728), .B(n3974), .Z(n3975) );
  CND2XL U4385 ( .A(n1351), .B(n1357), .Z(n4274) );
  CIVX2 U4386 ( .A(n48), .Z(n3892) );
  CIVXL U4387 ( .A(n48), .Z(n4058) );
  CENX2 U4388 ( .A(n3895), .B(n1143), .Z(n1139) );
  COR2XL U4389 ( .A(n2717), .B(n4510), .Z(n4247) );
  CND2IX2 U4390 ( .B(n3986), .A(n4251), .Z(n4252) );
  CIVX2 U4391 ( .A(n644), .Z(n646) );
  CND2XL U4392 ( .A(n1439), .B(n1441), .Z(n4035) );
  CEOX4 U4393 ( .A(a[30]), .B(n4603), .Z(n2812) );
  COND1X1 U4394 ( .A(n613), .B(n3843), .C(n3610), .Z(n3896) );
  COND1X1 U4395 ( .A(n613), .B(n630), .C(n614), .Z(n612) );
  CANR1X1 U4396 ( .A(n554), .B(n574), .C(n555), .Z(n553) );
  CNR2X2 U4397 ( .A(n353), .B(n261), .Z(n259) );
  COND1X2 U4398 ( .A(n3354), .B(net16471), .C(n3684), .Z(n459) );
  CND2X1 U4399 ( .A(n396), .B(n363), .Z(n361) );
  CND2X1 U4400 ( .A(n3897), .B(n3898), .Z(n1892) );
  CIVX1 U4401 ( .A(n2414), .Z(n3900) );
  CIVX1 U4402 ( .A(n2415), .Z(n3901) );
  CND2X1 U4403 ( .A(n3899), .B(n3900), .Z(n3897) );
  CND2X1 U4404 ( .A(n3901), .B(n3902), .Z(n3898) );
  CND2X1 U4405 ( .A(n1059), .B(n1082), .Z(n485) );
  CIVX2 U4406 ( .A(a[10]), .Z(n3992) );
  CNIVX2 U4407 ( .A(n57), .Z(n4466) );
  CND2XL U4408 ( .A(n1565), .B(n1567), .Z(n4516) );
  COND2X1 U4409 ( .A(n2691), .B(n27), .C(net16451), .D(n2690), .Z(n2165) );
  CEOX2 U4410 ( .A(n3785), .B(n4593), .Z(n2817) );
  CENX1 U4411 ( .A(n3815), .B(n4557), .Z(n2560) );
  CENX1 U4412 ( .A(net18828), .B(n4552), .Z(n2697) );
  CIVX2 U4413 ( .A(n3782), .Z(n4251) );
  CND2XL U4414 ( .A(n1389), .B(n1414), .Z(n4395) );
  CND2XL U4415 ( .A(n1389), .B(n1391), .Z(n4394) );
  CND3XL U4416 ( .A(n4537), .B(n4538), .C(n4539), .Z(n3905) );
  CIVX8 U4417 ( .A(n4596), .Z(n4595) );
  CIVXL U4418 ( .A(n674), .Z(n781) );
  CEO3XL U4419 ( .A(n1536), .B(n1521), .C(n1523), .Z(n4065) );
  CND3X1 U4420 ( .A(n3980), .B(n3981), .C(n3982), .Z(n1536) );
  COND2X1 U4421 ( .A(n81), .B(n2496), .C(net16413), .D(n2495), .Z(n1973) );
  CENXL U4422 ( .A(n4585), .B(n4556), .Z(n2495) );
  COND2X1 U4423 ( .A(n4012), .B(n2407), .C(n2406), .D(net16426), .Z(n1884) );
  COND2X1 U4424 ( .A(n4184), .B(n2595), .C(n4506), .D(n2594), .Z(n2070) );
  CENX1 U4425 ( .A(n4579), .B(n4556), .Z(n2594) );
  CND2X1 U4426 ( .A(n1409), .B(n1403), .Z(n4406) );
  CANR1X1 U4427 ( .A(n331), .B(n356), .C(n332), .Z(n330) );
  CIVXL U4428 ( .A(n334), .Z(n332) );
  CENX2 U4429 ( .A(n1283), .B(n1308), .Z(n3913) );
  CENX1 U4430 ( .A(n4579), .B(n4558), .Z(n2592) );
  CND2IX2 U4431 ( .B(net15988), .A(net17482), .Z(net17483) );
  CNIVX3 U4432 ( .A(n21), .Z(net18828) );
  CNIVX4 U4433 ( .A(n2792), .Z(n4556) );
  CIVX2 U4434 ( .A(n4476), .Z(n4212) );
  CIVXL U4435 ( .A(n529), .Z(n760) );
  CND2X1 U4436 ( .A(n1426), .B(n1403), .Z(n4407) );
  CANR1XL U4437 ( .A(n3896), .B(n3177), .C(n3875), .Z(n3911) );
  CENX2 U4438 ( .A(n4578), .B(n3992), .Z(n4462) );
  CENX2 U4439 ( .A(n3913), .B(n1281), .Z(n1277) );
  CND2X2 U4440 ( .A(net17483), .B(n3914), .Z(net16962) );
  CND2X2 U4441 ( .A(net17483), .B(n3914), .Z(net18261) );
  CIVX2 U4442 ( .A(n21), .Z(net15988) );
  CND2XL U4443 ( .A(n1145), .B(n1147), .Z(n3918) );
  CND2X1 U4444 ( .A(n1143), .B(n1147), .Z(n3917) );
  CND2XL U4445 ( .A(n1143), .B(n1145), .Z(n3916) );
  CND2X1 U4446 ( .A(n1166), .B(n1168), .Z(n3915) );
  CND2X1 U4447 ( .A(n1141), .B(n1166), .Z(net17989) );
  CND2X1 U4448 ( .A(n1141), .B(n1168), .Z(net17987) );
  CND2XL U4449 ( .A(n1089), .B(n1112), .Z(net18200) );
  CND2XL U4450 ( .A(n1150), .B(n1152), .Z(net18534) );
  CND2XL U4451 ( .A(n1148), .B(n1150), .Z(net18532) );
  CND3X2 U4452 ( .A(net17725), .B(net17723), .C(net17724), .Z(n1170) );
  CND2X1 U4453 ( .A(n1181), .B(n1208), .Z(net17724) );
  CND2X1 U4454 ( .A(n1181), .B(n1183), .Z(net17725) );
  CND2X1 U4455 ( .A(n1183), .B(n1208), .Z(net17723) );
  CEO3X1 U4456 ( .A(n1942), .B(n2033), .C(n2064), .Z(n1181) );
  CENXL U4457 ( .A(net15974), .B(net16104), .Z(n3920) );
  CIVX8 U4458 ( .A(n3921), .Z(net16433) );
  CIVX3 U4459 ( .A(n114), .Z(n3921) );
  CENX1 U4460 ( .A(a[24]), .B(n102), .Z(n114) );
  CNIVX4 U4461 ( .A(n2783), .Z(net16104) );
  COND2XL U4462 ( .A(net18896), .B(net15980), .C(n2680), .D(n3644), .Z(n1736)
         );
  CND2X2 U4463 ( .A(net18419), .B(a[8]), .Z(net18422) );
  CIVX2 U4464 ( .A(n3836), .Z(net18419) );
  CND2XL U4465 ( .A(net18419), .B(net18505), .Z(net18507) );
  CND2X1 U4466 ( .A(n3836), .B(net18420), .Z(n3926) );
  COND2X1 U4467 ( .A(net17728), .B(n2403), .C(n2402), .D(net17425), .Z(n1880)
         );
  CND2X1 U4468 ( .A(n1115), .B(n1140), .Z(net17756) );
  CND2X1 U4469 ( .A(n3143), .B(n1140), .Z(net17755) );
  CND2XL U4470 ( .A(n1173), .B(n1175), .Z(net17985) );
  CND2XL U4471 ( .A(n1200), .B(n1175), .Z(net17984) );
  CND2X1 U4472 ( .A(n2188), .B(n2096), .Z(n3930) );
  CND3X2 U4473 ( .A(n3931), .B(n3932), .C(n3933), .Z(n1172) );
  CND2X1 U4474 ( .A(n1210), .B(n1206), .Z(n3933) );
  CND2X1 U4475 ( .A(n1204), .B(n1206), .Z(n3932) );
  CND2X1 U4476 ( .A(n1204), .B(n1210), .Z(n3931) );
  CND3X1 U4477 ( .A(n3927), .B(net17984), .C(net17985), .Z(n1166) );
  CNIVXL U4478 ( .A(n1166), .Z(net18863) );
  CND2XL U4479 ( .A(n1200), .B(n1173), .Z(n3927) );
  CND2X1 U4480 ( .A(n1083), .B(n1106), .Z(n494) );
  COR2XL U4481 ( .A(n1132), .B(n1107), .Z(net18519) );
  CND2X1 U4482 ( .A(n1107), .B(n1132), .Z(n505) );
  COND1X1 U4483 ( .A(n512), .B(n504), .C(n505), .Z(n499) );
  CANR1X1 U4484 ( .A(n482), .B(n499), .C(n483), .Z(n481) );
  CND2X2 U4485 ( .A(n1133), .B(n1158), .Z(n512) );
  CIVXL U4486 ( .A(n512), .Z(n510) );
  CND2XL U4487 ( .A(n758), .B(n512), .Z(n176) );
  COAN1XL U4488 ( .A(n512), .B(n504), .C(n505), .Z(net18400) );
  CNR2X2 U4489 ( .A(n504), .B(n511), .Z(n498) );
  CND2XL U4490 ( .A(net18519), .B(n505), .Z(n175) );
  CNR2X2 U4491 ( .A(n3528), .B(n1133), .Z(n511) );
  CEO3X2 U4492 ( .A(n2156), .B(n1184), .C(n2125), .Z(n1157) );
  CND2XL U4493 ( .A(n1184), .B(n3723), .Z(net18593) );
  CND2XL U4494 ( .A(n1184), .B(n2125), .Z(net18592) );
  COND1X1 U4495 ( .A(n3397), .B(n515), .C(n481), .Z(n479) );
  COND1X1 U4496 ( .A(n484), .B(n494), .C(n485), .Z(n483) );
  COND1XL U4497 ( .A(n3757), .B(net18400), .C(n494), .Z(n490) );
  CAN2XL U4498 ( .A(n485), .B(net18527), .Z(net17136) );
  COR2XL U4499 ( .A(n1082), .B(n1059), .Z(net18527) );
  CNIVX4 U4500 ( .A(n149), .Z(net16471) );
  CANR1X1 U4501 ( .A(n478), .B(n546), .C(n479), .Z(n149) );
  CIVX2 U4502 ( .A(n468), .Z(n753) );
  CND2XL U4503 ( .A(n753), .B(n469), .Z(n171) );
  COND1X1 U4504 ( .A(n444), .B(n461), .C(n445), .Z(net19057) );
  COND1X1 U4505 ( .A(n444), .B(n3683), .C(n445), .Z(n439) );
  CIVX2 U4506 ( .A(n472), .Z(n474) );
  CNR2X1 U4507 ( .A(n514), .B(n3397), .Z(n478) );
  CANR1X1 U4508 ( .A(n478), .B(n546), .C(n479), .Z(net18832) );
  CANR1X1 U4509 ( .A(net17942), .B(n535), .C(n3409), .Z(n515) );
  CNR2X1 U4510 ( .A(n529), .B(n522), .Z(net17942) );
  CND2X1 U4511 ( .A(net17942), .B(n534), .Z(n514) );
  CANR1XL U4512 ( .A(n760), .B(n3695), .C(n528), .Z(n526) );
  CANR1XL U4513 ( .A(n520), .B(n3037), .C(n3234), .Z(net16274) );
  CIVXL U4514 ( .A(n3911), .Z(net18614) );
  CIVXL U4515 ( .A(n562), .Z(n564) );
  CNIVXL U4516 ( .A(n562), .Z(net18204) );
  CNR2X2 U4517 ( .A(n551), .B(n556), .Z(n549) );
  CNR2X2 U4518 ( .A(n1305), .B(n1332), .Z(n556) );
  CANR1X1 U4519 ( .A(n561), .B(n574), .C(net18204), .Z(n560) );
  CNR2IXL U4520 ( .B(n561), .A(n556), .Z(n554) );
  CND2XL U4521 ( .A(n3572), .B(n458), .Z(n170) );
  COR2X1 U4522 ( .A(n995), .B(n1014), .Z(n3937) );
  CND2XL U4523 ( .A(n462), .B(n3572), .Z(n451) );
  CANR1XL U4524 ( .A(n3572), .B(n3731), .C(n456), .Z(n452) );
  CND2X1 U4525 ( .A(n995), .B(n1014), .Z(n458) );
  CND2X1 U4526 ( .A(n3938), .B(net18507), .Z(n2650) );
  COR2X1 U4527 ( .A(net18610), .B(n2650), .Z(net18496) );
  CIVXL U4528 ( .A(net16102), .Z(net18505) );
  CNIVX4 U4529 ( .A(n2782), .Z(net16102) );
  COND2XL U4530 ( .A(n90), .B(n2465), .C(n2464), .D(net16512), .Z(n3939) );
  CND2XL U4531 ( .A(n1605), .B(n1616), .Z(n3940) );
  CND2XL U4532 ( .A(n1605), .B(n1603), .Z(n3941) );
  CND2XL U4533 ( .A(n1616), .B(n1603), .Z(n3942) );
  CND3X1 U4534 ( .A(n3940), .B(n3942), .C(n3941), .Z(n1598) );
  CND2XL U4535 ( .A(n1601), .B(n1614), .Z(n3943) );
  CND2XL U4536 ( .A(n1599), .B(n1601), .Z(n3944) );
  CND2XL U4537 ( .A(n1614), .B(n1599), .Z(n3945) );
  CND3X1 U4538 ( .A(n3943), .B(n3944), .C(n3945), .Z(n1596) );
  CEO3X2 U4539 ( .A(n1625), .B(n1621), .C(n1623), .Z(n1617) );
  CND2XL U4540 ( .A(n1625), .B(n1623), .Z(n3946) );
  CND2X1 U4541 ( .A(n1625), .B(n1621), .Z(n3947) );
  CND2X1 U4542 ( .A(n1623), .B(n1621), .Z(n3948) );
  CND3X2 U4543 ( .A(n3946), .B(n3947), .C(n3948), .Z(n1616) );
  CIVX3 U4544 ( .A(n4578), .Z(n4037) );
  CENX1 U4545 ( .A(net19060), .B(net16472), .Z(product[40]) );
  CND2X1 U4546 ( .A(n3461), .B(n4329), .Z(n4331) );
  COND1X1 U4547 ( .A(n268), .B(net16472), .C(n269), .Z(n267) );
  COND2XL U4548 ( .A(net17727), .B(n2388), .C(n2387), .D(net17425), .Z(n1870)
         );
  CFA1XL U4549 ( .A(n842), .B(n1868), .CI(n1837), .CO(n832), .S(n833) );
  CIVXL U4550 ( .A(n842), .Z(n843) );
  CIVX2 U4551 ( .A(n54), .Z(n4183) );
  CND2X2 U4552 ( .A(n3950), .B(n4397), .Z(n3952) );
  CND2X2 U4553 ( .A(n3951), .B(n3952), .Z(n87) );
  CNIVX4 U4554 ( .A(n87), .Z(net16511) );
  CENXL U4555 ( .A(n4121), .B(n4546), .Z(n2571) );
  CENXL U4556 ( .A(n4121), .B(n4549), .Z(n2568) );
  CENXL U4557 ( .A(n2809), .B(n4121), .Z(n2578) );
  CEO3X1 U4558 ( .A(n1761), .B(n1792), .C(n2093), .Z(n1127) );
  CND2XL U4559 ( .A(n1761), .B(n1792), .Z(n3953) );
  CND2XL U4560 ( .A(n1761), .B(n2093), .Z(n3954) );
  CND3X1 U4561 ( .A(n3953), .B(n3954), .C(n3955), .Z(n1126) );
  CND2XL U4562 ( .A(n1122), .B(n1124), .Z(n3956) );
  CND2XL U4563 ( .A(n1124), .B(n1126), .Z(n3957) );
  CND2XL U4564 ( .A(n1122), .B(n1126), .Z(n3958) );
  CND3X1 U4565 ( .A(n3956), .B(n3957), .C(n3958), .Z(n1094) );
  CIVX4 U4566 ( .A(net15916), .Z(net15912) );
  CNIVX4 U4567 ( .A(net15914), .Z(net17419) );
  CEO3X2 U4568 ( .A(n1269), .B(n1290), .C(n1263), .Z(n1255) );
  COR2XL U4569 ( .A(n2649), .B(n3644), .Z(n4096) );
  CND2IX2 U4570 ( .B(n1513), .A(n4019), .Z(n4021) );
  CND2XL U4571 ( .A(a[4]), .B(n3766), .Z(n3960) );
  CND2X2 U4572 ( .A(n3960), .B(n3961), .Z(n2825) );
  CIVXL U4573 ( .A(n3766), .Z(net19006) );
  CND2XL U4574 ( .A(n2170), .B(n2231), .Z(n4284) );
  CND2X1 U4575 ( .A(n3962), .B(n3173), .Z(n3964) );
  CND2X2 U4576 ( .A(n3963), .B(n3964), .Z(n4078) );
  CEOX2 U4577 ( .A(n1459), .B(n1478), .Z(n3965) );
  CEOX2 U4578 ( .A(n3965), .B(n1480), .Z(n1449) );
  CND2XL U4579 ( .A(n1480), .B(n1478), .Z(n3966) );
  CND2XL U4580 ( .A(n1480), .B(n3176), .Z(n3967) );
  CND2XL U4581 ( .A(n1478), .B(n1459), .Z(n3968) );
  CND3X1 U4582 ( .A(n3966), .B(n3967), .C(n3968), .Z(n1448) );
  CND2XL U4583 ( .A(n1505), .B(n1524), .Z(n3969) );
  CND2X1 U4584 ( .A(n4207), .B(n1528), .Z(n3972) );
  CND2X2 U4585 ( .A(n3970), .B(n3971), .Z(n3973) );
  CIVX2 U4586 ( .A(n4207), .Z(n3970) );
  CIVX1 U4587 ( .A(n1528), .Z(n3971) );
  CFA1XL U4588 ( .A(n1931), .B(n1872), .CI(n1900), .CO(n934), .S(n935) );
  CND2X1 U4589 ( .A(n3427), .B(n2084), .Z(n4361) );
  CND2X1 U4590 ( .A(n3975), .B(n3976), .Z(n1503) );
  CIVXL U4591 ( .A(n2138), .Z(n3974) );
  CNR2X1 U4592 ( .A(n665), .B(n660), .Z(n658) );
  CIVXL U4593 ( .A(n665), .Z(n779) );
  CENXL U4594 ( .A(n3165), .B(n2809), .Z(n2545) );
  CND2X1 U4595 ( .A(n1086), .B(n1065), .Z(n4054) );
  COND2X1 U4596 ( .A(n4461), .B(n2719), .C(n2718), .D(n4510), .Z(n2192) );
  CNR2X2 U4597 ( .A(n4266), .B(n1524), .Z(n622) );
  CND3X1 U4598 ( .A(n4103), .B(n4104), .C(n4105), .Z(n1524) );
  CND2X1 U4599 ( .A(n1372), .B(n1349), .Z(n4158) );
  CENX1 U4600 ( .A(n1225), .B(n1252), .Z(n3977) );
  CND2XL U4601 ( .A(n747), .B(n403), .Z(n165) );
  CEO3X2 U4602 ( .A(n1454), .B(n1433), .C(n1435), .Z(n1423) );
  CEOX1 U4603 ( .A(n2042), .B(n1920), .Z(n4219) );
  CENX2 U4604 ( .A(n3978), .B(n1385), .Z(n1373) );
  CNR2X2 U4605 ( .A(n333), .B(n324), .Z(n320) );
  CEOX2 U4606 ( .A(n190), .B(n624), .Z(product[22]) );
  CANR1X2 U4607 ( .A(n773), .B(n629), .C(n626), .Z(n624) );
  CND2X1 U4608 ( .A(n259), .B(n3759), .Z(n248) );
  CENX1 U4609 ( .A(n4085), .B(n4555), .Z(n2463) );
  CND2XL U4610 ( .A(n2018), .B(n2109), .Z(n3980) );
  CND2XL U4611 ( .A(n2018), .B(n1956), .Z(n3981) );
  CND2XL U4612 ( .A(n2109), .B(n1956), .Z(n3982) );
  COR2XL U4613 ( .A(n3122), .B(n2540), .Z(n3984) );
  CND2X2 U4614 ( .A(n3983), .B(n3984), .Z(n2018) );
  CND3X2 U4615 ( .A(n4405), .B(n4406), .C(n4407), .Z(n1396) );
  CND2X4 U4616 ( .A(n3115), .B(n2817), .Z(n99) );
  CIVX2 U4617 ( .A(n1511), .Z(n4019) );
  CENX1 U4618 ( .A(n3908), .B(n4554), .Z(n2662) );
  CND2X4 U4619 ( .A(n2815), .B(net16433), .Z(n117) );
  CND3X1 U4620 ( .A(n4381), .B(n4382), .C(n4383), .Z(n1274) );
  CIVXL U4621 ( .A(n664), .Z(n3987) );
  CIVXL U4622 ( .A(n659), .Z(n3988) );
  CIVXL U4623 ( .A(n3988), .Z(n3989) );
  CNR2X1 U4624 ( .A(n1274), .B(n1245), .Z(n543) );
  CFA1X2 U4625 ( .A(n1943), .B(n2157), .CI(n1912), .CO(n1210), .S(n1211) );
  CND3X1 U4626 ( .A(n4022), .B(n4023), .C(n4024), .Z(n1206) );
  CEO3X2 U4627 ( .A(n2195), .B(n1982), .C(n1951), .Z(n1431) );
  CND2X4 U4628 ( .A(n4399), .B(n4400), .Z(n2818) );
  COND2X1 U4629 ( .A(n27), .B(n2684), .C(net17297), .D(n2683), .Z(n2158) );
  CENXL U4630 ( .A(n4587), .B(n2785), .Z(n2455) );
  CENXL U4631 ( .A(n4587), .B(net16104), .Z(n2453) );
  CENXL U4632 ( .A(n4587), .B(n4563), .Z(n2454) );
  CENXL U4633 ( .A(n4587), .B(net16102), .Z(n2452) );
  CENXL U4634 ( .A(n4587), .B(n4562), .Z(n2456) );
  CENXL U4635 ( .A(n4587), .B(n4557), .Z(n2461) );
  CENXL U4636 ( .A(n4587), .B(n4561), .Z(n2457) );
  CENXL U4637 ( .A(n4587), .B(n4560), .Z(n2458) );
  CENXL U4638 ( .A(n4587), .B(n4558), .Z(n2460) );
  CENXL U4639 ( .A(n4587), .B(n4559), .Z(n2459) );
  CENX1 U4640 ( .A(n4587), .B(n4556), .Z(n2462) );
  CENX1 U4641 ( .A(n328), .B(n159), .Z(product[53]) );
  CND2X2 U4642 ( .A(n3994), .B(n3995), .Z(n2822) );
  COND2XL U4643 ( .A(net16309), .B(n2672), .C(n3644), .D(n2671), .Z(n2147) );
  COND2XL U4644 ( .A(net18897), .B(n2673), .C(net16490), .D(n2672), .Z(n2148)
         );
  COND1X1 U4645 ( .A(n678), .B(n3027), .C(n3997), .Z(n3996) );
  CANR1X1 U4646 ( .A(n686), .B(n4488), .C(n681), .Z(n3997) );
  COND2X1 U4647 ( .A(n27), .B(n2695), .C(net17297), .D(n2694), .Z(n2169) );
  CND2X1 U4648 ( .A(n1556), .B(n1558), .Z(n4191) );
  CEO3X1 U4649 ( .A(n2050), .B(n2021), .C(n1990), .Z(n1593) );
  CEO3X2 U4650 ( .A(n1282), .B(n1255), .C(n3365), .Z(n1249) );
  CEO3X2 U4651 ( .A(n1228), .B(n1203), .C(n1201), .Z(n1195) );
  CND2XL U4652 ( .A(n1201), .B(n1228), .Z(n4001) );
  CND2XL U4653 ( .A(n1228), .B(n1203), .Z(n4002) );
  CND2XL U4654 ( .A(n1201), .B(n1203), .Z(n4003) );
  CND3X1 U4655 ( .A(n4001), .B(n4003), .C(n4002), .Z(n1194) );
  CND2X1 U4656 ( .A(n4242), .B(n1135), .Z(n4006) );
  CND2X2 U4657 ( .A(n4004), .B(n4005), .Z(n4007) );
  CND2X2 U4658 ( .A(n4006), .B(n4007), .Z(n1133) );
  CIVX2 U4659 ( .A(n4242), .Z(n4004) );
  COND2XL U4660 ( .A(n4461), .B(n2745), .C(n2744), .D(n4510), .Z(n2218) );
  CND2X1 U4661 ( .A(n280), .B(n155), .Z(n4010) );
  CND2X2 U4662 ( .A(n4008), .B(n4009), .Z(n4011) );
  CND2X2 U4663 ( .A(n4010), .B(n4011), .Z(product[57]) );
  CIVX2 U4664 ( .A(n280), .Z(n4008) );
  CIVX2 U4665 ( .A(n155), .Z(n4009) );
  CND2XL U4666 ( .A(n4490), .B(n279), .Z(n155) );
  CND2XL U4667 ( .A(n2021), .B(n1990), .Z(n4178) );
  COND2X1 U4668 ( .A(n81), .B(n2486), .C(n4217), .D(n2485), .Z(n1963) );
  CIVXL U4669 ( .A(net16541), .Z(net18827) );
  CENXL U4670 ( .A(n4580), .B(n4558), .Z(n2559) );
  CENXL U4671 ( .A(n4580), .B(n4559), .Z(n2558) );
  CIVX3 U4672 ( .A(n102), .Z(net15916) );
  CND2X1 U4673 ( .A(n1190), .B(n1165), .Z(n4136) );
  CNIVXL U4674 ( .A(n3206), .Z(net18817) );
  CENXL U4675 ( .A(n3828), .B(net16102), .Z(n2386) );
  CENXL U4676 ( .A(net15910), .B(n4562), .Z(n2390) );
  CENXL U4677 ( .A(net15910), .B(net16104), .Z(n2387) );
  CND2XL U4678 ( .A(n1121), .B(n1127), .Z(n4290) );
  CND2XL U4679 ( .A(n1121), .B(n1146), .Z(n4292) );
  COND2X1 U4680 ( .A(n4461), .B(n2722), .C(n2721), .D(n4510), .Z(n2195) );
  CAOR1XL U4681 ( .A(n4217), .B(n81), .C(n2483), .Z(n1960) );
  COND2XL U4682 ( .A(n81), .B(n2513), .C(n3789), .D(n2512), .Z(n1990) );
  CNR2XL U4683 ( .A(n353), .B(n224), .Z(n222) );
  CENX1 U4684 ( .A(n4579), .B(n4553), .Z(n2597) );
  CND2X2 U4685 ( .A(n105), .B(n2816), .Z(n4012) );
  CND2X1 U4686 ( .A(n2816), .B(n3084), .Z(n4013) );
  CIVX1 U4687 ( .A(n120), .Z(n4311) );
  CND2XL U4688 ( .A(n760), .B(n3214), .Z(n178) );
  CIVXL U4689 ( .A(n417), .Z(n419) );
  CENXL U4690 ( .A(net15974), .B(n4564), .Z(n2649) );
  CND2X1 U4691 ( .A(n1425), .B(n1446), .Z(n4185) );
  CNIVX4 U4692 ( .A(n87), .Z(net16510) );
  CND3X2 U4693 ( .A(n4156), .B(n4157), .C(n4158), .Z(n1340) );
  CNR2XL U4694 ( .A(n522), .B(n529), .Z(n520) );
  CNR2IX1 U4695 ( .B(n3244), .A(n4505), .Z(n2056) );
  CND2X1 U4696 ( .A(n4267), .B(n4268), .Z(n4017) );
  CND2X2 U4697 ( .A(n4015), .B(n4016), .Z(n4018) );
  CIVX2 U4698 ( .A(n4268), .Z(n4016) );
  CND2X4 U4699 ( .A(n24), .B(n2825), .Z(net18772) );
  CND2X1 U4700 ( .A(n1513), .B(n1511), .Z(n4020) );
  CND2X2 U4701 ( .A(n4020), .B(n4021), .Z(n4207) );
  CND2XL U4702 ( .A(n2034), .B(n2127), .Z(n4022) );
  CIVX8 U4703 ( .A(n4520), .Z(n4579) );
  COND2X1 U4704 ( .A(n144), .B(n2281), .C(n2280), .D(n3277), .Z(n1765) );
  CIVXL U4705 ( .A(n3752), .Z(n4025) );
  CNIVXL U4706 ( .A(n3816), .Z(n4026) );
  CENXL U4707 ( .A(n4579), .B(n4544), .Z(n2606) );
  CENXL U4708 ( .A(n4579), .B(n4564), .Z(n2583) );
  CENX1 U4709 ( .A(n4579), .B(n4560), .Z(n2590) );
  CEO3X2 U4710 ( .A(n1354), .B(n1350), .C(n1352), .Z(n1319) );
  CND2XL U4711 ( .A(n1354), .B(n1352), .Z(n4027) );
  CND2XL U4712 ( .A(n1354), .B(n1350), .Z(n4028) );
  CND2X1 U4713 ( .A(n1352), .B(n1350), .Z(n4029) );
  CIVX3 U4714 ( .A(a[2]), .Z(n4422) );
  CND2X1 U4715 ( .A(n1244), .B(n1215), .Z(n541) );
  CENX1 U4716 ( .A(net15912), .B(n4550), .Z(n2402) );
  CIVXL U4717 ( .A(n864), .Z(n865) );
  CFA1XL U4718 ( .A(n864), .B(n1777), .CI(n1808), .CO(n852), .S(n853) );
  COND2XL U4719 ( .A(net17279), .B(n2535), .C(n3121), .D(n2534), .Z(n2012) );
  CHA1X1 U4720 ( .A(n2047), .B(n1729), .CO(n1542), .S(n1543) );
  COND2X1 U4721 ( .A(n4316), .B(n2572), .C(n2571), .D(n4505), .Z(n2047) );
  CIVXL U4722 ( .A(n397), .Z(n399) );
  CENX1 U4723 ( .A(n4153), .B(n1593), .Z(n1587) );
  CEO3X1 U4724 ( .A(n1462), .B(n1441), .C(n3787), .Z(n1437) );
  CND2XL U4725 ( .A(n3787), .B(n3320), .Z(n4033) );
  CND2XL U4726 ( .A(n3320), .B(n1441), .Z(n4034) );
  CND3X1 U4727 ( .A(n4033), .B(n4034), .C(n4035), .Z(n1436) );
  CIVXL U4728 ( .A(n102), .Z(net18718) );
  COND2X1 U4729 ( .A(net18310), .B(n2315), .C(net16439), .D(n2314), .Z(n1799)
         );
  CND2XL U4730 ( .A(n3603), .B(n3454), .Z(n4416) );
  CNR2X2 U4731 ( .A(n4350), .B(n4269), .Z(n4351) );
  CIVX3 U4732 ( .A(n39), .Z(n4578) );
  CENXL U4733 ( .A(n1528), .B(n4207), .Z(n4038) );
  CND2X1 U4734 ( .A(n12), .B(a[4]), .Z(n4039) );
  CENX1 U4735 ( .A(n1466), .B(n1464), .Z(n4151) );
  CNR2X2 U4736 ( .A(n1159), .B(n1186), .Z(n522) );
  CIVX3 U4737 ( .A(n3678), .Z(n4571) );
  CNR2X2 U4738 ( .A(n3196), .B(n385), .Z(n383) );
  CND2X1 U4739 ( .A(n658), .B(n4169), .Z(n651) );
  CFA1X1 U4740 ( .A(n1843), .B(n1871), .CI(n1812), .CO(n902), .S(n903) );
  COND2X1 U4741 ( .A(n3301), .B(n2390), .C(n2389), .D(net17425), .Z(n1871) );
  COND1X1 U4742 ( .A(n392), .B(n365), .C(n366), .Z(n364) );
  CND3X1 U4743 ( .A(n4516), .B(n4517), .C(n4518), .Z(n1562) );
  CEOX1 U4744 ( .A(n1725), .B(n2192), .Z(n1359) );
  CND3X2 U4745 ( .A(n4043), .B(n4044), .C(n4045), .Z(n1188) );
  CIVX2 U4746 ( .A(n1188), .Z(n4312) );
  CND2X1 U4747 ( .A(n1161), .B(n3603), .Z(n4414) );
  CIVX4 U4748 ( .A(n4124), .Z(n4509) );
  CEO3X1 U4749 ( .A(n1129), .B(n1125), .C(n1123), .Z(n1117) );
  CND2XL U4750 ( .A(n1129), .B(n1125), .Z(n4046) );
  CND2XL U4751 ( .A(n1129), .B(n1123), .Z(n4047) );
  CND2XL U4752 ( .A(n1125), .B(n1123), .Z(n4048) );
  CND3X1 U4753 ( .A(n4046), .B(n4047), .C(n4048), .Z(n1116) );
  CND2XL U4754 ( .A(n1095), .B(n1097), .Z(n4049) );
  CND2X1 U4755 ( .A(n1097), .B(n1116), .Z(n4050) );
  CND2XL U4756 ( .A(n1095), .B(n1116), .Z(n4051) );
  CND3X1 U4757 ( .A(n4049), .B(n4050), .C(n4051), .Z(n1088) );
  CND2X4 U4758 ( .A(n4374), .B(n4375), .Z(n4377) );
  CND2X1 U4759 ( .A(n699), .B(n691), .Z(n4373) );
  CND2X2 U4760 ( .A(n1088), .B(n1086), .Z(n4052) );
  CND2X1 U4761 ( .A(n1088), .B(n1065), .Z(n4053) );
  CND3X2 U4762 ( .A(n4052), .B(n4053), .C(n4054), .Z(n1060) );
  CND2XL U4763 ( .A(n1063), .B(n1084), .Z(n4055) );
  CND2XL U4764 ( .A(n1061), .B(n1063), .Z(n4056) );
  CND2XL U4765 ( .A(n1084), .B(n1061), .Z(n4057) );
  CND3X1 U4766 ( .A(n4055), .B(n4056), .C(n4057), .Z(n1058) );
  CND3X2 U4767 ( .A(n4087), .B(n4088), .C(n4089), .Z(n1152) );
  CND2X1 U4768 ( .A(n4026), .B(n2003), .Z(n4088) );
  CANR1X1 U4769 ( .A(n283), .B(n356), .C(n286), .Z(n282) );
  CND2X2 U4770 ( .A(n1091), .B(n1114), .Z(n4295) );
  CNR2X1 U4771 ( .A(n1581), .B(n1596), .Z(n643) );
  CENXL U4772 ( .A(n3908), .B(n4563), .Z(n4059) );
  CND2X4 U4773 ( .A(n2815), .B(net16433), .Z(net18628) );
  CENXL U4774 ( .A(net16541), .B(n4561), .Z(n2688) );
  CENXL U4775 ( .A(net16541), .B(n4557), .Z(n2692) );
  CENXL U4776 ( .A(net16541), .B(n4558), .Z(n2691) );
  CENXL U4777 ( .A(net16541), .B(n4556), .Z(n2693) );
  CENX1 U4778 ( .A(net16541), .B(n4555), .Z(n2694) );
  CND2X1 U4779 ( .A(n1908), .B(n1130), .Z(n4060) );
  CND2XL U4780 ( .A(n1908), .B(n2092), .Z(n4061) );
  CND2XL U4781 ( .A(n1130), .B(n2092), .Z(n4062) );
  CND3X1 U4782 ( .A(n4060), .B(n4061), .C(n4062), .Z(n1104) );
  CND2X4 U4783 ( .A(n96), .B(n3903), .Z(net18627) );
  CENX2 U4784 ( .A(a[0]), .B(n3678), .Z(n2827) );
  CENX1 U4785 ( .A(n4037), .B(n4564), .Z(n2616) );
  CND2X4 U4786 ( .A(n3328), .B(n2823), .Z(n4063) );
  CND2X4 U4787 ( .A(net16419), .B(n3309), .Z(n4064) );
  CIVXL U4788 ( .A(net18180), .Z(n574) );
  CEO3X2 U4789 ( .A(n1801), .B(n1887), .C(n2163), .Z(n1385) );
  CND2XL U4790 ( .A(n1801), .B(n1887), .Z(n4066) );
  CND2XL U4791 ( .A(n1801), .B(n2163), .Z(n4067) );
  CND2XL U4792 ( .A(n1887), .B(n2163), .Z(n4068) );
  CND3X1 U4793 ( .A(n4066), .B(n4067), .C(n4068), .Z(n1384) );
  CND2XL U4794 ( .A(n1404), .B(n1402), .Z(n4069) );
  CND2XL U4795 ( .A(n1404), .B(n1385), .Z(n4070) );
  CND2XL U4796 ( .A(n1402), .B(n1385), .Z(n4071) );
  CND3X1 U4797 ( .A(n4069), .B(n4070), .C(n4071), .Z(n1372) );
  CENXL U4798 ( .A(net15912), .B(n4543), .Z(n2409) );
  CENXL U4799 ( .A(net15912), .B(n4542), .Z(n2410) );
  CENXL U4800 ( .A(net15912), .B(n4548), .Z(n2404) );
  CENXL U4801 ( .A(n4547), .B(net15912), .Z(n2405) );
  CENXL U4802 ( .A(net15912), .B(n4565), .Z(n2384) );
  CND3X1 U4803 ( .A(net18592), .B(net18593), .C(n4072), .Z(n1156) );
  CND2X1 U4804 ( .A(net18496), .B(n4096), .Z(n2125) );
  CIVXL U4805 ( .A(n762), .Z(n4073) );
  CND2X1 U4806 ( .A(n4488), .B(n4489), .Z(n678) );
  CND2X1 U4807 ( .A(n1539), .B(n1537), .Z(n4286) );
  CIVXL U4808 ( .A(n356), .Z(n4074) );
  CENX2 U4809 ( .A(n168), .B(n435), .Z(product[44]) );
  COND1X2 U4810 ( .A(n3422), .B(net16471), .C(n441), .Z(n435) );
  CANR1X2 U4811 ( .A(n432), .B(n3257), .C(n3752), .Z(n417) );
  CND2X1 U4812 ( .A(n4238), .B(n1110), .Z(n4076) );
  CND2X2 U4813 ( .A(n4077), .B(n4076), .Z(n1085) );
  CND2X1 U4814 ( .A(n1442), .B(n1440), .Z(n4080) );
  CND2XL U4815 ( .A(n3174), .B(n1417), .Z(n4082) );
  CND2XL U4816 ( .A(n1417), .B(n1415), .Z(n4083) );
  CND2XL U4817 ( .A(n3173), .B(n1415), .Z(n4084) );
  CND3X1 U4818 ( .A(n4084), .B(n4083), .C(n4082), .Z(n1412) );
  CNIVX4 U4819 ( .A(n4588), .Z(n4085) );
  CND2XL U4820 ( .A(n4026), .B(n2063), .Z(n4087) );
  CND2X1 U4821 ( .A(n2063), .B(n2003), .Z(n4089) );
  CND2XL U4822 ( .A(n1148), .B(n1152), .Z(n4090) );
  CND3X1 U4823 ( .A(net18532), .B(n4090), .C(net18534), .Z(n1118) );
  COR2XL U4824 ( .A(n3121), .B(n2525), .Z(n4092) );
  CIVXL U4825 ( .A(n1130), .Z(n1131) );
  COND2X1 U4826 ( .A(n3301), .B(n2401), .C(n2400), .D(net17425), .Z(n1130) );
  CENXL U4827 ( .A(net15974), .B(n4557), .Z(n2659) );
  CENXL U4828 ( .A(n3908), .B(n4544), .Z(n2672) );
  CENXL U4829 ( .A(n3908), .B(n4563), .Z(n2652) );
  COND2XL U4830 ( .A(n4012), .B(n2387), .C(n2386), .D(net16426), .Z(n864) );
  COND2XL U4831 ( .A(n4012), .B(n2392), .C(n2391), .D(net17425), .Z(n1872) );
  CIVX2 U4832 ( .A(n470), .Z(n4449) );
  CND2IX2 U4833 ( .B(n4257), .A(n4216), .Z(n2096) );
  CND3X1 U4834 ( .A(n4384), .B(n4385), .C(n4386), .Z(n1132) );
  CANR1X1 U4835 ( .A(n3759), .B(n260), .C(n253), .Z(n249) );
  CEOX2 U4836 ( .A(n200), .B(n684), .Z(product[12]) );
  CANR1X1 U4837 ( .A(n4489), .B(n689), .C(n686), .Z(n684) );
  CNR2IX1 U4838 ( .B(n3244), .A(n3644), .Z(n2155) );
  CND2XL U4839 ( .A(n2166), .B(n1983), .Z(n4241) );
  CND2X4 U4840 ( .A(n4421), .B(n4422), .Z(n4424) );
  CENXL U4841 ( .A(n3909), .B(n4555), .Z(n2661) );
  COND2XL U4842 ( .A(net16309), .B(n2677), .C(n3644), .D(n2676), .Z(n2152) );
  CIVX2 U4843 ( .A(n4589), .Z(n4398) );
  CAOR1XL U4844 ( .A(n3122), .B(net17279), .C(n2516), .Z(n1993) );
  CND2XL U4845 ( .A(n1256), .B(n1231), .Z(n4425) );
  CND2XL U4846 ( .A(n1249), .B(n1276), .Z(n4099) );
  CND3X1 U4847 ( .A(n4097), .B(n4098), .C(n4099), .Z(n1244) );
  CND2XL U4848 ( .A(n1297), .B(n1301), .Z(n4102) );
  CND3X2 U4849 ( .A(n4100), .B(n4101), .C(n4102), .Z(n1284) );
  CND2XL U4850 ( .A(n1287), .B(n1314), .Z(n4539) );
  CND2XL U4851 ( .A(n1546), .B(n1527), .Z(n4103) );
  CND2XL U4852 ( .A(n1527), .B(n1529), .Z(n4104) );
  CND2XL U4853 ( .A(n1546), .B(n1529), .Z(n4105) );
  CNIVX4 U4854 ( .A(n2797), .Z(n4551) );
  CEOX1 U4855 ( .A(n2110), .B(n2141), .Z(n4106) );
  CEOX1 U4856 ( .A(n4106), .B(n1578), .Z(n1555) );
  CND2X1 U4857 ( .A(n2141), .B(n2110), .Z(n4109) );
  CEOX2 U4858 ( .A(n4188), .B(n1554), .Z(n1533) );
  CEO3X2 U4859 ( .A(n1207), .B(n1205), .C(n1213), .Z(n1199) );
  CND2X1 U4860 ( .A(n1207), .B(n1213), .Z(n4111) );
  CND2X1 U4861 ( .A(n1205), .B(n1213), .Z(n4112) );
  CND2XL U4862 ( .A(n1224), .B(n1199), .Z(n4115) );
  CEOX2 U4863 ( .A(n2228), .B(n2197), .Z(n4116) );
  CEOX2 U4864 ( .A(n4116), .B(n1984), .Z(n1477) );
  CND2X1 U4865 ( .A(n1984), .B(n2197), .Z(n4117) );
  CND2X4 U4866 ( .A(n2819), .B(n3789), .Z(n4120) );
  CND2X1 U4867 ( .A(n1537), .B(n1541), .Z(n4288) );
  CIVXL U4868 ( .A(n495), .Z(n4122) );
  CANR1X1 U4869 ( .A(n631), .B(n3512), .C(n3990), .Z(n4123) );
  CND2X1 U4870 ( .A(n3782), .B(n3986), .Z(n4253) );
  CNR2IXL U4871 ( .B(n3750), .A(net17297), .Z(n2187) );
  CND2X2 U4872 ( .A(n3709), .B(n4424), .Z(n4124) );
  CND2X1 U4873 ( .A(n1269), .B(n1263), .Z(n4126) );
  CND2X1 U4874 ( .A(n1290), .B(n1263), .Z(n4127) );
  CND3X2 U4875 ( .A(n4125), .B(n4126), .C(n4127), .Z(n1254) );
  CND2XL U4876 ( .A(n1229), .B(n1227), .Z(n4128) );
  CND2XL U4877 ( .A(n1229), .B(n1254), .Z(n4129) );
  CND2XL U4878 ( .A(n1227), .B(n1254), .Z(n4130) );
  CIVX1 U4879 ( .A(n4570), .Z(n4435) );
  CEO3X2 U4880 ( .A(n1446), .B(n1448), .C(n3294), .Z(n1419) );
  COND2X1 U4881 ( .A(n3302), .B(n2389), .C(n2388), .D(net16426), .Z(n890) );
  CENXL U4882 ( .A(n3828), .B(n4563), .Z(n2388) );
  CND2X1 U4883 ( .A(n1197), .B(n1222), .Z(n4132) );
  CND2X1 U4884 ( .A(n1195), .B(n1222), .Z(n4133) );
  CND3X2 U4885 ( .A(n4133), .B(n4132), .C(n4131), .Z(n1190) );
  CND2XL U4886 ( .A(n1165), .B(n1192), .Z(n4134) );
  COND2X1 U4887 ( .A(n3210), .B(n2755), .C(n6), .D(n2754), .Z(n2228) );
  CND2X2 U4888 ( .A(n767), .B(n768), .Z(n4155) );
  CEO3X2 U4889 ( .A(n1410), .B(n1406), .C(n1408), .Z(n1375) );
  CND2X1 U4890 ( .A(n1410), .B(n1406), .Z(n4137) );
  CND2X1 U4891 ( .A(n1410), .B(n1408), .Z(n4138) );
  CND2X1 U4892 ( .A(n1406), .B(n1408), .Z(n4139) );
  CND3X1 U4893 ( .A(n4137), .B(n4138), .C(n4139), .Z(n1374) );
  CND2X1 U4894 ( .A(n1373), .B(n1396), .Z(n4140) );
  CND2X1 U4895 ( .A(n1373), .B(n1375), .Z(n4141) );
  CND2X1 U4896 ( .A(n1396), .B(n1375), .Z(n4142) );
  CND3X2 U4897 ( .A(n4140), .B(n4141), .C(n4142), .Z(n1366) );
  CHA1X1 U4898 ( .A(n2172), .B(n1730), .CO(n1578), .S(n1579) );
  COND2XL U4899 ( .A(n4511), .B(n2256), .C(n2255), .D(n3277), .Z(n1742) );
  COND2XL U4900 ( .A(n4511), .B(n2254), .C(n2253), .D(n3277), .Z(n1741) );
  COND2XL U4901 ( .A(n4511), .B(n2255), .C(n2254), .D(n3277), .Z(n800) );
  COND2XL U4902 ( .A(n4511), .B(n2257), .C(n2256), .D(n3277), .Z(n810) );
  COND2XL U4903 ( .A(n4511), .B(n2258), .C(n2257), .D(n3277), .Z(n1743) );
  COND2XL U4904 ( .A(n4511), .B(n2259), .C(n2258), .D(n3277), .Z(n824) );
  COND2XL U4905 ( .A(n4511), .B(n2262), .C(n2261), .D(n3277), .Z(n1746) );
  CNIVXL U4906 ( .A(n1575), .Z(n4143) );
  CND2X1 U4907 ( .A(n1048), .B(n1027), .Z(n4144) );
  CND3X2 U4908 ( .A(n4144), .B(n4145), .C(n4146), .Z(n1020) );
  CND2XL U4909 ( .A(n1042), .B(n1040), .Z(n4147) );
  CND2X1 U4910 ( .A(n1042), .B(n1021), .Z(n4148) );
  CND2XL U4911 ( .A(n1040), .B(n1021), .Z(n4149) );
  CND3X1 U4912 ( .A(n4147), .B(n4148), .C(n4149), .Z(n1016) );
  CND2XL U4913 ( .A(n1413), .B(n1436), .Z(n4150) );
  CND2X2 U4914 ( .A(n4374), .B(n4375), .Z(n4152) );
  CEOX2 U4915 ( .A(n4404), .B(n1409), .Z(n1397) );
  CNR2X2 U4916 ( .A(n572), .B(n567), .Z(n561) );
  CANR1X2 U4917 ( .A(n620), .B(n629), .C(n4315), .Z(n619) );
  CENXL U4918 ( .A(n3815), .B(n4547), .Z(n2570) );
  CENXL U4919 ( .A(n4121), .B(n4540), .Z(n2579) );
  CENXL U4920 ( .A(n4542), .B(n4121), .Z(n2575) );
  CENXL U4921 ( .A(n4121), .B(n4553), .Z(n2564) );
  CENXL U4922 ( .A(n4121), .B(n4545), .Z(n2572) );
  CENXL U4923 ( .A(n4121), .B(n4543), .Z(n2574) );
  CENXL U4924 ( .A(n4568), .B(n3622), .Z(n2576) );
  COND2XL U4925 ( .A(n3301), .B(n2386), .C(n2385), .D(net16426), .Z(n1869) );
  CND2XL U4926 ( .A(n1306), .B(n3249), .Z(n4383) );
  CND2XL U4927 ( .A(n1307), .B(n1309), .Z(n4255) );
  CENX1 U4928 ( .A(n4595), .B(n4550), .Z(n2369) );
  CENX1 U4929 ( .A(n4595), .B(n4552), .Z(n2367) );
  CANR1X1 U4930 ( .A(n272), .B(n356), .C(n273), .Z(n269) );
  CEO3X2 U4931 ( .A(n1374), .B(n1372), .C(n1349), .Z(n1341) );
  CND2XL U4932 ( .A(n1374), .B(n1372), .Z(n4156) );
  CND2XL U4933 ( .A(n1374), .B(n1349), .Z(n4157) );
  CND2X1 U4934 ( .A(n1315), .B(n1340), .Z(n4160) );
  CND3X2 U4935 ( .A(n4159), .B(n4160), .C(n4161), .Z(n1308) );
  CND2X4 U4936 ( .A(n2813), .B(net16437), .Z(net18310) );
  CENXL U4937 ( .A(n3833), .B(n4550), .Z(n2435) );
  CENXL U4938 ( .A(n4568), .B(n3078), .Z(n2444) );
  CND2IXL U4939 ( .B(n3750), .A(net16541), .Z(n2713) );
  CENXL U4940 ( .A(n3244), .B(net16541), .Z(n2712) );
  CND2XL U4941 ( .A(n1257), .B(n1284), .Z(n4248) );
  CNIVX4 U4942 ( .A(n2793), .Z(n4555) );
  CEOX2 U4943 ( .A(n4165), .B(n977), .Z(n975) );
  CND2XL U4944 ( .A(n977), .B(n996), .Z(n4166) );
  CND2XL U4945 ( .A(n996), .B(n979), .Z(n4168) );
  CND3XL U4946 ( .A(n4166), .B(n4167), .C(n4168), .Z(n974) );
  CND2X1 U4947 ( .A(n957), .B(n974), .Z(n434) );
  CNR2X1 U4948 ( .A(n975), .B(n994), .Z(n448) );
  CND2X1 U4949 ( .A(n1335), .B(n1337), .Z(n4171) );
  CND2XL U4950 ( .A(n2195), .B(n1951), .Z(n4173) );
  CND2XL U4951 ( .A(n2195), .B(n1982), .Z(n4174) );
  CND3X1 U4952 ( .A(n4173), .B(n4174), .C(n4175), .Z(n1430) );
  CND2X1 U4953 ( .A(n387), .B(n418), .Z(n385) );
  CNR2IX1 U4954 ( .B(n396), .A(n389), .Z(n387) );
  CND2XL U4955 ( .A(n2050), .B(n2021), .Z(n4176) );
  CND2XL U4956 ( .A(n2050), .B(n1990), .Z(n4177) );
  CND2XL U4957 ( .A(n1606), .B(n1595), .Z(n4179) );
  CND2XL U4958 ( .A(n1606), .B(n1593), .Z(n4180) );
  CND2XL U4959 ( .A(n1595), .B(n1593), .Z(n4181) );
  CND3X1 U4960 ( .A(n4179), .B(n4180), .C(n4181), .Z(n1586) );
  CIVXL U4961 ( .A(n66), .Z(n4182) );
  CIVX2 U4962 ( .A(n66), .Z(n4584) );
  CNIVX4 U4963 ( .A(n2807), .Z(n4568) );
  CND2X1 U4964 ( .A(n1425), .B(n1448), .Z(n4187) );
  CNIVX4 U4965 ( .A(n2794), .Z(n4554) );
  CNIVX4 U4966 ( .A(n2788), .Z(n4560) );
  CEOX2 U4967 ( .A(n1558), .B(n1556), .Z(n4188) );
  CND2X1 U4968 ( .A(n1554), .B(n1556), .Z(n4189) );
  CND2X1 U4969 ( .A(n1554), .B(n1558), .Z(n4190) );
  CND3X2 U4970 ( .A(n4189), .B(n4190), .C(n4191), .Z(n1532) );
  CND3X2 U4971 ( .A(n4306), .B(n4307), .C(n4308), .Z(n1558) );
  COND2XL U4972 ( .A(net18772), .B(n2698), .C(net16451), .D(n2697), .Z(n2172)
         );
  CND2X1 U4973 ( .A(n1470), .B(n1472), .Z(n4193) );
  CND3X2 U4974 ( .A(n4192), .B(n4193), .C(n4194), .Z(n1442) );
  CND2XL U4975 ( .A(n1464), .B(n1466), .Z(n4195) );
  CND3X2 U4976 ( .A(n4335), .B(n4336), .C(n4337), .Z(n1312) );
  CND2X1 U4977 ( .A(n1346), .B(n1321), .Z(n4335) );
  CND2X1 U4978 ( .A(n1346), .B(n1344), .Z(n4336) );
  CND2X1 U4979 ( .A(n4198), .B(net15914), .Z(n4200) );
  CND2X1 U4980 ( .A(n1641), .B(n1652), .Z(n672) );
  COND2X1 U4981 ( .A(n4013), .B(n2408), .C(n2407), .D(net17425), .Z(n1885) );
  CND3X1 U4982 ( .A(n4296), .B(n4297), .C(n4298), .Z(n1468) );
  CIVX2 U4983 ( .A(n1089), .Z(net18199) );
  CENXL U4984 ( .A(n3893), .B(n4554), .Z(n2596) );
  CENX1 U4985 ( .A(n1638), .B(n1636), .Z(n4234) );
  COND2X1 U4986 ( .A(n4461), .B(n2733), .C(n2732), .D(n4510), .Z(n2206) );
  CEO3X1 U4987 ( .A(n1295), .B(n1293), .C(n1299), .Z(n1287) );
  CND2XL U4988 ( .A(n1135), .B(n3487), .Z(n4384) );
  CIVXL U4989 ( .A(n84), .Z(n4202) );
  CENX2 U4990 ( .A(n1256), .B(n4203), .Z(n1223) );
  CEOX2 U4991 ( .A(n189), .B(n619), .Z(product[23]) );
  CNR2IX1 U4992 ( .B(n3244), .A(net18914), .Z(n2122) );
  CIVX2 U4993 ( .A(n84), .Z(n4590) );
  CNIVX4 U4994 ( .A(n18), .Z(n4460) );
  CND2XL U4995 ( .A(n1452), .B(n1456), .Z(n4204) );
  CND2XL U4996 ( .A(n1452), .B(n1450), .Z(n4205) );
  CND2XL U4997 ( .A(n1456), .B(n1450), .Z(n4206) );
  CND3X1 U4998 ( .A(n4204), .B(n4205), .C(n4206), .Z(n1424) );
  CANR1XL U4999 ( .A(n3177), .B(n612), .C(n3875), .Z(net18180) );
  CANR1X1 U5000 ( .A(n576), .B(n612), .C(n577), .Z(n575) );
  CENXL U5001 ( .A(net18828), .B(n4543), .Z(n2706) );
  CENXL U5002 ( .A(net18828), .B(n4565), .Z(n2681) );
  CND2X1 U5003 ( .A(n661), .B(n778), .Z(n196) );
  CND2X1 U5004 ( .A(n1613), .B(n1626), .Z(n661) );
  CND2X2 U5005 ( .A(n3454), .B(n4312), .Z(n4313) );
  CIVXL U5006 ( .A(n3026), .Z(n4208) );
  CND2X1 U5007 ( .A(n1483), .B(n1504), .Z(n618) );
  CNIVX4 U5008 ( .A(n2800), .Z(n4548) );
  CEO3X2 U5009 ( .A(n1101), .B(n1120), .C(n1118), .Z(n1091) );
  CND2XL U5010 ( .A(n1120), .B(n1118), .Z(n4209) );
  CND2XL U5011 ( .A(n1120), .B(n1101), .Z(n4210) );
  CND2X1 U5012 ( .A(n1118), .B(n1101), .Z(n4211) );
  CND3X1 U5013 ( .A(n4209), .B(n4210), .C(n4211), .Z(n1090) );
  CND2X1 U5014 ( .A(n4476), .B(n1189), .Z(n4214) );
  CND2X2 U5015 ( .A(n4212), .B(n4213), .Z(n4215) );
  CND2X2 U5016 ( .A(n4215), .B(n4214), .Z(n1187) );
  CNR2X2 U5017 ( .A(n1214), .B(n1187), .Z(n529) );
  CND2X2 U5018 ( .A(n1187), .B(n1214), .Z(n530) );
  CIVXL U5019 ( .A(n573), .Z(n571) );
  CND2IX1 U5020 ( .B(n1163), .A(n1188), .Z(n4314) );
  COND2X1 U5021 ( .A(n99), .B(n2435), .C(net16416), .D(n2434), .Z(n1912) );
  CND2X4 U5022 ( .A(n4376), .B(n4152), .Z(n4217) );
  CND2X1 U5023 ( .A(n1216), .B(n1189), .Z(n4521) );
  COND1XL U5024 ( .A(n224), .B(n3732), .C(n225), .Z(n223) );
  CAOR1XL U5025 ( .A(n3277), .B(n4511), .C(n2252), .Z(n1740) );
  COND2XL U5026 ( .A(n4511), .B(n2253), .C(n2252), .D(n3277), .Z(n794) );
  CENX1 U5027 ( .A(n4582), .B(n4560), .Z(n2524) );
  CNR2X2 U5028 ( .A(n1275), .B(n1304), .Z(n551) );
  CENXL U5029 ( .A(n506), .B(n175), .Z(product[37]) );
  CENXL U5030 ( .A(n4570), .B(n4560), .Z(n2755) );
  CND2IXL U5031 ( .B(n3244), .A(n4600), .Z(n2317) );
  CIVXL U5032 ( .A(n646), .Z(n4218) );
  CND2XL U5033 ( .A(n1865), .B(n2042), .Z(n4220) );
  CND2XL U5034 ( .A(n1920), .B(n1865), .Z(n4221) );
  CND2XL U5035 ( .A(n2042), .B(n1920), .Z(n4222) );
  CND3X1 U5036 ( .A(n4220), .B(n4221), .C(n4222), .Z(n1432) );
  CIVXL U5037 ( .A(n1865), .Z(n4223) );
  CIVX1 U5038 ( .A(n4223), .Z(n4224) );
  COND2XL U5039 ( .A(net18628), .B(n2381), .C(net16433), .D(n2380), .Z(n1865)
         );
  CIVXL U5040 ( .A(n3790), .Z(n4225) );
  COND2X1 U5041 ( .A(net16309), .B(n2666), .C(n3644), .D(n2665), .Z(n2141) );
  CENXL U5042 ( .A(n3893), .B(n4547), .Z(n2603) );
  CENXL U5043 ( .A(n3893), .B(n4546), .Z(n2604) );
  CENXL U5044 ( .A(n3893), .B(n4555), .Z(n2595) );
  CENXL U5045 ( .A(n3753), .B(n4550), .Z(n2600) );
  CND2X1 U5046 ( .A(n1329), .B(n1331), .Z(n4227) );
  CND2XL U5047 ( .A(n1323), .B(n1329), .Z(n4228) );
  CND2XL U5048 ( .A(n1323), .B(n1331), .Z(n4229) );
  CND3X1 U5049 ( .A(n4227), .B(n4228), .C(n4229), .Z(n1316) );
  CND2X1 U5050 ( .A(n1345), .B(n1347), .Z(n4230) );
  CND2X1 U5051 ( .A(n1345), .B(n1370), .Z(n4231) );
  CND2X1 U5052 ( .A(n1347), .B(n1370), .Z(n4232) );
  CND3X2 U5053 ( .A(n4230), .B(n4231), .C(n4232), .Z(n1338) );
  CNIVX4 U5054 ( .A(n2801), .Z(n4547) );
  CNIVX4 U5055 ( .A(n2786), .Z(n4562) );
  CNIVX4 U5056 ( .A(n2795), .Z(n4553) );
  CENXL U5057 ( .A(n3026), .B(n4548), .Z(n2470) );
  CENXL U5058 ( .A(n4085), .B(n4541), .Z(n2478) );
  CENXL U5059 ( .A(n4085), .B(n4565), .Z(n2450) );
  CENXL U5060 ( .A(n4086), .B(n4547), .Z(n2471) );
  CIVXL U5061 ( .A(n222), .Z(n220) );
  CNIVX4 U5062 ( .A(n2790), .Z(n4558) );
  COND2X1 U5063 ( .A(n4063), .B(n2622), .C(net16420), .D(n2621), .Z(n2097) );
  CND2XL U5064 ( .A(n1306), .B(n1277), .Z(n4381) );
  CENXL U5065 ( .A(n4592), .B(n4546), .Z(n2439) );
  CENXL U5066 ( .A(n4592), .B(n4555), .Z(n2430) );
  CENXL U5067 ( .A(n4592), .B(n4545), .Z(n2440) );
  CENXL U5068 ( .A(n4592), .B(n2809), .Z(n2446) );
  CENXL U5069 ( .A(n4592), .B(n4549), .Z(n2436) );
  CND2X1 U5070 ( .A(n1528), .B(n4065), .Z(n4236) );
  CND2XL U5071 ( .A(n1511), .B(n4065), .Z(n4237) );
  CNIVX4 U5072 ( .A(n2784), .Z(n4563) );
  CIVXL U5073 ( .A(net18400), .Z(net18061) );
  CND2XL U5074 ( .A(n2227), .B(n2166), .Z(n4239) );
  CND2XL U5075 ( .A(n2227), .B(n1983), .Z(n4240) );
  CND3X1 U5076 ( .A(n4239), .B(n4240), .C(n4241), .Z(n1456) );
  CND3X2 U5077 ( .A(n4521), .B(n4522), .C(n4523), .Z(n1186) );
  CIVX4 U5078 ( .A(a[16]), .Z(n4375) );
  CND2X1 U5079 ( .A(n1317), .B(n1319), .Z(n4243) );
  CND2X1 U5080 ( .A(n1317), .B(n1342), .Z(n4244) );
  CND2X1 U5081 ( .A(n1319), .B(n1342), .Z(n4245) );
  CND3X2 U5082 ( .A(n4243), .B(n4244), .C(n4245), .Z(n1310) );
  CND2X2 U5083 ( .A(n4246), .B(n4247), .Z(n2191) );
  CENXL U5084 ( .A(n4512), .B(n4563), .Z(n2718) );
  CENXL U5085 ( .A(n4572), .B(net16104), .Z(n2717) );
  CNR2IX1 U5086 ( .B(n3750), .A(n3277), .Z(n1768) );
  CND2X1 U5087 ( .A(n1257), .B(n1286), .Z(n4249) );
  CND2XL U5088 ( .A(n1284), .B(n1286), .Z(n4250) );
  CNIVX4 U5089 ( .A(n2796), .Z(n4552) );
  CIVX2 U5090 ( .A(net15916), .Z(net15914) );
  COND1X1 U5091 ( .A(n4155), .B(n595), .C(n579), .Z(n577) );
  CND2XL U5092 ( .A(n1307), .B(n1334), .Z(n4254) );
  CND2XL U5093 ( .A(n1334), .B(n1309), .Z(n4256) );
  CND3X1 U5094 ( .A(n4254), .B(n4255), .C(n4256), .Z(n1304) );
  CNIVX8 U5095 ( .A(n2799), .Z(n4549) );
  CENXL U5096 ( .A(n635), .B(n192), .Z(product[20]) );
  CNIVX4 U5097 ( .A(n2798), .Z(n4550) );
  CENX1 U5098 ( .A(n4037), .B(n4562), .Z(n2621) );
  CENXL U5099 ( .A(n4037), .B(n2785), .Z(n2620) );
  CEO3X1 U5100 ( .A(n2049), .B(n2020), .C(n2233), .Z(n1575) );
  CND2XL U5101 ( .A(n3613), .B(n2020), .Z(n4258) );
  CND2XL U5102 ( .A(n3613), .B(n2233), .Z(n4259) );
  CND2X1 U5103 ( .A(n2020), .B(n2233), .Z(n4260) );
  CND2XL U5104 ( .A(n1590), .B(n1577), .Z(n4261) );
  CND2XL U5105 ( .A(n1590), .B(n1575), .Z(n4262) );
  CND2XL U5106 ( .A(n1577), .B(n1575), .Z(n4263) );
  COR2XL U5107 ( .A(n6), .B(n2759), .Z(n4265) );
  CND2X2 U5108 ( .A(n4264), .B(n4265), .Z(n2233) );
  CENXL U5109 ( .A(n4570), .B(n4555), .Z(n2760) );
  CENXL U5110 ( .A(n4570), .B(n4556), .Z(n2759) );
  CND2IXL U5111 ( .B(n3750), .A(n4579), .Z(n2614) );
  CENXL U5112 ( .A(n3893), .B(n4565), .Z(n2582) );
  CENXL U5113 ( .A(n3893), .B(n4545), .Z(n2605) );
  CENXL U5114 ( .A(n3893), .B(n4541), .Z(n2610) );
  CENXL U5115 ( .A(n3893), .B(n4552), .Z(n2598) );
  CENXL U5116 ( .A(n4121), .B(n4550), .Z(n2567) );
  CENXL U5117 ( .A(n3244), .B(n3790), .Z(n2580) );
  CENXL U5118 ( .A(n4592), .B(n4543), .Z(n2442) );
  CENXL U5119 ( .A(n4592), .B(n4542), .Z(n2443) );
  CENXL U5120 ( .A(n4591), .B(n4544), .Z(n2441) );
  CENXL U5121 ( .A(n4591), .B(n4561), .Z(n2424) );
  CENXL U5122 ( .A(n4591), .B(n4562), .Z(n2423) );
  CENXL U5123 ( .A(n4591), .B(net16102), .Z(n2419) );
  CENXL U5124 ( .A(n4591), .B(n2785), .Z(n2422) );
  CEO3XL U5125 ( .A(n1992), .B(n2205), .C(n2052), .Z(n1625) );
  CND2X1 U5126 ( .A(n4289), .B(n770), .Z(n594) );
  COND1X1 U5127 ( .A(n298), .B(net16472), .C(n299), .Z(n4267) );
  CND2XL U5128 ( .A(n738), .B(n296), .Z(n4268) );
  CNR2IX1 U5129 ( .B(n3244), .A(n123), .Z(n1834) );
  CIVX1 U5130 ( .A(n426), .Z(n4353) );
  CENXL U5131 ( .A(n4570), .B(n4562), .Z(n4270) );
  CENXL U5132 ( .A(n4570), .B(n4562), .Z(n2753) );
  CIVX8 U5133 ( .A(n3677), .Z(n4570) );
  CND2XL U5134 ( .A(n1289), .B(n1314), .Z(n4538) );
  CEO3X2 U5135 ( .A(n2162), .B(n1917), .C(n1800), .Z(n1353) );
  CND2X1 U5136 ( .A(n2162), .B(n1917), .Z(n4271) );
  CND2XL U5137 ( .A(n2162), .B(n1800), .Z(n4272) );
  CND2XL U5138 ( .A(n1917), .B(n1800), .Z(n4273) );
  CND3X1 U5139 ( .A(n4271), .B(n4272), .C(n4273), .Z(n1352) );
  CND2X1 U5140 ( .A(n1351), .B(n1353), .Z(n4275) );
  CND2X1 U5141 ( .A(n1357), .B(n1353), .Z(n4276) );
  CNR2XL U5142 ( .A(net16438), .B(n2315), .Z(n4278) );
  COR2X1 U5143 ( .A(n4277), .B(n4278), .Z(n1800) );
  CENXL U5144 ( .A(n4600), .B(n4540), .Z(n2315) );
  CEOX2 U5145 ( .A(n1164), .B(n1139), .Z(n4279) );
  CIVXL U5146 ( .A(n572), .Z(n766) );
  CNR2X4 U5147 ( .A(n4280), .B(n3907), .Z(net17930) );
  COND2X1 U5148 ( .A(n4013), .B(n2410), .C(n2409), .D(net17425), .Z(n1887) );
  CENXL U5149 ( .A(n4598), .B(n4554), .Z(n2332) );
  CENXL U5150 ( .A(n4598), .B(n4551), .Z(n2335) );
  CENXL U5151 ( .A(n4598), .B(n4550), .Z(n2336) );
  CIVXL U5152 ( .A(n4595), .Z(n4281) );
  CIVXL U5153 ( .A(n530), .Z(n528) );
  CIVXL U5154 ( .A(n622), .Z(n772) );
  CNR2X2 U5155 ( .A(n1613), .B(n1626), .Z(n660) );
  COND2X1 U5156 ( .A(n63), .B(n4225), .C(n2581), .D(n4505), .Z(n1733) );
  CENXL U5157 ( .A(n4592), .B(n4541), .Z(n2445) );
  CENXL U5158 ( .A(n4592), .B(n4540), .Z(n2447) );
  CNR2X1 U5159 ( .A(n1437), .B(n1460), .Z(n4282) );
  CND2X2 U5160 ( .A(n1525), .B(n1544), .Z(n628) );
  COAN1X1 U5161 ( .A(n606), .B(n4282), .C(n603), .Z(n595) );
  CND2X1 U5162 ( .A(n1310), .B(n1312), .Z(n4340) );
  CND2X1 U5163 ( .A(n1310), .B(n1285), .Z(n4338) );
  CIVXL U5164 ( .A(n4150), .Z(n590) );
  CENXL U5165 ( .A(n4582), .B(n4544), .Z(n2540) );
  CENXL U5166 ( .A(n4582), .B(n4558), .Z(n2526) );
  CENXL U5167 ( .A(n4582), .B(net16102), .Z(n2518) );
  CENXL U5168 ( .A(n4582), .B(n4563), .Z(n2520) );
  CENXL U5169 ( .A(n3078), .B(n4554), .Z(n2431) );
  CENXL U5170 ( .A(n3078), .B(n4552), .Z(n2433) );
  CENXL U5171 ( .A(n4589), .B(n4554), .Z(n2464) );
  CENXL U5172 ( .A(n4568), .B(n3026), .Z(n2477) );
  CENXL U5173 ( .A(n4550), .B(n4589), .Z(n2468) );
  CENXL U5174 ( .A(n4589), .B(n4551), .Z(n2467) );
  CENXL U5175 ( .A(n4589), .B(n4553), .Z(n2465) );
  CENXL U5176 ( .A(n4589), .B(n4552), .Z(n2466) );
  COND2X1 U5177 ( .A(net16309), .B(n2663), .C(net16490), .D(n2662), .Z(n2138)
         );
  CENXL U5178 ( .A(n4595), .B(n4561), .Z(n2358) );
  CENXL U5179 ( .A(n4595), .B(n4562), .Z(n2357) );
  CENXL U5180 ( .A(n4595), .B(n4559), .Z(n2360) );
  CENXL U5181 ( .A(n4595), .B(n4555), .Z(n2364) );
  CENXL U5182 ( .A(n4595), .B(n4558), .Z(n2361) );
  CENXL U5183 ( .A(n4595), .B(n4543), .Z(n2376) );
  CENXL U5184 ( .A(n4595), .B(n4557), .Z(n2362) );
  CENXL U5185 ( .A(n4595), .B(n2809), .Z(n2380) );
  COND1X2 U5186 ( .A(n471), .B(net16471), .C(n472), .Z(n470) );
  COND2X1 U5187 ( .A(n4013), .B(n2406), .C(n2405), .D(net17425), .Z(n1883) );
  CEO3X2 U5188 ( .A(n2170), .B(n2231), .C(n3979), .Z(n1541) );
  CND2XL U5189 ( .A(n2170), .B(n1987), .Z(n4283) );
  CND2X1 U5190 ( .A(n1987), .B(n2231), .Z(n4285) );
  CND2X1 U5191 ( .A(n1539), .B(n1541), .Z(n4287) );
  CIVXL U5192 ( .A(n543), .Z(n762) );
  CNR2IX1 U5193 ( .B(n3750), .A(net16426), .Z(n1893) );
  CAOR1XL U5194 ( .A(net17425), .B(net17728), .C(n2384), .Z(n1868) );
  COND2XL U5195 ( .A(n4012), .B(n2385), .C(n2384), .D(net17425), .Z(n842) );
  CENXL U5196 ( .A(n4592), .B(n4565), .Z(n2417) );
  COND2X1 U5197 ( .A(n3302), .B(n2405), .C(net17425), .D(n2404), .Z(n1882) );
  COR2XL U5198 ( .A(n1460), .B(n1437), .Z(n4289) );
  CND3X2 U5199 ( .A(n4290), .B(n4291), .C(n4292), .Z(n1114) );
  CND2X1 U5200 ( .A(n1093), .B(n1091), .Z(n4293) );
  CND2XL U5201 ( .A(n3360), .B(n1475), .Z(n4296) );
  CND2XL U5202 ( .A(n3360), .B(n1477), .Z(n4297) );
  CND2X1 U5203 ( .A(n1475), .B(n1477), .Z(n4298) );
  CND2X1 U5204 ( .A(n1445), .B(n1447), .Z(n4300) );
  CND2X1 U5205 ( .A(n1445), .B(n1468), .Z(n4301) );
  CND2X1 U5206 ( .A(n1447), .B(n1468), .Z(n4302) );
  CND3X2 U5207 ( .A(n4300), .B(n4301), .C(n4302), .Z(n1440) );
  COR2X1 U5208 ( .A(n4217), .B(n2506), .Z(n4304) );
  CND2X2 U5209 ( .A(n4303), .B(n4304), .Z(n1984) );
  CENXL U5210 ( .A(n4585), .B(n4544), .Z(n2507) );
  CENXL U5211 ( .A(n4585), .B(n4545), .Z(n2506) );
  CNR2X2 U5212 ( .A(n1685), .B(n1692), .Z(n693) );
  CIVX1 U5213 ( .A(n4561), .Z(n4358) );
  CIVXL U5214 ( .A(n567), .Z(n765) );
  CND2X1 U5215 ( .A(n1685), .B(n1692), .Z(n694) );
  CNIVX2 U5216 ( .A(n1988), .Z(n4309) );
  COND2XL U5217 ( .A(n4120), .B(n2511), .C(n4217), .D(n2510), .Z(n1988) );
  CENXL U5218 ( .A(n4577), .B(n4552), .Z(n2631) );
  CENXL U5219 ( .A(n4577), .B(n4551), .Z(n2632) );
  CENXL U5220 ( .A(n4568), .B(n4577), .Z(n2642) );
  CENXL U5221 ( .A(n4577), .B(n4550), .Z(n2633) );
  CENXL U5222 ( .A(n4577), .B(n4554), .Z(n2629) );
  CENXL U5223 ( .A(n4577), .B(n4553), .Z(n2630) );
  COND2X1 U5224 ( .A(n4461), .B(n2732), .C(n2731), .D(n4510), .Z(n2205) );
  CENXL U5225 ( .A(n3908), .B(n4556), .Z(n2660) );
  CND2X2 U5226 ( .A(n4313), .B(n4314), .Z(n4413) );
  COND2X1 U5227 ( .A(n3991), .B(n2480), .C(net16512), .D(n2479), .Z(n1957) );
  CENXL U5228 ( .A(n4568), .B(n3909), .Z(n2675) );
  CENXL U5229 ( .A(net15974), .B(n4551), .Z(n2665) );
  CENXL U5230 ( .A(n3909), .B(n4550), .Z(n2666) );
  CENXL U5231 ( .A(n3909), .B(n4553), .Z(n2663) );
  CIVXL U5232 ( .A(n4350), .Z(n4315) );
  CND2X4 U5233 ( .A(n2821), .B(n4504), .Z(n4316) );
  CNR2X2 U5234 ( .A(n4460), .B(n2715), .Z(n4464) );
  CND2XL U5235 ( .A(n4289), .B(n603), .Z(n187) );
  CND2X1 U5236 ( .A(n3143), .B(n1115), .Z(n4317) );
  CND3X2 U5237 ( .A(n4317), .B(net17756), .C(net17755), .Z(n1110) );
  COR2X1 U5238 ( .A(n2556), .B(n4505), .Z(n4320) );
  CND2X2 U5239 ( .A(n4319), .B(n4320), .Z(n2032) );
  CND2X1 U5240 ( .A(n4359), .B(n4360), .Z(n2556) );
  CENXL U5241 ( .A(net18828), .B(n4546), .Z(n2703) );
  CENXL U5242 ( .A(net18828), .B(n4547), .Z(n2702) );
  CENXL U5243 ( .A(net18828), .B(n4548), .Z(n2701) );
  CENXL U5244 ( .A(net18828), .B(n4549), .Z(n2700) );
  CENXL U5245 ( .A(net18828), .B(n4550), .Z(n2699) );
  CENXL U5246 ( .A(net18828), .B(n4545), .Z(n2704) );
  CENXL U5247 ( .A(net18828), .B(n4542), .Z(n2707) );
  CENXL U5248 ( .A(net18828), .B(n4540), .Z(n2711) );
  CENXL U5249 ( .A(n3747), .B(n4572), .Z(n2745) );
  CENXL U5250 ( .A(n3748), .B(n3909), .Z(n2679) );
  CENXL U5251 ( .A(n3747), .B(n3078), .Z(n2448) );
  CND2IXL U5252 ( .B(n3244), .A(n4572), .Z(n2746) );
  CENXL U5253 ( .A(n4568), .B(n4573), .Z(n2741) );
  CENXL U5254 ( .A(n2809), .B(n4512), .Z(n2743) );
  CENXL U5255 ( .A(n4572), .B(n4557), .Z(n2725) );
  CENXL U5256 ( .A(n4572), .B(n4561), .Z(n2721) );
  CIVXL U5257 ( .A(n666), .Z(n664) );
  COND2X1 U5258 ( .A(n3302), .B(net18209), .C(n2416), .D(net17425), .Z(n1728)
         );
  CENXL U5259 ( .A(n4595), .B(n4565), .Z(n2351) );
  CENXL U5260 ( .A(n4595), .B(net16104), .Z(n2354) );
  CENXL U5261 ( .A(n4595), .B(net16102), .Z(n2353) );
  CENXL U5262 ( .A(n4595), .B(n2785), .Z(n2356) );
  CENXL U5263 ( .A(n4595), .B(n4563), .Z(n2355) );
  CENXL U5264 ( .A(n4595), .B(n4560), .Z(n2359) );
  CENXL U5265 ( .A(n4595), .B(n4545), .Z(n2374) );
  CENXL U5266 ( .A(n4595), .B(n4542), .Z(n2377) );
  CENXL U5267 ( .A(n4595), .B(n4547), .Z(n2372) );
  CENXL U5268 ( .A(n4595), .B(n4546), .Z(n2373) );
  CENXL U5269 ( .A(n4595), .B(n4541), .Z(n2379) );
  CENXL U5270 ( .A(n4595), .B(n4540), .Z(n2381) );
  CENXL U5271 ( .A(n3908), .B(net16104), .Z(n2651) );
  CENXL U5272 ( .A(net15974), .B(n4558), .Z(n2658) );
  COND1X1 U5273 ( .A(n261), .B(n3732), .C(n262), .Z(n260) );
  CNIVX4 U5274 ( .A(n2810), .Z(n4540) );
  CENXL U5275 ( .A(n4540), .B(net15912), .Z(n2414) );
  CNIVX2 U5276 ( .A(n2809), .Z(n4567) );
  CEOX2 U5277 ( .A(n4413), .B(n1161), .Z(n1159) );
  CENX1 U5278 ( .A(n4579), .B(n4559), .Z(n2591) );
  CND2XL U5279 ( .A(n2064), .B(n2033), .Z(n4322) );
  CND2XL U5280 ( .A(n3939), .B(n2033), .Z(n4323) );
  CND2XL U5281 ( .A(n3939), .B(n2064), .Z(n4324) );
  CND3X1 U5282 ( .A(n4322), .B(n4323), .C(n4324), .Z(n1180) );
  COR2XL U5283 ( .A(n27), .B(n2709), .Z(n4326) );
  COR2X1 U5284 ( .A(net16451), .B(n2708), .Z(n4327) );
  CND2X2 U5285 ( .A(n4326), .B(n4327), .Z(n2183) );
  CENXL U5286 ( .A(net18828), .B(n4541), .Z(n2709) );
  CENXL U5287 ( .A(n4568), .B(net16541), .Z(n2708) );
  CND2XL U5288 ( .A(n4512), .B(n4544), .Z(n4330) );
  CIVXL U5289 ( .A(n4512), .Z(n4328) );
  CIVX1 U5290 ( .A(n4544), .Z(n4329) );
  COND2XL U5291 ( .A(n4461), .B(n2739), .C(n2738), .D(n4510), .Z(n2212) );
  COND2X1 U5292 ( .A(n4460), .B(n2738), .C(n2737), .D(n4510), .Z(n2211) );
  CND2X1 U5293 ( .A(n1321), .B(n1344), .Z(n4337) );
  CND3X2 U5294 ( .A(n4338), .B(n4340), .C(n4339), .Z(n1278) );
  COR2X1 U5295 ( .A(n710), .B(n708), .Z(n4341) );
  CND2X2 U5296 ( .A(n4341), .B(n709), .Z(n707) );
  CNR2X2 U5297 ( .A(n1713), .B(n1716), .Z(n708) );
  CND2X1 U5298 ( .A(n4600), .B(n2809), .Z(n4344) );
  CND2X2 U5299 ( .A(n4342), .B(n4343), .Z(n4345) );
  CND2X2 U5300 ( .A(n4344), .B(n4345), .Z(n2314) );
  CEOX2 U5301 ( .A(n4346), .B(n1481), .Z(n1471) );
  CND2X1 U5302 ( .A(n1481), .B(n1496), .Z(n4347) );
  CND2X1 U5303 ( .A(n1481), .B(n1498), .Z(n4348) );
  CND2XL U5304 ( .A(n1496), .B(n1498), .Z(n4349) );
  CND3X2 U5305 ( .A(n4347), .B(n4348), .C(n4349), .Z(n1470) );
  CIVX2 U5306 ( .A(n621), .Z(n4350) );
  CIVX2 U5307 ( .A(n4352), .Z(n1458) );
  CND2X1 U5308 ( .A(n1890), .B(n1727), .Z(n4352) );
  CND2X1 U5309 ( .A(n426), .B(n167), .Z(n4355) );
  CND2X2 U5310 ( .A(n4353), .B(n4354), .Z(n4356) );
  CND2X2 U5311 ( .A(n4356), .B(n4355), .Z(product[45]) );
  CIVX2 U5312 ( .A(n167), .Z(n4354) );
  CND2XL U5313 ( .A(n4580), .B(n4561), .Z(n4359) );
  CIVXL U5314 ( .A(n3815), .Z(n4357) );
  CEO3X1 U5315 ( .A(n2053), .B(n2084), .C(n2237), .Z(n1635) );
  CND2X1 U5316 ( .A(n2084), .B(n2237), .Z(n4363) );
  CND3X2 U5317 ( .A(n4361), .B(n4362), .C(n4363), .Z(n1634) );
  CND2XL U5318 ( .A(n1638), .B(n1636), .Z(n4364) );
  CND2XL U5319 ( .A(n1636), .B(n1634), .Z(n4366) );
  CND3X1 U5320 ( .A(n4364), .B(n4365), .C(n4366), .Z(n1618) );
  CND2XL U5321 ( .A(n1992), .B(n2052), .Z(n4367) );
  CND2XL U5322 ( .A(n1992), .B(n2205), .Z(n4368) );
  CND2XL U5323 ( .A(n2052), .B(n2205), .Z(n4369) );
  CND2X4 U5324 ( .A(n4371), .B(n4372), .Z(n4499) );
  CIVXL U5325 ( .A(n3027), .Z(n689) );
  CND2X2 U5326 ( .A(n4583), .B(a[16]), .Z(n4376) );
  CND2X4 U5327 ( .A(n4376), .B(n4377), .Z(net16413) );
  CND2X1 U5328 ( .A(n1217), .B(n1246), .Z(n4378) );
  CND2X1 U5329 ( .A(n1217), .B(n1219), .Z(n4379) );
  CND3X2 U5330 ( .A(n4378), .B(n4379), .C(n4380), .Z(n1214) );
  CND2XL U5331 ( .A(n3487), .B(n1137), .Z(n4386) );
  CEO3X2 U5332 ( .A(n1553), .B(n1566), .C(n1551), .Z(n1547) );
  CEOX2 U5333 ( .A(n4387), .B(n1547), .Z(n1545) );
  CND2X1 U5334 ( .A(n1553), .B(n1551), .Z(n4389) );
  CND2X1 U5335 ( .A(n1566), .B(n1551), .Z(n4390) );
  CND3X2 U5336 ( .A(n4388), .B(n4389), .C(n4390), .Z(n1546) );
  CND2XL U5337 ( .A(n1549), .B(n1547), .Z(n4392) );
  CND2XL U5338 ( .A(n1564), .B(n1547), .Z(n4393) );
  CND3X1 U5339 ( .A(n4391), .B(n4392), .C(n4393), .Z(n1544) );
  CND2XL U5340 ( .A(n1414), .B(n1391), .Z(n4396) );
  CND2X2 U5341 ( .A(n3099), .B(n4398), .Z(n4399) );
  CND2XL U5342 ( .A(n2024), .B(n2206), .Z(n4401) );
  CND2XL U5343 ( .A(n2024), .B(n2146), .Z(n4402) );
  CND2XL U5344 ( .A(n2206), .B(n2146), .Z(n4403) );
  CND3X1 U5345 ( .A(n4401), .B(n4402), .C(n4403), .Z(n1636) );
  CND2XL U5346 ( .A(n4583), .B(n4540), .Z(n4409) );
  CND2X1 U5347 ( .A(n3646), .B(n4408), .Z(n4410) );
  CND2X1 U5348 ( .A(n4409), .B(n4410), .Z(n2546) );
  CIVX1 U5349 ( .A(n4540), .Z(n4408) );
  CND2X1 U5350 ( .A(n1161), .B(n3114), .Z(n4415) );
  CIVXL U5351 ( .A(n4603), .Z(n4418) );
  CND2X2 U5352 ( .A(n4423), .B(n4424), .Z(n15) );
  CND2X2 U5353 ( .A(n15), .B(n2826), .Z(n18) );
  CND2XL U5354 ( .A(n1231), .B(n1258), .Z(n4427) );
  CND3X1 U5355 ( .A(n4425), .B(n4426), .C(n4427), .Z(n1222) );
  CND2X1 U5356 ( .A(n4474), .B(net17136), .Z(n4429) );
  CND2X2 U5357 ( .A(n4428), .B(net17512), .Z(n4430) );
  CND2X2 U5358 ( .A(n4429), .B(n4430), .Z(product[39]) );
  CIVX1 U5359 ( .A(n4474), .Z(n4428) );
  CIVX2 U5360 ( .A(net17136), .Z(net17512) );
  CND2X1 U5361 ( .A(n4432), .B(n183), .Z(n4433) );
  CND2XL U5362 ( .A(n4431), .B(n569), .Z(n4434) );
  CND2X2 U5363 ( .A(n4433), .B(n4434), .Z(product[29]) );
  CIVX2 U5364 ( .A(n183), .Z(n4431) );
  CIVXL U5365 ( .A(n569), .Z(n4432) );
  CND2X1 U5366 ( .A(n4570), .B(n4564), .Z(n4437) );
  CND2X2 U5367 ( .A(n4435), .B(n4436), .Z(n4438) );
  CND2X2 U5368 ( .A(n4437), .B(n4438), .Z(n2748) );
  CIVXL U5369 ( .A(n4564), .Z(n4436) );
  CND2X1 U5370 ( .A(n4439), .B(a[20]), .Z(n4442) );
  CIVXL U5371 ( .A(n4202), .Z(n4439) );
  CND2XL U5372 ( .A(n1454), .B(n1433), .Z(n4443) );
  CND2XL U5373 ( .A(n1454), .B(n1435), .Z(n4444) );
  CND2XL U5374 ( .A(n1433), .B(n1435), .Z(n4445) );
  CND3X1 U5375 ( .A(n4443), .B(n4444), .C(n4445), .Z(n1422) );
  CND2XL U5376 ( .A(n1401), .B(n1399), .Z(n4446) );
  CND2X1 U5377 ( .A(n1401), .B(n1422), .Z(n4447) );
  CND2XL U5378 ( .A(n1399), .B(n1422), .Z(n4448) );
  CND3X1 U5379 ( .A(n4446), .B(n4447), .C(n4448), .Z(n1392) );
  CND2X1 U5380 ( .A(n470), .B(n171), .Z(n4450) );
  CND2X2 U5381 ( .A(n4449), .B(net17451), .Z(n4451) );
  CND2X2 U5382 ( .A(n4450), .B(n4451), .Z(product[41]) );
  CIVX2 U5383 ( .A(n171), .Z(net17451) );
  CND2X1 U5384 ( .A(n371), .B(n162), .Z(n4454) );
  CND2X2 U5385 ( .A(n4452), .B(n4453), .Z(n4455) );
  CND2X2 U5386 ( .A(n4454), .B(n4455), .Z(product[50]) );
  CIVX2 U5387 ( .A(n162), .Z(n4453) );
  CND2XL U5388 ( .A(n513), .B(n176), .Z(n4456) );
  CND2X2 U5389 ( .A(net17438), .B(net17439), .Z(n4457) );
  CND2X2 U5390 ( .A(n4456), .B(n4457), .Z(product[36]) );
  CIVX1 U5391 ( .A(n3250), .Z(net17438) );
  CIVX2 U5392 ( .A(n176), .Z(net17439) );
  CIVXL U5393 ( .A(n594), .Z(n596) );
  COND2XL U5394 ( .A(n54), .B(n2611), .C(n4507), .D(n2610), .Z(n2086) );
  CND2IXL U5395 ( .B(n3244), .A(n4582), .Z(n2548) );
  CENXL U5396 ( .A(n4582), .B(n4550), .Z(n2534) );
  CENXL U5397 ( .A(n4568), .B(n4582), .Z(n2543) );
  CND2IXL U5398 ( .B(n3244), .A(n3760), .Z(n2515) );
  CENXL U5399 ( .A(n3760), .B(n4543), .Z(n2508) );
  CENXL U5400 ( .A(n3244), .B(n3760), .Z(n2514) );
  CENXL U5401 ( .A(n3760), .B(n4550), .Z(n2501) );
  CENXL U5402 ( .A(n3760), .B(n4551), .Z(n2500) );
  CENXL U5403 ( .A(n3760), .B(n4542), .Z(n2509) );
  CENXL U5404 ( .A(n4568), .B(n3760), .Z(n2510) );
  CENXL U5405 ( .A(n3760), .B(n4554), .Z(n2497) );
  CENXL U5406 ( .A(n4603), .B(n4564), .Z(n2253) );
  CENXL U5407 ( .A(n4597), .B(n4564), .Z(n2319) );
  CENXL U5408 ( .A(n4595), .B(n4564), .Z(n2352) );
  CENXL U5409 ( .A(n3828), .B(n4564), .Z(n2385) );
  CENXL U5410 ( .A(n4591), .B(n4564), .Z(n2418) );
  CENXL U5411 ( .A(n4587), .B(n4564), .Z(n2451) );
  CENXL U5412 ( .A(n4582), .B(n4564), .Z(n2517) );
  CENXL U5413 ( .A(n4580), .B(n4564), .Z(n2550) );
  CIVX2 U5414 ( .A(n4458), .Z(n4459) );
  CENXL U5415 ( .A(n3748), .B(n4582), .Z(n2547) );
  CENXL U5416 ( .A(n3748), .B(n4598), .Z(n2349) );
  CENXL U5417 ( .A(n3747), .B(n4600), .Z(n2316) );
  CENXL U5418 ( .A(n3747), .B(n4595), .Z(n2382) );
  CENXL U5419 ( .A(n3747), .B(n4575), .Z(n2646) );
  COND1X1 U5420 ( .A(n281), .B(net16472), .C(n282), .Z(n280) );
  COND1X1 U5421 ( .A(n248), .B(net16472), .C(n249), .Z(n247) );
  COND1X1 U5422 ( .A(n305), .B(net16472), .C(n306), .Z(n304) );
  COND2X1 U5423 ( .A(n63), .B(n2579), .C(n2578), .D(n4505), .Z(n2054) );
  CNIVX4 U5424 ( .A(n18), .Z(n4461) );
  CENXL U5425 ( .A(n4583), .B(n4565), .Z(n2516) );
  CENXL U5426 ( .A(n4583), .B(n4541), .Z(n2544) );
  CENXL U5427 ( .A(n4583), .B(n4545), .Z(n2539) );
  CENXL U5428 ( .A(n4583), .B(n4543), .Z(n2541) );
  CENXL U5429 ( .A(n4583), .B(n4549), .Z(n2535) );
  CENXL U5430 ( .A(n4583), .B(n4547), .Z(n2537) );
  CENXL U5431 ( .A(n3645), .B(n4546), .Z(n2538) );
  CENXL U5432 ( .A(n4548), .B(n4583), .Z(n2536) );
  CENXL U5433 ( .A(n3909), .B(n4541), .Z(n2676) );
  CENXL U5434 ( .A(n3909), .B(n4542), .Z(n2674) );
  CENXL U5435 ( .A(n4567), .B(n3909), .Z(n2677) );
  CENXL U5436 ( .A(n3909), .B(n4540), .Z(n2678) );
  CENXL U5437 ( .A(n3909), .B(n4546), .Z(n2670) );
  CENXL U5438 ( .A(n3909), .B(n4545), .Z(n2671) );
  CENXL U5439 ( .A(n3909), .B(n4548), .Z(n2668) );
  CENXL U5440 ( .A(n3909), .B(n4547), .Z(n2669) );
  CENXL U5441 ( .A(n3102), .B(n4543), .Z(n2673) );
  CENXL U5442 ( .A(n3909), .B(n4549), .Z(n2667) );
  CENXL U5443 ( .A(n4597), .B(n4565), .Z(n2318) );
  CENXL U5444 ( .A(n4597), .B(n4555), .Z(n2331) );
  CENXL U5445 ( .A(n4597), .B(n4549), .Z(n2337) );
  CENXL U5446 ( .A(n4597), .B(n4548), .Z(n2338) );
  CENXL U5447 ( .A(n4597), .B(n4547), .Z(n2339) );
  CENXL U5448 ( .A(n4597), .B(n4546), .Z(n2340) );
  CENXL U5449 ( .A(n4597), .B(n4545), .Z(n2341) );
  CENXL U5450 ( .A(n4597), .B(n4543), .Z(n2343) );
  CENXL U5451 ( .A(n4597), .B(n4540), .Z(n2348) );
  CIVX8 U5452 ( .A(n4586), .Z(n4585) );
  CENXL U5453 ( .A(n4585), .B(n4560), .Z(n2491) );
  CENXL U5454 ( .A(n4585), .B(n4561), .Z(n2490) );
  CENXL U5455 ( .A(n4591), .B(n4556), .Z(n2429) );
  CENXL U5456 ( .A(n4591), .B(n4557), .Z(n2428) );
  CENXL U5457 ( .A(n4591), .B(n4558), .Z(n2427) );
  CENXL U5458 ( .A(n4591), .B(n4563), .Z(n2421) );
  CENXL U5459 ( .A(n4591), .B(n4559), .Z(n2426) );
  CENXL U5460 ( .A(n4591), .B(net16104), .Z(n2420) );
  CIVX8 U5461 ( .A(a[0]), .Z(n6) );
  CNIVX1 U5462 ( .A(n2807), .Z(n4569) );
  COND2X1 U5463 ( .A(net18772), .B(n2683), .C(net17297), .D(n2682), .Z(n2157)
         );
  COND2X1 U5464 ( .A(n54), .B(n2612), .C(n4506), .D(n2611), .Z(n2087) );
  CENX2 U5465 ( .A(a[2]), .B(n4574), .Z(n2826) );
  COND2X1 U5466 ( .A(n4316), .B(n2563), .C(n2562), .D(n4505), .Z(n2038) );
  CIVXL U5467 ( .A(n57), .Z(n4581) );
  CND2XL U5468 ( .A(n516), .B(n758), .Z(n507) );
  CNR2X2 U5469 ( .A(n923), .B(n938), .Z(n409) );
  CND2XL U5470 ( .A(n1287), .B(n1289), .Z(n4537) );
  CNR2IX1 U5471 ( .B(n3750), .A(n3121), .Z(n2025) );
  CENXL U5472 ( .A(n3748), .B(n4571), .Z(n2778) );
  CENX1 U5473 ( .A(n4602), .B(n4555), .Z(n2265) );
  CIVXL U5474 ( .A(n266), .Z(n264) );
  CANR1XL U5475 ( .A(n4486), .B(n323), .C(n314), .Z(n310) );
  CNR2X1 U5476 ( .A(n302), .B(n295), .Z(n293) );
  CAN2XL U5477 ( .A(n785), .B(n697), .Z(n4473) );
  CND2X1 U5478 ( .A(n1665), .B(n1674), .Z(n683) );
  CND2XL U5479 ( .A(n788), .B(n709), .Z(n206) );
  CND2XL U5480 ( .A(n1348), .B(n1325), .Z(n4536) );
  CENX1 U5481 ( .A(n4602), .B(n4556), .Z(n2264) );
  CENX1 U5482 ( .A(n4602), .B(n4557), .Z(n2263) );
  CENX1 U5483 ( .A(n4602), .B(n4553), .Z(n2267) );
  CENX1 U5484 ( .A(n4602), .B(n4559), .Z(n2261) );
  CENX1 U5485 ( .A(n4602), .B(n4558), .Z(n2262) );
  CENX1 U5486 ( .A(n4602), .B(n4541), .Z(n2280) );
  CENX1 U5487 ( .A(n4037), .B(net16102), .Z(n2617) );
  CENX1 U5488 ( .A(n4585), .B(n4559), .Z(n2492) );
  COND2X1 U5489 ( .A(n9), .B(n2767), .C(n6), .D(n2766), .Z(n2240) );
  COND2XL U5490 ( .A(n27), .B(n2711), .C(net17297), .D(n2710), .Z(n2185) );
  COND2XL U5491 ( .A(n4461), .B(n4328), .C(n2746), .D(n4510), .Z(n1738) );
  CENX1 U5492 ( .A(n4602), .B(n4562), .Z(n2258) );
  CENX1 U5493 ( .A(n4602), .B(n2785), .Z(n2257) );
  CND2X2 U5494 ( .A(n4468), .B(n4469), .Z(n2821) );
  CND2X2 U5495 ( .A(n3420), .B(n359), .Z(n353) );
  CND2XL U5496 ( .A(n770), .B(n3172), .Z(n188) );
  CENXL U5497 ( .A(n545), .B(n4470), .Z(product[32]) );
  CAN2X1 U5498 ( .A(n762), .B(n544), .Z(n4470) );
  CND2XL U5499 ( .A(n4475), .B(n618), .Z(n189) );
  CND2XL U5500 ( .A(n541), .B(n761), .Z(n179) );
  CND2XL U5501 ( .A(n355), .B(n331), .Z(n329) );
  CENX1 U5502 ( .A(n4471), .B(n676), .Z(product[13]) );
  CAN2XL U5503 ( .A(n781), .B(n675), .Z(n4471) );
  CEOX1 U5504 ( .A(n194), .B(n3606), .Z(product[18]) );
  CND2XL U5505 ( .A(n776), .B(n4218), .Z(n194) );
  CNR2X2 U5506 ( .A(n353), .B(n309), .Z(n307) );
  CND2IXL U5507 ( .B(n556), .A(net17791), .Z(n182) );
  CND2XL U5508 ( .A(n568), .B(n765), .Z(n183) );
  CND2XL U5509 ( .A(n3969), .B(n772), .Z(n190) );
  CND2XL U5510 ( .A(n4169), .B(n656), .Z(n195) );
  CND2X2 U5511 ( .A(n3257), .B(n750), .Z(n416) );
  CAN2XL U5512 ( .A(n779), .B(n3987), .Z(n4472) );
  CNR2X2 U5513 ( .A(n333), .B(n4482), .Z(n283) );
  CENX1 U5514 ( .A(net17211), .B(n553), .Z(product[31]) );
  CIVXL U5515 ( .A(n389), .Z(n746) );
  CIVXL U5516 ( .A(n402), .Z(n747) );
  CND2XL U5517 ( .A(n3490), .B(n3372), .Z(n193) );
  CENX2 U5518 ( .A(n166), .B(n411), .Z(product[46]) );
  CND2X2 U5519 ( .A(n745), .B(n744), .Z(n365) );
  CENX1 U5520 ( .A(n698), .B(n4473), .Z(product[9]) );
  CND2XL U5521 ( .A(n4488), .B(n683), .Z(n200) );
  CND2XL U5522 ( .A(n786), .B(n701), .Z(n204) );
  CEOXL U5523 ( .A(n204), .B(n3245), .Z(product[8]) );
  CND2XL U5524 ( .A(n4489), .B(n688), .Z(n201) );
  CIVXL U5525 ( .A(n324), .Z(n741) );
  CND2X2 U5526 ( .A(n4479), .B(n742), .Z(n333) );
  CNR2X1 U5527 ( .A(n957), .B(n974), .Z(n433) );
  COAN1XL U5528 ( .A(n327), .B(n291), .C(n292), .Z(n4477) );
  CANR1XL U5529 ( .A(n314), .B(n293), .C(n294), .Z(n292) );
  COND1X1 U5530 ( .A(n724), .B(n722), .C(n723), .Z(n721) );
  COND1X1 U5531 ( .A(n257), .B(net16472), .C(n258), .Z(n256) );
  CANR1X1 U5532 ( .A(n729), .B(n4496), .C(n726), .Z(n724) );
  CND2XL U5533 ( .A(n4493), .B(n714), .Z(n207) );
  CND2XL U5534 ( .A(n4492), .B(n706), .Z(n205) );
  COR2X2 U5535 ( .A(n827), .B(n834), .Z(n4486) );
  CEOXL U5536 ( .A(n3297), .B(n206), .Z(product[6]) );
  COR2XL U5537 ( .A(n1740), .B(n794), .Z(n4491) );
  CND2XL U5538 ( .A(n1713), .B(n1716), .Z(n709) );
  CND2XL U5539 ( .A(n1723), .B(n2249), .Z(n723) );
  CENXL U5540 ( .A(n4463), .B(n4557), .Z(n2296) );
  CENXL U5541 ( .A(n4463), .B(n4556), .Z(n2297) );
  CENXL U5542 ( .A(n4600), .B(n4560), .Z(n2293) );
  CENXL U5543 ( .A(n4600), .B(n4558), .Z(n2295) );
  CENXL U5544 ( .A(n4600), .B(n4559), .Z(n2294) );
  CNR2IX1 U5545 ( .B(n3244), .A(n4507), .Z(n2089) );
  COND2XL U5546 ( .A(n4461), .B(n2743), .C(n2742), .D(n4510), .Z(n2216) );
  CENXL U5547 ( .A(n4580), .B(net16104), .Z(n2552) );
  CENXL U5548 ( .A(n4580), .B(net16102), .Z(n2551) );
  CENXL U5549 ( .A(n4582), .B(n4562), .Z(n2522) );
  CENXL U5550 ( .A(n4600), .B(n4561), .Z(n2292) );
  CENXL U5551 ( .A(n4600), .B(n4562), .Z(n2291) );
  CENXL U5552 ( .A(n4600), .B(n4564), .Z(n2286) );
  CENXL U5553 ( .A(n4600), .B(n4563), .Z(n2289) );
  CENXL U5554 ( .A(n4600), .B(n2785), .Z(n2290) );
  CENXL U5555 ( .A(n4600), .B(net16104), .Z(n2288) );
  CENXL U5556 ( .A(n4600), .B(net16102), .Z(n2287) );
  CENXL U5557 ( .A(n3622), .B(n4565), .Z(n2549) );
  CNIVX4 U5558 ( .A(n2791), .Z(n4557) );
  CND2XL U5559 ( .A(n534), .B(n760), .Z(n525) );
  CND2XL U5560 ( .A(n489), .B(n516), .Z(n487) );
  CNR2IXL U5561 ( .B(n498), .A(n3757), .Z(n489) );
  CND2XL U5562 ( .A(n751), .B(n449), .Z(n169) );
  COND1XL U5563 ( .A(n507), .B(n545), .C(n508), .Z(n506) );
  CENX1 U5564 ( .A(n524), .B(n177), .Z(product[35]) );
  COND1XL U5565 ( .A(n496), .B(n545), .C(n497), .Z(n495) );
  CENX1 U5566 ( .A(n531), .B(n178), .Z(product[34]) );
  COND1X1 U5567 ( .A(n532), .B(n545), .C(n533), .Z(n531) );
  CENX1 U5568 ( .A(n542), .B(n179), .Z(product[33]) );
  CENX1 U5569 ( .A(n584), .B(n185), .Z(product[27]) );
  CND2XL U5570 ( .A(n583), .B(n767), .Z(n185) );
  CND2XL U5571 ( .A(n596), .B(n768), .Z(n585) );
  CEOXL U5572 ( .A(n188), .B(n611), .Z(product[24]) );
  CND2XL U5573 ( .A(n4150), .B(n768), .Z(n186) );
  CANR1XL U5574 ( .A(n758), .B(n517), .C(n510), .Z(n508) );
  CANR1XL U5575 ( .A(n768), .B(n3770), .C(n590), .Z(n586) );
  CENX1 U5576 ( .A(n380), .B(n163), .Z(product[49]) );
  CND2XL U5577 ( .A(n745), .B(n379), .Z(n163) );
  CENX1 U5578 ( .A(n404), .B(n165), .Z(product[47]) );
  CENX1 U5579 ( .A(n673), .B(n198), .Z(product[14]) );
  CND2X1 U5580 ( .A(n774), .B(n634), .Z(n192) );
  COND1XL U5581 ( .A(n636), .B(n3606), .C(n4226), .Z(n635) );
  CENX1 U5582 ( .A(n629), .B(n191), .Z(product[21]) );
  CENX1 U5583 ( .A(n352), .B(n161), .Z(product[51]) );
  CND2XL U5584 ( .A(n4479), .B(n351), .Z(n161) );
  CND2XL U5585 ( .A(n3257), .B(n4025), .Z(n167) );
  CND2XL U5586 ( .A(n3420), .B(n750), .Z(n427) );
  CANR1XL U5587 ( .A(n766), .B(n574), .C(n571), .Z(n569) );
  COND1XL U5588 ( .A(n389), .B(n399), .C(n392), .Z(n388) );
  CND2XL U5589 ( .A(n750), .B(n434), .Z(n168) );
  CANR1XL U5590 ( .A(n750), .B(n439), .C(n432), .Z(n428) );
  CNR2X1 U5591 ( .A(n627), .B(n622), .Z(n620) );
  COR2X1 U5592 ( .A(n1483), .B(n1504), .Z(n4475) );
  CND2X1 U5593 ( .A(n1436), .B(n1413), .Z(n592) );
  CND2X1 U5594 ( .A(n1015), .B(n1036), .Z(n469) );
  CND2X1 U5595 ( .A(n1437), .B(n1460), .Z(n603) );
  CND2X1 U5596 ( .A(n3131), .B(n3829), .Z(n583) );
  CND2XL U5597 ( .A(n742), .B(n342), .Z(n160) );
  CND2XL U5598 ( .A(n355), .B(n4479), .Z(n344) );
  CENX1 U5599 ( .A(n202), .B(n695), .Z(product[10]) );
  CENX1 U5600 ( .A(n689), .B(n201), .Z(product[11]) );
  CND2XL U5601 ( .A(n4486), .B(n316), .Z(n158) );
  CENX1 U5602 ( .A(n304), .B(n157), .Z(product[55]) );
  CND2XL U5603 ( .A(n739), .B(n303), .Z(n157) );
  CND2XL U5604 ( .A(n736), .B(n266), .Z(n154) );
  CND2XL U5605 ( .A(n355), .B(n272), .Z(n268) );
  CND2XL U5606 ( .A(n355), .B(n283), .Z(n281) );
  CND2X1 U5607 ( .A(n4491), .B(n218), .Z(n150) );
  CNR2X1 U5608 ( .A(n1653), .B(n1664), .Z(n674) );
  COND1XL U5609 ( .A(n324), .B(n334), .C(n327), .Z(n323) );
  CANR1XL U5610 ( .A(n233), .B(n356), .C(n236), .Z(n232) );
  CNR2X1 U5611 ( .A(n1627), .B(n1640), .Z(n665) );
  CNR2X1 U5612 ( .A(n1525), .B(n1544), .Z(n627) );
  COND1XL U5613 ( .A(n295), .B(n303), .C(n296), .Z(n294) );
  COR2X1 U5614 ( .A(n1612), .B(n1597), .Z(n4480) );
  COR2X1 U5615 ( .A(n1563), .B(n1580), .Z(n4481) );
  CND2X1 U5616 ( .A(n1627), .B(n1640), .Z(n666) );
  CND2X1 U5617 ( .A(n1275), .B(n1304), .Z(n552) );
  CND2X1 U5618 ( .A(n893), .B(n906), .Z(n392) );
  CND2X1 U5619 ( .A(n1653), .B(n1664), .Z(n675) );
  CND2X1 U5620 ( .A(n1597), .B(n1612), .Z(n656) );
  CND2X1 U5621 ( .A(n1563), .B(n1580), .Z(n641) );
  CND2X1 U5622 ( .A(n907), .B(n922), .Z(n403) );
  CND2X1 U5623 ( .A(n1333), .B(n1360), .Z(n568) );
  COR2X1 U5624 ( .A(n291), .B(n324), .Z(n4482) );
  CND2X1 U5625 ( .A(n4486), .B(n293), .Z(n291) );
  COR2X1 U5626 ( .A(n265), .B(n241), .Z(n4483) );
  COND1XL U5627 ( .A(n213), .B(net16472), .C(n214), .Z(n212) );
  CND2XL U5628 ( .A(n222), .B(n4491), .Z(n213) );
  CANR1XL U5629 ( .A(n4491), .B(n223), .C(n216), .Z(n214) );
  CENX1 U5630 ( .A(n4570), .B(n2809), .Z(n2776) );
  CENX1 U5631 ( .A(n207), .B(n4485), .Z(product[5]) );
  CENX1 U5632 ( .A(n208), .B(n721), .Z(product[4]) );
  CND2X1 U5633 ( .A(n4495), .B(n720), .Z(n208) );
  CENX1 U5634 ( .A(n256), .B(n153), .Z(product[59]) );
  CND2XL U5635 ( .A(n3759), .B(n255), .Z(n153) );
  COND1XL U5636 ( .A(n231), .B(net16472), .C(n232), .Z(n230) );
  CND2XL U5637 ( .A(n355), .B(n233), .Z(n231) );
  CENX1 U5638 ( .A(n247), .B(n152), .Z(product[60]) );
  CND2X1 U5639 ( .A(n4497), .B(n246), .Z(n152) );
  CEOXL U5640 ( .A(n724), .B(n209), .Z(product[3]) );
  CND2X1 U5641 ( .A(n791), .B(n723), .Z(n209) );
  CANR1XL U5642 ( .A(n4498), .B(n236), .C(n227), .Z(n225) );
  CENX1 U5643 ( .A(n4484), .B(n1565), .Z(n1563) );
  CENX1 U5644 ( .A(n1582), .B(n1567), .Z(n4484) );
  COND1XL U5645 ( .A(n4483), .B(n275), .C(n3763), .Z(n236) );
  CENX1 U5646 ( .A(n4568), .B(n4579), .Z(n2609) );
  CENX1 U5647 ( .A(n4568), .B(n4571), .Z(n2774) );
  CNR2X1 U5648 ( .A(n1701), .B(n1706), .Z(n700) );
  CAOR1X1 U5649 ( .A(n721), .B(n4495), .C(n718), .Z(n4485) );
  CND2X1 U5650 ( .A(n1701), .B(n1706), .Z(n701) );
  COR2X1 U5651 ( .A(n1674), .B(n1665), .Z(n4488) );
  CND2X1 U5652 ( .A(n1693), .B(n1700), .Z(n697) );
  CND2X1 U5653 ( .A(n1675), .B(n1684), .Z(n688) );
  COR2X1 U5654 ( .A(n1675), .B(n1684), .Z(n4489) );
  CENX1 U5655 ( .A(n210), .B(n729), .Z(product[2]) );
  CND2X1 U5656 ( .A(n4496), .B(n728), .Z(n210) );
  CNR2X1 U5657 ( .A(n806), .B(n803), .Z(n265) );
  COR2X1 U5658 ( .A(n807), .B(n812), .Z(n4490) );
  CND2X1 U5659 ( .A(n806), .B(n803), .Z(n266) );
  CND2X1 U5660 ( .A(n835), .B(n844), .Z(n327) );
  CND2X1 U5661 ( .A(n807), .B(n812), .Z(n279) );
  CND2X1 U5662 ( .A(n813), .B(n818), .Z(n296) );
  CND2X1 U5663 ( .A(n3759), .B(n4497), .Z(n241) );
  CND2XL U5664 ( .A(n1740), .B(n794), .Z(n218) );
  CENX1 U5665 ( .A(n4585), .B(n2809), .Z(n2512) );
  CNR2IXL U5666 ( .B(n3244), .A(n4510), .Z(n2219) );
  CENX1 U5667 ( .A(n4569), .B(n4600), .Z(n2312) );
  CENX1 U5668 ( .A(n2809), .B(net16541), .Z(n2710) );
  CND3X1 U5669 ( .A(n4534), .B(n4535), .C(n4536), .Z(n1314) );
  CNR2X1 U5670 ( .A(n1723), .B(n2249), .Z(n722) );
  COR2X1 U5671 ( .A(n1707), .B(n1712), .Z(n4492) );
  COR2X1 U5672 ( .A(n1717), .B(n1720), .Z(n4493) );
  CENX1 U5673 ( .A(n2189), .B(n1883), .Z(n1273) );
  CAN2XL U5674 ( .A(n3764), .B(n731), .Z(product[1]) );
  CND2X1 U5675 ( .A(n1707), .B(n1712), .Z(n706) );
  CND2X1 U5676 ( .A(n1717), .B(n1720), .Z(n714) );
  CND2X1 U5677 ( .A(n1721), .B(n1722), .Z(n720) );
  CND2X1 U5678 ( .A(n2250), .B(n2219), .Z(n728) );
  COR2X1 U5679 ( .A(n1721), .B(n1722), .Z(n4495) );
  COR2X1 U5680 ( .A(n2250), .B(n2219), .Z(n4496) );
  COR2X1 U5681 ( .A(n798), .B(n797), .Z(n4497) );
  CND2X1 U5682 ( .A(n798), .B(n797), .Z(n246) );
  COR2X1 U5683 ( .A(n796), .B(n795), .Z(n4498) );
  CND2X1 U5684 ( .A(n796), .B(n795), .Z(n229) );
  CENX1 U5685 ( .A(net15912), .B(n4549), .Z(n2403) );
  CENX1 U5686 ( .A(net17419), .B(n4552), .Z(n2400) );
  CENX1 U5687 ( .A(net17419), .B(n4555), .Z(n2397) );
  CENX1 U5688 ( .A(net17411), .B(n4561), .Z(n2391) );
  CENX1 U5689 ( .A(n4585), .B(n4558), .Z(n2493) );
  CENX1 U5690 ( .A(n4585), .B(net16104), .Z(n2486) );
  CENX1 U5691 ( .A(n4585), .B(n4555), .Z(n2496) );
  CENX1 U5692 ( .A(n4037), .B(net16104), .Z(n2618) );
  CENX1 U5693 ( .A(n4585), .B(n4557), .Z(n2494) );
  CENX1 U5694 ( .A(n4585), .B(net16102), .Z(n2485) );
  CENX1 U5695 ( .A(n4585), .B(n2785), .Z(n2488) );
  CENX1 U5696 ( .A(n4585), .B(n4563), .Z(n2487) );
  CENX1 U5697 ( .A(n4575), .B(n4560), .Z(n2623) );
  CENX1 U5698 ( .A(n4037), .B(n4559), .Z(n2624) );
  CENX1 U5699 ( .A(n4575), .B(n4558), .Z(n2625) );
  CENX1 U5700 ( .A(n4037), .B(n4563), .Z(n2619) );
  CENX1 U5701 ( .A(n4585), .B(n4549), .Z(n2502) );
  CENX1 U5702 ( .A(n4585), .B(n4548), .Z(n2503) );
  CENX1 U5703 ( .A(n4575), .B(n4556), .Z(n2627) );
  CENX1 U5704 ( .A(n4585), .B(n4547), .Z(n2504) );
  CENX1 U5705 ( .A(n4587), .B(n4544), .Z(n2474) );
  CENX1 U5706 ( .A(n4585), .B(n4546), .Z(n2505) );
  CENX1 U5707 ( .A(n4585), .B(n4541), .Z(n2511) );
  CENX1 U5708 ( .A(n4585), .B(n4540), .Z(n2513) );
  CENX1 U5709 ( .A(n4570), .B(n4540), .Z(n2777) );
  CENX1 U5710 ( .A(n4570), .B(n4548), .Z(n2767) );
  CENX1 U5711 ( .A(n4570), .B(n4549), .Z(n2766) );
  CENX1 U5712 ( .A(n4570), .B(n4547), .Z(n2768) );
  CENX1 U5713 ( .A(n4570), .B(n4542), .Z(n2773) );
  CENX1 U5714 ( .A(n4576), .B(n4546), .Z(n2637) );
  CENX1 U5715 ( .A(n4570), .B(n4546), .Z(n2769) );
  CENX1 U5716 ( .A(n4570), .B(n4543), .Z(n2772) );
  CENX1 U5717 ( .A(n4570), .B(n4545), .Z(n2770) );
  CENX1 U5718 ( .A(n4585), .B(n4565), .Z(n2483) );
  CENX1 U5719 ( .A(n4576), .B(n4565), .Z(n2615) );
  CENX1 U5720 ( .A(n4570), .B(n4565), .Z(n2747) );
  CIVX2 U5721 ( .A(n4590), .Z(n4589) );
  CENX1 U5722 ( .A(n4602), .B(n4547), .Z(n2273) );
  CENX1 U5723 ( .A(n4602), .B(n4546), .Z(n2274) );
  CENX1 U5724 ( .A(n4602), .B(n4548), .Z(n2272) );
  CENX1 U5725 ( .A(n4602), .B(n4545), .Z(n2275) );
  CENX1 U5726 ( .A(n4602), .B(n4544), .Z(n2276) );
  CENX1 U5727 ( .A(n4602), .B(n4554), .Z(n2266) );
  CENX1 U5728 ( .A(n4602), .B(n4549), .Z(n2271) );
  CENX1 U5729 ( .A(n4602), .B(n4543), .Z(n2277) );
  CENX1 U5730 ( .A(n4602), .B(n4550), .Z(n2270) );
  CENX1 U5731 ( .A(n4602), .B(n4552), .Z(n2268) );
  CENX1 U5732 ( .A(n4602), .B(n4542), .Z(n2278) );
  CENX1 U5733 ( .A(n4602), .B(n4551), .Z(n2269) );
  CENX1 U5734 ( .A(n4602), .B(n4540), .Z(n2282) );
  CENX1 U5735 ( .A(n4512), .B(n4562), .Z(n2720) );
  CENX1 U5736 ( .A(n4600), .B(n4549), .Z(n2304) );
  CENX1 U5737 ( .A(n4600), .B(n4548), .Z(n2305) );
  CENX1 U5738 ( .A(n4600), .B(n4547), .Z(n2306) );
  CENX1 U5739 ( .A(n4600), .B(n4546), .Z(n2307) );
  CENX1 U5740 ( .A(n4600), .B(n4545), .Z(n2308) );
  CENX1 U5741 ( .A(n4600), .B(n4552), .Z(n2301) );
  CENX1 U5742 ( .A(n4600), .B(n4554), .Z(n2299) );
  CENX1 U5743 ( .A(n4600), .B(n4550), .Z(n2303) );
  CENX1 U5744 ( .A(n4600), .B(n4553), .Z(n2300) );
  CENX1 U5745 ( .A(n4600), .B(n4543), .Z(n2310) );
  CENX1 U5746 ( .A(n4600), .B(n4551), .Z(n2302) );
  CENX1 U5747 ( .A(n4600), .B(n4541), .Z(n2313) );
  CENX1 U5748 ( .A(net16541), .B(net16104), .Z(n2684) );
  CENX1 U5749 ( .A(n4600), .B(n4542), .Z(n2311) );
  CENX1 U5750 ( .A(n4579), .B(n4557), .Z(n2593) );
  CENX1 U5751 ( .A(n4570), .B(net16102), .Z(n2749) );
  CENX1 U5752 ( .A(n4570), .B(n4563), .Z(n2751) );
  CENX1 U5753 ( .A(n4570), .B(n4558), .Z(n2757) );
  CENX1 U5754 ( .A(n4570), .B(net16104), .Z(n2750) );
  CENX1 U5755 ( .A(n4570), .B(n4561), .Z(n2754) );
  CENX1 U5756 ( .A(n4570), .B(n2785), .Z(n2752) );
  CENX1 U5757 ( .A(n4570), .B(n4557), .Z(n2758) );
  CENX1 U5758 ( .A(n4571), .B(n4551), .Z(n2764) );
  CENX1 U5759 ( .A(n4571), .B(n4552), .Z(n2763) );
  CENX1 U5760 ( .A(n4570), .B(n4559), .Z(n2756) );
  CENX1 U5761 ( .A(n4571), .B(n4554), .Z(n2761) );
  CENX1 U5762 ( .A(n4571), .B(n4553), .Z(n2762) );
  CENX1 U5763 ( .A(n4571), .B(n4550), .Z(n2765) );
  CENX1 U5764 ( .A(n4570), .B(n4544), .Z(n2771) );
  CIVX2 U5765 ( .A(n4202), .Z(n4587) );
  CIVX2 U5766 ( .A(n4093), .Z(n4576) );
  CIVX2 U5767 ( .A(n4590), .Z(n4588) );
  CNR2IXL U5768 ( .B(n3244), .A(n6), .Z(product[0]) );
  CENX1 U5769 ( .A(n4600), .B(n4555), .Z(n2298) );
  CENX1 U5770 ( .A(n4600), .B(n4565), .Z(n2285) );
  CNIVX4 U5771 ( .A(n2781), .Z(n4564) );
  CNIVX4 U5772 ( .A(n2802), .Z(n4546) );
  CNIVX4 U5773 ( .A(n2803), .Z(n4545) );
  CNIVX4 U5774 ( .A(n2780), .Z(n4565) );
  CNIVX4 U5775 ( .A(n2805), .Z(n4543) );
  CNIVX4 U5776 ( .A(n2806), .Z(n4542) );
  CNIVX4 U5777 ( .A(n2808), .Z(n4541) );
  CENX1 U5778 ( .A(n343), .B(n160), .Z(product[52]) );
  CND2X1 U5779 ( .A(n2251), .B(n1739), .Z(n731) );
  COND2XL U5780 ( .A(n3210), .B(n3677), .C(n6), .D(n2779), .Z(n1739) );
  COND2X1 U5781 ( .A(net16309), .B(n2664), .C(n3644), .D(n2663), .Z(n2139) );
  CIVX1 U5782 ( .A(n4502), .Z(n4503) );
  CNIVX4 U5783 ( .A(net18832), .Z(net16472) );
  CENX4 U5784 ( .A(n4085), .B(n3785), .Z(n4508) );
  CENXL U5785 ( .A(n4595), .B(n4554), .Z(n2365) );
  CENXL U5786 ( .A(n4595), .B(n4551), .Z(n2368) );
  CENXL U5787 ( .A(n4595), .B(n4553), .Z(n2366) );
  CENX1 U5788 ( .A(n4568), .B(n4595), .Z(n2378) );
  COND2XL U5789 ( .A(net16309), .B(n2678), .C(n3644), .D(n2677), .Z(n2153) );
  COND2XL U5790 ( .A(net18610), .B(n2674), .C(n3644), .D(n2673), .Z(n2149) );
  COND2XL U5791 ( .A(net18896), .B(n2668), .C(n3644), .D(n2667), .Z(n2143) );
  COND2XL U5792 ( .A(net18610), .B(n2676), .C(n3644), .D(n2675), .Z(n2151) );
  COND2XL U5793 ( .A(net18896), .B(n2675), .C(n3644), .D(n2674), .Z(n2150) );
  COND2XL U5794 ( .A(net16309), .B(n2679), .C(n3644), .D(n2678), .Z(n2154) );
  COND2XL U5795 ( .A(net18897), .B(n2670), .C(n3644), .D(n2669), .Z(n2145) );
  CND2X4 U5796 ( .A(n2812), .B(net16496), .Z(n4511) );
  CENXL U5797 ( .A(n4597), .B(n4556), .Z(n2330) );
  CENXL U5798 ( .A(n4598), .B(n4563), .Z(n2322) );
  CENXL U5799 ( .A(n4598), .B(n2785), .Z(n2323) );
  CENXL U5800 ( .A(n4597), .B(n4562), .Z(n2324) );
  CENXL U5801 ( .A(n4598), .B(n4561), .Z(n2325) );
  CENXL U5802 ( .A(n4597), .B(n4560), .Z(n2326) );
  CENX1 U5803 ( .A(n4575), .B(n4557), .Z(n2626) );
  CENX1 U5804 ( .A(n4575), .B(n4544), .Z(n2639) );
  CND2IXL U5805 ( .B(n3751), .A(n3727), .Z(n2647) );
  CHA1X1 U5806 ( .A(n2210), .B(n1734), .CO(n1682), .S(n1683) );
  CND2XL U5807 ( .A(n1463), .B(n1484), .Z(n4513) );
  CND2XL U5808 ( .A(n1463), .B(n1465), .Z(n4514) );
  CND2XL U5809 ( .A(n1484), .B(n1465), .Z(n4515) );
  CND3X1 U5810 ( .A(n4513), .B(n4514), .C(n4515), .Z(n1460) );
  CND2XL U5811 ( .A(n1565), .B(n1582), .Z(n4517) );
  CND2XL U5812 ( .A(n1567), .B(n1582), .Z(n4518) );
  CENXL U5813 ( .A(n3748), .B(net17419), .Z(n2415) );
  CND2IXL U5814 ( .B(n3751), .A(net17419), .Z(n2416) );
  CNR2X1 U5815 ( .A(n1461), .B(n1482), .Z(n605) );
  CIVX1 U5816 ( .A(n4058), .Z(n4519) );
  CNR2X2 U5817 ( .A(n3518), .B(n543), .Z(n534) );
  CIVXL U5818 ( .A(n3518), .Z(n761) );
  CND2X1 U5819 ( .A(n1189), .B(n1191), .Z(n4522) );
  CEO3X2 U5820 ( .A(n2040), .B(n1863), .C(n1918), .Z(n1381) );
  CND2XL U5821 ( .A(n4530), .B(n1863), .Z(n4524) );
  CND2XL U5822 ( .A(n4530), .B(n1918), .Z(n4525) );
  CND2X1 U5823 ( .A(n1863), .B(n1918), .Z(n4526) );
  CND2X1 U5824 ( .A(n1377), .B(n1379), .Z(n4527) );
  CND2X1 U5825 ( .A(n1379), .B(n1381), .Z(n4528) );
  CND2X1 U5826 ( .A(n1377), .B(n1381), .Z(n4529) );
  CND2XL U5827 ( .A(n1295), .B(n1299), .Z(n4531) );
  CND2XL U5828 ( .A(n1295), .B(n1293), .Z(n4532) );
  CND2X1 U5829 ( .A(n1299), .B(n1293), .Z(n4533) );
  CND3X1 U5830 ( .A(n4531), .B(n4532), .C(n4533), .Z(n1286) );
  COND1XL U5831 ( .A(n556), .B(n564), .C(net17791), .Z(n555) );
  CND2IXL U5832 ( .B(n3750), .A(n3774), .Z(n2482) );
  CENX1 U5833 ( .A(n4501), .B(n4549), .Z(n2469) );
  COAN1X1 U5834 ( .A(n592), .B(n582), .C(n583), .Z(n579) );
  CENX1 U5835 ( .A(n450), .B(n169), .Z(product[43]) );
  CHA1X1 U5836 ( .A(n1731), .B(n2174), .CO(n1610), .S(n1611) );
  COND2X1 U5837 ( .A(n4120), .B(n3761), .C(n2515), .D(n4217), .Z(n1731) );
  CND2IXL U5838 ( .B(n3244), .A(n3909), .Z(n2680) );
  CEO3X2 U5839 ( .A(n1327), .B(n1348), .C(n1325), .Z(n1315) );
  CND2XL U5840 ( .A(n1327), .B(n1348), .Z(n4534) );
  CIVXL U5841 ( .A(n517), .Z(net16270) );
  CIVXL U5842 ( .A(net16274), .Z(n517) );
  CND2X1 U5843 ( .A(n1159), .B(n1186), .Z(n523) );
  CND2XL U5844 ( .A(n523), .B(n3840), .Z(n177) );
  CND2XL U5845 ( .A(n516), .B(net18817), .Z(n496) );
  CANR1XL U5846 ( .A(net18817), .B(n517), .C(net18061), .Z(n497) );
  COND2XL U5847 ( .A(n4063), .B(n3340), .C(n2647), .D(net16420), .Z(n1735) );
  COND1X2 U5848 ( .A(n412), .B(net16471), .C(n413), .Z(n411) );
  CIVX8 U5849 ( .A(n4604), .Z(n4602) );
  CND2X4 U5850 ( .A(n2822), .B(n4095), .Z(n54) );
  CND2X4 U5851 ( .A(n2821), .B(n4504), .Z(n63) );
  CND2X4 U5852 ( .A(n3252), .B(n78), .Z(n81) );
  CIVX2 U5853 ( .A(n212), .Z(product[63]) );
  CIVX2 U5854 ( .A(n890), .Z(n891) );
  CIVX2 U5855 ( .A(n824), .Z(n825) );
  CIVX2 U5856 ( .A(n810), .Z(n811) );
  CIVX2 U5857 ( .A(n800), .Z(n801) );
  CIVX2 U5858 ( .A(n794), .Z(n795) );
  CIVX2 U5859 ( .A(n722), .Z(n791) );
  CIVX2 U5860 ( .A(n700), .Z(n786) );
  CIVX2 U5861 ( .A(n693), .Z(n784) );
  CIVX2 U5862 ( .A(n633), .Z(n774) );
  CIVX2 U5863 ( .A(n295), .Z(n738) );
  CIVX2 U5864 ( .A(n731), .Z(n729) );
  CIVX2 U5865 ( .A(n728), .Z(n726) );
  CIVX2 U5866 ( .A(n714), .Z(n712) );
  CIVX2 U5867 ( .A(n706), .Z(n704) );
  CIVX2 U5868 ( .A(n688), .Z(n686) );
  CIVX2 U5869 ( .A(n683), .Z(n681) );
  CIVX2 U5870 ( .A(n656), .Z(n654) );
  CIVX2 U5871 ( .A(n627), .Z(n773) );
  CIVX2 U5872 ( .A(n618), .Z(n616) );
  CIVX2 U5873 ( .A(n591), .Z(n768) );
  CIVX2 U5874 ( .A(net19057), .Z(n441) );
  CIVX2 U5875 ( .A(n433), .Z(n750) );
  CIVX2 U5876 ( .A(n409), .Z(n748) );
  CIVX2 U5877 ( .A(n384), .Z(n382) );
  CIVX2 U5878 ( .A(n383), .Z(n381) );
  CIVX2 U5879 ( .A(n379), .Z(n377) );
  CIVX2 U5880 ( .A(n378), .Z(n745) );
  CIVX2 U5881 ( .A(n369), .Z(n744) );
  CIVX2 U5882 ( .A(n354), .Z(n356) );
  CIVX2 U5883 ( .A(n353), .Z(n355) );
  CIVX2 U5884 ( .A(n351), .Z(n349) );
  CIVX2 U5885 ( .A(n342), .Z(n340) );
  CIVX2 U5886 ( .A(n341), .Z(n742) );
  CIVX2 U5887 ( .A(n333), .Z(n331) );
  CIVX2 U5888 ( .A(n316), .Z(n314) );
  CIVX2 U5889 ( .A(n303), .Z(n301) );
  CIVX2 U5890 ( .A(n302), .Z(n739) );
  CIVX2 U5891 ( .A(n279), .Z(n277) );
  CIVX2 U5892 ( .A(n274), .Z(n272) );
  CIVX2 U5893 ( .A(n265), .Z(n736) );
  CIVX2 U5894 ( .A(n259), .Z(n257) );
  CIVX2 U5895 ( .A(n255), .Z(n253) );
  CIVX2 U5896 ( .A(n246), .Z(n244) );
  CIVX2 U5897 ( .A(n229), .Z(n227) );
  CIVX2 U5898 ( .A(n218), .Z(n216) );
endmodule


module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push0, _pushout_d, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, n147, n150, n152, n153, n156, n158,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, net6623, net13361, net13424, net13994,
         net14010, net14078, net14094, net16065, net16919, net16920, net16921,
         net17851, net17839, net17836, net14111, net26790, net14022, net14103,
         net14118, net14116, net14040, net13427, net13426, net13425, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] acc;
  wire   [1:0] cmd0;

  CFD2QX2 \q0_reg[31]  ( .D(n384), .CP(clk), .CD(n491), .Q(q0[31]) );
  CFD2QX2 \q0_reg[28]  ( .D(n323), .CP(clk), .CD(n491), .Q(q0[28]) );
  CFD2QX2 \q0_reg[26]  ( .D(n269), .CP(clk), .CD(n492), .Q(q0[26]) );
  CFD2QX2 \q0_reg[25]  ( .D(n383), .CP(clk), .CD(n491), .Q(q0[25]) );
  CFD2QX2 \q0_reg[24]  ( .D(n382), .CP(clk), .CD(n492), .Q(q0[24]) );
  CFD2QX2 \q0_reg[22]  ( .D(n322), .CP(clk), .CD(n492), .Q(q0[22]) );
  CFD2QX2 \q0_reg[0]  ( .D(n243), .CP(clk), .CD(n493), .Q(q0[0]) );
  CFD2QX2 \h0_reg[26]  ( .D(n371), .CP(clk), .CD(n494), .Q(h0[26]) );
  CFD2QX2 \h0_reg[5]  ( .D(n370), .CP(clk), .CD(n495), .Q(h0[5]) );
  CFD2QX2 \h0_reg[3]  ( .D(n369), .CP(clk), .CD(n495), .Q(h0[3]) );
  sfilt_DW01_add_2 add_43 ( .A({N272, N271, N270, N269, N268, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, 
        N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, 
        N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        N208}), .CI(1'b0), .SUM({N336, N335, N334, N333, N332, N331, N330, 
        N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, 
        N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, 
        N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, 
        N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280, N279, N278, N277, N276, N275, N274, N273}) );
  sfilt_DW01_add_6 add_39 ( .A({N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16}), .B(
        {n345, n328, n451, net17839, acc[59], n448, acc[57], n340, n449, n450, 
        n342, net17836, acc[51], net17851, acc[49], n333, acc[47:0]}), .CI(
        1'b0), .SUM({N207, N206, N205, N204, N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144}) );
  sfilt_DW_mult_tc_4 r300 ( .a(q0), .b({h0[31:3], n502, h0[1], n335}), 
        .product({N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, 
        N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, 
        N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23, N22, N21, N20, N19, N18, N17, N16}) );
  CFD2QX2 \q0_reg[3]  ( .D(n246), .CP(clk), .CD(n491), .Q(q0[3]) );
  CFD2QX1 \q0_reg[11]  ( .D(n254), .CP(clk), .CD(n493), .Q(q0[11]) );
  CFD2QX1 \q0_reg[19]  ( .D(n262), .CP(clk), .CD(n492), .Q(q0[19]) );
  CFD2QX1 \q0_reg[7]  ( .D(n250), .CP(clk), .CD(n493), .Q(q0[7]) );
  CFD2QXL \acc_reg[41]  ( .D(n168), .CP(clk), .CD(n497), .Q(acc[41]) );
  CFD2QXL \acc_reg[42]  ( .D(n167), .CP(clk), .CD(n497), .Q(acc[42]) );
  CFD2QXL \acc_reg[46]  ( .D(n163), .CP(clk), .CD(n497), .Q(acc[46]) );
  CFD2QXL \acc_reg[44]  ( .D(n165), .CP(clk), .CD(n497), .Q(acc[44]) );
  CFD2QXL \acc_reg[51]  ( .D(n158), .CP(clk), .CD(n497), .Q(acc[51]) );
  CFD2QXL \acc_reg[59]  ( .D(n150), .CP(clk), .CD(n496), .Q(acc[59]) );
  CFD2QXL \acc_reg[43]  ( .D(n166), .CP(clk), .CD(n497), .Q(acc[43]) );
  CFD2QXL \acc_reg[21]  ( .D(n188), .CP(clk), .CD(n499), .Q(acc[21]) );
  CFD2QXL \acc_reg[18]  ( .D(n191), .CP(clk), .CD(n499), .Q(acc[18]) );
  CFD2QXL \acc_reg[17]  ( .D(n192), .CP(clk), .CD(n499), .Q(acc[17]) );
  CFD2QXL \acc_reg[19]  ( .D(n190), .CP(clk), .CD(n499), .Q(acc[19]) );
  CFD2QXL \acc_reg[24]  ( .D(n185), .CP(clk), .CD(n499), .Q(acc[24]) );
  CFD2QXL \acc_reg[20]  ( .D(n189), .CP(clk), .CD(n499), .Q(acc[20]) );
  CFD2QXL \acc_reg[23]  ( .D(n186), .CP(clk), .CD(n499), .Q(acc[23]) );
  CFD2QXL \acc_reg[22]  ( .D(n187), .CP(clk), .CD(n499), .Q(acc[22]) );
  CFD2QXL \acc_reg[25]  ( .D(n184), .CP(clk), .CD(n499), .Q(acc[25]) );
  CFD2QXL \acc_reg[30]  ( .D(n179), .CP(clk), .CD(n498), .Q(acc[30]) );
  CFD2QXL \acc_reg[32]  ( .D(n177), .CP(clk), .CD(n498), .Q(acc[32]) );
  CFD2QXL \acc_reg[31]  ( .D(n178), .CP(clk), .CD(n498), .Q(acc[31]) );
  CFD2QXL \acc_reg[34]  ( .D(n175), .CP(clk), .CD(n498), .Q(acc[34]) );
  CFD2QXL \acc_reg[47]  ( .D(n162), .CP(clk), .CD(n497), .Q(acc[47]) );
  CFD2QXL \acc_reg[35]  ( .D(n174), .CP(clk), .CD(n498), .Q(acc[35]) );
  CFD2QXL \acc_reg[36]  ( .D(n173), .CP(clk), .CD(n498), .Q(acc[36]) );
  CFD2QXL \acc_reg[40]  ( .D(n169), .CP(clk), .CD(n498), .Q(acc[40]) );
  CFD2QXL \acc_reg[37]  ( .D(n172), .CP(clk), .CD(n498), .Q(acc[37]) );
  CFD2QXL \acc_reg[49]  ( .D(n160), .CP(clk), .CD(n497), .Q(acc[49]) );
  CFD2QXL \acc_reg[45]  ( .D(n164), .CP(clk), .CD(n497), .Q(acc[45]) );
  CFD2QXL \acc_reg[3]  ( .D(n206), .CP(clk), .CD(n500), .Q(acc[3]) );
  CFD2QX1 \q0_reg[5]  ( .D(n248), .CP(clk), .CD(n491), .Q(q0[5]) );
  CFD2QX1 \q0_reg[12]  ( .D(n319), .CP(clk), .CD(n492), .Q(q0[12]) );
  CFD2QXL \acc_reg[1]  ( .D(n208), .CP(clk), .CD(n501), .Q(acc[1]) );
  CFD2QXL \acc_reg[0]  ( .D(n209), .CP(clk), .CD(n501), .Q(acc[0]) );
  CFD2QXL \acc_reg[2]  ( .D(n207), .CP(clk), .CD(n500), .Q(acc[2]) );
  CFD2QX1 \q0_reg[13]  ( .D(n256), .CP(clk), .CD(n491), .Q(q0[13]) );
  CFD2QX1 \h0_reg[31]  ( .D(n360), .CP(clk), .CD(n493), .Q(h0[31]) );
  CFD2QX1 \h0_reg[30]  ( .D(n358), .CP(clk), .CD(n493), .Q(h0[30]) );
  CFD2QX2 \acc_reg[57]  ( .D(n152), .CP(clk), .CD(n496), .Q(acc[57]) );
  CFD2QX1 \h0_reg[1]  ( .D(n357), .CP(clk), .CD(n496), .Q(h0[1]) );
  CFD2QX1 \q0_reg[27]  ( .D(n359), .CP(clk), .CD(n491), .Q(q0[27]) );
  CFD2QX1 \h0_reg[28]  ( .D(n355), .CP(clk), .CD(n494), .Q(h0[28]) );
  CFD2QX1 \h0_reg[2]  ( .D(n213), .CP(clk), .CD(n496), .Q(h0[2]) );
  CFD2QX1 \q0_reg[15]  ( .D(n258), .CP(clk), .CD(n492), .Q(q0[15]) );
  CFD2QX1 \h0_reg[24]  ( .D(n361), .CP(clk), .CD(n494), .Q(h0[24]) );
  CFD2QX1 \h0_reg[8]  ( .D(n354), .CP(clk), .CD(n495), .Q(h0[8]) );
  CFD2QX1 \h0_reg[7]  ( .D(n363), .CP(clk), .CD(n495), .Q(h0[7]) );
  CFD2QX1 \h0_reg[13]  ( .D(n377), .CP(clk), .CD(n495), .Q(h0[13]) );
  CFD2QX1 \h0_reg[12]  ( .D(n347), .CP(clk), .CD(n495), .Q(h0[12]) );
  CFD2QX1 \h0_reg[15]  ( .D(n349), .CP(clk), .CD(n495), .Q(h0[15]) );
  CFD2QX1 \h0_reg[20]  ( .D(n373), .CP(clk), .CD(n494), .Q(h0[20]) );
  CFD2QX4 \q0_reg[16]  ( .D(n259), .CP(clk), .CD(n492), .Q(q0[16]) );
  CFD2QX1 \h0_reg[27]  ( .D(n353), .CP(clk), .CD(n494), .Q(h0[27]) );
  CFD2QX1 \h0_reg[19]  ( .D(n378), .CP(clk), .CD(n494), .Q(h0[19]) );
  CFD2QX1 \h0_reg[21]  ( .D(n352), .CP(clk), .CD(n494), .Q(h0[21]) );
  CFD2QX2 \q0_reg[23]  ( .D(n266), .CP(clk), .CD(n491), .Q(q0[23]) );
  CFD2QX1 \h0_reg[16]  ( .D(n379), .CP(clk), .CD(n494), .Q(h0[16]) );
  CFD2QX1 \h0_reg[25]  ( .D(n348), .CP(clk), .CD(n494), .Q(h0[25]) );
  CFD2QX1 \h0_reg[10]  ( .D(n381), .CP(clk), .CD(n495), .Q(h0[10]) );
  CFD2QX1 \h0_reg[22]  ( .D(n233), .CP(clk), .CD(n494), .Q(h0[22]) );
  CFD2QX1 \h0_reg[11]  ( .D(n350), .CP(clk), .CD(n495), .Q(h0[11]) );
  CFD2QX1 \h0_reg[9]  ( .D(n374), .CP(clk), .CD(n495), .Q(h0[9]) );
  CFD2QX1 \h0_reg[23]  ( .D(n351), .CP(clk), .CD(n494), .Q(h0[23]) );
  CFD2QX1 \h0_reg[17]  ( .D(n362), .CP(clk), .CD(n494), .Q(h0[17]) );
  CFD2QX1 \h0_reg[18]  ( .D(n380), .CP(clk), .CD(n494), .Q(h0[18]) );
  CFD2QX1 \q0_reg[18]  ( .D(n365), .CP(clk), .CD(n492), .Q(q0[18]) );
  CFD2QX1 \h0_reg[14]  ( .D(n368), .CP(clk), .CD(n495), .Q(h0[14]) );
  CFD2QX1 \h0_reg[29]  ( .D(n367), .CP(clk), .CD(n493), .Q(h0[29]) );
  CFD2QX2 \q0_reg[9]  ( .D(n252), .CP(clk), .CD(n493), .Q(q0[9]) );
  CFD2QX2 \q0_reg[21]  ( .D(n264), .CP(clk), .CD(n492), .Q(q0[21]) );
  CFD2QX2 \q0_reg[1]  ( .D(n316), .CP(clk), .CD(n493), .Q(q0[1]) );
  CFD2QX2 \q0_reg[2]  ( .D(n364), .CP(clk), .CD(n493), .Q(q0[2]) );
  CFD2XL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n1162), .Q(cmd0[1]), .QN(
        n426) );
  CFD2XL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n1162), .Q(cmd0[0]), .QN(
        n425) );
  CFD2XL push0_reg ( .D(pushin), .CP(clk), .CD(n1162), .Q(push0), .QN(net26790) );
  CFD2XL _pushout_reg ( .D(_pushout_d), .CP(clk), .CD(n1162), .Q(pushout) );
  CFD2XL \dout_reg[31]  ( .D(n307), .CP(clk), .CD(n1162), .Q(z[31]), .QN(n1161) );
  CFD2XL \dout_reg[30]  ( .D(n306), .CP(clk), .CD(n1162), .Q(z[30]), .QN(n1159) );
  CFD2XL \dout_reg[29]  ( .D(n305), .CP(clk), .CD(n1162), .Q(z[29]), .QN(n1157) );
  CFD2XL \dout_reg[28]  ( .D(n304), .CP(clk), .CD(n1162), .Q(z[28]), .QN(n1155) );
  CFD2XL \dout_reg[27]  ( .D(n303), .CP(clk), .CD(n1162), .Q(z[27]), .QN(n1153) );
  CFD2XL \dout_reg[26]  ( .D(n302), .CP(clk), .CD(n1162), .Q(z[26]), .QN(n1151) );
  CFD2XL \dout_reg[25]  ( .D(n301), .CP(clk), .CD(n1162), .Q(z[25]), .QN(n1149) );
  CFD2XL \dout_reg[24]  ( .D(n300), .CP(clk), .CD(n1162), .Q(z[24]), .QN(n1147) );
  CFD2XL \dout_reg[23]  ( .D(n299), .CP(clk), .CD(n1162), .Q(z[23]), .QN(n1145) );
  CFD2XL \dout_reg[22]  ( .D(n298), .CP(clk), .CD(n1162), .Q(z[22]), .QN(n1143) );
  CFD2XL \dout_reg[21]  ( .D(n297), .CP(clk), .CD(n1162), .Q(z[21]), .QN(n1141) );
  CFD2XL \dout_reg[20]  ( .D(n296), .CP(clk), .CD(n1162), .Q(z[20]), .QN(n1139) );
  CFD2XL \dout_reg[19]  ( .D(n295), .CP(clk), .CD(n1162), .Q(z[19]), .QN(n1137) );
  CFD2XL \dout_reg[18]  ( .D(n294), .CP(clk), .CD(n1162), .Q(z[18]), .QN(n1135) );
  CFD2XL \dout_reg[17]  ( .D(n293), .CP(clk), .CD(n1162), .Q(z[17]), .QN(n1133) );
  CFD2XL \dout_reg[16]  ( .D(n292), .CP(clk), .CD(n1162), .Q(z[16]), .QN(n1131) );
  CFD2XL \dout_reg[15]  ( .D(n291), .CP(clk), .CD(n1162), .Q(z[15]), .QN(n1129) );
  CFD2XL \dout_reg[14]  ( .D(n290), .CP(clk), .CD(n1162), .Q(z[14]), .QN(n1127) );
  CFD2XL \dout_reg[13]  ( .D(n289), .CP(clk), .CD(n1162), .Q(z[13]), .QN(n1125) );
  CFD2XL \dout_reg[12]  ( .D(n288), .CP(clk), .CD(n1162), .Q(z[12]), .QN(n1123) );
  CFD2XL \dout_reg[11]  ( .D(n287), .CP(clk), .CD(n1162), .Q(z[11]), .QN(n1121) );
  CFD2XL \dout_reg[10]  ( .D(n286), .CP(clk), .CD(n1162), .Q(z[10]), .QN(n1119) );
  CFD2XL \dout_reg[9]  ( .D(n285), .CP(clk), .CD(n1162), .Q(z[9]), .QN(n1117)
         );
  CFD2XL \dout_reg[8]  ( .D(n284), .CP(clk), .CD(n1162), .Q(z[8]), .QN(n1115)
         );
  CFD2XL \dout_reg[7]  ( .D(n283), .CP(clk), .CD(n1162), .Q(z[7]), .QN(n1113)
         );
  CFD2XL \dout_reg[6]  ( .D(n282), .CP(clk), .CD(n1162), .Q(z[6]), .QN(n1111)
         );
  CFD2XL \dout_reg[5]  ( .D(n281), .CP(clk), .CD(n1162), .Q(z[5]), .QN(n1109)
         );
  CFD2XL \dout_reg[4]  ( .D(n280), .CP(clk), .CD(n1162), .Q(z[4]), .QN(n1107)
         );
  CFD2XL \dout_reg[3]  ( .D(n279), .CP(clk), .CD(n1162), .Q(z[3]), .QN(n1105)
         );
  CFD2XL \dout_reg[1]  ( .D(n277), .CP(clk), .CD(n1162), .Q(z[1]), .QN(n1103)
         );
  CFD2XL \dout_reg[0]  ( .D(n276), .CP(clk), .CD(n1162), .Q(z[0]), .QN(n1101)
         );
  CFD2XL \dout_reg[2]  ( .D(n366), .CP(clk), .CD(n1162), .Q(z[2]) );
  CFD2XL \acc_reg[6]  ( .D(n203), .CP(clk), .CD(n1162), .Q(acc[6]), .QN(n1110)
         );
  CFD2XL \acc_reg[7]  ( .D(n202), .CP(clk), .CD(n1162), .Q(acc[7]), .QN(n1112)
         );
  CFD2XL \acc_reg[4]  ( .D(n205), .CP(clk), .CD(n1162), .Q(acc[4]), .QN(n1106)
         );
  CFD2XL \acc_reg[5]  ( .D(n204), .CP(clk), .CD(n1162), .Q(acc[5]), .QN(n1108)
         );
  CFD2XL \acc_reg[9]  ( .D(n200), .CP(clk), .CD(n1162), .Q(acc[9]), .QN(n1116)
         );
  CFD2XL \acc_reg[8]  ( .D(n201), .CP(clk), .CD(n1162), .Q(acc[8]), .QN(n1114)
         );
  CFD2XL \acc_reg[10]  ( .D(n199), .CP(clk), .CD(n1162), .Q(acc[10]), .QN(
        n1118) );
  CFD2XL \acc_reg[11]  ( .D(n198), .CP(clk), .CD(n1162), .Q(acc[11]), .QN(
        n1120) );
  CFD2XL \acc_reg[12]  ( .D(n197), .CP(clk), .CD(n1162), .Q(acc[12]), .QN(
        n1122) );
  CFD2XL \acc_reg[14]  ( .D(n195), .CP(clk), .CD(n1162), .Q(acc[14]), .QN(
        n1126) );
  CFD2XL \acc_reg[13]  ( .D(n196), .CP(clk), .CD(n1162), .Q(acc[13]), .QN(
        n1124) );
  CFD2XL \acc_reg[15]  ( .D(n194), .CP(clk), .CD(n1162), .Q(acc[15]), .QN(
        n1128) );
  CFD2XL \acc_reg[16]  ( .D(n193), .CP(clk), .CD(n1162), .Q(acc[16]), .QN(
        n1130) );
  CFD2XL \acc_reg[55]  ( .D(n407), .CP(clk), .CD(n1162), .Q(n449), .QN(n567)
         );
  CFD2XL \acc_reg[54]  ( .D(n395), .CP(clk), .CD(n1162), .Q(n450), .QN(n576)
         );
  CFD2XL \acc_reg[50]  ( .D(n417), .CP(clk), .CD(n1162), .Q(net17851), .QN(
        net13994) );
  CFD2XL \acc_reg[60]  ( .D(n421), .CP(clk), .CD(n1162), .Q(net17839), .QN(
        net14078) );
  CFD2XL \acc_reg[61]  ( .D(n399), .CP(clk), .CD(n1162), .Q(n451), .QN(n530)
         );
  CFD2XL \acc_reg[63]  ( .D(n210), .CP(clk), .CD(n501), .Q(n344), .QN(n343) );
  CFD2XL \acc_reg[53]  ( .D(n156), .CP(clk), .CD(n496), .QN(n341) );
  CFD2XL \acc_reg[56]  ( .D(n153), .CP(clk), .CD(n496), .QN(n339) );
  CFD2QX2 \q0_reg[20]  ( .D(n315), .CP(clk), .CD(n492), .Q(q0[20]) );
  CFD2X2 \acc_reg[58]  ( .D(n403), .CP(clk), .CD(n1162), .Q(n448), .QN(n548)
         );
  CFD2QX2 \acc_reg[38]  ( .D(n171), .CP(clk), .CD(n498), .Q(acc[38]) );
  CFD2X1 \acc_reg[52]  ( .D(n413), .CP(clk), .CD(n1162), .Q(net17836), .QN(
        net14010) );
  CFD2QX2 \acc_reg[39]  ( .D(n170), .CP(clk), .CD(n498), .Q(acc[39]) );
  CFD2QX2 \acc_reg[33]  ( .D(n176), .CP(clk), .CD(n498), .Q(acc[33]) );
  CFD2QX2 \acc_reg[27]  ( .D(n182), .CP(clk), .CD(n499), .Q(acc[27]) );
  CFD2QX2 \acc_reg[26]  ( .D(n318), .CP(clk), .CD(n499), .Q(acc[26]) );
  CFD2QX2 \acc_reg[28]  ( .D(n181), .CP(clk), .CD(n498), .Q(acc[28]) );
  CFD2QX2 \acc_reg[29]  ( .D(n180), .CP(clk), .CD(n498), .Q(acc[29]) );
  CFD2QX1 \q0_reg[4]  ( .D(n372), .CP(clk), .CD(n493), .Q(q0[4]) );
  CFD2QX1 \q0_reg[14]  ( .D(n257), .CP(clk), .CD(n492), .Q(q0[14]) );
  CFD2QX1 \h0_reg[4]  ( .D(n215), .CP(clk), .CD(n495), .Q(h0[4]) );
  CFD2QX1 \h0_reg[6]  ( .D(n356), .CP(clk), .CD(n495), .Q(h0[6]) );
  CFD2QX2 \q0_reg[6]  ( .D(n338), .CP(clk), .CD(n493), .Q(q0[6]) );
  CFD2X1 \h0_reg[0]  ( .D(n317), .CP(clk), .CD(n496), .Q(n335), .QN(n336) );
  CFD2XL \acc_reg[48]  ( .D(n161), .CP(clk), .CD(n497), .Q(n333), .QN(n334) );
  CFD2QX2 \q0_reg[29]  ( .D(n272), .CP(clk), .CD(n492), .Q(q0[29]) );
  CFD2QX4 \q0_reg[30]  ( .D(n273), .CP(clk), .CD(n491), .Q(q0[30]) );
  CFD2XL \acc_reg[62]  ( .D(n147), .CP(clk), .CD(n1162), .Q(n327), .QN(n326)
         );
  CFD2QX1 \q0_reg[10]  ( .D(n376), .CP(clk), .CD(n493), .Q(q0[10]) );
  CFD2QX2 \q0_reg[8]  ( .D(n375), .CP(clk), .CD(n493), .Q(q0[8]) );
  CFD2QX2 \q0_reg[17]  ( .D(n321), .CP(clk), .CD(n492), .Q(q0[17]) );
  CIVXL U308 ( .A(q0[17]), .Z(n308) );
  CIVX2 U309 ( .A(n308), .Z(n309) );
  CIVX1 U310 ( .A(n336), .Z(n310) );
  CDLY1XL U311 ( .A(q0[2]), .Z(n311) );
  CDLY1XL U312 ( .A(q0[18]), .Z(n312) );
  CIVXL U313 ( .A(q0[31]), .Z(n313) );
  CIVX2 U314 ( .A(n313), .Z(n314) );
  CANR2XL U315 ( .A(N78), .B(net16919), .C(N335), .D(net16920), .Z(net14111)
         );
  CANR2XL U316 ( .A(N167), .B(net16921), .C(N39), .D(net16919), .Z(n805) );
  CND2X1 U317 ( .A(n664), .B(n663), .Z(n170) );
  CANR2X1 U318 ( .A(N183), .B(net16921), .C(N55), .D(net16919), .Z(n664) );
  CNIVX1 U319 ( .A(n263), .Z(n315) );
  CNIVX1 U320 ( .A(n244), .Z(n316) );
  CNIVX1 U321 ( .A(n211), .Z(n317) );
  CNIVX1 U322 ( .A(n183), .Z(n318) );
  CNIVX1 U323 ( .A(n255), .Z(n319) );
  CNIVX1 U324 ( .A(n671), .Z(n320) );
  CNIVX1 U325 ( .A(n260), .Z(n321) );
  CNIVX1 U326 ( .A(n265), .Z(n322) );
  CNIVX1 U327 ( .A(n271), .Z(n323) );
  CDLY1XL U328 ( .A(q0[27]), .Z(n324) );
  CDLY1XL U329 ( .A(q0[8]), .Z(n325) );
  CMX2XL U330 ( .A0(q0[30]), .A1(q[30]), .S(n508), .Z(n273) );
  CMX2XL U331 ( .A0(q0[16]), .A1(q[16]), .S(n509), .Z(n259) );
  CMX2XL U332 ( .A0(q0[26]), .A1(q[26]), .S(n508), .Z(n269) );
  CIVX2 U333 ( .A(n326), .Z(n328) );
  CANR2XL U334 ( .A(n502), .B(n626), .C(h0[3]), .D(n629), .Z(n570) );
  CANR2XL U335 ( .A(n502), .B(n609), .C(h0[3]), .D(n612), .Z(n557) );
  CANR2XL U336 ( .A(n502), .B(n617), .C(h0[3]), .D(n620), .Z(n564) );
  CNIVXL U337 ( .A(N64), .Z(n329) );
  CDLY1XL U338 ( .A(q0[24]), .Z(n330) );
  CIVXL U339 ( .A(n330), .Z(n331) );
  CIVX2 U340 ( .A(n331), .Z(n332) );
  CANR2XL U341 ( .A(net16919), .B(N77), .C(N334), .D(net16920), .Z(n516) );
  CMX2XL U342 ( .A0(n312), .A1(q[18]), .S(n509), .Z(n261) );
  CMX2XL U343 ( .A0(q0[6]), .A1(q[6]), .S(n510), .Z(n249) );
  CND2X2 U344 ( .A(n877), .B(n504), .Z(n1060) );
  CND2X2 U345 ( .A(n735), .B(n1089), .Z(n1067) );
  CIVX3 U346 ( .A(n571), .Z(n877) );
  CIVX3 U347 ( .A(n582), .Z(n888) );
  CIVX3 U348 ( .A(n581), .Z(n893) );
  CND2X1 U349 ( .A(push0), .B(n423), .Z(n424) );
  CND4X1 U350 ( .A(net13425), .B(push0), .C(net13426), .D(net13427), .Z(
        net13424) );
  CNR3X1 U351 ( .A(n431), .B(net16921), .C(n432), .Z(n429) );
  CAOR2X1 U352 ( .A(N322), .B(net16920), .C(acc[49]), .D(net6623), .Z(n337) );
  CND2XL U353 ( .A(n797), .B(n796), .Z(n185) );
  CANR2XL U354 ( .A(N302), .B(net16920), .C(acc[29]), .D(net6623), .Z(n749) );
  CND2XL U355 ( .A(n750), .B(n749), .Z(n180) );
  CANR2XL U356 ( .A(N301), .B(net16920), .C(acc[28]), .D(net6623), .Z(n761) );
  CANR2XL U357 ( .A(N299), .B(net16920), .C(acc[26]), .D(net6623), .Z(n780) );
  CANR2XL U358 ( .A(N300), .B(net16920), .C(acc[27]), .D(net6623), .Z(n772) );
  CND2XL U359 ( .A(n762), .B(n761), .Z(n181) );
  CND2XL U360 ( .A(n781), .B(n780), .Z(n183) );
  CND2XL U361 ( .A(n773), .B(n772), .Z(n182) );
  CND2XL U362 ( .A(n738), .B(n737), .Z(n179) );
  CND2XL U363 ( .A(n720), .B(n719), .Z(n177) );
  CND2XL U364 ( .A(n728), .B(n727), .Z(n178) );
  CANR2XL U365 ( .A(N306), .B(net16920), .C(acc[33]), .D(net6623), .Z(n711) );
  CND2XL U366 ( .A(n712), .B(n711), .Z(n176) );
  CANR2XL U367 ( .A(N312), .B(net16920), .C(acc[39]), .D(net6623), .Z(n663) );
  CANR2XL U368 ( .A(N311), .B(net16920), .C(acc[38]), .D(net6623), .Z(n671) );
  CANR2XL U369 ( .A(N168), .B(net16921), .C(N40), .D(net16919), .Z(n797) );
  CND2X1 U370 ( .A(n422), .B(n412), .Z(n413) );
  CND2XL U371 ( .A(n428), .B(n416), .Z(n417) );
  CND2IX1 U372 ( .B(n424), .A(N194), .Z(n428) );
  CND2IX1 U373 ( .B(n424), .A(N196), .Z(n422) );
  CND2XL U374 ( .A(N199), .B(net16921), .Z(n545) );
  CND2XL U375 ( .A(n552), .B(n394), .Z(n395) );
  CND2XL U376 ( .A(N198), .B(net16921), .Z(n552) );
  CND2XL U377 ( .A(n672), .B(n320), .Z(n171) );
  CND2XL U378 ( .A(n545), .B(n406), .Z(n407) );
  CND2XL U379 ( .A(n648), .B(n647), .Z(n168) );
  CND2X1 U380 ( .A(N202), .B(net16921), .Z(n528) );
  CND2XL U381 ( .A(n515), .B(n398), .Z(n399) );
  CND2XL U382 ( .A(N205), .B(net16921), .Z(n515) );
  CND2XL U383 ( .A(n704), .B(n703), .Z(n175) );
  CND2XL U384 ( .A(n696), .B(n695), .Z(n174) );
  CND2XL U385 ( .A(n688), .B(n687), .Z(n173) );
  CND2XL U386 ( .A(N193), .B(net16921), .Z(n389) );
  CMX2XL U387 ( .A0(n314), .A1(q[31]), .S(n508), .Z(n274) );
  CNIVX1 U388 ( .A(n249), .Z(n338) );
  CND2XL U389 ( .A(N204), .B(net16921), .Z(n427) );
  CMX2XL U390 ( .A0(q0[22]), .A1(q[22]), .S(n508), .Z(n265) );
  CIVX2 U391 ( .A(n339), .Z(n340) );
  CIVX2 U392 ( .A(n341), .Z(n342) );
  CIVX2 U393 ( .A(n343), .Z(n345) );
  CND2IXL U394 ( .B(n346), .A(n523), .Z(n150) );
  COND1XL U395 ( .A(push0), .B(n541), .C(n524), .Z(n346) );
  CNIVX1 U396 ( .A(n223), .Z(n347) );
  CNIVX1 U397 ( .A(n236), .Z(n348) );
  CNIVX1 U398 ( .A(n226), .Z(n349) );
  CNIVX1 U399 ( .A(n222), .Z(n350) );
  CNIVX1 U400 ( .A(n234), .Z(n351) );
  CNIVX1 U401 ( .A(n232), .Z(n352) );
  CNIVX1 U402 ( .A(n238), .Z(n353) );
  CMXI2X2 U403 ( .A0(n1141), .A1(n1140), .S(net16065), .Z(n297) );
  CMXI2X2 U404 ( .A0(n1131), .A1(n1130), .S(net16065), .Z(n292) );
  CNIVX1 U405 ( .A(n219), .Z(n354) );
  CMXI2X2 U406 ( .A0(n1133), .A1(n1132), .S(net16065), .Z(n293) );
  CNIVX1 U407 ( .A(n239), .Z(n355) );
  CMXI2X2 U408 ( .A0(n1139), .A1(n1138), .S(net16065), .Z(n296) );
  CNIVX1 U409 ( .A(n217), .Z(n356) );
  CNIVX1 U410 ( .A(n212), .Z(n357) );
  CNIVX1 U411 ( .A(n241), .Z(n358) );
  CNIVX1 U412 ( .A(n270), .Z(n359) );
  CNIVX1 U413 ( .A(n242), .Z(n360) );
  CNIVX1 U414 ( .A(n235), .Z(n361) );
  CMXI2X2 U415 ( .A0(n1107), .A1(n1106), .S(net16065), .Z(n280) );
  CNIVX1 U416 ( .A(n228), .Z(n362) );
  CNIVX1 U417 ( .A(n218), .Z(n363) );
  CNIVX1 U418 ( .A(n245), .Z(n364) );
  CMXI2X2 U419 ( .A0(n1111), .A1(n1110), .S(net16065), .Z(n282) );
  CMXI2X2 U420 ( .A0(n1143), .A1(n1142), .S(net16065), .Z(n298) );
  CNIVX1 U421 ( .A(n261), .Z(n365) );
  CNIVX1 U422 ( .A(n278), .Z(n366) );
  CMXI2X2 U423 ( .A0(n1135), .A1(n1134), .S(net16065), .Z(n294) );
  CMXI2X2 U424 ( .A0(n1109), .A1(n1108), .S(net16065), .Z(n281) );
  CMXI2X2 U425 ( .A0(n1129), .A1(n1128), .S(net16065), .Z(n291) );
  CMXI2X2 U426 ( .A0(n1137), .A1(n1136), .S(net16065), .Z(n295) );
  CMXI2X2 U427 ( .A0(n1161), .A1(n1160), .S(net16065), .Z(n307) );
  CNIVX1 U428 ( .A(n240), .Z(n367) );
  CNIVX1 U429 ( .A(n225), .Z(n368) );
  CMXI2X2 U430 ( .A0(n1127), .A1(n1126), .S(net16065), .Z(n290) );
  CMXI2X2 U431 ( .A0(n1159), .A1(n1158), .S(net16065), .Z(n306) );
  CMXI2X2 U432 ( .A0(n1153), .A1(n1152), .S(net16065), .Z(n303) );
  CMXI2X2 U433 ( .A0(n1151), .A1(n1150), .S(net16065), .Z(n302) );
  CMXI2X2 U434 ( .A0(n1155), .A1(n1154), .S(net16065), .Z(n304) );
  CMXI2X2 U435 ( .A0(n1157), .A1(n1156), .S(net16065), .Z(n305) );
  CMXI2X2 U436 ( .A0(n1149), .A1(n1148), .S(net16065), .Z(n301) );
  CMXI2X2 U437 ( .A0(n1147), .A1(n1146), .S(net16065), .Z(n300) );
  CMXI2X2 U438 ( .A0(n1103), .A1(n1102), .S(net16065), .Z(n277) );
  CMXI2X2 U439 ( .A0(n1117), .A1(n1116), .S(net16065), .Z(n285) );
  CMXI2X2 U440 ( .A0(n1145), .A1(n1144), .S(net16065), .Z(n299) );
  CNIVX1 U441 ( .A(n214), .Z(n369) );
  CMX2XL U442 ( .A0(h0[3]), .A1(h[3]), .S(n513), .Z(n214) );
  CNIVX1 U443 ( .A(n216), .Z(n370) );
  CMX2XL U444 ( .A0(h0[5]), .A1(h[5]), .S(n512), .Z(n216) );
  CMXI2X2 U445 ( .A0(n1105), .A1(n1104), .S(net16065), .Z(n279) );
  CMXI2X2 U446 ( .A0(n1115), .A1(n1114), .S(net16065), .Z(n284) );
  CMXI2X2 U447 ( .A0(n1113), .A1(n1112), .S(net16065), .Z(n283) );
  CNIVX1 U448 ( .A(n237), .Z(n371) );
  CMX2XL U449 ( .A0(h0[26]), .A1(h[26]), .S(n511), .Z(n237) );
  CMXI2X2 U450 ( .A0(n1101), .A1(n1100), .S(net16065), .Z(n276) );
  CMXI2X2 U451 ( .A0(n1123), .A1(n1122), .S(net16065), .Z(n288) );
  CMXI2X2 U452 ( .A0(n1121), .A1(n1120), .S(net16065), .Z(n287) );
  CNIVX1 U453 ( .A(n247), .Z(n372) );
  CNIVX1 U454 ( .A(n231), .Z(n373) );
  CNIVX1 U455 ( .A(n220), .Z(n374) );
  CNIVX1 U456 ( .A(n251), .Z(n375) );
  CMX2XL U457 ( .A0(n325), .A1(q[8]), .S(n509), .Z(n251) );
  CMXI2X2 U458 ( .A0(n1119), .A1(n1118), .S(net16065), .Z(n286) );
  CNIVX1 U459 ( .A(n253), .Z(n376) );
  CNIVX1 U460 ( .A(n224), .Z(n377) );
  CNIVX1 U461 ( .A(n230), .Z(n378) );
  CMXI2X2 U462 ( .A0(n1125), .A1(n1124), .S(net16065), .Z(n289) );
  CNIVX1 U463 ( .A(n227), .Z(n379) );
  CNIVX1 U464 ( .A(n229), .Z(n380) );
  CNIVX1 U465 ( .A(n221), .Z(n381) );
  CNIVX1 U466 ( .A(n267), .Z(n382) );
  CNIVX1 U467 ( .A(n268), .Z(n383) );
  CNIVX1 U468 ( .A(n274), .Z(n384) );
  CANR2XL U469 ( .A(N190), .B(net16921), .C(net16919), .D(N62), .Z(n605) );
  CND2XL U470 ( .A(n605), .B(n604), .Z(n163) );
  CND2IXL U471 ( .B(n385), .A(n539), .Z(n153) );
  COND1XL U472 ( .A(push0), .B(n339), .C(n540), .Z(n385) );
  CND2IXL U473 ( .B(n386), .A(n560), .Z(n156) );
  COND1XL U474 ( .A(push0), .B(n341), .C(n561), .Z(n386) );
  CIVX1 U475 ( .A(net16919), .Z(n388) );
  CNR2X1 U476 ( .A(n388), .B(n445), .Z(n387) );
  CND2XL U477 ( .A(n389), .B(n390), .Z(n160) );
  CNR2X1 U478 ( .A(n387), .B(n337), .Z(n390) );
  CND2XL U479 ( .A(n427), .B(n420), .Z(n421) );
  CND2IXL U480 ( .B(n391), .A(n1095), .Z(n210) );
  COND1XL U481 ( .A(push0), .B(n1097), .C(n1096), .Z(n391) );
  CNR2X1 U482 ( .A(push0), .B(n576), .Z(n392) );
  CIVX1 U483 ( .A(n553), .Z(n393) );
  CNR2X1 U484 ( .A(n392), .B(n393), .Z(n394) );
  CNR2X1 U485 ( .A(push0), .B(n530), .Z(n396) );
  CIVX1 U486 ( .A(n516), .Z(n397) );
  CNR2X1 U487 ( .A(n396), .B(n397), .Z(n398) );
  CNR2X1 U488 ( .A(push0), .B(n548), .Z(n400) );
  CIVX1 U489 ( .A(n529), .Z(n401) );
  CNR2X1 U490 ( .A(n400), .B(n401), .Z(n402) );
  CND2X1 U491 ( .A(n528), .B(n402), .Z(n403) );
  CNR2X1 U492 ( .A(push0), .B(n567), .Z(n404) );
  CIVX1 U493 ( .A(n546), .Z(n405) );
  CNR2X1 U494 ( .A(n404), .B(n405), .Z(n406) );
  CND2IXL U495 ( .B(n408), .A(n591), .Z(n161) );
  CAOR2XL U496 ( .A(N321), .B(net16920), .C(n333), .D(net6623), .Z(n408) );
  CNR2XL U497 ( .A(N206), .B(n409), .Z(n430) );
  CND2XL U498 ( .A(net14111), .B(n434), .Z(n409) );
  CND2X1 U499 ( .A(n433), .B(net26790), .Z(n434) );
  CNR2X1 U500 ( .A(push0), .B(net14010), .Z(n410) );
  CIVX1 U501 ( .A(net14040), .Z(n411) );
  CNR2X1 U502 ( .A(n410), .B(n411), .Z(n412) );
  CNR2X1 U503 ( .A(push0), .B(net13994), .Z(n414) );
  CIVX1 U504 ( .A(net14022), .Z(n415) );
  CNR2X1 U505 ( .A(n414), .B(n415), .Z(n416) );
  CNR2X1 U506 ( .A(push0), .B(net14078), .Z(n418) );
  CIVX1 U507 ( .A(net14103), .Z(n419) );
  CNR2X1 U508 ( .A(n418), .B(n419), .Z(n420) );
  CIVX2 U509 ( .A(n424), .Z(net16921) );
  CIVX2 U510 ( .A(net13425), .Z(n423) );
  CND2X1 U511 ( .A(cmd0[0]), .B(n426), .Z(net13425) );
  CNR3XL U512 ( .A(net6623), .B(n426), .C(n425), .Z(_pushout_d) );
  CND2X1 U513 ( .A(n426), .B(n425), .Z(net13427) );
  CND2X1 U514 ( .A(cmd0[1]), .B(n425), .Z(net13426) );
  CANR2XL U515 ( .A(N68), .B(net16919), .C(N325), .D(net16920), .Z(net14040)
         );
  CAN2X1 U516 ( .A(net14118), .B(push0), .Z(net16919) );
  CIVX2 U517 ( .A(net13427), .Z(net14118) );
  CAN2X1 U518 ( .A(net14116), .B(push0), .Z(net16920) );
  CIVX2 U519 ( .A(net13426), .Z(net14116) );
  CANR2XL U520 ( .A(N76), .B(net16919), .C(N333), .D(net16920), .Z(net14103)
         );
  CANR2XL U521 ( .A(N66), .B(net16919), .C(N323), .D(net16920), .Z(net14022)
         );
  CIVX2 U522 ( .A(net14111), .Z(n431) );
  CIVX2 U523 ( .A(net14094), .Z(n433) );
  CIVX2 U524 ( .A(n434), .Z(n432) );
  CNR2XL U525 ( .A(n430), .B(n429), .Z(n147) );
  CIVX2 U526 ( .A(n327), .Z(net14094) );
  CND2XL U527 ( .A(n598), .B(n597), .Z(n162) );
  CIVXL U528 ( .A(n329), .Z(n435) );
  CIVXL U529 ( .A(n435), .Z(n436) );
  CIVX8 U530 ( .A(n503), .Z(n502) );
  CANR2XL U531 ( .A(N160), .B(net16921), .C(net16919), .D(N32), .Z(n864) );
  CANR2XL U532 ( .A(N161), .B(net16921), .C(N33), .D(net16919), .Z(n856) );
  CDLY1XL U533 ( .A(q0[29]), .Z(n437) );
  CMX2XL U534 ( .A0(n311), .A1(q[2]), .S(n510), .Z(n245) );
  CMX2XL U535 ( .A0(q0[28]), .A1(q[28]), .S(n508), .Z(n271) );
  CANR2XL U536 ( .A(N180), .B(net16921), .C(N52), .D(net16919), .Z(n688) );
  CDLY1XL U537 ( .A(q0[5]), .Z(n438) );
  CANR2XL U538 ( .A(N185), .B(net16921), .C(net16919), .D(N57), .Z(n648) );
  CANR2XL U539 ( .A(N174), .B(net16921), .C(N46), .D(net16919), .Z(n738) );
  CND2XL U540 ( .A(n622), .B(n621), .Z(n165) );
  CND2XL U541 ( .A(n640), .B(n639), .Z(n167) );
  CDLY1XL U542 ( .A(q0[14]), .Z(n439) );
  CMX2XL U543 ( .A0(h0[29]), .A1(h[29]), .S(n510), .Z(n240) );
  CMX2XL U544 ( .A0(h0[14]), .A1(h[14]), .S(n512), .Z(n225) );
  CDLY1XL U545 ( .A(q0[3]), .Z(n440) );
  CANR2XL U546 ( .A(net16921), .B(N191), .C(net16919), .D(N63), .Z(n598) );
  CMX2XL U547 ( .A0(q0[4]), .A1(q[4]), .S(n510), .Z(n247) );
  CDLY1XL U548 ( .A(q0[21]), .Z(n441) );
  CMX2XL U549 ( .A0(n439), .A1(q[14]), .S(n509), .Z(n257) );
  CIVXL U550 ( .A(h0[4]), .Z(n504) );
  CMX2XL U551 ( .A0(h0[9]), .A1(h[9]), .S(n512), .Z(n220) );
  CIVXL U552 ( .A(N65), .Z(n445) );
  CND2XL U553 ( .A(n632), .B(n631), .Z(n166) );
  CANR2XL U554 ( .A(N187), .B(net16921), .C(N59), .D(net16919), .Z(n632) );
  CMX2XL U555 ( .A0(h0[11]), .A1(h[11]), .S(n512), .Z(n222) );
  CANR2XL U556 ( .A(N164), .B(net16921), .C(net16919), .D(N36), .Z(n831) );
  CDLY1XL U557 ( .A(h0[22]), .Z(n446) );
  CMX2XL U558 ( .A0(n332), .A1(q[24]), .S(n508), .Z(n267) );
  CMX2XL U559 ( .A0(h0[10]), .A1(h[10]), .S(n512), .Z(n221) );
  CDLY1XL U560 ( .A(q0[7]), .Z(n490) );
  CDLY1XL U561 ( .A(q0[19]), .Z(n489) );
  CMX2XL U562 ( .A0(h0[20]), .A1(h[20]), .S(n511), .Z(n231) );
  CND2XL U563 ( .A(n680), .B(n679), .Z(n172) );
  CANR2XL U564 ( .A(N71), .B(net16919), .C(N328), .D(net16920), .Z(n546) );
  CMX2XL U565 ( .A0(h0[12]), .A1(h[12]), .S(n512), .Z(n223) );
  CDLY1XL U566 ( .A(q0[23]), .Z(n447) );
  CDLY1XL U567 ( .A(q0[11]), .Z(n487) );
  CMX2XL U568 ( .A0(n437), .A1(q[29]), .S(n508), .Z(n272) );
  CMX2XL U569 ( .A0(n442), .A1(h[4]), .S(n512), .Z(n215) );
  CMXI2XL U570 ( .A0(n1092), .A1(n1091), .S(n443), .Z(n1093) );
  COND2XL U571 ( .A(n442), .B(n745), .C(n630), .D(n612), .Z(n886) );
  CMXI2XL U572 ( .A0(n478), .A1(n837), .S(n442), .Z(n1010) );
  CMXI2XL U573 ( .A0(n481), .A1(n467), .S(n442), .Z(n933) );
  COND2XL U574 ( .A(n442), .B(n757), .C(n630), .D(n620), .Z(n901) );
  COND2XL U575 ( .A(n444), .B(n768), .C(n630), .D(n629), .Z(n913) );
  CMXI2XL U576 ( .A0(n474), .A1(n459), .S(n443), .Z(n977) );
  CND2XL U577 ( .A(n442), .B(n877), .Z(n630) );
  CIVDXL U578 ( .A(h0[4]), .Z0(n507), .Z1(n442) );
  CANR2XL U579 ( .A(n1081), .B(n1080), .C(n443), .D(n468), .Z(n1082) );
  CIVDXL U580 ( .A(h0[4]), .Z0(n506), .Z1(n443) );
  CIVDXL U581 ( .A(h0[4]), .Z0(n505), .Z1(n444) );
  CDLY1XL U582 ( .A(q0[15]), .Z(n486) );
  CANR2XL U583 ( .A(net16919), .B(N74), .C(N331), .D(net16920), .Z(n529) );
  CANR2XL U584 ( .A(N188), .B(net16921), .C(net16919), .D(N60), .Z(n622) );
  CDLY1XL U585 ( .A(q0[9]), .Z(n488) );
  CIVX3 U586 ( .A(h0[2]), .Z(n503) );
  CDLY1XL U587 ( .A(q0[13]), .Z(n452) );
  CMX2XL U588 ( .A0(n310), .A1(h[0]), .S(n513), .Z(n211) );
  CMXI2XL U589 ( .A0(net14094), .A1(n1097), .S(n310), .Z(n514) );
  CND2XL U590 ( .A(n310), .B(n519), .Z(n1071) );
  CND2XL U591 ( .A(n519), .B(n336), .Z(n518) );
  CND2XL U592 ( .A(n656), .B(n655), .Z(n169) );
  CANR2XL U593 ( .A(N184), .B(net16921), .C(net16919), .D(N56), .Z(n656) );
  CND2XL U594 ( .A(n580), .B(n503), .Z(n571) );
  CND2XL U595 ( .A(h0[3]), .B(n503), .Z(n581) );
  CND2XL U596 ( .A(n502), .B(h0[3]), .Z(n582) );
  CND2XL U597 ( .A(n614), .B(n613), .Z(n164) );
  CANR2XL U598 ( .A(N189), .B(net16921), .C(net16919), .D(N61), .Z(n614) );
  COAN1XL U599 ( .A(push0), .B(n554), .C(n535), .Z(n453) );
  CND2X1 U600 ( .A(n534), .B(n453), .Z(n152) );
  CANR2XL U601 ( .A(net16919), .B(N73), .C(N330), .D(net16920), .Z(n535) );
  COAN1XL U602 ( .A(push0), .B(n592), .C(n575), .Z(n454) );
  CND2XL U603 ( .A(n574), .B(n454), .Z(n158) );
  CIVX1 U604 ( .A(acc[51]), .Z(n592) );
  CANR2XL U605 ( .A(N67), .B(net16919), .C(N324), .D(net16920), .Z(n575) );
  CANR2XL U606 ( .A(N69), .B(net16919), .C(N326), .D(net16920), .Z(n561) );
  CIVX1 U607 ( .A(acc[59]), .Z(n541) );
  CANR2XL U608 ( .A(N75), .B(net16919), .C(N332), .D(net16920), .Z(n524) );
  CANR2XL U609 ( .A(net16919), .B(N72), .C(N329), .D(net16920), .Z(n540) );
  CIVX1 U610 ( .A(n344), .Z(n1097) );
  CANR2XL U611 ( .A(N79), .B(net16919), .C(N336), .D(net16920), .Z(n1096) );
  CMX2XL U612 ( .A0(h0[30]), .A1(h[30]), .S(n510), .Z(n241) );
  CND2XL U613 ( .A(N195), .B(net16921), .Z(n574) );
  CND2XL U614 ( .A(N197), .B(net16921), .Z(n560) );
  CND2XL U615 ( .A(N203), .B(net16921), .Z(n523) );
  CND2XL U616 ( .A(N200), .B(net16921), .Z(n539) );
  CND2XL U617 ( .A(N207), .B(net16921), .Z(n1095) );
  CMX2XL U618 ( .A0(h0[31]), .A1(h[31]), .S(n510), .Z(n242) );
  CMX2XL U619 ( .A0(h0[6]), .A1(h[6]), .S(n512), .Z(n217) );
  CIVXL U620 ( .A(h0[6]), .Z(n735) );
  CAN3XL U621 ( .A(h0[6]), .B(n466), .C(n1089), .Z(n1092) );
  CANR2XL U622 ( .A(net16919), .B(N70), .C(N327), .D(net16920), .Z(n553) );
  CMX2XL U623 ( .A0(h0[1]), .A1(h[1]), .S(n513), .Z(n212) );
  CANR2XL U624 ( .A(n310), .B(net14094), .C(h0[1]), .D(n1097), .Z(n517) );
  CND2XL U625 ( .A(h0[1]), .B(n310), .Z(n520) );
  CIVXL U626 ( .A(h0[1]), .Z(n519) );
  CND2XL U627 ( .A(h0[1]), .B(n336), .Z(n1072) );
  CNR2IXL U628 ( .B(n1087), .A(n883), .Z(N256) );
  CNR2IXL U629 ( .B(n1087), .A(n944), .Z(N251) );
  CNR2IXL U630 ( .B(n1087), .A(n955), .Z(N250) );
  CNR2IXL U631 ( .B(n1087), .A(n966), .Z(N249) );
  CNR2IXL U632 ( .B(n1087), .A(n999), .Z(N246) );
  CNR2IXL U633 ( .B(n1087), .A(n988), .Z(N247) );
  CANR2XL U634 ( .A(n888), .B(n660), .C(n877), .D(n765), .Z(n661) );
  CAN2XL U635 ( .A(n662), .B(n661), .Z(n475) );
  CANR2XL U636 ( .A(n888), .B(n684), .C(n877), .D(n792), .Z(n685) );
  CAN2XL U637 ( .A(n686), .B(n685), .Z(n473) );
  CNR2IX1 U638 ( .B(n1087), .A(n933), .Z(N252) );
  CIVX1 U639 ( .A(n757), .Z(n758) );
  COND1X1 U640 ( .A(n883), .B(n1069), .C(n882), .Z(N224) );
  CAN2XL U641 ( .A(n484), .B(n580), .Z(n467) );
  CANR2XL U642 ( .A(n888), .B(n668), .C(n877), .D(n776), .Z(n669) );
  CAN2XL U643 ( .A(n670), .B(n669), .Z(n474) );
  CNR2IX1 U644 ( .B(n1087), .A(n977), .Z(N248) );
  CNR2IX1 U645 ( .B(n1087), .A(n1035), .Z(N243) );
  CNR2IX1 U646 ( .B(n1087), .A(n1010), .Z(N245) );
  COND1XL U647 ( .A(n1040), .B(n871), .C(n862), .Z(N226) );
  COND1XL U648 ( .A(n905), .B(n871), .C(n760), .Z(N238) );
  CAN2X1 U649 ( .A(n483), .B(n580), .Z(n466) );
  COAN1X1 U650 ( .A(n484), .B(n580), .C(n579), .Z(n460) );
  COAN1X1 U651 ( .A(n483), .B(n580), .C(n551), .Z(n459) );
  CAN2X1 U652 ( .A(n544), .B(n580), .Z(n463) );
  CAN2X1 U653 ( .A(n533), .B(n580), .Z(n461) );
  CAN2X1 U654 ( .A(n538), .B(n580), .Z(n462) );
  CANR2X1 U655 ( .A(n888), .B(n716), .C(n877), .D(n825), .Z(n717) );
  CAN2XL U656 ( .A(n702), .B(n701), .Z(n477) );
  CANR2X1 U657 ( .A(n888), .B(n708), .C(n877), .D(n816), .Z(n709) );
  CAN2XL U658 ( .A(n638), .B(n637), .Z(n481) );
  CAN2XL U659 ( .A(n654), .B(n653), .Z(n472) );
  CAN2XL U660 ( .A(n678), .B(n677), .Z(n476) );
  CAN2XL U661 ( .A(n646), .B(n645), .Z(n471) );
  CAN2XL U662 ( .A(n694), .B(n693), .Z(n478) );
  CANR2XL U663 ( .A(N186), .B(net16921), .C(net16919), .D(N58), .Z(n640) );
  CNR2IX1 U664 ( .B(n1087), .A(n1070), .Z(N241) );
  CAN2XL U665 ( .A(n881), .B(n877), .Z(n455) );
  CAN2XL U666 ( .A(n455), .B(n747), .Z(N271) );
  COND1X1 U667 ( .A(n874), .B(n871), .C(n736), .Z(N240) );
  CIVXL U668 ( .A(n768), .Z(n769) );
  CIVXL U669 ( .A(n745), .Z(n746) );
  CAN2X2 U670 ( .A(n1090), .B(n505), .Z(n458) );
  CIVX4 U671 ( .A(n547), .Z(n892) );
  CANR2XL U672 ( .A(n888), .B(n700), .C(n877), .D(n808), .Z(n701) );
  CANR2XL U673 ( .A(n888), .B(n652), .C(n877), .D(n754), .Z(n653) );
  CANR2XL U674 ( .A(n888), .B(n644), .C(n877), .D(n742), .Z(n645) );
  CANR2XL U675 ( .A(n888), .B(n636), .C(n877), .D(n732), .Z(n637) );
  CANR2XL U676 ( .A(n888), .B(n676), .C(n877), .D(n784), .Z(n677) );
  CANR2XL U677 ( .A(n888), .B(n692), .C(n877), .D(n800), .Z(n693) );
  CMX2XL U678 ( .A0(n527), .A1(n485), .S(n502), .Z(n484) );
  CANR2XL U679 ( .A(N176), .B(net16921), .C(net16919), .D(N48), .Z(n720) );
  CANR2XL U680 ( .A(N175), .B(net16921), .C(N47), .D(net16919), .Z(n728) );
  CANR2XL U681 ( .A(N173), .B(net16921), .C(net16919), .D(N45), .Z(n750) );
  CANR2XL U682 ( .A(N172), .B(net16921), .C(net16919), .D(N44), .Z(n762) );
  CANR2XL U683 ( .A(N182), .B(net16921), .C(net16919), .D(N54), .Z(n672) );
  CANR2XL U684 ( .A(N181), .B(net16921), .C(N53), .D(net16919), .Z(n680) );
  CANR2XL U685 ( .A(N179), .B(net16921), .C(N51), .D(net16919), .Z(n696) );
  CANR2XL U686 ( .A(net16921), .B(N178), .C(N50), .D(net16919), .Z(n704) );
  CANR2XL U687 ( .A(N171), .B(net16921), .C(N43), .D(net16919), .Z(n773) );
  CANR2XL U688 ( .A(N170), .B(net16921), .C(net16919), .D(N42), .Z(n781) );
  CANR2XL U689 ( .A(N177), .B(net16921), .C(N49), .D(net16919), .Z(n712) );
  CANR2XL U690 ( .A(N169), .B(net16921), .C(N41), .D(net16919), .Z(n789) );
  CANR2XL U691 ( .A(N165), .B(net16921), .C(N37), .D(net16919), .Z(n822) );
  CANR2XL U692 ( .A(N163), .B(net16921), .C(net16919), .D(N35), .Z(n840) );
  CANR2XL U693 ( .A(N159), .B(net16921), .C(N31), .D(net16919), .Z(n873) );
  CANR2XL U694 ( .A(N158), .B(net16921), .C(N30), .D(net16919), .Z(n885) );
  CANR2XL U695 ( .A(N157), .B(net16921), .C(N29), .D(net16919), .Z(n900) );
  CANR2XL U696 ( .A(N156), .B(net16921), .C(N28), .D(net16919), .Z(n912) );
  CANR2XL U697 ( .A(N155), .B(net16921), .C(N27), .D(net16919), .Z(n924) );
  CANR2XL U698 ( .A(N154), .B(net16921), .C(N26), .D(net16919), .Z(n935) );
  CANR2XL U699 ( .A(N153), .B(net16921), .C(N25), .D(net16919), .Z(n946) );
  CANR2XL U700 ( .A(N152), .B(net16921), .C(N24), .D(net16919), .Z(n957) );
  CANR2XL U701 ( .A(N275), .B(net16920), .C(acc[2]), .D(net6623), .Z(n1022) );
  CANR2XL U702 ( .A(N276), .B(net16920), .C(acc[3]), .D(net6623), .Z(n1011) );
  CANR2XL U703 ( .A(N151), .B(net16921), .C(N23), .D(net16919), .Z(n968) );
  CANR2XL U704 ( .A(N150), .B(net16921), .C(N22), .D(net16919), .Z(n979) );
  CANR2XL U705 ( .A(N149), .B(net16921), .C(N21), .D(net16919), .Z(n990) );
  CANR2XL U706 ( .A(N277), .B(net16920), .C(acc[4]), .D(net6623), .Z(n1000) );
  CANR2XL U707 ( .A(N274), .B(net16920), .C(acc[1]), .D(net6623), .Z(n1036) );
  CMX2XL U708 ( .A0(z[2]), .A1(acc[2]), .S(net16065), .Z(n278) );
  CNR2IXL U709 ( .B(n1087), .A(n1021), .Z(N244) );
  CNR2IX1 U710 ( .B(n1087), .A(n1049), .Z(N242) );
  COND1XL U711 ( .A(n972), .B(n871), .C(n811), .Z(N232) );
  COND1XL U712 ( .A(n1016), .B(n871), .C(n846), .Z(N228) );
  COND1XL U713 ( .A(n939), .B(n871), .C(n787), .Z(N235) );
  COND1XL U714 ( .A(n891), .B(n871), .C(n748), .Z(N239) );
  COND1XL U715 ( .A(n917), .B(n871), .C(n771), .Z(N237) );
  COND1XL U716 ( .A(n1026), .B(n871), .C(n854), .Z(N227) );
  COND1XL U717 ( .A(n1053), .B(n871), .C(n870), .Z(N225) );
  COND1XL U718 ( .A(n950), .B(n871), .C(n795), .Z(N234) );
  COND1XL U719 ( .A(n961), .B(n871), .C(n803), .Z(N233) );
  COND1XL U720 ( .A(n928), .B(n871), .C(n779), .Z(N236) );
  CIVX4 U721 ( .A(n518), .Z(n1056) );
  CIVX4 U722 ( .A(n1071), .Z(n1055) );
  CAN2XL U723 ( .A(n1087), .B(n442), .Z(n456) );
  CIVX2 U724 ( .A(n1052), .Z(n1081) );
  CIVX2 U725 ( .A(n1067), .Z(n1087) );
  CIVX2 U726 ( .A(n871), .Z(n881) );
  CND2IX1 U727 ( .B(n1057), .A(n1058), .Z(n1059) );
  CND2IX1 U728 ( .B(n1027), .A(n1058), .Z(n1028) );
  CND2IX1 U729 ( .B(n1041), .A(n1058), .Z(n1042) );
  CAN2XL U730 ( .A(n1073), .B(n1090), .Z(n457) );
  COND1XL U731 ( .A(n994), .B(n871), .C(n829), .Z(N230) );
  CND2XL U732 ( .A(n1087), .B(n507), .Z(n871) );
  COND1XL U733 ( .A(n983), .B(n871), .C(n820), .Z(N231) );
  COND1XL U734 ( .A(n1005), .B(n871), .C(n838), .Z(N229) );
  CIVX4 U735 ( .A(n1072), .Z(n1054) );
  CIVX4 U736 ( .A(n520), .Z(n1075) );
  CND2X1 U737 ( .A(n893), .B(n507), .Z(n1077) );
  CND2X1 U738 ( .A(n892), .B(n506), .Z(n1084) );
  CAN2X1 U739 ( .A(n590), .B(n589), .Z(n464) );
  CAN2X1 U740 ( .A(n596), .B(n595), .Z(n465) );
  CAN2X1 U741 ( .A(n880), .B(n879), .Z(n468) );
  CAN2X1 U742 ( .A(n586), .B(n585), .Z(n469) );
  CAN2X1 U743 ( .A(n603), .B(n602), .Z(n470) );
  CAN2X1 U744 ( .A(n718), .B(n717), .Z(n479) );
  CAN2X1 U745 ( .A(n726), .B(n725), .Z(n480) );
  CAN2X1 U746 ( .A(n710), .B(n709), .Z(n482) );
  CAN2XL U747 ( .A(n485), .B(n503), .Z(n483) );
  CNIVX1 U748 ( .A(n1162), .Z(n498) );
  CNIVX1 U749 ( .A(n1162), .Z(n499) );
  CNIVX1 U750 ( .A(n1162), .Z(n500) );
  CNIVX1 U751 ( .A(n1162), .Z(n501) );
  CNIVX1 U752 ( .A(n1162), .Z(n496) );
  CNIVX1 U753 ( .A(n1162), .Z(n495) );
  CNIVX1 U754 ( .A(n1162), .Z(n494) );
  CNIVX1 U755 ( .A(n1162), .Z(n491) );
  CNIVX1 U756 ( .A(n1162), .Z(n492) );
  CNIVX1 U757 ( .A(n1162), .Z(n493) );
  CNIVX1 U758 ( .A(n1162), .Z(n497) );
  CND2XL U759 ( .A(h0[5]), .B(n735), .Z(n1069) );
  CNIVX1 U760 ( .A(pushin), .Z(n513) );
  CIVXL U761 ( .A(h0[3]), .Z(n580) );
  CAN2XL U762 ( .A(n1056), .B(n345), .Z(n485) );
  CIVX2 U763 ( .A(push0), .Z(net6623) );
  CNIVX1 U764 ( .A(pushin), .Z(n512) );
  CNIVX1 U765 ( .A(pushin), .Z(n511) );
  CNIVX1 U766 ( .A(pushin), .Z(n510) );
  CNIVX1 U767 ( .A(pushin), .Z(n508) );
  CNIVX1 U768 ( .A(pushin), .Z(n509) );
  CNIVX1 U769 ( .A(net13361), .Z(net16065) );
  CIVX2 U770 ( .A(rst), .Z(n1162) );
  CMX2XL U771 ( .A0(n441), .A1(q[21]), .S(n508), .Z(n264) );
  CMX2XL U772 ( .A0(n447), .A1(q[23]), .S(n508), .Z(n266) );
  CMX2XL U773 ( .A0(n486), .A1(q[15]), .S(n509), .Z(n258) );
  CMX2XL U774 ( .A0(n487), .A1(q[11]), .S(n509), .Z(n254) );
  CMX2XL U775 ( .A0(n488), .A1(q[9]), .S(n509), .Z(n252) );
  CMX2XL U776 ( .A0(n438), .A1(q[5]), .S(n510), .Z(n248) );
  CMX2XL U777 ( .A0(q0[25]), .A1(q[25]), .S(n508), .Z(n268) );
  CMX2XL U778 ( .A0(n324), .A1(q[27]), .S(n508), .Z(n270) );
  CMX2XL U779 ( .A0(n309), .A1(q[17]), .S(n509), .Z(n260) );
  CMX2XL U780 ( .A0(n452), .A1(q[13]), .S(n509), .Z(n256) );
  CMX2XL U781 ( .A0(n490), .A1(q[7]), .S(n510), .Z(n250) );
  CMX2XL U782 ( .A0(n440), .A1(q[3]), .S(n510), .Z(n246) );
  CMX2XL U783 ( .A0(q0[1]), .A1(q[1]), .S(n510), .Z(n244) );
  CMX2X1 U784 ( .A0(q0[20]), .A1(q[20]), .S(n508), .Z(n263) );
  CMX2X1 U785 ( .A0(n489), .A1(q[19]), .S(n509), .Z(n262) );
  CMX2X1 U786 ( .A0(q0[12]), .A1(q[12]), .S(n509), .Z(n255) );
  CMX2X1 U787 ( .A0(q0[10]), .A1(q[10]), .S(n509), .Z(n253) );
  CMX2X1 U788 ( .A0(q0[0]), .A1(q[0]), .S(n510), .Z(n243) );
  CMX2X1 U789 ( .A0(h0[28]), .A1(h[28]), .S(n510), .Z(n239) );
  CMX2X1 U790 ( .A0(h0[27]), .A1(h[27]), .S(n511), .Z(n238) );
  CMX2X1 U791 ( .A0(h0[25]), .A1(h[25]), .S(n511), .Z(n236) );
  CMX2X1 U792 ( .A0(h0[24]), .A1(h[24]), .S(n511), .Z(n235) );
  CMX2X1 U793 ( .A0(h0[23]), .A1(h[23]), .S(n511), .Z(n234) );
  CMX2X1 U794 ( .A0(n446), .A1(h[22]), .S(n511), .Z(n233) );
  CMX2X1 U795 ( .A0(h0[21]), .A1(h[21]), .S(n511), .Z(n232) );
  CMX2X1 U796 ( .A0(h0[19]), .A1(h[19]), .S(n511), .Z(n230) );
  CMX2X1 U797 ( .A0(h0[18]), .A1(h[18]), .S(n511), .Z(n229) );
  CMX2X1 U798 ( .A0(h0[17]), .A1(h[17]), .S(n511), .Z(n228) );
  CMX2X1 U799 ( .A0(h0[16]), .A1(h[16]), .S(n511), .Z(n227) );
  CMX2X1 U800 ( .A0(h0[15]), .A1(h[15]), .S(n512), .Z(n226) );
  CMX2X1 U801 ( .A0(h0[13]), .A1(h[13]), .S(n512), .Z(n224) );
  CMX2X1 U802 ( .A0(h0[8]), .A1(h[8]), .S(n512), .Z(n219) );
  CMX2X1 U803 ( .A0(h0[7]), .A1(h[7]), .S(n512), .Z(n218) );
  CMX2X1 U804 ( .A0(n502), .A1(h[2]), .S(n513), .Z(n213) );
  CIVX2 U805 ( .A(h0[5]), .Z(n1089) );
  CAN2X1 U806 ( .A(n881), .B(n466), .Z(N272) );
  CND2X1 U807 ( .A(n514), .B(n519), .Z(n612) );
  CIVX2 U808 ( .A(n612), .Z(n747) );
  COND3X1 U809 ( .A(n451), .B(n518), .C(n520), .D(n517), .Z(n620) );
  CIVX2 U810 ( .A(n620), .Z(n759) );
  CAN2X1 U811 ( .A(n455), .B(n759), .Z(N270) );
  CANR2X1 U812 ( .A(n1055), .B(n530), .C(n1054), .D(net14094), .Z(n522) );
  CANR2X1 U813 ( .A(n1075), .B(n1097), .C(n1056), .D(net14078), .Z(n521) );
  CND2X1 U814 ( .A(n522), .B(n521), .Z(n629) );
  CIVX2 U815 ( .A(n629), .Z(n770) );
  CAN2X1 U816 ( .A(n455), .B(n770), .Z(N269) );
  CANR2X1 U817 ( .A(n1055), .B(net14078), .C(n1054), .D(n530), .Z(n526) );
  CANR2X1 U818 ( .A(n1075), .B(net14094), .C(n1056), .D(n541), .Z(n525) );
  CND2X1 U819 ( .A(n526), .B(n525), .Z(n601) );
  CIVX2 U820 ( .A(n601), .Z(n527) );
  CAN2X1 U821 ( .A(n467), .B(n881), .Z(N268) );
  CANR2X1 U822 ( .A(n1055), .B(n541), .C(n1054), .D(net14078), .Z(n532) );
  CANR2X1 U823 ( .A(n1075), .B(n530), .C(n1056), .D(n548), .Z(n531) );
  CND2X1 U824 ( .A(n532), .B(n531), .Z(n609) );
  CMXI2X1 U825 ( .A0(n609), .A1(n612), .S(n502), .Z(n533) );
  CAN2X1 U826 ( .A(n461), .B(n881), .Z(N267) );
  CIVX2 U827 ( .A(acc[57]), .Z(n554) );
  CND2X1 U828 ( .A(N201), .B(net16921), .Z(n534) );
  CANR2X1 U829 ( .A(n1055), .B(n548), .C(n1054), .D(n541), .Z(n537) );
  CANR2X1 U830 ( .A(n1075), .B(net14078), .C(n1056), .D(n554), .Z(n536) );
  CND2X1 U831 ( .A(n537), .B(n536), .Z(n617) );
  CMXI2X1 U832 ( .A0(n617), .A1(n620), .S(n502), .Z(n538) );
  CAN2X1 U833 ( .A(n462), .B(n881), .Z(N266) );
  CANR2X1 U834 ( .A(n1055), .B(n554), .C(n1054), .D(n548), .Z(n543) );
  CANR2X1 U835 ( .A(n1075), .B(n541), .C(n1056), .D(n339), .Z(n542) );
  CND2X1 U836 ( .A(n543), .B(n542), .Z(n626) );
  CMXI2X1 U837 ( .A0(n626), .A1(n629), .S(n502), .Z(n544) );
  CAN2X1 U838 ( .A(n463), .B(n881), .Z(N265) );
  CND2X1 U839 ( .A(n502), .B(n580), .Z(n547) );
  CANR2X1 U840 ( .A(n1055), .B(n339), .C(n1054), .D(n554), .Z(n550) );
  CANR2X1 U841 ( .A(n1075), .B(n548), .C(n1056), .D(n567), .Z(n549) );
  CND2X1 U842 ( .A(n550), .B(n549), .Z(n636) );
  CANR2X1 U843 ( .A(n892), .B(n601), .C(n877), .D(n636), .Z(n551) );
  CAN2X1 U844 ( .A(n459), .B(n881), .Z(N264) );
  CANR2X1 U845 ( .A(n1055), .B(n567), .C(n1054), .D(n339), .Z(n556) );
  CANR2X1 U846 ( .A(n1075), .B(n554), .C(n1056), .D(n576), .Z(n555) );
  CND2X1 U847 ( .A(n556), .B(n555), .Z(n644) );
  CIVX2 U848 ( .A(n644), .Z(n558) );
  COND3X1 U849 ( .A(n558), .B(n571), .C(n582), .D(n557), .Z(n559) );
  CIVX2 U850 ( .A(n559), .Z(n819) );
  CAN2X1 U851 ( .A(n819), .B(n881), .Z(N263) );
  CANR2X1 U852 ( .A(n1055), .B(n576), .C(n1054), .D(n567), .Z(n563) );
  CANR2X1 U853 ( .A(n1075), .B(n339), .C(n1056), .D(n341), .Z(n562) );
  CND2X1 U854 ( .A(n563), .B(n562), .Z(n652) );
  CIVX2 U855 ( .A(n652), .Z(n565) );
  COND3X1 U856 ( .A(n565), .B(n571), .C(n582), .D(n564), .Z(n566) );
  CIVX2 U857 ( .A(n566), .Z(n828) );
  CAN2X1 U858 ( .A(n828), .B(n881), .Z(N262) );
  CANR2X1 U859 ( .A(n1055), .B(n341), .C(n1054), .D(n576), .Z(n569) );
  CANR2X1 U860 ( .A(n1075), .B(n567), .C(n1056), .D(net14010), .Z(n568) );
  CND2X1 U861 ( .A(n569), .B(n568), .Z(n660) );
  CIVX2 U862 ( .A(n660), .Z(n572) );
  COND3X1 U863 ( .A(n572), .B(n571), .C(n582), .D(n570), .Z(n573) );
  CIVX2 U864 ( .A(n573), .Z(n837) );
  CAN2X1 U865 ( .A(n837), .B(n881), .Z(N261) );
  CANR2X1 U866 ( .A(n1055), .B(net14010), .C(n1054), .D(n341), .Z(n578) );
  CANR2X1 U867 ( .A(n1075), .B(n576), .C(n1056), .D(n592), .Z(n577) );
  CND2X1 U868 ( .A(n578), .B(n577), .Z(n668) );
  CANR2X1 U869 ( .A(n892), .B(n636), .C(n877), .D(n668), .Z(n579) );
  CAN2X1 U870 ( .A(n460), .B(n881), .Z(N260) );
  CANR2X1 U871 ( .A(n893), .B(n609), .C(n892), .D(n644), .Z(n586) );
  CANR2X1 U872 ( .A(n1055), .B(n592), .C(n1054), .D(net14010), .Z(n584) );
  CANR2X1 U873 ( .A(n1075), .B(n341), .C(n1056), .D(net13994), .Z(n583) );
  CND2X1 U874 ( .A(n584), .B(n583), .Z(n676) );
  CANR2X1 U875 ( .A(n888), .B(n612), .C(n877), .D(n676), .Z(n585) );
  CAN2X1 U876 ( .A(n469), .B(n881), .Z(N259) );
  CANR2X1 U877 ( .A(n893), .B(n617), .C(n892), .D(n652), .Z(n590) );
  CANR2X1 U878 ( .A(n1055), .B(net13994), .C(n1054), .D(n592), .Z(n588) );
  CIVX2 U879 ( .A(acc[49]), .Z(n606) );
  CANR2X1 U880 ( .A(n1075), .B(net14010), .C(n1056), .D(n606), .Z(n587) );
  CND2X1 U881 ( .A(n588), .B(n587), .Z(n684) );
  CANR2X1 U882 ( .A(n888), .B(n620), .C(n877), .D(n684), .Z(n589) );
  CAN2X1 U883 ( .A(n464), .B(n881), .Z(N258) );
  CANR2X1 U884 ( .A(N192), .B(net16921), .C(n436), .D(net16919), .Z(n591) );
  CANR2X1 U885 ( .A(n893), .B(n626), .C(n892), .D(n660), .Z(n596) );
  CANR2X1 U886 ( .A(n1055), .B(n606), .C(n1054), .D(net13994), .Z(n594) );
  CANR2X1 U887 ( .A(n1075), .B(n592), .C(n1056), .D(n334), .Z(n593) );
  CND2X1 U888 ( .A(n594), .B(n593), .Z(n692) );
  CANR2X1 U889 ( .A(n888), .B(n629), .C(n877), .D(n692), .Z(n595) );
  CAN2X1 U890 ( .A(n465), .B(n881), .Z(N257) );
  CANR2X1 U891 ( .A(N320), .B(net16920), .C(acc[47]), .D(net6623), .Z(n597) );
  CANR2X1 U892 ( .A(n893), .B(n636), .C(n892), .D(n668), .Z(n603) );
  CANR2X1 U893 ( .A(n1055), .B(n334), .C(n1054), .D(n606), .Z(n600) );
  CIVX2 U894 ( .A(acc[47]), .Z(n623) );
  CANR2X1 U895 ( .A(n1075), .B(net13994), .C(n1056), .D(n623), .Z(n599) );
  CND2X1 U896 ( .A(n600), .B(n599), .Z(n700) );
  CANR2X1 U897 ( .A(n888), .B(n601), .C(n877), .D(n700), .Z(n602) );
  CMXI2X1 U898 ( .A0(n470), .A1(n466), .S(n442), .Z(n883) );
  CANR2X1 U899 ( .A(N319), .B(net16920), .C(acc[46]), .D(net6623), .Z(n604) );
  CANR2X1 U900 ( .A(n893), .B(n644), .C(n892), .D(n676), .Z(n611) );
  CANR2X1 U901 ( .A(n1055), .B(n623), .C(n1054), .D(n334), .Z(n608) );
  CIVX2 U902 ( .A(acc[46]), .Z(n633) );
  CANR2X1 U903 ( .A(n1075), .B(n606), .C(n1056), .D(n633), .Z(n607) );
  CND2X1 U904 ( .A(n608), .B(n607), .Z(n708) );
  CANR2X1 U905 ( .A(n888), .B(n609), .C(n877), .D(n708), .Z(n610) );
  CND2X1 U906 ( .A(n611), .B(n610), .Z(n745) );
  CAN2X1 U907 ( .A(n1087), .B(n886), .Z(N255) );
  CANR2X1 U908 ( .A(N318), .B(net16920), .C(acc[45]), .D(net6623), .Z(n613) );
  CANR2X1 U909 ( .A(n893), .B(n652), .C(n892), .D(n684), .Z(n619) );
  CANR2X1 U910 ( .A(n1055), .B(n633), .C(n1054), .D(n623), .Z(n616) );
  CIVX2 U911 ( .A(acc[45]), .Z(n641) );
  CANR2X1 U912 ( .A(n1075), .B(n334), .C(n1056), .D(n641), .Z(n615) );
  CND2X1 U913 ( .A(n616), .B(n615), .Z(n716) );
  CANR2X1 U914 ( .A(n888), .B(n617), .C(n877), .D(n716), .Z(n618) );
  CND2X1 U915 ( .A(n619), .B(n618), .Z(n757) );
  CAN2X1 U916 ( .A(n1087), .B(n901), .Z(N254) );
  CANR2X1 U917 ( .A(N317), .B(net16920), .C(acc[44]), .D(net6623), .Z(n621) );
  CANR2X1 U918 ( .A(n893), .B(n660), .C(n892), .D(n692), .Z(n628) );
  CANR2X1 U919 ( .A(n1055), .B(n641), .C(n1054), .D(n633), .Z(n625) );
  CIVX2 U920 ( .A(acc[44]), .Z(n649) );
  CANR2X1 U921 ( .A(n1075), .B(n623), .C(n1056), .D(n649), .Z(n624) );
  CND2X1 U922 ( .A(n625), .B(n624), .Z(n724) );
  CANR2X1 U923 ( .A(n888), .B(n626), .C(n877), .D(n724), .Z(n627) );
  CND2X1 U924 ( .A(n628), .B(n627), .Z(n768) );
  CAN2X1 U925 ( .A(n1087), .B(n913), .Z(N253) );
  CANR2X1 U926 ( .A(N316), .B(net16920), .C(acc[43]), .D(net6623), .Z(n631) );
  CANR2X1 U927 ( .A(n893), .B(n668), .C(n892), .D(n700), .Z(n638) );
  CANR2X1 U928 ( .A(n1055), .B(n649), .C(n1054), .D(n641), .Z(n635) );
  CIVX2 U929 ( .A(acc[43]), .Z(n657) );
  CANR2X1 U930 ( .A(n1075), .B(n633), .C(n1056), .D(n657), .Z(n634) );
  CND2X1 U931 ( .A(n635), .B(n634), .Z(n732) );
  CANR2X1 U932 ( .A(N315), .B(net16920), .C(acc[42]), .D(net6623), .Z(n639) );
  CANR2X1 U933 ( .A(n893), .B(n676), .C(n892), .D(n708), .Z(n646) );
  CANR2X1 U934 ( .A(n1055), .B(n657), .C(n1054), .D(n649), .Z(n643) );
  CIVX2 U935 ( .A(acc[42]), .Z(n665) );
  CANR2X1 U936 ( .A(n1075), .B(n641), .C(n1056), .D(n665), .Z(n642) );
  CND2X1 U937 ( .A(n643), .B(n642), .Z(n742) );
  CMXI2X1 U938 ( .A0(n471), .A1(n461), .S(n444), .Z(n944) );
  CANR2X1 U939 ( .A(N314), .B(net16920), .C(acc[41]), .D(net6623), .Z(n647) );
  CANR2X1 U940 ( .A(n893), .B(n684), .C(n892), .D(n716), .Z(n654) );
  CANR2X1 U941 ( .A(n1055), .B(n665), .C(n1054), .D(n657), .Z(n651) );
  CIVX2 U942 ( .A(acc[41]), .Z(n673) );
  CANR2X1 U943 ( .A(n1075), .B(n649), .C(n1056), .D(n673), .Z(n650) );
  CND2X1 U944 ( .A(n651), .B(n650), .Z(n754) );
  CMXI2X1 U945 ( .A0(n472), .A1(n462), .S(n443), .Z(n955) );
  CANR2X1 U946 ( .A(N313), .B(net16920), .C(acc[40]), .D(net6623), .Z(n655) );
  CANR2X1 U947 ( .A(n893), .B(n692), .C(n892), .D(n724), .Z(n662) );
  CANR2X1 U948 ( .A(n1055), .B(n673), .C(n1054), .D(n665), .Z(n659) );
  CIVX2 U949 ( .A(acc[40]), .Z(n681) );
  CANR2X1 U950 ( .A(n1075), .B(n657), .C(n1056), .D(n681), .Z(n658) );
  CND2X1 U951 ( .A(n659), .B(n658), .Z(n765) );
  CMXI2X1 U952 ( .A0(n475), .A1(n463), .S(n444), .Z(n966) );
  CANR2X1 U953 ( .A(n893), .B(n700), .C(n892), .D(n732), .Z(n670) );
  CANR2X1 U954 ( .A(n1055), .B(n681), .C(n1054), .D(n673), .Z(n667) );
  CIVX2 U955 ( .A(acc[39]), .Z(n689) );
  CANR2X1 U956 ( .A(n1075), .B(n665), .C(n1056), .D(n689), .Z(n666) );
  CND2X1 U957 ( .A(n667), .B(n666), .Z(n776) );
  CANR2X1 U958 ( .A(n893), .B(n708), .C(n892), .D(n742), .Z(n678) );
  CANR2X1 U959 ( .A(n1055), .B(n689), .C(n1054), .D(n681), .Z(n675) );
  CIVX2 U960 ( .A(acc[38]), .Z(n697) );
  CANR2X1 U961 ( .A(n1075), .B(n673), .C(n1056), .D(n697), .Z(n674) );
  CND2X1 U962 ( .A(n675), .B(n674), .Z(n784) );
  CMXI2X1 U963 ( .A0(n476), .A1(n819), .S(n443), .Z(n988) );
  CANR2X1 U964 ( .A(N310), .B(net16920), .C(acc[37]), .D(net6623), .Z(n679) );
  CANR2X1 U965 ( .A(n893), .B(n716), .C(n892), .D(n754), .Z(n686) );
  CANR2X1 U966 ( .A(n1055), .B(n697), .C(n1054), .D(n689), .Z(n683) );
  CIVX2 U967 ( .A(acc[37]), .Z(n705) );
  CANR2X1 U968 ( .A(n1075), .B(n681), .C(n1056), .D(n705), .Z(n682) );
  CND2X1 U969 ( .A(n683), .B(n682), .Z(n792) );
  CMXI2X1 U970 ( .A0(n473), .A1(n828), .S(n444), .Z(n999) );
  CANR2X1 U971 ( .A(N309), .B(net16920), .C(acc[36]), .D(net6623), .Z(n687) );
  CANR2X1 U972 ( .A(n893), .B(n724), .C(n892), .D(n765), .Z(n694) );
  CANR2X1 U973 ( .A(n1055), .B(n705), .C(n1054), .D(n697), .Z(n691) );
  CIVX2 U974 ( .A(acc[36]), .Z(n713) );
  CANR2X1 U975 ( .A(n1075), .B(n689), .C(n1056), .D(n713), .Z(n690) );
  CND2X1 U976 ( .A(n691), .B(n690), .Z(n800) );
  CANR2X1 U977 ( .A(N308), .B(net16920), .C(acc[35]), .D(net6623), .Z(n695) );
  CANR2X1 U978 ( .A(n893), .B(n732), .C(n892), .D(n776), .Z(n702) );
  CANR2X1 U979 ( .A(n1055), .B(n713), .C(n1054), .D(n705), .Z(n699) );
  CIVX2 U980 ( .A(acc[35]), .Z(n721) );
  CANR2X1 U981 ( .A(n1075), .B(n697), .C(n1056), .D(n721), .Z(n698) );
  CND2X1 U982 ( .A(n699), .B(n698), .Z(n808) );
  CMXI2X1 U983 ( .A0(n477), .A1(n460), .S(n444), .Z(n1021) );
  CANR2X1 U984 ( .A(N307), .B(net16920), .C(acc[34]), .D(net6623), .Z(n703) );
  CANR2X1 U985 ( .A(n893), .B(n742), .C(n892), .D(n784), .Z(n710) );
  CANR2X1 U986 ( .A(n1055), .B(n721), .C(n1054), .D(n713), .Z(n707) );
  CIVX2 U987 ( .A(acc[34]), .Z(n729) );
  CANR2X1 U988 ( .A(n1075), .B(n705), .C(n1056), .D(n729), .Z(n706) );
  CND2X1 U989 ( .A(n707), .B(n706), .Z(n816) );
  CMXI2X1 U990 ( .A0(n482), .A1(n469), .S(n444), .Z(n1035) );
  CANR2X1 U991 ( .A(n893), .B(n754), .C(n892), .D(n792), .Z(n718) );
  CANR2X1 U992 ( .A(n1055), .B(n729), .C(n1054), .D(n721), .Z(n715) );
  CIVX2 U993 ( .A(acc[33]), .Z(n739) );
  CANR2X1 U994 ( .A(n1075), .B(n713), .C(n1056), .D(n739), .Z(n714) );
  CND2X1 U995 ( .A(n715), .B(n714), .Z(n825) );
  CMXI2X1 U996 ( .A0(n479), .A1(n464), .S(n443), .Z(n1049) );
  CANR2X1 U997 ( .A(N305), .B(net16920), .C(acc[32]), .D(net6623), .Z(n719) );
  CANR2X1 U998 ( .A(n893), .B(n765), .C(n892), .D(n800), .Z(n726) );
  CANR2X1 U999 ( .A(n1055), .B(n739), .C(n1054), .D(n729), .Z(n723) );
  CIVX2 U1000 ( .A(acc[32]), .Z(n751) );
  CANR2X1 U1001 ( .A(n1075), .B(n721), .C(n1056), .D(n751), .Z(n722) );
  CND2X1 U1002 ( .A(n723), .B(n722), .Z(n834) );
  CANR2X1 U1003 ( .A(n888), .B(n724), .C(n877), .D(n834), .Z(n725) );
  CMXI2X1 U1004 ( .A0(n480), .A1(n465), .S(n444), .Z(n1070) );
  CANR2X1 U1005 ( .A(N304), .B(net16920), .C(acc[31]), .D(net6623), .Z(n727)
         );
  CANR2X1 U1006 ( .A(n893), .B(n776), .C(n892), .D(n808), .Z(n734) );
  CANR2X1 U1007 ( .A(n1055), .B(n751), .C(n1054), .D(n739), .Z(n731) );
  CIVX2 U1008 ( .A(acc[31]), .Z(n1160) );
  CANR2X1 U1009 ( .A(n1075), .B(n729), .C(n1056), .D(n1160), .Z(n730) );
  CND2X1 U1010 ( .A(n731), .B(n730), .Z(n843) );
  CANR2X1 U1011 ( .A(n888), .B(n732), .C(n877), .D(n843), .Z(n733) );
  CND2X1 U1012 ( .A(n734), .B(n733), .Z(n874) );
  CIVX2 U1013 ( .A(n1069), .Z(n1090) );
  CANR2X1 U1014 ( .A(n466), .B(n458), .C(n456), .D(n470), .Z(n736) );
  CANR2X1 U1015 ( .A(N303), .B(net16920), .C(acc[30]), .D(net6623), .Z(n737)
         );
  CANR2X1 U1016 ( .A(n893), .B(n784), .C(n892), .D(n816), .Z(n744) );
  CANR2X1 U1017 ( .A(n1055), .B(n1160), .C(n1054), .D(n751), .Z(n741) );
  CIVX2 U1018 ( .A(acc[30]), .Z(n1158) );
  CANR2X1 U1019 ( .A(n1075), .B(n739), .C(n1056), .D(n1158), .Z(n740) );
  CND2X1 U1020 ( .A(n741), .B(n740), .Z(n851) );
  CANR2X1 U1021 ( .A(n888), .B(n742), .C(n877), .D(n851), .Z(n743) );
  CND2X1 U1022 ( .A(n744), .B(n743), .Z(n891) );
  CIVX2 U1023 ( .A(n1060), .Z(n1073) );
  CANR2X1 U1024 ( .A(n457), .B(n747), .C(n456), .D(n746), .Z(n748) );
  CANR2X1 U1025 ( .A(n893), .B(n792), .C(n892), .D(n825), .Z(n756) );
  CANR2X1 U1026 ( .A(n1055), .B(n1158), .C(n1054), .D(n1160), .Z(n753) );
  CIVX2 U1027 ( .A(acc[29]), .Z(n1156) );
  CANR2X1 U1028 ( .A(n1075), .B(n751), .C(n1056), .D(n1156), .Z(n752) );
  CND2X1 U1029 ( .A(n753), .B(n752), .Z(n859) );
  CANR2X1 U1030 ( .A(n888), .B(n754), .C(n877), .D(n859), .Z(n755) );
  CND2X1 U1031 ( .A(n756), .B(n755), .Z(n905) );
  CANR2X1 U1032 ( .A(n457), .B(n759), .C(n456), .D(n758), .Z(n760) );
  CANR2X1 U1033 ( .A(n893), .B(n800), .C(n892), .D(n834), .Z(n767) );
  CANR2X1 U1034 ( .A(n1055), .B(n1156), .C(n1054), .D(n1158), .Z(n764) );
  CIVX2 U1035 ( .A(acc[28]), .Z(n1154) );
  CANR2X1 U1036 ( .A(n1075), .B(n1160), .C(n1056), .D(n1154), .Z(n763) );
  CND2X1 U1037 ( .A(n764), .B(n763), .Z(n867) );
  CANR2X1 U1038 ( .A(n888), .B(n765), .C(n877), .D(n867), .Z(n766) );
  CND2X1 U1039 ( .A(n767), .B(n766), .Z(n917) );
  CANR2X1 U1040 ( .A(n457), .B(n770), .C(n456), .D(n769), .Z(n771) );
  CANR2X1 U1041 ( .A(n893), .B(n808), .C(n892), .D(n843), .Z(n778) );
  CANR2X1 U1042 ( .A(n1055), .B(n1154), .C(n1054), .D(n1156), .Z(n775) );
  CIVX2 U1043 ( .A(acc[27]), .Z(n1152) );
  CANR2X1 U1044 ( .A(n1075), .B(n1158), .C(n1056), .D(n1152), .Z(n774) );
  CND2X1 U1045 ( .A(n775), .B(n774), .Z(n878) );
  CANR2X1 U1046 ( .A(n888), .B(n776), .C(n877), .D(n878), .Z(n777) );
  CND2X1 U1047 ( .A(n778), .B(n777), .Z(n928) );
  CANR2X1 U1048 ( .A(n467), .B(n458), .C(n481), .D(n456), .Z(n779) );
  CANR2X1 U1049 ( .A(n893), .B(n816), .C(n892), .D(n851), .Z(n786) );
  CANR2X1 U1050 ( .A(n1055), .B(n1152), .C(n1054), .D(n1154), .Z(n783) );
  CIVX2 U1051 ( .A(acc[26]), .Z(n1150) );
  CANR2X1 U1052 ( .A(n1075), .B(n1156), .C(n1056), .D(n1150), .Z(n782) );
  CND2X1 U1053 ( .A(n783), .B(n782), .Z(n887) );
  CANR2X1 U1054 ( .A(n888), .B(n784), .C(n877), .D(n887), .Z(n785) );
  CND2X1 U1055 ( .A(n786), .B(n785), .Z(n939) );
  CANR2X1 U1056 ( .A(n461), .B(n458), .C(n471), .D(n456), .Z(n787) );
  CANR2X1 U1057 ( .A(N298), .B(net16920), .C(acc[25]), .D(net6623), .Z(n788)
         );
  CND2X1 U1058 ( .A(n789), .B(n788), .Z(n184) );
  CANR2X1 U1059 ( .A(n893), .B(n825), .C(n892), .D(n859), .Z(n794) );
  CANR2X1 U1060 ( .A(n1055), .B(n1150), .C(n1054), .D(n1152), .Z(n791) );
  CIVX2 U1061 ( .A(acc[25]), .Z(n1148) );
  CANR2X1 U1062 ( .A(n1075), .B(n1154), .C(n1056), .D(n1148), .Z(n790) );
  CND2X1 U1063 ( .A(n791), .B(n790), .Z(n902) );
  CANR2X1 U1064 ( .A(n888), .B(n792), .C(n877), .D(n902), .Z(n793) );
  CND2X1 U1065 ( .A(n794), .B(n793), .Z(n950) );
  CANR2X1 U1066 ( .A(n462), .B(n458), .C(n472), .D(n456), .Z(n795) );
  CANR2X1 U1067 ( .A(N297), .B(net16920), .C(acc[24]), .D(net6623), .Z(n796)
         );
  CANR2X1 U1068 ( .A(n893), .B(n834), .C(n892), .D(n867), .Z(n802) );
  CANR2X1 U1069 ( .A(n1055), .B(n1148), .C(n1054), .D(n1150), .Z(n799) );
  CIVX2 U1070 ( .A(acc[24]), .Z(n1146) );
  CANR2X1 U1071 ( .A(n1075), .B(n1152), .C(n1056), .D(n1146), .Z(n798) );
  CND2X1 U1072 ( .A(n799), .B(n798), .Z(n914) );
  CANR2X1 U1073 ( .A(n888), .B(n800), .C(n877), .D(n914), .Z(n801) );
  CND2X1 U1074 ( .A(n802), .B(n801), .Z(n961) );
  CANR2X1 U1075 ( .A(n463), .B(n458), .C(n475), .D(n456), .Z(n803) );
  CANR2X1 U1076 ( .A(N296), .B(net16920), .C(acc[23]), .D(net6623), .Z(n804)
         );
  CND2X1 U1077 ( .A(n805), .B(n804), .Z(n186) );
  CANR2X1 U1078 ( .A(n893), .B(n843), .C(n892), .D(n878), .Z(n810) );
  CANR2X1 U1079 ( .A(n1055), .B(n1146), .C(n1054), .D(n1148), .Z(n807) );
  CIVX2 U1080 ( .A(acc[23]), .Z(n1144) );
  CANR2X1 U1081 ( .A(n1075), .B(n1150), .C(n1056), .D(n1144), .Z(n806) );
  CND2X1 U1082 ( .A(n807), .B(n806), .Z(n925) );
  CANR2X1 U1083 ( .A(n888), .B(n808), .C(n877), .D(n925), .Z(n809) );
  CND2X1 U1084 ( .A(n810), .B(n809), .Z(n972) );
  CANR2X1 U1085 ( .A(n459), .B(n458), .C(n474), .D(n456), .Z(n811) );
  CANR2X1 U1086 ( .A(N166), .B(net16921), .C(N38), .D(net16919), .Z(n813) );
  CANR2X1 U1087 ( .A(N295), .B(net16920), .C(acc[22]), .D(net6623), .Z(n812)
         );
  CND2X1 U1088 ( .A(n813), .B(n812), .Z(n187) );
  CANR2X1 U1089 ( .A(n893), .B(n851), .C(n892), .D(n887), .Z(n818) );
  CANR2X1 U1090 ( .A(n1055), .B(n1144), .C(n1054), .D(n1146), .Z(n815) );
  CIVX2 U1091 ( .A(acc[22]), .Z(n1142) );
  CANR2X1 U1092 ( .A(n1075), .B(n1148), .C(n1056), .D(n1142), .Z(n814) );
  CND2X1 U1093 ( .A(n815), .B(n814), .Z(n936) );
  CANR2X1 U1094 ( .A(n888), .B(n816), .C(n877), .D(n936), .Z(n817) );
  CND2X1 U1095 ( .A(n818), .B(n817), .Z(n983) );
  CANR2X1 U1096 ( .A(n819), .B(n458), .C(n476), .D(n456), .Z(n820) );
  CANR2X1 U1097 ( .A(N294), .B(net16920), .C(acc[21]), .D(net6623), .Z(n821)
         );
  CND2X1 U1098 ( .A(n822), .B(n821), .Z(n188) );
  CANR2X1 U1099 ( .A(n893), .B(n859), .C(n892), .D(n902), .Z(n827) );
  CANR2X1 U1100 ( .A(n1055), .B(n1142), .C(n1054), .D(n1144), .Z(n824) );
  CIVX2 U1101 ( .A(acc[21]), .Z(n1140) );
  CANR2X1 U1102 ( .A(n1075), .B(n1146), .C(n1056), .D(n1140), .Z(n823) );
  CND2X1 U1103 ( .A(n824), .B(n823), .Z(n947) );
  CANR2X1 U1104 ( .A(n888), .B(n825), .C(n877), .D(n947), .Z(n826) );
  CND2X1 U1105 ( .A(n827), .B(n826), .Z(n994) );
  CANR2X1 U1106 ( .A(n828), .B(n458), .C(n473), .D(n456), .Z(n829) );
  CANR2X1 U1107 ( .A(N293), .B(net16920), .C(acc[20]), .D(net6623), .Z(n830)
         );
  CND2X1 U1108 ( .A(n831), .B(n830), .Z(n189) );
  CANR2X1 U1109 ( .A(n893), .B(n867), .C(n892), .D(n914), .Z(n836) );
  CANR2X1 U1110 ( .A(n1055), .B(n1140), .C(n1054), .D(n1142), .Z(n833) );
  CIVX2 U1111 ( .A(acc[20]), .Z(n1138) );
  CANR2X1 U1112 ( .A(n1075), .B(n1144), .C(n1056), .D(n1138), .Z(n832) );
  CND2X1 U1113 ( .A(n833), .B(n832), .Z(n958) );
  CANR2X1 U1114 ( .A(n888), .B(n834), .C(n877), .D(n958), .Z(n835) );
  CND2X1 U1115 ( .A(n836), .B(n835), .Z(n1005) );
  CANR2X1 U1116 ( .A(n837), .B(n458), .C(n478), .D(n456), .Z(n838) );
  CANR2X1 U1117 ( .A(N292), .B(net16920), .C(acc[19]), .D(net6623), .Z(n839)
         );
  CND2X1 U1118 ( .A(n840), .B(n839), .Z(n190) );
  CANR2X1 U1119 ( .A(n893), .B(n878), .C(n892), .D(n925), .Z(n845) );
  CANR2X1 U1120 ( .A(n1055), .B(n1138), .C(n1054), .D(n1140), .Z(n842) );
  CIVX2 U1121 ( .A(acc[19]), .Z(n1136) );
  CANR2X1 U1122 ( .A(n1075), .B(n1142), .C(n1056), .D(n1136), .Z(n841) );
  CND2X1 U1123 ( .A(n842), .B(n841), .Z(n969) );
  CANR2X1 U1124 ( .A(n888), .B(n843), .C(n877), .D(n969), .Z(n844) );
  CND2X1 U1125 ( .A(n845), .B(n844), .Z(n1016) );
  CANR2X1 U1126 ( .A(n460), .B(n458), .C(n477), .D(n456), .Z(n846) );
  CANR2X1 U1127 ( .A(N162), .B(net16921), .C(N34), .D(net16919), .Z(n848) );
  CANR2X1 U1128 ( .A(N291), .B(net16920), .C(acc[18]), .D(net6623), .Z(n847)
         );
  CND2X1 U1129 ( .A(n848), .B(n847), .Z(n191) );
  CANR2X1 U1130 ( .A(n893), .B(n887), .C(n892), .D(n936), .Z(n853) );
  CANR2X1 U1131 ( .A(n1055), .B(n1136), .C(n1054), .D(n1138), .Z(n850) );
  CIVX2 U1132 ( .A(acc[18]), .Z(n1134) );
  CANR2X1 U1133 ( .A(n1075), .B(n1140), .C(n1056), .D(n1134), .Z(n849) );
  CND2X1 U1134 ( .A(n850), .B(n849), .Z(n980) );
  CANR2X1 U1135 ( .A(n888), .B(n851), .C(n877), .D(n980), .Z(n852) );
  CND2X1 U1136 ( .A(n853), .B(n852), .Z(n1026) );
  CANR2X1 U1137 ( .A(n469), .B(n458), .C(n482), .D(n456), .Z(n854) );
  CANR2X1 U1138 ( .A(N290), .B(net16920), .C(acc[17]), .D(net6623), .Z(n855)
         );
  CND2X1 U1139 ( .A(n856), .B(n855), .Z(n192) );
  CANR2X1 U1140 ( .A(n893), .B(n902), .C(n892), .D(n947), .Z(n861) );
  CANR2X1 U1141 ( .A(n1055), .B(n1134), .C(n1054), .D(n1136), .Z(n858) );
  CIVX2 U1142 ( .A(acc[17]), .Z(n1132) );
  CANR2X1 U1143 ( .A(n1075), .B(n1138), .C(n1056), .D(n1132), .Z(n857) );
  CND2X1 U1144 ( .A(n858), .B(n857), .Z(n991) );
  CANR2X1 U1145 ( .A(n888), .B(n859), .C(n877), .D(n991), .Z(n860) );
  CND2X1 U1146 ( .A(n861), .B(n860), .Z(n1040) );
  CANR2X1 U1147 ( .A(n464), .B(n458), .C(n479), .D(n456), .Z(n862) );
  CANR2X1 U1148 ( .A(N289), .B(net16920), .C(acc[16]), .D(net6623), .Z(n863)
         );
  CND2X1 U1149 ( .A(n864), .B(n863), .Z(n193) );
  CANR2X1 U1150 ( .A(n893), .B(n914), .C(n892), .D(n958), .Z(n869) );
  CANR2X1 U1151 ( .A(n1055), .B(n1132), .C(n1054), .D(n1134), .Z(n866) );
  CANR2X1 U1152 ( .A(n1075), .B(n1136), .C(n1056), .D(n1130), .Z(n865) );
  CND2X1 U1153 ( .A(n866), .B(n865), .Z(n1002) );
  CANR2X1 U1154 ( .A(n888), .B(n867), .C(n877), .D(n1002), .Z(n868) );
  CND2X1 U1155 ( .A(n869), .B(n868), .Z(n1053) );
  CANR2X1 U1156 ( .A(n465), .B(n458), .C(n480), .D(n456), .Z(n870) );
  CANR2X1 U1157 ( .A(N288), .B(net16920), .C(acc[15]), .D(net6623), .Z(n872)
         );
  CND2X1 U1158 ( .A(n873), .B(n872), .Z(n194) );
  CIVX2 U1159 ( .A(n874), .Z(n1088) );
  CANR2X1 U1160 ( .A(n893), .B(n925), .C(n892), .D(n969), .Z(n880) );
  CANR2X1 U1161 ( .A(n1055), .B(n1130), .C(n1054), .D(n1132), .Z(n876) );
  CANR2X1 U1162 ( .A(n1075), .B(n1134), .C(n1056), .D(n1128), .Z(n875) );
  CND2X1 U1163 ( .A(n876), .B(n875), .Z(n1013) );
  CANR2X1 U1164 ( .A(n888), .B(n878), .C(n877), .D(n1013), .Z(n879) );
  CANR2X1 U1165 ( .A(n456), .B(n1088), .C(n881), .D(n468), .Z(n882) );
  CANR2X1 U1166 ( .A(N287), .B(net16920), .C(acc[14]), .D(net6623), .Z(n884)
         );
  CND2X1 U1167 ( .A(n885), .B(n884), .Z(n195) );
  CIVX2 U1168 ( .A(n886), .Z(n898) );
  CIVX2 U1169 ( .A(n887), .Z(n896) );
  CND2X1 U1170 ( .A(n888), .B(n507), .Z(n1052) );
  CANR2X1 U1171 ( .A(n1055), .B(n1128), .C(n1054), .D(n1130), .Z(n890) );
  CANR2X1 U1172 ( .A(n1075), .B(n1132), .C(n1056), .D(n1126), .Z(n889) );
  CND2X1 U1173 ( .A(n890), .B(n889), .Z(n1025) );
  COND2X1 U1174 ( .A(n507), .B(n891), .C(n1060), .D(n1025), .Z(n895) );
  COND2X1 U1175 ( .A(n1084), .B(n980), .C(n1077), .D(n936), .Z(n894) );
  CANR3X1 U1176 ( .A(n896), .B(n1081), .C(n895), .D(n894), .Z(n897) );
  COND2X1 U1177 ( .A(n898), .B(n1069), .C(n897), .D(n1067), .Z(N223) );
  CANR2X1 U1178 ( .A(N286), .B(net16920), .C(acc[13]), .D(net6623), .Z(n899)
         );
  CND2X1 U1179 ( .A(n900), .B(n899), .Z(n196) );
  CIVX2 U1180 ( .A(n901), .Z(n910) );
  CIVX2 U1181 ( .A(n902), .Z(n908) );
  CANR2X1 U1182 ( .A(n1055), .B(n1126), .C(n1054), .D(n1128), .Z(n904) );
  CANR2X1 U1183 ( .A(n1075), .B(n1130), .C(n1056), .D(n1124), .Z(n903) );
  CND2X1 U1184 ( .A(n904), .B(n903), .Z(n1039) );
  COND2X1 U1185 ( .A(n504), .B(n905), .C(n1060), .D(n1039), .Z(n907) );
  COND2X1 U1186 ( .A(n1084), .B(n991), .C(n1077), .D(n947), .Z(n906) );
  CANR3X1 U1187 ( .A(n908), .B(n1081), .C(n907), .D(n906), .Z(n909) );
  COND2X1 U1188 ( .A(n910), .B(n1069), .C(n909), .D(n1067), .Z(N222) );
  CANR2X1 U1189 ( .A(N285), .B(net16920), .C(acc[12]), .D(net6623), .Z(n911)
         );
  CND2X1 U1190 ( .A(n912), .B(n911), .Z(n197) );
  CIVX2 U1191 ( .A(n913), .Z(n922) );
  CIVX2 U1192 ( .A(n914), .Z(n920) );
  CANR2X1 U1193 ( .A(n1055), .B(n1124), .C(n1054), .D(n1126), .Z(n916) );
  CANR2X1 U1194 ( .A(n1075), .B(n1128), .C(n1056), .D(n1122), .Z(n915) );
  CND2X1 U1195 ( .A(n916), .B(n915), .Z(n1051) );
  COND2X1 U1196 ( .A(n505), .B(n917), .C(n1060), .D(n1051), .Z(n919) );
  COND2X1 U1197 ( .A(n1084), .B(n1002), .C(n1077), .D(n958), .Z(n918) );
  CANR3X1 U1198 ( .A(n920), .B(n1081), .C(n919), .D(n918), .Z(n921) );
  COND2X1 U1199 ( .A(n922), .B(n1069), .C(n921), .D(n1067), .Z(N221) );
  CANR2X1 U1200 ( .A(N284), .B(net16920), .C(acc[11]), .D(net6623), .Z(n923)
         );
  CND2X1 U1201 ( .A(n924), .B(n923), .Z(n198) );
  CIVX2 U1202 ( .A(n925), .Z(n931) );
  CANR2X1 U1203 ( .A(n1055), .B(n1122), .C(n1054), .D(n1124), .Z(n927) );
  CANR2X1 U1204 ( .A(n1075), .B(n1126), .C(n1056), .D(n1120), .Z(n926) );
  CND2X1 U1205 ( .A(n927), .B(n926), .Z(n1079) );
  COND2X1 U1206 ( .A(n504), .B(n928), .C(n1060), .D(n1079), .Z(n930) );
  COND2X1 U1207 ( .A(n1084), .B(n1013), .C(n1077), .D(n969), .Z(n929) );
  CANR3X1 U1208 ( .A(n931), .B(n1081), .C(n930), .D(n929), .Z(n932) );
  COND2X1 U1209 ( .A(n933), .B(n1069), .C(n932), .D(n1067), .Z(N220) );
  CANR2X1 U1210 ( .A(N283), .B(net16920), .C(acc[10]), .D(net6623), .Z(n934)
         );
  CND2X1 U1211 ( .A(n935), .B(n934), .Z(n199) );
  CIVX2 U1212 ( .A(n936), .Z(n942) );
  CANR2X1 U1213 ( .A(n1055), .B(n1120), .C(n1054), .D(n1122), .Z(n938) );
  CANR2X1 U1214 ( .A(n1075), .B(n1124), .C(n1056), .D(n1118), .Z(n937) );
  CND2X1 U1215 ( .A(n938), .B(n937), .Z(n1027) );
  COND2X1 U1216 ( .A(n504), .B(n939), .C(n1060), .D(n1027), .Z(n941) );
  COND2X1 U1217 ( .A(n1084), .B(n1025), .C(n1077), .D(n980), .Z(n940) );
  CANR3X1 U1218 ( .A(n942), .B(n1081), .C(n941), .D(n940), .Z(n943) );
  COND2X1 U1219 ( .A(n944), .B(n1069), .C(n943), .D(n1067), .Z(N219) );
  CANR2X1 U1220 ( .A(N282), .B(net16920), .C(acc[9]), .D(net6623), .Z(n945) );
  CND2X1 U1221 ( .A(n946), .B(n945), .Z(n200) );
  CIVX2 U1222 ( .A(n947), .Z(n953) );
  CANR2X1 U1223 ( .A(n1055), .B(n1118), .C(n1054), .D(n1120), .Z(n949) );
  CANR2X1 U1224 ( .A(n1075), .B(n1122), .C(n1056), .D(n1116), .Z(n948) );
  CND2X1 U1225 ( .A(n949), .B(n948), .Z(n1041) );
  COND2X1 U1226 ( .A(n506), .B(n950), .C(n1060), .D(n1041), .Z(n952) );
  COND2X1 U1227 ( .A(n1084), .B(n1039), .C(n1077), .D(n991), .Z(n951) );
  CANR3X1 U1228 ( .A(n953), .B(n1081), .C(n952), .D(n951), .Z(n954) );
  COND2X1 U1229 ( .A(n955), .B(n1069), .C(n954), .D(n1067), .Z(N218) );
  CANR2X1 U1230 ( .A(N281), .B(net16920), .C(acc[8]), .D(net6623), .Z(n956) );
  CND2X1 U1231 ( .A(n957), .B(n956), .Z(n201) );
  CIVX2 U1232 ( .A(n958), .Z(n964) );
  CANR2X1 U1233 ( .A(n1055), .B(n1116), .C(n1054), .D(n1118), .Z(n960) );
  CANR2X1 U1234 ( .A(n1075), .B(n1120), .C(n1056), .D(n1114), .Z(n959) );
  CND2X1 U1235 ( .A(n960), .B(n959), .Z(n1057) );
  COND2X1 U1236 ( .A(n504), .B(n961), .C(n1060), .D(n1057), .Z(n963) );
  COND2X1 U1237 ( .A(n1084), .B(n1051), .C(n1077), .D(n1002), .Z(n962) );
  CANR3X1 U1238 ( .A(n964), .B(n1081), .C(n963), .D(n962), .Z(n965) );
  COND2X1 U1239 ( .A(n966), .B(n1069), .C(n965), .D(n1067), .Z(N217) );
  CANR2X1 U1240 ( .A(N280), .B(net16920), .C(acc[7]), .D(net6623), .Z(n967) );
  CND2X1 U1241 ( .A(n968), .B(n967), .Z(n202) );
  CIVX2 U1242 ( .A(n969), .Z(n975) );
  CANR2X1 U1243 ( .A(n1055), .B(n1114), .C(n1054), .D(n1116), .Z(n971) );
  CANR2X1 U1244 ( .A(n1075), .B(n1118), .C(n1056), .D(n1112), .Z(n970) );
  CND2X1 U1245 ( .A(n971), .B(n970), .Z(n1078) );
  COND2X1 U1246 ( .A(n504), .B(n972), .C(n1060), .D(n1078), .Z(n974) );
  COND2X1 U1247 ( .A(n1084), .B(n1079), .C(n1077), .D(n1013), .Z(n973) );
  CANR3X1 U1248 ( .A(n975), .B(n1081), .C(n974), .D(n973), .Z(n976) );
  COND2X1 U1249 ( .A(n977), .B(n1069), .C(n976), .D(n1067), .Z(N216) );
  CANR2X1 U1250 ( .A(N279), .B(net16920), .C(acc[6]), .D(net6623), .Z(n978) );
  CND2X1 U1251 ( .A(n979), .B(n978), .Z(n203) );
  CIVX2 U1252 ( .A(n980), .Z(n986) );
  CANR2X1 U1253 ( .A(n1055), .B(n1112), .C(n1054), .D(n1114), .Z(n982) );
  CANR2X1 U1254 ( .A(n1075), .B(n1116), .C(n1056), .D(n1110), .Z(n981) );
  CND2X1 U1255 ( .A(n982), .B(n981), .Z(n1024) );
  COND2X1 U1256 ( .A(n504), .B(n983), .C(n1060), .D(n1024), .Z(n985) );
  COND2X1 U1257 ( .A(n1084), .B(n1027), .C(n1077), .D(n1025), .Z(n984) );
  CANR3X1 U1258 ( .A(n986), .B(n1081), .C(n985), .D(n984), .Z(n987) );
  COND2X1 U1259 ( .A(n988), .B(n1069), .C(n987), .D(n1067), .Z(N215) );
  CANR2X1 U1260 ( .A(N278), .B(net16920), .C(acc[5]), .D(net6623), .Z(n989) );
  CND2X1 U1261 ( .A(n990), .B(n989), .Z(n204) );
  CIVX2 U1262 ( .A(n991), .Z(n997) );
  CANR2X1 U1263 ( .A(n1055), .B(n1110), .C(n1054), .D(n1112), .Z(n993) );
  CANR2X1 U1264 ( .A(n1075), .B(n1114), .C(n1056), .D(n1108), .Z(n992) );
  CND2X1 U1265 ( .A(n993), .B(n992), .Z(n1038) );
  COND2X1 U1266 ( .A(n505), .B(n994), .C(n1060), .D(n1038), .Z(n996) );
  COND2X1 U1267 ( .A(n1084), .B(n1041), .C(n1077), .D(n1039), .Z(n995) );
  CANR3X1 U1268 ( .A(n997), .B(n1081), .C(n996), .D(n995), .Z(n998) );
  COND2X1 U1269 ( .A(n999), .B(n1069), .C(n998), .D(n1067), .Z(N214) );
  CANR2X1 U1270 ( .A(N148), .B(net16921), .C(N20), .D(net16919), .Z(n1001) );
  CND2X1 U1271 ( .A(n1001), .B(n1000), .Z(n205) );
  CIVX2 U1272 ( .A(n1002), .Z(n1008) );
  CANR2X1 U1273 ( .A(n1055), .B(n1108), .C(n1054), .D(n1110), .Z(n1004) );
  CANR2X1 U1274 ( .A(n1075), .B(n1112), .C(n1056), .D(n1106), .Z(n1003) );
  CND2X1 U1275 ( .A(n1004), .B(n1003), .Z(n1050) );
  COND2X1 U1276 ( .A(n504), .B(n1005), .C(n1060), .D(n1050), .Z(n1007) );
  COND2X1 U1277 ( .A(n1084), .B(n1057), .C(n1077), .D(n1051), .Z(n1006) );
  CANR3X1 U1278 ( .A(n1008), .B(n1081), .C(n1007), .D(n1006), .Z(n1009) );
  COND2X1 U1279 ( .A(n1010), .B(n1069), .C(n1009), .D(n1067), .Z(N213) );
  CANR2X1 U1280 ( .A(N147), .B(net16921), .C(N19), .D(net16919), .Z(n1012) );
  CND2X1 U1281 ( .A(n1012), .B(n1011), .Z(n206) );
  CIVX2 U1282 ( .A(n1013), .Z(n1019) );
  CANR2X1 U1283 ( .A(n1055), .B(n1106), .C(n1054), .D(n1108), .Z(n1015) );
  CIVX2 U1284 ( .A(acc[3]), .Z(n1104) );
  CANR2X1 U1285 ( .A(n1075), .B(n1110), .C(n1056), .D(n1104), .Z(n1014) );
  CND2X1 U1286 ( .A(n1015), .B(n1014), .Z(n1085) );
  COND2X1 U1287 ( .A(n506), .B(n1016), .C(n1060), .D(n1085), .Z(n1018) );
  COND2X1 U1288 ( .A(n1078), .B(n1084), .C(n1077), .D(n1079), .Z(n1017) );
  CANR3X1 U1289 ( .A(n1019), .B(n1081), .C(n1018), .D(n1017), .Z(n1020) );
  COND2X1 U1290 ( .A(n1021), .B(n1069), .C(n1020), .D(n1067), .Z(N212) );
  CANR2X1 U1291 ( .A(N146), .B(net16921), .C(N18), .D(net16919), .Z(n1023) );
  CND2X1 U1292 ( .A(n1023), .B(n1022), .Z(n207) );
  CIVX2 U1293 ( .A(n1024), .Z(n1033) );
  CIVX2 U1294 ( .A(n1084), .Z(n1065) );
  COND2X1 U1295 ( .A(n505), .B(n1026), .C(n1052), .D(n1025), .Z(n1032) );
  CANR2X1 U1296 ( .A(acc[3]), .B(n1055), .C(acc[4]), .D(n1054), .Z(n1030) );
  CANR2X1 U1297 ( .A(acc[5]), .B(n1075), .C(acc[2]), .D(n1056), .Z(n1029) );
  CIVX2 U1298 ( .A(n1077), .Z(n1058) );
  COND4CX1 U1299 ( .A(n1030), .B(n1029), .C(n1060), .D(n1028), .Z(n1031) );
  CANR3X1 U1300 ( .A(n1033), .B(n1065), .C(n1032), .D(n1031), .Z(n1034) );
  COND2X1 U1301 ( .A(n1035), .B(n1069), .C(n1034), .D(n1067), .Z(N211) );
  CANR2X1 U1302 ( .A(N145), .B(net16921), .C(N17), .D(net16919), .Z(n1037) );
  CND2X1 U1303 ( .A(n1037), .B(n1036), .Z(n208) );
  CIVX2 U1304 ( .A(n1038), .Z(n1047) );
  COND2X1 U1305 ( .A(n505), .B(n1040), .C(n1052), .D(n1039), .Z(n1046) );
  CANR2X1 U1306 ( .A(acc[2]), .B(n1055), .C(acc[3]), .D(n1054), .Z(n1044) );
  CANR2X1 U1307 ( .A(acc[4]), .B(n1075), .C(acc[1]), .D(n1056), .Z(n1043) );
  COND4CX1 U1308 ( .A(n1044), .B(n1043), .C(n1060), .D(n1042), .Z(n1045) );
  CANR3X1 U1309 ( .A(n1047), .B(n1065), .C(n1046), .D(n1045), .Z(n1048) );
  COND2X1 U1310 ( .A(n1049), .B(n1069), .C(n1048), .D(n1067), .Z(N210) );
  CIVX2 U1311 ( .A(n1050), .Z(n1066) );
  COND2X1 U1312 ( .A(n505), .B(n1053), .C(n1052), .D(n1051), .Z(n1064) );
  CANR2X1 U1313 ( .A(acc[1]), .B(n1055), .C(acc[2]), .D(n1054), .Z(n1062) );
  CANR2X1 U1314 ( .A(acc[3]), .B(n1075), .C(n1056), .D(acc[0]), .Z(n1061) );
  COND4CX1 U1315 ( .A(n1062), .B(n1061), .C(n1060), .D(n1059), .Z(n1063) );
  CANR3X1 U1316 ( .A(n1066), .B(n1065), .C(n1064), .D(n1063), .Z(n1068) );
  COND2X1 U1317 ( .A(n1070), .B(n1069), .C(n1068), .D(n1067), .Z(N209) );
  CIVX2 U1318 ( .A(acc[1]), .Z(n1102) );
  CIVX2 U1319 ( .A(acc[0]), .Z(n1100) );
  COND2X1 U1320 ( .A(n1072), .B(n1102), .C(n1100), .D(n1071), .Z(n1074) );
  COND4CX1 U1321 ( .A(acc[2]), .B(n1075), .C(n1074), .D(n1073), .Z(n1076) );
  COAN1X1 U1322 ( .A(n1078), .B(n1077), .C(n1076), .Z(n1083) );
  CIVX2 U1323 ( .A(n1079), .Z(n1080) );
  COND3X1 U1324 ( .A(n1085), .B(n1084), .C(n1083), .D(n1082), .Z(n1086) );
  CANR2X1 U1325 ( .A(n458), .B(n1088), .C(n1087), .D(n1086), .Z(n1094) );
  CAN2X1 U1326 ( .A(n470), .B(n1090), .Z(n1091) );
  CND2X1 U1327 ( .A(n1094), .B(n1093), .Z(N208) );
  CANR2X1 U1328 ( .A(N144), .B(net16921), .C(N16), .D(net16919), .Z(n1099) );
  CANR2X1 U1329 ( .A(N273), .B(net16920), .C(acc[0]), .D(net6623), .Z(n1098)
         );
  CND2X1 U1330 ( .A(n1099), .B(n1098), .Z(n209) );
  CIVX2 U1331 ( .A(net13424), .Z(net13361) );
endmodule

