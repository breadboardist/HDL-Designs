
module sfilt_DW01_add_2 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n83, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n133, n134, n135, n136, n137, n138, n139,
         n140, n142, n145, n146, n147, n148, n149, n150, n151, n153, n154,
         n155, n156, n157, n158, n159, n160, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n179, n180,
         n181, n182, n183, n184, n185, n186, n188, n191, n192, n193, n194,
         n195, n196, n197, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n235,
         n236, n237, n238, n239, n240, n243, n244, n245, n246, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n267, n268, n269, n270, n271, n272, n273, n274,
         n276, n279, n280, n281, n282, n283, n284, n285, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n323, n324, n325, n326, n327, n328, n331,
         n332, n333, n334, n335, n336, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n351, n352, n353, n354, n355, n356, n357,
         n360, n361, n362, n363, n364, n365, n366, n369, n370, n373, n374,
         n375, n376, n379, n380, n381, n382, n383, n384, n385, n386, n389,
         n390, n391, n392, n394, n397, n398, n399, n401, n402, n403, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n425, n426, n427, n428, n429,
         n430, n431, n432, n434, n437, n438, n439, n440, n441, n442, n443,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n481, n482, n483, n484,
         n485, n486, n489, n490, n491, n492, n493, n494, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n509, n510, n511, n512,
         n513, n514, n515, n518, n519, n520, n521, n522, n523, n524, n527,
         n528, n531, n532, n533, n534, n537, n538, n539, n540, n541, n542,
         n543, n544, n547, n548, n549, n550, n552, n555, n556, n557, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n574, n575, n576, n577, n578, n579, n580, n583, n584,
         n585, n586, n588, n589, n590, n591, n592, n593, n594, n595, n598,
         n599, n600, n601, n602, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n915, n916, n917;

  COND1X1 U123 ( .A(n163), .B(n206), .C(n164), .Z(n5) );
  COND1X1 U347 ( .A(n339), .B(n374), .C(n340), .Z(n334) );
  COND1X1 U553 ( .A(n497), .B(n532), .C(n498), .Z(n492) );
  CNR2XL U784 ( .A(n486), .B(n481), .Z(n475) );
  CNR2XL U785 ( .A(n544), .B(n539), .Z(n537) );
  CNR2XL U786 ( .A(n222), .B(n213), .Z(n211) );
  CNR2XL U787 ( .A(B[24]), .B(A[24]), .Z(n486) );
  CND2XL U788 ( .A(B[2]), .B(A[2]), .Z(n646) );
  CND2X1 U789 ( .A(B[36]), .B(A[36]), .Z(n369) );
  CNR2XL U790 ( .A(n560), .B(n555), .Z(n549) );
  CNR2XL U791 ( .A(B[28]), .B(A[28]), .Z(n446) );
  CNR2XL U792 ( .A(B[16]), .B(A[16]), .Z(n560) );
  CND2XL U793 ( .A(n580), .B(n568), .Z(n566) );
  CNR2X1 U794 ( .A(n589), .B(n584), .Z(n580) );
  CANR1XL U795 ( .A(n140), .B(n119), .C(n120), .Z(n118) );
  CANR1XL U796 ( .A(n648), .B(n640), .C(n641), .Z(n639) );
  COND1XL U797 ( .A(n561), .B(n555), .C(n556), .Z(n550) );
  COND1XL U798 ( .A(n447), .B(n437), .C(n438), .Z(n432) );
  CNR2X1 U799 ( .A(B[40]), .B(A[40]), .Z(n328) );
  CNR2X1 U800 ( .A(B[44]), .B(A[44]), .Z(n288) );
  CNR2XL U801 ( .A(n4), .B(n159), .Z(n157) );
  CNR2XL U802 ( .A(n4), .B(n89), .Z(n87) );
  CNR2XL U803 ( .A(n4), .B(n113), .Z(n111) );
  CND2XL U804 ( .A(n6), .B(n91), .Z(n89) );
  CND2XL U805 ( .A(n6), .B(n115), .Z(n113) );
  CNR2XL U806 ( .A(n335), .B(n260), .Z(n258) );
  CNR2XL U807 ( .A(n493), .B(n418), .Z(n416) );
  CANR1X1 U808 ( .A(n618), .B(n564), .C(n565), .Z(n563) );
  CNIVX2 U809 ( .A(n2), .Z(n917) );
  CND2XL U810 ( .A(n375), .B(n357), .Z(n355) );
  CND2XL U811 ( .A(n533), .B(n515), .Z(n513) );
  CND2XL U812 ( .A(n6), .B(n128), .Z(n126) );
  CND2XL U813 ( .A(n6), .B(n139), .Z(n137) );
  CND2XL U814 ( .A(n6), .B(n660), .Z(n150) );
  CND2XL U815 ( .A(n229), .B(n666), .Z(n218) );
  CND2XL U816 ( .A(n174), .B(n207), .Z(n172) );
  CND2XL U817 ( .A(n207), .B(n185), .Z(n183) );
  CND2XL U818 ( .A(n453), .B(n431), .Z(n429) );
  CANR1X1 U819 ( .A(n230), .B(n211), .C(n212), .Z(n206) );
  CANR1X1 U820 ( .A(n392), .B(n379), .C(n380), .Z(n374) );
  CANR1X1 U821 ( .A(n550), .B(n537), .C(n538), .Z(n532) );
  CANR1X1 U822 ( .A(n611), .B(n598), .C(n599), .Z(n593) );
  CANR1X1 U823 ( .A(n476), .B(n457), .C(n458), .Z(n452) );
  CANR1X1 U824 ( .A(n318), .B(n299), .C(n300), .Z(n294) );
  CNR2XL U825 ( .A(n645), .B(n642), .Z(n640) );
  COND1X1 U826 ( .A(n619), .B(n639), .C(n620), .Z(n618) );
  CND2XL U827 ( .A(n629), .B(n621), .Z(n619) );
  CNR2XL U828 ( .A(n626), .B(n623), .Z(n621) );
  CNR2XL U829 ( .A(n513), .B(n506), .Z(n504) );
  CNR2XL U830 ( .A(n328), .B(n323), .Z(n317) );
  CNR2XL U831 ( .A(n154), .B(n145), .Z(n139) );
  CNR2XL U832 ( .A(n288), .B(n279), .Z(n273) );
  CNR2XL U833 ( .A(n615), .B(n612), .Z(n610) );
  CNR2XL U834 ( .A(n106), .B(n97), .Z(n95) );
  CNR2XL U835 ( .A(n402), .B(n397), .Z(n391) );
  CNR2XL U836 ( .A(n605), .B(n600), .Z(n598) );
  CNR2XL U837 ( .A(n468), .B(n459), .Z(n457) );
  CNR2XL U838 ( .A(n575), .B(n570), .Z(n568) );
  CNR2XL U839 ( .A(n386), .B(n381), .Z(n379) );
  CNR2XL U840 ( .A(n310), .B(n301), .Z(n299) );
  CNR2XL U841 ( .A(n422), .B(n413), .Z(n411) );
  CNR2XL U842 ( .A(n348), .B(n343), .Z(n341) );
  CNR2XL U843 ( .A(n264), .B(n255), .Z(n253) );
  CNR2XL U844 ( .A(n130), .B(n121), .Z(n119) );
  CNR2IXL U845 ( .B(n139), .A(n130), .Z(n128) );
  CNR2XL U846 ( .A(n355), .B(n348), .Z(n346) );
  CNR2XL U847 ( .A(B[8]), .B(A[8]), .Z(n615) );
  CNR2XL U848 ( .A(B[32]), .B(A[32]), .Z(n402) );
  CNR2XL U849 ( .A(B[56]), .B(A[56]), .Z(n154) );
  CND2XL U850 ( .A(B[18]), .B(A[18]), .Z(n547) );
  CND2XL U851 ( .A(B[22]), .B(A[22]), .Z(n509) );
  CND2XL U852 ( .A(B[6]), .B(A[6]), .Z(n627) );
  CND2XL U853 ( .A(B[30]), .B(A[30]), .Z(n425) );
  CND2XL U854 ( .A(B[34]), .B(A[34]), .Z(n389) );
  CND2XL U855 ( .A(B[58]), .B(A[58]), .Z(n133) );
  CND2XL U856 ( .A(B[46]), .B(A[46]), .Z(n267) );
  CND2XL U857 ( .A(B[38]), .B(A[38]), .Z(n351) );
  CND2XL U858 ( .A(B[1]), .B(A[1]), .Z(n650) );
  CEOXL U859 ( .A(n22), .B(n244), .Z(SUM[48]) );
  CEOXL U860 ( .A(n23), .B(n257), .Z(SUM[47]) );
  CEOXL U861 ( .A(n24), .B(n268), .Z(SUM[46]) );
  CEOXL U862 ( .A(n25), .B(n281), .Z(SUM[45]) );
  CEOXL U863 ( .A(n26), .B(n290), .Z(SUM[44]) );
  CEOXL U864 ( .A(n27), .B(n303), .Z(SUM[43]) );
  CEOXL U865 ( .A(n28), .B(n312), .Z(SUM[42]) );
  CEOXL U866 ( .A(n29), .B(n325), .Z(SUM[41]) );
  CEOXL U867 ( .A(n30), .B(n332), .Z(SUM[40]) );
  CEOXL U868 ( .A(n31), .B(n345), .Z(SUM[39]) );
  CEOXL U869 ( .A(n32), .B(n352), .Z(SUM[38]) );
  CEOXL U870 ( .A(n33), .B(n363), .Z(SUM[37]) );
  CEOXL U871 ( .A(n34), .B(n370), .Z(SUM[36]) );
  CEOXL U872 ( .A(n35), .B(n383), .Z(SUM[35]) );
  CEOXL U873 ( .A(n36), .B(n390), .Z(SUM[34]) );
  CEOXL U874 ( .A(n37), .B(n399), .Z(SUM[33]) );
  CEOXL U875 ( .A(n7), .B(n73), .Z(SUM[63]) );
  CEOXL U876 ( .A(n8), .B(n86), .Z(SUM[62]) );
  CEOXL U877 ( .A(n9), .B(n99), .Z(SUM[61]) );
  CEOXL U878 ( .A(n10), .B(n110), .Z(SUM[60]) );
  CEOXL U879 ( .A(n11), .B(n123), .Z(SUM[59]) );
  CEOXL U880 ( .A(n12), .B(n134), .Z(SUM[58]) );
  CEOXL U881 ( .A(n13), .B(n147), .Z(SUM[57]) );
  CEOXL U882 ( .A(n14), .B(n156), .Z(SUM[56]) );
  CEOXL U883 ( .A(n15), .B(n169), .Z(SUM[55]) );
  CEOXL U884 ( .A(n16), .B(n180), .Z(SUM[54]) );
  CEOXL U885 ( .A(n17), .B(n193), .Z(SUM[53]) );
  CEOXL U886 ( .A(n18), .B(n202), .Z(SUM[52]) );
  CEOXL U887 ( .A(n19), .B(n215), .Z(SUM[51]) );
  CEOXL U888 ( .A(n20), .B(n224), .Z(SUM[50]) );
  CEOXL U889 ( .A(n21), .B(n237), .Z(SUM[49]) );
  CEOXL U890 ( .A(n39), .B(n415), .Z(SUM[31]) );
  CEOXL U891 ( .A(n40), .B(n426), .Z(SUM[30]) );
  CEOXL U892 ( .A(n41), .B(n439), .Z(SUM[29]) );
  CEOXL U893 ( .A(n42), .B(n448), .Z(SUM[28]) );
  CEOXL U894 ( .A(n43), .B(n461), .Z(SUM[27]) );
  CEOXL U895 ( .A(n44), .B(n470), .Z(SUM[26]) );
  CEOXL U896 ( .A(n45), .B(n483), .Z(SUM[25]) );
  CEOXL U897 ( .A(n46), .B(n490), .Z(SUM[24]) );
  CEOXL U898 ( .A(n47), .B(n503), .Z(SUM[23]) );
  CEOXL U899 ( .A(n48), .B(n510), .Z(SUM[22]) );
  CEOXL U900 ( .A(n49), .B(n521), .Z(SUM[21]) );
  CEOXL U901 ( .A(n50), .B(n528), .Z(SUM[20]) );
  CEOXL U902 ( .A(n51), .B(n541), .Z(SUM[19]) );
  CEOXL U903 ( .A(n52), .B(n548), .Z(SUM[18]) );
  CEOXL U904 ( .A(n53), .B(n557), .Z(SUM[17]) );
  CEOXL U905 ( .A(n55), .B(n572), .Z(SUM[15]) );
  CEOXL U906 ( .A(n57), .B(n586), .Z(SUM[13]) );
  CEOXL U907 ( .A(n59), .B(n602), .Z(SUM[11]) );
  CEOXL U908 ( .A(n64), .B(n628), .Z(SUM[6]) );
  CND2IXL U909 ( .B(n651), .A(n652), .Z(n70) );
  CND2X1 U910 ( .A(n333), .B(n249), .Z(n4) );
  CNR2XL U911 ( .A(n4), .B(n76), .Z(n74) );
  CNR2X1 U912 ( .A(n205), .B(n163), .Z(n6) );
  CNR2X1 U913 ( .A(n373), .B(n339), .Z(n333) );
  CNR2X1 U914 ( .A(n293), .B(n251), .Z(n249) );
  CIVX2 U915 ( .A(n563), .Z(n562) );
  CNR2X1 U916 ( .A(n531), .B(n497), .Z(n491) );
  CNR2X1 U917 ( .A(n117), .B(n93), .Z(n91) );
  CNR2X1 U918 ( .A(n451), .B(n409), .Z(n407) );
  CNR2XL U919 ( .A(n4), .B(n102), .Z(n100) );
  CNR2XL U920 ( .A(n4), .B(n126), .Z(n124) );
  CNR2XL U921 ( .A(n4), .B(n137), .Z(n135) );
  CNR2XL U922 ( .A(n4), .B(n150), .Z(n148) );
  CNR2XL U923 ( .A(n4), .B(n172), .Z(n170) );
  CNR2XL U924 ( .A(n4), .B(n183), .Z(n181) );
  CNR2XL U925 ( .A(n4), .B(n196), .Z(n194) );
  CNR2XL U926 ( .A(n4), .B(n205), .Z(n203) );
  CNR2XL U927 ( .A(n4), .B(n218), .Z(n216) );
  CNR2XL U928 ( .A(n4), .B(n227), .Z(n225) );
  CNR2XL U929 ( .A(n335), .B(n271), .Z(n269) );
  CNR2XL U930 ( .A(n335), .B(n284), .Z(n282) );
  CNR2XL U931 ( .A(n335), .B(n293), .Z(n291) );
  CNR2XL U932 ( .A(n335), .B(n306), .Z(n304) );
  CNR2XL U933 ( .A(n335), .B(n315), .Z(n313) );
  CNR2XL U934 ( .A(n493), .B(n429), .Z(n427) );
  CNR2XL U935 ( .A(n493), .B(n442), .Z(n440) );
  CNR2XL U936 ( .A(n493), .B(n451), .Z(n449) );
  CNR2XL U937 ( .A(n493), .B(n464), .Z(n462) );
  CNR2XL U938 ( .A(n493), .B(n473), .Z(n471) );
  CND2XL U939 ( .A(n6), .B(n78), .Z(n76) );
  CANR1XL U940 ( .A(n629), .B(n638), .C(n630), .Z(n628) );
  COND1XL U941 ( .A(n578), .B(n617), .C(n579), .Z(n577) );
  CND2X1 U942 ( .A(n594), .B(n580), .Z(n578) );
  CANR1XL U943 ( .A(n580), .B(n595), .C(n583), .Z(n579) );
  COND1XL U944 ( .A(n592), .B(n617), .C(n593), .Z(n591) );
  COND1XL U945 ( .A(n608), .B(n617), .C(n609), .Z(n607) );
  CANR1XL U946 ( .A(n491), .B(n562), .C(n492), .Z(n490) );
  CNR2X1 U947 ( .A(n592), .B(n566), .Z(n564) );
  COND1XL U948 ( .A(n566), .B(n593), .C(n567), .Z(n565) );
  CANR1XL U949 ( .A(n357), .B(n376), .C(n360), .Z(n356) );
  CANR1XL U950 ( .A(n515), .B(n534), .C(n518), .Z(n514) );
  COND1XL U951 ( .A(n405), .B(n563), .C(n406), .Z(n2) );
  CND2XL U952 ( .A(n491), .B(n407), .Z(n405) );
  CANR1XL U953 ( .A(n492), .B(n407), .C(n408), .Z(n406) );
  CNR2X1 U954 ( .A(n117), .B(n80), .Z(n78) );
  CND2X1 U955 ( .A(n139), .B(n119), .Z(n117) );
  COND1XL U956 ( .A(n89), .B(n3), .C(n90), .Z(n88) );
  CANR1XL U957 ( .A(n91), .B(n5), .C(n92), .Z(n90) );
  COND1XL U958 ( .A(n93), .B(n118), .C(n94), .Z(n92) );
  COND1XL U959 ( .A(n113), .B(n3), .C(n114), .Z(n112) );
  CANR1XL U960 ( .A(n115), .B(n5), .C(n116), .Z(n114) );
  COND1XL U961 ( .A(n137), .B(n3), .C(n138), .Z(n136) );
  CANR1XL U962 ( .A(n139), .B(n5), .C(n140), .Z(n138) );
  COND1XL U963 ( .A(n159), .B(n3), .C(n160), .Z(n158) );
  COND1XL U964 ( .A(n183), .B(n3), .C(n184), .Z(n182) );
  CANR1XL U965 ( .A(n185), .B(n208), .C(n186), .Z(n184) );
  COND1XL U966 ( .A(n205), .B(n3), .C(n206), .Z(n204) );
  COND1XL U967 ( .A(n227), .B(n3), .C(n228), .Z(n226) );
  COND1XL U968 ( .A(n271), .B(n336), .C(n272), .Z(n270) );
  CANR1XL U969 ( .A(n273), .B(n296), .C(n274), .Z(n272) );
  COND1XL U970 ( .A(n293), .B(n336), .C(n294), .Z(n292) );
  COND1XL U971 ( .A(n315), .B(n336), .C(n316), .Z(n314) );
  COND1XL U972 ( .A(n429), .B(n494), .C(n430), .Z(n428) );
  CANR1XL U973 ( .A(n431), .B(n454), .C(n432), .Z(n430) );
  COND1XL U974 ( .A(n451), .B(n494), .C(n452), .Z(n450) );
  COND1XL U975 ( .A(n473), .B(n494), .C(n474), .Z(n472) );
  CND2X1 U976 ( .A(n229), .B(n211), .Z(n205) );
  CND2X1 U977 ( .A(n475), .B(n457), .Z(n451) );
  CND2X1 U978 ( .A(n317), .B(n299), .Z(n293) );
  CND2X1 U979 ( .A(n549), .B(n537), .Z(n531) );
  CND2X1 U980 ( .A(n391), .B(n379), .Z(n373) );
  CND2X1 U981 ( .A(n610), .B(n598), .Z(n592) );
  CND2X1 U982 ( .A(n515), .B(n499), .Z(n497) );
  CND2X1 U983 ( .A(n185), .B(n165), .Z(n163) );
  CND2X1 U984 ( .A(n273), .B(n253), .Z(n251) );
  CND2X1 U985 ( .A(n357), .B(n341), .Z(n339) );
  CND2X1 U986 ( .A(n431), .B(n411), .Z(n409) );
  CND2X1 U987 ( .A(n317), .B(n674), .Z(n306) );
  CND2X1 U988 ( .A(n475), .B(n690), .Z(n464) );
  CND2XL U989 ( .A(n6), .B(n104), .Z(n102) );
  CND2X1 U990 ( .A(n207), .B(n664), .Z(n196) );
  CND2X1 U991 ( .A(n295), .B(n273), .Z(n271) );
  CND2X1 U992 ( .A(n295), .B(n672), .Z(n284) );
  CND2X1 U993 ( .A(n453), .B(n688), .Z(n442) );
  CND2X1 U994 ( .A(n262), .B(n295), .Z(n260) );
  CND2X1 U995 ( .A(n420), .B(n453), .Z(n418) );
  COND1XL U996 ( .A(n251), .B(n294), .C(n252), .Z(n250) );
  CANR1XL U997 ( .A(n274), .B(n253), .C(n254), .Z(n252) );
  COND1XL U998 ( .A(n267), .B(n255), .C(n256), .Z(n254) );
  CANR1XL U999 ( .A(n186), .B(n165), .C(n166), .Z(n164) );
  COND1XL U1000 ( .A(n179), .B(n167), .C(n168), .Z(n166) );
  COND1XL U1001 ( .A(n133), .B(n121), .C(n122), .Z(n120) );
  CANR1XL U1002 ( .A(n360), .B(n341), .C(n342), .Z(n340) );
  COND1XL U1003 ( .A(n351), .B(n343), .C(n344), .Z(n342) );
  CANR1XL U1004 ( .A(n484), .B(n562), .C(n485), .Z(n483) );
  CNR2XL U1005 ( .A(n493), .B(n486), .Z(n484) );
  COND1XL U1006 ( .A(n486), .B(n494), .C(n489), .Z(n485) );
  CANR1XL U1007 ( .A(n504), .B(n562), .C(n505), .Z(n503) );
  COND1XL U1008 ( .A(n506), .B(n514), .C(n509), .Z(n505) );
  COND1XL U1009 ( .A(n606), .B(n600), .C(n601), .Z(n599) );
  COND1XL U1010 ( .A(n311), .B(n301), .C(n302), .Z(n300) );
  COND1XL U1011 ( .A(n469), .B(n459), .C(n460), .Z(n458) );
  COND1XL U1012 ( .A(n223), .B(n213), .C(n214), .Z(n212) );
  COND1XL U1013 ( .A(n547), .B(n539), .C(n540), .Z(n538) );
  COND1XL U1014 ( .A(n389), .B(n381), .C(n382), .Z(n380) );
  CANR1XL U1015 ( .A(n518), .B(n499), .C(n500), .Z(n498) );
  COND1XL U1016 ( .A(n509), .B(n501), .C(n502), .Z(n500) );
  COND1XL U1017 ( .A(n289), .B(n279), .C(n280), .Z(n274) );
  COND1XL U1018 ( .A(n403), .B(n397), .C(n398), .Z(n392) );
  COND1XL U1019 ( .A(n201), .B(n191), .C(n192), .Z(n186) );
  COND1XL U1020 ( .A(n155), .B(n145), .C(n146), .Z(n140) );
  COND1XL U1021 ( .A(n331), .B(n323), .C(n324), .Z(n318) );
  COND1XL U1022 ( .A(n489), .B(n481), .C(n482), .Z(n476) );
  COND1XL U1023 ( .A(n243), .B(n235), .C(n236), .Z(n230) );
  COND1XL U1024 ( .A(n646), .B(n642), .C(n643), .Z(n641) );
  CNR2X1 U1025 ( .A(n200), .B(n191), .Z(n185) );
  CNR2X1 U1026 ( .A(n446), .B(n437), .Z(n431) );
  CANR1XL U1027 ( .A(n630), .B(n621), .C(n622), .Z(n620) );
  COND1XL U1028 ( .A(n616), .B(n612), .C(n613), .Z(n611) );
  COND1XL U1029 ( .A(n652), .B(n649), .C(n650), .Z(n648) );
  COND1XL U1030 ( .A(n109), .B(n97), .C(n98), .Z(n96) );
  CNR2X1 U1031 ( .A(n240), .B(n235), .Z(n229) );
  CNR2X1 U1032 ( .A(n524), .B(n519), .Z(n515) );
  CNR2X1 U1033 ( .A(n366), .B(n361), .Z(n357) );
  COND1XL U1034 ( .A(n527), .B(n519), .C(n520), .Z(n518) );
  COND1XL U1035 ( .A(n637), .B(n631), .C(n632), .Z(n630) );
  COND1XL U1036 ( .A(n369), .B(n361), .C(n362), .Z(n360) );
  COND1XL U1037 ( .A(n590), .B(n584), .C(n585), .Z(n583) );
  CANR1XL U1038 ( .A(n583), .B(n568), .C(n569), .Z(n567) );
  COND1XL U1039 ( .A(n576), .B(n570), .C(n571), .Z(n569) );
  CNR2X1 U1040 ( .A(n117), .B(n106), .Z(n104) );
  CNR2X1 U1041 ( .A(n506), .B(n501), .Z(n499) );
  CNR2X1 U1042 ( .A(n176), .B(n167), .Z(n165) );
  COND1XL U1043 ( .A(n409), .B(n452), .C(n410), .Z(n408) );
  CANR1XL U1044 ( .A(n432), .B(n411), .C(n412), .Z(n410) );
  COND1XL U1045 ( .A(n425), .B(n413), .C(n414), .Z(n412) );
  COND1XL U1046 ( .A(n627), .B(n623), .C(n624), .Z(n622) );
  COND1XL U1047 ( .A(n76), .B(n3), .C(n77), .Z(n75) );
  CANR1XL U1048 ( .A(n78), .B(n5), .C(n79), .Z(n77) );
  COND1XL U1049 ( .A(n80), .B(n118), .C(n81), .Z(n79) );
  CANR1XL U1050 ( .A(n915), .B(n96), .C(n83), .Z(n81) );
  COND1XL U1051 ( .A(n102), .B(n3), .C(n103), .Z(n101) );
  CANR1XL U1052 ( .A(n104), .B(n5), .C(n105), .Z(n103) );
  COND1XL U1053 ( .A(n106), .B(n118), .C(n109), .Z(n105) );
  COND1XL U1054 ( .A(n126), .B(n3), .C(n127), .Z(n125) );
  CANR1XL U1055 ( .A(n128), .B(n5), .C(n129), .Z(n127) );
  COND1XL U1056 ( .A(n130), .B(n142), .C(n133), .Z(n129) );
  COND1XL U1057 ( .A(n150), .B(n3), .C(n151), .Z(n149) );
  CANR1XL U1058 ( .A(n660), .B(n5), .C(n153), .Z(n151) );
  COND1XL U1059 ( .A(n172), .B(n3), .C(n173), .Z(n171) );
  CANR1XL U1060 ( .A(n208), .B(n174), .C(n175), .Z(n173) );
  COND1XL U1061 ( .A(n176), .B(n188), .C(n179), .Z(n175) );
  COND1XL U1062 ( .A(n196), .B(n3), .C(n197), .Z(n195) );
  CANR1XL U1063 ( .A(n664), .B(n208), .C(n199), .Z(n197) );
  COND1XL U1064 ( .A(n218), .B(n3), .C(n219), .Z(n217) );
  CANR1XL U1065 ( .A(n666), .B(n230), .C(n221), .Z(n219) );
  COND1XL U1066 ( .A(n240), .B(n3), .C(n243), .Z(n239) );
  COND1XL U1067 ( .A(n366), .B(n374), .C(n369), .Z(n365) );
  COND1XL U1068 ( .A(n386), .B(n394), .C(n389), .Z(n385) );
  COND1XL U1069 ( .A(n524), .B(n532), .C(n527), .Z(n523) );
  COND1XL U1070 ( .A(n544), .B(n552), .C(n547), .Z(n543) );
  COND1XL U1071 ( .A(n260), .B(n336), .C(n261), .Z(n259) );
  CANR1XL U1072 ( .A(n296), .B(n262), .C(n263), .Z(n261) );
  COND1XL U1073 ( .A(n264), .B(n276), .C(n267), .Z(n263) );
  COND1XL U1074 ( .A(n284), .B(n336), .C(n285), .Z(n283) );
  CANR1XL U1075 ( .A(n672), .B(n296), .C(n287), .Z(n285) );
  COND1XL U1076 ( .A(n306), .B(n336), .C(n307), .Z(n305) );
  CANR1XL U1077 ( .A(n674), .B(n318), .C(n309), .Z(n307) );
  COND1XL U1078 ( .A(n328), .B(n336), .C(n331), .Z(n327) );
  COND1XL U1079 ( .A(n418), .B(n494), .C(n419), .Z(n417) );
  CANR1XL U1080 ( .A(n454), .B(n420), .C(n421), .Z(n419) );
  COND1XL U1081 ( .A(n422), .B(n434), .C(n425), .Z(n421) );
  COND1XL U1082 ( .A(n442), .B(n494), .C(n443), .Z(n441) );
  CANR1XL U1083 ( .A(n688), .B(n454), .C(n445), .Z(n443) );
  COND1XL U1084 ( .A(n464), .B(n494), .C(n465), .Z(n463) );
  CANR1XL U1085 ( .A(n690), .B(n476), .C(n467), .Z(n465) );
  COND1XL U1086 ( .A(n348), .B(n356), .C(n351), .Z(n347) );
  CNR2X1 U1087 ( .A(n636), .B(n631), .Z(n629) );
  CNR2IXL U1088 ( .B(n185), .A(n176), .Z(n174) );
  CNR2IXL U1089 ( .B(n273), .A(n264), .Z(n262) );
  CNR2IXL U1090 ( .B(n431), .A(n422), .Z(n420) );
  CNR2XL U1091 ( .A(n4), .B(n240), .Z(n238) );
  CNR2XL U1092 ( .A(n335), .B(n328), .Z(n326) );
  CNR2XL U1093 ( .A(n373), .B(n366), .Z(n364) );
  CNR2IXL U1094 ( .B(n391), .A(n386), .Z(n384) );
  CNR2XL U1095 ( .A(n531), .B(n524), .Z(n522) );
  CNR2IXL U1096 ( .B(n549), .A(n544), .Z(n542) );
  CND2X1 U1097 ( .A(n95), .B(n915), .Z(n80) );
  CNR2X1 U1098 ( .A(B[48]), .B(A[48]), .Z(n240) );
  CNR2X1 U1099 ( .A(B[20]), .B(A[20]), .Z(n524) );
  CNR2X1 U1100 ( .A(B[34]), .B(A[34]), .Z(n386) );
  CNR2X1 U1101 ( .A(B[18]), .B(A[18]), .Z(n544) );
  CNR2X1 U1102 ( .A(B[46]), .B(A[46]), .Z(n264) );
  CNR2X1 U1103 ( .A(B[38]), .B(A[38]), .Z(n348) );
  CNR2X1 U1104 ( .A(B[22]), .B(A[22]), .Z(n506) );
  CNR2X1 U1105 ( .A(B[36]), .B(A[36]), .Z(n366) );
  CNR2X1 U1106 ( .A(B[30]), .B(A[30]), .Z(n422) );
  CNR2X1 U1107 ( .A(B[54]), .B(A[54]), .Z(n176) );
  CNR2X1 U1108 ( .A(B[58]), .B(A[58]), .Z(n130) );
  CNR2X1 U1109 ( .A(B[60]), .B(A[60]), .Z(n106) );
  CNR2X1 U1110 ( .A(B[47]), .B(A[47]), .Z(n255) );
  CNR2X1 U1111 ( .A(B[23]), .B(A[23]), .Z(n501) );
  CNR2X1 U1112 ( .A(B[41]), .B(A[41]), .Z(n323) );
  CNR2X1 U1113 ( .A(B[45]), .B(A[45]), .Z(n279) );
  CNR2X1 U1114 ( .A(B[25]), .B(A[25]), .Z(n481) );
  CNR2X1 U1115 ( .A(B[17]), .B(A[17]), .Z(n555) );
  CNR2X1 U1116 ( .A(B[49]), .B(A[49]), .Z(n235) );
  CNR2X1 U1117 ( .A(B[35]), .B(A[35]), .Z(n381) );
  CNR2X1 U1118 ( .A(B[11]), .B(A[11]), .Z(n600) );
  CNR2X1 U1119 ( .A(B[53]), .B(A[53]), .Z(n191) );
  CNR2X1 U1120 ( .A(B[19]), .B(A[19]), .Z(n539) );
  CNR2X1 U1121 ( .A(B[21]), .B(A[21]), .Z(n519) );
  CNR2X1 U1122 ( .A(B[29]), .B(A[29]), .Z(n437) );
  CNR2X1 U1123 ( .A(B[43]), .B(A[43]), .Z(n301) );
  CNR2X1 U1124 ( .A(B[39]), .B(A[39]), .Z(n343) );
  CNR2X1 U1125 ( .A(B[33]), .B(A[33]), .Z(n397) );
  CNR2X1 U1126 ( .A(B[15]), .B(A[15]), .Z(n570) );
  CNR2X1 U1127 ( .A(B[27]), .B(A[27]), .Z(n459) );
  CNR2X1 U1128 ( .A(B[13]), .B(A[13]), .Z(n584) );
  CNR2X1 U1129 ( .A(B[37]), .B(A[37]), .Z(n361) );
  CNR2X1 U1130 ( .A(B[9]), .B(A[9]), .Z(n612) );
  CNR2X1 U1131 ( .A(B[51]), .B(A[51]), .Z(n213) );
  CNR2X1 U1132 ( .A(B[31]), .B(A[31]), .Z(n413) );
  CNR2X1 U1133 ( .A(B[7]), .B(A[7]), .Z(n623) );
  CNR2X1 U1134 ( .A(B[55]), .B(A[55]), .Z(n167) );
  CNR2X1 U1135 ( .A(B[5]), .B(A[5]), .Z(n631) );
  CNR2X1 U1136 ( .A(B[57]), .B(A[57]), .Z(n145) );
  CNR2X1 U1137 ( .A(B[3]), .B(A[3]), .Z(n642) );
  CNR2X1 U1138 ( .A(B[59]), .B(A[59]), .Z(n121) );
  CNR2X1 U1139 ( .A(B[61]), .B(A[61]), .Z(n97) );
  CNR2X1 U1140 ( .A(B[6]), .B(A[6]), .Z(n626) );
  CNR2X1 U1141 ( .A(B[2]), .B(A[2]), .Z(n645) );
  CNR2X1 U1142 ( .A(B[52]), .B(A[52]), .Z(n200) );
  CNR2X1 U1143 ( .A(B[42]), .B(A[42]), .Z(n310) );
  CNR2X1 U1144 ( .A(B[26]), .B(A[26]), .Z(n468) );
  CNR2X1 U1145 ( .A(B[50]), .B(A[50]), .Z(n222) );
  CNR2X1 U1146 ( .A(B[10]), .B(A[10]), .Z(n605) );
  CNR2X1 U1147 ( .A(B[12]), .B(A[12]), .Z(n589) );
  CNR2X1 U1148 ( .A(B[14]), .B(A[14]), .Z(n575) );
  CNR2X1 U1149 ( .A(B[4]), .B(A[4]), .Z(n636) );
  CND2X1 U1150 ( .A(B[0]), .B(A[0]), .Z(n652) );
  CNR2X1 U1151 ( .A(B[1]), .B(A[1]), .Z(n649) );
  COR2X1 U1152 ( .A(B[62]), .B(A[62]), .Z(n915) );
  CNR2XL U1153 ( .A(B[0]), .B(A[0]), .Z(n651) );
  COR2X1 U1154 ( .A(B[63]), .B(A[63]), .Z(n916) );
  CND2X1 U1155 ( .A(B[16]), .B(A[16]), .Z(n561) );
  CND2X1 U1156 ( .A(B[10]), .B(A[10]), .Z(n606) );
  CND2X1 U1157 ( .A(B[32]), .B(A[32]), .Z(n403) );
  CND2X1 U1158 ( .A(B[44]), .B(A[44]), .Z(n289) );
  CND2X1 U1159 ( .A(B[42]), .B(A[42]), .Z(n311) );
  CND2X1 U1160 ( .A(B[4]), .B(A[4]), .Z(n637) );
  CND2X1 U1161 ( .A(B[26]), .B(A[26]), .Z(n469) );
  CND2X1 U1162 ( .A(B[14]), .B(A[14]), .Z(n576) );
  CND2X1 U1163 ( .A(B[28]), .B(A[28]), .Z(n447) );
  CND2X1 U1164 ( .A(B[12]), .B(A[12]), .Z(n590) );
  CND2X1 U1165 ( .A(B[50]), .B(A[50]), .Z(n223) );
  CND2X1 U1166 ( .A(B[52]), .B(A[52]), .Z(n201) );
  CND2X1 U1167 ( .A(B[56]), .B(A[56]), .Z(n155) );
  CND2X1 U1168 ( .A(B[40]), .B(A[40]), .Z(n331) );
  CND2X1 U1169 ( .A(B[8]), .B(A[8]), .Z(n616) );
  CND2X1 U1170 ( .A(B[24]), .B(A[24]), .Z(n489) );
  CND2X1 U1171 ( .A(B[48]), .B(A[48]), .Z(n243) );
  CND2XL U1172 ( .A(B[20]), .B(A[20]), .Z(n527) );
  CND2XL U1173 ( .A(B[54]), .B(A[54]), .Z(n179) );
  CND2X1 U1174 ( .A(B[60]), .B(A[60]), .Z(n109) );
  CND2X1 U1175 ( .A(B[62]), .B(A[62]), .Z(n85) );
  CND2XL U1176 ( .A(B[47]), .B(A[47]), .Z(n256) );
  CND2XL U1177 ( .A(B[23]), .B(A[23]), .Z(n502) );
  CND2XL U1178 ( .A(B[11]), .B(A[11]), .Z(n601) );
  CND2XL U1179 ( .A(B[33]), .B(A[33]), .Z(n398) );
  CND2XL U1180 ( .A(B[45]), .B(A[45]), .Z(n280) );
  CND2XL U1181 ( .A(B[41]), .B(A[41]), .Z(n324) );
  CND2XL U1182 ( .A(B[9]), .B(A[9]), .Z(n613) );
  CND2XL U1183 ( .A(B[17]), .B(A[17]), .Z(n556) );
  CND2XL U1184 ( .A(B[35]), .B(A[35]), .Z(n382) );
  CND2XL U1185 ( .A(B[39]), .B(A[39]), .Z(n344) );
  CND2XL U1186 ( .A(B[43]), .B(A[43]), .Z(n302) );
  CND2XL U1187 ( .A(B[3]), .B(A[3]), .Z(n643) );
  CND2XL U1188 ( .A(B[25]), .B(A[25]), .Z(n482) );
  CND2XL U1189 ( .A(B[19]), .B(A[19]), .Z(n540) );
  CND2XL U1190 ( .A(B[27]), .B(A[27]), .Z(n460) );
  CND2XL U1191 ( .A(B[15]), .B(A[15]), .Z(n571) );
  CND2XL U1192 ( .A(B[7]), .B(A[7]), .Z(n624) );
  CND2XL U1193 ( .A(B[31]), .B(A[31]), .Z(n414) );
  CND2XL U1194 ( .A(B[13]), .B(A[13]), .Z(n585) );
  CND2XL U1195 ( .A(B[29]), .B(A[29]), .Z(n438) );
  CND2XL U1196 ( .A(B[5]), .B(A[5]), .Z(n632) );
  CND2XL U1197 ( .A(B[37]), .B(A[37]), .Z(n362) );
  CND2XL U1198 ( .A(B[21]), .B(A[21]), .Z(n520) );
  CND2XL U1199 ( .A(B[49]), .B(A[49]), .Z(n236) );
  CND2XL U1200 ( .A(B[51]), .B(A[51]), .Z(n214) );
  CND2XL U1201 ( .A(B[55]), .B(A[55]), .Z(n168) );
  CND2XL U1202 ( .A(B[57]), .B(A[57]), .Z(n146) );
  CND2XL U1203 ( .A(B[53]), .B(A[53]), .Z(n192) );
  CND2XL U1204 ( .A(B[59]), .B(A[59]), .Z(n122) );
  CND2XL U1205 ( .A(B[61]), .B(A[61]), .Z(n98) );
  CND2X1 U1206 ( .A(B[63]), .B(A[63]), .Z(n72) );
  CND2X1 U1207 ( .A(n916), .B(n72), .Z(n7) );
  CANR1XL U1208 ( .A(n74), .B(n917), .C(n75), .Z(n73) );
  CND2XL U1209 ( .A(n915), .B(n85), .Z(n8) );
  CANR1XL U1210 ( .A(n87), .B(n917), .C(n88), .Z(n86) );
  CND2XL U1211 ( .A(n655), .B(n98), .Z(n9) );
  CANR1XL U1212 ( .A(n100), .B(n917), .C(n101), .Z(n99) );
  CND2XL U1213 ( .A(n656), .B(n109), .Z(n10) );
  CANR1XL U1214 ( .A(n111), .B(n917), .C(n112), .Z(n110) );
  CND2XL U1215 ( .A(n657), .B(n122), .Z(n11) );
  CANR1XL U1216 ( .A(n124), .B(n917), .C(n125), .Z(n123) );
  CND2XL U1217 ( .A(n658), .B(n133), .Z(n12) );
  CANR1XL U1218 ( .A(n135), .B(n917), .C(n136), .Z(n134) );
  CND2XL U1219 ( .A(n659), .B(n146), .Z(n13) );
  CANR1XL U1220 ( .A(n148), .B(n917), .C(n149), .Z(n147) );
  CND2XL U1221 ( .A(n660), .B(n155), .Z(n14) );
  CANR1XL U1222 ( .A(n157), .B(n917), .C(n158), .Z(n156) );
  CND2XL U1223 ( .A(n661), .B(n168), .Z(n15) );
  CANR1XL U1224 ( .A(n170), .B(n917), .C(n171), .Z(n169) );
  CND2XL U1225 ( .A(n662), .B(n179), .Z(n16) );
  CANR1XL U1226 ( .A(n181), .B(n917), .C(n182), .Z(n180) );
  CND2XL U1227 ( .A(n663), .B(n192), .Z(n17) );
  CANR1XL U1228 ( .A(n194), .B(n917), .C(n195), .Z(n193) );
  CND2XL U1229 ( .A(n664), .B(n201), .Z(n18) );
  CANR1XL U1230 ( .A(n203), .B(n917), .C(n204), .Z(n202) );
  CND2XL U1231 ( .A(n665), .B(n214), .Z(n19) );
  CANR1XL U1232 ( .A(n216), .B(n917), .C(n217), .Z(n215) );
  CND2XL U1233 ( .A(n666), .B(n223), .Z(n20) );
  CANR1XL U1234 ( .A(n225), .B(n917), .C(n226), .Z(n224) );
  CND2XL U1235 ( .A(n667), .B(n236), .Z(n21) );
  CANR1XL U1236 ( .A(n238), .B(n917), .C(n239), .Z(n237) );
  CND2XL U1237 ( .A(n668), .B(n243), .Z(n22) );
  CANR1XL U1238 ( .A(n245), .B(n917), .C(n246), .Z(n244) );
  CND2XL U1239 ( .A(n669), .B(n256), .Z(n23) );
  CANR1XL U1240 ( .A(n258), .B(n917), .C(n259), .Z(n257) );
  CND2XL U1241 ( .A(n670), .B(n267), .Z(n24) );
  CANR1XL U1242 ( .A(n269), .B(n917), .C(n270), .Z(n268) );
  CND2XL U1243 ( .A(n671), .B(n280), .Z(n25) );
  CANR1XL U1244 ( .A(n282), .B(n917), .C(n283), .Z(n281) );
  CND2XL U1245 ( .A(n672), .B(n289), .Z(n26) );
  CANR1XL U1246 ( .A(n291), .B(n917), .C(n292), .Z(n290) );
  CND2XL U1247 ( .A(n673), .B(n302), .Z(n27) );
  CANR1XL U1248 ( .A(n304), .B(n917), .C(n305), .Z(n303) );
  CND2XL U1249 ( .A(n674), .B(n311), .Z(n28) );
  CANR1XL U1250 ( .A(n313), .B(n917), .C(n314), .Z(n312) );
  CND2XL U1251 ( .A(n675), .B(n324), .Z(n29) );
  CANR1XL U1252 ( .A(n326), .B(n917), .C(n327), .Z(n325) );
  CND2XL U1253 ( .A(n676), .B(n331), .Z(n30) );
  CANR1XL U1254 ( .A(n333), .B(n917), .C(n334), .Z(n332) );
  CND2XL U1255 ( .A(n677), .B(n344), .Z(n31) );
  CANR1XL U1256 ( .A(n346), .B(n917), .C(n347), .Z(n345) );
  CND2XL U1257 ( .A(n678), .B(n351), .Z(n32) );
  CANR1XL U1258 ( .A(n353), .B(n917), .C(n354), .Z(n352) );
  CND2XL U1259 ( .A(n679), .B(n362), .Z(n33) );
  CANR1XL U1260 ( .A(n364), .B(n917), .C(n365), .Z(n363) );
  CND2XL U1261 ( .A(n680), .B(n369), .Z(n34) );
  CANR1XL U1262 ( .A(n375), .B(n917), .C(n376), .Z(n370) );
  CND2XL U1263 ( .A(n681), .B(n382), .Z(n35) );
  CANR1XL U1264 ( .A(n384), .B(n917), .C(n385), .Z(n383) );
  CND2XL U1265 ( .A(n682), .B(n389), .Z(n36) );
  CANR1XL U1266 ( .A(n391), .B(n917), .C(n392), .Z(n390) );
  CND2XL U1267 ( .A(n683), .B(n398), .Z(n37) );
  CANR1XL U1268 ( .A(n684), .B(n917), .C(n401), .Z(n399) );
  CEOXL U1269 ( .A(n62), .B(n617), .Z(SUM[8]) );
  CND2XL U1270 ( .A(n708), .B(n616), .Z(n62) );
  CND2XL U1271 ( .A(n710), .B(n627), .Z(n64) );
  CEOX1 U1272 ( .A(n65), .B(n633), .Z(SUM[5]) );
  CND2XL U1273 ( .A(n711), .B(n632), .Z(n65) );
  CANR1XL U1274 ( .A(n712), .B(n638), .C(n635), .Z(n633) );
  CND2XL U1275 ( .A(n701), .B(n571), .Z(n55) );
  CANR1XL U1276 ( .A(n702), .B(n577), .C(n574), .Z(n572) );
  CND2XL U1277 ( .A(n703), .B(n585), .Z(n57) );
  CANR1XL U1278 ( .A(n704), .B(n591), .C(n588), .Z(n586) );
  CND2XL U1279 ( .A(n705), .B(n601), .Z(n59) );
  CANR1XL U1280 ( .A(n706), .B(n607), .C(n604), .Z(n602) );
  CENX1 U1281 ( .A(n917), .B(n38), .Z(SUM[32]) );
  CND2XL U1282 ( .A(n684), .B(n403), .Z(n38) );
  CND2XL U1283 ( .A(n685), .B(n414), .Z(n39) );
  CANR1XL U1284 ( .A(n416), .B(n562), .C(n417), .Z(n415) );
  CND2XL U1285 ( .A(n686), .B(n425), .Z(n40) );
  CANR1XL U1286 ( .A(n427), .B(n562), .C(n428), .Z(n426) );
  CND2XL U1287 ( .A(n687), .B(n438), .Z(n41) );
  CANR1XL U1288 ( .A(n440), .B(n562), .C(n441), .Z(n439) );
  CND2XL U1289 ( .A(n688), .B(n447), .Z(n42) );
  CANR1XL U1290 ( .A(n449), .B(n562), .C(n450), .Z(n448) );
  CND2XL U1291 ( .A(n689), .B(n460), .Z(n43) );
  CANR1XL U1292 ( .A(n462), .B(n562), .C(n463), .Z(n461) );
  CND2XL U1293 ( .A(n690), .B(n469), .Z(n44) );
  CANR1XL U1294 ( .A(n471), .B(n562), .C(n472), .Z(n470) );
  CND2XL U1295 ( .A(n691), .B(n482), .Z(n45) );
  CND2XL U1296 ( .A(n692), .B(n489), .Z(n46) );
  CND2XL U1297 ( .A(n693), .B(n502), .Z(n47) );
  CND2XL U1298 ( .A(n694), .B(n509), .Z(n48) );
  CANR1XL U1299 ( .A(n511), .B(n562), .C(n512), .Z(n510) );
  CND2XL U1300 ( .A(n695), .B(n520), .Z(n49) );
  CANR1XL U1301 ( .A(n522), .B(n562), .C(n523), .Z(n521) );
  CND2XL U1302 ( .A(n696), .B(n527), .Z(n50) );
  CANR1XL U1303 ( .A(n533), .B(n562), .C(n534), .Z(n528) );
  CND2XL U1304 ( .A(n697), .B(n540), .Z(n51) );
  CANR1XL U1305 ( .A(n542), .B(n562), .C(n543), .Z(n541) );
  CND2XL U1306 ( .A(n698), .B(n547), .Z(n52) );
  CANR1XL U1307 ( .A(n549), .B(n562), .C(n550), .Z(n548) );
  CND2XL U1308 ( .A(n699), .B(n556), .Z(n53) );
  CANR1XL U1309 ( .A(n700), .B(n562), .C(n559), .Z(n557) );
  CENX1 U1310 ( .A(n562), .B(n54), .Z(SUM[16]) );
  CND2XL U1311 ( .A(n700), .B(n561), .Z(n54) );
  CENX1 U1312 ( .A(n577), .B(n56), .Z(SUM[14]) );
  CND2XL U1313 ( .A(n702), .B(n576), .Z(n56) );
  CENX1 U1314 ( .A(n591), .B(n58), .Z(SUM[12]) );
  CND2XL U1315 ( .A(n704), .B(n590), .Z(n58) );
  CENX1 U1316 ( .A(n607), .B(n60), .Z(SUM[10]) );
  CND2XL U1317 ( .A(n706), .B(n606), .Z(n60) );
  CENX1 U1318 ( .A(n625), .B(n63), .Z(SUM[7]) );
  CND2XL U1319 ( .A(n709), .B(n624), .Z(n63) );
  COND1XL U1320 ( .A(n626), .B(n628), .C(n627), .Z(n625) );
  CENX1 U1321 ( .A(n614), .B(n61), .Z(SUM[9]) );
  CND2XL U1322 ( .A(n707), .B(n613), .Z(n61) );
  COND1XL U1323 ( .A(n615), .B(n617), .C(n616), .Z(n614) );
  CENX1 U1324 ( .A(n638), .B(n66), .Z(SUM[4]) );
  CND2XL U1325 ( .A(n712), .B(n637), .Z(n66) );
  CENX1 U1326 ( .A(n644), .B(n67), .Z(SUM[3]) );
  CND2XL U1327 ( .A(n713), .B(n643), .Z(n67) );
  COND1XL U1328 ( .A(n645), .B(n647), .C(n646), .Z(n644) );
  CEOX1 U1329 ( .A(n68), .B(n647), .Z(SUM[2]) );
  CND2XL U1330 ( .A(n714), .B(n646), .Z(n68) );
  CEOXL U1331 ( .A(n652), .B(n69), .Z(SUM[1]) );
  CND2XL U1332 ( .A(n715), .B(n650), .Z(n69) );
  CANR1X2 U1333 ( .A(n334), .B(n249), .C(n250), .Z(n3) );
  CIVX2 U1334 ( .A(n96), .Z(n94) );
  CIVX2 U1335 ( .A(n95), .Z(n93) );
  CIVX2 U1336 ( .A(n85), .Z(n83) );
  CIVX2 U1337 ( .A(n649), .Z(n715) );
  CIVX2 U1338 ( .A(n645), .Z(n714) );
  CIVX2 U1339 ( .A(n642), .Z(n713) );
  CIVX2 U1340 ( .A(n631), .Z(n711) );
  CIVX2 U1341 ( .A(n626), .Z(n710) );
  CIVX2 U1342 ( .A(n623), .Z(n709) );
  CIVX2 U1343 ( .A(n615), .Z(n708) );
  CIVX2 U1344 ( .A(n612), .Z(n707) );
  CIVX2 U1345 ( .A(n600), .Z(n705) );
  CIVX2 U1346 ( .A(n584), .Z(n703) );
  CIVX2 U1347 ( .A(n570), .Z(n701) );
  CIVX2 U1348 ( .A(n555), .Z(n699) );
  CIVX2 U1349 ( .A(n544), .Z(n698) );
  CIVX2 U1350 ( .A(n539), .Z(n697) );
  CIVX2 U1351 ( .A(n524), .Z(n696) );
  CIVX2 U1352 ( .A(n519), .Z(n695) );
  CIVX2 U1353 ( .A(n506), .Z(n694) );
  CIVX2 U1354 ( .A(n501), .Z(n693) );
  CIVX2 U1355 ( .A(n486), .Z(n692) );
  CIVX2 U1356 ( .A(n481), .Z(n691) );
  CIVX2 U1357 ( .A(n459), .Z(n689) );
  CIVX2 U1358 ( .A(n437), .Z(n687) );
  CIVX2 U1359 ( .A(n422), .Z(n686) );
  CIVX2 U1360 ( .A(n413), .Z(n685) );
  CIVX2 U1361 ( .A(n397), .Z(n683) );
  CIVX2 U1362 ( .A(n386), .Z(n682) );
  CIVX2 U1363 ( .A(n381), .Z(n681) );
  CIVX2 U1364 ( .A(n366), .Z(n680) );
  CIVX2 U1365 ( .A(n361), .Z(n679) );
  CIVX2 U1366 ( .A(n348), .Z(n678) );
  CIVX2 U1367 ( .A(n343), .Z(n677) );
  CIVX2 U1368 ( .A(n328), .Z(n676) );
  CIVX2 U1369 ( .A(n323), .Z(n675) );
  CIVX2 U1370 ( .A(n301), .Z(n673) );
  CIVX2 U1371 ( .A(n279), .Z(n671) );
  CIVX2 U1372 ( .A(n264), .Z(n670) );
  CIVX2 U1373 ( .A(n255), .Z(n669) );
  CIVX2 U1374 ( .A(n240), .Z(n668) );
  CIVX2 U1375 ( .A(n235), .Z(n667) );
  CIVX2 U1376 ( .A(n213), .Z(n665) );
  CIVX2 U1377 ( .A(n191), .Z(n663) );
  CIVX2 U1378 ( .A(n176), .Z(n662) );
  CIVX2 U1379 ( .A(n167), .Z(n661) );
  CIVX2 U1380 ( .A(n145), .Z(n659) );
  CIVX2 U1381 ( .A(n130), .Z(n658) );
  CIVX2 U1382 ( .A(n121), .Z(n657) );
  CIVX2 U1383 ( .A(n106), .Z(n656) );
  CIVX2 U1384 ( .A(n97), .Z(n655) );
  CIVX2 U1385 ( .A(n648), .Z(n647) );
  CIVX2 U1386 ( .A(n639), .Z(n638) );
  CIVX2 U1387 ( .A(n637), .Z(n635) );
  CIVX2 U1388 ( .A(n636), .Z(n712) );
  CIVX2 U1389 ( .A(n618), .Z(n617) );
  CIVX2 U1390 ( .A(n611), .Z(n609) );
  CIVX2 U1391 ( .A(n610), .Z(n608) );
  CIVX2 U1392 ( .A(n606), .Z(n604) );
  CIVX2 U1393 ( .A(n605), .Z(n706) );
  CIVX2 U1394 ( .A(n593), .Z(n595) );
  CIVX2 U1395 ( .A(n592), .Z(n594) );
  CIVX2 U1396 ( .A(n590), .Z(n588) );
  CIVX2 U1397 ( .A(n589), .Z(n704) );
  CIVX2 U1398 ( .A(n576), .Z(n574) );
  CIVX2 U1399 ( .A(n575), .Z(n702) );
  CIVX2 U1400 ( .A(n561), .Z(n559) );
  CIVX2 U1401 ( .A(n560), .Z(n700) );
  CIVX2 U1402 ( .A(n550), .Z(n552) );
  CIVX2 U1403 ( .A(n532), .Z(n534) );
  CIVX2 U1404 ( .A(n531), .Z(n533) );
  CIVX2 U1405 ( .A(n514), .Z(n512) );
  CIVX2 U1406 ( .A(n513), .Z(n511) );
  CIVX2 U1407 ( .A(n492), .Z(n494) );
  CIVX2 U1408 ( .A(n491), .Z(n493) );
  CIVX2 U1409 ( .A(n476), .Z(n474) );
  CIVX2 U1410 ( .A(n475), .Z(n473) );
  CIVX2 U1411 ( .A(n469), .Z(n467) );
  CIVX2 U1412 ( .A(n468), .Z(n690) );
  CIVX2 U1413 ( .A(n452), .Z(n454) );
  CIVX2 U1414 ( .A(n451), .Z(n453) );
  CIVX2 U1415 ( .A(n447), .Z(n445) );
  CIVX2 U1416 ( .A(n446), .Z(n688) );
  CIVX2 U1417 ( .A(n432), .Z(n434) );
  CIVX2 U1418 ( .A(n403), .Z(n401) );
  CIVX2 U1419 ( .A(n402), .Z(n684) );
  CIVX2 U1420 ( .A(n392), .Z(n394) );
  CIVX2 U1421 ( .A(n374), .Z(n376) );
  CIVX2 U1422 ( .A(n373), .Z(n375) );
  CIVX2 U1423 ( .A(n356), .Z(n354) );
  CIVX2 U1424 ( .A(n355), .Z(n353) );
  CIVX2 U1425 ( .A(n334), .Z(n336) );
  CIVX2 U1426 ( .A(n333), .Z(n335) );
  CIVX2 U1427 ( .A(n318), .Z(n316) );
  CIVX2 U1428 ( .A(n317), .Z(n315) );
  CIVX2 U1429 ( .A(n311), .Z(n309) );
  CIVX2 U1430 ( .A(n310), .Z(n674) );
  CIVX2 U1431 ( .A(n294), .Z(n296) );
  CIVX2 U1432 ( .A(n293), .Z(n295) );
  CIVX2 U1433 ( .A(n289), .Z(n287) );
  CIVX2 U1434 ( .A(n288), .Z(n672) );
  CIVX2 U1435 ( .A(n274), .Z(n276) );
  CIVX2 U1436 ( .A(n3), .Z(n246) );
  CIVX2 U1437 ( .A(n4), .Z(n245) );
  CIVX2 U1438 ( .A(n230), .Z(n228) );
  CIVX2 U1439 ( .A(n229), .Z(n227) );
  CIVX2 U1440 ( .A(n223), .Z(n221) );
  CIVX2 U1441 ( .A(n222), .Z(n666) );
  CIVX2 U1442 ( .A(n206), .Z(n208) );
  CIVX2 U1443 ( .A(n205), .Z(n207) );
  CIVX2 U1444 ( .A(n201), .Z(n199) );
  CIVX2 U1445 ( .A(n200), .Z(n664) );
  CIVX2 U1446 ( .A(n186), .Z(n188) );
  CIVX2 U1447 ( .A(n5), .Z(n160) );
  CIVX2 U1448 ( .A(n6), .Z(n159) );
  CIVX2 U1449 ( .A(n155), .Z(n153) );
  CIVX2 U1450 ( .A(n154), .Z(n660) );
  CIVX2 U1451 ( .A(n140), .Z(n142) );
  CIVX2 U1452 ( .A(n118), .Z(n116) );
  CIVX2 U1453 ( .A(n117), .Z(n115) );
  CIVX2 U1454 ( .A(n70), .Z(SUM[0]) );
endmodule


module sfilt_DW01_add_3 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31, n32,
         n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n68, n69, n70, n71, n72, n73, n74, n75, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108,
         n109, n110, n111, n112, n113, n114, n115, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n216, n217, n218, n219, n220, n221, n222,
         n223, n225, n226, n227, n228, n229, n230, n231, n232, n233, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n260, n261, n262, n263, n264, n265, n266, n267, n269, n270,
         n271;
  assign n13 = A[56];
  assign n17 = A[55];
  assign n24 = A[54];
  assign n28 = A[53];
  assign n33 = A[52];
  assign n37 = A[51];
  assign n43 = A[50];
  assign n47 = A[49];
  assign n52 = A[48];
  assign n56 = A[47];
  assign n64 = A[46];
  assign n68 = A[45];
  assign n73 = A[44];
  assign n77 = A[43];
  assign n83 = A[42];
  assign n87 = A[41];
  assign n92 = A[40];
  assign n96 = A[39];
  assign n104 = A[38];
  assign n108 = A[37];
  assign n113 = A[36];
  assign n117 = A[35];
  assign n123 = A[34];
  assign n127 = A[33];
  assign n132 = A[32];
  assign n135 = A[31];
  assign n143 = A[30];
  assign n146 = A[29];
  assign n150 = A[28];
  assign n153 = A[27];
  assign n160 = A[26];
  assign n163 = A[25];
  assign n167 = A[24];
  assign n170 = A[23];
  assign n177 = A[22];
  assign n180 = A[21];
  assign n184 = A[20];
  assign n187 = A[19];
  assign n194 = A[18];
  assign n197 = A[17];
  assign n201 = A[16];
  assign n205 = A[15];
  assign n212 = A[14];
  assign n216 = A[13];
  assign n221 = A[12];
  assign n225 = A[11];
  assign n231 = A[10];
  assign n235 = A[9];
  assign n240 = A[8];
  assign n243 = A[7];
  assign n249 = A[6];
  assign n252 = A[5];
  assign n256 = A[4];
  assign n260 = A[3];
  assign n265 = A[2];
  assign n269 = A[1];

  CHA1X1 U2 ( .A(A[62]), .B(n4), .CO(n3), .S(SUM[62]) );
  CHA1X1 U3 ( .A(A[61]), .B(n5), .CO(n4), .S(SUM[61]) );
  CHA1X1 U4 ( .A(A[60]), .B(n6), .CO(n5), .S(SUM[60]) );
  CHA1X1 U5 ( .A(A[59]), .B(n7), .CO(n6), .S(SUM[59]) );
  CHA1X1 U6 ( .A(A[58]), .B(n8), .CO(n7), .S(SUM[58]) );
  CHA1X1 U7 ( .A(A[57]), .B(n9), .CO(n8), .S(SUM[57]) );
  CIVXL U334 ( .A(n138), .Z(n137) );
  CIVX1 U335 ( .A(n208), .Z(n207) );
  CIVXL U336 ( .A(n246), .Z(n245) );
  CIVX1 U337 ( .A(n263), .Z(n262) );
  CNR2XL U338 ( .A(n1), .B(n270), .Z(n267) );
  CEOXL U339 ( .A(n1), .B(n270), .Z(SUM[1]) );
  CNR2XL U340 ( .A(A[0]), .B(B[0]), .Z(n271) );
  CNR2X1 U341 ( .A(n155), .B(n149), .Z(n148) );
  CNR2X1 U342 ( .A(n172), .B(n166), .Z(n165) );
  CNR2X1 U343 ( .A(n189), .B(n183), .Z(n182) );
  CNR2X1 U344 ( .A(n19), .B(n18), .Z(n15) );
  CNR2X1 U345 ( .A(n30), .B(n29), .Z(n26) );
  CNR2X1 U346 ( .A(n40), .B(n38), .Z(n35) );
  CNR2X1 U347 ( .A(n49), .B(n48), .Z(n45) );
  CNR2X1 U348 ( .A(n70), .B(n69), .Z(n66) );
  CNR2X1 U349 ( .A(n80), .B(n78), .Z(n75) );
  CNR2X1 U350 ( .A(n89), .B(n88), .Z(n85) );
  CNR2X1 U351 ( .A(n110), .B(n109), .Z(n106) );
  CNR2X1 U352 ( .A(n129), .B(n128), .Z(n125) );
  CNR2X1 U353 ( .A(n172), .B(n157), .Z(n156) );
  CNR2X1 U354 ( .A(n207), .B(n174), .Z(n173) );
  CNR2X1 U355 ( .A(n207), .B(n191), .Z(n190) );
  CND2X1 U356 ( .A(n58), .B(n20), .Z(n19) );
  CND2X1 U357 ( .A(n39), .B(n31), .Z(n30) );
  CND2X1 U358 ( .A(n58), .B(n50), .Z(n49) );
  CND2X1 U359 ( .A(n79), .B(n71), .Z(n70) );
  CND2X1 U360 ( .A(n98), .B(n90), .Z(n89) );
  CND2X1 U361 ( .A(n119), .B(n111), .Z(n110) );
  CND2X1 U362 ( .A(n137), .B(n130), .Z(n129) );
  CND2X1 U363 ( .A(n139), .B(n208), .Z(n138) );
  CNR2X1 U364 ( .A(n174), .B(n140), .Z(n139) );
  CND2X1 U365 ( .A(n158), .B(n141), .Z(n140) );
  CNR2X1 U366 ( .A(n149), .B(n142), .Z(n141) );
  CND2X1 U367 ( .A(n58), .B(n41), .Z(n40) );
  CND2X1 U368 ( .A(n137), .B(n60), .Z(n59) );
  CND2X1 U369 ( .A(n98), .B(n81), .Z(n80) );
  CND2X1 U370 ( .A(n137), .B(n100), .Z(n99) );
  CND2X1 U371 ( .A(n137), .B(n121), .Z(n120) );
  CNR2X1 U372 ( .A(n207), .B(n200), .Z(n199) );
  CNR2X1 U373 ( .A(n262), .B(n255), .Z(n254) );
  CNR2X1 U374 ( .A(n59), .B(n57), .Z(n54) );
  CNR2X1 U375 ( .A(n99), .B(n97), .Z(n94) );
  CNR2X1 U376 ( .A(n120), .B(n118), .Z(n115) );
  CNR2X1 U377 ( .A(n207), .B(n206), .Z(n203) );
  CNR2X1 U378 ( .A(n218), .B(n217), .Z(n214) );
  CNR2X1 U379 ( .A(n228), .B(n226), .Z(n223) );
  CNR2X1 U380 ( .A(n237), .B(n236), .Z(n233) );
  CNR2X1 U381 ( .A(n262), .B(n261), .Z(n258) );
  CND2X1 U382 ( .A(n227), .B(n219), .Z(n218) );
  CND2X1 U383 ( .A(n245), .B(n238), .Z(n237) );
  CND2X1 U384 ( .A(n245), .B(n229), .Z(n228) );
  CENX1 U385 ( .A(n15), .B(n14), .Z(SUM[56]) );
  CEOX1 U386 ( .A(n18), .B(n19), .Z(SUM[55]) );
  CENX1 U387 ( .A(n26), .B(n25), .Z(SUM[54]) );
  CEOX1 U388 ( .A(n29), .B(n30), .Z(SUM[53]) );
  CENX1 U389 ( .A(n35), .B(n34), .Z(SUM[52]) );
  CENX1 U390 ( .A(n39), .B(n38), .Z(SUM[51]) );
  CENX1 U391 ( .A(n45), .B(n44), .Z(SUM[50]) );
  CEOX1 U392 ( .A(n48), .B(n49), .Z(SUM[49]) );
  CENX1 U393 ( .A(n58), .B(n57), .Z(SUM[47]) );
  CENX1 U394 ( .A(n66), .B(n65), .Z(SUM[46]) );
  CEOX1 U395 ( .A(n69), .B(n70), .Z(SUM[45]) );
  CENX1 U396 ( .A(n75), .B(n74), .Z(SUM[44]) );
  CENX1 U397 ( .A(n79), .B(n78), .Z(SUM[43]) );
  CENX1 U398 ( .A(n85), .B(n84), .Z(SUM[42]) );
  CEOX1 U399 ( .A(n88), .B(n89), .Z(SUM[41]) );
  CENX1 U400 ( .A(n106), .B(n105), .Z(SUM[38]) );
  CEOX1 U401 ( .A(n109), .B(n110), .Z(SUM[37]) );
  CENX1 U402 ( .A(n125), .B(n124), .Z(SUM[34]) );
  CEOX1 U403 ( .A(n144), .B(n145), .Z(SUM[30]) );
  CENX1 U404 ( .A(n148), .B(n147), .Z(SUM[29]) );
  CEOX1 U405 ( .A(n151), .B(n152), .Z(SUM[28]) );
  CEOX1 U406 ( .A(n154), .B(n155), .Z(SUM[27]) );
  CEOX1 U407 ( .A(n161), .B(n162), .Z(SUM[26]) );
  CENX1 U408 ( .A(n165), .B(n164), .Z(SUM[25]) );
  CEOX1 U409 ( .A(n178), .B(n179), .Z(SUM[22]) );
  CENX1 U410 ( .A(n182), .B(n181), .Z(SUM[21]) );
  CND2X1 U411 ( .A(A[0]), .B(B[0]), .Z(n1) );
  CNR2X1 U412 ( .A(n239), .B(n230), .Z(n229) );
  CND2X1 U413 ( .A(n235), .B(n231), .Z(n230) );
  CNR2X1 U414 ( .A(n131), .B(n122), .Z(n121) );
  CND2X1 U415 ( .A(n127), .B(n123), .Z(n122) );
  CNR2X1 U416 ( .A(n91), .B(n82), .Z(n81) );
  CND2X1 U417 ( .A(n87), .B(n83), .Z(n82) );
  CNR2X1 U418 ( .A(n51), .B(n42), .Z(n41) );
  CND2X1 U419 ( .A(n47), .B(n43), .Z(n42) );
  CNR2X1 U420 ( .A(n101), .B(n61), .Z(n60) );
  CND2X1 U421 ( .A(n81), .B(n62), .Z(n61) );
  CNR2X1 U422 ( .A(n72), .B(n63), .Z(n62) );
  CND2X1 U423 ( .A(n68), .B(n64), .Z(n63) );
  CNR2X1 U424 ( .A(n264), .B(n1), .Z(n263) );
  CND2X1 U425 ( .A(n269), .B(n265), .Z(n264) );
  CNR2X1 U426 ( .A(n209), .B(n246), .Z(n208) );
  CND2X1 U427 ( .A(n229), .B(n210), .Z(n209) );
  CNR2X1 U428 ( .A(n220), .B(n211), .Z(n210) );
  CND2X1 U429 ( .A(n216), .B(n212), .Z(n211) );
  CNR2X1 U430 ( .A(n166), .B(n159), .Z(n158) );
  CND2X1 U431 ( .A(n163), .B(n160), .Z(n159) );
  CNR2X1 U432 ( .A(n10), .B(n138), .Z(n9) );
  CND2X1 U433 ( .A(n60), .B(n11), .Z(n10) );
  CNR2X1 U434 ( .A(n21), .B(n12), .Z(n11) );
  CND2X1 U435 ( .A(n260), .B(n256), .Z(n255) );
  CND2X1 U436 ( .A(n205), .B(n201), .Z(n200) );
  CND2X1 U437 ( .A(n187), .B(n184), .Z(n183) );
  CND2X1 U438 ( .A(n170), .B(n167), .Z(n166) );
  CND2X1 U439 ( .A(n153), .B(n150), .Z(n149) );
  CND2X1 U440 ( .A(n192), .B(n175), .Z(n174) );
  CNR2X1 U441 ( .A(n183), .B(n176), .Z(n175) );
  CND2X1 U442 ( .A(n180), .B(n177), .Z(n176) );
  CND2X1 U443 ( .A(n247), .B(n263), .Z(n246) );
  CNR2X1 U444 ( .A(n255), .B(n248), .Z(n247) );
  CND2X1 U445 ( .A(n252), .B(n249), .Z(n248) );
  CND2X1 U446 ( .A(n243), .B(n240), .Z(n239) );
  CND2X1 U447 ( .A(n225), .B(n221), .Z(n220) );
  CND2X1 U448 ( .A(n135), .B(n132), .Z(n131) );
  CND2X1 U449 ( .A(n117), .B(n113), .Z(n112) );
  CND2X1 U450 ( .A(n96), .B(n92), .Z(n91) );
  CND2X1 U451 ( .A(n77), .B(n73), .Z(n72) );
  CND2X1 U452 ( .A(n56), .B(n52), .Z(n51) );
  CND2X1 U453 ( .A(n37), .B(n33), .Z(n32) );
  CND2X1 U454 ( .A(n121), .B(n102), .Z(n101) );
  CNR2X1 U455 ( .A(n112), .B(n103), .Z(n102) );
  CND2X1 U456 ( .A(n108), .B(n104), .Z(n103) );
  CND2X1 U457 ( .A(n41), .B(n22), .Z(n21) );
  CNR2X1 U458 ( .A(n32), .B(n23), .Z(n22) );
  CND2X1 U459 ( .A(n28), .B(n24), .Z(n23) );
  CND2X1 U460 ( .A(n148), .B(n146), .Z(n145) );
  CND2X1 U461 ( .A(n156), .B(n153), .Z(n152) );
  CND2X1 U462 ( .A(n165), .B(n163), .Z(n162) );
  CND2X1 U463 ( .A(n182), .B(n180), .Z(n179) );
  CEOX1 U464 ( .A(A[63]), .B(n3), .Z(SUM[63]) );
  CND2X1 U465 ( .A(n146), .B(n143), .Z(n142) );
  CNR2X1 U466 ( .A(n200), .B(n193), .Z(n192) );
  CND2X1 U467 ( .A(n197), .B(n194), .Z(n193) );
  CND2X1 U468 ( .A(n17), .B(n13), .Z(n12) );
  CENX1 U469 ( .A(n54), .B(n53), .Z(SUM[48]) );
  CENX1 U470 ( .A(n94), .B(n93), .Z(SUM[40]) );
  CENX1 U471 ( .A(n98), .B(n97), .Z(SUM[39]) );
  CENX1 U472 ( .A(n115), .B(n114), .Z(SUM[36]) );
  CENX1 U473 ( .A(n119), .B(n118), .Z(SUM[35]) );
  CEOX1 U474 ( .A(n128), .B(n129), .Z(SUM[33]) );
  CEOX1 U475 ( .A(n133), .B(n134), .Z(SUM[32]) );
  CENX1 U476 ( .A(n137), .B(n136), .Z(SUM[31]) );
  CEOX1 U477 ( .A(n168), .B(n169), .Z(SUM[24]) );
  CEOX1 U478 ( .A(n171), .B(n172), .Z(SUM[23]) );
  CEOX1 U479 ( .A(n185), .B(n186), .Z(SUM[20]) );
  CEOX1 U480 ( .A(n188), .B(n189), .Z(SUM[19]) );
  CEOX1 U481 ( .A(n195), .B(n196), .Z(SUM[18]) );
  CENX1 U482 ( .A(n199), .B(n198), .Z(SUM[17]) );
  CENX1 U483 ( .A(n203), .B(n202), .Z(SUM[16]) );
  CEOX1 U484 ( .A(n206), .B(n207), .Z(SUM[15]) );
  CENX1 U485 ( .A(n214), .B(n213), .Z(SUM[14]) );
  CEOX1 U486 ( .A(n217), .B(n218), .Z(SUM[13]) );
  CENX1 U487 ( .A(n223), .B(n222), .Z(SUM[12]) );
  CENX1 U488 ( .A(n227), .B(n226), .Z(SUM[11]) );
  CENX1 U489 ( .A(n233), .B(n232), .Z(SUM[10]) );
  CEOX1 U490 ( .A(n236), .B(n237), .Z(SUM[9]) );
  CEOX1 U491 ( .A(n241), .B(n242), .Z(SUM[8]) );
  CENX1 U492 ( .A(n245), .B(n244), .Z(SUM[7]) );
  CEOX1 U493 ( .A(n250), .B(n251), .Z(SUM[6]) );
  CENX1 U494 ( .A(n258), .B(n257), .Z(SUM[4]) );
  CENX1 U495 ( .A(n267), .B(n266), .Z(SUM[2]) );
  CENX1 U496 ( .A(n254), .B(n253), .Z(SUM[5]) );
  CND2X1 U497 ( .A(n137), .B(n135), .Z(n134) );
  CND2X1 U498 ( .A(n173), .B(n170), .Z(n169) );
  CND2X1 U499 ( .A(n190), .B(n187), .Z(n186) );
  CND2X1 U500 ( .A(n199), .B(n197), .Z(n196) );
  CND2X1 U501 ( .A(n245), .B(n243), .Z(n242) );
  CND2X1 U502 ( .A(n254), .B(n252), .Z(n251) );
  CEOX1 U503 ( .A(n261), .B(n262), .Z(SUM[3]) );
  CND2IX1 U504 ( .B(n271), .A(n1), .Z(n2) );
  CIVX2 U505 ( .A(n99), .Z(n98) );
  CIVX2 U506 ( .A(n96), .Z(n97) );
  CIVX2 U507 ( .A(n92), .Z(n93) );
  CIVX2 U508 ( .A(n91), .Z(n90) );
  CIVX2 U509 ( .A(n87), .Z(n88) );
  CIVX2 U510 ( .A(n83), .Z(n84) );
  CIVX2 U511 ( .A(n80), .Z(n79) );
  CIVX2 U512 ( .A(n77), .Z(n78) );
  CIVX2 U513 ( .A(n73), .Z(n74) );
  CIVX2 U514 ( .A(n72), .Z(n71) );
  CIVX2 U515 ( .A(n68), .Z(n69) );
  CIVX2 U516 ( .A(n64), .Z(n65) );
  CIVX2 U517 ( .A(n59), .Z(n58) );
  CIVX2 U518 ( .A(n56), .Z(n57) );
  CIVX2 U519 ( .A(n52), .Z(n53) );
  CIVX2 U520 ( .A(n51), .Z(n50) );
  CIVX2 U521 ( .A(n47), .Z(n48) );
  CIVX2 U522 ( .A(n43), .Z(n44) );
  CIVX2 U523 ( .A(n40), .Z(n39) );
  CIVX2 U524 ( .A(n37), .Z(n38) );
  CIVX2 U525 ( .A(n33), .Z(n34) );
  CIVX2 U526 ( .A(n32), .Z(n31) );
  CIVX2 U527 ( .A(n28), .Z(n29) );
  CIVX2 U528 ( .A(n269), .Z(n270) );
  CIVX2 U529 ( .A(n265), .Z(n266) );
  CIVX2 U530 ( .A(n260), .Z(n261) );
  CIVX2 U531 ( .A(n256), .Z(n257) );
  CIVX2 U532 ( .A(n252), .Z(n253) );
  CIVX2 U533 ( .A(n249), .Z(n250) );
  CIVX2 U534 ( .A(n24), .Z(n25) );
  CIVX2 U535 ( .A(n243), .Z(n244) );
  CIVX2 U536 ( .A(n240), .Z(n241) );
  CIVX2 U537 ( .A(n239), .Z(n238) );
  CIVX2 U538 ( .A(n235), .Z(n236) );
  CIVX2 U539 ( .A(n231), .Z(n232) );
  CIVX2 U540 ( .A(n228), .Z(n227) );
  CIVX2 U541 ( .A(n225), .Z(n226) );
  CIVX2 U542 ( .A(n221), .Z(n222) );
  CIVX2 U543 ( .A(n220), .Z(n219) );
  CIVX2 U544 ( .A(n216), .Z(n217) );
  CIVX2 U545 ( .A(n212), .Z(n213) );
  CIVX2 U546 ( .A(n205), .Z(n206) );
  CIVX2 U547 ( .A(n201), .Z(n202) );
  CIVX2 U548 ( .A(n21), .Z(n20) );
  CIVX2 U549 ( .A(n197), .Z(n198) );
  CIVX2 U550 ( .A(n194), .Z(n195) );
  CIVX2 U551 ( .A(n192), .Z(n191) );
  CIVX2 U552 ( .A(n190), .Z(n189) );
  CIVX2 U553 ( .A(n187), .Z(n188) );
  CIVX2 U554 ( .A(n184), .Z(n185) );
  CIVX2 U555 ( .A(n180), .Z(n181) );
  CIVX2 U556 ( .A(n177), .Z(n178) );
  CIVX2 U557 ( .A(n173), .Z(n172) );
  CIVX2 U558 ( .A(n170), .Z(n171) );
  CIVX2 U559 ( .A(n167), .Z(n168) );
  CIVX2 U560 ( .A(n163), .Z(n164) );
  CIVX2 U561 ( .A(n160), .Z(n161) );
  CIVX2 U562 ( .A(n17), .Z(n18) );
  CIVX2 U563 ( .A(n158), .Z(n157) );
  CIVX2 U564 ( .A(n156), .Z(n155) );
  CIVX2 U565 ( .A(n153), .Z(n154) );
  CIVX2 U566 ( .A(n150), .Z(n151) );
  CIVX2 U567 ( .A(n146), .Z(n147) );
  CIVX2 U568 ( .A(n143), .Z(n144) );
  CIVX2 U569 ( .A(n13), .Z(n14) );
  CIVX2 U570 ( .A(n135), .Z(n136) );
  CIVX2 U571 ( .A(n132), .Z(n133) );
  CIVX2 U572 ( .A(n131), .Z(n130) );
  CIVX2 U573 ( .A(n127), .Z(n128) );
  CIVX2 U574 ( .A(n123), .Z(n124) );
  CIVX2 U575 ( .A(n120), .Z(n119) );
  CIVX2 U576 ( .A(n117), .Z(n118) );
  CIVX2 U577 ( .A(n113), .Z(n114) );
  CIVX2 U578 ( .A(n112), .Z(n111) );
  CIVX2 U579 ( .A(n108), .Z(n109) );
  CIVX2 U580 ( .A(n104), .Z(n105) );
  CIVX2 U581 ( .A(n101), .Z(n100) );
  CIVX2 U582 ( .A(n2), .Z(SUM[0]) );
endmodule


module sfilt_DW_mult_tc_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n9, n12, n18, n21, n24, n27, n30, n33, n36, n39, n42, n45,
         n48, n54, n57, n63, n66, n72, n75, n78, n81, n84, n87, n90, n93, n99,
         n102, n105, n108, n111, n114, n117, n120, n126, n129, n132, n135,
         n136, n141, n144, n145, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n173, n174, n175, n176, n177, n178, n179, n181, n184,
         n185, n186, n187, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n212, n213, n214, n222, n224, n241, n246, n247, n248,
         n249, n254, n255, n256, n258, n260, n261, n262, n264, n265, n266,
         n267, n268, n269, n272, n273, n274, n275, n277, n279, n280, n281,
         n282, n283, n286, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n301, n302, n303, n304, n306, n308, n309, n310, n314, n316,
         n317, n318, n319, n320, n323, n324, n327, n328, n329, n330, n331,
         n332, n333, n334, n340, n342, n343, n344, n345, n349, n351, n352,
         n353, n355, n356, n360, n362, n363, n364, n365, n366, n369, n370,
         n371, n372, n373, n377, n378, n379, n380, n381, n383, n384, n385,
         n386, n387, n388, n389, n392, n393, n394, n395, n396, n397, n402,
         n403, n404, n405, n406, n408, n409, n410, n411, n413, n414, n415,
         n416, n417, n418, n419, n423, n425, n426, n427, n428, n432, n434,
         n435, n438, n440, n444, n445, n448, n449, n450, n451, n452, n456,
         n458, n459, n460, n461, n462, n467, n468, n469, n470, n472, n482,
         n485, n486, n487, n488, n489, n490, n491, n494, n495, n496, n497,
         n504, n505, n506, n507, n508, n510, n511, n512, n513, n514, n516,
         n520, n521, n522, n523, n524, n525, n526, n528, n529, n530, n531,
         n532, n534, n535, n540, n541, n542, n543, n554, n555, n560, n564,
         n569, n571, n572, n574, n578, n582, n583, n584, n585, n586, n590,
         n593, n594, n595, n596, n597, n601, n603, n604, n605, n611, n612,
         n614, n616, n618, n619, n620, n621, n622, n623, n626, n627, n628,
         n629, n632, n633, n634, n635, n636, n637, n639, n641, n642, n643,
         n644, n649, n650, n651, n654, n656, n657, n658, n659, n660, n661,
         n662, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n681, n683, n684, n686, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n704, n706, n707, n708, n709, n710, n712, n714,
         n718, n720, n721, n722, n723, n724, n726, n728, n729, n731, n735,
         n736, n738, n739, n741, n744, n745, n746, n747, n748, n751, n753,
         n756, n757, n758, n766, n767, n770, n773, n774, n776, n779, n780,
         n781, n784, n785, n786, n788, n791, n794, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1336, n1338, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1359, n1370, n1371, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1386, n1389, n1390, n1391, n1392, n1393,
         n1397, n1402, n1403, n1406, n1407, n1409, n1412, n1413, n1414, n1415,
         n1417, n1418, n1419, n1420, n1421, n1423, n1426, n1427, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2070, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2812, n2813, n2814, n2815, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2826, n2827, net15997, net15995,
         net16027, net16037, net16065, net16063, net16059, net16069, net16067,
         net16089, net16087, net16083, net16093, net16091, net16109, net16107,
         net16544, net16548, net16550, net16558, net16570, net16759, net16771,
         net16772, net16784, net16788, net16791, net16793, net16802, net16801,
         net16800, net16812, net16817, net16816, net16824, net16839, net16838,
         net16844, net16843, net16850, net16849, net18254, net18260, net18422,
         net18543, net18593, net18592, net18609, net18608, net18607, net18618,
         net18643, net18670, net18731, net18730, net18736, net18743, net18742,
         net18817, net18875, net18897, net18905, net18937, net18936, net18948,
         net18953, net18982, net18981, net19016, net19048, net19047, net19061,
         net19060, net19076, net19089, net19108, net19122, net19151, net19168,
         net19200, net19205, net19204, net19203, net19269, net19268, net19267,
         net19292, net19307, net19316, net19384, net19388, net19401, net19409,
         net19417, net19462, net19505, net19508, net19517, net19518, net19521,
         net19522, net19531, net19530, net19555, n2825, n2690, n2691, n480,
         net19127, net18739, net18620, n764, n763, n559, n556, n552, n551,
         n1305, n1304, net18420, n218, n216, n150, net19133, n765, n573, n568,
         n562, n1361, n2505, n2504, n2164, n2009, n1979, n1429, n1428, n546,
         n515, n499, n484, n483, n481, n479, n478, n225, n223, n221, n220,
         n219, net18451, n630, n579, n577, n576, n548, n547, net18816, n2069,
         n1408, n1396, n1385, n1384, n1373, n1372, n1367, n1366, n1363, n1362,
         n1360, n1337, n1333, n1332, n2041, n1451, net19500, n2226, n2195,
         n2040, n1949, n1920, n1861, n1433, n1432, n1431, n1430, n1399, n1398,
         net16644, n96, n2163, n1948, n1919, n1450, n1425, n1424, n1416, n1405,
         n1404, n1395, n1394, n1388, n1365, n1364, n1339, n1335, n1334,
         net16658, n2350, n2349, n2071, n1890, n1832, n1726, n1435, n1434,
         n1422, n1411, n1410, n1401, n1400, n1369, n1368, net18421, n795, n229,
         n227, n151, net19465, n447, n359, n354, n253, n244, n242, n236, n233,
         n232, n231, n230, n149, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n57 = a[13];
  assign n66 = a[15];
  assign n75 = a[17];
  assign n84 = a[19];
  assign n93 = a[21];
  assign n102 = a[23];
  assign n111 = a[25];
  assign n120 = a[27];
  assign n129 = a[29];
  assign n136 = a[31];
  assign n145 = b[0];
  assign n2780 = b[31];
  assign n2781 = b[30];
  assign n2782 = b[29];
  assign n2783 = b[28];
  assign n2784 = b[27];
  assign n2785 = b[26];
  assign n2786 = b[25];
  assign n2787 = b[24];
  assign n2788 = b[23];
  assign n2789 = b[22];
  assign n2790 = b[21];
  assign n2791 = b[20];
  assign n2792 = b[19];
  assign n2793 = b[18];
  assign n2794 = b[17];
  assign n2795 = b[16];
  assign n2796 = b[15];
  assign n2797 = b[14];
  assign n2798 = b[13];
  assign n2799 = b[12];
  assign n2800 = b[11];
  assign n2801 = b[10];
  assign n2802 = b[9];
  assign n2803 = b[8];
  assign n2804 = b[7];
  assign n2805 = b[6];
  assign n2806 = b[5];
  assign n2807 = b[4];
  assign n2808 = b[3];
  assign n2809 = b[2];
  assign n2810 = b[1];

  CND2X2 U187 ( .A(n735), .B(net18422), .Z(n241) );
  COND1X1 U208 ( .A(n3658), .B(n149), .C(n258), .Z(n256) );
  CND2X2 U213 ( .A(n272), .B(n736), .Z(n261) );
  COND1X1 U222 ( .A(n268), .B(n3279), .C(n269), .Z(n267) );
  CND2X2 U229 ( .A(n283), .B(n4282), .Z(n274) );
  COND1X1 U238 ( .A(n281), .B(n3280), .C(n282), .Z(n280) );
  CNR2X2 U243 ( .A(n333), .B(n3716), .Z(n283) );
  CANR1X1 U250 ( .A(n314), .B(n293), .C(n294), .Z(n292) );
  COND1X1 U252 ( .A(n295), .B(n303), .C(n296), .Z(n294) );
  CNR2X2 U255 ( .A(n813), .B(n818), .Z(n295) );
  COND1X1 U258 ( .A(n298), .B(net19409), .C(n299), .Z(n297) );
  CNR2X2 U265 ( .A(n826), .B(n819), .Z(n302) );
  COND1X1 U268 ( .A(n3628), .B(n149), .C(n306), .Z(n304) );
  COND1X1 U284 ( .A(n318), .B(net19409), .C(n319), .Z(n317) );
  CNR2X2 U295 ( .A(n835), .B(n844), .Z(n324) );
  COND1X1 U298 ( .A(n329), .B(n149), .C(n330), .Z(n328) );
  COND1X1 U316 ( .A(n344), .B(net19409), .C(n345), .Z(n343) );
  COND1X1 U328 ( .A(n353), .B(n3279), .C(n3705), .Z(n352) );
  CNR2X2 U339 ( .A(n365), .B(n389), .Z(n363) );
  CNR2X2 U347 ( .A(n867), .B(n878), .Z(n369) );
  CNR2X2 U375 ( .A(n893), .B(n906), .Z(n389) );
  COND1X1 U378 ( .A(n394), .B(net19409), .C(n395), .Z(n393) );
  CNR2X2 U385 ( .A(n409), .B(n3212), .Z(n396) );
  CNR2X2 U389 ( .A(n907), .B(n922), .Z(n402) );
  COND1X1 U392 ( .A(n405), .B(n149), .C(n406), .Z(n404) );
  CND2X2 U400 ( .A(n923), .B(n938), .Z(n410) );
  COND1X1 U402 ( .A(n3135), .B(net19409), .C(n413), .Z(n411) );
  COND1X1 U420 ( .A(n427), .B(n3279), .C(n428), .Z(n426) );
  COND1X1 U432 ( .A(n440), .B(net19409), .C(n3632), .Z(n435) );
  COND1X1 U450 ( .A(n451), .B(n3280), .C(n452), .Z(n450) );
  COND1X1 U462 ( .A(n3134), .B(net19409), .C(n3718), .Z(n459) );
  CNR2X2 U507 ( .A(n1083), .B(n1106), .Z(n491) );
  COND1X1 U725 ( .A(n651), .B(n668), .C(n3696), .Z(n650) );
  CFA1X1 U858 ( .A(n800), .B(n1771), .CI(n1741), .CO(n796), .S(n797) );
  CFA1X1 U859 ( .A(n1772), .B(n804), .CI(n801), .CO(n798), .S(n799) );
  CFA1X1 U861 ( .A(n1803), .B(n805), .CI(n808), .CO(n802), .S(n803) );
  CFA1X1 U862 ( .A(n810), .B(n1773), .CI(n1742), .CO(n804), .S(n805) );
  CFA1X1 U863 ( .A(n816), .B(n814), .CI(n809), .CO(n806), .S(n807) );
  CFA1X1 U864 ( .A(n1743), .B(n811), .CI(n1804), .CO(n808), .S(n809) );
  CFA1X1 U866 ( .A(n817), .B(n815), .CI(n820), .CO(n812), .S(n813) );
  CFA1X1 U867 ( .A(n1744), .B(n822), .CI(n1834), .CO(n814), .S(n815) );
  CFA1X1 U868 ( .A(n824), .B(n1805), .CI(n1774), .CO(n816), .S(n817) );
  CFA1X1 U869 ( .A(n823), .B(n821), .CI(n828), .CO(n818), .S(n819) );
  CFA1X1 U870 ( .A(n825), .B(n830), .CI(n832), .CO(n820), .S(n821) );
  CFA1X1 U873 ( .A(n838), .B(n829), .CI(n836), .CO(n826), .S(n827) );
  CFA1X1 U874 ( .A(n840), .B(n831), .CI(n833), .CO(n828), .S(n829) );
  CFA1X1 U877 ( .A(n839), .B(n837), .CI(n846), .CO(n834), .S(n835) );
  CFA1X1 U878 ( .A(n850), .B(n848), .CI(n841), .CO(n836), .S(n837) );
  CFA1X1 U879 ( .A(n1837), .B(n852), .CI(n843), .CO(n838), .S(n839) );
  CFA1X1 U880 ( .A(n1777), .B(n1865), .CI(n1747), .CO(n840), .S(n841) );
  CFA1X1 U882 ( .A(n849), .B(n847), .CI(n856), .CO(n844), .S(n845) );
  CFA1X1 U883 ( .A(n851), .B(n858), .CI(n853), .CO(n846), .S(n847) );
  CFA1X1 U884 ( .A(n1895), .B(n860), .CI(n862), .CO(n848), .S(n849) );
  CFA1X1 U886 ( .A(n4034), .B(n1866), .CI(n1807), .CO(n852), .S(n853) );
  CFA1X1 U887 ( .A(n859), .B(n868), .CI(n857), .CO(n854), .S(n855) );
  CFA1X1 U888 ( .A(n861), .B(n870), .CI(n872), .CO(n856), .S(n857) );
  CFA1X1 U889 ( .A(n876), .B(n863), .CI(n874), .CO(n858), .S(n859) );
  CFA1X1 U890 ( .A(n1867), .B(n865), .CI(n1779), .CO(n860), .S(n861) );
  CFA1X1 U894 ( .A(n884), .B(n882), .CI(n873), .CO(n868), .S(n869) );
  CFA1X1 U895 ( .A(n886), .B(n877), .CI(n875), .CO(n870), .S(n871) );
  CFA1X1 U896 ( .A(n1780), .B(n888), .CI(n1927), .CO(n872), .S(n873) );
  CFA1X1 U897 ( .A(n1839), .B(n1868), .CI(n1750), .CO(n874), .S(n875) );
  CFA1X1 U899 ( .A(n883), .B(n881), .CI(n894), .CO(n878), .S(n879) );
  CFA1X1 U900 ( .A(n885), .B(n896), .CI(n898), .CO(n880), .S(n881) );
  CFA1X1 U901 ( .A(n900), .B(n889), .CI(n887), .CO(n882), .S(n883) );
  CFA1X1 U902 ( .A(n891), .B(n902), .CI(n904), .CO(n884), .S(n885) );
  CFA1X1 U904 ( .A(n1810), .B(n1928), .CI(n1781), .CO(n888), .S(n889) );
  CFA1X1 U910 ( .A(n920), .B(n1958), .CI(n1899), .CO(n900), .S(n901) );
  CFA1X1 U916 ( .A(n934), .B(n917), .CI(n932), .CO(n912), .S(n913) );
  CFA1X1 U921 ( .A(n927), .B(n925), .CI(n940), .CO(n922), .S(n923) );
  CFA1X1 U922 ( .A(n944), .B(n942), .CI(n929), .CO(n924), .S(n925) );
  CFA1X1 U923 ( .A(n937), .B(n931), .CI(n946), .CO(n926), .S(n927) );
  CFA1X1 U924 ( .A(n948), .B(n935), .CI(n933), .CO(n928), .S(n929) );
  CFA1X1 U925 ( .A(n1990), .B(n950), .CI(n952), .CO(n930), .S(n931) );
  CFA1X1 U926 ( .A(n1841), .B(n1931), .CI(n1901), .CO(n932), .S(n933) );
  CFA1X1 U927 ( .A(n1872), .B(n1813), .CI(n1784), .CO(n934), .S(n935) );
  CFA1X1 U932 ( .A(n951), .B(n949), .CI(n953), .CO(n944), .S(n945) );
  CFA1X1 U934 ( .A(n3712), .B(n955), .CI(n1932), .CO(n948), .S(n949) );
  CFA1X1 U938 ( .A(n961), .B(n959), .CI(n976), .CO(n956), .S(n957) );
  CFA1X1 U939 ( .A(n980), .B(n978), .CI(n963), .CO(n958), .S(n959) );
  CFA1X1 U940 ( .A(n982), .B(n965), .CI(n967), .CO(n960), .S(n961) );
  CFA1X1 U941 ( .A(n971), .B(n984), .CI(n973), .CO(n962), .S(n963) );
  CFA1X1 U943 ( .A(n1962), .B(n990), .CI(n2022), .CO(n966), .S(n967) );
  CFA1X1 U944 ( .A(n1933), .B(n1873), .CI(n1843), .CO(n968), .S(n969) );
  CFA1X1 U948 ( .A(n1000), .B(n998), .CI(n981), .CO(n976), .S(n977) );
  CFA1X1 U950 ( .A(n989), .B(n1004), .CI(n991), .CO(n980), .S(n981) );
  CFA1X1 U952 ( .A(n993), .B(n1010), .CI(n1012), .CO(n984), .S(n985) );
  CFA1X1 U953 ( .A(n1963), .B(n1934), .CI(n1904), .CO(n986), .S(n987) );
  CFA1X1 U954 ( .A(n1816), .B(n1787), .CI(n1993), .CO(n988), .S(n989) );
  CFA1X1 U955 ( .A(n1844), .B(n2023), .CI(n1757), .CO(n990), .S(n991) );
  CFA1X1 U957 ( .A(n999), .B(n997), .CI(n1016), .CO(n994), .S(n995) );
  CFA1X1 U959 ( .A(n1005), .B(n1003), .CI(n1022), .CO(n998), .S(n999) );
  CFA1X1 U960 ( .A(n1007), .B(n1024), .CI(n1026), .CO(n1000), .S(n1001) );
  CFA1X1 U962 ( .A(n1032), .B(n1028), .CI(n1030), .CO(n1004), .S(n1005) );
  CFA1X1 U964 ( .A(n1817), .B(n1874), .CI(n1935), .CO(n1008), .S(n1009) );
  CFA1X1 U965 ( .A(n1845), .B(n1905), .CI(n1788), .CO(n1010), .S(n1011) );
  CFA1X1 U971 ( .A(n1029), .B(n1031), .CI(n1033), .CO(n1022), .S(n1023) );
  CFA1X1 U972 ( .A(n1054), .B(n1052), .CI(n1050), .CO(n1024), .S(n1025) );
  CFA1X1 U973 ( .A(n1965), .B(n1056), .CI(n1035), .CO(n1026), .S(n1027) );
  CFA1X1 U978 ( .A(n1041), .B(n1039), .CI(n1060), .CO(n1036), .S(n1037) );
  CFA1X1 U980 ( .A(n1047), .B(n1045), .CI(n1066), .CO(n1040), .S(n1041) );
  CFA1X1 U984 ( .A(n2088), .B(n1076), .CI(n1078), .CO(n1048), .S(n1049) );
  CFA1X1 U987 ( .A(n1819), .B(n1790), .CI(n1937), .CO(n1054), .S(n1055) );
  CFA1X1 U988 ( .A(n2057), .B(n1080), .CI(n1760), .CO(n1056), .S(n1057) );
  CFA1X1 U990 ( .A(n1088), .B(n1086), .CI(n1065), .CO(n1060), .S(n1061) );
  CFA1X1 U996 ( .A(n1967), .B(n1081), .CI(n1848), .CO(n1072), .S(n1073) );
  CFA1X1 U998 ( .A(n2058), .B(n2027), .CI(n1877), .CO(n1076), .S(n1077) );
  CFA1X1 U999 ( .A(n1907), .B(n1791), .CI(n2089), .CO(n1078), .S(n1079) );
  CFA1X1 U1006 ( .A(n1105), .B(n1103), .CI(n1099), .CO(n1092), .S(n1093) );
  CFA1X1 U1008 ( .A(n2028), .B(n1128), .CI(n2121), .CO(n1096), .S(n1097) );
  CFA1X1 U1010 ( .A(n1878), .B(n1938), .CI(n1849), .CO(n1100), .S(n1101) );
  CFA1X1 U1011 ( .A(n1908), .B(n4023), .CI(n1792), .CO(n1102), .S(n1103) );
  CFA1X1 U1012 ( .A(n1762), .B(n2090), .CI(n2059), .CO(n1104), .S(n1105) );
  CFA1X1 U1016 ( .A(n1144), .B(n1142), .CI(n1119), .CO(n1112), .S(n1113) );
  CFA1X1 U1018 ( .A(n1123), .B(n1127), .CI(n1129), .CO(n1116), .S(n1117) );
  CFA1X1 U1021 ( .A(n2060), .B(n1999), .CI(n2029), .CO(n1122), .S(n1123) );
  CFA1X1 U1022 ( .A(n2091), .B(n4005), .CI(n1850), .CO(n1124), .S(n1125) );
  CFA1X1 U1023 ( .A(n1879), .B(n1822), .CI(n1763), .CO(n1126), .S(n1127) );
  CFA1X1 U1024 ( .A(n1909), .B(n1793), .CI(n2122), .CO(n1128), .S(n1129) );
  CFA1X1 U1031 ( .A(n1155), .B(n1149), .CI(n1157), .CO(n1142), .S(n1143) );
  CFA1X1 U1035 ( .A(n1910), .B(n2000), .CI(n1880), .CO(n1150), .S(n1151) );
  CFA1X1 U1042 ( .A(n1173), .B(n1196), .CI(n1171), .CO(n1164), .S(n1165) );
  CFA1X1 U1043 ( .A(n1175), .B(n1198), .CI(n1200), .CO(n1166), .S(n1167) );
  CFA1X1 U1046 ( .A(n1206), .B(n1204), .CI(n1210), .CO(n1172), .S(n1173) );
  CFA1X1 U1048 ( .A(n2062), .B(n2031), .CI(n2124), .CO(n1176), .S(n1177) );
  CFA1X1 U1049 ( .A(n1852), .B(n2001), .CI(n1881), .CO(n1178), .S(n1179) );
  CFA1X1 U1050 ( .A(n1911), .B(n1824), .CI(n1795), .CO(n1180), .S(n1181) );
  CFA1X1 U1051 ( .A(n1765), .B(n1940), .CI(n2155), .CO(n1182), .S(n1183) );
  CFA1X1 U1056 ( .A(n1201), .B(n1224), .CI(n1199), .CO(n1192), .S(n1193) );
  CFA1X1 U1058 ( .A(n1207), .B(n1230), .CI(n1209), .CO(n1196), .S(n1197) );
  CFA1X1 U1062 ( .A(n1941), .B(n2094), .CI(n2125), .CO(n1204), .S(n1205) );
  CFA1X1 U1064 ( .A(n2002), .B(n1912), .CI(n1882), .CO(n1208), .S(n1209) );
  CFA1X1 U1070 ( .A(n1229), .B(n1227), .CI(n1254), .CO(n1220), .S(n1221) );
  CFA1X1 U1078 ( .A(n1826), .B(n1854), .CI(n2126), .CO(n1236), .S(n1237) );
  CFA1X1 U1086 ( .A(n1288), .B(n1286), .CI(n1261), .CO(n1252), .S(n1253) );
  CFA1X1 U1092 ( .A(n2065), .B(n2127), .CI(n2158), .CO(n1264), .S(n1265) );
  CFA1X1 U1095 ( .A(n2189), .B(n1973), .CI(n1768), .CO(n1270), .S(n1271) );
  COR2X1 U1097 ( .A(n1798), .B(n2034), .Z(n1272) );
  CFA1X1 U1102 ( .A(n1318), .B(n1316), .CI(n1291), .CO(n1282), .S(n1283) );
  CFA1X1 U1105 ( .A(n1322), .B(n1324), .CI(n1326), .CO(n1288), .S(n1289) );
  CFA1X1 U1109 ( .A(n2097), .B(n2128), .CI(n1915), .CO(n1296), .S(n1297) );
  CFA1X1 U1111 ( .A(n1799), .B(n2004), .CI(n2221), .CO(n1300), .S(n1301) );
  CHA1X1 U1112 ( .A(n1769), .B(n1724), .CO(n1302), .S(n1303) );
  CFA1X1 U1119 ( .A(n1331), .B(n1327), .CI(n1329), .CO(n1316), .S(n1317) );
  CFA1X1 U1120 ( .A(n1352), .B(n1354), .CI(n1356), .CO(n1318), .S(n1319) );
  CFA1X1 U1121 ( .A(n2129), .B(n1350), .CI(n4288), .CO(n1320), .S(n1321) );
  CFA1X1 U1122 ( .A(n2160), .B(n2098), .CI(n2067), .CO(n1322), .S(n1323) );
  CFA1X1 U1124 ( .A(n2191), .B(n1886), .CI(n1857), .CO(n1326), .S(n1327) );
  CFA1X1 U1125 ( .A(n2222), .B(n2005), .CI(n1800), .CO(n1328), .S(n1329) );
  CFA1X1 U1126 ( .A(n1770), .B(n2036), .CI(n1829), .CO(n1330), .S(n1331) );
  CFA1X1 U1132 ( .A(n1355), .B(n1357), .CI(n1353), .CO(n1342), .S(n1343) );
  CFA1X1 U1135 ( .A(n2006), .B(n1359), .CI(n4028), .CO(n1348), .S(n1349) );
  CFA1X1 U1137 ( .A(n1830), .B(n1858), .CI(n1887), .CO(n1352), .S(n1353) );
  CFA1X1 U1139 ( .A(n2223), .B(n2037), .CI(n2192), .CO(n1356), .S(n1357) );
  CFA1X1 U1150 ( .A(n2131), .B(n1947), .CI(n1918), .CO(n1378), .S(n1379) );
  CFA1X1 U1151 ( .A(n2162), .B(n1888), .CI(n1831), .CO(n1380), .S(n1381) );
  CFA1X1 U1152 ( .A(n2007), .B(n2193), .CI(n2224), .CO(n1382), .S(n1383) );
  CFA1X1 U1156 ( .A(n1420), .B(n1418), .CI(n1397), .CO(n1390), .S(n1391) );
  CFA1X1 U1164 ( .A(n2194), .B(n2008), .CI(n1889), .CO(n1406), .S(n1407) );
  CFA1X1 U1167 ( .A(n3382), .B(n1415), .CI(n1438), .CO(n1412), .S(n1413) );
  CFA1X1 U1170 ( .A(n1446), .B(n1444), .CI(n1448), .CO(n1418), .S(n1419) );
  CFA1X1 U1174 ( .A(n2133), .B(n1458), .CI(n2102), .CO(n1426), .S(n1427) );
  CFA1X1 U1185 ( .A(n1459), .B(n1478), .CI(n1480), .CO(n1448), .S(n1449) );
  CFA1X1 U1188 ( .A(n1891), .B(n1980), .CI(n1921), .CO(n1454), .S(n1455) );
  CFA1X1 U1189 ( .A(n2072), .B(n2196), .CI(n2227), .CO(n1456), .S(n1457) );
  CFA1X1 U1191 ( .A(n1465), .B(n1463), .CI(n1484), .CO(n1460), .S(n1461) );
  CFA1X1 U1192 ( .A(n1488), .B(n1486), .CI(n1467), .CO(n1462), .S(n1463) );
  CFA1X1 U1196 ( .A(n1498), .B(n1481), .CI(n1496), .CO(n1470), .S(n1471) );
  CFA1X1 U1197 ( .A(n2104), .B(n1500), .CI(n1502), .CO(n1472), .S(n1473) );
  CFA1X1 U1198 ( .A(n2135), .B(n4024), .CI(n1981), .CO(n1474), .S(n1475) );
  CFA1X1 U1199 ( .A(n2197), .B(n1951), .CI(n2166), .CO(n1476), .S(n1477) );
  CFA1X1 U1200 ( .A(n2042), .B(n2228), .CI(n1892), .CO(n1478), .S(n1479) );
  CFA1X1 U1201 ( .A(n1863), .B(n1922), .CI(n2073), .CO(n1480), .S(n1481) );
  CFA1X1 U1205 ( .A(n1501), .B(n1495), .CI(n1514), .CO(n1488), .S(n1489) );
  CFA1X1 U1206 ( .A(n1520), .B(n1499), .CI(n1497), .CO(n1490), .S(n1491) );
  CFA1X1 U1208 ( .A(n2105), .B(n1503), .CI(n2043), .CO(n1494), .S(n1495) );
  CFA1X1 U1209 ( .A(n2136), .B(n3404), .CI(n1952), .CO(n1496), .S(n1497) );
  CFA1X1 U1210 ( .A(n2012), .B(n2167), .CI(n2198), .CO(n1498), .S(n1499) );
  CFA1X1 U1211 ( .A(n2074), .B(n1923), .CI(n2229), .CO(n1500), .S(n1501) );
  CFA1X1 U1218 ( .A(n3711), .B(n1538), .CI(n1540), .CO(n1514), .S(n1515) );
  CFA1X1 U1221 ( .A(n2230), .B(n2044), .CI(n1924), .CO(n1520), .S(n1521) );
  CFA1X1 U1223 ( .A(n3128), .B(n1527), .CI(n1546), .CO(n1524), .S(n1525) );
  CFA1X1 U1224 ( .A(n1533), .B(n1548), .CI(n1531), .CO(n1526), .S(n1527) );
  CFA1X1 U1225 ( .A(n1552), .B(n1550), .CI(n1535), .CO(n1528), .S(n1529) );
  CFA1X1 U1226 ( .A(n1539), .B(n1554), .CI(n1541), .CO(n1530), .S(n1531) );
  CFA1X1 U1227 ( .A(n1558), .B(n1537), .CI(n1556), .CO(n1532), .S(n1533) );
  CFA1X1 U1228 ( .A(n2045), .B(n1560), .CI(n1543), .CO(n1534), .S(n1535) );
  CFA1X1 U1229 ( .A(n2107), .B(n1984), .CI(n1954), .CO(n1536), .S(n1537) );
  CFA1X1 U1230 ( .A(n2169), .B(n2138), .CI(n2014), .CO(n1538), .S(n1539) );
  CFA1X1 U1231 ( .A(n2231), .B(n2200), .CI(n2076), .CO(n1540), .S(n1541) );
  CFA1X1 U1233 ( .A(n1549), .B(n1547), .CI(n1564), .CO(n1544) );
  CFA1X1 U1235 ( .A(n1555), .B(n1568), .CI(n1570), .CO(n1548), .S(n1549) );
  CFA1X1 U1236 ( .A(n1561), .B(n1557), .CI(n1559), .CO(n1550), .S(n1551) );
  CFA1X1 U1237 ( .A(n1576), .B(n1574), .CI(n1572), .CO(n1552), .S(n1553) );
  CFA1X1 U1238 ( .A(n3608), .B(n1578), .CI(n2139), .CO(n1554), .S(n1555) );
  CFA1X1 U1239 ( .A(n2201), .B(n2046), .CI(n2015), .CO(n1556), .S(n1557) );
  CFA1X1 U1240 ( .A(n2077), .B(n2232), .CI(n1955), .CO(n1558), .S(n1559) );
  CFA1X1 U1244 ( .A(n1577), .B(n1586), .CI(n1588), .CO(n1566), .S(n1567) );
  CFA1X1 U1246 ( .A(n1579), .B(n1592), .CI(n1594), .CO(n1570), .S(n1571) );
  CFA1X1 U1248 ( .A(n2078), .B(n2016), .CI(n2202), .CO(n1574), .S(n1575) );
  CFA1X1 U1249 ( .A(n2109), .B(n2233), .CI(n1986), .CO(n1576), .S(n1577) );
  CFA1X1 U1253 ( .A(n1593), .B(n1602), .CI(n1604), .CO(n1584), .S(n1585) );
  CFA1X1 U1254 ( .A(n1606), .B(n1591), .CI(n1595), .CO(n1586), .S(n1587) );
  CFA1X1 U1255 ( .A(n2172), .B(n1608), .CI(n1610), .CO(n1588), .S(n1589) );
  CFA1X1 U1256 ( .A(n2079), .B(n2048), .CI(n2203), .CO(n1590), .S(n1591) );
  CFA1X1 U1257 ( .A(n2234), .B(n2110), .CI(n1987), .CO(n1592), .S(n1593) );
  CFA1X1 U1258 ( .A(n1957), .B(n2017), .CI(n2141), .CO(n1594), .S(n1595) );
  CFA1X1 U1259 ( .A(n1601), .B(n1599), .CI(n1614), .CO(n1596), .S(n1597) );
  CFA1X1 U1262 ( .A(n1620), .B(n1624), .CI(n1622), .CO(n1602), .S(n1603) );
  CFA1X1 U1264 ( .A(n2049), .B(n2080), .CI(n2018), .CO(n1606), .S(n1607) );
  CFA1X1 U1265 ( .A(n2111), .B(n2235), .CI(n2204), .CO(n1608), .S(n1609) );
  CFA1X1 U1267 ( .A(n1617), .B(n1615), .CI(n1628), .CO(n1612), .S(n1613) );
  CFA1X1 U1268 ( .A(n1632), .B(n1630), .CI(n1619), .CO(n1614), .S(n1615) );
  CFA1X1 U1271 ( .A(n2081), .B(n2205), .CI(n2174), .CO(n1620), .S(n1621) );
  CFA1X1 U1272 ( .A(n2112), .B(n2236), .CI(n2019), .CO(n1622), .S(n1623) );
  CFA1X1 U1274 ( .A(n1631), .B(n1629), .CI(n1642), .CO(n1626), .S(n1627) );
  CFA1X1 U1275 ( .A(n1646), .B(n1633), .CI(n1644), .CO(n1628), .S(n1629) );
  CFA1X1 U1276 ( .A(n1648), .B(n1637), .CI(n1635), .CO(n1630), .S(n1631) );
  CFA1X1 U1277 ( .A(n2175), .B(n1639), .CI(n1650), .CO(n1632), .S(n1633) );
  CFA1X1 U1278 ( .A(n2113), .B(n2206), .CI(n2082), .CO(n1634), .S(n1635) );
  CFA1X1 U1281 ( .A(n1645), .B(n1643), .CI(n1654), .CO(n1640), .S(n1641) );
  CFA1X1 U1282 ( .A(n1649), .B(n1656), .CI(n1647), .CO(n1642), .S(n1643) );
  CFA1X1 U1284 ( .A(n2207), .B(n1662), .CI(n2114), .CO(n1646), .S(n1647) );
  CFA1X1 U1285 ( .A(n2145), .B(n2052), .CI(n2238), .CO(n1648), .S(n1649) );
  CFA1X1 U1287 ( .A(n1657), .B(n1655), .CI(n1666), .CO(n1652), .S(n1653) );
  CFA1X1 U1288 ( .A(n1659), .B(n1668), .CI(n1661), .CO(n1654), .S(n1655) );
  CFA1X1 U1289 ( .A(n1663), .B(n1670), .CI(n1672), .CO(n1656), .S(n1657) );
  CFA1X1 U1290 ( .A(n3687), .B(n1733), .CI(n3437), .CO(n1658), .S(n1659) );
  CFA1X1 U1291 ( .A(n2146), .B(n2239), .CI(n2208), .CO(n1660), .S(n1661) );
  CFA1X1 U1293 ( .A(n1676), .B(n1667), .CI(n1669), .CO(n1664), .S(n1665) );
  CFA1X1 U1294 ( .A(n1673), .B(n1678), .CI(n1671), .CO(n1666), .S(n1667) );
  CFA1X1 U1295 ( .A(n2209), .B(n1680), .CI(n1682), .CO(n1668), .S(n1669) );
  CFA1X1 U1296 ( .A(n2147), .B(n2085), .CI(n2240), .CO(n1670), .S(n1671) );
  CFA1X1 U1298 ( .A(n1679), .B(n1677), .CI(n1686), .CO(n1674), .S(n1675) );
  CFA1X1 U1299 ( .A(n1690), .B(n1681), .CI(n1688), .CO(n1676), .S(n1677) );
  CFA1X1 U1300 ( .A(n2148), .B(n1683), .CI(n1734), .CO(n1678), .S(n1679) );
  CFA1X1 U1301 ( .A(n2179), .B(n2241), .CI(n2210), .CO(n1680), .S(n1681) );
  CFA1X1 U1303 ( .A(n1689), .B(n1687), .CI(n1694), .CO(n1684), .S(n1685) );
  CFA1X1 U1304 ( .A(n1698), .B(n1696), .CI(n1691), .CO(n1686), .S(n1687) );
  CFA1X1 U1307 ( .A(n1697), .B(n1695), .CI(n1702), .CO(n1692), .S(n1693) );
  CFA1X1 U1308 ( .A(n2212), .B(n1704), .CI(n1699), .CO(n1694), .S(n1695) );
  CHA1X1 U1310 ( .A(n2150), .B(n2119), .CO(n1698), .S(n1699) );
  CFA1X1 U1311 ( .A(n1708), .B(n1703), .CI(n1705), .CO(n1700), .S(n1701) );
  CFA1X1 U1312 ( .A(n2182), .B(n1710), .CI(n2244), .CO(n1702), .S(n1703) );
  CFA1X1 U1313 ( .A(n2120), .B(n2213), .CI(n2151), .CO(n1704), .S(n1705) );
  CFA1X1 U1314 ( .A(n1711), .B(n1709), .CI(n1714), .CO(n1706), .S(n1707) );
  CFA1X1 U1315 ( .A(n2214), .B(n2245), .CI(n2183), .CO(n1708), .S(n1709) );
  CHA1X1 U1316 ( .A(n1736), .B(n2152), .CO(n1710), .S(n1711) );
  CFA1X1 U1317 ( .A(n2246), .B(n1715), .CI(n1718), .CO(n1712), .S(n1713) );
  CFA1X1 U1318 ( .A(n2215), .B(n2153), .CI(n2184), .CO(n1714), .S(n1715) );
  CFA1X1 U1319 ( .A(n2216), .B(n1719), .CI(n2247), .CO(n1716), .S(n1717) );
  CHA1X1 U1320 ( .A(n1737), .B(n2185), .CO(n1718), .S(n1719) );
  CFA1X1 U1321 ( .A(n2186), .B(n2248), .CI(n2217), .CO(n1720), .S(n1721) );
  CHA1X1 U1322 ( .A(n1738), .B(n2249), .CO(n1722), .S(n1723) );
  COND2X1 U1323 ( .A(n4261), .B(n4263), .C(n3576), .D(n2284), .Z(n1724) );
  COND2X1 U1336 ( .A(n4260), .B(n2264), .C(n3576), .D(n2263), .Z(n1750) );
  COND2X1 U1338 ( .A(n144), .B(n2266), .C(n3576), .D(n2265), .Z(n1752) );
  COND2X1 U1340 ( .A(n4261), .B(n2268), .C(n3577), .D(n2267), .Z(n1754) );
  COND2X1 U1341 ( .A(n144), .B(n2269), .C(n3576), .D(n2268), .Z(n1755) );
  COND2X1 U1343 ( .A(n4260), .B(n2271), .C(n3576), .D(n2270), .Z(n1757) );
  COND2X1 U1344 ( .A(n144), .B(n2272), .C(n3576), .D(n2271), .Z(n1758) );
  COND2X1 U1346 ( .A(n144), .B(n2274), .C(n3577), .D(n2273), .Z(n1760) );
  COND2X1 U1347 ( .A(n4260), .B(n2275), .C(n3577), .D(n2274), .Z(n1761) );
  COND2X1 U1349 ( .A(n4260), .B(n2277), .C(n3577), .D(n2276), .Z(n1763) );
  COND2X1 U1352 ( .A(n4260), .B(n2280), .C(n3577), .D(n2279), .Z(n1766) );
  COND2X1 U1354 ( .A(n144), .B(n2282), .C(n3576), .D(n2281), .Z(n1768) );
  COND2X1 U1355 ( .A(n2283), .B(n4261), .C(n3577), .D(n2282), .Z(n1769) );
  CND2IX1 U1389 ( .B(net16109), .A(n4262), .Z(n2284) );
  COND2X1 U1400 ( .A(n3116), .B(n2294), .C(n3709), .D(n2293), .Z(n1779) );
  COND2X1 U1403 ( .A(n4136), .B(n2297), .C(n3709), .D(n2296), .Z(n1782) );
  COND2X1 U1404 ( .A(n3116), .B(n2298), .C(n3709), .D(n2297), .Z(n1783) );
  COND2X1 U1405 ( .A(n3116), .B(n2299), .C(n3709), .D(n2298), .Z(n1784) );
  COND2X1 U1407 ( .A(n4136), .B(n2301), .C(n3709), .D(n2300), .Z(n1786) );
  COND2X1 U1408 ( .A(n3116), .B(n2302), .C(n3709), .D(n2301), .Z(n1787) );
  COND2X1 U1409 ( .A(n4136), .B(n2303), .C(n132), .D(n2302), .Z(n1788) );
  COND2X1 U1410 ( .A(n4136), .B(n2304), .C(n3709), .D(n2303), .Z(n1789) );
  COND2X1 U1411 ( .A(n3116), .B(n2305), .C(n3709), .D(n2304), .Z(n1790) );
  COND2X1 U1412 ( .A(n3116), .B(n2306), .C(n3709), .D(n2305), .Z(n1791) );
  COND2X1 U1413 ( .A(n3116), .B(n2307), .C(n3709), .D(n2306), .Z(n1792) );
  COND2X1 U1414 ( .A(n3116), .B(n2308), .C(n3709), .D(n2307), .Z(n1793) );
  COND2X1 U1415 ( .A(n135), .B(n2309), .C(n132), .D(n2308), .Z(n1794) );
  COND2X1 U1416 ( .A(n3116), .B(n2310), .C(n132), .D(n2309), .Z(n1795) );
  COND2X1 U1417 ( .A(n135), .B(n2311), .C(n132), .D(n2310), .Z(n1796) );
  COND2X1 U1418 ( .A(n4136), .B(n2312), .C(n132), .D(n2311), .Z(n1797) );
  COND2X1 U1419 ( .A(n135), .B(n2313), .C(n3709), .D(n2312), .Z(n1798) );
  COND2X1 U1420 ( .A(n135), .B(n2314), .C(n132), .D(n2313), .Z(n1799) );
  COND2X1 U1421 ( .A(n135), .B(n2315), .C(n132), .D(n2314), .Z(n1800) );
  COND2X1 U1468 ( .A(n3607), .B(n2328), .C(net16802), .D(n2327), .Z(n1811) );
  COND2X1 U1471 ( .A(n3607), .B(n2331), .C(net16802), .D(n2330), .Z(n1814) );
  COND2X1 U1472 ( .A(n3606), .B(n2332), .C(net16802), .D(n2331), .Z(n1815) );
  COND2X1 U1473 ( .A(n3607), .B(n2333), .C(net16802), .D(n2332), .Z(n1816) );
  COND2X1 U1474 ( .A(n3606), .B(n2334), .C(net16801), .D(n2333), .Z(n1817) );
  COND2X1 U1475 ( .A(n3607), .B(n2335), .C(net16802), .D(n2334), .Z(n1818) );
  COND2X1 U1476 ( .A(n3606), .B(n2336), .C(net16802), .D(n2335), .Z(n1819) );
  COND2X1 U1477 ( .A(n3607), .B(n2337), .C(net16802), .D(n2336), .Z(n1820) );
  COND2X1 U1480 ( .A(n126), .B(n2340), .C(net16802), .D(n2339), .Z(n1823) );
  COND2X1 U1483 ( .A(n3606), .B(n2343), .C(net16802), .D(n2342), .Z(n1826) );
  COND2X1 U1484 ( .A(n3606), .B(n2344), .C(net16801), .D(n2343), .Z(n1827) );
  COND2X1 U1487 ( .A(n126), .B(n2347), .C(net16801), .D(n3575), .Z(n1830) );
  COND2X1 U1488 ( .A(n3606), .B(n2348), .C(net16801), .D(n2347), .Z(n1831) );
  COND2X1 U1531 ( .A(n4033), .B(n2357), .C(net16784), .D(n2356), .Z(n1839) );
  COND2X1 U1532 ( .A(n4033), .B(n2358), .C(net16784), .D(n2357), .Z(n890) );
  COND2X1 U1534 ( .A(net19417), .B(n2360), .C(net16784), .D(n2359), .Z(n920)
         );
  COND2X1 U1535 ( .A(n4033), .B(n2361), .C(net16784), .D(n2360), .Z(n1841) );
  COND2X1 U1536 ( .A(net19417), .B(n2362), .C(net16784), .D(n2361), .Z(n1842)
         );
  COND2X1 U1537 ( .A(n117), .B(n2363), .C(net16784), .D(n2362), .Z(n1843) );
  COND2X1 U1538 ( .A(n4033), .B(n2364), .C(net16784), .D(n2363), .Z(n1844) );
  COND2X1 U1539 ( .A(n4033), .B(n2365), .C(n4295), .D(n2364), .Z(n1845) );
  COND2X1 U1540 ( .A(n4033), .B(n2366), .C(net16784), .D(n2365), .Z(n1846) );
  COND2X1 U1542 ( .A(n4033), .B(n2368), .C(n4295), .D(n2367), .Z(n1848) );
  COND2X1 U1543 ( .A(n117), .B(n2369), .C(net16784), .D(n2368), .Z(n1849) );
  COND2X1 U1544 ( .A(n4033), .B(n2370), .C(n3032), .D(n2369), .Z(n1850) );
  COND2X1 U1545 ( .A(n117), .B(n2371), .C(net16784), .D(n2370), .Z(n1851) );
  COND2X1 U1547 ( .A(net19417), .B(n2373), .C(net16784), .D(n2372), .Z(n1853)
         );
  COND2X1 U1548 ( .A(n4033), .B(n2374), .C(n4295), .D(n2373), .Z(n1854) );
  COND2X1 U1550 ( .A(n4033), .B(n2376), .C(net16784), .D(n2375), .Z(n1856) );
  COND2X1 U1551 ( .A(n2377), .B(n117), .C(net16784), .D(n2376), .Z(n1857) );
  COND2X1 U1552 ( .A(n3364), .B(net19417), .C(net16784), .D(n2377), .Z(n1858)
         );
  COND2X1 U1553 ( .A(n2379), .B(net19417), .C(net16784), .D(n2378), .Z(n1859)
         );
  CND2IX1 U1590 ( .B(net16109), .A(n4291), .Z(n2383) );
  COND2X1 U1598 ( .A(net19122), .B(n2390), .C(net16839), .D(n2389), .Z(n1870)
         );
  COND2X1 U1600 ( .A(n4188), .B(n2392), .C(net16839), .D(n2391), .Z(n1872) );
  COND2X1 U1602 ( .A(n4188), .B(n2394), .C(net19462), .D(n2393), .Z(n1873) );
  COND2X1 U1603 ( .A(net19122), .B(n2395), .C(net16839), .D(n2394), .Z(n992)
         );
  COND2X1 U1604 ( .A(n2396), .B(n4188), .C(net19462), .D(n2395), .Z(n1874) );
  COND2X1 U1608 ( .A(net19122), .B(n2400), .C(net19462), .D(n2399), .Z(n1878)
         );
  COND2X1 U1609 ( .A(n4188), .B(n2401), .C(net16839), .D(n2400), .Z(n1879) );
  COND2X1 U1610 ( .A(net19122), .B(n2402), .C(net19462), .D(n2401), .Z(n1880)
         );
  COND2X1 U1612 ( .A(n4188), .B(n2404), .C(net19462), .D(n2403), .Z(n1882) );
  COND2X1 U1613 ( .A(net19122), .B(n2405), .C(net19462), .D(n2404), .Z(n1883)
         );
  COND2X1 U1614 ( .A(n108), .B(n2406), .C(net19462), .D(n2405), .Z(n1884) );
  COND2X1 U1615 ( .A(net19122), .B(n2407), .C(net19462), .D(n2406), .Z(n1885)
         );
  COND2X1 U1616 ( .A(n4188), .B(n2408), .C(net16839), .D(n2407), .Z(n1886) );
  COND2X1 U1618 ( .A(net19122), .B(n2410), .C(net16839), .D(n2409), .Z(n1888)
         );
  COND2X1 U1619 ( .A(n4188), .B(n2411), .C(net19462), .D(n2410), .Z(n1889) );
  COND2X1 U1621 ( .A(n4188), .B(n2413), .C(net16839), .D(n2412), .Z(n1891) );
  COND2X1 U1622 ( .A(n4188), .B(n2414), .C(net19462), .D(n2413), .Z(n1892) );
  COND2X1 U1623 ( .A(n4188), .B(n2415), .C(net19462), .D(n2414), .Z(n1893) );
  COND2X1 U1658 ( .A(n99), .B(n3948), .C(n3919), .D(n2449), .Z(n1729) );
  COND2X1 U1660 ( .A(n2418), .B(n99), .C(n3920), .D(n2417), .Z(n1896) );
  COND2X1 U1663 ( .A(n99), .B(n2421), .C(n3920), .D(n2420), .Z(n1899) );
  COND2X1 U1664 ( .A(n99), .B(n2422), .C(n3919), .D(n2421), .Z(n1900) );
  COND2X1 U1665 ( .A(n99), .B(n2423), .C(n3919), .D(n2422), .Z(n1901) );
  COND2X1 U1666 ( .A(n99), .B(n2424), .C(n3919), .D(n2423), .Z(n1902) );
  COND2X1 U1667 ( .A(n99), .B(n2425), .C(n3919), .D(n2424), .Z(n1903) );
  COND2X1 U1669 ( .A(n99), .B(n2427), .C(n3920), .D(n2426), .Z(n1905) );
  COND2X1 U1672 ( .A(net18897), .B(n2430), .C(n3919), .D(n2429), .Z(n1907) );
  COND2X1 U1673 ( .A(n99), .B(n2431), .C(n3920), .D(n2430), .Z(n1908) );
  COND2X1 U1675 ( .A(net18897), .B(n2433), .C(n3920), .D(n2432), .Z(n1910) );
  COND2X1 U1676 ( .A(net18897), .B(n2434), .C(n3919), .D(n2433), .Z(n1911) );
  COND2X1 U1677 ( .A(n99), .B(n2435), .C(n3919), .D(n2434), .Z(n1912) );
  COND2X1 U1678 ( .A(net18897), .B(n2436), .C(n3919), .D(n2435), .Z(n1913) );
  COND2X1 U1679 ( .A(n99), .B(n2437), .C(n3919), .D(n2436), .Z(n1914) );
  COND2X1 U1680 ( .A(n99), .B(n2438), .C(n3920), .D(n2437), .Z(n1915) );
  COND2X1 U1681 ( .A(n99), .B(n2439), .C(n3920), .D(n2438), .Z(n1916) );
  COND2X1 U1682 ( .A(net18897), .B(n2440), .C(n3919), .D(n2439), .Z(n1917) );
  COND2X1 U1683 ( .A(n99), .B(n2441), .C(n3919), .D(n2440), .Z(n1918) );
  COND2X1 U1686 ( .A(net18897), .B(n2444), .C(n3919), .D(n2443), .Z(n1921) );
  COND2X1 U1687 ( .A(n99), .B(n2445), .C(n3919), .D(n2444), .Z(n1922) );
  COND2X1 U1688 ( .A(n99), .B(n2446), .C(n3919), .D(n2445), .Z(n1923) );
  COND2X1 U1689 ( .A(n99), .B(n2447), .C(n3920), .D(n2446), .Z(n1924) );
  COND2X1 U1690 ( .A(n2448), .B(net18897), .C(n3920), .D(n2447), .Z(n1925) );
  CAOR1X1 U1726 ( .A(n3277), .B(net18593), .C(n2450), .Z(n1927) );
  COND2X1 U1729 ( .A(net18592), .B(n2453), .C(n3278), .D(n2452), .Z(n1930) );
  COND2X1 U1731 ( .A(net18592), .B(n2455), .C(n3278), .D(n2454), .Z(n1932) );
  COND2X1 U1732 ( .A(n90), .B(n2456), .C(n3278), .D(n2455), .Z(n1933) );
  COND2X1 U1733 ( .A(net18592), .B(n2457), .C(n3278), .D(n2456), .Z(n1934) );
  COND2X1 U1734 ( .A(net18592), .B(n2458), .C(n3277), .D(n2457), .Z(n1935) );
  COND2X1 U1735 ( .A(net18593), .B(n2459), .C(n87), .D(n2458), .Z(n1936) );
  COND2X1 U1736 ( .A(net18593), .B(n2460), .C(n3278), .D(n2459), .Z(n1937) );
  COND2X1 U1737 ( .A(n90), .B(n2461), .C(n87), .D(n2460), .Z(n1080) );
  COND2X1 U1738 ( .A(n2462), .B(net18592), .C(n3277), .D(n2461), .Z(n1938) );
  COND2X1 U1739 ( .A(net18592), .B(n2463), .C(n3277), .D(n2462), .Z(n1130) );
  COND2X1 U1742 ( .A(net18593), .B(n3742), .C(n3277), .D(n2465), .Z(n1941) );
  COND2X1 U1744 ( .A(net18593), .B(n2468), .C(n3278), .D(n2467), .Z(n1943) );
  COND2X1 U1745 ( .A(net18593), .B(n2469), .C(n3278), .D(n2468), .Z(n1944) );
  COND2X1 U1748 ( .A(net18592), .B(n2472), .C(n3278), .D(n2471), .Z(n1947) );
  COND2X1 U1751 ( .A(net18593), .B(n2475), .C(n3277), .D(n2474), .Z(n1950) );
  COND2X1 U1752 ( .A(n2476), .B(net18593), .C(n3277), .D(n2475), .Z(n1951) );
  COND2X1 U1753 ( .A(net18592), .B(n2477), .C(n3277), .D(n2476), .Z(n1952) );
  COND2X1 U1754 ( .A(n2478), .B(net18593), .C(n3277), .D(n2477), .Z(n1953) );
  COND2X1 U1755 ( .A(net18592), .B(n2479), .C(n3278), .D(n2478), .Z(n1954) );
  COND2X1 U1756 ( .A(net18592), .B(n2480), .C(n3278), .D(n2479), .Z(n1955) );
  COND2X1 U1795 ( .A(n2484), .B(net19060), .C(n2485), .D(net18607), .Z(n1960)
         );
  COND2X1 U1802 ( .A(net18607), .B(n2492), .C(net19061), .D(n2491), .Z(n1967)
         );
  COND2X1 U1803 ( .A(n81), .B(n2493), .C(net19060), .D(n2492), .Z(n1968) );
  COND2X1 U1806 ( .A(n81), .B(n2496), .C(n2495), .D(net19060), .Z(n1184) );
  COND2X1 U1808 ( .A(net18607), .B(n2498), .C(net19060), .D(n2497), .Z(n1972)
         );
  COND2X1 U1809 ( .A(n4174), .B(net18607), .C(net19061), .D(n2498), .Z(n1973)
         );
  COND2X1 U1811 ( .A(net18607), .B(n2501), .C(net19060), .D(n4189), .Z(n1975)
         );
  COND2X1 U1819 ( .A(net18607), .B(n2509), .C(net19061), .D(n2508), .Z(n1983)
         );
  COND2X1 U1822 ( .A(n81), .B(n2512), .C(n78), .D(n2511), .Z(n1986) );
  COND2X1 U1823 ( .A(net18607), .B(n2513), .C(net19060), .D(n2512), .Z(n1987)
         );
  COND2X1 U1863 ( .A(net19518), .B(n2519), .C(net16771), .D(n2518), .Z(n1993)
         );
  COND2X1 U1866 ( .A(net19518), .B(n2522), .C(n4289), .D(n2521), .Z(n1996) );
  COND2X1 U1869 ( .A(net19518), .B(n2525), .C(n4289), .D(n2524), .Z(n1999) );
  COND2X1 U1870 ( .A(net19518), .B(n2526), .C(n4289), .D(n2525), .Z(n2000) );
  COND2X1 U1871 ( .A(net18670), .B(n2527), .C(net16771), .D(n2526), .Z(n2001)
         );
  COND2X1 U1872 ( .A(net19518), .B(n2528), .C(net16771), .D(n2527), .Z(n2002)
         );
  COND2X1 U1873 ( .A(n3075), .B(n2529), .C(n2528), .D(n4289), .Z(n1242) );
  COND2X1 U1875 ( .A(net19518), .B(n2531), .C(n4144), .D(n2530), .Z(n2004) );
  COND2X1 U1876 ( .A(n3415), .B(n2532), .C(net16771), .D(n2531), .Z(n2005) );
  COND2X1 U1878 ( .A(n3415), .B(n2534), .C(n4289), .D(n2533), .Z(n2007) );
  COND2X1 U1879 ( .A(net19518), .B(n2535), .C(net16771), .D(n2534), .Z(n2008)
         );
  COND2X1 U1881 ( .A(net19518), .B(n2537), .C(net16771), .D(n3876), .Z(n2010)
         );
  COND2X1 U1883 ( .A(net19518), .B(n2539), .C(n4289), .D(n2538), .Z(n2012) );
  COND2X1 U1885 ( .A(net18670), .B(n2541), .C(n4144), .D(n2540), .Z(n2014) );
  COND2X1 U1886 ( .A(n3757), .B(n2542), .C(n4289), .D(n2541), .Z(n2015) );
  COND2X1 U1888 ( .A(net18670), .B(n2544), .C(net16771), .D(n2543), .Z(n2017)
         );
  COND2X1 U1889 ( .A(net19518), .B(n2545), .C(net16771), .D(n2544), .Z(n2018)
         );
  COND2X1 U1890 ( .A(net18670), .B(n2546), .C(net16771), .D(n2545), .Z(n2019)
         );
  COND2X1 U1928 ( .A(n2550), .B(net19168), .C(net19151), .D(n2549), .Z(n2023)
         );
  COND2X1 U1929 ( .A(n2550), .B(net19151), .C(n4135), .D(n2551), .Z(n2024) );
  COND2X1 U1931 ( .A(n63), .B(n2553), .C(net19151), .D(n2552), .Z(n2026) );
  COND2X1 U1932 ( .A(net19168), .B(n2554), .C(net19151), .D(n2553), .Z(n2027)
         );
  COND2X1 U1934 ( .A(n2556), .B(n4135), .C(net19500), .D(n2555), .Z(n2029) );
  COND2X1 U1935 ( .A(net19168), .B(n4030), .C(net19500), .D(n2556), .Z(n2030)
         );
  COND2X1 U1936 ( .A(n2558), .B(n63), .C(net19151), .D(n4030), .Z(n2031) );
  COND2X1 U1937 ( .A(n2559), .B(net19168), .C(net19500), .D(n2558), .Z(n2032)
         );
  COND2X1 U1938 ( .A(n2560), .B(n3139), .C(net19500), .D(n2559), .Z(n2033) );
  COND2X1 U1939 ( .A(n2561), .B(n3139), .C(net19151), .D(n2560), .Z(n2034) );
  COND2X1 U1941 ( .A(n2563), .B(n63), .C(net19500), .D(n2562), .Z(n2036) );
  COND2X1 U1942 ( .A(net19168), .B(n2564), .C(net19151), .D(n2563), .Z(n2037)
         );
  COND2X1 U1943 ( .A(n2565), .B(n3139), .C(net19500), .D(n2564), .Z(n2038) );
  COND2X1 U1944 ( .A(n3139), .B(n2566), .C(net19151), .D(n2565), .Z(n2039) );
  COND2X1 U1947 ( .A(n3139), .B(n2569), .C(net19151), .D(n3873), .Z(n2042) );
  COND2X1 U1948 ( .A(n3139), .B(n2570), .C(net19151), .D(n2569), .Z(n2043) );
  COND2X1 U1949 ( .A(n3139), .B(n2571), .C(net19500), .D(n2570), .Z(n2044) );
  COND2X1 U1951 ( .A(net19168), .B(n2573), .C(net19151), .D(n2572), .Z(n2046)
         );
  COND2X1 U1953 ( .A(n2575), .B(n4135), .C(net19500), .D(n2574), .Z(n2048) );
  COND2X1 U1954 ( .A(n2576), .B(n3139), .C(net19151), .D(n2575), .Z(n2049) );
  COND2X1 U1955 ( .A(net19168), .B(n2577), .C(net19151), .D(n2576), .Z(n2050)
         );
  COND2X1 U1996 ( .A(n2583), .B(n3839), .C(n2584), .D(n54), .Z(n2057) );
  COND2X1 U1997 ( .A(n3877), .B(n2585), .C(n3839), .D(n2584), .Z(n2058) );
  COND2X1 U1998 ( .A(n3877), .B(n2586), .C(n3839), .D(n2585), .Z(n2059) );
  COND2X1 U1999 ( .A(n3877), .B(n2587), .C(net18736), .D(n2586), .Z(n2060) );
  COND2X1 U2001 ( .A(n54), .B(n2589), .C(n3839), .D(n2588), .Z(n2062) );
  COND2X1 U2002 ( .A(n3877), .B(n2590), .C(n3839), .D(n2589), .Z(n2063) );
  COND2X1 U2003 ( .A(n3877), .B(n2591), .C(n3839), .D(n2590), .Z(n2064) );
  COND2X1 U2005 ( .A(n54), .B(n2593), .C(n3839), .D(n2592), .Z(n2066) );
  COND2X1 U2006 ( .A(n3877), .B(n2594), .C(n3839), .D(n2593), .Z(n2067) );
  COND2X1 U2009 ( .A(n3877), .B(n2597), .C(n3839), .D(n2596), .Z(n2070) );
  COND2X1 U2011 ( .A(n54), .B(n2599), .C(net18736), .D(n2598), .Z(n2072) );
  COND2X1 U2012 ( .A(n3877), .B(n2600), .C(n3839), .D(n2599), .Z(n2073) );
  COND2X1 U2013 ( .A(n54), .B(n2601), .C(net18736), .D(n2600), .Z(n2074) );
  COND2X1 U2016 ( .A(n3877), .B(n2604), .C(n3839), .D(n2603), .Z(n2077) );
  COND2X1 U2017 ( .A(n3877), .B(n3443), .C(n3839), .D(n2604), .Z(n2078) );
  COND2X1 U2018 ( .A(n54), .B(n2606), .C(n3839), .D(n2605), .Z(n2079) );
  COND2X1 U2020 ( .A(n54), .B(n2608), .C(n3839), .D(n2607), .Z(n2081) );
  COND2X1 U2021 ( .A(n54), .B(n2609), .C(n3839), .D(n2608), .Z(n2082) );
  COND2X1 U2022 ( .A(n3877), .B(n2610), .C(n3839), .D(n2609), .Z(n2083) );
  COND2X1 U2025 ( .A(n2613), .B(n3877), .C(n3839), .D(n2612), .Z(n2086) );
  COND2X1 U2062 ( .A(n2616), .B(n45), .C(net16793), .D(n2615), .Z(n2089) );
  COND2X1 U2067 ( .A(n3092), .B(n2621), .C(net16793), .D(n2620), .Z(n2094) );
  COND2X1 U2068 ( .A(n45), .B(n2622), .C(n4017), .D(n2621), .Z(n2095) );
  COND2X1 U2070 ( .A(n45), .B(n2624), .C(net16793), .D(n2623), .Z(n2097) );
  COND2X1 U2072 ( .A(n45), .B(n2626), .C(n4018), .D(n2625), .Z(n2099) );
  COND2X1 U2076 ( .A(n45), .B(n2630), .C(n4018), .D(n2629), .Z(n2103) );
  COND2X1 U2079 ( .A(n45), .B(n2633), .C(net16793), .D(n2632), .Z(n2106) );
  COND2X1 U2080 ( .A(n3092), .B(n2634), .C(net16793), .D(n2633), .Z(n2107) );
  COND2X1 U2081 ( .A(n45), .B(n2635), .C(net16793), .D(n2634), .Z(n2108) );
  COND2X1 U2084 ( .A(n3092), .B(n2638), .C(net16793), .D(n2637), .Z(n2111) );
  COND2X1 U2086 ( .A(n3963), .B(n2640), .C(net16793), .D(n2639), .Z(n2113) );
  COND2X1 U2129 ( .A(n2649), .B(n36), .C(net16791), .D(n2648), .Z(n2122) );
  COND2X1 U2132 ( .A(n4002), .B(n2652), .C(net19508), .D(n2651), .Z(n2125) );
  COND2X1 U2133 ( .A(n4003), .B(n2653), .C(net19508), .D(n2652), .Z(n2126) );
  COND2X1 U2135 ( .A(n4002), .B(n2655), .C(net19508), .D(n2654), .Z(n2128) );
  COND2X1 U2138 ( .A(n4003), .B(n2658), .C(net19508), .D(n2657), .Z(n2131) );
  COND2X1 U2140 ( .A(n4003), .B(n2660), .C(net19508), .D(n2659), .Z(n2133) );
  COND2X1 U2141 ( .A(n4002), .B(n2661), .C(net19508), .D(n2660), .Z(n2134) );
  COND2X1 U2142 ( .A(n4003), .B(n2662), .C(net19508), .D(n2661), .Z(n2135) );
  COND2X1 U2143 ( .A(n4002), .B(n2663), .C(net19508), .D(n2662), .Z(n2136) );
  COND2X1 U2144 ( .A(n4003), .B(n2664), .C(net19508), .D(n2663), .Z(n2137) );
  COND2X1 U2145 ( .A(n4003), .B(n2665), .C(net19508), .D(n2664), .Z(n2138) );
  COND2X1 U2146 ( .A(n4002), .B(n2666), .C(net19508), .D(n2665), .Z(n2139) );
  COND2X1 U2147 ( .A(n4003), .B(n2667), .C(net19508), .D(n2666), .Z(n2140) );
  COND2X1 U2150 ( .A(n4002), .B(n2670), .C(net19508), .D(n2669), .Z(n2143) );
  COND2X1 U2153 ( .A(n4002), .B(n2673), .C(net19508), .D(n2672), .Z(n2146) );
  COND2X1 U2154 ( .A(n4003), .B(n2674), .C(net19508), .D(n2673), .Z(n2147) );
  COND2X1 U2156 ( .A(n4003), .B(n2676), .C(net19508), .D(n2675), .Z(n2149) );
  COND2X1 U2159 ( .A(n2679), .B(n4002), .C(net19508), .D(n2678), .Z(n2152) );
  COND2X1 U2196 ( .A(n4040), .B(net18743), .C(n3678), .D(n2681), .Z(n2155) );
  COND2X1 U2198 ( .A(n27), .B(n2684), .C(n3678), .D(n2683), .Z(n2157) );
  COND2X1 U2199 ( .A(n3593), .B(n2685), .C(net16772), .D(n2684), .Z(n2158) );
  COND2X1 U2200 ( .A(net18743), .B(n2686), .C(net16772), .D(n4141), .Z(n2159)
         );
  COND2X1 U2201 ( .A(net18742), .B(n2687), .C(net16772), .D(n2686), .Z(n2160)
         );
  COND2X1 U2202 ( .A(n3024), .B(n2688), .C(net16772), .D(n2687), .Z(n2161) );
  COND2X1 U2203 ( .A(net18742), .B(n2689), .C(net16772), .D(n2688), .Z(n2162)
         );
  COND2X1 U2207 ( .A(n3024), .B(n2693), .C(net16772), .D(n2692), .Z(n2166) );
  COND2X1 U2209 ( .A(n3024), .B(n2695), .C(net16772), .D(n2694), .Z(n2168) );
  COND2X1 U2210 ( .A(net18742), .B(n2696), .C(net16772), .D(n2695), .Z(n2169)
         );
  COND2X1 U2212 ( .A(n3024), .B(n2698), .C(net16772), .D(n2697), .Z(n2171) );
  COND2X1 U2215 ( .A(net18742), .B(n2701), .C(n3678), .D(n2700), .Z(n2174) );
  COND2X1 U2219 ( .A(net18743), .B(n2705), .C(net16772), .D(n2704), .Z(n2178)
         );
  COND2X1 U2225 ( .A(n3024), .B(n2711), .C(net16772), .D(n2710), .Z(n2184) );
  COND2X1 U2263 ( .A(n4221), .B(n18), .C(net16816), .D(n2714), .Z(n2188) );
  COND2X1 U2265 ( .A(n4001), .B(n2717), .C(net16816), .D(n2716), .Z(n2190) );
  COND2X1 U2266 ( .A(n18), .B(n2718), .C(net16817), .D(n2717), .Z(n2191) );
  COND2X1 U2267 ( .A(n4001), .B(n2719), .C(net16817), .D(n2718), .Z(n2192) );
  COND2X1 U2268 ( .A(n18), .B(n2720), .C(net16817), .D(n2719), .Z(n2193) );
  COND2X1 U2269 ( .A(n4001), .B(n2721), .C(net16816), .D(n2720), .Z(n2194) );
  COND2X1 U2271 ( .A(n4001), .B(n2723), .C(net16816), .D(n2722), .Z(n2196) );
  COND2X1 U2272 ( .A(n4001), .B(n2724), .C(net16816), .D(n2723), .Z(n2197) );
  COND2X1 U2273 ( .A(n4001), .B(n2725), .C(net16816), .D(n2724), .Z(n2198) );
  COND2X1 U2274 ( .A(n18), .B(n2726), .C(net16817), .D(n2725), .Z(n2199) );
  COND2X1 U2275 ( .A(n18), .B(n2727), .C(net16816), .D(n2726), .Z(n2200) );
  COND2X1 U2276 ( .A(n4001), .B(n2728), .C(net16816), .D(n2727), .Z(n2201) );
  COND2X1 U2277 ( .A(n4001), .B(n2729), .C(net16816), .D(n2728), .Z(n2202) );
  COND2X1 U2278 ( .A(n18), .B(n2730), .C(net16816), .D(n2729), .Z(n2203) );
  COND2X1 U2279 ( .A(n4001), .B(n2731), .C(net16817), .D(n2730), .Z(n2204) );
  COND2X1 U2280 ( .A(n18), .B(n2732), .C(net16816), .D(n2731), .Z(n2205) );
  COND2X1 U2281 ( .A(n18), .B(n2733), .C(net16816), .D(n2732), .Z(n2206) );
  COND2X1 U2282 ( .A(n4001), .B(n2734), .C(net16816), .D(n2733), .Z(n2207) );
  COND2X1 U2283 ( .A(n4001), .B(n2735), .C(net16817), .D(n2734), .Z(n2208) );
  COND2X1 U2285 ( .A(n4001), .B(n2737), .C(net16816), .D(n2736), .Z(n2210) );
  COND2X1 U2292 ( .A(n4001), .B(n2744), .C(net16816), .D(n2743), .Z(n2217) );
  COND2X1 U2330 ( .A(n2748), .B(net19555), .C(n6), .D(n2747), .Z(n2221) );
  COND2X1 U2332 ( .A(net19555), .B(n2750), .C(n6), .D(n2749), .Z(n2223) );
  COND2X1 U2333 ( .A(net19555), .B(n2751), .C(n6), .D(n2750), .Z(n2224) );
  COND2X1 U2334 ( .A(net19555), .B(n2752), .C(n6), .D(n2751), .Z(n2225) );
  COND2X1 U2336 ( .A(n9), .B(n2754), .C(n6), .D(n2753), .Z(n2227) );
  COND2X1 U2337 ( .A(net19555), .B(n2755), .C(n6), .D(n2754), .Z(n2228) );
  COND2X1 U2338 ( .A(net19555), .B(n2756), .C(n6), .D(n2755), .Z(n2229) );
  COND2X1 U2339 ( .A(n9), .B(n2757), .C(n6), .D(n2756), .Z(n2230) );
  COND2X1 U2340 ( .A(n9), .B(n2758), .C(n6), .D(n2757), .Z(n2231) );
  COND2X1 U2341 ( .A(net19555), .B(n2759), .C(n6), .D(n2758), .Z(n2232) );
  COND2X1 U2342 ( .A(net19555), .B(n2760), .C(n6), .D(n2759), .Z(n2233) );
  COND2X1 U2343 ( .A(net19555), .B(n2761), .C(n6), .D(n2760), .Z(n2234) );
  COND2X1 U2344 ( .A(net19555), .B(n2762), .C(n6), .D(n2761), .Z(n2235) );
  COND2X1 U2346 ( .A(n9), .B(n2764), .C(n6), .D(n2763), .Z(n2237) );
  COND2X1 U2347 ( .A(net19555), .B(n2765), .C(n6), .D(n2764), .Z(n2238) );
  COND2X1 U2348 ( .A(net19555), .B(n2766), .C(n6), .D(n2765), .Z(n2239) );
  COND2X1 U2349 ( .A(net19555), .B(n2767), .C(n6), .D(n2766), .Z(n2240) );
  COND2X1 U2350 ( .A(net19555), .B(n2768), .C(n6), .D(n2767), .Z(n2241) );
  COND2X1 U2351 ( .A(net19555), .B(n2769), .C(n6), .D(n2768), .Z(n2242) );
  COND2X1 U2352 ( .A(net19555), .B(n2770), .C(n6), .D(n2769), .Z(n2243) );
  COND2X1 U2353 ( .A(net19555), .B(n2771), .C(n6), .D(n2770), .Z(n2244) );
  COND2X1 U2354 ( .A(net19555), .B(n2772), .C(n6), .D(n2771), .Z(n2245) );
  COND2X1 U2355 ( .A(net19555), .B(n2773), .C(n6), .D(n2772), .Z(n2246) );
  COND2X1 U2356 ( .A(net19555), .B(n2774), .C(n6), .D(n2773), .Z(n2247) );
  COND2X1 U2357 ( .A(net19555), .B(n2775), .C(n6), .D(n2774), .Z(n2248) );
  COND2X1 U2358 ( .A(net19555), .B(n2776), .C(n6), .D(n2775), .Z(n2249) );
  COND2X1 U2359 ( .A(net19555), .B(n2777), .C(n6), .D(n2776), .Z(n2250) );
  COND2X1 U2360 ( .A(n2778), .B(net19555), .C(n6), .D(n2777), .Z(n2251) );
  CEOX2 U2473 ( .A(n4351), .B(a[20]), .Z(n2817) );
  COND2X1 U1814 ( .A(net18607), .B(n2504), .C(n78), .D(n2503), .Z(n1978) );
  COND2X1 U1816 ( .A(net18607), .B(n2506), .C(net19061), .D(n2505), .Z(n1980)
         );
  COND2X1 U2205 ( .A(net18742), .B(n2691), .C(n3678), .D(n2690), .Z(n2164) );
  COND2X1 U1880 ( .A(net18670), .B(n2536), .C(net16771), .D(n2535), .Z(n2009)
         );
  COND2X1 U1805 ( .A(n81), .B(n2495), .C(net19060), .D(n2494), .Z(n1970) );
  COND2X1 U1815 ( .A(n81), .B(n2505), .C(net19060), .D(n2504), .Z(n1979) );
  CFA1X1 U1175 ( .A(n2009), .B(n1979), .CI(n2164), .CO(n1428), .S(n1429) );
  CNR2X2 U487 ( .A(n514), .B(n480), .Z(n478) );
  COND1X1 U162 ( .A(n220), .B(n3280), .C(n221), .Z(n219) );
  CFA1X1 U1134 ( .A(n1384), .B(n1380), .CI(n1382), .CO(n1346), .S(n1347) );
  CFA1X1 U1153 ( .A(n1802), .B(n1859), .CI(n2069), .CO(n1384), .S(n1385) );
  CFA1X1 U1131 ( .A(n1374), .B(n1372), .CI(n1349), .CO(n1340), .S(n1341) );
  CFA1X1 U1147 ( .A(n1406), .B(n1385), .CI(n1408), .CO(n1372), .S(n1373) );
  CFA1X1 U1144 ( .A(n1396), .B(n1373), .CI(n1375), .CO(n1366), .S(n1367) );
  CNR2X2 U596 ( .A(net19127), .B(n1332), .Z(n556) );
  COND2X1 U1946 ( .A(n3873), .B(n63), .C(net19500), .D(n2567), .Z(n2041) );
  COND2X1 U1945 ( .A(n3139), .B(n3617), .C(net19151), .D(n2566), .Z(n2040) );
  COND2X1 U2335 ( .A(net19555), .B(n2753), .C(n6), .D(n2752), .Z(n2226) );
  COND2X1 U1555 ( .A(n4033), .B(n3878), .C(net16784), .D(n2380), .Z(n1861) );
  CFA1X1 U1177 ( .A(n1861), .B(n2040), .CI(n2226), .CO(n1432), .S(n1433) );
  COND2X1 U2270 ( .A(n18), .B(n2722), .C(net16816), .D(n2721), .Z(n2195) );
  COND2X1 U1750 ( .A(net18593), .B(n2474), .C(n3277), .D(n2473), .Z(n1949) );
  CFA1X1 U1176 ( .A(n2195), .B(n1949), .CI(n1920), .CO(n1430), .S(n1431) );
  CFA1X1 U1160 ( .A(n1430), .B(n1432), .CI(n1428), .CO(n1398), .S(n1399) );
  CFA1X1 U1186 ( .A(n2103), .B(n2134), .CI(n2041), .CO(n1450), .S(n1451) );
  CFA1X1 U1173 ( .A(n1456), .B(n1452), .CI(n1450), .CO(n1424), .S(n1425) );
  COND2X1 U2204 ( .A(net18743), .B(n2690), .C(net16772), .D(n2689), .Z(n2163)
         );
  COND2X1 U1684 ( .A(n99), .B(n2442), .C(n3920), .D(n2441), .Z(n1919) );
  CFA1X1 U1158 ( .A(n1407), .B(n1424), .CI(n1405), .CO(n1394), .S(n1395) );
  CFA1X1 U1141 ( .A(n1365), .B(n1363), .CI(n1388), .CO(n1360), .S(n1361) );
  CFA1X1 U1127 ( .A(n1337), .B(n1335), .CI(n1362), .CO(n1332), .S(n1333) );
  CFA1X1 U1113 ( .A(n1309), .B(n1307), .CI(n1334), .CO(n1304), .S(n1305) );
  COND2X1 U1620 ( .A(net19122), .B(n2412), .C(net16839), .D(n2411), .Z(n1890)
         );
  CFA1X1 U1178 ( .A(n2071), .B(n1890), .CI(n1833), .CO(n1434), .S(n1435) );
  COND2X1 U1489 ( .A(n2349), .B(n3607), .C(net16801), .D(n2348), .Z(n1832) );
  CFA1X1 U1157 ( .A(n1401), .B(n1399), .CI(n1422), .CO(n1392), .S(n1393) );
  CFA1X1 U1161 ( .A(n2101), .B(n1434), .CI(n1411), .CO(n1400), .S(n1401) );
  CFA1X1 U1145 ( .A(n1379), .B(n1398), .CI(n1400), .CO(n1368), .S(n1369) );
  CND2X2 U333 ( .A(n438), .B(n3240), .Z(n353) );
  CANR1X1 U188 ( .A(net18422), .B(n253), .C(n244), .Z(n242) );
  CNR2X2 U181 ( .A(n274), .B(n3710), .Z(n233) );
  COND1X1 U176 ( .A(n231), .B(n3280), .C(n232), .Z(n230) );
  CNIVX1 U2507 ( .A(n1997), .Z(n3022) );
  CIVXL U2508 ( .A(net18608), .Z(n3023) );
  COND2X1 U2509 ( .A(net18593), .B(n2454), .C(n87), .D(n2453), .Z(n1931) );
  CND2X2 U2510 ( .A(n2825), .B(n24), .Z(n3024) );
  CNR2XL U2511 ( .A(n636), .B(n3102), .Z(n3025) );
  CENX1 U2512 ( .A(n1101), .B(n1120), .Z(n4015) );
  CNIVXL U2513 ( .A(net19518), .Z(n3026) );
  CND3X1 U2514 ( .A(n3769), .B(n3770), .C(n3771), .Z(n1280) );
  CND2XL U2515 ( .A(n1280), .B(n1255), .Z(n3631) );
  CND2X1 U2516 ( .A(n3749), .B(n3750), .Z(n3027) );
  CEOXL U2517 ( .A(n4324), .B(n3290), .Z(n2343) );
  CENX1 U2518 ( .A(n4328), .B(net16850), .Z(n2469) );
  CIVX3 U2519 ( .A(n3763), .Z(n3764) );
  CENXL U2520 ( .A(n1894), .B(n2106), .Z(n3463) );
  COND2XL U2521 ( .A(n99), .B(n3948), .C(n3919), .D(n2449), .Z(n3028) );
  CANR1XL U2522 ( .A(net18420), .B(n3613), .C(n216), .Z(n214) );
  CIVXL U2523 ( .A(n659), .Z(n3029) );
  CIVXL U2524 ( .A(n3029), .Z(n3030) );
  COND2XL U2525 ( .A(n144), .B(n2270), .C(n3576), .D(n2269), .Z(n3031) );
  CNIVX1 U2526 ( .A(net16784), .Z(n3032) );
  CIVXL U2527 ( .A(a[18]), .Z(n3488) );
  CENX2 U2528 ( .A(n1020), .B(n1001), .Z(n3113) );
  CNIVXL U2529 ( .A(n1468), .Z(n3033) );
  CND3X1 U2530 ( .A(n4112), .B(n4113), .C(n4114), .Z(n1468) );
  CENX1 U2531 ( .A(n4338), .B(n4343), .Z(n2751) );
  CENX1 U2532 ( .A(n4338), .B(net16843), .Z(n2685) );
  CIVXL U2533 ( .A(n409), .Z(n748) );
  CND2XL U2534 ( .A(n1275), .B(n1304), .Z(n3034) );
  CIVX1 U2535 ( .A(n521), .Z(n3534) );
  COND2X1 U2536 ( .A(net18592), .B(n2473), .C(n3278), .D(n2472), .Z(n1948) );
  CENX1 U2537 ( .A(n4326), .B(net16850), .Z(n2473) );
  CIVXL U2538 ( .A(n1341), .Z(n3422) );
  CIVX1 U2539 ( .A(n2567), .Z(n3616) );
  COND2X2 U2540 ( .A(net18607), .B(n2497), .C(net19060), .D(n2496), .Z(n1971)
         );
  CND3X2 U2541 ( .A(n3243), .B(n3244), .C(n3245), .Z(n904) );
  CND2X1 U2542 ( .A(n1752), .B(n1929), .Z(n3243) );
  CIVXL U2543 ( .A(n1248), .Z(n3035) );
  CIVX1 U2544 ( .A(n3035), .Z(n3036) );
  CND3X1 U2545 ( .A(n3629), .B(n3630), .C(n3631), .Z(n1248) );
  CND2XL U2546 ( .A(n1280), .B(n1282), .Z(n3629) );
  CNIVX1 U2547 ( .A(n1611), .Z(n3037) );
  CDLY1XL U2548 ( .A(n1159), .Z(n3661) );
  CENX2 U2549 ( .A(n3113), .B(n1018), .Z(n997) );
  CIVDX3 U2550 ( .A(n4293), .Z0(n3577) );
  CANR1XL U2551 ( .A(n3824), .B(n535), .C(n521), .Z(n3038) );
  CENX1 U2552 ( .A(n4327), .B(n4349), .Z(n2569) );
  CENX1 U2553 ( .A(n4340), .B(n4343), .Z(n2749) );
  CANR1XL U2554 ( .A(n4277), .B(n3030), .C(n654), .Z(n3039) );
  CANR1X1 U2555 ( .A(n4277), .B(n659), .C(n654), .Z(n3696) );
  CND2X2 U2556 ( .A(n3440), .B(n3441), .Z(n3040) );
  CND2X1 U2557 ( .A(n3440), .B(n3441), .Z(n1275) );
  CND2XL U2558 ( .A(n968), .B(n972), .Z(n3740) );
  CIVX1 U2559 ( .A(n968), .Z(n3571) );
  CNR2X1 U2560 ( .A(net18742), .B(n2703), .Z(n3924) );
  CENX1 U2561 ( .A(n4337), .B(net16844), .Z(n2686) );
  CENX1 U2562 ( .A(n4329), .B(net15995), .Z(n2336) );
  CENX1 U2563 ( .A(n3041), .B(n869), .Z(n867) );
  CENX2 U2564 ( .A(n871), .B(n880), .Z(n3041) );
  CND2XL U2565 ( .A(n987), .B(n1006), .Z(n4070) );
  CND3XL U2566 ( .A(n3697), .B(n3699), .C(n3698), .Z(n3042) );
  CND2X1 U2567 ( .A(net19076), .B(a[10]), .Z(n3541) );
  CENXL U2568 ( .A(n3363), .B(n1136), .Z(n3043) );
  COND2X1 U2569 ( .A(n4260), .B(n2278), .C(n3576), .D(n2277), .Z(n3044) );
  CENXL U2570 ( .A(n3363), .B(n1136), .Z(n1109) );
  COND2XL U2571 ( .A(n4260), .B(n2278), .C(n3576), .D(n2277), .Z(n1764) );
  CND2XL U2572 ( .A(n1551), .B(n1553), .Z(n3101) );
  CFA1X2 U2573 ( .A(n919), .B(n915), .CI(n930), .CO(n910), .S(n911) );
  CEO3X1 U2574 ( .A(n1600), .B(n1589), .C(n1587), .Z(n1583) );
  CND2XL U2575 ( .A(n1600), .B(n1587), .Z(n3045) );
  CND2XL U2576 ( .A(n1600), .B(n1589), .Z(n3046) );
  CND2X1 U2577 ( .A(n1587), .B(n1589), .Z(n3047) );
  CND3X2 U2578 ( .A(n3045), .B(n3046), .C(n3047), .Z(n1582) );
  CND3XL U2579 ( .A(n3688), .B(n3689), .C(n3690), .Z(n3048) );
  CND3X1 U2580 ( .A(n3692), .B(n3693), .C(n3694), .Z(n1600) );
  CND2X1 U2581 ( .A(n1565), .B(n1582), .Z(n3668) );
  CENX1 U2582 ( .A(n4329), .B(net16850), .Z(n2468) );
  CIVX2 U2583 ( .A(n641), .Z(n639) );
  CIVX3 U2584 ( .A(n96), .Z(n3988) );
  CNIVX1 U2585 ( .A(net18670), .Z(n3757) );
  CFA1X1 U2586 ( .A(n1660), .B(n1651), .CI(n1658), .CO(n1644), .S(n1645) );
  CDLY1XL U2587 ( .A(n665), .Z(n3049) );
  CND2X1 U2588 ( .A(n988), .B(n969), .Z(n3301) );
  CENXL U2589 ( .A(n4324), .B(n4000), .Z(n2574) );
  CND2X1 U2590 ( .A(n1121), .B(n1125), .Z(n3394) );
  CENX2 U2591 ( .A(n3050), .B(n1238), .Z(n1203) );
  CENX2 U2592 ( .A(n2187), .B(n1240), .Z(n3050) );
  CIVX2 U2593 ( .A(n1339), .Z(n3423) );
  CND2X2 U2594 ( .A(n1091), .B(n1093), .Z(n4185) );
  CIVX3 U2595 ( .A(a[6]), .Z(n3662) );
  CENX2 U2596 ( .A(n3051), .B(n2130), .Z(n1355) );
  CENX1 U2597 ( .A(n2161), .B(n1946), .Z(n3051) );
  CND2X1 U2598 ( .A(n3368), .B(n3053), .Z(n3054) );
  CND2X1 U2599 ( .A(n3052), .B(n3372), .Z(n3055) );
  CND2X2 U2600 ( .A(n3054), .B(n3055), .Z(n1033) );
  CIVX2 U2601 ( .A(n3368), .Z(n3052) );
  CIVXL U2602 ( .A(n3372), .Z(n3053) );
  CIVXL U2603 ( .A(n3356), .Z(n3056) );
  CIVX2 U2604 ( .A(n1875), .Z(n3356) );
  CENX2 U2605 ( .A(n3057), .B(n1429), .Z(n1423) );
  CENX2 U2606 ( .A(n1454), .B(n1435), .Z(n3057) );
  CND2XL U2607 ( .A(n1566), .B(n1551), .Z(n3099) );
  CND3X2 U2608 ( .A(n3184), .B(n3185), .C(n3186), .Z(n916) );
  CIVX1 U2609 ( .A(n1492), .Z(n3680) );
  CIVXL U2610 ( .A(n4356), .Z(n3058) );
  CENX1 U2611 ( .A(n1220), .B(n1193), .Z(n3639) );
  COND2XL U2612 ( .A(n3607), .B(n2327), .C(net16801), .D(n2326), .Z(n1810) );
  CND2X4 U2613 ( .A(n2813), .B(n132), .Z(n135) );
  CIVXL U2614 ( .A(net19316), .Z(n3059) );
  CIVXL U2615 ( .A(n3059), .Z(n3060) );
  CEOX2 U2616 ( .A(n1267), .B(n1290), .Z(n3952) );
  COR2XL U2617 ( .A(n1613), .B(n1626), .Z(n3061) );
  CENX2 U2618 ( .A(n1569), .B(n4006), .Z(n1565) );
  COND2XL U2619 ( .A(n99), .B(n2429), .C(n3920), .D(n2428), .Z(n1906) );
  CHA1X1 U2620 ( .A(n1726), .B(n1832), .CO(n1410), .S(n1411) );
  COND2X1 U2621 ( .A(n126), .B(n3984), .C(net16802), .D(n2350), .Z(n1726) );
  CENX1 U2622 ( .A(n2810), .B(n3393), .Z(n2414) );
  CND2XL U2623 ( .A(n2130), .B(n1946), .Z(n3062) );
  CND2XL U2624 ( .A(n2130), .B(n2161), .Z(n3063) );
  CND2XL U2625 ( .A(n1946), .B(n2161), .Z(n3064) );
  CND3X1 U2626 ( .A(n3062), .B(n3063), .C(n3064), .Z(n1354) );
  COR2X1 U2627 ( .A(n4002), .B(n2657), .Z(n3065) );
  COR2XL U2628 ( .A(net19508), .B(n2656), .Z(n3066) );
  CND2X2 U2629 ( .A(n3065), .B(n3066), .Z(n2130) );
  CENXL U2630 ( .A(n2789), .B(n4255), .Z(n2657) );
  CENXL U2631 ( .A(net16544), .B(n4254), .Z(n2656) );
  CEO3X2 U2632 ( .A(n1337), .B(n1335), .C(n1362), .Z(n3892) );
  CIVXL U2633 ( .A(n4088), .Z(n3067) );
  CIVXL U2634 ( .A(n3067), .Z(n3068) );
  COND2X1 U2635 ( .A(net19122), .B(n2399), .C(net19462), .D(n2398), .Z(n1877)
         );
  CND2X2 U2636 ( .A(n1223), .B(n1225), .Z(n3849) );
  CANR1XL U2637 ( .A(n419), .B(n387), .C(n388), .Z(n3069) );
  COND1X1 U2638 ( .A(n389), .B(n4011), .C(n392), .Z(n388) );
  CND2XL U2639 ( .A(n102), .B(a[22]), .Z(n3072) );
  CND2X1 U2640 ( .A(n3070), .B(n3071), .Z(n3073) );
  CND2X1 U2641 ( .A(n3072), .B(n3073), .Z(n4187) );
  CIVXL U2642 ( .A(a[22]), .Z(n3070) );
  CIVXL U2643 ( .A(n102), .Z(n3071) );
  CND2X1 U2644 ( .A(n1218), .B(n1220), .Z(n3960) );
  CENX2 U2645 ( .A(n1092), .B(n3218), .Z(n1065) );
  CIVX1 U2646 ( .A(n572), .Z(n766) );
  CENX2 U2647 ( .A(n1234), .B(n1232), .Z(n3448) );
  CIVX2 U2648 ( .A(n4025), .Z(n3968) );
  CND2X1 U2649 ( .A(n1394), .B(n1371), .Z(n3194) );
  CENX1 U2650 ( .A(n4325), .B(net18643), .Z(n2540) );
  COND2X2 U2651 ( .A(n54), .B(n2603), .C(n3839), .D(n2602), .Z(n2076) );
  CND2XL U2652 ( .A(n1404), .B(n1410), .Z(n3205) );
  CND2XL U2653 ( .A(n1338), .B(n1340), .Z(n4215) );
  CAN2XL U2654 ( .A(n1769), .B(n1724), .Z(n3074) );
  CENX2 U2655 ( .A(n4323), .B(net16788), .Z(n2608) );
  CIVXL U2656 ( .A(n3414), .Z(n3075) );
  CIVX1 U2657 ( .A(n3414), .Z(n3415) );
  CENX1 U2658 ( .A(n4331), .B(n4253), .Z(n2400) );
  CIVX4 U2659 ( .A(net16089), .Z(net16083) );
  CIVX1 U2660 ( .A(n3397), .Z(n3398) );
  CEO3X2 U2661 ( .A(n1976), .B(n1917), .C(n2099), .Z(n1351) );
  CND2XL U2662 ( .A(n1976), .B(n2099), .Z(n3076) );
  CND2XL U2663 ( .A(n1976), .B(n1917), .Z(n3077) );
  CND2XL U2664 ( .A(n2099), .B(n1917), .Z(n3078) );
  CND3X1 U2665 ( .A(n3076), .B(n3077), .C(n3078), .Z(n1350) );
  CEO3X2 U2666 ( .A(n1297), .B(n1295), .C(n1320), .Z(n1285) );
  CND2X1 U2667 ( .A(n1297), .B(n1320), .Z(n3079) );
  CND2XL U2668 ( .A(n1297), .B(n1295), .Z(n3080) );
  CND2X2 U2669 ( .A(n1320), .B(n1295), .Z(n3081) );
  CND3X2 U2670 ( .A(n3079), .B(n3080), .C(n3081), .Z(n1284) );
  COND2X1 U2671 ( .A(n2502), .B(net18607), .C(n78), .D(n2501), .Z(n1976) );
  CEO3X2 U2672 ( .A(n2066), .B(n1828), .C(n1856), .Z(n1295) );
  CIVXL U2673 ( .A(n1638), .Z(n3082) );
  CIVXL U2674 ( .A(n3082), .Z(n3083) );
  CIVX2 U2675 ( .A(n3768), .Z(n3207) );
  CENXL U2676 ( .A(n4339), .B(n4254), .Z(n2651) );
  CND2XL U2677 ( .A(n1943), .B(n1827), .Z(n4300) );
  CND3X2 U2678 ( .A(n4183), .B(n4184), .C(n4185), .Z(n1086) );
  CND2X1 U2679 ( .A(n1114), .B(n1091), .Z(n4183) );
  CND2X1 U2680 ( .A(n1114), .B(n1093), .Z(n4184) );
  CEO3X1 U2681 ( .A(n1378), .B(n1351), .C(n1376), .Z(n1345) );
  CND2XL U2682 ( .A(n1378), .B(n1351), .Z(n3084) );
  CND2XL U2683 ( .A(n1378), .B(n1376), .Z(n3085) );
  CND2X1 U2684 ( .A(n1351), .B(n1376), .Z(n3086) );
  CND3X2 U2685 ( .A(n3084), .B(n3085), .C(n3086), .Z(n1344) );
  CEOX2 U2686 ( .A(n1346), .B(n1321), .Z(n3087) );
  CEOX2 U2687 ( .A(n3087), .B(n1344), .Z(n1313) );
  CND2XL U2688 ( .A(n1346), .B(n1321), .Z(n3088) );
  CND2X1 U2689 ( .A(n1346), .B(n1344), .Z(n3089) );
  CND2X1 U2690 ( .A(n1321), .B(n1344), .Z(n3090) );
  CND3X1 U2691 ( .A(n3088), .B(n3089), .C(n3090), .Z(n1312) );
  CND2X1 U2692 ( .A(n1995), .B(n1936), .Z(n3506) );
  CIVX1 U2693 ( .A(n416), .Z(n418) );
  CEO3X2 U2694 ( .A(n1201), .B(n1224), .C(n1199), .Z(n3091) );
  CND3X2 U2695 ( .A(n3321), .B(n3322), .C(n3323), .Z(n1224) );
  CND2X2 U2696 ( .A(n2823), .B(n42), .Z(n3092) );
  CND2X1 U2697 ( .A(n2823), .B(n42), .Z(n3963) );
  COND1X1 U2698 ( .A(n666), .B(n660), .C(n661), .Z(n659) );
  CENX2 U2699 ( .A(n3093), .B(n3122), .Z(n1447) );
  CENX1 U2700 ( .A(n1476), .B(n1474), .Z(n3093) );
  CIVX3 U2701 ( .A(n39), .Z(net18817) );
  COR2X1 U2702 ( .A(n36), .B(n2671), .Z(n3094) );
  COR2X1 U2703 ( .A(n4175), .B(n2670), .Z(n3095) );
  CND2X2 U2704 ( .A(n3094), .B(n3095), .Z(n2144) );
  CNIVX1 U2705 ( .A(n33), .Z(n4175) );
  CAN2XL U2706 ( .A(n3028), .B(n1925), .Z(n3711) );
  CND2XL U2707 ( .A(n1203), .B(n1228), .Z(n4245) );
  CNIVXL U2708 ( .A(n3220), .Z(n3403) );
  CIVXL U2709 ( .A(n1280), .Z(n3096) );
  CIVX1 U2710 ( .A(n3096), .Z(n3097) );
  CND2X4 U2711 ( .A(n2822), .B(net18953), .Z(n54) );
  CENX1 U2712 ( .A(n4332), .B(net16063), .Z(n2596) );
  CEOX2 U2713 ( .A(n1553), .B(n1551), .Z(n3098) );
  CEOX2 U2714 ( .A(n3098), .B(n1566), .Z(n1547) );
  CND2X1 U2715 ( .A(n1566), .B(n1553), .Z(n3100) );
  CND3X2 U2716 ( .A(n3099), .B(n3100), .C(n3101), .Z(n1546) );
  CNR2XL U2717 ( .A(n1545), .B(n1562), .Z(n3102) );
  CNR2XL U2718 ( .A(n1545), .B(n1562), .Z(n3103) );
  CEO3X1 U2719 ( .A(n1529), .B(n1546), .C(n1527), .Z(n4089) );
  CNR2X1 U2720 ( .A(n1545), .B(n1562), .Z(n633) );
  CIVXL U2721 ( .A(n632), .Z(n3104) );
  CIVXL U2722 ( .A(n3104), .Z(n3105) );
  CND2X2 U2723 ( .A(n3635), .B(n3636), .Z(n1163) );
  CND2X2 U2724 ( .A(n3633), .B(n3527), .Z(n3636) );
  CENX2 U2725 ( .A(net16558), .B(net16850), .Z(n2465) );
  CENX2 U2726 ( .A(n1203), .B(n1228), .Z(n4234) );
  CENX2 U2727 ( .A(n1147), .B(n1168), .Z(n3449) );
  CND3XL U2728 ( .A(n3913), .B(n3914), .C(n3915), .Z(n3106) );
  CND3XL U2729 ( .A(n3913), .B(n3914), .C(n3915), .Z(n3107) );
  CND3XL U2730 ( .A(n3913), .B(n3914), .C(n3915), .Z(n1162) );
  CND2X2 U2731 ( .A(n4172), .B(n33), .Z(n36) );
  CNIVX2 U2732 ( .A(n30), .Z(n3574) );
  CIVXL U2733 ( .A(n3788), .Z(n3108) );
  CIVX1 U2734 ( .A(n612), .Z(n611) );
  CFA1XL U2735 ( .A(n2180), .B(n2242), .CI(n2118), .CO(n1688), .S(n1689) );
  CENXL U2736 ( .A(n673), .B(n198), .Z(product[14]) );
  CHA1X1 U2737 ( .A(n2084), .B(n2053), .CO(n1662), .S(n1663) );
  COND1XL U2738 ( .A(n585), .B(n611), .C(n586), .Z(n584) );
  CENXL U2739 ( .A(n190), .B(n3109), .Z(product[22]) );
  CAOR1X1 U2740 ( .A(n773), .B(n629), .C(n626), .Z(n3109) );
  CND3X1 U2741 ( .A(n3305), .B(n3306), .C(n3307), .Z(n942) );
  CND2IX2 U2742 ( .B(n3110), .A(n3249), .Z(n1929) );
  CNR2XL U2743 ( .A(n2451), .B(n3277), .Z(n3110) );
  COND2X1 U2744 ( .A(n4188), .B(n2387), .C(net19462), .D(n2386), .Z(n1867) );
  CENX1 U2745 ( .A(n4334), .B(n4251), .Z(n2297) );
  CANR1X1 U2746 ( .A(n4282), .B(n286), .C(n277), .Z(n3111) );
  CANR1XL U2747 ( .A(n4282), .B(n286), .C(n277), .Z(n3112) );
  CANR1X1 U2748 ( .A(n4282), .B(n286), .C(n277), .Z(n275) );
  CENXL U2749 ( .A(n181), .B(n3114), .Z(product[31]) );
  CAOR1X1 U2750 ( .A(n554), .B(n574), .C(n555), .Z(n3114) );
  COR2X1 U2751 ( .A(n974), .B(n957), .Z(n4276) );
  CENX1 U2752 ( .A(n1013), .B(n3182), .Z(n1003) );
  CND2X1 U2753 ( .A(n658), .B(n4277), .Z(n651) );
  CND2X2 U2754 ( .A(n3508), .B(n3509), .Z(n1995) );
  CANR1X1 U2755 ( .A(n397), .B(n363), .C(n364), .Z(n3797) );
  CEN3X2 U2756 ( .A(n1213), .B(n1211), .C(n3410), .Z(n1199) );
  CENX1 U2757 ( .A(n3115), .B(n2176), .Z(n1651) );
  CENX1 U2758 ( .A(n2021), .B(n2083), .Z(n3115) );
  CIVXL U2759 ( .A(n410), .Z(n408) );
  CND2XL U2760 ( .A(n1473), .B(n1494), .Z(n3813) );
  CND2X4 U2761 ( .A(n3890), .B(n132), .Z(n3116) );
  CND2X2 U2762 ( .A(n3890), .B(n132), .Z(n4136) );
  CIVXL U2763 ( .A(n582), .Z(n3117) );
  CND2XL U2764 ( .A(n1008), .B(n987), .Z(n4068) );
  CND2X1 U2765 ( .A(n3912), .B(n3634), .Z(n3635) );
  CNIVX16 U2766 ( .A(n4351), .Z(n4292) );
  CND2X1 U2767 ( .A(n1253), .B(n1278), .Z(n4181) );
  COND1X1 U2768 ( .A(n675), .B(n671), .C(n672), .Z(n670) );
  CIVXL U2769 ( .A(n671), .Z(n780) );
  CENX1 U2770 ( .A(n1177), .B(n3118), .Z(n1171) );
  CENX1 U2771 ( .A(n1208), .B(n1179), .Z(n3118) );
  CAOR1X1 U2772 ( .A(net16772), .B(net18743), .C(n2681), .Z(n2154) );
  CND2XL U2773 ( .A(n1148), .B(n1152), .Z(n3436) );
  CND2XL U2774 ( .A(n1150), .B(n1148), .Z(n3434) );
  CEO3XL U2775 ( .A(n1631), .B(n1642), .C(n1629), .Z(n3119) );
  CND3XL U2776 ( .A(n3701), .B(n3702), .C(n3703), .Z(n3120) );
  CND3XL U2777 ( .A(n3701), .B(n3702), .C(n3703), .Z(n3121) );
  CND3XL U2778 ( .A(n3701), .B(n3702), .C(n3703), .Z(n1464) );
  CNIVX2 U2779 ( .A(n1451), .Z(n3122) );
  CENX1 U2780 ( .A(n3123), .B(n3121), .Z(n1439) );
  CENX1 U2781 ( .A(n1443), .B(n1466), .Z(n3123) );
  CENX2 U2782 ( .A(a[20]), .B(n3987), .Z(n3124) );
  CENX2 U2783 ( .A(a[20]), .B(n3987), .Z(n96) );
  CIVX4 U2784 ( .A(n3988), .Z(net16812) );
  CENX1 U2785 ( .A(n3125), .B(n1469), .Z(n1465) );
  CENX1 U2786 ( .A(n1471), .B(n1490), .Z(n3125) );
  CEOX4 U2787 ( .A(a[16]), .B(n3997), .Z(n3126) );
  CENX1 U2788 ( .A(n4322), .B(net18643), .Z(n2543) );
  CNIVX3 U2789 ( .A(net19401), .Z(net16824) );
  CNIVXL U2790 ( .A(n983), .Z(n3127) );
  CNIVX1 U2791 ( .A(n1529), .Z(n3128) );
  CIVXL U2792 ( .A(n1584), .Z(n3695) );
  COND1X2 U2793 ( .A(n559), .B(net18620), .C(n552), .Z(n3174) );
  CNR2X2 U2794 ( .A(n3892), .B(n1360), .Z(n3544) );
  COR2X1 U2795 ( .A(n939), .B(n956), .Z(n3129) );
  CND2X2 U2796 ( .A(n1245), .B(n1274), .Z(n4088) );
  CAN2X1 U2797 ( .A(n3856), .B(n3857), .Z(n3130) );
  CND2XL U2798 ( .A(n1215), .B(n1244), .Z(n3131) );
  CND2X1 U2799 ( .A(net19521), .B(n1436), .Z(net19292) );
  CEO3XL U2800 ( .A(n1114), .B(n1093), .C(n1091), .Z(n3132) );
  COAN1XL U2801 ( .A(n385), .B(n4020), .C(n3069), .Z(n3133) );
  CIVX2 U2802 ( .A(n472), .Z(n3602) );
  CNIVXL U2803 ( .A(n460), .Z(n3134) );
  COR2XL U2804 ( .A(n440), .B(n416), .Z(n3135) );
  COR2XL U2805 ( .A(n1059), .B(n3405), .Z(n3136) );
  COR2X1 U2806 ( .A(n1483), .B(n1504), .Z(n3620) );
  CND2X2 U2807 ( .A(n620), .B(n3621), .Z(n3442) );
  CNR2X2 U2808 ( .A(n627), .B(n622), .Z(n620) );
  CIVXL U2809 ( .A(net19200), .Z(n629) );
  CENX2 U2810 ( .A(a[16]), .B(net18937), .Z(n78) );
  CENX1 U2811 ( .A(n4333), .B(n4306), .Z(n2562) );
  CIVXL U2812 ( .A(n3178), .Z(n3137) );
  CIVX1 U2813 ( .A(n1853), .Z(n3178) );
  CEOX1 U2814 ( .A(n1383), .B(n1381), .Z(n4226) );
  CENX2 U2815 ( .A(n4323), .B(n4292), .Z(n2443) );
  CEOXL U2816 ( .A(n4107), .B(n3361), .Z(n3138) );
  CIVX2 U2817 ( .A(n3360), .Z(n3361) );
  CND2X2 U2818 ( .A(n4012), .B(net19500), .Z(n3139) );
  CENX1 U2819 ( .A(n4329), .B(n4145), .Z(n2567) );
  COND1X2 U2820 ( .A(n410), .B(n402), .C(n403), .Z(n397) );
  CENX1 U2821 ( .A(n3140), .B(n1235), .Z(n1229) );
  CENX1 U2822 ( .A(n1270), .B(n1268), .Z(n3140) );
  CND2XL U2823 ( .A(n1139), .B(n1164), .Z(n4039) );
  CENX2 U2824 ( .A(n3141), .B(n1121), .Z(n1115) );
  CENX2 U2825 ( .A(n1146), .B(n1125), .Z(n3141) );
  CND2X1 U2826 ( .A(n1442), .B(n3744), .Z(n3745) );
  CND2X2 U2827 ( .A(n1605), .B(n3143), .Z(n3144) );
  CND2X1 U2828 ( .A(n3142), .B(n1603), .Z(n3145) );
  CND2X2 U2829 ( .A(n3144), .B(n3145), .Z(n3648) );
  CIVX2 U2830 ( .A(n1605), .Z(n3142) );
  CIVX1 U2831 ( .A(n1603), .Z(n3143) );
  CENX1 U2832 ( .A(n4327), .B(net18982), .Z(n2701) );
  CENXL U2833 ( .A(n4338), .B(n4306), .Z(n2553) );
  CIVX4 U2834 ( .A(n3126), .Z(net19061) );
  CEOX2 U2835 ( .A(n962), .B(n945), .Z(n3146) );
  CEOX2 U2836 ( .A(n3146), .B(n960), .Z(n941) );
  CND2X1 U2837 ( .A(n960), .B(n945), .Z(n3147) );
  CND2X1 U2838 ( .A(n960), .B(n962), .Z(n3148) );
  CND2XL U2839 ( .A(n945), .B(n962), .Z(n3149) );
  CND3X2 U2840 ( .A(n3147), .B(n3148), .C(n3149), .Z(n940) );
  CND2X1 U2841 ( .A(n1121), .B(n1146), .Z(n3395) );
  CND2XL U2842 ( .A(n2024), .B(n1034), .Z(n3295) );
  COND2XL U2843 ( .A(net18607), .B(n2494), .C(net19061), .D(n2493), .Z(n1969)
         );
  COND2XL U2844 ( .A(net18670), .B(n3733), .C(n4289), .D(n2522), .Z(n1997) );
  CND3X1 U2845 ( .A(n4163), .B(n4164), .C(n4165), .Z(n1158) );
  COND2XL U2846 ( .A(n3963), .B(n2625), .C(net16793), .D(n2624), .Z(n2098) );
  CND2X1 U2847 ( .A(net16027), .B(n3488), .Z(n3489) );
  CANR1XL U2848 ( .A(net18739), .B(n562), .C(n3174), .Z(n3150) );
  CANR1X1 U2849 ( .A(net18739), .B(n562), .C(n3174), .Z(n548) );
  CIVX4 U2850 ( .A(n4361), .Z(n3151) );
  CIVX1 U2851 ( .A(n4361), .Z(n3152) );
  CEOX2 U2852 ( .A(n1048), .B(n1046), .Z(n3153) );
  CEOX1 U2853 ( .A(n3153), .B(n1027), .Z(n1021) );
  CND2XL U2854 ( .A(n1027), .B(n1046), .Z(n3154) );
  CND2X1 U2855 ( .A(n1027), .B(n1048), .Z(n3155) );
  CND2XL U2856 ( .A(n1046), .B(n1048), .Z(n3156) );
  CND3X1 U2857 ( .A(n3154), .B(n3155), .C(n3156), .Z(n1020) );
  CEO3X2 U2858 ( .A(n1021), .B(n1042), .C(n1040), .Z(n1017) );
  CND2XL U2859 ( .A(n1021), .B(n1040), .Z(n3157) );
  CND2XL U2860 ( .A(n1021), .B(n1042), .Z(n3158) );
  CND2X1 U2861 ( .A(n1040), .B(n1042), .Z(n3159) );
  CND3X1 U2862 ( .A(n3157), .B(n3158), .C(n3159), .Z(n1016) );
  CIVX2 U2863 ( .A(n4361), .Z(n4359) );
  CND2X1 U2864 ( .A(n1020), .B(n1018), .Z(n3254) );
  CND2X2 U2865 ( .A(n1115), .B(n1140), .Z(n3784) );
  CND3X2 U2866 ( .A(n3939), .B(n3940), .C(n3941), .Z(n1228) );
  CND2X1 U2867 ( .A(n1130), .B(n1154), .Z(n3162) );
  CND2X2 U2868 ( .A(n3160), .B(n3161), .Z(n3163) );
  CND2X2 U2869 ( .A(n3162), .B(n3163), .Z(n4058) );
  CIVXL U2870 ( .A(n1130), .Z(n3160) );
  CIVX2 U2871 ( .A(n1154), .Z(n3161) );
  CFA1X1 U2872 ( .A(n1794), .B(n1939), .CI(n1823), .CO(n1154), .S(n1155) );
  CNR2X2 U2873 ( .A(n1187), .B(n1214), .Z(n529) );
  CND2X1 U2874 ( .A(n1299), .B(n1301), .Z(n3166) );
  CND2X2 U2875 ( .A(n3164), .B(n3165), .Z(n3167) );
  CND2X2 U2876 ( .A(n3166), .B(n3167), .Z(n3514) );
  CIVX2 U2877 ( .A(n1299), .Z(n3164) );
  CIVX2 U2878 ( .A(n1301), .Z(n3165) );
  CENX2 U2879 ( .A(n3449), .B(n1145), .Z(n1139) );
  CENX1 U2880 ( .A(n3168), .B(n1053), .Z(n1045) );
  CENX2 U2881 ( .A(n1055), .B(n1057), .Z(n3168) );
  CEOX2 U2882 ( .A(n916), .B(n903), .Z(n3169) );
  CEOX2 U2883 ( .A(n3169), .B(n918), .Z(n899) );
  CND2XL U2884 ( .A(n918), .B(n903), .Z(n3170) );
  CND2X1 U2885 ( .A(n918), .B(n916), .Z(n3171) );
  CND2XL U2886 ( .A(n903), .B(n916), .Z(n3172) );
  CND3X1 U2887 ( .A(n3170), .B(n3171), .C(n3172), .Z(n898) );
  CFA1X1 U2888 ( .A(n1122), .B(n1126), .CI(n1124), .CO(n1094), .S(n1095) );
  CNIVX2 U2889 ( .A(n1969), .Z(n4005) );
  COND2XL U2890 ( .A(n4003), .B(n2675), .C(net19508), .D(n2674), .Z(n2148) );
  COND2XL U2891 ( .A(n4003), .B(n2677), .C(net19508), .D(n2676), .Z(n2150) );
  COND2X1 U2892 ( .A(n4003), .B(n2659), .C(net16791), .D(n2658), .Z(n2132) );
  CIVXL U2893 ( .A(n4356), .Z(n3173) );
  CENX2 U2894 ( .A(n1135), .B(n4272), .Z(n1133) );
  CEO3X2 U2895 ( .A(n1116), .B(n1097), .C(n1095), .Z(n1089) );
  CENX2 U2896 ( .A(n1112), .B(n1089), .Z(n3614) );
  CND2XL U2897 ( .A(n1767), .B(n1942), .Z(n4168) );
  CIVXL U2898 ( .A(n432), .Z(n3175) );
  CND2XL U2899 ( .A(n1170), .B(n1172), .Z(n3780) );
  CEO3X1 U2900 ( .A(n1475), .B(n1477), .C(n1479), .Z(n1469) );
  CND3X2 U2901 ( .A(n3369), .B(n3370), .C(n3371), .Z(n1032) );
  CND2X1 U2902 ( .A(n3372), .B(n3056), .Z(n3370) );
  COND2XL U2903 ( .A(n4260), .B(n2273), .C(n3577), .D(n2272), .Z(n1759) );
  COND2X1 U2904 ( .A(n3877), .B(n2588), .C(n3839), .D(n2587), .Z(n2061) );
  CENX2 U2905 ( .A(n3409), .B(n3640), .Z(n3176) );
  CENXL U2906 ( .A(n3409), .B(n3640), .Z(n1161) );
  CND2X1 U2907 ( .A(n1796), .B(n3178), .Z(n3179) );
  CND2X1 U2908 ( .A(n3177), .B(n1853), .Z(n3180) );
  CND2X2 U2909 ( .A(n3179), .B(n3180), .Z(n3221) );
  CIVXL U2910 ( .A(n1796), .Z(n3177) );
  CENXL U2911 ( .A(n4323), .B(n4360), .Z(n2311) );
  CENXL U2912 ( .A(n2802), .B(net16850), .Z(n2472) );
  CENXL U2913 ( .A(n2810), .B(net16850), .Z(n2480) );
  CENXL U2914 ( .A(n4323), .B(net16850), .Z(n2476) );
  CENXL U2915 ( .A(n4321), .B(net16850), .Z(n2479) );
  CENXL U2916 ( .A(n4331), .B(net16850), .Z(n2466) );
  CENX1 U2917 ( .A(n4330), .B(net16850), .Z(n2467) );
  CENX1 U2918 ( .A(n4332), .B(net16850), .Z(n2464) );
  COND2X2 U2919 ( .A(n117), .B(n2372), .C(net16784), .D(n2371), .Z(n1852) );
  CENX2 U2920 ( .A(n3181), .B(n1256), .Z(n1223) );
  CENX2 U2921 ( .A(n1258), .B(n1231), .Z(n3181) );
  CND3X2 U2922 ( .A(n4296), .B(n4297), .C(n4298), .Z(n1132) );
  CENX2 U2923 ( .A(n1009), .B(n1011), .Z(n3182) );
  CEOX2 U2924 ( .A(n1930), .B(n1783), .Z(n3183) );
  CEOX2 U2925 ( .A(n3183), .B(n3234), .Z(n917) );
  CND2XL U2926 ( .A(n3234), .B(n1783), .Z(n3184) );
  CND2X1 U2927 ( .A(n3234), .B(n1930), .Z(n3185) );
  CND2XL U2928 ( .A(n1783), .B(n1930), .Z(n3186) );
  CIVX2 U2929 ( .A(n3233), .Z(n3234) );
  CND3X1 U2930 ( .A(n3965), .B(n3966), .C(n3967), .Z(n1058) );
  CENX1 U2931 ( .A(n4336), .B(n4253), .Z(n2390) );
  CENX2 U2932 ( .A(n3187), .B(n1062), .Z(n1039) );
  CENX2 U2933 ( .A(n1064), .B(n1043), .Z(n3187) );
  CIVX1 U2934 ( .A(n4358), .Z(n3263) );
  CANR1X2 U2935 ( .A(net18739), .B(n562), .C(n3174), .Z(n3946) );
  CND3X2 U2936 ( .A(n3387), .B(n3388), .C(n3389), .Z(n1238) );
  CIVX1 U2937 ( .A(n3124), .Z(n3377) );
  CEO3X2 U2938 ( .A(n2064), .B(n1243), .C(n2033), .Z(n1233) );
  CND2XL U2939 ( .A(n1243), .B(n2033), .Z(n3188) );
  CND2XL U2940 ( .A(n1243), .B(n2064), .Z(n3189) );
  CND2X1 U2941 ( .A(n2033), .B(n2064), .Z(n3190) );
  CND3X1 U2942 ( .A(n3188), .B(n3189), .C(n3190), .Z(n1232) );
  CND2X1 U2943 ( .A(n1252), .B(n1225), .Z(n3850) );
  CEOX2 U2944 ( .A(n1225), .B(n1252), .Z(n3847) );
  CND2X1 U2945 ( .A(n3827), .B(n3828), .Z(n3762) );
  COAN1X1 U2946 ( .A(n547), .B(n3866), .C(n3150), .Z(n3731) );
  CENX1 U2947 ( .A(n2802), .B(net18982), .Z(n2703) );
  CEOX2 U2948 ( .A(n1371), .B(n1394), .Z(n3191) );
  CEOX2 U2949 ( .A(n3191), .B(n1369), .Z(n1365) );
  CND2X1 U2950 ( .A(n1369), .B(n1394), .Z(n3192) );
  CND2X1 U2951 ( .A(n1369), .B(n1371), .Z(n3193) );
  CND3X2 U2952 ( .A(n3192), .B(n3193), .C(n3194), .Z(n1364) );
  CIVX1 U2953 ( .A(n1364), .Z(n3344) );
  CIVXL U2954 ( .A(n3487), .Z(n3195) );
  CEO3X1 U2955 ( .A(n1069), .B(n1067), .C(n1090), .Z(n1063) );
  CND2X1 U2956 ( .A(n1069), .B(n1067), .Z(n3196) );
  CND2X1 U2957 ( .A(n1069), .B(n1090), .Z(n3197) );
  CND2X1 U2958 ( .A(n1067), .B(n1090), .Z(n3198) );
  CND3X2 U2959 ( .A(n3196), .B(n3197), .C(n3198), .Z(n1062) );
  CND2XL U2960 ( .A(n1064), .B(n1043), .Z(n3199) );
  CND2X1 U2961 ( .A(n1064), .B(n1062), .Z(n3200) );
  CND2XL U2962 ( .A(n1043), .B(n1062), .Z(n3201) );
  CND3X1 U2963 ( .A(n3199), .B(n3200), .C(n3201), .Z(n1038) );
  COR2X1 U2964 ( .A(n1058), .B(n1037), .Z(n3202) );
  CENX1 U2965 ( .A(n3482), .B(n1096), .Z(n1067) );
  CENX1 U2966 ( .A(n1079), .B(n1073), .Z(n3482) );
  CENX2 U2967 ( .A(net16570), .B(n4291), .Z(n2372) );
  COND2X1 U2968 ( .A(net19122), .B(n2397), .C(net16839), .D(n2396), .Z(n1875)
         );
  COND1X1 U2969 ( .A(n3710), .B(n275), .C(n3981), .Z(n236) );
  CIVX1 U2970 ( .A(n3111), .Z(n273) );
  COND2X1 U2971 ( .A(net19122), .B(n2388), .C(net16839), .D(n2387), .Z(n1868)
         );
  CNR2X1 U2972 ( .A(n81), .B(n2507), .Z(n3870) );
  CND2X2 U2973 ( .A(n4123), .B(n1308), .Z(n4126) );
  CEOX2 U2974 ( .A(n1410), .B(n1402), .Z(n3203) );
  CEOX2 U2975 ( .A(n3203), .B(n1404), .Z(n1375) );
  CND2XL U2976 ( .A(n1404), .B(n1402), .Z(n3204) );
  CND2XL U2977 ( .A(n1402), .B(n1410), .Z(n3206) );
  CND3X1 U2978 ( .A(n3204), .B(n3205), .C(n3206), .Z(n1374) );
  CFA1X1 U2979 ( .A(n2163), .B(n1948), .CI(n1919), .CO(n1404), .S(n1405) );
  CND2X1 U2980 ( .A(n1281), .B(n4205), .Z(n4207) );
  CND2XL U2981 ( .A(n3768), .B(n3208), .Z(n3209) );
  CND2X2 U2982 ( .A(n3207), .B(n1314), .Z(n3210) );
  CND2X2 U2983 ( .A(n3209), .B(n3210), .Z(n1281) );
  CIVXL U2984 ( .A(n1314), .Z(n3208) );
  CENX1 U2985 ( .A(n1110), .B(n3614), .Z(n1085) );
  COND2X2 U2986 ( .A(n81), .B(n2488), .C(net19060), .D(n2487), .Z(n1963) );
  CIVX1 U2987 ( .A(n378), .Z(n745) );
  CIVXL U2988 ( .A(n1308), .Z(n4124) );
  CIVX2 U2989 ( .A(net16644), .Z(n87) );
  CENX1 U2990 ( .A(n4326), .B(n3393), .Z(n2407) );
  COND1X1 U2991 ( .A(n547), .B(n3869), .C(n3946), .Z(n3211) );
  COND1XL U2992 ( .A(n547), .B(n3869), .C(n3946), .Z(n546) );
  CENXL U2993 ( .A(n635), .B(n192), .Z(product[20]) );
  CIVX3 U2994 ( .A(n747), .Z(n3212) );
  CIVX2 U2995 ( .A(n402), .Z(n747) );
  CND3XL U2996 ( .A(n3581), .B(n3583), .C(n3582), .Z(n3213) );
  CND3XL U2997 ( .A(n3581), .B(n3583), .C(n3582), .Z(n1522) );
  CNIVX2 U2998 ( .A(n30), .Z(n3962) );
  CND2X1 U2999 ( .A(n1447), .B(n3215), .Z(n3216) );
  CND2XL U3000 ( .A(n3027), .B(n3214), .Z(n3217) );
  CND2X1 U3001 ( .A(n3216), .B(n3217), .Z(n4115) );
  CIVXL U3002 ( .A(n1447), .Z(n3214) );
  CIVXL U3003 ( .A(n3027), .Z(n3215) );
  CND2X1 U3004 ( .A(n3749), .B(n3750), .Z(n1445) );
  CND2XL U3005 ( .A(n897), .B(n895), .Z(n3274) );
  CND2XL U3006 ( .A(n895), .B(n908), .Z(n3276) );
  CENXL U3007 ( .A(n4325), .B(net18618), .Z(n2507) );
  COND2XL U3008 ( .A(n2745), .B(n4001), .C(net16816), .D(n2744), .Z(n2218) );
  COND2XL U3009 ( .A(n4001), .B(n2739), .C(net16816), .D(n2738), .Z(n2212) );
  COND2XL U3010 ( .A(n4001), .B(n2743), .C(net16816), .D(n2742), .Z(n2216) );
  COND2XL U3011 ( .A(n4001), .B(n2736), .C(net16817), .D(n2735), .Z(n2209) );
  CAOR1XL U3012 ( .A(net16816), .B(n4001), .C(n2714), .Z(n2187) );
  COND2XL U3013 ( .A(n4001), .B(n2741), .C(net16816), .D(n2740), .Z(n2214) );
  COND2XL U3014 ( .A(n4001), .B(n2740), .C(net16816), .D(n2739), .Z(n2213) );
  CND2IX1 U3015 ( .B(n3495), .A(n1189), .Z(n4127) );
  CND2X1 U3016 ( .A(n1215), .B(n1244), .Z(n541) );
  CIVXL U3017 ( .A(n556), .Z(n764) );
  CND2XL U3018 ( .A(n3819), .B(n3880), .Z(n3821) );
  CENX1 U3019 ( .A(n1094), .B(n1071), .Z(n3218) );
  CEOXL U3020 ( .A(n2808), .B(n3384), .Z(n2544) );
  CENX1 U3021 ( .A(net16550), .B(net16824), .Z(n2527) );
  CNIVX2 U3022 ( .A(a[8]), .Z(n4101) );
  CNIVX4 U3023 ( .A(n12), .Z(n3219) );
  CIVX1 U3024 ( .A(n12), .Z(n3999) );
  CNR2X2 U3025 ( .A(n409), .B(n3212), .Z(n3220) );
  CEOX1 U3026 ( .A(n3373), .B(n1583), .Z(n1581) );
  CIVX3 U3027 ( .A(n4359), .Z(n4170) );
  CEOX2 U3028 ( .A(n3221), .B(n1971), .Z(n1211) );
  CND2XL U3029 ( .A(n1971), .B(n3137), .Z(n3222) );
  CND2XL U3030 ( .A(n1971), .B(n1796), .Z(n3223) );
  CND2XL U3031 ( .A(n1853), .B(n1796), .Z(n3224) );
  CND3X1 U3032 ( .A(n3222), .B(n3223), .C(n3224), .Z(n1210) );
  CIVXL U3033 ( .A(net18643), .Z(net18905) );
  CIVX1 U3034 ( .A(n4014), .Z(n4360) );
  CND3XL U3035 ( .A(n4245), .B(n4246), .C(n4247), .Z(n3225) );
  CND2IX1 U3036 ( .B(net16027), .A(a[18]), .Z(n3490) );
  CENX1 U3037 ( .A(n4325), .B(n4254), .Z(n2672) );
  CEO3X1 U3038 ( .A(n1303), .B(n1328), .C(n1330), .Z(n1291) );
  CND2XL U3039 ( .A(n1303), .B(n1330), .Z(n3226) );
  CND2X1 U3040 ( .A(n1303), .B(n1328), .Z(n3227) );
  CND2X1 U3041 ( .A(n1330), .B(n1328), .Z(n3228) );
  CND3X2 U3042 ( .A(n3226), .B(n3227), .C(n3228), .Z(n1290) );
  CEOX1 U3043 ( .A(n1074), .B(n1072), .Z(n4155) );
  CEOX2 U3044 ( .A(n912), .B(n899), .Z(n3229) );
  CEOX2 U3045 ( .A(n910), .B(n3229), .Z(n895) );
  CND2X2 U3046 ( .A(n910), .B(n899), .Z(n3230) );
  CND2X2 U3047 ( .A(n910), .B(n912), .Z(n3231) );
  CND2X1 U3048 ( .A(n899), .B(n912), .Z(n3232) );
  CND3X2 U3049 ( .A(n3230), .B(n3231), .C(n3232), .Z(n894) );
  CIVX1 U3050 ( .A(n1871), .Z(n3233) );
  CIVX3 U3051 ( .A(n3408), .Z(n3822) );
  CENX1 U3052 ( .A(n4171), .B(n3962), .Z(n3235) );
  CENX2 U3053 ( .A(n4171), .B(n3962), .Z(n42) );
  CANR1X2 U3054 ( .A(n3620), .B(n621), .C(n616), .Z(n614) );
  CENX1 U3055 ( .A(n4321), .B(net18643), .Z(n2545) );
  CND2X1 U3056 ( .A(n1125), .B(n1146), .Z(n3396) );
  CND2X1 U3057 ( .A(n1182), .B(n1178), .Z(n3927) );
  CND2X1 U3058 ( .A(n1182), .B(n1180), .Z(n3928) );
  CND2X1 U3059 ( .A(n3461), .B(n1516), .Z(n3457) );
  CEOX1 U3060 ( .A(n2142), .B(n2173), .Z(n3236) );
  CEOX2 U3061 ( .A(n3236), .B(n3037), .Z(n1605) );
  CND2XL U3062 ( .A(n1611), .B(n2173), .Z(n3237) );
  CND2X1 U3063 ( .A(n1611), .B(n2142), .Z(n3238) );
  CND2XL U3064 ( .A(n2173), .B(n2142), .Z(n3239) );
  CND3X1 U3065 ( .A(n3237), .B(n3238), .C(n3239), .Z(n1604) );
  COND2XL U3066 ( .A(n4002), .B(n2669), .C(net19508), .D(n2668), .Z(n2142) );
  COND1XL U3067 ( .A(n385), .B(n4020), .C(n386), .Z(n384) );
  CENX1 U3068 ( .A(n4325), .B(net16067), .Z(n2639) );
  CIVXL U3069 ( .A(n627), .Z(n773) );
  CHA1X1 U3070 ( .A(n1730), .B(n1956), .CO(n1578), .S(n1579) );
  CENXL U3071 ( .A(n4340), .B(n4000), .Z(n2551) );
  CFA1X1 U3072 ( .A(n1808), .B(n1749), .CI(n1896), .CO(n862), .S(n863) );
  COND2X1 U3073 ( .A(n144), .B(n2263), .C(n3576), .D(n2262), .Z(n1749) );
  CNR2X2 U3074 ( .A(n3421), .B(n416), .Z(n3240) );
  COND1X1 U3075 ( .A(n512), .B(n504), .C(n505), .Z(n499) );
  CND2X1 U3076 ( .A(n3881), .B(n767), .Z(n3241) );
  CENXL U3077 ( .A(n4336), .B(net18936), .Z(n2522) );
  CENXL U3078 ( .A(n2789), .B(net16824), .Z(n2525) );
  CENXL U3079 ( .A(net16558), .B(net18936), .Z(n2531) );
  CENX1 U3080 ( .A(n4342), .B(net16824), .Z(n2516) );
  CANR1XL U3081 ( .A(n363), .B(n397), .C(n3468), .Z(n362) );
  CND2XL U3082 ( .A(n3213), .B(n1518), .Z(n3455) );
  CND3X2 U3083 ( .A(n3909), .B(n3910), .C(n3911), .Z(n1066) );
  CENX1 U3084 ( .A(n4326), .B(net18982), .Z(n2704) );
  CND2X1 U3085 ( .A(n3798), .B(n4317), .Z(n177) );
  CIVX2 U3086 ( .A(n1442), .Z(n3743) );
  CEO3X2 U3087 ( .A(n1752), .B(n1929), .C(n1811), .Z(n905) );
  CEOX2 U3088 ( .A(n901), .B(n914), .Z(n3242) );
  CEOX2 U3089 ( .A(n3242), .B(n905), .Z(n897) );
  CND2XL U3090 ( .A(n1752), .B(n1811), .Z(n3244) );
  CND2X1 U3091 ( .A(n1929), .B(n1811), .Z(n3245) );
  CND2XL U3092 ( .A(n901), .B(n914), .Z(n3246) );
  CND2X1 U3093 ( .A(n901), .B(n905), .Z(n3247) );
  CND2X1 U3094 ( .A(n914), .B(n905), .Z(n3248) );
  CND3X1 U3095 ( .A(n3246), .B(n3247), .C(n3248), .Z(n896) );
  COR2X1 U3096 ( .A(n2452), .B(net18592), .Z(n3249) );
  CANR1X2 U3097 ( .A(n686), .B(n4281), .C(n681), .Z(n679) );
  CIVXL U3098 ( .A(net18730), .Z(net18731) );
  COND2X1 U3099 ( .A(n2418), .B(n3920), .C(n2419), .D(n99), .Z(n1897) );
  CND2X1 U3100 ( .A(n396), .B(n363), .Z(n3420) );
  CENX2 U3101 ( .A(n4324), .B(n3729), .Z(n2607) );
  COND2XL U3102 ( .A(n3116), .B(n2290), .C(n3709), .D(n2289), .Z(n1775) );
  CFA1XL U3103 ( .A(n1746), .B(n1864), .CI(n1776), .CO(n830), .S(n831) );
  CEO3X2 U3104 ( .A(n1044), .B(n1023), .C(n1025), .Z(n1019) );
  CND2X1 U3105 ( .A(n1023), .B(n1044), .Z(n3250) );
  CND2X1 U3106 ( .A(n1044), .B(n1025), .Z(n3251) );
  CND2X1 U3107 ( .A(n1023), .B(n1025), .Z(n3252) );
  CND3X2 U3108 ( .A(n3250), .B(n3251), .C(n3252), .Z(n1018) );
  CND2XL U3109 ( .A(n1020), .B(n1001), .Z(n3253) );
  CND2XL U3110 ( .A(n1001), .B(n1018), .Z(n3255) );
  CND3X1 U3111 ( .A(n3253), .B(n3254), .C(n3255), .Z(n996) );
  CEOX1 U3112 ( .A(n1185), .B(n2093), .Z(n3256) );
  CEOX1 U3113 ( .A(n3256), .B(n1212), .Z(n1175) );
  CND2XL U3114 ( .A(n1212), .B(n2093), .Z(n3257) );
  CND2X1 U3115 ( .A(n1212), .B(n1185), .Z(n3258) );
  CND2XL U3116 ( .A(n2093), .B(n1185), .Z(n3259) );
  CND3XL U3117 ( .A(n3257), .B(n3258), .C(n3259), .Z(n1174) );
  COND1X1 U3118 ( .A(n480), .B(n3871), .C(n3834), .Z(n3260) );
  COND1XL U3119 ( .A(n480), .B(n3038), .C(n3834), .Z(n3879) );
  CANR1XL U3120 ( .A(n419), .B(n387), .C(n388), .Z(n386) );
  CANR1XL U3121 ( .A(n478), .B(n546), .C(n3879), .Z(net18543) );
  CEO3XL U3122 ( .A(n1041), .B(n1039), .C(n1060), .Z(n3261) );
  COND2X1 U3123 ( .A(n3877), .B(n2612), .C(net18731), .D(n2611), .Z(n2085) );
  COND1X2 U3124 ( .A(n480), .B(n515), .C(n481), .Z(n479) );
  CND2X4 U3125 ( .A(n114), .B(n4010), .Z(n117) );
  COND2XL U3126 ( .A(n2286), .B(n3709), .C(n2287), .D(n3116), .Z(n1773) );
  COND2XL U3127 ( .A(n3116), .B(n2288), .C(n3709), .D(n2287), .Z(n810) );
  COND2XL U3128 ( .A(n3116), .B(n2289), .C(n3709), .D(n2288), .Z(n1774) );
  COND2XL U3129 ( .A(n3116), .B(n2292), .C(n3709), .D(n2291), .Z(n1777) );
  COND2XL U3130 ( .A(n3116), .B(n2293), .C(n3709), .D(n2292), .Z(n1778) );
  COND2XL U3131 ( .A(n3116), .B(n2291), .C(n3709), .D(n2290), .Z(n1776) );
  COND2XL U3132 ( .A(n4136), .B(n2296), .C(n3709), .D(n2295), .Z(n1781) );
  CND2X1 U3133 ( .A(a[26]), .B(n4358), .Z(n3264) );
  CND2X2 U3134 ( .A(n3263), .B(n3262), .Z(n3265) );
  CND2X4 U3135 ( .A(n3264), .B(n3265), .Z(net18254) );
  CIVX1 U3136 ( .A(a[26]), .Z(n3262) );
  CIVX3 U3137 ( .A(net18254), .Z(net16800) );
  CIVX3 U3138 ( .A(net18254), .Z(net16801) );
  CIVXL U3139 ( .A(n745), .Z(n3266) );
  CIVXL U3140 ( .A(n3266), .Z(n3267) );
  CANR1XL U3141 ( .A(n432), .B(n3129), .C(n423), .Z(n3268) );
  CANR1X1 U3142 ( .A(n432), .B(n3129), .C(n423), .Z(n3269) );
  CANR1X1 U3143 ( .A(n432), .B(n3129), .C(n423), .Z(n417) );
  CEO3X2 U3144 ( .A(n928), .B(n926), .C(n913), .Z(n909) );
  CND2XL U3145 ( .A(n928), .B(n926), .Z(n3270) );
  CND2X1 U3146 ( .A(n928), .B(n913), .Z(n3271) );
  CND2XL U3147 ( .A(n926), .B(n913), .Z(n3272) );
  CND3X1 U3148 ( .A(n3270), .B(n3271), .C(n3272), .Z(n908) );
  CEOX2 U3149 ( .A(n897), .B(n895), .Z(n3273) );
  CEOX2 U3150 ( .A(n3273), .B(n908), .Z(n893) );
  CND2X1 U3151 ( .A(n897), .B(n908), .Z(n3275) );
  CND3X1 U3152 ( .A(n3274), .B(n3275), .C(n3276), .Z(n892) );
  CIVX4 U3153 ( .A(net16644), .Z(n3277) );
  CIVX4 U3154 ( .A(net16644), .Z(n3278) );
  CENX2 U3155 ( .A(n4340), .B(n3730), .Z(n2584) );
  CANR1X1 U3156 ( .A(n478), .B(net19465), .C(n479), .Z(n3279) );
  CANR1X1 U3157 ( .A(n478), .B(net19465), .C(n479), .Z(n3280) );
  CANR1X1 U3158 ( .A(n478), .B(net19465), .C(n479), .Z(n149) );
  CIVX1 U3159 ( .A(n1080), .Z(n1081) );
  CNR2X2 U3160 ( .A(n923), .B(n938), .Z(n409) );
  CNIVX4 U3161 ( .A(net19048), .Z(net16788) );
  CIVXL U3162 ( .A(n440), .Z(n3281) );
  CIVXL U3163 ( .A(n3202), .Z(n3282) );
  CENX1 U3164 ( .A(n4341), .B(net16824), .Z(n2517) );
  CIVX1 U3165 ( .A(n2056), .Z(n3357) );
  COND2X2 U3166 ( .A(n2583), .B(n3877), .C(n3839), .D(n2582), .Z(n2056) );
  CEO3X2 U3167 ( .A(n1994), .B(n2055), .C(n1964), .Z(n1007) );
  CND2XL U3168 ( .A(n1994), .B(n1964), .Z(n3283) );
  CND2XL U3169 ( .A(n1994), .B(n2055), .Z(n3284) );
  CND2XL U3170 ( .A(n1964), .B(n2055), .Z(n3285) );
  CND3X1 U3171 ( .A(n3283), .B(n3284), .C(n3285), .Z(n1006) );
  CNR2XL U3172 ( .A(net18670), .B(n2520), .Z(n3286) );
  CNR2XL U3173 ( .A(n4144), .B(n2519), .Z(n3287) );
  COR2X1 U3174 ( .A(n3286), .B(n3287), .Z(n1994) );
  COND2XL U3175 ( .A(n81), .B(n2489), .C(net19060), .D(n2488), .Z(n1964) );
  CND2XL U3176 ( .A(n1277), .B(n1279), .Z(n4091) );
  CND2X1 U3177 ( .A(n776), .B(n4274), .Z(n636) );
  CANR1X2 U3178 ( .A(n349), .B(n4279), .C(n340), .Z(n334) );
  CIVXL U3179 ( .A(n334), .Z(n332) );
  CANR1X2 U3180 ( .A(n576), .B(net18451), .C(n577), .Z(n3869) );
  CANR1XL U3181 ( .A(n576), .B(net18451), .C(n577), .Z(n3866) );
  CND2X1 U3182 ( .A(n1311), .B(n1336), .Z(n4122) );
  COND2XL U3183 ( .A(n4033), .B(n2367), .C(net16784), .D(n2366), .Z(n1847) );
  COND2X1 U3184 ( .A(n2578), .B(n4135), .C(net19500), .D(n2577), .Z(n2051) );
  CIVX1 U3185 ( .A(net19505), .Z(n3288) );
  CND2X1 U3186 ( .A(a[28]), .B(net15997), .Z(n3291) );
  CND2X2 U3187 ( .A(n3289), .B(n3290), .Z(n3292) );
  CND2X4 U3188 ( .A(n3291), .B(n3292), .Z(n132) );
  CIVX2 U3189 ( .A(a[28]), .Z(n3289) );
  CIVX2 U3190 ( .A(net15997), .Z(n3290) );
  CIVX2 U3191 ( .A(net19505), .Z(net15997) );
  CNR2IX2 U3192 ( .B(net16109), .A(n132), .Z(n1802) );
  CNR2X1 U3193 ( .A(n636), .B(n3102), .Z(n3480) );
  CND2IX2 U3194 ( .B(n1313), .A(n3444), .Z(n3446) );
  COND1X2 U3195 ( .A(n628), .B(n622), .C(n623), .Z(n621) );
  CEO3X2 U3196 ( .A(n1068), .B(n1049), .C(n1070), .Z(n1043) );
  COR2XL U3197 ( .A(n1580), .B(n1563), .Z(n3756) );
  CAOR1XL U3198 ( .A(n3839), .B(n3877), .C(n2582), .Z(n2055) );
  CEO3X2 U3199 ( .A(n1758), .B(n1034), .C(n2024), .Z(n1013) );
  CND2XL U3200 ( .A(n1758), .B(n2024), .Z(n3293) );
  CND2XL U3201 ( .A(n1758), .B(n1034), .Z(n3294) );
  CND3X1 U3202 ( .A(n3293), .B(n3294), .C(n3295), .Z(n1012) );
  CND2XL U3203 ( .A(n1009), .B(n1011), .Z(n3296) );
  CND2XL U3204 ( .A(n1009), .B(n1013), .Z(n3297) );
  CND2XL U3205 ( .A(n1011), .B(n1013), .Z(n3298) );
  CND3X1 U3206 ( .A(n3296), .B(n3297), .C(n3298), .Z(n1002) );
  CIVXL U3207 ( .A(n559), .Z(n3299) );
  CIVXL U3208 ( .A(n3299), .Z(n3300) );
  CIVX2 U3209 ( .A(n1336), .Z(n3763) );
  CAOR1X1 U3210 ( .A(n520), .B(n3829), .C(n3535), .Z(n4053) );
  CEO3X1 U3211 ( .A(n988), .B(n969), .C(n986), .Z(n965) );
  CND2XL U3212 ( .A(n988), .B(n986), .Z(n3302) );
  CND2X1 U3213 ( .A(n969), .B(n986), .Z(n3303) );
  CND3X2 U3214 ( .A(n3301), .B(n3302), .C(n3303), .Z(n964) );
  CEOX2 U3215 ( .A(n966), .B(n947), .Z(n3304) );
  CEOX2 U3216 ( .A(n3304), .B(n964), .Z(n943) );
  CND2X1 U3217 ( .A(n966), .B(n947), .Z(n3305) );
  CND2X1 U3218 ( .A(n966), .B(n964), .Z(n3306) );
  CND2X1 U3219 ( .A(n947), .B(n964), .Z(n3307) );
  CIVXL U3220 ( .A(n4356), .Z(n3308) );
  CND2X1 U3221 ( .A(n1071), .B(n1094), .Z(n3525) );
  CND2X4 U3222 ( .A(n114), .B(n2815), .Z(n4033) );
  COND2XL U3223 ( .A(n99), .B(n2428), .C(n3920), .D(n2427), .Z(n3309) );
  CANR1X2 U3224 ( .A(n736), .B(n273), .C(n264), .Z(n262) );
  CFA1X1 U3225 ( .A(n1815), .B(n1903), .CI(n1786), .CO(n970), .S(n971) );
  CND2X1 U3226 ( .A(n1761), .B(n3022), .Z(n3589) );
  CANR1X2 U3227 ( .A(n478), .B(n3211), .C(n3260), .Z(net19409) );
  CENXL U3228 ( .A(n1110), .B(n3614), .Z(n3310) );
  COND2XL U3229 ( .A(n2385), .B(net16839), .C(n2386), .D(net19122), .Z(n1866)
         );
  CAOR1XL U3230 ( .A(net16839), .B(net19122), .C(n2384), .Z(n1864) );
  CDLY1XL U3231 ( .A(n3030), .Z(n3311) );
  CANR1XL U3232 ( .A(n669), .B(n677), .C(n670), .Z(n3312) );
  CANR1XL U3233 ( .A(n669), .B(n677), .C(n670), .Z(n3313) );
  CANR1X1 U3234 ( .A(n669), .B(n677), .C(n670), .Z(n668) );
  COND2XL U3235 ( .A(n2451), .B(net18593), .C(n3278), .D(n2450), .Z(n1928) );
  CENXL U3236 ( .A(n4322), .B(n3487), .Z(n2477) );
  CND2X1 U3237 ( .A(n1474), .B(n1476), .Z(n3513) );
  CND3XL U3238 ( .A(n3697), .B(n3699), .C(n3698), .Z(n3314) );
  CND3XL U3239 ( .A(n3697), .B(n3699), .C(n3698), .Z(n1510) );
  CND2XL U3240 ( .A(n1312), .B(n1285), .Z(n4178) );
  CND2X1 U3241 ( .A(n3737), .B(n3316), .Z(n3317) );
  CND2X2 U3242 ( .A(n3315), .B(n972), .Z(n3318) );
  CND2X2 U3243 ( .A(n3317), .B(n3318), .Z(n947) );
  CIVX2 U3244 ( .A(n3737), .Z(n3315) );
  CIVXL U3245 ( .A(n972), .Z(n3316) );
  CIVXL U3246 ( .A(n4268), .Z(n3319) );
  CIVXL U3247 ( .A(n3319), .Z(n3320) );
  CEO3X1 U3248 ( .A(n1241), .B(n1237), .C(n1260), .Z(n1225) );
  CND2XL U3249 ( .A(n1241), .B(n1260), .Z(n3321) );
  CND2XL U3250 ( .A(n1241), .B(n1237), .Z(n3322) );
  CND2X1 U3251 ( .A(n1260), .B(n1237), .Z(n3323) );
  CEO3X1 U3252 ( .A(n1201), .B(n1224), .C(n3398), .Z(n3615) );
  CEOX2 U3253 ( .A(n1183), .B(n1181), .Z(n3324) );
  CEOX2 U3254 ( .A(n3324), .B(n1202), .Z(n1169) );
  CND2X1 U3255 ( .A(n1202), .B(n1181), .Z(n3325) );
  CND2X1 U3256 ( .A(n1202), .B(n1183), .Z(n3326) );
  CND2XL U3257 ( .A(n1181), .B(n1183), .Z(n3327) );
  CND3X2 U3258 ( .A(n3325), .B(n3326), .C(n3327), .Z(n1168) );
  CND3X2 U3259 ( .A(n3390), .B(n3391), .C(n3392), .Z(n1202) );
  CND2X1 U3260 ( .A(n1168), .B(n1147), .Z(n3475) );
  CND3X2 U3261 ( .A(net19203), .B(net19205), .C(net19204), .Z(n1336) );
  CIVXL U3262 ( .A(n534), .Z(n532) );
  CND2X1 U3263 ( .A(n3490), .B(n3489), .Z(n3328) );
  CND2X1 U3264 ( .A(n3489), .B(n3490), .Z(n3872) );
  CEOX1 U3265 ( .A(n2030), .B(n2061), .Z(n3329) );
  CEOX1 U3266 ( .A(n3329), .B(n2154), .Z(n1149) );
  CND2XL U3267 ( .A(n2154), .B(n2030), .Z(n3330) );
  CND2XL U3268 ( .A(n2154), .B(n2061), .Z(n3331) );
  CND2XL U3269 ( .A(n2030), .B(n2061), .Z(n3332) );
  CND3X1 U3270 ( .A(n3330), .B(n3331), .C(n3332), .Z(n1148) );
  CEO3XL U3271 ( .A(n1116), .B(n1097), .C(n1095), .Z(n3333) );
  COND2X2 U3272 ( .A(n2682), .B(n3678), .C(n2683), .D(n27), .Z(n2156) );
  CEO3X2 U3273 ( .A(n1309), .B(n1334), .C(n3625), .Z(net19127) );
  CNR2X1 U3274 ( .A(n3854), .B(n3853), .Z(n3864) );
  CIVX1 U3275 ( .A(n1259), .Z(n3854) );
  CND2X1 U3276 ( .A(n1251), .B(n1278), .Z(n4182) );
  CND2XL U3277 ( .A(n1162), .B(n1164), .Z(n4038) );
  CIVXL U3278 ( .A(n102), .Z(n3334) );
  CIVX2 U3279 ( .A(n102), .Z(n4356) );
  COR2X1 U3280 ( .A(n4144), .B(n2539), .Z(n3806) );
  CENX1 U3281 ( .A(n2808), .B(n4000), .Z(n2577) );
  CND2X1 U3282 ( .A(n2003), .B(n1884), .Z(n4131) );
  CND3X2 U3283 ( .A(n3848), .B(n3849), .C(n3850), .Z(n1218) );
  CND2X1 U3284 ( .A(n3466), .B(n3467), .Z(n3637) );
  CIVX1 U3285 ( .A(net19076), .Z(n3539) );
  CND2X1 U3286 ( .A(n4170), .B(a[28]), .Z(n3337) );
  CND2X2 U3287 ( .A(n3335), .B(n3336), .Z(n3338) );
  CND2X2 U3288 ( .A(n3337), .B(n3338), .Z(n3890) );
  CIVX2 U3289 ( .A(n4170), .Z(n3335) );
  CIVX1 U3290 ( .A(a[28]), .Z(n3336) );
  CND2X2 U3291 ( .A(n4075), .B(n4074), .Z(n1904) );
  CND2X1 U3292 ( .A(n3830), .B(n3138), .Z(n3340) );
  CND2X2 U3293 ( .A(n3339), .B(n1247), .Z(n3341) );
  CND2X2 U3294 ( .A(n3340), .B(n3341), .Z(n1245) );
  CIVX2 U3295 ( .A(n3830), .Z(n3339) );
  COR2XL U3296 ( .A(n1245), .B(n1274), .Z(n3342) );
  CND2X1 U3297 ( .A(n3807), .B(n3344), .Z(n3345) );
  CND2X2 U3298 ( .A(n3343), .B(n1364), .Z(n3346) );
  CND2X2 U3299 ( .A(n3345), .B(n3346), .Z(n1335) );
  CIVX2 U3300 ( .A(n3807), .Z(n3343) );
  CND2XL U3301 ( .A(n869), .B(n880), .Z(n3347) );
  CND2X1 U3302 ( .A(n869), .B(n871), .Z(n3348) );
  CND2XL U3303 ( .A(n880), .B(n871), .Z(n3349) );
  CND3XL U3304 ( .A(n3347), .B(n3348), .C(n3349), .Z(n866) );
  CEO3X1 U3305 ( .A(n1898), .B(n1869), .C(n1751), .Z(n887) );
  CND2XL U3306 ( .A(n1898), .B(n1751), .Z(n3350) );
  CND2XL U3307 ( .A(n1898), .B(n1869), .Z(n3351) );
  CND2XL U3308 ( .A(n1751), .B(n1869), .Z(n3352) );
  CND3X1 U3309 ( .A(n3350), .B(n3351), .C(n3352), .Z(n886) );
  COR2X2 U3310 ( .A(n855), .B(n866), .Z(n4275) );
  COND2XL U3311 ( .A(n144), .B(n2265), .C(n3577), .D(n2264), .Z(n1751) );
  COND2XL U3312 ( .A(n2389), .B(n4188), .C(net19462), .D(n2388), .Z(n1869) );
  COND2XL U3313 ( .A(n99), .B(n2420), .C(n3919), .D(n2419), .Z(n1898) );
  CND2XL U3314 ( .A(n1205), .B(n1211), .Z(n4140) );
  CNR2X2 U3315 ( .A(n1505), .B(n1524), .Z(n622) );
  CENX2 U3316 ( .A(n2789), .B(n4253), .Z(n2393) );
  CND2XL U3317 ( .A(n1068), .B(n1070), .Z(n3353) );
  CND2XL U3318 ( .A(n1068), .B(n1049), .Z(n3354) );
  CND2X1 U3319 ( .A(n1070), .B(n1049), .Z(n3355) );
  CND3XL U3320 ( .A(n3353), .B(n3354), .C(n3355), .Z(n1042) );
  CND3XL U3321 ( .A(n4048), .B(n4049), .C(n4050), .Z(n1070) );
  CIVX2 U3322 ( .A(n354), .Z(n356) );
  CND3X2 U3323 ( .A(n3956), .B(n3958), .C(n3957), .Z(n1254) );
  CND2X1 U3324 ( .A(n1875), .B(n3357), .Z(n3358) );
  CND2X1 U3325 ( .A(n3356), .B(n2056), .Z(n3359) );
  CND2X2 U3326 ( .A(n3358), .B(n3359), .Z(n3368) );
  COND1X2 U3327 ( .A(n444), .B(n461), .C(n3982), .Z(n3659) );
  COND2X1 U3328 ( .A(n117), .B(n2359), .C(net16784), .D(n2358), .Z(n1840) );
  COND2X1 U3329 ( .A(n2514), .B(n81), .C(net19060), .D(n2513), .Z(n1988) );
  CENX1 U3330 ( .A(net16544), .B(n3730), .Z(n2590) );
  CIVXL U3331 ( .A(n1278), .Z(n3360) );
  CND3X1 U3332 ( .A(n4177), .B(n4178), .C(n4179), .Z(n1278) );
  CNIVX2 U3333 ( .A(n1217), .Z(n4032) );
  CND3X1 U3334 ( .A(n4247), .B(n4246), .C(n4245), .Z(n1194) );
  CIVX4 U3335 ( .A(n3377), .Z(n3920) );
  CENXL U3336 ( .A(n1306), .B(n1279), .Z(n3362) );
  CENX1 U3337 ( .A(n4321), .B(n4291), .Z(n2380) );
  CENX1 U3338 ( .A(n1113), .B(n1138), .Z(n3363) );
  CND2XL U3339 ( .A(n2188), .B(n1942), .Z(n4167) );
  CND3X1 U3340 ( .A(n3667), .B(n3668), .C(n3669), .Z(n1562) );
  CEO3X1 U3341 ( .A(n1564), .B(n1549), .C(n1547), .Z(n1545) );
  CND3X2 U3342 ( .A(n4082), .B(n4084), .C(n4083), .Z(n1564) );
  CND2X1 U3343 ( .A(n1584), .B(n1571), .Z(n4082) );
  COND2XL U3344 ( .A(n3024), .B(n2710), .C(net16772), .D(n2709), .Z(n2183) );
  COND2XL U3345 ( .A(n2712), .B(net18743), .C(net16772), .D(n2711), .Z(n2185)
         );
  COND2XL U3346 ( .A(net18743), .B(n2707), .C(net16772), .D(n2706), .Z(n2180)
         );
  CENXL U3347 ( .A(n4322), .B(n4291), .Z(n3364) );
  CND2XL U3348 ( .A(n1828), .B(n1856), .Z(n3365) );
  CND2XL U3349 ( .A(n1828), .B(n2066), .Z(n3366) );
  CND2X1 U3350 ( .A(n1856), .B(n2066), .Z(n3367) );
  CND3X2 U3351 ( .A(n3365), .B(n3366), .C(n3367), .Z(n1294) );
  CND2X1 U3352 ( .A(n3372), .B(n2056), .Z(n3369) );
  CND2XL U3353 ( .A(n1875), .B(n2056), .Z(n3371) );
  CNIVX2 U3354 ( .A(n1759), .Z(n3372) );
  COR2X1 U3355 ( .A(n3919), .B(n2425), .Z(n4075) );
  CEOX2 U3356 ( .A(n1598), .B(n1585), .Z(n3373) );
  CND2XL U3357 ( .A(n1583), .B(n1585), .Z(n3374) );
  CND2XL U3358 ( .A(n1583), .B(n1598), .Z(n3375) );
  CND2XL U3359 ( .A(n1585), .B(n1598), .Z(n3376) );
  CND3X1 U3360 ( .A(n3374), .B(n3375), .C(n3376), .Z(n1580) );
  CND2X1 U3361 ( .A(n1581), .B(n1596), .Z(n644) );
  CND3X2 U3362 ( .A(n3511), .B(n3512), .C(n3513), .Z(n1446) );
  CIVX2 U3363 ( .A(n3124), .Z(n3378) );
  CND2X1 U3364 ( .A(n1429), .B(n1435), .Z(n3379) );
  CND2X1 U3365 ( .A(n1429), .B(n1454), .Z(n3380) );
  CND2XL U3366 ( .A(n1435), .B(n1454), .Z(n3381) );
  CND3X1 U3367 ( .A(n3379), .B(n3380), .C(n3381), .Z(n1422) );
  CEOX1 U3368 ( .A(n3683), .B(n1421), .Z(n3382) );
  CIVX1 U3369 ( .A(n1423), .Z(n3610) );
  CEOXL U3370 ( .A(n3683), .B(n1421), .Z(n1417) );
  CIVX2 U3371 ( .A(n1311), .Z(n3444) );
  CND2XL U3372 ( .A(a[16]), .B(n3868), .Z(n3385) );
  CND2X1 U3373 ( .A(n3383), .B(n3384), .Z(n3386) );
  CND2X2 U3374 ( .A(n3385), .B(n3386), .Z(n3867) );
  CIVXL U3375 ( .A(a[16]), .Z(n3383) );
  CIVX1 U3376 ( .A(n3868), .Z(n3384) );
  CEO3X1 U3377 ( .A(n1913), .B(n1797), .C(n2157), .Z(n1239) );
  CND2XL U3378 ( .A(n1913), .B(n1797), .Z(n3387) );
  CND2XL U3379 ( .A(n1913), .B(n2157), .Z(n3388) );
  CND2X1 U3380 ( .A(n1797), .B(n2157), .Z(n3389) );
  CND2XL U3381 ( .A(n2187), .B(n1240), .Z(n3390) );
  CND2XL U3382 ( .A(n2187), .B(n1238), .Z(n3391) );
  CND2XL U3383 ( .A(n1240), .B(n1238), .Z(n3392) );
  CIVX2 U3384 ( .A(n4087), .Z(n3393) );
  CIVX4 U3385 ( .A(n4354), .Z(n4087) );
  CIVX1 U3386 ( .A(n3416), .Z(n3417) );
  CND3X1 U3387 ( .A(n3394), .B(n3395), .C(n3396), .Z(n1114) );
  CND3X2 U3388 ( .A(n3927), .B(n3928), .C(n3929), .Z(n1146) );
  CIVXL U3389 ( .A(n1199), .Z(n3397) );
  CENX2 U3390 ( .A(n1441), .B(n1462), .Z(n4271) );
  COND2X2 U3391 ( .A(n126), .B(n2346), .C(net16801), .D(n2345), .Z(n1829) );
  CIVX2 U3392 ( .A(n3912), .Z(n3633) );
  COR2X1 U3393 ( .A(n1437), .B(n1460), .Z(n4267) );
  CEOX2 U3394 ( .A(n911), .B(n924), .Z(n3399) );
  CEOX2 U3395 ( .A(n3399), .B(n909), .Z(n907) );
  CND2XL U3396 ( .A(n909), .B(n924), .Z(n3400) );
  CND2X1 U3397 ( .A(n909), .B(n911), .Z(n3401) );
  CND2XL U3398 ( .A(n924), .B(n911), .Z(n3402) );
  CND3X1 U3399 ( .A(n3400), .B(n3401), .C(n3402), .Z(n906) );
  CFA1X1 U3400 ( .A(n1785), .B(n1902), .CI(n1814), .CO(n950), .S(n951) );
  CIVX2 U3401 ( .A(net18981), .Z(net18982) );
  CND3X1 U3402 ( .A(n3517), .B(n3518), .C(n3519), .Z(n974) );
  CND2IX1 U3403 ( .B(n3695), .A(n1569), .Z(n4084) );
  CNIVX1 U3404 ( .A(n1982), .Z(n3404) );
  COND2XL U3405 ( .A(n2352), .B(n4033), .C(n3032), .D(n2351), .Z(n1835) );
  COND2XL U3406 ( .A(n4033), .B(n2354), .C(n3032), .D(n2353), .Z(n1837) );
  CFA1XL U3407 ( .A(n842), .B(n1836), .CI(n1806), .CO(n832), .S(n833) );
  CFA1XL U3408 ( .A(n1745), .B(n1835), .CI(n1775), .CO(n822), .S(n823) );
  CFA1XL U3409 ( .A(n1778), .B(n1838), .CI(n1748), .CO(n850), .S(n851) );
  CEO3X1 U3410 ( .A(n1820), .B(n1761), .C(n3022), .Z(n1075) );
  CND3X1 U3411 ( .A(n4222), .B(n4223), .C(n4224), .Z(n3405) );
  CND3XL U3412 ( .A(n4223), .B(n4222), .C(n4224), .Z(n1082) );
  CENX1 U3413 ( .A(n2802), .B(n3730), .Z(n2604) );
  CND2X1 U3414 ( .A(n1325), .B(n1348), .Z(n3765) );
  COND2XL U3415 ( .A(n2385), .B(n4188), .C(net19462), .D(n2384), .Z(n1865) );
  COND2XL U3416 ( .A(net18607), .B(n2508), .C(net19061), .D(n2507), .Z(n1982)
         );
  CENX1 U3417 ( .A(n2808), .B(n3729), .Z(n2610) );
  CENX1 U3418 ( .A(net16550), .B(net16067), .Z(n2626) );
  CND2XL U3419 ( .A(n3446), .B(n3445), .Z(n3406) );
  CIVXL U3420 ( .A(n3891), .Z(n3407) );
  CENX1 U3421 ( .A(a[18]), .B(n3986), .Z(n3408) );
  CIVX1 U3422 ( .A(n448), .Z(n751) );
  CND2XL U3423 ( .A(n462), .B(n3320), .Z(n451) );
  CNIVX2 U3424 ( .A(n1190), .Z(n3409) );
  CENXL U3425 ( .A(n4338), .B(n4254), .Z(n2652) );
  CENX1 U3426 ( .A(n4340), .B(n4254), .Z(n2650) );
  CENX2 U3427 ( .A(n1389), .B(n4269), .Z(n3481) );
  CIVXL U3428 ( .A(n1205), .Z(n3410) );
  CIVX2 U3429 ( .A(n644), .Z(n3411) );
  CND2X1 U3430 ( .A(n1251), .B(n1253), .Z(n4180) );
  CND2X4 U3431 ( .A(n4256), .B(n4257), .Z(n3412) );
  CFA1XL U3432 ( .A(n2243), .B(n2181), .CI(n1735), .CO(n1696), .S(n1697) );
  CND2IX1 U3433 ( .B(n3494), .A(n1189), .Z(n4128) );
  CENX2 U3434 ( .A(n1414), .B(n1391), .Z(n4269) );
  CIVXL U3435 ( .A(n389), .Z(n746) );
  CND2IX1 U3436 ( .B(n4305), .A(n3413), .Z(n1855) );
  COR2XL U3437 ( .A(net16784), .B(n2374), .Z(n3413) );
  CIVX1 U3438 ( .A(n4008), .Z(n3414) );
  CIVXL U3439 ( .A(n1262), .Z(n3416) );
  CNIVX1 U3440 ( .A(n1296), .Z(n3418) );
  CENX1 U3441 ( .A(n1995), .B(n3419), .Z(n1029) );
  CENX1 U3442 ( .A(n1936), .B(n1818), .Z(n3419) );
  CIVX2 U3443 ( .A(n643), .Z(n776) );
  CNR2X2 U3444 ( .A(n1015), .B(n1036), .Z(n468) );
  COR2X1 U3445 ( .A(n1665), .B(n1674), .Z(n4281) );
  CND2X1 U3446 ( .A(n396), .B(n363), .Z(n3421) );
  CIVX2 U3447 ( .A(n970), .Z(n3570) );
  CND2X2 U3448 ( .A(n1341), .B(n3423), .Z(n3424) );
  CND2X1 U3449 ( .A(n3422), .B(n1339), .Z(n3425) );
  CND2X2 U3450 ( .A(n3425), .B(n3424), .Z(n3807) );
  CND2XL U3451 ( .A(n1345), .B(n3776), .Z(n3428) );
  CND2X2 U3452 ( .A(n3426), .B(n3427), .Z(n3429) );
  CND2X2 U3453 ( .A(n3428), .B(n3429), .Z(n1339) );
  CIVXL U3454 ( .A(n1345), .Z(n3426) );
  CIVX1 U3455 ( .A(n3776), .Z(n3427) );
  CND2X1 U3456 ( .A(n1339), .B(n1341), .Z(n3810) );
  CEO3X1 U3457 ( .A(n1851), .B(n1970), .C(n1184), .Z(n1153) );
  CND2XL U3458 ( .A(n1851), .B(n1970), .Z(n3430) );
  CND2XL U3459 ( .A(n1851), .B(n1184), .Z(n3431) );
  CND2X1 U3460 ( .A(n1970), .B(n1184), .Z(n3432) );
  CND3X1 U3461 ( .A(n3430), .B(n3431), .C(n3432), .Z(n1152) );
  CEOX2 U3462 ( .A(n1150), .B(n1148), .Z(n3433) );
  CEOX2 U3463 ( .A(n3433), .B(n1152), .Z(n1119) );
  CND2X1 U3464 ( .A(n1150), .B(n1152), .Z(n3435) );
  CND3X1 U3465 ( .A(n3434), .B(n3436), .C(n3435), .Z(n1118) );
  CFA1X1 U3466 ( .A(n2087), .B(n2211), .CI(n2149), .CO(n1690), .S(n1691) );
  CNIVX2 U3467 ( .A(n2115), .Z(n3437) );
  CND2XL U3468 ( .A(n3225), .B(n1169), .Z(n3915) );
  CND2X1 U3469 ( .A(n1290), .B(n1263), .Z(n3958) );
  CND2X1 U3470 ( .A(n1290), .B(n1267), .Z(n3956) );
  CIVX3 U3471 ( .A(n4346), .Z(n4344) );
  CND2X1 U3472 ( .A(n3362), .B(n1277), .Z(n3440) );
  CND2X2 U3473 ( .A(n3439), .B(n3438), .Z(n3441) );
  CIVX2 U3474 ( .A(n3964), .Z(n3438) );
  CIVX1 U3475 ( .A(n1277), .Z(n3439) );
  CENX1 U3476 ( .A(n1306), .B(n1279), .Z(n3964) );
  CENX1 U3477 ( .A(n4334), .B(n4253), .Z(n2396) );
  CENX2 U3478 ( .A(a[16]), .B(net18937), .Z(n3875) );
  CND2X4 U3479 ( .A(net18608), .B(a[16]), .Z(n4257) );
  CEO3X1 U3480 ( .A(n1008), .B(n987), .C(n1006), .Z(n983) );
  CEOX1 U3481 ( .A(n3882), .B(n941), .Z(n939) );
  CENX1 U3482 ( .A(n1108), .B(n3132), .Z(n3865) );
  CND2X1 U3483 ( .A(n1166), .B(n1143), .Z(n3585) );
  CENXL U3484 ( .A(n4326), .B(n3730), .Z(n3443) );
  CNIVX2 U3485 ( .A(n72), .Z(net19518) );
  CIVX4 U3486 ( .A(n3), .Z(n4346) );
  CIVX4 U3487 ( .A(net18618), .Z(net18608) );
  CENX2 U3488 ( .A(n3361), .B(n4107), .Z(n1247) );
  CNR2X2 U3489 ( .A(n333), .B(n324), .Z(n320) );
  CND2X2 U3490 ( .A(n4275), .B(n4279), .Z(n333) );
  COND2XL U3491 ( .A(net18670), .B(n2529), .C(n4289), .D(n2528), .Z(n4044) );
  CND2X1 U3492 ( .A(n1311), .B(n1313), .Z(n3445) );
  CND2X2 U3493 ( .A(n3445), .B(n3446), .Z(n3932) );
  CENX1 U3494 ( .A(n4322), .B(net15995), .Z(n2345) );
  CENX2 U3495 ( .A(n3447), .B(n1390), .Z(n1363) );
  CENX2 U3496 ( .A(n1392), .B(n1367), .Z(n3447) );
  CNR2X1 U3497 ( .A(n975), .B(n994), .Z(n448) );
  CIVXL U3498 ( .A(n3313), .Z(n667) );
  CENX1 U3499 ( .A(n4015), .B(n3752), .Z(n1091) );
  CENX2 U3500 ( .A(n3448), .B(n1236), .Z(n1201) );
  CEOX2 U3501 ( .A(n1395), .B(n1416), .Z(n3450) );
  CEOX2 U3502 ( .A(n3450), .B(n1393), .Z(n1389) );
  CND2XL U3503 ( .A(n1393), .B(n1416), .Z(n3451) );
  CND2X1 U3504 ( .A(n1393), .B(n1395), .Z(n3452) );
  CND2XL U3505 ( .A(n1416), .B(n1395), .Z(n3453) );
  CND3X1 U3506 ( .A(n3451), .B(n3452), .C(n3453), .Z(n1388) );
  CND2XL U3507 ( .A(n1820), .B(n1997), .Z(n3588) );
  CND2XL U3508 ( .A(n1565), .B(n1567), .Z(n3667) );
  CIVX2 U3509 ( .A(n434), .Z(n432) );
  CEO3X2 U3510 ( .A(n1522), .B(n1516), .C(n3462), .Z(n1493) );
  CEOX1 U3511 ( .A(n1512), .B(n3042), .Z(n3454) );
  CEOX2 U3512 ( .A(n3454), .B(n1493), .Z(n1487) );
  CND2X1 U3513 ( .A(n3213), .B(n1516), .Z(n3456) );
  CND3X2 U3514 ( .A(n3455), .B(n3456), .C(n3457), .Z(n1492) );
  CND2XL U3515 ( .A(n3314), .B(n1512), .Z(n3458) );
  CND2X1 U3516 ( .A(n1512), .B(n1493), .Z(n3459) );
  CND2XL U3517 ( .A(n1510), .B(n1493), .Z(n3460) );
  CND3X1 U3518 ( .A(n3458), .B(n3460), .C(n3459), .Z(n1486) );
  CND3XL U3519 ( .A(n3802), .B(n3803), .C(n3804), .Z(n3461) );
  CND3XL U3520 ( .A(n3802), .B(n3803), .C(n3804), .Z(n3462) );
  CND3XL U3521 ( .A(n3802), .B(n3803), .C(n3804), .Z(n1518) );
  CENX1 U3522 ( .A(n3463), .B(n1953), .Z(n1523) );
  CND2X2 U3523 ( .A(n1220), .B(n3465), .Z(n3466) );
  CND2XL U3524 ( .A(n3091), .B(n3464), .Z(n3467) );
  CIVXL U3525 ( .A(n1220), .Z(n3464) );
  CIVX1 U3526 ( .A(n3091), .Z(n3465) );
  COND1XL U3527 ( .A(n392), .B(n365), .C(n366), .Z(n3468) );
  CND2X1 U3528 ( .A(a[10]), .B(n3470), .Z(n3471) );
  CND2X1 U3529 ( .A(n3469), .B(net18816), .Z(n3472) );
  CND2X2 U3530 ( .A(n3471), .B(n3472), .Z(net18953) );
  CIVXL U3531 ( .A(a[10]), .Z(n3469) );
  CIVX1 U3532 ( .A(net18816), .Z(n3470) );
  CND3X2 U3533 ( .A(n3782), .B(n3783), .C(n3784), .Z(n1110) );
  CND2X1 U3534 ( .A(n1110), .B(n1112), .Z(n4105) );
  CND2XL U3535 ( .A(n1145), .B(n1168), .Z(n3473) );
  CND2X1 U3536 ( .A(n1145), .B(n1147), .Z(n3474) );
  CND3X1 U3537 ( .A(n3473), .B(n3474), .C(n3475), .Z(n1138) );
  CND2X1 U3538 ( .A(n3555), .B(n3556), .Z(n1145) );
  CND2XL U3539 ( .A(n3775), .B(n1151), .Z(n3555) );
  CENX1 U3540 ( .A(n1176), .B(n1153), .Z(n3775) );
  CND2X2 U3541 ( .A(n1249), .B(n3477), .Z(n3478) );
  CND2X1 U3542 ( .A(n3476), .B(n1276), .Z(n3479) );
  CND2X2 U3543 ( .A(n3478), .B(n3479), .Z(n3830) );
  CIVXL U3544 ( .A(n1249), .Z(n3476) );
  CIVX1 U3545 ( .A(n1276), .Z(n3477) );
  CND3X1 U3546 ( .A(n4219), .B(n4218), .C(n4217), .Z(n1276) );
  CND2X2 U3547 ( .A(n3906), .B(n3905), .Z(n3908) );
  CNR2X2 U3548 ( .A(n3241), .B(n594), .Z(n576) );
  CNIVX2 U3549 ( .A(n21), .Z(n3543) );
  CNIVX2 U3550 ( .A(n21), .Z(n3998) );
  COND2X1 U3551 ( .A(n4002), .B(n2678), .C(net19508), .D(n2677), .Z(n2151) );
  CND3X2 U3552 ( .A(n3523), .B(n3524), .C(n3525), .Z(n1064) );
  CND2X1 U3553 ( .A(n1092), .B(n1094), .Z(n3524) );
  CND2XL U3554 ( .A(n2825), .B(n3678), .Z(n3593) );
  CIVXL U3555 ( .A(n3049), .Z(n779) );
  CNIVX4 U3556 ( .A(n2177), .Z(n3687) );
  COND2X1 U3557 ( .A(net18742), .B(n2704), .C(net16772), .D(n2703), .Z(n2177)
         );
  CAOR1XL U3558 ( .A(n3722), .B(n4260), .C(n2252), .Z(n1740) );
  COND2XL U3559 ( .A(n4260), .B(n2256), .C(n3577), .D(n2255), .Z(n1742) );
  COND2XL U3560 ( .A(n4260), .B(n2262), .C(n3576), .D(n2261), .Z(n1748) );
  COAN1X1 U3561 ( .A(n458), .B(n448), .C(n449), .Z(n3982) );
  CND2X1 U3562 ( .A(n1083), .B(n1106), .Z(n494) );
  CIVX3 U3563 ( .A(net18254), .Z(net16802) );
  CENX1 U3564 ( .A(n2802), .B(n4291), .Z(n2373) );
  COND2XL U3565 ( .A(n3877), .B(n2607), .C(n3839), .D(n2606), .Z(n2080) );
  CENXL U3566 ( .A(n4334), .B(net16063), .Z(n2594) );
  CENXL U3567 ( .A(n4329), .B(net16063), .Z(n2600) );
  CEO3X2 U3568 ( .A(n1753), .B(n1812), .C(n1959), .Z(n919) );
  CND2XL U3569 ( .A(n1753), .B(n1959), .Z(n3483) );
  CND2XL U3570 ( .A(n1753), .B(n1812), .Z(n3484) );
  CND2XL U3571 ( .A(n1959), .B(n1812), .Z(n3485) );
  CND3X1 U3572 ( .A(n3483), .B(n3484), .C(n3485), .Z(n918) );
  CFA1X1 U3573 ( .A(n1197), .B(n1195), .CI(n1222), .CO(n1190), .S(n1191) );
  CND3X2 U3574 ( .A(n3765), .B(n3766), .C(n3767), .Z(n1314) );
  CND3X2 U3575 ( .A(n4304), .B(n4303), .C(n4302), .Z(n1256) );
  CIVX2 U3576 ( .A(net16759), .Z(n3486) );
  CIVX2 U3577 ( .A(net16759), .Z(n3487) );
  CIVXL U3578 ( .A(net16759), .Z(net16027) );
  COR2XL U3579 ( .A(n2521), .B(net19518), .Z(n3508) );
  CEO3X1 U3580 ( .A(n2168), .B(n2137), .C(n2075), .Z(n1517) );
  CND2XL U3581 ( .A(n2168), .B(n2075), .Z(n3491) );
  CND2XL U3582 ( .A(n2168), .B(n2137), .Z(n3492) );
  CND2X1 U3583 ( .A(n2075), .B(n2137), .Z(n3493) );
  CND3X1 U3584 ( .A(n3491), .B(n3492), .C(n3493), .Z(n1516) );
  COND2X1 U3585 ( .A(n3877), .B(n2602), .C(n3839), .D(n2601), .Z(n2075) );
  CND2X1 U3586 ( .A(n1216), .B(n1191), .Z(n3496) );
  CND2X2 U3587 ( .A(n3494), .B(n3495), .Z(n3497) );
  CND2X2 U3588 ( .A(n3496), .B(n3497), .Z(n4009) );
  CIVX2 U3589 ( .A(n1191), .Z(n3494) );
  CIVX2 U3590 ( .A(n1216), .Z(n3495) );
  CND3X1 U3591 ( .A(n4191), .B(n4192), .C(n4193), .Z(n1216) );
  CEO3XL U3592 ( .A(n2188), .B(n1942), .C(n1767), .Z(n1241) );
  CIVXL U3593 ( .A(n4029), .Z(n3498) );
  CIVXL U3594 ( .A(n3498), .Z(n3499) );
  CIVXL U3595 ( .A(n3528), .Z(n3500) );
  CEOX2 U3596 ( .A(n1433), .B(n1431), .Z(n3501) );
  CEOX2 U3597 ( .A(n3501), .B(n1427), .Z(n1421) );
  CND2X1 U3598 ( .A(n1427), .B(n1431), .Z(n3502) );
  CND2XL U3599 ( .A(n1427), .B(n1433), .Z(n3503) );
  CND2XL U3600 ( .A(n1431), .B(n1433), .Z(n3504) );
  CND3XL U3601 ( .A(n3502), .B(n3503), .C(n3504), .Z(n1420) );
  CND2XL U3602 ( .A(n756), .B(n494), .Z(n174) );
  CND3X1 U3603 ( .A(n4109), .B(n4110), .C(n4111), .Z(n1108) );
  CND2XL U3604 ( .A(n1995), .B(n1818), .Z(n3505) );
  CND2XL U3605 ( .A(n1818), .B(n1936), .Z(n3507) );
  CND3X1 U3606 ( .A(n3505), .B(n3506), .C(n3507), .Z(n1028) );
  COR2XL U3607 ( .A(net16771), .B(n2520), .Z(n3509) );
  CENXL U3608 ( .A(n4337), .B(net16824), .Z(n2521) );
  COND1XL U3609 ( .A(n3269), .B(n3420), .C(n362), .Z(n360) );
  COND2XL U3610 ( .A(n81), .B(n2496), .C(n2495), .D(net19061), .Z(n3510) );
  CND2X1 U3611 ( .A(n1451), .B(n1474), .Z(n3511) );
  CND2X1 U3612 ( .A(n1451), .B(n1476), .Z(n3512) );
  CENX2 U3613 ( .A(n3514), .B(n1293), .Z(n1287) );
  COND2X1 U3614 ( .A(n4003), .B(n2672), .C(net19508), .D(n2671), .Z(n2145) );
  CENX1 U3615 ( .A(n3515), .B(n1075), .Z(n1069) );
  CENX1 U3616 ( .A(n1102), .B(n1077), .Z(n3515) );
  CEOX2 U3617 ( .A(n979), .B(n996), .Z(n3516) );
  CEOX2 U3618 ( .A(n3516), .B(n977), .Z(n975) );
  CND2XL U3619 ( .A(n977), .B(n996), .Z(n3517) );
  CND2X1 U3620 ( .A(n977), .B(n979), .Z(n3518) );
  CND2XL U3621 ( .A(n996), .B(n979), .Z(n3519) );
  CND2X1 U3622 ( .A(n1231), .B(n1256), .Z(n3520) );
  CND2X1 U3623 ( .A(n1256), .B(n1258), .Z(n3521) );
  CND2XL U3624 ( .A(n1231), .B(n1258), .Z(n3522) );
  CND3X1 U3625 ( .A(n3520), .B(n3521), .C(n3522), .Z(n1222) );
  CND2X1 U3626 ( .A(n1092), .B(n1071), .Z(n3523) );
  CENX2 U3627 ( .A(n4346), .B(a[2]), .Z(n3526) );
  CENX2 U3628 ( .A(n4346), .B(a[2]), .Z(net18260) );
  CIVX1 U3629 ( .A(n3634), .Z(n3527) );
  CIVX1 U3630 ( .A(n1167), .Z(n3634) );
  COR2XL U3631 ( .A(n1244), .B(n1215), .Z(n3528) );
  CND2X2 U3632 ( .A(net16091), .B(n3530), .Z(n3531) );
  CND2X2 U3633 ( .A(n3529), .B(a[2]), .Z(n3532) );
  CND2X4 U3634 ( .A(n3531), .B(n3532), .Z(n2826) );
  CIVX4 U3635 ( .A(net16091), .Z(n3529) );
  CIVXL U3636 ( .A(a[2]), .Z(n3530) );
  CDLY1XL U3637 ( .A(n1186), .Z(n3533) );
  CIVXL U3638 ( .A(n3534), .Z(n3535) );
  COND2X2 U3639 ( .A(n90), .B(n2464), .C(n3278), .D(n2463), .Z(n1939) );
  CIVX2 U3640 ( .A(n1266), .Z(n3897) );
  CND2X1 U3641 ( .A(n1177), .B(n1179), .Z(n3536) );
  CND2X1 U3642 ( .A(n1177), .B(n1208), .Z(n3537) );
  CND2X1 U3643 ( .A(n1179), .B(n1208), .Z(n3538) );
  CND3X2 U3644 ( .A(n3536), .B(n3537), .C(n3538), .Z(n1170) );
  CENXL U3645 ( .A(n4333), .B(n4360), .Z(n2298) );
  CENXL U3646 ( .A(n4331), .B(n4360), .Z(n2301) );
  CENXL U3647 ( .A(n4332), .B(n4360), .Z(n2299) );
  CENXL U3648 ( .A(net16558), .B(n4360), .Z(n2300) );
  CND2IXL U3649 ( .B(net16109), .A(n3152), .Z(n2317) );
  CENXL U3650 ( .A(n4330), .B(n4360), .Z(n2302) );
  CENXL U3651 ( .A(n4329), .B(n4360), .Z(n2303) );
  CND2X1 U3652 ( .A(n3539), .B(n3540), .Z(n3542) );
  CND2X2 U3653 ( .A(n3541), .B(n3542), .Z(n2822) );
  CIVXL U3654 ( .A(a[10]), .Z(n3540) );
  COND1X1 U3655 ( .A(n487), .B(n3731), .C(n488), .Z(n486) );
  CND2X1 U3656 ( .A(n1607), .B(n1609), .Z(n3692) );
  CANR1X1 U3657 ( .A(n4276), .B(n4027), .C(n432), .Z(n428) );
  CND2X2 U3658 ( .A(n4133), .B(n4134), .Z(n2003) );
  CENX1 U3659 ( .A(n4035), .B(n2003), .Z(n1267) );
  CND2X1 U3660 ( .A(n1248), .B(n1250), .Z(n4192) );
  CENX1 U3661 ( .A(n1347), .B(n1370), .Z(n3776) );
  CND3X1 U3662 ( .A(n4227), .B(n4228), .C(n4229), .Z(n1370) );
  CND3X2 U3663 ( .A(n3778), .B(n3780), .C(n3779), .Z(n1140) );
  CIVX1 U3664 ( .A(n369), .Z(n744) );
  CND2XL U3665 ( .A(n2013), .B(n1983), .Z(n3803) );
  CENX1 U3666 ( .A(n4326), .B(n4291), .Z(n2374) );
  CEO3X2 U3667 ( .A(n1906), .B(n1966), .C(n1847), .Z(n1053) );
  CND2XL U3668 ( .A(n1906), .B(n1966), .Z(n3545) );
  CND2XL U3669 ( .A(n1906), .B(n1847), .Z(n3546) );
  CND2XL U3670 ( .A(n1966), .B(n1847), .Z(n3547) );
  CND3X1 U3671 ( .A(n3545), .B(n3546), .C(n3547), .Z(n1052) );
  CND2XL U3672 ( .A(n1055), .B(n1057), .Z(n3548) );
  CND2XL U3673 ( .A(n1055), .B(n1053), .Z(n3549) );
  CND2XL U3674 ( .A(n1057), .B(n1053), .Z(n3550) );
  CND3X1 U3675 ( .A(n3548), .B(n3549), .C(n3550), .Z(n1044) );
  CNR2XL U3676 ( .A(net18607), .B(n2491), .Z(n3551) );
  CNR2XL U3677 ( .A(net19061), .B(n2490), .Z(n3552) );
  COR2X1 U3678 ( .A(n3551), .B(n3552), .Z(n1966) );
  CND2X2 U3679 ( .A(n3553), .B(n3554), .Z(n3556) );
  CIVXL U3680 ( .A(n1151), .Z(n3553) );
  CIVX2 U3681 ( .A(n3775), .Z(n3554) );
  CND3X2 U3682 ( .A(n3684), .B(n3685), .C(n3686), .Z(n1416) );
  CEO3X1 U3683 ( .A(n1506), .B(n1487), .C(n1485), .Z(n1483) );
  CND2XL U3684 ( .A(n1506), .B(n1485), .Z(n3557) );
  CND2XL U3685 ( .A(n1506), .B(n1487), .Z(n3558) );
  CND2X1 U3686 ( .A(n1485), .B(n1487), .Z(n3559) );
  CND3XL U3687 ( .A(n3557), .B(n3558), .C(n3559), .Z(n1482) );
  CEOX2 U3688 ( .A(n1511), .B(n1513), .Z(n3560) );
  CEOX1 U3689 ( .A(n3560), .B(n1528), .Z(n1507) );
  CND2X1 U3690 ( .A(n1528), .B(n1513), .Z(n3561) );
  CND2X1 U3691 ( .A(n1528), .B(n1511), .Z(n3562) );
  CND2XL U3692 ( .A(n1513), .B(n1511), .Z(n3563) );
  CND3X1 U3693 ( .A(n3561), .B(n3562), .C(n3563), .Z(n1506) );
  CND2X1 U3694 ( .A(n3760), .B(n3761), .Z(n1485) );
  CIVXL U3695 ( .A(n1342), .Z(n3564) );
  CIVXL U3696 ( .A(n3564), .Z(n3565) );
  CIVX4 U3697 ( .A(n4354), .Z(n3943) );
  CIVXL U3698 ( .A(n1534), .Z(n3566) );
  CIVX1 U3699 ( .A(n3566), .Z(n3567) );
  CIVXL U3700 ( .A(n1391), .Z(n3568) );
  CIVXL U3701 ( .A(n3568), .Z(n3569) );
  CND2IXL U3702 ( .B(net16109), .A(net18643), .Z(n2548) );
  COR2X1 U3703 ( .A(n2540), .B(net18670), .Z(n3805) );
  CIVX8 U3704 ( .A(n4293), .Z(n4294) );
  CIVX4 U3705 ( .A(n4293), .Z(n3576) );
  CND2X2 U3706 ( .A(n2825), .B(n24), .Z(net18742) );
  CIVX4 U3707 ( .A(n75), .Z(n3986) );
  COR2X1 U3708 ( .A(n2530), .B(n3415), .Z(n4133) );
  CEOX2 U3709 ( .A(n3952), .B(n1263), .Z(n1255) );
  COND1X1 U3710 ( .A(n710), .B(n708), .C(n709), .Z(n707) );
  CANR1X1 U3711 ( .A(n4278), .B(n4284), .C(n712), .Z(n710) );
  COND1X1 U3712 ( .A(n724), .B(n722), .C(n723), .Z(n721) );
  CND2X1 U3713 ( .A(n970), .B(n3571), .Z(n3572) );
  CND2X1 U3714 ( .A(n3570), .B(n968), .Z(n3573) );
  CND2X2 U3715 ( .A(n3572), .B(n3573), .Z(n3737) );
  COND2XL U3716 ( .A(n3877), .B(n2611), .C(n3839), .D(n2610), .Z(n2084) );
  CND2XL U3717 ( .A(n2083), .B(n2021), .Z(n3923) );
  CFA1X1 U3718 ( .A(n1991), .B(n1755), .CI(n1842), .CO(n952), .S(n953) );
  COND1X2 U3719 ( .A(n3716), .B(n334), .C(n4273), .Z(n286) );
  COND2X1 U3720 ( .A(n3606), .B(n2325), .C(net16801), .D(n2324), .Z(n1808) );
  CND2X2 U3721 ( .A(n2814), .B(net16800), .Z(n126) );
  CND2XL U3722 ( .A(n1473), .B(n1492), .Z(n3812) );
  CEOX2 U3723 ( .A(n3843), .B(n1017), .Z(n1015) );
  CENXL U3724 ( .A(n2808), .B(net15995), .Z(n3575) );
  CND2X1 U3725 ( .A(n3120), .B(n1466), .Z(n3578) );
  CND2X1 U3726 ( .A(n1464), .B(n1443), .Z(n3579) );
  CND2XL U3727 ( .A(n1466), .B(n1443), .Z(n3580) );
  CND3X2 U3728 ( .A(n3578), .B(n3579), .C(n3580), .Z(n1438) );
  CND3X1 U3729 ( .A(n3812), .B(n3813), .C(n3814), .Z(n1466) );
  CEO3X2 U3730 ( .A(n1472), .B(n1470), .C(n1449), .Z(n1443) );
  CND2XL U3731 ( .A(n2106), .B(n1953), .Z(n3581) );
  CND2X1 U3732 ( .A(n1953), .B(n1894), .Z(n3582) );
  CND2XL U3733 ( .A(n2106), .B(n1894), .Z(n3583) );
  CND2X2 U3734 ( .A(n4089), .B(n1544), .Z(n628) );
  CEO3X2 U3735 ( .A(n1166), .B(n1143), .C(n1141), .Z(n1137) );
  CND2X1 U3736 ( .A(n1166), .B(n1141), .Z(n3584) );
  CND2X1 U3737 ( .A(n1141), .B(n1143), .Z(n3586) );
  CND3X2 U3738 ( .A(n3584), .B(n3585), .C(n3586), .Z(n1136) );
  CEO3X2 U3739 ( .A(n1174), .B(n1170), .C(n1172), .Z(n1141) );
  CND2XL U3740 ( .A(n1136), .B(n1113), .Z(n4110) );
  CNIVX8 U3741 ( .A(n111), .Z(n3704) );
  CIVXL U3742 ( .A(n4044), .Z(n1243) );
  CHA1X1 U3743 ( .A(n2117), .B(n2086), .CO(n1682), .S(n1683) );
  COND2X1 U3744 ( .A(n45), .B(n2644), .C(n4017), .D(n2643), .Z(n2117) );
  CND2X1 U3745 ( .A(n878), .B(n867), .Z(n370) );
  CND2X1 U3746 ( .A(n2013), .B(n2199), .Z(n3802) );
  CND2XL U3747 ( .A(n1161), .B(n1163), .Z(n4164) );
  CENX2 U3748 ( .A(n1192), .B(n1165), .Z(n3640) );
  CNIVX4 U3749 ( .A(n4359), .Z(n4251) );
  CND3X2 U3750 ( .A(n3831), .B(n3832), .C(n3833), .Z(n1244) );
  CND2XL U3751 ( .A(n1820), .B(n1761), .Z(n3587) );
  CND3X1 U3752 ( .A(n3587), .B(n3588), .C(n3589), .Z(n1074) );
  CND2XL U3753 ( .A(n1077), .B(n1102), .Z(n3590) );
  CND2XL U3754 ( .A(n1102), .B(n1075), .Z(n3591) );
  CND2XL U3755 ( .A(n1077), .B(n1075), .Z(n3592) );
  CND3X1 U3756 ( .A(n3590), .B(n3592), .C(n3591), .Z(n1068) );
  CND2X1 U3757 ( .A(n2825), .B(n3678), .Z(n27) );
  CIVX1 U3758 ( .A(n460), .Z(n462) );
  CEOX2 U3759 ( .A(n2140), .B(n2171), .Z(n3594) );
  CEOX2 U3760 ( .A(n3594), .B(n2047), .Z(n1573) );
  CND2XL U3761 ( .A(n2047), .B(n2171), .Z(n3595) );
  CND2X1 U3762 ( .A(n2047), .B(n2140), .Z(n3596) );
  CND2XL U3763 ( .A(n2171), .B(n2140), .Z(n3597) );
  CND3X1 U3764 ( .A(n3595), .B(n3596), .C(n3597), .Z(n1572) );
  COR2XL U3765 ( .A(net19500), .B(n2573), .Z(n4086) );
  COND2X2 U3766 ( .A(n2409), .B(net19122), .C(net16839), .D(n2408), .Z(n1887)
         );
  CND2X1 U3767 ( .A(a[10]), .B(net18816), .Z(n3600) );
  CND2X2 U3768 ( .A(n3598), .B(n3599), .Z(n3601) );
  CND2X4 U3769 ( .A(n3600), .B(n3601), .Z(net16658) );
  CIVX1 U3770 ( .A(a[10]), .Z(n3598) );
  CIVX2 U3771 ( .A(net18816), .Z(n3599) );
  CIVX1 U3772 ( .A(net16658), .Z(net18736) );
  CIVX8 U3773 ( .A(net16658), .Z(n3839) );
  CENX1 U3774 ( .A(n4337), .B(n4255), .Z(n2653) );
  CENX2 U3775 ( .A(net16570), .B(net16850), .Z(n2471) );
  CNIVX2 U3776 ( .A(n1517), .Z(n3603) );
  CIVXL U3777 ( .A(n1084), .Z(n3604) );
  CIVXL U3778 ( .A(n3604), .Z(n3605) );
  CND2X2 U3779 ( .A(n2814), .B(net16800), .Z(n3606) );
  CND2X2 U3780 ( .A(n2814), .B(net16800), .Z(n3607) );
  CND3X1 U3781 ( .A(n4311), .B(n4312), .C(n4313), .Z(n1436) );
  CEOX1 U3782 ( .A(n3652), .B(n2050), .Z(n1625) );
  CNR2IX1 U3783 ( .B(net16109), .A(net19060), .Z(n1989) );
  CENX2 U3784 ( .A(n1219), .B(n1246), .Z(n4031) );
  CND2X2 U3785 ( .A(n3641), .B(n1419), .Z(n3644) );
  CND2X2 U3786 ( .A(n1447), .B(n1468), .Z(n4118) );
  CNIVX2 U3787 ( .A(n2170), .Z(n3608) );
  CNR2X1 U3788 ( .A(n879), .B(n892), .Z(n378) );
  CIVXL U3789 ( .A(n379), .Z(n377) );
  CND3X1 U3790 ( .A(n4230), .B(n4231), .C(n4232), .Z(n1376) );
  CND2X1 U3791 ( .A(n1421), .B(n1423), .Z(n3684) );
  CND2XL U3792 ( .A(n1061), .B(n1063), .Z(n3967) );
  CIVX1 U3793 ( .A(n4169), .Z(n4093) );
  CENX2 U3794 ( .A(n1137), .B(n1160), .Z(n4272) );
  CND2XL U3795 ( .A(n3117), .B(n583), .Z(n185) );
  COND2X1 U3796 ( .A(net18592), .B(n2465), .C(n3277), .D(n2464), .Z(n1940) );
  CND2X2 U3797 ( .A(n1425), .B(n3610), .Z(n3611) );
  CND2X1 U3798 ( .A(n3609), .B(n1423), .Z(n3612) );
  CND2X2 U3799 ( .A(n3611), .B(n3612), .Z(n3683) );
  CIVXL U3800 ( .A(n1425), .Z(n3609) );
  COND1XL U3801 ( .A(n224), .B(net19531), .C(n225), .Z(n3613) );
  CND2X2 U3802 ( .A(n4125), .B(n4126), .Z(n1277) );
  COND2X2 U3803 ( .A(net18593), .B(n2471), .C(n3277), .D(n2470), .Z(n1946) );
  CIVX1 U3804 ( .A(n3616), .Z(n3617) );
  CENX2 U3805 ( .A(n4334), .B(n4255), .Z(n2660) );
  CIVXL U3806 ( .A(n3107), .Z(n3618) );
  CIVX1 U3807 ( .A(n3618), .Z(n3619) );
  COR2X2 U3808 ( .A(n1483), .B(n1504), .Z(n3621) );
  CND3X1 U3809 ( .A(n3973), .B(n3974), .C(n3975), .Z(n1504) );
  CENX1 U3810 ( .A(n4328), .B(n4000), .Z(n3873) );
  CIVXL U3811 ( .A(n3411), .Z(n3622) );
  CNR2XL U3812 ( .A(n440), .B(n416), .Z(n3623) );
  CNR2XL U3813 ( .A(n440), .B(n416), .Z(n414) );
  CIVX2 U3814 ( .A(n438), .Z(n440) );
  COND2X1 U3815 ( .A(n3026), .B(n2533), .C(net16771), .D(n2532), .Z(n2006) );
  CENX2 U3816 ( .A(a[12]), .B(net19047), .Z(n3624) );
  CIVX4 U3817 ( .A(n3624), .Z(net19500) );
  CENXL U3818 ( .A(n3406), .B(n3764), .Z(n3625) );
  CANR1X1 U3819 ( .A(n4275), .B(n356), .C(n349), .Z(n345) );
  CANR1X1 U3820 ( .A(n331), .B(n356), .C(n332), .Z(n330) );
  CANR1X1 U3821 ( .A(n320), .B(n356), .C(n323), .Z(n319) );
  CANR1X1 U3822 ( .A(n283), .B(n356), .C(n286), .Z(n282) );
  CANR1X1 U3823 ( .A(n233), .B(n356), .C(n236), .Z(n232) );
  CAN2XL U3824 ( .A(n739), .B(n3626), .Z(n3627) );
  CIVX1 U3825 ( .A(n309), .Z(n3626) );
  CND2XL U3826 ( .A(n355), .B(n3626), .Z(n3628) );
  CIVX3 U3827 ( .A(n353), .Z(n355) );
  CND2X1 U3828 ( .A(n320), .B(n3713), .Z(n309) );
  CEO3X2 U3829 ( .A(n1282), .B(n1255), .C(n3097), .Z(n1249) );
  CND2X1 U3830 ( .A(n1282), .B(n1255), .Z(n3630) );
  CND2XL U3831 ( .A(n1248), .B(n1221), .Z(n4191) );
  CIVXL U3832 ( .A(n308), .Z(n306) );
  CIVXL U3833 ( .A(n260), .Z(n258) );
  COND2XL U3834 ( .A(n126), .B(n2339), .C(net16802), .D(n2338), .Z(n1822) );
  CENXL U3835 ( .A(n2808), .B(net15995), .Z(n2346) );
  CND2X1 U3836 ( .A(n1364), .B(n1339), .Z(n3808) );
  CND2XL U3837 ( .A(n1419), .B(n1442), .Z(n3837) );
  COND2X1 U3838 ( .A(net18607), .B(n2510), .C(n78), .D(n2509), .Z(n1984) );
  COND1XL U3839 ( .A(n224), .B(net19530), .C(n225), .Z(n223) );
  CIVXL U3840 ( .A(n4027), .Z(n3632) );
  CENX1 U3841 ( .A(n4335), .B(n4255), .Z(n2655) );
  CIVX2 U3842 ( .A(n1163), .Z(n4097) );
  CFA1X1 U3843 ( .A(n2054), .B(n2178), .CI(n2116), .CO(n1672), .S(n1673) );
  CNR2IX1 U3844 ( .B(net16109), .A(net19151), .Z(n2054) );
  CENX1 U3845 ( .A(n4325), .B(net16844), .Z(n2705) );
  CIVXL U3846 ( .A(n1998), .Z(n4051) );
  CNR2X2 U3847 ( .A(n1107), .B(n1132), .Z(n504) );
  CNR2XL U3848 ( .A(n1107), .B(n1132), .Z(n3660) );
  CIVXL U3849 ( .A(n4011), .Z(n3638) );
  CND2X1 U3850 ( .A(n3835), .B(n3642), .Z(n3643) );
  CND2X2 U3851 ( .A(n3644), .B(n3643), .Z(n1415) );
  CIVX2 U3852 ( .A(n3835), .Z(n3641) );
  CIVXL U3853 ( .A(n1419), .Z(n3642) );
  CENX1 U3854 ( .A(n4333), .B(n4253), .Z(n2397) );
  CND2X1 U3855 ( .A(n1247), .B(n1249), .Z(n3832) );
  CEO3X2 U3856 ( .A(n1625), .B(n1621), .C(n1623), .Z(n1617) );
  CND2X1 U3857 ( .A(n1625), .B(n1621), .Z(n3645) );
  CND2X1 U3858 ( .A(n1625), .B(n1623), .Z(n3646) );
  CND2X1 U3859 ( .A(n1621), .B(n1623), .Z(n3647) );
  CND3X2 U3860 ( .A(n3645), .B(n3646), .C(n3647), .Z(n1616) );
  CEOX2 U3861 ( .A(n1616), .B(n3648), .Z(n1599) );
  CND2XL U3862 ( .A(n1605), .B(n1603), .Z(n3649) );
  CND2X1 U3863 ( .A(n1605), .B(n1616), .Z(n3650) );
  CND2XL U3864 ( .A(n1603), .B(n1616), .Z(n3651) );
  CND3X1 U3865 ( .A(n3649), .B(n3650), .C(n3651), .Z(n1598) );
  CEOX1 U3866 ( .A(n2143), .B(n1989), .Z(n3652) );
  CND2XL U3867 ( .A(n2050), .B(n1989), .Z(n3653) );
  CND2X1 U3868 ( .A(n2050), .B(n2143), .Z(n3654) );
  CND2XL U3869 ( .A(n1989), .B(n2143), .Z(n3655) );
  CND3X1 U3870 ( .A(n3653), .B(n3654), .C(n3655), .Z(n1624) );
  CND2IX2 U3871 ( .B(n4097), .A(n4098), .Z(n4099) );
  CAN2X1 U3872 ( .A(n735), .B(n3656), .Z(n3657) );
  CIVX2 U3873 ( .A(n261), .Z(n3656) );
  CND2X1 U3874 ( .A(n355), .B(n3656), .Z(n3658) );
  CND2X1 U3875 ( .A(n3627), .B(n355), .Z(n298) );
  CND2X1 U3876 ( .A(n3657), .B(n355), .Z(n248) );
  CENXL U3877 ( .A(n4323), .B(net16093), .Z(n2740) );
  CENXL U3878 ( .A(n4324), .B(net16093), .Z(n2739) );
  CENXL U3879 ( .A(n2808), .B(net16093), .Z(n2742) );
  CENXL U3880 ( .A(n2810), .B(net16093), .Z(n2744) );
  CENXL U3881 ( .A(n2802), .B(net16093), .Z(n2736) );
  CENXL U3882 ( .A(n4322), .B(net16093), .Z(n2741) );
  CENXL U3883 ( .A(n4327), .B(net16093), .Z(n2734) );
  CENXL U3884 ( .A(net16570), .B(net16093), .Z(n2735) );
  CENXL U3885 ( .A(n4321), .B(net16093), .Z(n2743) );
  CENXL U3886 ( .A(n4326), .B(net16093), .Z(n2737) );
  CENXL U3887 ( .A(n4342), .B(net16093), .Z(n2714) );
  CENXL U3888 ( .A(n4328), .B(net16093), .Z(n2733) );
  CENXL U3889 ( .A(n4329), .B(net16093), .Z(n2732) );
  CENXL U3890 ( .A(net16558), .B(net16093), .Z(n2729) );
  CENXL U3891 ( .A(n4333), .B(net16093), .Z(n2727) );
  CND2X2 U3892 ( .A(a[6]), .B(n3663), .Z(n3664) );
  CND2X1 U3893 ( .A(n4348), .B(n3662), .Z(n3665) );
  CND2X2 U3894 ( .A(n3664), .B(n3665), .Z(n4172) );
  CIVX2 U3895 ( .A(n4348), .Z(n3663) );
  CEOX2 U3896 ( .A(n1567), .B(n1582), .Z(n3666) );
  CEOX2 U3897 ( .A(n1565), .B(n3666), .Z(n1563) );
  CND2XL U3898 ( .A(n1567), .B(n1582), .Z(n3669) );
  CND2XL U3899 ( .A(n3261), .B(n1058), .Z(n3670) );
  CEOX2 U3900 ( .A(n1536), .B(n1523), .Z(n3671) );
  CEOX2 U3901 ( .A(n3671), .B(n3603), .Z(n1513) );
  CND2X1 U3902 ( .A(n1517), .B(n1523), .Z(n3672) );
  CND2X1 U3903 ( .A(n1517), .B(n1536), .Z(n3673) );
  CND2XL U3904 ( .A(n1523), .B(n1536), .Z(n3674) );
  CND3X1 U3905 ( .A(n3672), .B(n3673), .C(n3674), .Z(n1512) );
  CND2XL U3906 ( .A(net16544), .B(n4000), .Z(n3676) );
  CND2X1 U3907 ( .A(n3675), .B(n3880), .Z(n3677) );
  CND2X1 U3908 ( .A(n3676), .B(n3677), .Z(n4030) );
  CIVXL U3909 ( .A(net16544), .Z(n3675) );
  CENX2 U3910 ( .A(a[4]), .B(n3219), .Z(n3678) );
  CENX2 U3911 ( .A(a[4]), .B(n3219), .Z(n24) );
  CIVX1 U3912 ( .A(n84), .Z(n3985) );
  CENXL U3913 ( .A(n642), .B(n193), .Z(product[19]) );
  CENX1 U3914 ( .A(n4332), .B(n4000), .Z(n2563) );
  CENX2 U3915 ( .A(n1491), .B(n1489), .Z(n3934) );
  CND2X1 U3916 ( .A(n1494), .B(n3680), .Z(n3681) );
  CND2X1 U3917 ( .A(n3679), .B(n1492), .Z(n3682) );
  CND2X2 U3918 ( .A(n3681), .B(n3682), .Z(n3811) );
  CIVXL U3919 ( .A(n1494), .Z(n3679) );
  COND2X1 U3920 ( .A(n3092), .B(n2623), .C(net16793), .D(n2622), .Z(n2096) );
  COND2X1 U3921 ( .A(n3092), .B(n2618), .C(net16793), .D(n2617), .Z(n2091) );
  COND2X1 U3922 ( .A(n18), .B(n2738), .C(net16816), .D(n2737), .Z(n2211) );
  CND2X1 U3923 ( .A(n1421), .B(n1425), .Z(n3685) );
  CND2XL U3924 ( .A(n1423), .B(n1425), .Z(n3686) );
  CENXL U3925 ( .A(n4332), .B(net16067), .Z(n2629) );
  CENXL U3926 ( .A(net16548), .B(net16067), .Z(n2625) );
  CND2XL U3927 ( .A(n1439), .B(n1441), .Z(n4312) );
  CEO3X1 U3928 ( .A(n1638), .B(n1634), .C(n1636), .Z(n1619) );
  CND2XL U3929 ( .A(n3083), .B(n1634), .Z(n3688) );
  CND2XL U3930 ( .A(n3083), .B(n1636), .Z(n3689) );
  CND2XL U3931 ( .A(n1634), .B(n1636), .Z(n3690) );
  CND3X1 U3932 ( .A(n3688), .B(n3689), .C(n3690), .Z(n1618) );
  CEOX2 U3933 ( .A(n1607), .B(n1609), .Z(n3691) );
  CEOX1 U3934 ( .A(n3691), .B(n3048), .Z(n1601) );
  CND2X1 U3935 ( .A(n1607), .B(n1618), .Z(n3693) );
  CND2X1 U3936 ( .A(n1609), .B(n1618), .Z(n3694) );
  CND2X2 U3937 ( .A(n975), .B(n994), .Z(n449) );
  COND2XL U3938 ( .A(n144), .B(n2270), .C(n3576), .D(n2269), .Z(n1756) );
  CENX1 U3939 ( .A(a[24]), .B(n4354), .Z(n4295) );
  CEO3X2 U3940 ( .A(n1521), .B(n1519), .C(n3567), .Z(n1511) );
  CND2XL U3941 ( .A(n1534), .B(n1521), .Z(n3697) );
  CND2XL U3942 ( .A(n1521), .B(n1519), .Z(n3698) );
  CND2XL U3943 ( .A(n1534), .B(n1519), .Z(n3699) );
  CDLY1XL U3944 ( .A(n677), .Z(n3700) );
  CDLY1XL U3945 ( .A(n3576), .Z(n3722) );
  CND2X4 U3946 ( .A(n2812), .B(n4294), .Z(n4261) );
  CND2XL U3947 ( .A(n1469), .B(n1490), .Z(n3701) );
  CND2XL U3948 ( .A(n1469), .B(n1471), .Z(n3702) );
  CND2XL U3949 ( .A(n1490), .B(n1471), .Z(n3703) );
  CNIVXL U3950 ( .A(net19531), .Z(n3705) );
  CIVX2 U3951 ( .A(n111), .Z(n4358) );
  COND1X1 U3952 ( .A(n417), .B(n3420), .C(n3797), .Z(n3823) );
  CND2X1 U3953 ( .A(n1165), .B(n1190), .Z(n3706) );
  CND2X1 U3954 ( .A(n1190), .B(n1192), .Z(n3707) );
  CND2X1 U3955 ( .A(n1165), .B(n1192), .Z(n3708) );
  CND3X2 U3956 ( .A(n3706), .B(n3707), .C(n3708), .Z(n1160) );
  CND2X1 U3957 ( .A(n1135), .B(n1160), .Z(n4296) );
  CENX2 U3958 ( .A(a[0]), .B(n4346), .Z(n2827) );
  CIVX4 U3959 ( .A(n4346), .Z(n4343) );
  COR2X2 U3960 ( .A(net19061), .B(n2506), .Z(n4119) );
  CANR1X1 U3961 ( .A(n3403), .B(n415), .C(n3638), .Z(n395) );
  CIVXL U3962 ( .A(n3309), .Z(n1035) );
  CIVX8 U3963 ( .A(n4263), .Z(n4362) );
  CND2X1 U3964 ( .A(n1575), .B(n1573), .Z(n4081) );
  CNIVX4 U3965 ( .A(n2792), .Z(n4334) );
  CHA1X1 U3966 ( .A(n1727), .B(n1862), .CO(n1458), .S(n1459) );
  CND2X1 U3967 ( .A(n4085), .B(n4086), .Z(n2047) );
  CENX1 U3968 ( .A(n4337), .B(n4344), .Z(n2752) );
  CENX1 U3969 ( .A(n4325), .B(n4253), .Z(n2408) );
  CENX1 U3970 ( .A(n4327), .B(n4292), .Z(n2437) );
  CNIVX4 U3971 ( .A(n2795), .Z(net16558) );
  CNIVX4 U3972 ( .A(n2799), .Z(n4328) );
  CNIVX12 U3973 ( .A(n2794), .Z(n4332) );
  CIVX2 U3974 ( .A(a[16]), .Z(net18609) );
  CNIVX4 U3975 ( .A(n2798), .Z(n4329) );
  CENX1 U3976 ( .A(n4321), .B(n4362), .Z(n2281) );
  CNIVX4 U3977 ( .A(n2796), .Z(n4331) );
  CENX1 U3978 ( .A(n4340), .B(net19089), .Z(n2683) );
  CND3X1 U3979 ( .A(n4202), .B(n4203), .C(n4204), .Z(n1298) );
  CENX1 U3980 ( .A(n4334), .B(net18936), .Z(n2528) );
  CNIVX4 U3981 ( .A(n2787), .Z(n4335) );
  CNIVX4 U3982 ( .A(n2785), .Z(n4337) );
  CNIVX4 U3983 ( .A(n2784), .Z(n4338) );
  CNIVX4 U3984 ( .A(n2783), .Z(n4339) );
  COND2X1 U3985 ( .A(n99), .B(n2428), .C(n3920), .D(n2427), .Z(n1034) );
  CNIVX4 U3986 ( .A(n2805), .Z(n4324) );
  CNIVX4 U3987 ( .A(n2782), .Z(n4340) );
  CIVDX3 U3988 ( .A(n136), .Z0(n4263), .Z1(n4262) );
  CND3X1 U3989 ( .A(n3734), .B(n3735), .C(n3736), .Z(n972) );
  CND2X1 U3990 ( .A(n1590), .B(n1575), .Z(n4079) );
  CND2X1 U3991 ( .A(n1590), .B(n1573), .Z(n4080) );
  CEOX1 U3992 ( .A(n4220), .B(n1409), .Z(n1397) );
  CND3X1 U3993 ( .A(n4242), .B(n4243), .C(n4244), .Z(n1226) );
  CNR2X1 U3994 ( .A(n302), .B(n295), .Z(n293) );
  CND2X1 U3995 ( .A(n293), .B(n3713), .Z(n291) );
  CND2X1 U3996 ( .A(n233), .B(net18421), .Z(n224) );
  CEOX1 U3997 ( .A(n4067), .B(n3127), .Z(n979) );
  CNIVX4 U3998 ( .A(n145), .Z(net16109) );
  CND2X1 U3999 ( .A(n826), .B(n819), .Z(n303) );
  CENX4 U4000 ( .A(a[28]), .B(n3288), .Z(n3709) );
  COR2X1 U4001 ( .A(n265), .B(n241), .Z(n3710) );
  CNIVX1 U4002 ( .A(n1961), .Z(n3712) );
  COR2X1 U4003 ( .A(n827), .B(n834), .Z(n3713) );
  CIVDXL U4004 ( .A(n1725), .Z0(n3714), .Z1(n3715) );
  COR2X1 U4005 ( .A(n291), .B(n324), .Z(n3716) );
  COR2XL U4006 ( .A(n1214), .B(n1187), .Z(n3717) );
  CANR1XL U4007 ( .A(n753), .B(n3602), .C(n467), .Z(n3718) );
  CAN2X1 U4008 ( .A(n3860), .B(n3861), .Z(n3719) );
  CAN2XL U4009 ( .A(n1257), .B(n3853), .Z(n3720) );
  CAN2XL U4010 ( .A(n1259), .B(n3853), .Z(n3721) );
  CNR2X1 U4011 ( .A(n1386), .B(n1361), .Z(n572) );
  COR2XL U4012 ( .A(n2251), .B(n1739), .Z(n3723) );
  CENXL U4013 ( .A(n3724), .B(n619), .Z(product[23]) );
  CAN2XL U4014 ( .A(n3620), .B(n618), .Z(n3724) );
  CENXL U4015 ( .A(n3725), .B(n3731), .Z(product[32]) );
  CAN2XL U4016 ( .A(n3342), .B(n3068), .Z(n3725) );
  CENXL U4017 ( .A(n611), .B(n3726), .Z(product[24]) );
  CAN2XL U4018 ( .A(n770), .B(n4108), .Z(n3726) );
  COND2X1 U4019 ( .A(n3606), .B(n2323), .C(net16801), .D(n2322), .Z(n842) );
  CENXL U4020 ( .A(n486), .B(n173), .Z(product[39]) );
  CENXL U4021 ( .A(n584), .B(n185), .Z(product[27]) );
  CENXL U4022 ( .A(n3727), .B(n560), .Z(product[30]) );
  CAN2XL U4023 ( .A(n3300), .B(n764), .Z(n3727) );
  CENXL U4024 ( .A(n3728), .B(n569), .Z(product[29]) );
  CAN2XL U4025 ( .A(n568), .B(n765), .Z(n3728) );
  CNR2IX1 U4026 ( .B(n3220), .A(n389), .Z(n387) );
  COND2XL U4027 ( .A(n2555), .B(net19168), .C(net19151), .D(n2554), .Z(n2028)
         );
  CIVXL U4028 ( .A(n458), .Z(n456) );
  COND1X1 U4029 ( .A(n611), .B(n594), .C(net19384), .Z(n593) );
  CNIVX4 U4030 ( .A(net19048), .Z(n3729) );
  CNIVX4 U4031 ( .A(net19048), .Z(n3730) );
  CENXL U4032 ( .A(n629), .B(n191), .Z(product[21]) );
  CIVXL U4033 ( .A(n212), .Z(product[63]) );
  CENXL U4034 ( .A(n3732), .B(net19409), .Z(product[40]) );
  CAN2XL U4035 ( .A(n3202), .B(n3670), .Z(n3732) );
  CNR2X1 U4036 ( .A(n440), .B(n385), .Z(n383) );
  CIVXL U4037 ( .A(n383), .Z(n381) );
  CENXL U4038 ( .A(n4335), .B(net18643), .Z(n3733) );
  CIVXL U4039 ( .A(n666), .Z(n664) );
  CND2X1 U4040 ( .A(n779), .B(n666), .Z(n197) );
  CEO3X1 U4041 ( .A(n1756), .B(n992), .C(n3741), .Z(n973) );
  CND2XL U4042 ( .A(n1756), .B(n992), .Z(n3734) );
  CND2XL U4043 ( .A(n3031), .B(n1992), .Z(n3735) );
  CND2XL U4044 ( .A(n992), .B(n1992), .Z(n3736) );
  CND2XL U4045 ( .A(n970), .B(n968), .Z(n3738) );
  CND2XL U4046 ( .A(n970), .B(n972), .Z(n3739) );
  CND3X1 U4047 ( .A(n3738), .B(n3739), .C(n3740), .Z(n946) );
  CNIVX1 U4048 ( .A(n1992), .Z(n3741) );
  COND2XL U4049 ( .A(n2517), .B(net16771), .C(n2518), .D(net19518), .Z(n1992)
         );
  COND2X1 U4050 ( .A(n2580), .B(n3139), .C(net19500), .D(n2579), .Z(n2053) );
  CENX1 U4051 ( .A(n4321), .B(n3729), .Z(n2611) );
  CIVX2 U4052 ( .A(n4176), .Z(n4348) );
  CIVX2 U4053 ( .A(n1188), .Z(n4098) );
  CENXL U4054 ( .A(net16109), .B(net16037), .Z(n2514) );
  CENXL U4055 ( .A(n2802), .B(net16037), .Z(n2505) );
  CENXL U4056 ( .A(n4342), .B(net16037), .Z(n2483) );
  CENXL U4057 ( .A(n4324), .B(net16037), .Z(n2508) );
  CENXL U4058 ( .A(n4323), .B(net16037), .Z(n2509) );
  CENXL U4059 ( .A(n4321), .B(net16037), .Z(n2512) );
  CENXL U4060 ( .A(n4322), .B(net16037), .Z(n2510) );
  CENXL U4061 ( .A(n2808), .B(net16037), .Z(n2511) );
  CENXL U4062 ( .A(n4327), .B(net16037), .Z(n2503) );
  CENXL U4063 ( .A(net16558), .B(net16037), .Z(n2498) );
  CENXL U4064 ( .A(n4332), .B(net16037), .Z(n2497) );
  CND2IXL U4065 ( .B(net16109), .A(net16037), .Z(n2515) );
  CENX1 U4066 ( .A(n4329), .B(net16037), .Z(n2501) );
  CENXL U4067 ( .A(n4326), .B(net16037), .Z(n2506) );
  CENX1 U4068 ( .A(n4328), .B(net16037), .Z(n2502) );
  CENXL U4069 ( .A(n4331), .B(net16850), .Z(n3742) );
  CND2X1 U4070 ( .A(n3743), .B(n1440), .Z(n3746) );
  CND2X2 U4071 ( .A(n3745), .B(n3746), .Z(n3835) );
  CIVX2 U4072 ( .A(n1440), .Z(n3744) );
  CND2XL U4073 ( .A(n4013), .B(n1453), .Z(n3749) );
  CND2X1 U4074 ( .A(n3747), .B(n3748), .Z(n3750) );
  CIVX1 U4075 ( .A(n4013), .Z(n3747) );
  CIVXL U4076 ( .A(n1453), .Z(n3748) );
  CIVXL U4077 ( .A(n1118), .Z(n3751) );
  CIVXL U4078 ( .A(n3751), .Z(n3752) );
  CND2X1 U4079 ( .A(n1015), .B(n1036), .Z(n469) );
  CENX1 U4080 ( .A(n4326), .B(net16059), .Z(n2605) );
  CENX1 U4081 ( .A(n4328), .B(n3730), .Z(n2601) );
  CND2X1 U4082 ( .A(n1390), .B(n1367), .Z(n3753) );
  CND2X1 U4083 ( .A(n1390), .B(n1392), .Z(n3754) );
  CND2XL U4084 ( .A(n1367), .B(n1392), .Z(n3755) );
  CND3X2 U4085 ( .A(n3753), .B(n3754), .C(n3755), .Z(n1362) );
  CIVX4 U4086 ( .A(n3526), .Z(net16816) );
  CIVX8 U4087 ( .A(n4290), .Z(n4291) );
  CIVX4 U4088 ( .A(n4357), .Z(n4290) );
  CENX1 U4089 ( .A(n2810), .B(n4291), .Z(n2381) );
  CND2X1 U4090 ( .A(n3934), .B(n1508), .Z(n3760) );
  CND2X2 U4091 ( .A(n3758), .B(n3759), .Z(n3761) );
  CIVXL U4092 ( .A(n1508), .Z(n3758) );
  CIVX2 U4093 ( .A(n3934), .Z(n3759) );
  CND3X1 U4094 ( .A(n4149), .B(n4150), .C(n4151), .Z(n1508) );
  CIVXL U4095 ( .A(n93), .Z(n4353) );
  CIVX2 U4096 ( .A(n93), .Z(n4264) );
  CENX1 U4097 ( .A(n4334), .B(net16843), .Z(n2693) );
  CENX1 U4098 ( .A(n2802), .B(net18937), .Z(n2538) );
  CENXL U4099 ( .A(net16570), .B(net16037), .Z(n2504) );
  CEO3X1 U4100 ( .A(n1325), .B(n1348), .C(n1323), .Z(n1315) );
  CND2XL U4101 ( .A(n1325), .B(n1323), .Z(n3766) );
  CND2X1 U4102 ( .A(n1348), .B(n1323), .Z(n3767) );
  CEOX2 U4103 ( .A(n1289), .B(n1287), .Z(n3768) );
  CND2X1 U4104 ( .A(n1287), .B(n1289), .Z(n3769) );
  CND2X1 U4105 ( .A(n1289), .B(n1314), .Z(n3770) );
  CND2X1 U4106 ( .A(n1287), .B(n1314), .Z(n3771) );
  CEO3X1 U4107 ( .A(n1945), .B(n1975), .C(n1916), .Z(n1325) );
  CND2XL U4108 ( .A(n1945), .B(n1916), .Z(n3772) );
  CND2XL U4109 ( .A(n1945), .B(n1975), .Z(n3773) );
  CND2XL U4110 ( .A(n1916), .B(n1975), .Z(n3774) );
  CND3X1 U4111 ( .A(n3772), .B(n3773), .C(n3774), .Z(n1324) );
  COND2X1 U4112 ( .A(net18592), .B(n2470), .C(n3278), .D(n2469), .Z(n1945) );
  COND2X1 U4113 ( .A(n54), .B(n2592), .C(n3839), .D(n2591), .Z(n2065) );
  CAOR1XL U4114 ( .A(n3919), .B(n99), .C(n2417), .Z(n1895) );
  COND2X1 U4115 ( .A(net18897), .B(n2443), .C(n3920), .D(n2442), .Z(n1920) );
  COND2X1 U4116 ( .A(net18897), .B(n2432), .C(n3920), .D(n2431), .Z(n1909) );
  CEOXL U4117 ( .A(n1900), .B(n921), .Z(n3792) );
  CEO3X2 U4118 ( .A(n2108), .B(n1985), .C(n1926), .Z(n1561) );
  CND2XL U4119 ( .A(n1926), .B(n2108), .Z(n3918) );
  CFA1XL U4120 ( .A(n890), .B(n1897), .CI(n1809), .CO(n876), .S(n877) );
  CIVX4 U4121 ( .A(n3126), .Z(net19060) );
  CENXL U4122 ( .A(n4336), .B(n4145), .Z(n2555) );
  CENXL U4123 ( .A(n4339), .B(n4349), .Z(n2552) );
  CENX1 U4124 ( .A(n4341), .B(net16843), .Z(n2682) );
  CNR2X2 U4125 ( .A(n511), .B(n504), .Z(n4029) );
  CIVXL U4126 ( .A(n530), .Z(n528) );
  CANR1X1 U4127 ( .A(n359), .B(n3659), .C(n3823), .Z(n3777) );
  CANR1XL U4128 ( .A(n359), .B(n3659), .C(n3823), .Z(net19531) );
  CND2XL U4129 ( .A(n1174), .B(n1170), .Z(n3778) );
  CND2X1 U4130 ( .A(n1174), .B(n1172), .Z(n3779) );
  CEOX2 U4131 ( .A(n1117), .B(n1115), .Z(n3781) );
  CEOX2 U4132 ( .A(n3781), .B(n1140), .Z(n1111) );
  CND2X1 U4133 ( .A(n1117), .B(n1115), .Z(n3782) );
  CND2X1 U4134 ( .A(n1117), .B(n1140), .Z(n3783) );
  CEO3X2 U4135 ( .A(n2063), .B(n2032), .C(n1825), .Z(n1207) );
  CND2XL U4136 ( .A(n2032), .B(n1825), .Z(n3785) );
  CND2XL U4137 ( .A(n2032), .B(n2063), .Z(n3786) );
  CND2XL U4138 ( .A(n1825), .B(n2063), .Z(n3787) );
  CND3X1 U4139 ( .A(n3785), .B(n3786), .C(n3787), .Z(n1206) );
  COND2XL U4140 ( .A(n3607), .B(n2342), .C(net16801), .D(n2341), .Z(n1825) );
  COND2X1 U4141 ( .A(n2398), .B(n4188), .C(net19462), .D(n2397), .Z(n1876) );
  CIVXL U4142 ( .A(n4108), .Z(n3788) );
  CND2X4 U4143 ( .A(n4103), .B(net19269), .Z(n33) );
  CND2X2 U4144 ( .A(n3998), .B(a[6]), .Z(net19269) );
  CANR1X1 U4145 ( .A(net18421), .B(n236), .C(n227), .Z(n225) );
  CIVX2 U4146 ( .A(n48), .Z(net19047) );
  COND2X1 U4147 ( .A(n3092), .B(n2632), .C(net16793), .D(n2631), .Z(n2105) );
  CEO3X2 U4148 ( .A(n1754), .B(n1960), .C(n954), .Z(n937) );
  CND2X1 U4149 ( .A(n1754), .B(n1960), .Z(n3789) );
  CND2X1 U4150 ( .A(n1754), .B(n954), .Z(n3790) );
  CND2X1 U4151 ( .A(n1960), .B(n954), .Z(n3791) );
  CND3X2 U4152 ( .A(n3789), .B(n3790), .C(n3791), .Z(n936) );
  CEOX1 U4153 ( .A(n3792), .B(n936), .Z(n915) );
  CND2X1 U4154 ( .A(n1900), .B(n921), .Z(n3793) );
  CND2X1 U4155 ( .A(n1900), .B(n936), .Z(n3794) );
  CND2X1 U4156 ( .A(n921), .B(n936), .Z(n3795) );
  CND3X2 U4157 ( .A(n3793), .B(n3794), .C(n3795), .Z(n914) );
  CIVX1 U4158 ( .A(n4170), .Z(n3796) );
  CND2X1 U4159 ( .A(n1613), .B(n1626), .Z(n661) );
  CND2XL U4160 ( .A(n3661), .B(n3533), .Z(n3798) );
  CENXL U4161 ( .A(net16544), .B(net16824), .Z(n2524) );
  CENXL U4162 ( .A(n4339), .B(net18643), .Z(n2519) );
  CENXL U4163 ( .A(n4340), .B(net18643), .Z(n2518) );
  CENXL U4164 ( .A(n4338), .B(net18643), .Z(n2520) );
  CIVX1 U4165 ( .A(n1860), .Z(n3799) );
  CIVX2 U4166 ( .A(n3799), .Z(n3800) );
  CEOX1 U4167 ( .A(n1983), .B(n2199), .Z(n3801) );
  CEOX1 U4168 ( .A(n3801), .B(n2013), .Z(n1519) );
  CND2XL U4169 ( .A(n2199), .B(n1983), .Z(n3804) );
  CND2X2 U4170 ( .A(n3805), .B(n3806), .Z(n2013) );
  CHA1XL U4171 ( .A(n2020), .B(n2051), .CO(n1638), .S(n1639) );
  CND2X1 U4172 ( .A(n1364), .B(n1341), .Z(n3809) );
  CND3X2 U4173 ( .A(n3808), .B(n3809), .C(n3810), .Z(n1334) );
  CEOX2 U4174 ( .A(n3811), .B(n1473), .Z(n1467) );
  CND2XL U4175 ( .A(n1492), .B(n1494), .Z(n3814) );
  CENXL U4176 ( .A(n4332), .B(n4259), .Z(n2431) );
  CENXL U4177 ( .A(n4331), .B(n4259), .Z(n2433) );
  CENXL U4178 ( .A(n4329), .B(n4259), .Z(n2435) );
  CENX1 U4179 ( .A(n4333), .B(n4259), .Z(n2430) );
  COND2X1 U4180 ( .A(net18670), .B(n2517), .C(n4144), .D(n2516), .Z(n1991) );
  CND2XL U4181 ( .A(n2010), .B(n1950), .Z(n4198) );
  CENX1 U4182 ( .A(n3865), .B(n3310), .Z(n1083) );
  COND2XL U4183 ( .A(net19417), .B(n2380), .C(n4295), .D(n2379), .Z(n1860) );
  CND3X2 U4184 ( .A(n766), .B(net18739), .C(n765), .Z(n547) );
  CIVX1 U4185 ( .A(n3544), .Z(n765) );
  CND2X1 U4186 ( .A(net16548), .B(net16843), .Z(n3817) );
  CND2X2 U4187 ( .A(n3815), .B(n3816), .Z(n3818) );
  CND2X2 U4188 ( .A(n3817), .B(n3818), .Z(n2691) );
  CIVXL U4189 ( .A(net16548), .Z(n3815) );
  CIVX1 U4190 ( .A(net16843), .Z(n3816) );
  CNIVX4 U4191 ( .A(n2790), .Z(net16548) );
  COND2X1 U4192 ( .A(n3024), .B(n2692), .C(net16772), .D(n2691), .Z(n2165) );
  CND2XL U4193 ( .A(n4306), .B(n4330), .Z(n3820) );
  CND2X1 U4194 ( .A(n3820), .B(n3821), .Z(n2566) );
  CIVXL U4195 ( .A(n4330), .Z(n3819) );
  CNIVX4 U4196 ( .A(n2797), .Z(n4330) );
  CIVX1 U4197 ( .A(n582), .Z(n767) );
  CENX1 U4198 ( .A(n4336), .B(n4255), .Z(n2654) );
  COND2XL U4199 ( .A(net18670), .B(n2524), .C(n4144), .D(n3733), .Z(n1998) );
  COND1X1 U4200 ( .A(n484), .B(n494), .C(n485), .Z(n483) );
  CENX2 U4201 ( .A(n4170), .B(a[28]), .Z(n2813) );
  CENX1 U4202 ( .A(n4325), .B(n4360), .Z(n2309) );
  CENX1 U4203 ( .A(n2808), .B(n4291), .Z(n2379) );
  CENX1 U4204 ( .A(n4322), .B(n4291), .Z(n2378) );
  CNR2XL U4205 ( .A(n522), .B(n529), .Z(n3824) );
  CNR2XL U4206 ( .A(n522), .B(n529), .Z(n3825) );
  CND2X1 U4207 ( .A(n3639), .B(n1218), .Z(n3827) );
  CND2X2 U4208 ( .A(n3637), .B(n3826), .Z(n3828) );
  CND2X2 U4209 ( .A(n3827), .B(n3828), .Z(n1189) );
  CIVXL U4210 ( .A(n1218), .Z(n3826) );
  CNR2XL U4211 ( .A(n522), .B(n529), .Z(n520) );
  COND1X1 U4212 ( .A(n4088), .B(n540), .C(n541), .Z(n3829) );
  CND2X1 U4213 ( .A(n1247), .B(n1276), .Z(n3831) );
  CND2XL U4214 ( .A(n1276), .B(n1249), .Z(n3833) );
  COND1X1 U4215 ( .A(n4088), .B(n540), .C(n541), .Z(n535) );
  CNR2X1 U4216 ( .A(n1245), .B(n1274), .Z(n543) );
  CANR1X1 U4217 ( .A(n482), .B(n499), .C(n483), .Z(n3834) );
  CANR1X1 U4218 ( .A(n482), .B(n499), .C(n483), .Z(n481) );
  CENXL U4219 ( .A(n4341), .B(n4251), .Z(n2286) );
  CENXL U4220 ( .A(n4340), .B(n4251), .Z(n2287) );
  CENXL U4221 ( .A(n4339), .B(n4251), .Z(n2288) );
  CENXL U4222 ( .A(n4336), .B(n4251), .Z(n2291) );
  CENXL U4223 ( .A(n4335), .B(n4251), .Z(n2292) );
  CENXL U4224 ( .A(n4338), .B(n4251), .Z(n2289) );
  CENXL U4225 ( .A(n4337), .B(n4251), .Z(n2290) );
  CENXL U4226 ( .A(net16544), .B(n4251), .Z(n2293) );
  CENXL U4227 ( .A(n2789), .B(n4251), .Z(n2294) );
  CND2XL U4228 ( .A(n1419), .B(n1440), .Z(n3836) );
  CND2XL U4229 ( .A(n1440), .B(n1442), .Z(n3838) );
  CND3X1 U4230 ( .A(n3836), .B(n3837), .C(n3838), .Z(n1414) );
  CND2XL U4231 ( .A(n3569), .B(n1414), .Z(n4316) );
  CND2XL U4232 ( .A(n1151), .B(n1153), .Z(n3840) );
  CND2X1 U4233 ( .A(n1151), .B(n1176), .Z(n3841) );
  CND2XL U4234 ( .A(n1153), .B(n1176), .Z(n3842) );
  CND3X1 U4235 ( .A(n3840), .B(n3841), .C(n3842), .Z(n1144) );
  CEOX2 U4236 ( .A(n1019), .B(n1038), .Z(n3843) );
  CND2XL U4237 ( .A(n1017), .B(n1038), .Z(n3844) );
  CND2X1 U4238 ( .A(n1017), .B(n1019), .Z(n3845) );
  CND2XL U4239 ( .A(n1038), .B(n1019), .Z(n3846) );
  CND3XL U4240 ( .A(n3844), .B(n3845), .C(n3846), .Z(n1014) );
  CEOX1 U4241 ( .A(n3847), .B(n1223), .Z(n1219) );
  CND2X1 U4242 ( .A(n1223), .B(n1252), .Z(n3848) );
  CND2X2 U4243 ( .A(n3130), .B(n3851), .Z(n1251) );
  CND2X1 U4244 ( .A(n3852), .B(n3719), .Z(n1250) );
  CIVX2 U4245 ( .A(n1284), .Z(n3853) );
  CIVXL U4246 ( .A(n1257), .Z(n3855) );
  CND2X1 U4247 ( .A(n3854), .B(n3720), .Z(n3856) );
  CND2X1 U4248 ( .A(n3855), .B(n3721), .Z(n3857) );
  CND2X1 U4249 ( .A(n3855), .B(n3863), .Z(n3858) );
  CND2XL U4250 ( .A(n1259), .B(n1284), .Z(n3860) );
  CND2XL U4251 ( .A(n1257), .B(n1284), .Z(n3861) );
  CND2XL U4252 ( .A(n1257), .B(n1259), .Z(n3852) );
  CND2X1 U4253 ( .A(n3858), .B(n3859), .Z(n3862) );
  CIVX2 U4254 ( .A(n3862), .Z(n3851) );
  CNR2XL U4255 ( .A(n3853), .B(n1259), .Z(n3863) );
  CND2XL U4256 ( .A(n1257), .B(n3864), .Z(n3859) );
  COND2XL U4257 ( .A(n3116), .B(n2295), .C(n3709), .D(n2294), .Z(n1780) );
  CFA1X1 U4258 ( .A(n2132), .B(n1978), .CI(n2070), .CO(n1402), .S(n1403) );
  COND2X1 U4259 ( .A(n3963), .B(n2627), .C(net16793), .D(n2626), .Z(n2100) );
  CND2X2 U4260 ( .A(n745), .B(n744), .Z(n365) );
  CIVXL U4261 ( .A(n3996), .Z(n3868) );
  CNIVX4 U4262 ( .A(net19401), .Z(net18643) );
  CEOX4 U4263 ( .A(n3704), .B(a[24]), .Z(n2815) );
  CND2IX2 U4264 ( .B(n3870), .A(n4119), .Z(n1981) );
  CHA1X1 U4265 ( .A(n1988), .B(n1731), .CO(n1610), .S(n1611) );
  CENXL U4266 ( .A(net16544), .B(n4343), .Z(n2755) );
  CANR1X1 U4267 ( .A(n3824), .B(n535), .C(n521), .Z(n3871) );
  CANR1X1 U4268 ( .A(n520), .B(n3829), .C(n521), .Z(n515) );
  CIVX3 U4269 ( .A(n3624), .Z(net19151) );
  CEOX2 U4270 ( .A(n3487), .B(a[18]), .Z(n2818) );
  CAN2X1 U4271 ( .A(n3715), .B(n1801), .Z(n4288) );
  CIVX3 U4272 ( .A(n3985), .Z(n3987) );
  CIVX1 U4273 ( .A(n30), .Z(n4176) );
  COND1X2 U4274 ( .A(n530), .B(n522), .C(n523), .Z(n521) );
  COND2X1 U4275 ( .A(n81), .B(n3986), .C(n2515), .D(n3875), .Z(n1731) );
  CEOXL U4276 ( .A(n4341), .B(n3663), .Z(n2649) );
  CND2X2 U4277 ( .A(net18618), .B(net18609), .Z(n4256) );
  CENX1 U4278 ( .A(n4324), .B(net16824), .Z(n2541) );
  CND2XL U4279 ( .A(n1271), .B(n1269), .Z(n4304) );
  CND2XL U4280 ( .A(n1265), .B(n1269), .Z(n4303) );
  CEO3X1 U4281 ( .A(n1827), .B(n1855), .C(n1943), .Z(n1269) );
  CIVX4 U4282 ( .A(n3378), .Z(n3919) );
  COND2X1 U4283 ( .A(net19518), .B(n2543), .C(n4144), .D(n2542), .Z(n2016) );
  COND2X2 U4284 ( .A(n2715), .B(net16816), .C(n2716), .D(n18), .Z(n2189) );
  COND1X2 U4285 ( .A(n573), .B(n3544), .C(n568), .Z(n562) );
  CND2X2 U4286 ( .A(n1333), .B(n1360), .Z(n568) );
  CAN2X1 U4287 ( .A(n1461), .B(n1482), .Z(n3874) );
  CIVX2 U4288 ( .A(n469), .Z(n467) );
  CANR1X1 U4289 ( .A(n748), .B(n415), .C(n408), .Z(n406) );
  CIVX1 U4290 ( .A(n594), .Z(n596) );
  CND2X2 U4291 ( .A(n770), .B(n4267), .Z(n594) );
  COND2X1 U4292 ( .A(n2616), .B(net16793), .C(n2617), .D(n3092), .Z(n2090) );
  COR2XL U4293 ( .A(n1436), .B(n1413), .Z(n3881) );
  CND2X4 U4294 ( .A(net16817), .B(n2826), .Z(n18) );
  CIVX4 U4295 ( .A(net18260), .Z(net16817) );
  CENXL U4296 ( .A(n4327), .B(net18643), .Z(n3876) );
  CND2X4 U4297 ( .A(n2822), .B(net18953), .Z(n3877) );
  CENXL U4298 ( .A(n2810), .B(n4291), .Z(n3878) );
  CNR2X2 U4299 ( .A(n1215), .B(n1244), .Z(n540) );
  CIVXL U4300 ( .A(n3906), .Z(n3880) );
  CENXL U4301 ( .A(n2810), .B(net15995), .Z(n2348) );
  CENXL U4302 ( .A(net16558), .B(n3983), .Z(n2333) );
  CENXL U4303 ( .A(net16550), .B(n3983), .Z(n2329) );
  CEOX2 U4304 ( .A(n943), .B(n958), .Z(n3882) );
  CND2XL U4305 ( .A(n941), .B(n958), .Z(n3883) );
  CND2X1 U4306 ( .A(n941), .B(n943), .Z(n3884) );
  CND2XL U4307 ( .A(n958), .B(n943), .Z(n3885) );
  CND3X1 U4308 ( .A(n3883), .B(n3884), .C(n3885), .Z(n938) );
  CNR2X1 U4309 ( .A(n353), .B(n224), .Z(n222) );
  COR2X1 U4310 ( .A(n3577), .B(n2278), .Z(n3931) );
  CENXL U4311 ( .A(n4342), .B(net16850), .Z(n2450) );
  CND2IXL U4312 ( .B(net16109), .A(net16850), .Z(n2482) );
  COR2XL U4313 ( .A(n63), .B(n2574), .Z(n4085) );
  CEO3X2 U4314 ( .A(n1342), .B(n1319), .C(n1317), .Z(n1311) );
  CND2X1 U4315 ( .A(n3565), .B(n1317), .Z(n3886) );
  CND2XL U4316 ( .A(n1342), .B(n1319), .Z(n3887) );
  CND2X1 U4317 ( .A(n1317), .B(n1319), .Z(n3888) );
  CND3X2 U4318 ( .A(n3886), .B(n3887), .C(n3888), .Z(n1310) );
  CIVXL U4319 ( .A(n3985), .Z(n3889) );
  CENX1 U4320 ( .A(a[26]), .B(net19505), .Z(n2814) );
  CAOR1XL U4321 ( .A(n3709), .B(n3116), .C(n2285), .Z(n1771) );
  COND2XL U4322 ( .A(n2286), .B(n3116), .C(n3709), .D(n2285), .Z(n1772) );
  COND2X1 U4323 ( .A(n4136), .B(n2300), .C(n3709), .D(n2299), .Z(n1785) );
  COND2X1 U4324 ( .A(net18592), .B(n2467), .C(n3278), .D(n2466), .Z(n1942) );
  CIVXL U4325 ( .A(n3263), .Z(n3891) );
  COND2X1 U4326 ( .A(n3092), .B(n2629), .C(net16793), .D(n2628), .Z(n2102) );
  CND2XL U4327 ( .A(n4333), .B(n3894), .Z(n3895) );
  CND2XL U4328 ( .A(n3893), .B(n3195), .Z(n3896) );
  CND2X1 U4329 ( .A(n3895), .B(n3896), .Z(n2463) );
  CIVXL U4330 ( .A(n4333), .Z(n3893) );
  CIVXL U4331 ( .A(net16849), .Z(n3894) );
  CNIVX4 U4332 ( .A(n2793), .Z(n4333) );
  CND2X1 U4333 ( .A(n1266), .B(n3898), .Z(n3899) );
  CND2X2 U4334 ( .A(n3897), .B(n1272), .Z(n3900) );
  CND2X2 U4335 ( .A(n3899), .B(n3900), .Z(n3901) );
  CIVX1 U4336 ( .A(n1272), .Z(n3898) );
  CEOX2 U4337 ( .A(n3901), .B(n1264), .Z(n1231) );
  CND2XL U4338 ( .A(n1264), .B(n1272), .Z(n3902) );
  CND2XL U4339 ( .A(n1264), .B(n1266), .Z(n3903) );
  CND2XL U4340 ( .A(n1272), .B(n1266), .Z(n3904) );
  CND3X1 U4341 ( .A(n3902), .B(n3903), .C(n3904), .Z(n1230) );
  CFA1X1 U4342 ( .A(n1840), .B(n1870), .CI(n1782), .CO(n902), .S(n903) );
  CIVX2 U4343 ( .A(n4346), .Z(n4345) );
  CND2X2 U4344 ( .A(n2827), .B(n6), .Z(n9) );
  CEOX2 U4345 ( .A(n1403), .B(n1426), .Z(n4220) );
  COND2XL U4346 ( .A(n3024), .B(n2702), .C(net16772), .D(n2701), .Z(n2175) );
  COND2XL U4347 ( .A(n2253), .B(n3577), .C(n2254), .D(n144), .Z(n1741) );
  COND2XL U4348 ( .A(n144), .B(n2258), .C(n3577), .D(n2257), .Z(n1744) );
  COND2XL U4349 ( .A(n144), .B(n2259), .C(n3577), .D(n2258), .Z(n1745) );
  CND2XL U4350 ( .A(a[12]), .B(n4307), .Z(n3907) );
  CND2X2 U4351 ( .A(n3907), .B(n3908), .Z(n4012) );
  CIVXL U4352 ( .A(a[12]), .Z(n3905) );
  CIVX1 U4353 ( .A(n4307), .Z(n3906) );
  CIVX1 U4354 ( .A(n4307), .Z(n4145) );
  CIVX1 U4355 ( .A(n4307), .Z(n4349) );
  CND2X1 U4356 ( .A(n1096), .B(n1073), .Z(n3909) );
  CND2X1 U4357 ( .A(n1096), .B(n1079), .Z(n3910) );
  CND2XL U4358 ( .A(n1073), .B(n1079), .Z(n3911) );
  CEOX2 U4359 ( .A(n1169), .B(n1194), .Z(n3912) );
  CND2X1 U4360 ( .A(n1167), .B(n3225), .Z(n3913) );
  CND2X1 U4361 ( .A(n1167), .B(n1169), .Z(n3914) );
  CEOX2 U4362 ( .A(n4036), .B(n3619), .Z(n1135) );
  CEO3X1 U4363 ( .A(n2165), .B(n2010), .C(n1950), .Z(n1453) );
  CND2XL U4364 ( .A(n1985), .B(n1926), .Z(n3916) );
  CND2XL U4365 ( .A(n1985), .B(n2108), .Z(n3917) );
  CND3X1 U4366 ( .A(n3916), .B(n3917), .C(n3918), .Z(n1560) );
  CNR2IXL U4367 ( .B(n145), .A(n3920), .Z(n1926) );
  COND2X1 U4368 ( .A(n81), .B(n2511), .C(n78), .D(n2510), .Z(n1985) );
  COND2X1 U4369 ( .A(n54), .B(n2596), .C(n3839), .D(n2595), .Z(n2069) );
  CND2X1 U4370 ( .A(n1271), .B(n1265), .Z(n4302) );
  CND2XL U4371 ( .A(n2176), .B(n2083), .Z(n3921) );
  CND2XL U4372 ( .A(n2176), .B(n2021), .Z(n3922) );
  CND3X1 U4373 ( .A(n3921), .B(n3922), .C(n3923), .Z(n1650) );
  CNR2XL U4374 ( .A(net16772), .B(n2702), .Z(n3925) );
  COR2X1 U4375 ( .A(n3924), .B(n3925), .Z(n2176) );
  CND2X1 U4376 ( .A(n1641), .B(n1652), .Z(n672) );
  CANR1XL U4377 ( .A(n4267), .B(n3788), .C(n601), .Z(n3926) );
  CIVX2 U4378 ( .A(n4355), .Z(n4252) );
  CIVX1 U4379 ( .A(n3334), .Z(n4355) );
  CENX1 U4380 ( .A(net16558), .B(n4253), .Z(n2399) );
  CND2IXL U4381 ( .B(net16109), .A(net16093), .Z(n2746) );
  CENXL U4382 ( .A(n4332), .B(net16093), .Z(n2728) );
  CENXL U4383 ( .A(n4330), .B(net16093), .Z(n2731) );
  CENXL U4384 ( .A(n4331), .B(net16093), .Z(n2730) );
  CEO3X2 U4385 ( .A(n1182), .B(n1180), .C(n1178), .Z(n1147) );
  CND2X1 U4386 ( .A(n1178), .B(n1180), .Z(n3929) );
  COR2X1 U4387 ( .A(n4261), .B(n2279), .Z(n3930) );
  CND2X2 U4388 ( .A(n3930), .B(n3931), .Z(n1765) );
  CENXL U4389 ( .A(n4322), .B(n4362), .Z(n2279) );
  CENXL U4390 ( .A(n4323), .B(n4362), .Z(n2278) );
  COND2X2 U4391 ( .A(n4188), .B(n2403), .C(net16839), .D(n2402), .Z(n1881) );
  CEOX1 U4392 ( .A(n4329), .B(n4087), .Z(n2402) );
  CENX2 U4393 ( .A(n3764), .B(n3932), .Z(n1307) );
  CND2X2 U4394 ( .A(n4354), .B(a[24]), .Z(n3944) );
  CIVXL U4395 ( .A(n770), .Z(n3933) );
  CIVX1 U4396 ( .A(n605), .Z(n770) );
  CIVXL U4397 ( .A(n3510), .Z(n1185) );
  CENX1 U4398 ( .A(n4171), .B(n3574), .Z(n4018) );
  CANR1XL U4399 ( .A(n3621), .B(n621), .C(n616), .Z(n3935) );
  CEO3X2 U4400 ( .A(n1883), .B(n1972), .C(n2095), .Z(n1235) );
  CND2XL U4401 ( .A(n1883), .B(n1972), .Z(n3936) );
  CND2XL U4402 ( .A(n1883), .B(n2095), .Z(n3937) );
  CND2XL U4403 ( .A(n1972), .B(n2095), .Z(n3938) );
  CND3X1 U4404 ( .A(n3936), .B(n3937), .C(n3938), .Z(n1234) );
  CND2XL U4405 ( .A(n1270), .B(n1268), .Z(n3939) );
  CND2X1 U4406 ( .A(n1270), .B(n1235), .Z(n3940) );
  CND2X1 U4407 ( .A(n1268), .B(n1235), .Z(n3941) );
  CENX1 U4408 ( .A(n4234), .B(n1226), .Z(n1195) );
  COAN1X1 U4409 ( .A(n369), .B(n379), .C(n370), .Z(n366) );
  CIVX4 U4410 ( .A(n4026), .Z(n4347) );
  CFA1X1 U4411 ( .A(n1846), .B(n2025), .CI(n1789), .CO(n1030), .S(n1031) );
  COND2X1 U4412 ( .A(n2552), .B(n63), .C(net19500), .D(n2551), .Z(n2025) );
  CND2X4 U4413 ( .A(n3942), .B(n3943), .Z(n3945) );
  CND2X4 U4414 ( .A(n3944), .B(n3945), .Z(n114) );
  CIVX2 U4415 ( .A(a[24]), .Z(n3942) );
  CND2X4 U4416 ( .A(n114), .B(n2815), .Z(net19417) );
  CENXL U4417 ( .A(n4338), .B(net16843), .Z(n4141) );
  CENXL U4418 ( .A(n4330), .B(net16087), .Z(n2698) );
  CENXL U4419 ( .A(n4331), .B(net16087), .Z(n2697) );
  CENXL U4420 ( .A(n4332), .B(net16087), .Z(n2695) );
  CENXL U4421 ( .A(net16558), .B(net16087), .Z(n2696) );
  CENXL U4422 ( .A(n4333), .B(net16087), .Z(n2694) );
  CENXL U4423 ( .A(n4329), .B(net16087), .Z(n2699) );
  CND2IXL U4424 ( .B(net16109), .A(net16087), .Z(n2713) );
  CAOR1XL U4425 ( .A(n78), .B(n81), .C(n2483), .Z(n1958) );
  CND2XL U4426 ( .A(n1283), .B(n1308), .Z(n4218) );
  CEOX2 U4427 ( .A(n1164), .B(n1139), .Z(n4036) );
  COND1XL U4428 ( .A(n3312), .B(n651), .C(n3039), .Z(n3947) );
  CIVXL U4429 ( .A(n415), .Z(n413) );
  CIVXL U4430 ( .A(n3269), .Z(n419) );
  CIVXL U4431 ( .A(n4292), .Z(n3948) );
  CENX1 U4432 ( .A(n4323), .B(n4291), .Z(n2377) );
  COND2X1 U4433 ( .A(n2481), .B(net18593), .C(n3277), .D(n2480), .Z(n1956) );
  CIVX2 U4434 ( .A(net19047), .Z(net19048) );
  COND2X1 U4435 ( .A(n117), .B(n3891), .C(net16784), .D(n2383), .Z(n1727) );
  CND2XL U4436 ( .A(n1470), .B(n1449), .Z(n3949) );
  CND2XL U4437 ( .A(n1470), .B(n1472), .Z(n3950) );
  CND2X1 U4438 ( .A(n1449), .B(n1472), .Z(n3951) );
  CND3X1 U4439 ( .A(n3949), .B(n3950), .C(n3951), .Z(n1442) );
  COND2XL U4440 ( .A(n3092), .B(n2645), .C(net16793), .D(n2644), .Z(n2118) );
  COND2XL U4441 ( .A(n3092), .B(n2641), .C(net16793), .D(n2640), .Z(n2114) );
  COND2XL U4442 ( .A(n3092), .B(n2628), .C(net16793), .D(n2627), .Z(n2101) );
  COND2XL U4443 ( .A(n3963), .B(n2642), .C(net16793), .D(n2641), .Z(n2115) );
  COND2XL U4444 ( .A(n3092), .B(n2631), .C(net16793), .D(n2630), .Z(n2104) );
  COND2XL U4445 ( .A(n3092), .B(n2636), .C(net16793), .D(n2635), .Z(n2109) );
  COND2XL U4446 ( .A(n3092), .B(n2637), .C(net16793), .D(n2636), .Z(n2110) );
  COND2X1 U4447 ( .A(n45), .B(n2639), .C(net16793), .D(n2638), .Z(n2112) );
  CNIVX4 U4448 ( .A(net16083), .Z(net16844) );
  CEO3X2 U4449 ( .A(n2096), .B(n2220), .C(n3074), .Z(n1263) );
  CND2XL U4450 ( .A(n1302), .B(n2096), .Z(n3953) );
  CND2X1 U4451 ( .A(n2096), .B(n2220), .Z(n3954) );
  CND2X1 U4452 ( .A(n1302), .B(n2220), .Z(n3955) );
  CND3X1 U4453 ( .A(n3953), .B(n3954), .C(n3955), .Z(n1262) );
  CND2X1 U4454 ( .A(n1267), .B(n1263), .Z(n3957) );
  CND2X1 U4455 ( .A(n1218), .B(n3615), .Z(n3959) );
  CND2X1 U4456 ( .A(n3615), .B(n1220), .Z(n3961) );
  CND3X2 U4457 ( .A(n3959), .B(n3960), .C(n3961), .Z(n1188) );
  CND2X2 U4458 ( .A(n3202), .B(n753), .Z(n460) );
  CENX1 U4459 ( .A(n4332), .B(n4253), .Z(n2398) );
  CND2X2 U4460 ( .A(n2823), .B(n3235), .Z(n45) );
  CEO3X2 U4461 ( .A(n1063), .B(n1084), .C(n1061), .Z(n1059) );
  CND2XL U4462 ( .A(n3605), .B(n1061), .Z(n3965) );
  CND2XL U4463 ( .A(n3605), .B(n1063), .Z(n3966) );
  CNR2IX1 U4464 ( .B(net16109), .A(net16838), .Z(n1894) );
  CND2X1 U4465 ( .A(n4025), .B(n1098), .Z(n3970) );
  CND2X2 U4466 ( .A(n3968), .B(n3969), .Z(n3971) );
  CND2X2 U4467 ( .A(n3970), .B(n3971), .Z(n1071) );
  CIVXL U4468 ( .A(n1098), .Z(n3969) );
  CENX1 U4469 ( .A(n1104), .B(n1100), .Z(n4025) );
  CEOX2 U4470 ( .A(n1509), .B(n1526), .Z(n3972) );
  CEOX2 U4471 ( .A(n3972), .B(n1507), .Z(n1505) );
  CND2XL U4472 ( .A(n1507), .B(n1526), .Z(n3973) );
  CND2X1 U4473 ( .A(n1507), .B(n1509), .Z(n3974) );
  CND2XL U4474 ( .A(n1526), .B(n1509), .Z(n3975) );
  CEOX2 U4475 ( .A(n1294), .B(n1273), .Z(n3976) );
  CEOX2 U4476 ( .A(n3976), .B(n3418), .Z(n1261) );
  CND2XL U4477 ( .A(n1296), .B(n1273), .Z(n3977) );
  CND2XL U4478 ( .A(n1296), .B(n1294), .Z(n3978) );
  CND2XL U4479 ( .A(n1273), .B(n1294), .Z(n3979) );
  CND3X1 U4480 ( .A(n3977), .B(n3978), .C(n3979), .Z(n1260) );
  CENX1 U4481 ( .A(a[12]), .B(n4307), .Z(n2821) );
  CND2X4 U4482 ( .A(n3875), .B(n3412), .Z(n81) );
  COR2XL U4483 ( .A(n1505), .B(n1524), .Z(n3980) );
  CENX1 U4484 ( .A(n4333), .B(net18936), .Z(n2529) );
  CENXL U4485 ( .A(n230), .B(n151), .Z(product[61]) );
  CANR1X1 U4486 ( .A(n359), .B(n3659), .C(n360), .Z(n354) );
  COND1X1 U4487 ( .A(n547), .B(n3869), .C(n548), .Z(net19465) );
  CND2XL U4488 ( .A(n355), .B(n233), .Z(n231) );
  COAN1X1 U4489 ( .A(n266), .B(n241), .C(n242), .Z(n3981) );
  CIVX2 U4490 ( .A(n246), .Z(n244) );
  CIVX2 U4491 ( .A(n255), .Z(n253) );
  CANR1X1 U4492 ( .A(n735), .B(n260), .C(n253), .Z(n249) );
  CNR2X2 U4493 ( .A(n3421), .B(n416), .Z(n359) );
  CANR1X1 U4494 ( .A(n359), .B(n3659), .C(n3823), .Z(net19530) );
  CIVX2 U4495 ( .A(n449), .Z(n447) );
  CANR1X1 U4496 ( .A(n456), .B(n751), .C(n447), .Z(n445) );
  CND2X1 U4497 ( .A(net18421), .B(n229), .Z(n151) );
  COR2X1 U4498 ( .A(n796), .B(n795), .Z(net18421) );
  CIVX2 U4499 ( .A(n794), .Z(n795) );
  CND2X1 U4500 ( .A(n796), .B(n795), .Z(n229) );
  CIVX2 U4501 ( .A(n229), .Z(n227) );
  CND2X1 U4502 ( .A(n1343), .B(n1368), .Z(net19204) );
  CEO3X2 U4503 ( .A(n1343), .B(n1368), .C(n1366), .Z(n1337) );
  CND2X1 U4504 ( .A(n1366), .B(n1368), .Z(net19205) );
  CENXL U4505 ( .A(net16107), .B(net15995), .Z(n2349) );
  CIVX4 U4506 ( .A(n3984), .Z(net15995) );
  CIVX1 U4507 ( .A(n120), .Z(n3984) );
  CIVXL U4508 ( .A(n3984), .Z(n3983) );
  CNIVX1 U4509 ( .A(n145), .Z(net16107) );
  CND2IXL U4510 ( .B(net16109), .A(n3983), .Z(n2350) );
  CENXL U4511 ( .A(net16544), .B(n3983), .Z(n2326) );
  CNIVX4 U4512 ( .A(n105), .Z(net16839) );
  COND2X1 U4513 ( .A(n3877), .B(n2598), .C(n3839), .D(n2597), .Z(n2071) );
  CEO3XL U4514 ( .A(n1365), .B(n1388), .C(n1363), .Z(net19133) );
  CENX4 U4515 ( .A(a[18]), .B(n3986), .Z(net16644) );
  CIVX4 U4516 ( .A(n3986), .Z(net16037) );
  CIVX4 U4517 ( .A(a[0]), .Z(n6) );
  CND2X2 U4518 ( .A(n1305), .B(n1332), .Z(n559) );
  CND2X1 U4519 ( .A(n1366), .B(n1343), .Z(net19203) );
  CND3X2 U4520 ( .A(n3992), .B(n3993), .C(n3994), .Z(n1396) );
  CND2X1 U4521 ( .A(n1426), .B(n1409), .Z(n3994) );
  CND2X1 U4522 ( .A(n1403), .B(n1409), .Z(n3993) );
  CND2X1 U4523 ( .A(n1403), .B(n1426), .Z(n3992) );
  CND3X1 U4524 ( .A(n3991), .B(n3990), .C(n3989), .Z(n1408) );
  CND2XL U4525 ( .A(n2225), .B(n3800), .Z(n3991) );
  CND2XL U4526 ( .A(n2039), .B(n3800), .Z(n3990) );
  CND2XL U4527 ( .A(n2039), .B(n2225), .Z(n3989) );
  CIVX2 U4528 ( .A(n39), .Z(net18816) );
  COND2XL U4529 ( .A(n3092), .B(net18817), .C(net16793), .D(n2647), .Z(n1735)
         );
  CIVXL U4530 ( .A(n3866), .Z(n574) );
  COND1X2 U4531 ( .A(n578), .B(n595), .C(n579), .Z(n577) );
  COAN1X1 U4532 ( .A(net19292), .B(n582), .C(n583), .Z(n579) );
  COND1X2 U4533 ( .A(n3442), .B(n630), .C(n614), .Z(net18451) );
  CANR1X2 U4534 ( .A(n3480), .B(n650), .C(n632), .Z(n630) );
  CNR2XL U4535 ( .A(n572), .B(n3544), .Z(net19307) );
  CIVXL U4536 ( .A(n3926), .Z(n597) );
  COR2X1 U4537 ( .A(n1436), .B(n1413), .Z(net19316) );
  COND1X1 U4538 ( .A(n3442), .B(net19200), .C(n3935), .Z(n612) );
  CANR1XL U4539 ( .A(n3947), .B(n3025), .C(n3105), .Z(net19200) );
  CIVXL U4540 ( .A(n3947), .Z(n649) );
  CENXL U4541 ( .A(n219), .B(n150), .Z(product[62]) );
  CIVXL U4542 ( .A(n223), .Z(n221) );
  CIVXL U4543 ( .A(n222), .Z(n220) );
  CNR2X2 U4544 ( .A(n1059), .B(n3405), .Z(n484) );
  CNIVX4 U4545 ( .A(n3995), .Z(n3997) );
  CIVX2 U4546 ( .A(n3996), .Z(n3995) );
  CNIVX4 U4547 ( .A(n3995), .Z(net18937) );
  CIVX2 U4548 ( .A(n66), .Z(n3996) );
  CENXL U4549 ( .A(a[14]), .B(n3996), .Z(n2820) );
  CIVX2 U4550 ( .A(n3996), .Z(net19401) );
  CNIVX8 U4551 ( .A(n2801), .Z(net16570) );
  CIVXL U4552 ( .A(n562), .Z(n564) );
  CND2X1 U4553 ( .A(net19133), .B(n1386), .Z(n573) );
  CND2XL U4554 ( .A(n766), .B(n573), .Z(n184) );
  CIVX1 U4555 ( .A(n573), .Z(n571) );
  CND2X1 U4556 ( .A(net18420), .B(n218), .Z(n150) );
  COR2X1 U4557 ( .A(n1740), .B(n794), .Z(net18420) );
  CND2XL U4558 ( .A(n222), .B(net18420), .Z(n213) );
  CND2X1 U4559 ( .A(n1740), .B(n794), .Z(n218) );
  CIVX2 U4560 ( .A(n218), .Z(n216) );
  CNR2X2 U4561 ( .A(n551), .B(n556), .Z(net18739) );
  CNR2X1 U4562 ( .A(n3040), .B(n1304), .Z(n551) );
  COND1XL U4563 ( .A(n556), .B(n564), .C(n3300), .Z(n555) );
  CNR2X2 U4564 ( .A(n3040), .B(n1304), .Z(net18620) );
  CND2X1 U4565 ( .A(n1275), .B(n1304), .Z(n552) );
  CIVX1 U4566 ( .A(net18620), .Z(n763) );
  CND2XL U4567 ( .A(n3034), .B(n763), .Z(n181) );
  CNR2IXL U4568 ( .B(net19307), .A(n556), .Z(n554) );
  CIVXL U4569 ( .A(n514), .Z(n516) );
  CND2X2 U4570 ( .A(n4029), .B(n482), .Z(n480) );
  COND1XL U4571 ( .A(n491), .B(net19517), .C(n494), .Z(n490) );
  COND2XL U4572 ( .A(net18743), .B(n2692), .C(net16772), .D(n2691), .Z(
        net18875) );
  CNIVX4 U4573 ( .A(n3998), .Z(net16843) );
  CENX4 U4574 ( .A(a[6]), .B(n3543), .Z(net19508) );
  CENX1 U4575 ( .A(a[6]), .B(n3543), .Z(net16791) );
  CIVX2 U4576 ( .A(n21), .Z(net16089) );
  CIVXL U4577 ( .A(n21), .Z(net18981) );
  CND2X2 U4578 ( .A(n2825), .B(n24), .Z(net18743) );
  CENX4 U4579 ( .A(a[4]), .B(n3219), .Z(net16772) );
  CIVX4 U4580 ( .A(n3999), .Z(net16091) );
  CENX1 U4581 ( .A(n2789), .B(net16843), .Z(n2690) );
  CEOX2 U4582 ( .A(a[4]), .B(net16083), .Z(n2825) );
  CIVX1 U4583 ( .A(n12), .Z(net19016) );
  CIVX3 U4584 ( .A(n4307), .Z(n4000) );
  CEOX1 U4585 ( .A(n4327), .B(n4290), .Z(n2371) );
  CND2X4 U4586 ( .A(net16817), .B(n2826), .Z(n4001) );
  CENX2 U4587 ( .A(n3762), .B(n4009), .Z(n1187) );
  CND2X2 U4588 ( .A(n4172), .B(n33), .Z(n4002) );
  CND2X2 U4589 ( .A(n4172), .B(n33), .Z(n4003) );
  CND2X4 U4590 ( .A(n2827), .B(n6), .Z(net19555) );
  CIVX2 U4591 ( .A(n120), .Z(net19505) );
  CIVX2 U4592 ( .A(n4087), .Z(n4004) );
  CND2IX1 U4593 ( .B(a[22]), .A(n4264), .Z(n4266) );
  CIVX2 U4594 ( .A(net16065), .Z(net16063) );
  CIVX3 U4595 ( .A(net19076), .Z(net16059) );
  CENX1 U4596 ( .A(n1571), .B(n1584), .Z(n4006) );
  CND2XL U4597 ( .A(n1109), .B(n1111), .Z(n4319) );
  CNIVX1 U4598 ( .A(n2123), .Z(n4007) );
  COAN1XL U4599 ( .A(n274), .B(n3777), .C(n3112), .Z(n269) );
  CND2XL U4600 ( .A(n3623), .B(n748), .Z(n405) );
  CND2XL U4601 ( .A(n414), .B(n3220), .Z(n394) );
  CIVX2 U4602 ( .A(n4143), .Z(n4144) );
  CENXL U4603 ( .A(n2802), .B(n3308), .Z(n2406) );
  CND2XL U4604 ( .A(n4233), .B(n2820), .Z(n4008) );
  CIVXL U4605 ( .A(net19517), .Z(net19522) );
  CEO3XL U4606 ( .A(n1417), .B(n1438), .C(n1415), .Z(net19521) );
  COAN1XL U4607 ( .A(n512), .B(n3660), .C(n505), .Z(net19517) );
  CEOX2 U4608 ( .A(a[24]), .B(n3704), .Z(n4010) );
  CEOX1 U4609 ( .A(n4155), .B(n1051), .Z(n1047) );
  COAN1XL U4610 ( .A(n410), .B(n402), .C(n403), .Z(n4011) );
  CEO3X2 U4611 ( .A(n4051), .B(n1968), .C(n1131), .Z(n1099) );
  CENX1 U4612 ( .A(n1455), .B(n1457), .Z(n4013) );
  CIVXL U4613 ( .A(n129), .Z(n4014) );
  CND2XL U4614 ( .A(n1108), .B(n3132), .Z(n4224) );
  COND2XL U4615 ( .A(net19122), .B(n2391), .C(net19462), .D(n2390), .Z(n1871)
         );
  COND2XL U4616 ( .A(net19122), .B(n2393), .C(net16839), .D(n2392), .Z(n4016)
         );
  COND2X1 U4617 ( .A(n2393), .B(net19122), .C(net16839), .D(n2392), .Z(n954)
         );
  CENXL U4618 ( .A(n4171), .B(n3574), .Z(n4017) );
  CAOR1XL U4619 ( .A(n753), .B(n3602), .C(n467), .Z(n4019) );
  CENX2 U4620 ( .A(n4327), .B(net16059), .Z(n2602) );
  CENX2 U4621 ( .A(net16570), .B(n3729), .Z(n2603) );
  CNIVX4 U4622 ( .A(n105), .Z(net19462) );
  COAN1X1 U4623 ( .A(n444), .B(n461), .C(n445), .Z(n4020) );
  CIVXL U4624 ( .A(n4098), .Z(n4021) );
  CIVXL U4625 ( .A(n511), .Z(n758) );
  CENX2 U4626 ( .A(n4022), .B(n1300), .Z(n1259) );
  CENX1 U4627 ( .A(n1298), .B(n1292), .Z(n4022) );
  CNIVX1 U4628 ( .A(n1821), .Z(n4023) );
  CNIVX1 U4629 ( .A(n2011), .Z(n4024) );
  CND2XL U4630 ( .A(n2123), .B(n2092), .Z(n4057) );
  CENXL U4631 ( .A(net16544), .B(net18618), .Z(n2491) );
  CENXL U4632 ( .A(n4337), .B(net18618), .Z(n2488) );
  CENXL U4633 ( .A(n2789), .B(net18618), .Z(n2492) );
  CENXL U4634 ( .A(n4340), .B(net18618), .Z(n2485) );
  CENXL U4635 ( .A(n4339), .B(n3023), .Z(n2486) );
  CENXL U4636 ( .A(n4334), .B(net18618), .Z(n2495) );
  CENXL U4637 ( .A(net16550), .B(net18618), .Z(n2494) );
  CENXL U4638 ( .A(n4335), .B(net18618), .Z(n2490) );
  CENXL U4639 ( .A(n4338), .B(net18618), .Z(n2487) );
  CENXL U4640 ( .A(net16548), .B(net18618), .Z(n2493) );
  CENXL U4641 ( .A(n4336), .B(n3023), .Z(n2489) );
  CENXL U4642 ( .A(n4341), .B(net18618), .Z(n2484) );
  CIVXL U4643 ( .A(n512), .Z(n510) );
  CIVX2 U4644 ( .A(n30), .Z(n4026) );
  CIVXL U4645 ( .A(n4020), .Z(n4027) );
  CENX1 U4646 ( .A(n4328), .B(n4291), .Z(n2370) );
  CNIVX2 U4647 ( .A(n2068), .Z(n4028) );
  CENX2 U4648 ( .A(n4031), .B(n4032), .Z(n1215) );
  COND2X1 U4649 ( .A(n9), .B(n2763), .C(n6), .D(n2762), .Z(n2236) );
  CND2IX1 U4650 ( .B(n1163), .A(n1188), .Z(n4100) );
  COND1XL U4651 ( .A(n372), .B(net18543), .C(n373), .Z(n371) );
  CIVX1 U4652 ( .A(n865), .Z(n4034) );
  CIVX1 U4653 ( .A(n864), .Z(n865) );
  CENXL U4654 ( .A(n1884), .B(n1914), .Z(n4035) );
  CND2XL U4655 ( .A(n3106), .B(n1139), .Z(n4037) );
  CND3X1 U4656 ( .A(n4037), .B(n4038), .C(n4039), .Z(n1134) );
  COND2X1 U4657 ( .A(n2654), .B(n36), .C(net16791), .D(n2653), .Z(n2127) );
  CENXL U4658 ( .A(n4341), .B(net16843), .Z(n4040) );
  CAOR1XL U4659 ( .A(n4289), .B(n3757), .C(n2516), .Z(n1990) );
  CNR2X1 U4660 ( .A(n671), .B(n674), .Z(n669) );
  COND2X1 U4661 ( .A(net18743), .B(n2706), .C(net16772), .D(n2705), .Z(n2179)
         );
  CND2XL U4662 ( .A(n1236), .B(n1232), .Z(n4041) );
  CND2X1 U4663 ( .A(n1236), .B(n1234), .Z(n4042) );
  CND2XL U4664 ( .A(n1232), .B(n1234), .Z(n4043) );
  CND3X1 U4665 ( .A(n4041), .B(n4042), .C(n4043), .Z(n1200) );
  CIVX2 U4666 ( .A(n4358), .Z(n4357) );
  CIVXL U4667 ( .A(n564), .Z(net19388) );
  CENXL U4668 ( .A(n4325), .B(net16091), .Z(n2738) );
  CENXL U4669 ( .A(net16548), .B(net16091), .Z(n2724) );
  CENXL U4670 ( .A(n2789), .B(net16091), .Z(n2723) );
  CENXL U4671 ( .A(n4340), .B(net16091), .Z(n2716) );
  CENXL U4672 ( .A(net16550), .B(net16091), .Z(n2725) );
  CENXL U4673 ( .A(n4339), .B(net16091), .Z(n2717) );
  CENXL U4674 ( .A(n4338), .B(net16091), .Z(n2718) );
  CENXL U4675 ( .A(n4337), .B(net16091), .Z(n2719) );
  CENXL U4676 ( .A(n4334), .B(net16091), .Z(n2726) );
  CENXL U4677 ( .A(n4336), .B(net16091), .Z(n2720) );
  CENXL U4678 ( .A(n4335), .B(net16091), .Z(n2721) );
  CENXL U4679 ( .A(net16544), .B(net16091), .Z(n2722) );
  CIVXL U4680 ( .A(n597), .Z(net19384) );
  CND2XL U4681 ( .A(n4052), .B(n1968), .Z(n4045) );
  CND2XL U4682 ( .A(n4052), .B(n1130), .Z(n4046) );
  CND2XL U4683 ( .A(n1968), .B(n1130), .Z(n4047) );
  CND3X1 U4684 ( .A(n4045), .B(n4046), .C(n4047), .Z(n1098) );
  CND2XL U4685 ( .A(n1104), .B(n1100), .Z(n4048) );
  CND2XL U4686 ( .A(n1104), .B(n1098), .Z(n4049) );
  CND2XL U4687 ( .A(n1100), .B(n1098), .Z(n4050) );
  CIVXL U4688 ( .A(n4051), .Z(n4052) );
  CND3XL U4689 ( .A(n4181), .B(n4180), .C(n4182), .Z(n4054) );
  CEO3X1 U4690 ( .A(n3044), .B(n4007), .C(n4063), .Z(n1157) );
  CND2XL U4691 ( .A(n3044), .B(n2123), .Z(n4055) );
  CND2XL U4692 ( .A(n1764), .B(n2092), .Z(n4056) );
  CND3X1 U4693 ( .A(n4055), .B(n4056), .C(n4057), .Z(n1156) );
  CEOX2 U4694 ( .A(n1156), .B(n4058), .Z(n1121) );
  CND2XL U4695 ( .A(n1131), .B(n1154), .Z(n4059) );
  CND2X1 U4696 ( .A(n1131), .B(n1156), .Z(n4060) );
  CND2XL U4697 ( .A(n1154), .B(n1156), .Z(n4061) );
  CND3X1 U4698 ( .A(n4059), .B(n4060), .C(n4061), .Z(n1120) );
  CIVXL U4699 ( .A(n2092), .Z(n4062) );
  CIVX1 U4700 ( .A(n4062), .Z(n4063) );
  COND2XL U4701 ( .A(n3963), .B(n2619), .C(n4018), .D(n2618), .Z(n2092) );
  CND2XL U4702 ( .A(n1118), .B(n1120), .Z(n4064) );
  CND2XL U4703 ( .A(n1118), .B(n1101), .Z(n4065) );
  CND2XL U4704 ( .A(n1120), .B(n1101), .Z(n4066) );
  CND3X1 U4705 ( .A(n4064), .B(n4065), .C(n4066), .Z(n1090) );
  CEOX1 U4706 ( .A(n985), .B(n1002), .Z(n4067) );
  CND2X1 U4707 ( .A(n1008), .B(n1006), .Z(n4069) );
  CND3X2 U4708 ( .A(n4068), .B(n4069), .C(n4070), .Z(n982) );
  CND2X1 U4709 ( .A(n985), .B(n1002), .Z(n4071) );
  CND2X1 U4710 ( .A(n983), .B(n985), .Z(n4072) );
  CND2X1 U4711 ( .A(n1002), .B(n983), .Z(n4073) );
  CND3X2 U4712 ( .A(n4073), .B(n4072), .C(n4071), .Z(n978) );
  COR2X1 U4713 ( .A(net18897), .B(n2426), .Z(n4074) );
  CENXL U4714 ( .A(n2789), .B(n4352), .Z(n2426) );
  CIVX4 U4715 ( .A(n129), .Z(n4361) );
  CND2XL U4716 ( .A(n1116), .B(n1095), .Z(n4076) );
  CND2XL U4717 ( .A(n1116), .B(n1097), .Z(n4077) );
  CND2X1 U4718 ( .A(n1095), .B(n1097), .Z(n4078) );
  CND3X1 U4719 ( .A(n4076), .B(n4077), .C(n4078), .Z(n1088) );
  CEO3X2 U4720 ( .A(n1590), .B(n1575), .C(n1573), .Z(n1569) );
  CND3X2 U4721 ( .A(n4079), .B(n4080), .C(n4081), .Z(n1568) );
  CND2X1 U4722 ( .A(n1571), .B(n1569), .Z(n4083) );
  COND2XL U4723 ( .A(n3415), .B(n2538), .C(n4144), .D(n2537), .Z(n2011) );
  CNR2IXL U4724 ( .B(n4029), .A(n491), .Z(n489) );
  CND2XL U4725 ( .A(n505), .B(n757), .Z(n175) );
  CND2X2 U4726 ( .A(n1187), .B(n1214), .Z(n530) );
  COND2XL U4727 ( .A(n2319), .B(n3606), .C(net16802), .D(n2318), .Z(n1804) );
  COND2XL U4728 ( .A(n3607), .B(n2321), .C(net16802), .D(n2320), .Z(n824) );
  COND2XL U4729 ( .A(n3607), .B(n2322), .C(net16802), .D(n2321), .Z(n1806) );
  COND2XL U4730 ( .A(n3606), .B(n2326), .C(net16802), .D(n2325), .Z(n1809) );
  COND2XL U4731 ( .A(n3606), .B(n2330), .C(net16802), .D(n2329), .Z(n1813) );
  COND2XL U4732 ( .A(n126), .B(n2341), .C(net16802), .D(n2340), .Z(n1824) );
  CHA1X1 U4733 ( .A(n1728), .B(n1893), .CO(n1502), .S(n1503) );
  COND2X1 U4734 ( .A(n4188), .B(n4087), .C(net16839), .D(n2416), .Z(n1728) );
  CNIVX4 U4735 ( .A(n4348), .Z(n4254) );
  CENXL U4736 ( .A(n4342), .B(net15995), .Z(n2318) );
  CENXL U4737 ( .A(n4341), .B(net15995), .Z(n2319) );
  CENXL U4738 ( .A(n4340), .B(net15995), .Z(n2320) );
  CENXL U4739 ( .A(n4339), .B(net15995), .Z(n2321) );
  CENXL U4740 ( .A(n2789), .B(net15995), .Z(n2327) );
  CENXL U4741 ( .A(n4337), .B(net15995), .Z(n2323) );
  CENXL U4742 ( .A(n4332), .B(net15995), .Z(n2332) );
  CENXL U4743 ( .A(n4330), .B(net15995), .Z(n2335) );
  CENXL U4744 ( .A(n4335), .B(net15995), .Z(n2325) );
  CENXL U4745 ( .A(n4333), .B(net15995), .Z(n2331) );
  CENXL U4746 ( .A(n4338), .B(net15995), .Z(n2322) );
  CENXL U4747 ( .A(n4326), .B(net15995), .Z(n2341) );
  CENXL U4748 ( .A(net16548), .B(net15995), .Z(n2328) );
  CENXL U4749 ( .A(n4336), .B(net15995), .Z(n2324) );
  CENXL U4750 ( .A(n4325), .B(net15995), .Z(n2342) );
  CENXL U4751 ( .A(n4334), .B(net15995), .Z(n2330) );
  CENXL U4752 ( .A(n4321), .B(net15995), .Z(n2347) );
  CENXL U4753 ( .A(n4331), .B(net15995), .Z(n2334) );
  CENXL U4754 ( .A(n4327), .B(net15995), .Z(n2338) );
  CENXL U4755 ( .A(net16570), .B(net15995), .Z(n2339) );
  CENXL U4756 ( .A(n2802), .B(net15995), .Z(n2340) );
  CENXL U4757 ( .A(n4328), .B(net15995), .Z(n2337) );
  CENXL U4758 ( .A(n4323), .B(net15995), .Z(n2344) );
  CIVXL U4759 ( .A(n3103), .Z(n774) );
  CIVX2 U4760 ( .A(n4353), .Z(n4258) );
  CND2X1 U4761 ( .A(n1310), .B(n1312), .Z(n4179) );
  COND2X1 U4762 ( .A(n2382), .B(net19417), .C(n4295), .D(n2381), .Z(n1862) );
  CND2X2 U4763 ( .A(n4276), .B(n3129), .Z(n416) );
  CENXL U4764 ( .A(n4333), .B(net16067), .Z(n2628) );
  CENXL U4765 ( .A(n4331), .B(net16067), .Z(n2631) );
  CND2IXL U4766 ( .B(net16109), .A(net16067), .Z(n2647) );
  CENXL U4767 ( .A(n4337), .B(net16067), .Z(n2620) );
  CENXL U4768 ( .A(net16544), .B(net16067), .Z(n2623) );
  CENXL U4769 ( .A(n2789), .B(net16067), .Z(n2624) );
  CENXL U4770 ( .A(n4329), .B(net16067), .Z(n2633) );
  CENXL U4771 ( .A(net16558), .B(net16067), .Z(n2630) );
  CENXL U4772 ( .A(n4341), .B(net16067), .Z(n2616) );
  CENXL U4773 ( .A(n4330), .B(net16067), .Z(n2632) );
  CENXL U4774 ( .A(n4340), .B(net16067), .Z(n2617) );
  CENXL U4775 ( .A(n4335), .B(net16067), .Z(n2622) );
  CENXL U4776 ( .A(n4339), .B(net16067), .Z(n2618) );
  CNIVX4 U4777 ( .A(n2780), .Z(n4342) );
  CAOR1XL U4778 ( .A(net19508), .B(n4002), .C(n2648), .Z(n2121) );
  CENXL U4779 ( .A(n4338), .B(n4259), .Z(n2421) );
  CENXL U4780 ( .A(n4339), .B(n4259), .Z(n2420) );
  CENXL U4781 ( .A(n4340), .B(n4259), .Z(n2419) );
  CENXL U4782 ( .A(n4325), .B(n4259), .Z(n2441) );
  CENXL U4783 ( .A(net16544), .B(n4259), .Z(n2425) );
  COND2XL U4784 ( .A(n4260), .B(n2267), .C(n3576), .D(n2266), .Z(n1753) );
  COND2XL U4785 ( .A(n144), .B(n2260), .C(n3577), .D(n2259), .Z(n1746) );
  COND2XL U4786 ( .A(n4260), .B(n2261), .C(n3576), .D(n2260), .Z(n1747) );
  COND2XL U4787 ( .A(n144), .B(n2255), .C(n3576), .D(n2254), .Z(n800) );
  COND2XL U4788 ( .A(n2253), .B(n4260), .C(n3722), .D(n2252), .Z(n794) );
  COND2XL U4789 ( .A(n144), .B(n2257), .C(n3576), .D(n2256), .Z(n1743) );
  CND2XL U4790 ( .A(n1110), .B(n3333), .Z(n4104) );
  COND2XL U4791 ( .A(net18670), .B(n2547), .C(net16771), .D(n2546), .Z(n2020)
         );
  CND3X2 U4792 ( .A(n4127), .B(n4128), .C(n4129), .Z(n1186) );
  COND2X1 U4793 ( .A(n4261), .B(n2276), .C(n3577), .D(n2275), .Z(n1762) );
  CNR2IX1 U4794 ( .B(net16109), .A(n4295), .Z(n1863) );
  COND2XL U4795 ( .A(net18607), .B(n2487), .C(net19060), .D(n2486), .Z(n1962)
         );
  COND2XL U4796 ( .A(net18607), .B(n2490), .C(net19060), .D(n2489), .Z(n1965)
         );
  COND2XL U4797 ( .A(n2484), .B(net18607), .C(net19060), .D(n2483), .Z(n1959)
         );
  COND2XL U4798 ( .A(net18607), .B(n2486), .C(net19061), .D(n2485), .Z(n1961)
         );
  CNR2X2 U4799 ( .A(n3481), .B(n1412), .Z(n582) );
  CND2XL U4800 ( .A(n1277), .B(n1306), .Z(n4090) );
  CND2XL U4801 ( .A(n1306), .B(n1279), .Z(n4092) );
  CND3X1 U4802 ( .A(n4090), .B(n4091), .C(n4092), .Z(n1274) );
  CND2XL U4803 ( .A(n4169), .B(n1974), .Z(n4095) );
  CND2X2 U4804 ( .A(n4093), .B(n4094), .Z(n4096) );
  CND2X2 U4805 ( .A(n4095), .B(n4096), .Z(n1299) );
  CIVXL U4806 ( .A(n1974), .Z(n4094) );
  CND2X1 U4807 ( .A(n1299), .B(n1293), .Z(n4239) );
  CND2X2 U4808 ( .A(n4099), .B(n4100), .Z(n4162) );
  CNIVX4 U4809 ( .A(a[8]), .Z(n4102) );
  CENXL U4810 ( .A(n4331), .B(n4349), .Z(n2565) );
  CENXL U4811 ( .A(n4335), .B(n4000), .Z(n2556) );
  CENXL U4812 ( .A(net16550), .B(n4000), .Z(n2560) );
  COND1X1 U4813 ( .A(n697), .B(n693), .C(n694), .Z(n692) );
  CND2X1 U4814 ( .A(n1685), .B(n1692), .Z(n694) );
  CIVX4 U4815 ( .A(net19016), .Z(net16093) );
  CND2X2 U4816 ( .A(net19267), .B(net19268), .Z(n4103) );
  CIVX2 U4817 ( .A(net16083), .Z(net19267) );
  CIVX2 U4818 ( .A(a[6]), .Z(net19268) );
  CAOR1XL U4819 ( .A(net19500), .B(net19168), .C(n2549), .Z(n2022) );
  COND2XL U4820 ( .A(net19168), .B(n2572), .C(net19151), .D(n2571), .Z(n2045)
         );
  COND2XL U4821 ( .A(n4135), .B(n2579), .C(net19151), .D(n2578), .Z(n2052) );
  CND2XL U4822 ( .A(n3333), .B(n1112), .Z(n4106) );
  CND3X1 U4823 ( .A(n4104), .B(n4106), .C(n4105), .Z(n1084) );
  CENX2 U4824 ( .A(n1253), .B(n1251), .Z(n4107) );
  CNR2X2 U4825 ( .A(n1525), .B(n1544), .Z(n627) );
  CNIVX3 U4826 ( .A(n4233), .Z(n4289) );
  CENXL U4827 ( .A(n4341), .B(n4253), .Z(n2385) );
  CENXL U4828 ( .A(n4340), .B(n4253), .Z(n2386) );
  CENXL U4829 ( .A(n4339), .B(n4253), .Z(n2387) );
  CENXL U4830 ( .A(n4335), .B(n4253), .Z(n2391) );
  CENXL U4831 ( .A(n4337), .B(n4253), .Z(n2389) );
  CENXL U4832 ( .A(n4338), .B(n4253), .Z(n2388) );
  CIVX4 U4833 ( .A(n4252), .Z(n4253) );
  CIVXL U4834 ( .A(n3874), .Z(n4108) );
  CEOX1 U4835 ( .A(n1729), .B(n1925), .Z(n1543) );
  CND2X1 U4836 ( .A(n1136), .B(n1138), .Z(n4109) );
  CND2XL U4837 ( .A(n1138), .B(n1113), .Z(n4111) );
  CIVX1 U4838 ( .A(n4307), .Z(n4306) );
  CNR2X2 U4839 ( .A(n1159), .B(n1186), .Z(n522) );
  CND2X1 U4840 ( .A(n1159), .B(n1186), .Z(n523) );
  CAOR1XL U4841 ( .A(n4295), .B(n4033), .C(n2351), .Z(n1834) );
  COND2XL U4842 ( .A(n4033), .B(n2355), .C(n4295), .D(n2354), .Z(n1838) );
  COND2XL U4843 ( .A(n2352), .B(n4295), .C(n2353), .D(net19417), .Z(n1836) );
  COND2XL U4844 ( .A(n4033), .B(n2356), .C(n4295), .D(n2355), .Z(n864) );
  CENXL U4845 ( .A(n4339), .B(n3407), .Z(n2354) );
  CENXL U4846 ( .A(n4341), .B(n3407), .Z(n2352) );
  CENXL U4847 ( .A(n4338), .B(n3704), .Z(n2355) );
  CENXL U4848 ( .A(n4337), .B(n3704), .Z(n2356) );
  CENXL U4849 ( .A(n4336), .B(n3704), .Z(n2357) );
  CENXL U4850 ( .A(n4335), .B(n3704), .Z(n2358) );
  CENXL U4851 ( .A(n2789), .B(n3704), .Z(n2360) );
  CENXL U4852 ( .A(net16544), .B(n3704), .Z(n2359) );
  CENXL U4853 ( .A(net16548), .B(n3704), .Z(n2361) );
  CENXL U4854 ( .A(net16550), .B(n3704), .Z(n2362) );
  CENXL U4855 ( .A(n4325), .B(n3704), .Z(n2375) );
  CENXL U4856 ( .A(n4334), .B(n3704), .Z(n2363) );
  CENXL U4857 ( .A(n4330), .B(n3574), .Z(n2665) );
  CIVXL U4858 ( .A(n693), .Z(n784) );
  CNR2X2 U4859 ( .A(n1641), .B(n1652), .Z(n671) );
  CND2XL U4860 ( .A(n1475), .B(n1477), .Z(n4112) );
  CND2XL U4861 ( .A(n1475), .B(n1479), .Z(n4113) );
  CND2X1 U4862 ( .A(n1477), .B(n1479), .Z(n4114) );
  CEOX2 U4863 ( .A(n4115), .B(n3033), .Z(n1441) );
  CND2X1 U4864 ( .A(n3027), .B(n1447), .Z(n4116) );
  CND2X1 U4865 ( .A(n1445), .B(n1468), .Z(n4117) );
  CND3X2 U4866 ( .A(n4116), .B(n4117), .C(n4118), .Z(n1440) );
  CFA1X1 U4867 ( .A(n2144), .B(n1732), .CI(n2237), .CO(n1636), .S(n1637) );
  CND2XL U4868 ( .A(n641), .B(n3756), .Z(n193) );
  COND2X1 U4869 ( .A(net18670), .B(net18905), .C(net16771), .D(n2548), .Z(
        n1732) );
  CND2XL U4870 ( .A(n1311), .B(n1313), .Z(n4120) );
  CND2XL U4871 ( .A(n1336), .B(n1313), .Z(n4121) );
  CND3X1 U4872 ( .A(n4121), .B(n4120), .C(n4122), .Z(n1306) );
  CAOR1XL U4873 ( .A(n4017), .B(n3092), .C(n2615), .Z(n2088) );
  CND2X1 U4874 ( .A(n4216), .B(n4124), .Z(n4125) );
  CIVX2 U4875 ( .A(n4216), .Z(n4123) );
  CND3X1 U4876 ( .A(n4213), .B(n4214), .C(n4215), .Z(n1308) );
  CENX1 U4877 ( .A(n1265), .B(n1271), .Z(n4194) );
  COND2XL U4878 ( .A(n3877), .B(n2595), .C(net18731), .D(n2594), .Z(n2068) );
  CND2IXL U4879 ( .B(net16109), .A(net16063), .Z(n2614) );
  CENXL U4880 ( .A(n4325), .B(net16063), .Z(n2606) );
  CENXL U4881 ( .A(n4339), .B(net16063), .Z(n2585) );
  CENXL U4882 ( .A(net16558), .B(net16063), .Z(n2597) );
  CENXL U4883 ( .A(n4330), .B(net16063), .Z(n2599) );
  CENXL U4884 ( .A(n4331), .B(net16063), .Z(n2598) );
  CENXL U4885 ( .A(n4333), .B(net16063), .Z(n2595) );
  CND2XL U4886 ( .A(n1216), .B(n1191), .Z(n4129) );
  COND2X1 U4887 ( .A(n3606), .B(n2345), .C(net16802), .D(n2344), .Z(n1828) );
  CENX1 U4888 ( .A(n4324), .B(n4291), .Z(n2376) );
  CNIVX4 U4889 ( .A(n2788), .Z(net16544) );
  CND2XL U4890 ( .A(n2003), .B(n1914), .Z(n4130) );
  CND2XL U4891 ( .A(n1914), .B(n1884), .Z(n4132) );
  CND3X1 U4892 ( .A(n4130), .B(n4131), .C(n4132), .Z(n1266) );
  COR2XL U4893 ( .A(net16771), .B(n2529), .Z(n4134) );
  CENXL U4894 ( .A(n4332), .B(net18936), .Z(n2530) );
  CND2X2 U4895 ( .A(n4012), .B(net19500), .Z(n4135) );
  CND2X2 U4896 ( .A(n4012), .B(net19500), .Z(net19168) );
  CND2X2 U4897 ( .A(n2821), .B(net19500), .Z(n63) );
  CND2XL U4898 ( .A(n1300), .B(n1292), .Z(n4146) );
  CENXL U4899 ( .A(n2802), .B(n4347), .Z(n2670) );
  CENXL U4900 ( .A(n4333), .B(n4347), .Z(n2661) );
  CENXL U4901 ( .A(n4332), .B(n4347), .Z(n2662) );
  CENXL U4902 ( .A(n4329), .B(n4347), .Z(n2666) );
  CENX1 U4903 ( .A(n3036), .B(n4137), .Z(n1217) );
  CENX1 U4904 ( .A(n1250), .B(n1221), .Z(n4137) );
  CIVX1 U4905 ( .A(n84), .Z(net16759) );
  CENXL U4906 ( .A(net16558), .B(n4345), .Z(n2762) );
  CND2XL U4907 ( .A(n1213), .B(n1205), .Z(n4138) );
  CND2XL U4908 ( .A(n1213), .B(n1211), .Z(n4139) );
  CND3X1 U4909 ( .A(n4138), .B(n4140), .C(n4139), .Z(n1198) );
  CND2X4 U4910 ( .A(n2817), .B(net16812), .Z(n99) );
  CIVXL U4911 ( .A(n4345), .Z(n4142) );
  CNR2X2 U4912 ( .A(n540), .B(n543), .Z(n534) );
  CND2IX4 U4913 ( .B(n4187), .A(net16838), .Z(net19122) );
  CND2IXL U4914 ( .B(n4187), .A(net16839), .Z(n108) );
  CNIVX4 U4915 ( .A(n75), .Z(net18618) );
  CIVXL U4916 ( .A(n48), .Z(net16065) );
  CND2X1 U4917 ( .A(n1310), .B(n1285), .Z(n4177) );
  CIVXL U4918 ( .A(n4233), .Z(n4143) );
  CIVXL U4919 ( .A(n516), .Z(net19108) );
  CNIVX4 U4920 ( .A(net19401), .Z(net18936) );
  CND2XL U4921 ( .A(n1300), .B(n1298), .Z(n4147) );
  CND2XL U4922 ( .A(n1292), .B(n1298), .Z(n4148) );
  CND3X1 U4923 ( .A(n4146), .B(n4147), .C(n4148), .Z(n1258) );
  CIVXL U4924 ( .A(net18981), .Z(net19089) );
  CEO3X2 U4925 ( .A(n1532), .B(n1530), .C(n1515), .Z(n1509) );
  CND2XL U4926 ( .A(n1532), .B(n1530), .Z(n4149) );
  CND2XL U4927 ( .A(n1532), .B(n1515), .Z(n4150) );
  CND2X1 U4928 ( .A(n1530), .B(n1515), .Z(n4151) );
  CND2XL U4929 ( .A(n1491), .B(n1489), .Z(n4152) );
  CND2X1 U4930 ( .A(n1491), .B(n1508), .Z(n4153) );
  CND2XL U4931 ( .A(n1489), .B(n1508), .Z(n4154) );
  CND3X1 U4932 ( .A(n4152), .B(n4153), .C(n4154), .Z(n1484) );
  CIVX1 U4933 ( .A(n48), .Z(net19076) );
  CENX1 U4934 ( .A(net16544), .B(net16843), .Z(n2689) );
  COND2XL U4935 ( .A(net18743), .B(n2709), .C(net16772), .D(n2708), .Z(n2182)
         );
  COND2XL U4936 ( .A(n3024), .B(n2699), .C(net16772), .D(n2698), .Z(n2172) );
  COND2XL U4937 ( .A(net18743), .B(n2700), .C(net16772), .D(n2699), .Z(n2173)
         );
  COND2XL U4938 ( .A(net18743), .B(n2708), .C(net16772), .D(n2707), .Z(n2181)
         );
  COND2XL U4939 ( .A(n3024), .B(n2694), .C(net16772), .D(n2693), .Z(n2167) );
  COND2XL U4940 ( .A(n3024), .B(n2697), .C(net16772), .D(n2696), .Z(n2170) );
  CEO3X2 U4941 ( .A(n1876), .B(n1996), .C(n2026), .Z(n1051) );
  CND2XL U4942 ( .A(n2026), .B(n1996), .Z(n4156) );
  CND2XL U4943 ( .A(n2026), .B(n1876), .Z(n4157) );
  CND2XL U4944 ( .A(n1876), .B(n1996), .Z(n4158) );
  CND3X1 U4945 ( .A(n4156), .B(n4157), .C(n4158), .Z(n1050) );
  CND2XL U4946 ( .A(n1074), .B(n1072), .Z(n4159) );
  CND2X1 U4947 ( .A(n1074), .B(n1051), .Z(n4160) );
  CND2X1 U4948 ( .A(n1072), .B(n1051), .Z(n4161) );
  CND3X2 U4949 ( .A(n4159), .B(n4160), .C(n4161), .Z(n1046) );
  CIVX4 U4950 ( .A(net18817), .Z(net16069) );
  CIVXL U4951 ( .A(n3700), .Z(n676) );
  CENX4 U4952 ( .A(a[24]), .B(n4354), .Z(net16784) );
  CND2XL U4953 ( .A(n1217), .B(n1219), .Z(n4249) );
  CENXL U4954 ( .A(n574), .B(n184), .Z(product[28]) );
  CEOX2 U4955 ( .A(n3176), .B(n4162), .Z(n1159) );
  CND2XL U4956 ( .A(n3176), .B(n4021), .Z(n4163) );
  CND2XL U4957 ( .A(n4021), .B(n1163), .Z(n4165) );
  CND2XL U4958 ( .A(n2188), .B(n1767), .Z(n4166) );
  CND3X1 U4959 ( .A(n4166), .B(n4167), .C(n4168), .Z(n1240) );
  CENX1 U4960 ( .A(n2159), .B(n2190), .Z(n4169) );
  CIVX1 U4961 ( .A(n425), .Z(n423) );
  CND2X4 U4962 ( .A(n2812), .B(n4294), .Z(n144) );
  CNR2X2 U4963 ( .A(n444), .B(n460), .Z(n438) );
  CENX2 U4964 ( .A(net18817), .B(n4101), .Z(n2823) );
  CIVX4 U4965 ( .A(net18817), .Z(net16067) );
  CENX2 U4966 ( .A(a[14]), .B(n4308), .Z(n4233) );
  CENXL U4967 ( .A(n4336), .B(net16067), .Z(n2621) );
  CENXL U4968 ( .A(n4341), .B(n3889), .Z(n2451) );
  CENXL U4969 ( .A(n4338), .B(n3889), .Z(n2454) );
  CENXL U4970 ( .A(n4340), .B(n3889), .Z(n2452) );
  CENXL U4971 ( .A(n4339), .B(n3889), .Z(n2453) );
  CENXL U4972 ( .A(n2789), .B(n3487), .Z(n2459) );
  CENXL U4973 ( .A(net16544), .B(n3487), .Z(n2458) );
  CENXL U4974 ( .A(n4325), .B(n3486), .Z(n2474) );
  CENXL U4975 ( .A(n4335), .B(n3889), .Z(n2457) );
  CENXL U4976 ( .A(net16550), .B(n3486), .Z(n2461) );
  CENXL U4977 ( .A(n4337), .B(n3487), .Z(n2455) );
  CENXL U4978 ( .A(n4336), .B(n3486), .Z(n2456) );
  CENXL U4979 ( .A(n4334), .B(n3889), .Z(n2462) );
  CENXL U4980 ( .A(net16548), .B(n3486), .Z(n2460) );
  COND2X1 U4981 ( .A(n2649), .B(net16791), .C(n2650), .D(n4003), .Z(n2123) );
  CND2X1 U4982 ( .A(n2820), .B(n4233), .Z(n72) );
  CNIVX4 U4983 ( .A(n2786), .Z(n4336) );
  CND2X2 U4984 ( .A(n4266), .B(n4265), .Z(n105) );
  CND2IXL U4985 ( .B(net16109), .A(n4253), .Z(n2416) );
  CENXL U4986 ( .A(net16544), .B(n4362), .Z(n2260) );
  CENXL U4987 ( .A(n2789), .B(n4262), .Z(n2261) );
  CENXL U4988 ( .A(n4336), .B(n4362), .Z(n2258) );
  CENXL U4989 ( .A(n4335), .B(n4262), .Z(n2259) );
  CENXL U4990 ( .A(net16548), .B(n4362), .Z(n2262) );
  CENXL U4991 ( .A(net16550), .B(n4362), .Z(n2263) );
  CENXL U4992 ( .A(n4332), .B(n4262), .Z(n2266) );
  CENXL U4993 ( .A(n4333), .B(n4262), .Z(n2265) );
  CENXL U4994 ( .A(n4334), .B(n4262), .Z(n2264) );
  CENXL U4995 ( .A(net16558), .B(n4262), .Z(n2267) );
  CENXL U4996 ( .A(n4331), .B(n4262), .Z(n2268) );
  CENXL U4997 ( .A(n4330), .B(n4262), .Z(n2269) );
  CENXL U4998 ( .A(n4329), .B(n4262), .Z(n2270) );
  CENX1 U4999 ( .A(n2808), .B(n4262), .Z(n2280) );
  CNIVX4 U5000 ( .A(a[8]), .Z(n4171) );
  CIVX4 U5001 ( .A(n3486), .Z(net16849) );
  CEOX4 U5002 ( .A(n4362), .B(a[30]), .Z(n2812) );
  CENX1 U5003 ( .A(n4194), .B(n1269), .Z(n1257) );
  CENXL U5004 ( .A(n604), .B(n187), .Z(product[25]) );
  CIVXL U5005 ( .A(n4053), .Z(n4173) );
  COR2X1 U5006 ( .A(n4205), .B(n1281), .Z(n4206) );
  CIVX1 U5007 ( .A(n1283), .Z(n4205) );
  CENXL U5008 ( .A(n4338), .B(net16067), .Z(n2619) );
  COND2XL U5009 ( .A(n3963), .B(n2620), .C(net16793), .D(n2619), .Z(n2093) );
  COND1X1 U5010 ( .A(n416), .B(n4020), .C(n3268), .Z(n415) );
  CANR1X1 U5011 ( .A(n739), .B(n308), .C(n301), .Z(n299) );
  CIVXL U5012 ( .A(net16089), .Z(net18948) );
  CENXL U5013 ( .A(n176), .B(n513), .Z(product[36]) );
  CENXL U5014 ( .A(n177), .B(n524), .Z(product[35]) );
  COND1X1 U5015 ( .A(n392), .B(n365), .C(n366), .Z(n364) );
  CENXL U5016 ( .A(n4331), .B(net16037), .Z(n4174) );
  CENXL U5017 ( .A(n178), .B(n531), .Z(product[34]) );
  CENXL U5018 ( .A(n179), .B(n542), .Z(product[33]) );
  CENXL U5019 ( .A(n174), .B(n495), .Z(product[38]) );
  CENXL U5020 ( .A(n175), .B(n506), .Z(product[37]) );
  CNIVX4 U5021 ( .A(n2800), .Z(n4327) );
  CEO3X2 U5022 ( .A(n1312), .B(n1285), .C(n1310), .Z(n1279) );
  CND3X1 U5023 ( .A(n4182), .B(n4181), .C(n4180), .Z(n1246) );
  COND2X1 U5024 ( .A(n144), .B(n2281), .C(n3576), .D(n2280), .Z(n1767) );
  CND2IX1 U5025 ( .B(n4241), .A(n4186), .Z(n2035) );
  COR2XL U5026 ( .A(net19500), .B(n2561), .Z(n4186) );
  CND2IX4 U5027 ( .B(n4187), .A(net16838), .Z(n4188) );
  CENXL U5028 ( .A(n4330), .B(net16037), .Z(n4189) );
  CENXL U5029 ( .A(n459), .B(n170), .Z(product[42]) );
  CENXL U5030 ( .A(n435), .B(n168), .Z(product[44]) );
  CENXL U5031 ( .A(n411), .B(n166), .Z(product[46]) );
  CENXL U5032 ( .A(n393), .B(n164), .Z(product[48]) );
  CENXL U5033 ( .A(n343), .B(n160), .Z(product[52]) );
  CENXL U5034 ( .A(n317), .B(n158), .Z(product[54]) );
  CAOR1XL U5035 ( .A(net16801), .B(n3607), .C(n2318), .Z(n1803) );
  COND2XL U5036 ( .A(n2319), .B(net16801), .C(n2320), .D(n3607), .Z(n1805) );
  COND2XL U5037 ( .A(n3607), .B(n2324), .C(net16801), .D(n2323), .Z(n1807) );
  COND2XL U5038 ( .A(n3606), .B(n2329), .C(net16801), .D(n2328), .Z(n1812) );
  COND2XL U5039 ( .A(n3607), .B(n2338), .C(net16801), .D(n2337), .Z(n1821) );
  CNR2IX1 U5040 ( .B(net16109), .A(net16801), .Z(n1833) );
  CIVXL U5041 ( .A(n4254), .Z(n4190) );
  CND2XL U5042 ( .A(n1203), .B(n1226), .Z(n4246) );
  CENXL U5043 ( .A(n4322), .B(n4145), .Z(n2576) );
  CENXL U5044 ( .A(n4323), .B(n4349), .Z(n2575) );
  CENXL U5045 ( .A(n4326), .B(n4306), .Z(n2572) );
  CENXL U5046 ( .A(n4342), .B(n4145), .Z(n2549) );
  CENXL U5047 ( .A(n2802), .B(n4000), .Z(n2571) );
  CENXL U5048 ( .A(n4321), .B(n4000), .Z(n2578) );
  CENXL U5049 ( .A(net16558), .B(n4000), .Z(n2564) );
  CENXL U5050 ( .A(net16570), .B(n4145), .Z(n2570) );
  CND2X4 U5051 ( .A(n2817), .B(net16812), .Z(net18897) );
  CENXL U5052 ( .A(n4342), .B(n4343), .Z(n2747) );
  CND2XL U5053 ( .A(n1221), .B(n1250), .Z(n4193) );
  CENXL U5054 ( .A(n4326), .B(net18643), .Z(n2539) );
  CENXL U5055 ( .A(n4327), .B(net18643), .Z(n2536) );
  CENXL U5056 ( .A(n2810), .B(net18936), .Z(n2546) );
  CENXL U5057 ( .A(n4328), .B(net18936), .Z(n2535) );
  CENXL U5058 ( .A(net16570), .B(net18937), .Z(n2537) );
  CENXL U5059 ( .A(n4323), .B(net18643), .Z(n2542) );
  CNIVX4 U5060 ( .A(n4347), .Z(n4255) );
  CANR1XL U5061 ( .A(n3756), .B(n3411), .C(n639), .Z(n4195) );
  COND1X1 U5062 ( .A(n678), .B(n690), .C(n679), .Z(n677) );
  CIVXL U5063 ( .A(n690), .Z(n689) );
  CND2XL U5064 ( .A(n1085), .B(n3132), .Z(n4223) );
  CAOR1XL U5065 ( .A(n6), .B(net19555), .C(n2747), .Z(n2220) );
  CND2XL U5066 ( .A(net18875), .B(n2010), .Z(n4196) );
  CND2XL U5067 ( .A(net18875), .B(n1950), .Z(n4197) );
  CND3X1 U5068 ( .A(n4196), .B(n4197), .C(n4198), .Z(n1452) );
  CND2XL U5069 ( .A(n1455), .B(n1457), .Z(n4199) );
  CND2XL U5070 ( .A(n1455), .B(n1453), .Z(n4200) );
  CND2XL U5071 ( .A(n1457), .B(n1453), .Z(n4201) );
  CND3X1 U5072 ( .A(n4199), .B(n4200), .C(n4201), .Z(n1444) );
  CND2XL U5073 ( .A(n1974), .B(n2190), .Z(n4202) );
  CND2XL U5074 ( .A(n1974), .B(n2159), .Z(n4203) );
  CND2XL U5075 ( .A(n2190), .B(n2159), .Z(n4204) );
  CND2X2 U5076 ( .A(n4206), .B(n4207), .Z(n4216) );
  CNR2XL U5077 ( .A(n81), .B(n2500), .Z(n4208) );
  CNR2XL U5078 ( .A(net19060), .B(n2499), .Z(n4209) );
  COR2X1 U5079 ( .A(n4208), .B(n4209), .Z(n1974) );
  CENXL U5080 ( .A(n4330), .B(net16037), .Z(n2500) );
  CENXL U5081 ( .A(n4331), .B(net16037), .Z(n2499) );
  CND2X1 U5082 ( .A(n1345), .B(n1370), .Z(n4210) );
  CND2X1 U5083 ( .A(n1345), .B(n1347), .Z(n4211) );
  CND2X1 U5084 ( .A(n1370), .B(n1347), .Z(n4212) );
  CND3X2 U5085 ( .A(n4210), .B(n4211), .C(n4212), .Z(n1338) );
  CEO3X2 U5086 ( .A(n1315), .B(n1338), .C(n1340), .Z(n1309) );
  CND2XL U5087 ( .A(n1315), .B(n1338), .Z(n4213) );
  CND2XL U5088 ( .A(n1315), .B(n1340), .Z(n4214) );
  CND2XL U5089 ( .A(n1283), .B(n1281), .Z(n4217) );
  CND2XL U5090 ( .A(n1281), .B(n1308), .Z(n4219) );
  CEO3X2 U5091 ( .A(n2225), .B(n2039), .C(n3800), .Z(n1409) );
  COND1X1 U5092 ( .A(n309), .B(net19530), .C(n310), .Z(n308) );
  CENXL U5093 ( .A(n4341), .B(n3219), .Z(n4221) );
  CIVXL U5094 ( .A(net19292), .Z(n590) );
  CND2X1 U5095 ( .A(n1107), .B(n1132), .Z(n505) );
  COND2X1 U5096 ( .A(n81), .B(n2503), .C(net19060), .D(n2502), .Z(n1977) );
  CND2XL U5097 ( .A(n1085), .B(n1108), .Z(n4222) );
  CNR2X1 U5098 ( .A(n3405), .B(n1059), .Z(n4225) );
  CEOX2 U5099 ( .A(n4226), .B(n1377), .Z(n1371) );
  CND2XL U5100 ( .A(n1377), .B(n1381), .Z(n4227) );
  CND2XL U5101 ( .A(n1377), .B(n1383), .Z(n4228) );
  CND2XL U5102 ( .A(n1381), .B(n1383), .Z(n4229) );
  CEO3X2 U5103 ( .A(n2100), .B(n2038), .C(n1977), .Z(n1377) );
  CND2XL U5104 ( .A(n2100), .B(n1977), .Z(n4230) );
  CND2XL U5105 ( .A(n2100), .B(n2038), .Z(n4231) );
  CND2XL U5106 ( .A(n1977), .B(n2038), .Z(n4232) );
  COND2X1 U5107 ( .A(n36), .B(n2651), .C(net19508), .D(n2650), .Z(n2124) );
  CENXL U5108 ( .A(n4334), .B(net16067), .Z(n2627) );
  CND2XL U5109 ( .A(n3136), .B(n485), .Z(n173) );
  CND2XL U5110 ( .A(n3061), .B(n661), .Z(n196) );
  CANR1X2 U5111 ( .A(n3874), .B(n4267), .C(n601), .Z(n595) );
  CIVDX2 U5112 ( .A(n4350), .Z0(n4308), .Z1(n4307) );
  COND2X1 U5113 ( .A(n2748), .B(n6), .C(n2749), .D(n9), .Z(n2222) );
  CENXL U5114 ( .A(n4342), .B(n3796), .Z(n2285) );
  CENXL U5115 ( .A(n4328), .B(n3152), .Z(n2304) );
  CENXL U5116 ( .A(net16570), .B(n3152), .Z(n2306) );
  CENXL U5117 ( .A(n4327), .B(n3151), .Z(n2305) );
  CENXL U5118 ( .A(n2802), .B(n4251), .Z(n2307) );
  CENXL U5119 ( .A(n4324), .B(n3152), .Z(n2310) );
  CENXL U5120 ( .A(n4322), .B(n3151), .Z(n2312) );
  CENXL U5121 ( .A(n4321), .B(n3151), .Z(n2314) );
  CENXL U5122 ( .A(n2810), .B(n3151), .Z(n2315) );
  CENXL U5123 ( .A(n2808), .B(n3152), .Z(n2313) );
  CEO3X2 U5124 ( .A(n1885), .B(n1944), .C(n2035), .Z(n1293) );
  CND2XL U5125 ( .A(n1885), .B(n1944), .Z(n4235) );
  CND2X1 U5126 ( .A(n1885), .B(n2035), .Z(n4236) );
  CND2X1 U5127 ( .A(n1944), .B(n2035), .Z(n4237) );
  CND3X2 U5128 ( .A(n4235), .B(n4236), .C(n4237), .Z(n1292) );
  CND2XL U5129 ( .A(n1301), .B(n1299), .Z(n4238) );
  CND2XL U5130 ( .A(n1301), .B(n1293), .Z(n4240) );
  CND3X1 U5131 ( .A(n4238), .B(n4240), .C(n4239), .Z(n1286) );
  CNR2XL U5132 ( .A(n2562), .B(net19168), .Z(n4241) );
  CIVXL U5133 ( .A(n491), .Z(n756) );
  CND3X1 U5134 ( .A(n4318), .B(n4319), .C(n4320), .Z(n1106) );
  CENXL U5135 ( .A(n297), .B(n156), .Z(product[56]) );
  CIVXL U5136 ( .A(n3839), .Z(net18730) );
  CIVX4 U5137 ( .A(n4356), .Z(n4354) );
  CFA1X1 U5138 ( .A(n1242), .B(n1766), .CI(n2156), .CO(n1212), .S(n1213) );
  CENXL U5139 ( .A(n4342), .B(n4291), .Z(n2351) );
  COND1X2 U5140 ( .A(n633), .B(n637), .C(n634), .Z(n632) );
  CENXL U5141 ( .A(net16558), .B(n4347), .Z(n2663) );
  CENXL U5142 ( .A(n4331), .B(n3574), .Z(n2664) );
  CEO3X1 U5143 ( .A(n1262), .B(n1233), .C(n1239), .Z(n1227) );
  CND2X1 U5144 ( .A(n1233), .B(n3417), .Z(n4242) );
  CND2XL U5145 ( .A(n3417), .B(n1239), .Z(n4243) );
  CND2X1 U5146 ( .A(n1233), .B(n1239), .Z(n4244) );
  CND2XL U5147 ( .A(n1228), .B(n1226), .Z(n4247) );
  CND2XL U5148 ( .A(n1217), .B(n4054), .Z(n4248) );
  CND2XL U5149 ( .A(n4054), .B(n1219), .Z(n4250) );
  CND3X1 U5150 ( .A(n4248), .B(n4249), .C(n4250), .Z(n1214) );
  CENX1 U5151 ( .A(n3714), .B(n1801), .Z(n1359) );
  CND2X1 U5152 ( .A(n1158), .B(n1133), .Z(n512) );
  CNR2X1 U5153 ( .A(n1158), .B(n1133), .Z(n511) );
  CENXL U5154 ( .A(n4321), .B(net16069), .Z(n2644) );
  CNIVX4 U5155 ( .A(n2806), .Z(n4323) );
  CNR2X2 U5156 ( .A(n4225), .B(n491), .Z(n482) );
  CENX4 U5157 ( .A(a[30]), .B(n3151), .Z(n141) );
  CANR1X2 U5158 ( .A(n753), .B(n3602), .C(n467), .Z(n461) );
  CENXL U5159 ( .A(n4341), .B(n4000), .Z(n2550) );
  CENXL U5160 ( .A(net16109), .B(n4306), .Z(n2580) );
  CENXL U5161 ( .A(n4337), .B(n4000), .Z(n2554) );
  CENXL U5162 ( .A(n4325), .B(n4000), .Z(n2573) );
  CENXL U5163 ( .A(n2810), .B(n4000), .Z(n2579) );
  CENXL U5164 ( .A(n2789), .B(n4306), .Z(n2558) );
  CENXL U5165 ( .A(n4334), .B(n4306), .Z(n2561) );
  CENXL U5166 ( .A(net16548), .B(n4349), .Z(n2559) );
  CENXL U5167 ( .A(n163), .B(n380), .Z(product[49]) );
  CENXL U5168 ( .A(n162), .B(n371), .Z(product[50]) );
  CENXL U5169 ( .A(n171), .B(n470), .Z(product[41]) );
  CENXL U5170 ( .A(n450), .B(n169), .Z(product[43]) );
  CENXL U5171 ( .A(n426), .B(n167), .Z(product[45]) );
  CENXL U5172 ( .A(n404), .B(n165), .Z(product[47]) );
  CENXL U5173 ( .A(n352), .B(n161), .Z(product[51]) );
  CENXL U5174 ( .A(n328), .B(n159), .Z(product[53]) );
  CNR2IX1 U5175 ( .B(net16109), .A(n3577), .Z(n1770) );
  CNIVX4 U5176 ( .A(n72), .Z(net18670) );
  CANR1X2 U5177 ( .A(n3411), .B(n4274), .C(n639), .Z(n637) );
  CENXL U5178 ( .A(net16107), .B(net16093), .Z(n2745) );
  CENXL U5179 ( .A(net16107), .B(n4344), .Z(n2778) );
  CENXL U5180 ( .A(net16107), .B(net16069), .Z(n2646) );
  CENXL U5181 ( .A(net16107), .B(net18643), .Z(n2547) );
  CENXL U5182 ( .A(net16107), .B(net16850), .Z(n2481) );
  CENXL U5183 ( .A(net16107), .B(n3730), .Z(n2613) );
  CENXL U5184 ( .A(net16107), .B(n4291), .Z(n2382) );
  CENXL U5185 ( .A(net16107), .B(n4292), .Z(n2448) );
  CENXL U5186 ( .A(net16107), .B(n4362), .Z(n2283) );
  COND1X1 U5187 ( .A(n248), .B(net19409), .C(n249), .Z(n247) );
  CNR2X1 U5188 ( .A(n1596), .B(n1581), .Z(n643) );
  CNR2X2 U5189 ( .A(n1613), .B(n1626), .Z(n660) );
  CENX1 U5190 ( .A(n4335), .B(net16844), .Z(n2688) );
  CENX1 U5191 ( .A(n4336), .B(net16844), .Z(n2687) );
  CENXL U5192 ( .A(n4342), .B(n4004), .Z(n2384) );
  CENXL U5193 ( .A(net16107), .B(n4004), .Z(n2415) );
  CENXL U5194 ( .A(n4323), .B(n3308), .Z(n2410) );
  CENXL U5195 ( .A(n4322), .B(n3308), .Z(n2411) );
  CENXL U5196 ( .A(n2808), .B(n3173), .Z(n2412) );
  CENXL U5197 ( .A(n4321), .B(n3058), .Z(n2413) );
  CENXL U5198 ( .A(n4324), .B(n3058), .Z(n2409) );
  CENXL U5199 ( .A(n4327), .B(n3173), .Z(n2404) );
  CENXL U5200 ( .A(n4328), .B(n4354), .Z(n2403) );
  CENXL U5201 ( .A(net16570), .B(n3173), .Z(n2405) );
  CND2X2 U5202 ( .A(n3872), .B(n3822), .Z(n90) );
  CND2X4 U5203 ( .A(n3328), .B(n3277), .Z(net18592) );
  CND2X4 U5204 ( .A(n2818), .B(n3822), .Z(net18593) );
  CENXL U5205 ( .A(net16107), .B(n3796), .Z(n2316) );
  CENXL U5206 ( .A(n4326), .B(n3152), .Z(n2308) );
  CENXL U5207 ( .A(net16107), .B(n4255), .Z(n2679) );
  CENXL U5208 ( .A(n4323), .B(n3574), .Z(n2674) );
  CENXL U5209 ( .A(n4324), .B(n4347), .Z(n2673) );
  CENXL U5210 ( .A(n2810), .B(n3574), .Z(n2678) );
  CENXL U5211 ( .A(n4327), .B(n3574), .Z(n2668) );
  CENXL U5212 ( .A(n2808), .B(n4347), .Z(n2676) );
  CENXL U5213 ( .A(n4321), .B(n3574), .Z(n2677) );
  CENXL U5214 ( .A(net16570), .B(n3574), .Z(n2669) );
  CENXL U5215 ( .A(n4328), .B(n3574), .Z(n2667) );
  CENXL U5216 ( .A(n4322), .B(n3574), .Z(n2675) );
  CENXL U5217 ( .A(n4342), .B(n4347), .Z(n2648) );
  CENXL U5218 ( .A(n4326), .B(n3574), .Z(n2671) );
  CENXL U5219 ( .A(n4341), .B(n4343), .Z(n2748) );
  CENXL U5220 ( .A(n4339), .B(n4343), .Z(n2750) );
  CENXL U5221 ( .A(n2808), .B(net16843), .Z(n2709) );
  CENXL U5222 ( .A(n4321), .B(net18948), .Z(n2710) );
  CENXL U5223 ( .A(net16109), .B(net18948), .Z(n2712) );
  CENXL U5224 ( .A(n4324), .B(net18982), .Z(n2706) );
  CENXL U5225 ( .A(n2810), .B(net18948), .Z(n2711) );
  CENXL U5226 ( .A(n4323), .B(net16844), .Z(n2707) );
  CENXL U5227 ( .A(n4322), .B(net18982), .Z(n2708) );
  CENXL U5228 ( .A(n4328), .B(net18982), .Z(n2700) );
  CENXL U5229 ( .A(n4342), .B(net18982), .Z(n2681) );
  CENXL U5230 ( .A(net16570), .B(net18982), .Z(n2702) );
  CND2X4 U5231 ( .A(n2819), .B(n3867), .Z(net18607) );
  CND2X4 U5232 ( .A(n4256), .B(n4257), .Z(n2819) );
  CIVX1 U5233 ( .A(n4264), .Z(n4259) );
  CIVX3 U5234 ( .A(n4264), .Z(n4351) );
  CENXL U5235 ( .A(n205), .B(n707), .Z(product[7]) );
  COR2XL U5236 ( .A(n2250), .B(n2219), .Z(n4286) );
  COND2X1 U5237 ( .A(n4001), .B(n2742), .C(net16816), .D(n2741), .Z(n2215) );
  COND2X1 U5238 ( .A(n2316), .B(n4136), .C(n3709), .D(n2315), .Z(n1801) );
  CND2X4 U5239 ( .A(n2812), .B(n4294), .Z(n4260) );
  CND2X1 U5240 ( .A(n799), .B(n802), .Z(n255) );
  CNIVX4 U5241 ( .A(n105), .Z(net16838) );
  CANR1XL U5242 ( .A(n3713), .B(n323), .C(n314), .Z(n310) );
  COAN1X1 U5243 ( .A(n327), .B(n291), .C(n292), .Z(n4273) );
  CANR1X1 U5244 ( .A(n4283), .B(n707), .C(n704), .Z(n702) );
  COND2X1 U5245 ( .A(n3092), .B(n2643), .C(net16793), .D(n2642), .Z(n2116) );
  CND2XL U5246 ( .A(n93), .B(a[22]), .Z(n4265) );
  CND2X2 U5247 ( .A(net19316), .B(n767), .Z(n578) );
  CND2XL U5248 ( .A(n355), .B(n331), .Z(n329) );
  CND2X1 U5249 ( .A(n879), .B(n892), .Z(n379) );
  CND2XL U5250 ( .A(n786), .B(n701), .Z(n204) );
  CND2X1 U5251 ( .A(n827), .B(n834), .Z(n316) );
  CENX1 U5252 ( .A(n208), .B(n721), .Z(product[4]) );
  CENX1 U5253 ( .A(n4339), .B(net16844), .Z(n2684) );
  CENX1 U5254 ( .A(n4342), .B(n4292), .Z(n2417) );
  COND2XL U5255 ( .A(net18743), .B(net18981), .C(net16772), .D(n2713), .Z(
        n1737) );
  CNIVX8 U5256 ( .A(n2809), .Z(n4321) );
  COND2X1 U5257 ( .A(n36), .B(n2668), .C(net16791), .D(n2667), .Z(n2141) );
  CND2XL U5258 ( .A(n516), .B(n758), .Z(n507) );
  CND2XL U5259 ( .A(n3320), .B(n458), .Z(n170) );
  CND2X2 U5260 ( .A(n4268), .B(n751), .Z(n444) );
  CENXL U5261 ( .A(n593), .B(n186), .Z(product[26]) );
  CND2XL U5262 ( .A(n746), .B(n392), .Z(n164) );
  CND2XL U5263 ( .A(n3175), .B(n4276), .Z(n168) );
  CND2XL U5264 ( .A(n4275), .B(n351), .Z(n161) );
  CND2XL U5265 ( .A(n747), .B(n403), .Z(n165) );
  CND2XL U5266 ( .A(n383), .B(n3267), .Z(n372) );
  CEOXL U5267 ( .A(n196), .B(n662), .Z(product[16]) );
  CEOXL U5268 ( .A(n195), .B(n657), .Z(product[17]) );
  CND2XL U5269 ( .A(n4277), .B(n656), .Z(n195) );
  CNR2XL U5270 ( .A(n1461), .B(n1482), .Z(n605) );
  CND2XL U5271 ( .A(n3980), .B(n623), .Z(n190) );
  CANR1X1 U5272 ( .A(n699), .B(n691), .C(n692), .Z(n690) );
  CNR2XL U5273 ( .A(n693), .B(n696), .Z(n691) );
  COND1X1 U5274 ( .A(n700), .B(n702), .C(n701), .Z(n699) );
  CND2XL U5275 ( .A(n4281), .B(n4280), .Z(n678) );
  CND2XL U5276 ( .A(n738), .B(n296), .Z(n156) );
  CND2XL U5277 ( .A(n355), .B(n320), .Z(n318) );
  CND2XL U5278 ( .A(n355), .B(n4275), .Z(n344) );
  CND2XL U5279 ( .A(n4279), .B(n342), .Z(n160) );
  CND2XL U5280 ( .A(n741), .B(n327), .Z(n159) );
  CND2XL U5281 ( .A(n355), .B(n283), .Z(n281) );
  CND2XL U5282 ( .A(n4282), .B(n279), .Z(n155) );
  CEOXL U5283 ( .A(n200), .B(n684), .Z(product[12]) );
  CND2XL U5284 ( .A(n4281), .B(n683), .Z(n200) );
  CND2XL U5285 ( .A(n781), .B(n675), .Z(n199) );
  CND2XL U5286 ( .A(n785), .B(n697), .Z(n203) );
  CEOXL U5287 ( .A(n702), .B(n204), .Z(product[8]) );
  CND2XL U5288 ( .A(n4280), .B(n688), .Z(n201) );
  CANR1X1 U5289 ( .A(n729), .B(n4286), .C(n726), .Z(n724) );
  CND2XL U5290 ( .A(n355), .B(n272), .Z(n268) );
  CENXL U5291 ( .A(n247), .B(n152), .Z(product[60]) );
  CND2XL U5292 ( .A(net18422), .B(n246), .Z(n152) );
  CND2XL U5293 ( .A(n1701), .B(n1706), .Z(n701) );
  COND1X1 U5294 ( .A(n261), .B(n3777), .C(n262), .Z(n260) );
  CIVX1 U5295 ( .A(n266), .Z(n264) );
  CND2XL U5296 ( .A(n4283), .B(n706), .Z(n205) );
  CND2XL U5297 ( .A(n4286), .B(n728), .Z(n210) );
  CND2XL U5298 ( .A(n4285), .B(n720), .Z(n208) );
  CND2XL U5299 ( .A(n4284), .B(n714), .Z(n207) );
  CND2XL U5300 ( .A(n1713), .B(n1716), .Z(n709) );
  CND2XL U5301 ( .A(n1723), .B(n2218), .Z(n723) );
  COND2XL U5302 ( .A(n2646), .B(n3092), .C(net16793), .D(n2645), .Z(n2119) );
  CNR2IX1 U5303 ( .B(net16109), .A(net16772), .Z(n2186) );
  CENXL U5304 ( .A(n4328), .B(n4352), .Z(n2436) );
  COND2XL U5305 ( .A(n4002), .B(n2656), .C(net19508), .D(n2655), .Z(n2129) );
  CENXL U5306 ( .A(n4340), .B(n3704), .Z(n2353) );
  CANR1XL U5307 ( .A(n3499), .B(n4053), .C(net19522), .Z(n497) );
  CND2XL U5308 ( .A(n534), .B(n3717), .Z(n525) );
  CND2XL U5309 ( .A(n3499), .B(n516), .Z(n496) );
  CND2XL U5310 ( .A(n489), .B(n516), .Z(n487) );
  CANR1XL U5311 ( .A(n758), .B(n4053), .C(n510), .Z(n508) );
  CANR1XL U5312 ( .A(n489), .B(n4053), .C(n490), .Z(n488) );
  CANR1XL U5313 ( .A(n3320), .B(n4019), .C(n456), .Z(n452) );
  CND2XL U5314 ( .A(n753), .B(n469), .Z(n171) );
  COND1XL U5315 ( .A(n3282), .B(net18543), .C(n3670), .Z(n470) );
  CND2XL U5316 ( .A(n751), .B(n449), .Z(n169) );
  COND1XL U5317 ( .A(n507), .B(n3731), .C(n508), .Z(n506) );
  COND1XL U5318 ( .A(n496), .B(n3731), .C(n497), .Z(n495) );
  CND2XL U5319 ( .A(n3131), .B(n3528), .Z(n179) );
  COND1XL U5320 ( .A(n543), .B(n3731), .C(n3068), .Z(n542) );
  CND2XL U5321 ( .A(n530), .B(n3717), .Z(n178) );
  COND1XL U5322 ( .A(n532), .B(n3731), .C(n4309), .Z(n531) );
  CND2XL U5323 ( .A(n512), .B(n758), .Z(n176) );
  COND1XL U5324 ( .A(net19108), .B(n3731), .C(n4173), .Z(n513) );
  CND2XL U5325 ( .A(n3060), .B(net19292), .Z(n186) );
  CND2X1 U5326 ( .A(n4267), .B(n603), .Z(n187) );
  COND1XL U5327 ( .A(n3933), .B(n611), .C(n3108), .Z(n604) );
  CND2XL U5328 ( .A(n3881), .B(n596), .Z(n585) );
  CANR1XL U5329 ( .A(n766), .B(n574), .C(n571), .Z(n569) );
  CANR1XL U5330 ( .A(net19307), .B(n574), .C(net19388), .Z(n560) );
  CANR1XL U5331 ( .A(n620), .B(n629), .C(n621), .Z(n619) );
  CND2X1 U5332 ( .A(n387), .B(n418), .Z(n385) );
  CANR1XL U5333 ( .A(n3060), .B(n597), .C(n590), .Z(n586) );
  CANR1XL U5334 ( .A(n3267), .B(n384), .C(n377), .Z(n373) );
  CND2XL U5335 ( .A(n3129), .B(n425), .Z(n167) );
  CND2XL U5336 ( .A(n3281), .B(n4276), .Z(n427) );
  CND2XL U5337 ( .A(n748), .B(n410), .Z(n166) );
  COND1XL U5338 ( .A(n525), .B(n3731), .C(n526), .Z(n524) );
  CNR2X1 U5339 ( .A(n660), .B(n665), .Z(n658) );
  CND2XL U5340 ( .A(n744), .B(n370), .Z(n162) );
  CND2XL U5341 ( .A(n3267), .B(n379), .Z(n163) );
  COND1XL U5342 ( .A(n381), .B(net18543), .C(n3133), .Z(n380) );
  COR2X1 U5343 ( .A(n995), .B(n1014), .Z(n4268) );
  CND2X1 U5344 ( .A(n3261), .B(n1058), .Z(n472) );
  CND2X1 U5345 ( .A(n995), .B(n1014), .Z(n458) );
  CND2X1 U5346 ( .A(n1437), .B(n1460), .Z(n603) );
  CND2X1 U5347 ( .A(n1483), .B(n1504), .Z(n618) );
  CND2X1 U5348 ( .A(n1059), .B(n1082), .Z(n485) );
  CND2X1 U5349 ( .A(n3481), .B(n1412), .Z(n583) );
  CND2XL U5350 ( .A(n773), .B(n628), .Z(n191) );
  COND1XL U5351 ( .A(n643), .B(n649), .C(n3622), .Z(n642) );
  CND2X1 U5352 ( .A(n774), .B(n634), .Z(n192) );
  COND1XL U5353 ( .A(n649), .B(n636), .C(n4195), .Z(n635) );
  CENX1 U5354 ( .A(n667), .B(n197), .Z(product[15]) );
  CANR1XL U5355 ( .A(n779), .B(n667), .C(n664), .Z(n662) );
  CANR1XL U5356 ( .A(n667), .B(n658), .C(n3311), .Z(n657) );
  CEOXL U5357 ( .A(n194), .B(n649), .Z(product[18]) );
  CND2XL U5358 ( .A(n776), .B(n3622), .Z(n194) );
  CENX1 U5359 ( .A(n4270), .B(n3043), .Z(n1107) );
  CENX1 U5360 ( .A(n1111), .B(n1134), .Z(n4270) );
  CENX1 U5361 ( .A(n4271), .B(n1439), .Z(n1437) );
  CND2XL U5362 ( .A(n739), .B(n303), .Z(n157) );
  CND2XL U5363 ( .A(n3713), .B(n316), .Z(n158) );
  CNR2X1 U5364 ( .A(n1627), .B(n1640), .Z(n665) );
  COR2X1 U5365 ( .A(n1580), .B(n1563), .Z(n4274) );
  COR2X1 U5366 ( .A(n1597), .B(n1612), .Z(n4277) );
  CND2X1 U5367 ( .A(n3119), .B(n1640), .Z(n666) );
  CND2X1 U5368 ( .A(n893), .B(n906), .Z(n392) );
  CND2X1 U5369 ( .A(n957), .B(n974), .Z(n434) );
  CND2X1 U5370 ( .A(n939), .B(n956), .Z(n425) );
  CND2X1 U5371 ( .A(n855), .B(n866), .Z(n351) );
  CND2X1 U5372 ( .A(n1563), .B(n1580), .Z(n641) );
  CND2X1 U5373 ( .A(n1597), .B(n1612), .Z(n656) );
  CND2X1 U5374 ( .A(n907), .B(n922), .Z(n403) );
  CND2X1 U5375 ( .A(n1505), .B(n1524), .Z(n623) );
  CND2X1 U5376 ( .A(n1545), .B(n1562), .Z(n634) );
  COND1XL U5377 ( .A(n324), .B(n334), .C(n327), .Z(n323) );
  CND2XL U5378 ( .A(n780), .B(n672), .Z(n198) );
  COND1XL U5379 ( .A(n674), .B(n676), .C(n675), .Z(n673) );
  CENX1 U5380 ( .A(n689), .B(n201), .Z(product[11]) );
  CENX1 U5381 ( .A(n202), .B(n695), .Z(product[10]) );
  CND2X1 U5382 ( .A(n784), .B(n694), .Z(n202) );
  COND1XL U5383 ( .A(n696), .B(n698), .C(n697), .Z(n695) );
  CANR1XL U5384 ( .A(n4280), .B(n689), .C(n686), .Z(n684) );
  CEOXL U5385 ( .A(n199), .B(n676), .Z(product[13]) );
  CEOXL U5386 ( .A(n698), .B(n203), .Z(product[9]) );
  CNR2X1 U5387 ( .A(n1653), .B(n1664), .Z(n674) );
  CNR2X1 U5388 ( .A(n1693), .B(n1700), .Z(n696) );
  CNR2X1 U5389 ( .A(n1685), .B(n1692), .Z(n693) );
  CND2XL U5390 ( .A(n735), .B(n255), .Z(n153) );
  CND2XL U5391 ( .A(n736), .B(n266), .Z(n154) );
  CAOR1X1 U5392 ( .A(n721), .B(n4285), .C(n718), .Z(n4278) );
  CNR2X1 U5393 ( .A(n1701), .B(n1706), .Z(n700) );
  COR2X1 U5394 ( .A(n845), .B(n854), .Z(n4279) );
  COR2X1 U5395 ( .A(n1675), .B(n1684), .Z(n4280) );
  CND2X1 U5396 ( .A(n1653), .B(n1664), .Z(n675) );
  CND2X1 U5397 ( .A(n1693), .B(n1700), .Z(n697) );
  CND2X1 U5398 ( .A(n845), .B(n854), .Z(n342) );
  CND2X1 U5399 ( .A(n1675), .B(n1684), .Z(n688) );
  CND2X1 U5400 ( .A(n1665), .B(n1674), .Z(n683) );
  CENX1 U5401 ( .A(n207), .B(n4278), .Z(product[5]) );
  CEOXL U5402 ( .A(n724), .B(n209), .Z(product[3]) );
  CND2X1 U5403 ( .A(n791), .B(n723), .Z(n209) );
  CEOXL U5404 ( .A(n710), .B(n206), .Z(product[6]) );
  CND2X1 U5405 ( .A(n788), .B(n709), .Z(n206) );
  COR2X1 U5406 ( .A(n807), .B(n812), .Z(n4282) );
  CND2X1 U5407 ( .A(n835), .B(n844), .Z(n327) );
  CND2X1 U5408 ( .A(n807), .B(n812), .Z(n279) );
  CND2X1 U5409 ( .A(n813), .B(n818), .Z(n296) );
  CENX1 U5410 ( .A(n210), .B(n729), .Z(product[2]) );
  CNR2X1 U5411 ( .A(n1713), .B(n1716), .Z(n708) );
  CNR2X1 U5412 ( .A(n1723), .B(n2218), .Z(n722) );
  COR2X1 U5413 ( .A(n1707), .B(n1712), .Z(n4283) );
  COR2X1 U5414 ( .A(n1717), .B(n1720), .Z(n4284) );
  CENX1 U5415 ( .A(n1798), .B(n2034), .Z(n1273) );
  CND2X1 U5416 ( .A(n1721), .B(n1722), .Z(n720) );
  CND2X1 U5417 ( .A(n1717), .B(n1720), .Z(n714) );
  CND2X1 U5418 ( .A(n2250), .B(n2219), .Z(n728) );
  CND2X1 U5419 ( .A(n1707), .B(n1712), .Z(n706) );
  COR2X1 U5420 ( .A(n1721), .B(n1722), .Z(n4285) );
  CNR2X1 U5421 ( .A(n806), .B(n803), .Z(n265) );
  CNR2X1 U5422 ( .A(n799), .B(n802), .Z(n254) );
  COR2X1 U5423 ( .A(n798), .B(n797), .Z(net18422) );
  CND2X1 U5424 ( .A(n806), .B(n803), .Z(n266) );
  CND2X1 U5425 ( .A(n798), .B(n797), .Z(n246) );
  CAN2XL U5426 ( .A(n3723), .B(n731), .Z(product[1]) );
  CENX1 U5427 ( .A(n2789), .B(net16059), .Z(n2591) );
  CENX1 U5428 ( .A(n4330), .B(n4258), .Z(n2434) );
  CENX1 U5429 ( .A(net16548), .B(net16059), .Z(n2592) );
  CENX1 U5430 ( .A(n4335), .B(net16059), .Z(n2589) );
  CENX1 U5431 ( .A(net16550), .B(net16059), .Z(n2593) );
  CENX1 U5432 ( .A(n4336), .B(net16059), .Z(n2588) );
  CENX1 U5433 ( .A(n4337), .B(net16059), .Z(n2587) );
  CENX1 U5434 ( .A(net16558), .B(n4258), .Z(n2432) );
  CENX1 U5435 ( .A(net16548), .B(n4258), .Z(n2427) );
  CENX1 U5436 ( .A(n4334), .B(n4258), .Z(n2429) );
  CENX1 U5437 ( .A(net16550), .B(n4258), .Z(n2428) );
  CENX1 U5438 ( .A(n4335), .B(n4258), .Z(n2424) );
  CENX1 U5439 ( .A(n4338), .B(net16059), .Z(n2586) );
  CENX1 U5440 ( .A(n2808), .B(n4292), .Z(n2445) );
  CENX1 U5441 ( .A(n4324), .B(net16850), .Z(n2475) );
  CENX1 U5442 ( .A(n2808), .B(net16850), .Z(n2478) );
  CENX1 U5443 ( .A(n4330), .B(n4345), .Z(n2764) );
  CENX1 U5444 ( .A(n4331), .B(n4345), .Z(n2763) );
  CENX1 U5445 ( .A(n4336), .B(n4343), .Z(n2753) );
  CENX1 U5446 ( .A(n2810), .B(n4344), .Z(n2777) );
  CENX1 U5447 ( .A(n4321), .B(n4344), .Z(n2776) );
  CENX1 U5448 ( .A(n4326), .B(n4344), .Z(n2770) );
  CENX1 U5449 ( .A(n2789), .B(n4343), .Z(n2756) );
  CENX1 U5450 ( .A(n2802), .B(n4344), .Z(n2769) );
  CENX1 U5451 ( .A(net16550), .B(n4343), .Z(n2758) );
  CENX1 U5452 ( .A(n4335), .B(n4343), .Z(n2754) );
  CENX1 U5453 ( .A(n4327), .B(n4344), .Z(n2767) );
  CENX1 U5454 ( .A(n4322), .B(n4344), .Z(n2774) );
  CENX1 U5455 ( .A(n4328), .B(n4344), .Z(n2766) );
  CENX1 U5456 ( .A(net16548), .B(n4343), .Z(n2757) );
  CENX1 U5457 ( .A(n2808), .B(n4344), .Z(n2775) );
  CENX1 U5458 ( .A(n4334), .B(n4343), .Z(n2759) );
  CENX1 U5459 ( .A(net16570), .B(n4344), .Z(n2768) );
  CENX1 U5460 ( .A(n4324), .B(n4344), .Z(n2772) );
  CENX1 U5461 ( .A(n4325), .B(n4344), .Z(n2771) );
  CENX1 U5462 ( .A(n4329), .B(n4345), .Z(n2765) );
  CENX2 U5463 ( .A(a[14]), .B(n4308), .Z(net16771) );
  CENX1 U5464 ( .A(n4341), .B(net16059), .Z(n2583) );
  CENXL U5465 ( .A(n4341), .B(net16091), .Z(n2715) );
  CNR2IXL U5466 ( .B(net16109), .A(net16816), .Z(n2219) );
  CENX1 U5467 ( .A(n4333), .B(net16037), .Z(n2496) );
  CENX1 U5468 ( .A(net16570), .B(n4292), .Z(n2438) );
  CENX1 U5469 ( .A(n4331), .B(net18643), .Z(n2532) );
  CENX1 U5470 ( .A(n2802), .B(n4292), .Z(n2439) );
  CENX1 U5471 ( .A(n4330), .B(n4291), .Z(n2368) );
  CENX1 U5472 ( .A(n4329), .B(n4291), .Z(n2369) );
  CENX1 U5473 ( .A(n4331), .B(n4291), .Z(n2367) );
  CENX1 U5474 ( .A(n4330), .B(net18643), .Z(n2533) );
  CENX1 U5475 ( .A(net16550), .B(n4253), .Z(n2395) );
  CENX1 U5476 ( .A(net16548), .B(n4253), .Z(n2394) );
  CENX1 U5477 ( .A(net16558), .B(n4291), .Z(n2366) );
  CENX1 U5478 ( .A(n4332), .B(n4291), .Z(n2365) );
  CENX1 U5479 ( .A(n4330), .B(n4253), .Z(n2401) );
  CENX1 U5480 ( .A(n4326), .B(n4292), .Z(n2440) );
  CENX1 U5481 ( .A(net16544), .B(n4253), .Z(n2392) );
  CENX1 U5482 ( .A(n4333), .B(n4291), .Z(n2364) );
  CENX1 U5483 ( .A(n4329), .B(net18936), .Z(n2534) );
  CENX1 U5484 ( .A(n4324), .B(n4292), .Z(n2442) );
  CENX1 U5485 ( .A(n2810), .B(n4292), .Z(n2447) );
  CENX1 U5486 ( .A(n4321), .B(n4292), .Z(n2446) );
  CENX1 U5487 ( .A(n4322), .B(net16788), .Z(n2609) );
  CENX1 U5488 ( .A(n2810), .B(net16037), .Z(n2513) );
  CENX1 U5489 ( .A(n4322), .B(n4292), .Z(n2444) );
  CENX1 U5490 ( .A(n2810), .B(n3730), .Z(n2612) );
  CENX1 U5491 ( .A(n4324), .B(n4362), .Z(n2277) );
  CENX1 U5492 ( .A(n2810), .B(n4362), .Z(n2282) );
  CENX1 U5493 ( .A(net16550), .B(net16844), .Z(n2692) );
  CENX1 U5494 ( .A(n4328), .B(net16069), .Z(n2634) );
  CENX1 U5495 ( .A(n4326), .B(net16069), .Z(n2638) );
  CENX1 U5496 ( .A(n4326), .B(n4362), .Z(n2275) );
  CENX1 U5497 ( .A(n2808), .B(net16069), .Z(n2643) );
  CENX1 U5498 ( .A(n4327), .B(net16069), .Z(n2635) );
  CENX1 U5499 ( .A(n4322), .B(net16069), .Z(n2642) );
  CENX1 U5500 ( .A(n4325), .B(n4362), .Z(n2276) );
  CENX1 U5501 ( .A(net16570), .B(net16069), .Z(n2636) );
  CENX1 U5502 ( .A(n4328), .B(n4362), .Z(n2271) );
  CENX1 U5503 ( .A(n2802), .B(n4362), .Z(n2274) );
  CENX1 U5504 ( .A(net16570), .B(n4362), .Z(n2273) );
  CENX1 U5505 ( .A(n4324), .B(net16069), .Z(n2640) );
  CENX1 U5506 ( .A(n2802), .B(net16069), .Z(n2637) );
  CENX1 U5507 ( .A(n4327), .B(n4362), .Z(n2272) );
  CENX1 U5508 ( .A(n4342), .B(net16069), .Z(n2615) );
  CENX1 U5509 ( .A(n4342), .B(n3729), .Z(n2582) );
  CNR2IX1 U5510 ( .B(net16109), .A(n3277), .Z(n1957) );
  CNR2IXL U5511 ( .B(net16109), .A(net16793), .Z(n2120) );
  CNR2IX1 U5512 ( .B(net16109), .A(n3839), .Z(n2087) );
  CNR2IXL U5513 ( .B(net16109), .A(net19508), .Z(n2153) );
  CNR2IXL U5514 ( .B(net16109), .A(net16771), .Z(n2021) );
  CENX1 U5515 ( .A(net16548), .B(n4251), .Z(n2295) );
  CENX1 U5516 ( .A(n4337), .B(n4258), .Z(n2422) );
  CENX1 U5517 ( .A(net16550), .B(n4251), .Z(n2296) );
  CENX1 U5518 ( .A(n4336), .B(n4258), .Z(n2423) );
  CENX1 U5519 ( .A(n4323), .B(n4344), .Z(n2773) );
  CENX1 U5520 ( .A(n4341), .B(n4258), .Z(n2418) );
  CENX1 U5521 ( .A(n4340), .B(n4262), .Z(n2254) );
  CENX1 U5522 ( .A(n2810), .B(net16069), .Z(n2645) );
  CENX1 U5523 ( .A(n4323), .B(net16069), .Z(n2641) );
  CENX1 U5524 ( .A(n4337), .B(n4262), .Z(n2257) );
  CENX1 U5525 ( .A(n4338), .B(n4262), .Z(n2256) );
  CENX1 U5526 ( .A(n4339), .B(n4262), .Z(n2255) );
  CENX1 U5527 ( .A(n4341), .B(n4262), .Z(n2253) );
  CENX1 U5528 ( .A(n4342), .B(n4362), .Z(n2252) );
  CNR2IX1 U5529 ( .B(net16109), .A(n6), .Z(product[0]) );
  CIVX2 U5530 ( .A(n57), .Z(n4350) );
  CNIVX8 U5531 ( .A(n2791), .Z(net16550) );
  CNIVX8 U5532 ( .A(n2781), .Z(n4341) );
  CNIVX4 U5533 ( .A(n2804), .Z(n4325) );
  CNIVX4 U5534 ( .A(n2807), .Z(n4322) );
  CNIVX4 U5535 ( .A(n2803), .Z(n4326) );
  COND1XL U5536 ( .A(n213), .B(net19409), .C(n214), .Z(n212) );
  CENXL U5537 ( .A(n304), .B(n157), .Z(product[55]) );
  CENXL U5538 ( .A(n154), .B(n267), .Z(product[58]) );
  CIVX8 U5539 ( .A(net16849), .Z(net16850) );
  CND2IXL U5540 ( .B(net16109), .A(n4352), .Z(n2449) );
  CND2X1 U5541 ( .A(n3825), .B(n534), .Z(n514) );
  CIVXL U5542 ( .A(n4353), .Z(n4352) );
  CENX1 U5543 ( .A(n4327), .B(net16850), .Z(n2470) );
  CIVX8 U5544 ( .A(n141), .Z(n4293) );
  CENX4 U5545 ( .A(n4102), .B(n4347), .Z(net16793) );
  CENXL U5546 ( .A(n256), .B(n153), .Z(product[59]) );
  CENXL U5547 ( .A(n280), .B(n155), .Z(product[57]) );
  CND2IXL U5548 ( .B(net16109), .A(n4349), .Z(n2581) );
  CND2X1 U5549 ( .A(n1135), .B(n1137), .Z(n4297) );
  CND2XL U5550 ( .A(n1160), .B(n1137), .Z(n4298) );
  CENX1 U5551 ( .A(net16548), .B(net18643), .Z(n2526) );
  CND2IXL U5552 ( .B(net16109), .A(n3574), .Z(n2680) );
  CENX1 U5553 ( .A(net16548), .B(n4254), .Z(n2658) );
  CENX1 U5554 ( .A(net16550), .B(n4254), .Z(n2659) );
  CND2XL U5555 ( .A(n1943), .B(n1855), .Z(n4299) );
  CND2XL U5556 ( .A(n1855), .B(n1827), .Z(n4301) );
  CND3X1 U5557 ( .A(n4299), .B(n4301), .C(n4300), .Z(n1268) );
  CNR2XL U5558 ( .A(n4033), .B(n2375), .Z(n4305) );
  COAN1XL U5559 ( .A(n4088), .B(n3500), .C(n3131), .Z(n4309) );
  CIVXL U5560 ( .A(n4309), .Z(n4310) );
  CANR1XL U5561 ( .A(n3717), .B(n4310), .C(n528), .Z(n526) );
  CND2XL U5562 ( .A(n1439), .B(n1462), .Z(n4311) );
  CND2XL U5563 ( .A(n1462), .B(n1441), .Z(n4313) );
  CND2XL U5564 ( .A(n1389), .B(n3569), .Z(n4314) );
  CND2XL U5565 ( .A(n1389), .B(n1414), .Z(n4315) );
  CND3XL U5566 ( .A(n4314), .B(n4315), .C(n4316), .Z(n1386) );
  COND2XL U5567 ( .A(net19555), .B(n4142), .C(n6), .D(n2779), .Z(n1739) );
  CENX1 U5568 ( .A(n4332), .B(n4345), .Z(n2761) );
  CENX1 U5569 ( .A(n4333), .B(n4345), .Z(n2760) );
  CND2IXL U5570 ( .B(net16109), .A(n4345), .Z(n2779) );
  CND2X1 U5571 ( .A(n2251), .B(n1739), .Z(n731) );
  COR2XL U5572 ( .A(n3533), .B(n3661), .Z(n4317) );
  CND2XL U5573 ( .A(n1134), .B(n1109), .Z(n4318) );
  CND2XL U5574 ( .A(n1134), .B(n1111), .Z(n4320) );
  COND2XL U5575 ( .A(n4135), .B(n3880), .C(net19151), .D(n2581), .Z(n1733) );
  COND2XL U5576 ( .A(n3877), .B(net19076), .C(n3839), .D(n2614), .Z(n1734) );
  COND2XL U5577 ( .A(n4001), .B(net19016), .C(net16816), .D(n2746), .Z(n1738)
         );
  COND2XL U5578 ( .A(n90), .B(n3195), .C(n3278), .D(n2482), .Z(n1730) );
  COND2XL U5579 ( .A(n4003), .B(n4190), .C(net19508), .D(n2680), .Z(n1736) );
  COND2XL U5580 ( .A(n135), .B(n4014), .C(n132), .D(n2317), .Z(n1725) );
  CIVXL U5581 ( .A(n3660), .Z(n757) );
  CIVX1 U5582 ( .A(net16089), .Z(net16087) );
  CIVX2 U5583 ( .A(n992), .Z(n993) );
  CIVX2 U5584 ( .A(n4016), .Z(n955) );
  CIVX2 U5585 ( .A(n920), .Z(n921) );
  CIVX2 U5586 ( .A(n890), .Z(n891) );
  CIVX2 U5587 ( .A(n842), .Z(n843) );
  CIVX2 U5588 ( .A(n824), .Z(n825) );
  CIVX2 U5589 ( .A(n810), .Z(n811) );
  CIVX2 U5590 ( .A(n800), .Z(n801) );
  CIVX2 U5591 ( .A(n722), .Z(n791) );
  CIVX2 U5592 ( .A(n708), .Z(n788) );
  CIVX2 U5593 ( .A(n700), .Z(n786) );
  CIVX2 U5594 ( .A(n696), .Z(n785) );
  CIVX2 U5595 ( .A(n674), .Z(n781) );
  CIVX2 U5596 ( .A(n324), .Z(n741) );
  CIVX2 U5597 ( .A(n295), .Z(n738) );
  CIVX2 U5598 ( .A(n731), .Z(n729) );
  CIVX2 U5599 ( .A(n728), .Z(n726) );
  CIVX2 U5600 ( .A(n720), .Z(n718) );
  CIVX2 U5601 ( .A(n714), .Z(n712) );
  CIVX2 U5602 ( .A(n706), .Z(n704) );
  CIVX2 U5603 ( .A(n699), .Z(n698) );
  CIVX2 U5604 ( .A(n688), .Z(n686) );
  CIVX2 U5605 ( .A(n683), .Z(n681) );
  CIVX2 U5606 ( .A(n656), .Z(n654) );
  CIVX2 U5607 ( .A(n628), .Z(n626) );
  CIVX2 U5608 ( .A(n618), .Z(n616) );
  CIVX2 U5609 ( .A(n603), .Z(n601) );
  CIVX2 U5610 ( .A(n468), .Z(n753) );
  CIVX2 U5611 ( .A(n351), .Z(n349) );
  CIVX2 U5612 ( .A(n342), .Z(n340) );
  CIVX2 U5613 ( .A(n333), .Z(n331) );
  CIVX2 U5614 ( .A(n316), .Z(n314) );
  CIVX2 U5615 ( .A(n303), .Z(n301) );
  CIVX2 U5616 ( .A(n302), .Z(n739) );
  CIVX2 U5617 ( .A(n279), .Z(n277) );
  CIVX2 U5618 ( .A(n274), .Z(n272) );
  CIVX2 U5619 ( .A(n265), .Z(n736) );
  CIVX2 U5620 ( .A(n254), .Z(n735) );
  CIVX2 U5621 ( .A(n1130), .Z(n1131) );
endmodule


module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push0, cmd0_en_stg0, cmd1_en_stg0, cmd0_en_stg1, cmd1_en_stg1,
         push0_stg0, cmd0_en_stg2_d, cmd1_en_stg2_d, push0_stg2, push0_stg1,
         cmd2_en_stg1, cmd2_en_stg2, cmd0_en_stg2, cmd1_en_stg2, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59,
         N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73,
         N74, N75, N76, N77, N78, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
         N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248,
         N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N399, N400, N401, N402, N403, N404, N405, N406, roundit,
         _pushout_d, N418, N419, N420, N421, N422, N423, N424, N425, N426,
         N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437,
         N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, n12,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312;
  wire   [1:0] cmd0;
  wire   [1:0] cmd0_stg0;
  wire   [1:0] cmd0_stg2;
  wire   [1:0] cmd0_stg1;
  wire   [63:0] out0_stg0;
  wire   [63:0] out0_stg2;
  wire   [63:0] out0_stg1;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] acc_cmd1;
  wire   [63:0] acc;
  wire   [63:0] out1_stg2;
  wire   [63:0] out1_stg0;
  wire   [63:0] out1_stg1;
  wire   [63:0] acc_cmd2;
  wire   [63:0] out2_stg2;
  wire   [6:0] h0_stg1;
  wire   [6:0] h0_stg0;

  CAOR2X1 U369 ( .A(h0_stg0[0]), .B(cmd2_en_stg1), .C(n1362), .D(n1985), .Z(
        n612) );
  CAOR2X1 U372 ( .A(h0_stg0[1]), .B(cmd2_en_stg1), .C(n1369), .D(n1985), .Z(
        n615) );
  CAOR2X1 U375 ( .A(h0_stg0[2]), .B(cmd2_en_stg1), .C(n1213), .D(n1985), .Z(
        n618) );
  CAOR2X1 U378 ( .A(h0_stg0[3]), .B(cmd2_en_stg1), .C(n1375), .D(n1985), .Z(
        n621) );
  CAOR2X1 U381 ( .A(h0_stg0[4]), .B(cmd2_en_stg1), .C(n1218), .D(n1985), .Z(
        n624) );
  CAOR2X1 U384 ( .A(h0_stg0[5]), .B(cmd2_en_stg1), .C(n1224), .D(n1985), .Z(
        n627) );
  CAOR2X1 U387 ( .A(h0_stg0[6]), .B(cmd2_en_stg1), .C(n1225), .D(n1985), .Z(
        n630) );
  CFD2QX2 \q0_reg[30]  ( .D(n688), .CP(clk), .CD(n1307), .Q(q0[30]) );
  CFD2QX2 \q0_reg[20]  ( .D(n678), .CP(clk), .CD(n1319), .Q(q0[20]) );
  CFD2QX2 \q0_reg[2]  ( .D(n791), .CP(clk), .CD(n1321), .Q(q0[2]) );
  CFD2QX2 \q0_reg[0]  ( .D(n790), .CP(clk), .CD(n1321), .Q(q0[0]) );
  sfilt_DW01_add_2 add_121 ( .A(out1_stg1), .B(acc_cmd1), .CI(1'b0), .SUM({
        N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, 
        N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, 
        N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, 
        N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, 
        N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, 
        N212, N211, N210, N209}) );
  sfilt_DW01_add_3 add_187 ( .A(out2_stg2), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, roundit}), 
        .CI(1'b0), .SUM({N481, N480, N479, N478, N477, N476, N475, N474, N473, 
        N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, 
        N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, 
        N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, 
        N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, 
        N424, N423, N422, N421, N420, N419, N418}) );
  sfilt_DW_mult_tc_1 r304 ( .a({q0[31:19], n804, q0[17], n1127, q0[15:0]}), 
        .b(h0), .product({N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15}) );
  CFD2QX1 \q0_reg[27]  ( .D(n685), .CP(clk), .CD(n1307), .Q(q0[27]) );
  CFD2QX1 \q0_reg[15]  ( .D(n673), .CP(clk), .CD(n1320), .Q(q0[15]) );
  CFD2QX1 \q0_reg[13]  ( .D(n671), .CP(clk), .CD(n1320), .Q(q0[13]) );
  CFD2QX1 \q0_reg[19]  ( .D(n677), .CP(clk), .CD(n1319), .Q(q0[19]) );
  CFD2QXL \out0_stg0_reg[42]  ( .D(N57), .CP(clk), .CD(n1347), .Q(
        out0_stg0[42]) );
  CFD2QXL \out1_stg0_reg[42]  ( .D(N57), .CP(clk), .CD(n1308), .Q(
        out1_stg0[42]) );
  CFD2QXL \out0_stg0_reg[43]  ( .D(N58), .CP(clk), .CD(n1346), .Q(
        out0_stg0[43]) );
  CFD2QXL \out1_stg0_reg[43]  ( .D(N58), .CP(clk), .CD(n1308), .Q(
        out1_stg0[43]) );
  CFD2QXL \out0_stg0_reg[44]  ( .D(N59), .CP(clk), .CD(n1346), .Q(
        out0_stg0[44]) );
  CFD2QXL \out1_stg0_reg[44]  ( .D(N59), .CP(clk), .CD(n1307), .Q(
        out1_stg0[44]) );
  CFD2QXL \out0_stg0_reg[45]  ( .D(N60), .CP(clk), .CD(n1346), .Q(
        out0_stg0[45]) );
  CFD2QXL \out1_stg0_reg[45]  ( .D(N60), .CP(clk), .CD(n1307), .Q(
        out1_stg0[45]) );
  CFD2QXL \out0_stg0_reg[46]  ( .D(N61), .CP(clk), .CD(n1345), .Q(
        out0_stg0[46]) );
  CFD2QXL \out1_stg0_reg[46]  ( .D(N61), .CP(clk), .CD(n1307), .Q(
        out1_stg0[46]) );
  CFD2QXL \out0_stg0_reg[47]  ( .D(N62), .CP(clk), .CD(n1345), .Q(
        out0_stg0[47]) );
  CFD2QXL \out1_stg0_reg[47]  ( .D(N62), .CP(clk), .CD(n1313), .Q(
        out1_stg0[47]) );
  CFD2QXL \out0_stg0_reg[48]  ( .D(N63), .CP(clk), .CD(n1344), .Q(
        out0_stg0[48]) );
  CFD2QXL \out1_stg0_reg[48]  ( .D(N63), .CP(clk), .CD(n1331), .Q(
        out1_stg0[48]) );
  CFD2QXL \out0_stg0_reg[49]  ( .D(N64), .CP(clk), .CD(n1344), .Q(
        out0_stg0[49]) );
  CFD2QXL \out1_stg0_reg[49]  ( .D(N64), .CP(clk), .CD(n1331), .Q(
        out1_stg0[49]) );
  CFD2QXL \out0_stg0_reg[50]  ( .D(N65), .CP(clk), .CD(n1344), .Q(
        out0_stg0[50]) );
  CFD2QXL \out1_stg0_reg[50]  ( .D(N65), .CP(clk), .CD(n1331), .Q(
        out1_stg0[50]) );
  CFD2QXL \out0_stg0_reg[51]  ( .D(N66), .CP(clk), .CD(n1319), .Q(
        out0_stg0[51]) );
  CFD2QXL \out1_stg0_reg[51]  ( .D(N66), .CP(clk), .CD(n1331), .Q(
        out1_stg0[51]) );
  CFD2QXL \out0_stg0_reg[52]  ( .D(N67), .CP(clk), .CD(n1318), .Q(
        out0_stg0[52]) );
  CFD2QXL \out1_stg0_reg[52]  ( .D(N67), .CP(clk), .CD(n1330), .Q(
        out1_stg0[52]) );
  CFD2QXL \out0_stg0_reg[53]  ( .D(N68), .CP(clk), .CD(n1318), .Q(
        out0_stg0[53]) );
  CFD2QXL \out1_stg0_reg[53]  ( .D(N68), .CP(clk), .CD(n1330), .Q(
        out1_stg0[53]) );
  CFD2QXL \out0_stg0_reg[54]  ( .D(N69), .CP(clk), .CD(n1318), .Q(
        out0_stg0[54]) );
  CFD2QXL \out1_stg0_reg[54]  ( .D(N69), .CP(clk), .CD(n1330), .Q(
        out1_stg0[54]) );
  CFD2QXL \out0_stg0_reg[55]  ( .D(N70), .CP(clk), .CD(n1317), .Q(
        out0_stg0[55]) );
  CFD2QXL \out1_stg0_reg[55]  ( .D(N70), .CP(clk), .CD(n1330), .Q(
        out1_stg0[55]) );
  CFD2QXL \out0_stg0_reg[56]  ( .D(N71), .CP(clk), .CD(n1317), .Q(
        out0_stg0[56]) );
  CFD2QXL \out1_stg0_reg[56]  ( .D(N71), .CP(clk), .CD(n1330), .Q(
        out1_stg0[56]) );
  CFD2QXL \out0_stg0_reg[57]  ( .D(N72), .CP(clk), .CD(n1317), .Q(
        out0_stg0[57]) );
  CFD2QXL \out1_stg0_reg[57]  ( .D(N72), .CP(clk), .CD(n1330), .Q(
        out1_stg0[57]) );
  CFD2QXL \out0_stg0_reg[58]  ( .D(N73), .CP(clk), .CD(n1316), .Q(
        out0_stg0[58]) );
  CFD2QXL \out1_stg0_reg[58]  ( .D(N73), .CP(clk), .CD(n1329), .Q(
        out1_stg0[58]) );
  CFD2QXL \out0_stg0_reg[59]  ( .D(N74), .CP(clk), .CD(n1316), .Q(
        out0_stg0[59]) );
  CFD2QXL \out1_stg0_reg[59]  ( .D(N74), .CP(clk), .CD(n1329), .Q(
        out1_stg0[59]) );
  CFD2QXL \out0_stg0_reg[60]  ( .D(N75), .CP(clk), .CD(n1315), .Q(
        out0_stg0[60]) );
  CFD2QXL \out1_stg0_reg[60]  ( .D(N75), .CP(clk), .CD(n1329), .Q(
        out1_stg0[60]) );
  CFD2QXL \out0_stg0_reg[61]  ( .D(N76), .CP(clk), .CD(n1315), .Q(
        out0_stg0[61]) );
  CFD2QXL \out1_stg0_reg[61]  ( .D(N76), .CP(clk), .CD(n1329), .Q(
        out1_stg0[61]) );
  CFD2QXL \out0_stg0_reg[62]  ( .D(N77), .CP(clk), .CD(n1315), .Q(
        out0_stg0[62]) );
  CFD2QXL \out1_stg0_reg[62]  ( .D(N77), .CP(clk), .CD(n1329), .Q(
        out1_stg0[62]) );
  CFD2QXL \out0_stg1_reg[63]  ( .D(n1096), .CP(clk), .CD(n1323), .Q(
        out0_stg1[63]) );
  CFD2QXL \out0_stg1_reg[62]  ( .D(n1094), .CP(clk), .CD(n1315), .Q(
        out0_stg1[62]) );
  CFD2QXL \out0_stg1_reg[61]  ( .D(n1092), .CP(clk), .CD(n1315), .Q(
        out0_stg1[61]) );
  CFD2QXL \out0_stg1_reg[60]  ( .D(n1090), .CP(clk), .CD(n1315), .Q(
        out0_stg1[60]) );
  CFD2QXL \out0_stg1_reg[59]  ( .D(n1088), .CP(clk), .CD(n1316), .Q(
        out0_stg1[59]) );
  CFD2QXL \out0_stg1_reg[58]  ( .D(n1086), .CP(clk), .CD(n1316), .Q(
        out0_stg1[58]) );
  CFD2QXL \out0_stg1_reg[57]  ( .D(n1084), .CP(clk), .CD(n1317), .Q(
        out0_stg1[57]) );
  CFD2QXL \out0_stg1_reg[56]  ( .D(n1082), .CP(clk), .CD(n1317), .Q(
        out0_stg1[56]) );
  CFD2QXL \out0_stg1_reg[55]  ( .D(n1080), .CP(clk), .CD(n1317), .Q(
        out0_stg1[55]) );
  CFD2QXL \out0_stg1_reg[54]  ( .D(n1078), .CP(clk), .CD(n1318), .Q(
        out0_stg1[54]) );
  CFD2QXL \out0_stg1_reg[53]  ( .D(n1076), .CP(clk), .CD(n1318), .Q(
        out0_stg1[53]) );
  CFD2QXL \out0_stg1_reg[52]  ( .D(n1074), .CP(clk), .CD(n1319), .Q(
        out0_stg1[52]) );
  CFD2QXL \out0_stg1_reg[51]  ( .D(n1072), .CP(clk), .CD(n1319), .Q(
        out0_stg1[51]) );
  CFD2QXL \out0_stg1_reg[50]  ( .D(n1070), .CP(clk), .CD(n1344), .Q(
        out0_stg1[50]) );
  CFD2QXL \out0_stg1_reg[49]  ( .D(n1068), .CP(clk), .CD(n1344), .Q(
        out0_stg1[49]) );
  CFD2QXL \out0_stg1_reg[48]  ( .D(n1066), .CP(clk), .CD(n1344), .Q(
        out0_stg1[48]) );
  CFD2QXL \out0_stg1_reg[47]  ( .D(n1064), .CP(clk), .CD(n1345), .Q(
        out0_stg1[47]) );
  CFD2QXL \out0_stg1_reg[46]  ( .D(n1062), .CP(clk), .CD(n1345), .Q(
        out0_stg1[46]) );
  CFD2QXL \out0_stg1_reg[45]  ( .D(n1060), .CP(clk), .CD(n1346), .Q(
        out0_stg1[45]) );
  CFD2QXL \out0_stg1_reg[44]  ( .D(n1058), .CP(clk), .CD(n1346), .Q(
        out0_stg1[44]) );
  CFD2QXL \out0_stg1_reg[43]  ( .D(n1056), .CP(clk), .CD(n1346), .Q(
        out0_stg1[43]) );
  CFD2QXL \out0_stg1_reg[42]  ( .D(n1054), .CP(clk), .CD(n1347), .Q(
        out0_stg1[42]) );
  CFD2QXL \out0_stg1_reg[41]  ( .D(n1052), .CP(clk), .CD(n1347), .Q(
        out0_stg1[41]) );
  CFD2QXL \out0_stg1_reg[40]  ( .D(n1050), .CP(clk), .CD(n1348), .Q(
        out0_stg1[40]) );
  CFD2QXL \out0_stg1_reg[39]  ( .D(n1048), .CP(clk), .CD(n1348), .Q(
        out0_stg1[39]) );
  CFD2QXL \out0_stg1_reg[38]  ( .D(n1046), .CP(clk), .CD(n1348), .Q(
        out0_stg1[38]) );
  CFD2QXL \out0_stg1_reg[37]  ( .D(n1044), .CP(clk), .CD(n1349), .Q(
        out0_stg1[37]) );
  CFD2QXL \out0_stg1_reg[36]  ( .D(n1042), .CP(clk), .CD(n1349), .Q(
        out0_stg1[36]) );
  CFD2QXL \out0_stg1_reg[35]  ( .D(n1040), .CP(clk), .CD(n1349), .Q(
        out0_stg1[35]) );
  CFD2QXL \out0_stg1_reg[34]  ( .D(n1038), .CP(clk), .CD(n1350), .Q(
        out0_stg1[34]) );
  CFD2QXL \out0_stg1_reg[33]  ( .D(n1036), .CP(clk), .CD(n1350), .Q(
        out0_stg1[33]) );
  CFD2QXL \out0_stg1_reg[32]  ( .D(n1034), .CP(clk), .CD(n1351), .Q(
        out0_stg1[32]) );
  CFD2QXL \out0_stg1_reg[31]  ( .D(n1032), .CP(clk), .CD(n1351), .Q(
        out0_stg1[31]) );
  CFD2QXL \out0_stg1_reg[30]  ( .D(n1030), .CP(clk), .CD(n1351), .Q(
        out0_stg1[30]) );
  CFD2QXL \out0_stg1_reg[29]  ( .D(n1028), .CP(clk), .CD(n1352), .Q(
        out0_stg1[29]) );
  CFD2QXL \out0_stg1_reg[28]  ( .D(n1026), .CP(clk), .CD(n1352), .Q(
        out0_stg1[28]) );
  CFD2QXL \out0_stg1_reg[27]  ( .D(n1024), .CP(clk), .CD(n1353), .Q(
        out0_stg1[27]) );
  CFD2QXL \out0_stg1_reg[26]  ( .D(n1022), .CP(clk), .CD(n1353), .Q(
        out0_stg1[26]) );
  CFD2QXL \out0_stg1_reg[25]  ( .D(n1020), .CP(clk), .CD(n1353), .Q(
        out0_stg1[25]) );
  CFD2QXL \out0_stg1_reg[24]  ( .D(n1018), .CP(clk), .CD(n1354), .Q(
        out0_stg1[24]) );
  CFD2QXL \out0_stg1_reg[23]  ( .D(n1016), .CP(clk), .CD(n1354), .Q(
        out0_stg1[23]) );
  CFD2QXL \out0_stg1_reg[22]  ( .D(n1014), .CP(clk), .CD(n1355), .Q(
        out0_stg1[22]) );
  CFD2QXL \out0_stg1_reg[21]  ( .D(n1012), .CP(clk), .CD(n1355), .Q(
        out0_stg1[21]) );
  CFD2QXL \out0_stg1_reg[20]  ( .D(n1010), .CP(clk), .CD(n1355), .Q(
        out0_stg1[20]) );
  CFD2QXL \out0_stg1_reg[19]  ( .D(n1008), .CP(clk), .CD(n1356), .Q(
        out0_stg1[19]) );
  CFD2QXL \out0_stg1_reg[18]  ( .D(n1006), .CP(clk), .CD(n1331), .Q(
        out0_stg1[18]) );
  CFD2QXL \out0_stg1_reg[17]  ( .D(n1004), .CP(clk), .CD(n1332), .Q(
        out0_stg1[17]) );
  CFD2QXL \out0_stg1_reg[16]  ( .D(n1002), .CP(clk), .CD(n1332), .Q(
        out0_stg1[16]) );
  CFD2QXL \out0_stg1_reg[15]  ( .D(n1000), .CP(clk), .CD(n1333), .Q(
        out0_stg1[15]) );
  CFD2QXL \out0_stg1_reg[14]  ( .D(n998), .CP(clk), .CD(n1333), .Q(
        out0_stg1[14]) );
  CFD2QXL \out0_stg1_reg[13]  ( .D(n996), .CP(clk), .CD(n1333), .Q(
        out0_stg1[13]) );
  CFD2QXL \out0_stg1_reg[12]  ( .D(n994), .CP(clk), .CD(n1334), .Q(
        out0_stg1[12]) );
  CFD2QXL \out0_stg1_reg[11]  ( .D(n992), .CP(clk), .CD(n1334), .Q(
        out0_stg1[11]) );
  CFD2QXL \out0_stg1_reg[10]  ( .D(n990), .CP(clk), .CD(n1335), .Q(
        out0_stg1[10]) );
  CFD2QXL \out0_stg1_reg[9]  ( .D(n988), .CP(clk), .CD(n1335), .Q(out0_stg1[9]) );
  CFD2QXL \out0_stg1_reg[8]  ( .D(n986), .CP(clk), .CD(n1335), .Q(out0_stg1[8]) );
  CFD2QXL \out0_stg1_reg[7]  ( .D(n984), .CP(clk), .CD(n1336), .Q(out0_stg1[7]) );
  CFD2QXL \out0_stg1_reg[6]  ( .D(n982), .CP(clk), .CD(n1336), .Q(out0_stg1[6]) );
  CFD2QXL \out0_stg1_reg[5]  ( .D(n980), .CP(clk), .CD(n1336), .Q(out0_stg1[5]) );
  CFD2QXL \out0_stg1_reg[4]  ( .D(n978), .CP(clk), .CD(n1337), .Q(out0_stg1[4]) );
  CFD2QXL \out0_stg1_reg[3]  ( .D(n976), .CP(clk), .CD(n1337), .Q(out0_stg1[3]) );
  CFD2QXL \out0_stg1_reg[2]  ( .D(n974), .CP(clk), .CD(n1338), .Q(out0_stg1[2]) );
  CFD2QXL \out0_stg1_reg[1]  ( .D(n972), .CP(clk), .CD(n1338), .Q(out0_stg1[1]) );
  CFD2QXL \out0_stg1_reg[0]  ( .D(n970), .CP(clk), .CD(n1338), .Q(out0_stg1[0]) );
  CFD2QXL cmd1_en_stg1_reg ( .D(cmd1_en_stg0), .CP(clk), .CD(n1314), .Q(
        cmd1_en_stg1) );
  CFD2QXL cmd0_en_stg1_reg ( .D(cmd0_en_stg0), .CP(clk), .CD(n1339), .Q(
        cmd0_en_stg1) );
  CFD2QXL \dout_reg[31]  ( .D(n789), .CP(clk), .CD(n1343), .Q(z[31]) );
  CFD2QXL \dout_reg[30]  ( .D(n788), .CP(clk), .CD(n1343), .Q(z[30]) );
  CFD2QXL \dout_reg[29]  ( .D(n787), .CP(clk), .CD(n1343), .Q(z[29]) );
  CFD2QXL \dout_reg[28]  ( .D(n786), .CP(clk), .CD(n1343), .Q(z[28]) );
  CFD2QXL \dout_reg[27]  ( .D(n785), .CP(clk), .CD(n1343), .Q(z[27]) );
  CFD2QXL \dout_reg[26]  ( .D(n784), .CP(clk), .CD(n1343), .Q(z[26]) );
  CFD2QXL \dout_reg[25]  ( .D(n783), .CP(clk), .CD(n1343), .Q(z[25]) );
  CFD2QXL \dout_reg[24]  ( .D(n782), .CP(clk), .CD(n1343), .Q(z[24]) );
  CFD2QXL \dout_reg[23]  ( .D(n781), .CP(clk), .CD(n1343), .Q(z[23]) );
  CFD2QXL \dout_reg[22]  ( .D(n780), .CP(clk), .CD(n1343), .Q(z[22]) );
  CFD2QXL \dout_reg[21]  ( .D(n779), .CP(clk), .CD(n1343), .Q(z[21]) );
  CFD2QXL \dout_reg[20]  ( .D(n778), .CP(clk), .CD(n1343), .Q(z[20]) );
  CFD2QXL \dout_reg[19]  ( .D(n777), .CP(clk), .CD(n1342), .Q(z[19]) );
  CFD2QXL \dout_reg[18]  ( .D(n776), .CP(clk), .CD(n1342), .Q(z[18]) );
  CFD2QXL \dout_reg[17]  ( .D(n775), .CP(clk), .CD(n1342), .Q(z[17]) );
  CFD2QXL \dout_reg[16]  ( .D(n774), .CP(clk), .CD(n1342), .Q(z[16]) );
  CFD2QXL \dout_reg[15]  ( .D(n773), .CP(clk), .CD(n1342), .Q(z[15]) );
  CFD2QXL \dout_reg[14]  ( .D(n772), .CP(clk), .CD(n1342), .Q(z[14]) );
  CFD2QXL \dout_reg[13]  ( .D(n771), .CP(clk), .CD(n1342), .Q(z[13]) );
  CFD2QXL \dout_reg[12]  ( .D(n770), .CP(clk), .CD(n1342), .Q(z[12]) );
  CFD2QXL \dout_reg[11]  ( .D(n769), .CP(clk), .CD(n1342), .Q(z[11]) );
  CFD2QXL \dout_reg[10]  ( .D(n768), .CP(clk), .CD(n1342), .Q(z[10]) );
  CFD2QXL \dout_reg[9]  ( .D(n767), .CP(clk), .CD(n1342), .Q(z[9]) );
  CFD2QXL \dout_reg[8]  ( .D(n766), .CP(clk), .CD(n1342), .Q(z[8]) );
  CFD2QXL \dout_reg[7]  ( .D(n765), .CP(clk), .CD(n1342), .Q(z[7]) );
  CFD2QXL \dout_reg[6]  ( .D(n764), .CP(clk), .CD(n1341), .Q(z[6]) );
  CFD2QXL \dout_reg[5]  ( .D(n763), .CP(clk), .CD(n1341), .Q(z[5]) );
  CFD2QXL \dout_reg[4]  ( .D(n762), .CP(clk), .CD(n1341), .Q(z[4]) );
  CFD2QXL \dout_reg[3]  ( .D(n761), .CP(clk), .CD(n1341), .Q(z[3]) );
  CFD2QXL \dout_reg[2]  ( .D(n760), .CP(clk), .CD(n1341), .Q(z[2]) );
  CFD2QXL \dout_reg[1]  ( .D(n759), .CP(clk), .CD(n1341), .Q(z[1]) );
  CFD2QXL \dout_reg[0]  ( .D(n758), .CP(clk), .CD(n1341), .Q(z[0]) );
  CFD2QXL \out2_stg2_reg[58]  ( .D(n552), .CP(clk), .CD(n1324), .Q(
        out2_stg2[58]) );
  CFD2QXL \out2_stg2_reg[59]  ( .D(n551), .CP(clk), .CD(n1324), .Q(
        out2_stg2[59]) );
  CFD2QXL \out2_stg2_reg[60]  ( .D(n550), .CP(clk), .CD(n1324), .Q(
        out2_stg2[60]) );
  CFD2QXL \out2_stg2_reg[61]  ( .D(n549), .CP(clk), .CD(n1324), .Q(
        out2_stg2[61]) );
  CFD2QXL \out2_stg2_reg[62]  ( .D(n548), .CP(clk), .CD(n1324), .Q(
        out2_stg2[62]) );
  CFD2QXL \h0_stg0_reg[6]  ( .D(n968), .CP(clk), .CD(n1340), .Q(h0_stg0[6]) );
  CFD2QXL \h0_stg0_reg[5]  ( .D(n967), .CP(clk), .CD(n1341), .Q(h0_stg0[5]) );
  CFD2QXL \h0_stg0_reg[4]  ( .D(n966), .CP(clk), .CD(n1341), .Q(h0_stg0[4]) );
  CFD2QXL \h0_stg0_reg[3]  ( .D(n964), .CP(clk), .CD(n1341), .Q(h0_stg0[3]) );
  CFD2QXL \h0_stg0_reg[2]  ( .D(n963), .CP(clk), .CD(n1341), .Q(h0_stg0[2]) );
  CFD2QXL \h0_stg0_reg[1]  ( .D(n962), .CP(clk), .CD(n1341), .Q(h0_stg0[1]) );
  CFD2QXL \h0_stg0_reg[0]  ( .D(n961), .CP(clk), .CD(n1341), .Q(h0_stg0[0]) );
  CFD2QXL \h0_stg1_reg[6]  ( .D(n630), .CP(clk), .CD(n1339), .Q(h0_stg1[6]) );
  CFD2QXL \h0_stg1_reg[5]  ( .D(n627), .CP(clk), .CD(n1339), .Q(h0_stg1[5]) );
  CFD2QXL \out1_stg1_reg[63]  ( .D(n959), .CP(clk), .CD(n1329), .Q(
        out1_stg1[63]) );
  CFD2QXL \out1_stg1_reg[62]  ( .D(n957), .CP(clk), .CD(n1329), .Q(
        out1_stg1[62]) );
  CFD2QXL \out1_stg1_reg[61]  ( .D(n955), .CP(clk), .CD(n1329), .Q(
        out1_stg1[61]) );
  CFD2QXL \out1_stg1_reg[60]  ( .D(n953), .CP(clk), .CD(n1329), .Q(
        out1_stg1[60]) );
  CFD2QXL \out1_stg1_reg[54]  ( .D(n951), .CP(clk), .CD(n1330), .Q(
        out1_stg1[54]) );
  CFD2QXL \out0_stg2_reg[63]  ( .D(n691), .CP(clk), .CD(n1324), .Q(
        out0_stg2[63]) );
  CFD2QXL \cmd0_stg2_reg[0]  ( .D(n949), .CP(clk), .CD(n1340), .Q(cmd0_stg2[0]) );
  CFD2QXL \cmd0_stg2_reg[1]  ( .D(n947), .CP(clk), .CD(n1340), .Q(cmd0_stg2[1]) );
  CFD2QXL push0_reg ( .D(n1385), .CP(clk), .CD(n1340), .Q(push0) );
  CFD2QXL \out2_stg2_reg[63]  ( .D(n547), .CP(clk), .CD(n1324), .Q(
        out2_stg2[63]) );
  CFD2QXL \h0_stg1_reg[3]  ( .D(n621), .CP(clk), .CD(n1339), .Q(h0_stg1[3]) );
  CFD2QXL cmd2_en_stg1_reg ( .D(n799), .CP(clk), .CD(n1339), .Q(cmd2_en_stg1)
         );
  CFD2QXL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n1340), .Q(cmd0[0]) );
  CFD2QXL \h0_stg1_reg[2]  ( .D(n618), .CP(clk), .CD(n1339), .Q(h0_stg1[2]) );
  CFD2QXL \h0_stg1_reg[4]  ( .D(n624), .CP(clk), .CD(n1339), .Q(h0_stg1[4]) );
  CFD2QXL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n1340), .Q(cmd0[1]) );
  CFD2QXL \h0_stg1_reg[1]  ( .D(n615), .CP(clk), .CD(n1339), .Q(h0_stg1[1]) );
  CFD2QXL \out2_stg2_reg[57]  ( .D(n553), .CP(clk), .CD(n1324), .Q(
        out2_stg2[57]) );
  CFD2QXL \acc_reg[63]  ( .D(n546), .CP(clk), .CD(n1339), .Q(acc[63]) );
  CFD2QXL \acc_reg[32]  ( .D(n480), .CP(clk), .CD(n1351), .Q(acc[32]) );
  CFD2QXL \acc_reg[33]  ( .D(n478), .CP(clk), .CD(n1351), .Q(acc[33]) );
  CFD2QXL \acc_reg[34]  ( .D(n476), .CP(clk), .CD(n1350), .Q(acc[34]) );
  CFD2QXL \acc_reg[35]  ( .D(n474), .CP(clk), .CD(n1350), .Q(acc[35]) );
  CFD2QXL \acc_reg[36]  ( .D(n472), .CP(clk), .CD(n1349), .Q(acc[36]) );
  CFD2QXL \acc_reg[37]  ( .D(n470), .CP(clk), .CD(n1349), .Q(acc[37]) );
  CFD2QXL \acc_reg[38]  ( .D(n468), .CP(clk), .CD(n1349), .Q(acc[38]) );
  CFD2QXL \acc_reg[39]  ( .D(n466), .CP(clk), .CD(n1348), .Q(acc[39]) );
  CFD2QXL \acc_reg[40]  ( .D(n464), .CP(clk), .CD(n1348), .Q(acc[40]) );
  CFD2QXL \acc_reg[41]  ( .D(n462), .CP(clk), .CD(n1347), .Q(acc[41]) );
  CFD2QXL \acc_reg[42]  ( .D(n460), .CP(clk), .CD(n1347), .Q(acc[42]) );
  CFD2QXL \acc_reg[43]  ( .D(n458), .CP(clk), .CD(n1347), .Q(acc[43]) );
  CFD2QXL \acc_reg[44]  ( .D(n456), .CP(clk), .CD(n1346), .Q(acc[44]) );
  CFD2QXL \acc_reg[45]  ( .D(n454), .CP(clk), .CD(n1346), .Q(acc[45]) );
  CFD2QXL \acc_reg[46]  ( .D(n452), .CP(clk), .CD(n1345), .Q(acc[46]) );
  CFD2QXL \acc_reg[47]  ( .D(n450), .CP(clk), .CD(n1345), .Q(acc[47]) );
  CFD2QXL \acc_reg[48]  ( .D(n448), .CP(clk), .CD(n1345), .Q(acc[48]) );
  CFD2QXL \acc_reg[49]  ( .D(n446), .CP(clk), .CD(n1344), .Q(acc[49]) );
  CFD2QXL \acc_reg[50]  ( .D(n444), .CP(clk), .CD(n1344), .Q(acc[50]) );
  CFD2QXL \acc_reg[51]  ( .D(n442), .CP(clk), .CD(n1344), .Q(acc[51]) );
  CFD2QXL \acc_reg[52]  ( .D(n440), .CP(clk), .CD(n1319), .Q(acc[52]) );
  CFD2QXL \acc_reg[53]  ( .D(n438), .CP(clk), .CD(n1318), .Q(acc[53]) );
  CFD2QXL \acc_reg[54]  ( .D(n436), .CP(clk), .CD(n1318), .Q(acc[54]) );
  CFD2QXL \acc_reg[55]  ( .D(n434), .CP(clk), .CD(n1318), .Q(acc[55]) );
  CFD2QXL \acc_reg[56]  ( .D(n432), .CP(clk), .CD(n1317), .Q(acc[56]) );
  CFD2QXL \acc_reg[57]  ( .D(n430), .CP(clk), .CD(n1317), .Q(acc[57]) );
  CFD2QXL \acc_reg[58]  ( .D(n428), .CP(clk), .CD(n1316), .Q(acc[58]) );
  CFD2QXL \acc_reg[59]  ( .D(n426), .CP(clk), .CD(n1316), .Q(acc[59]) );
  CFD2QXL \acc_reg[60]  ( .D(n424), .CP(clk), .CD(n1316), .Q(acc[60]) );
  CFD2QXL \acc_reg[61]  ( .D(n422), .CP(clk), .CD(n1315), .Q(acc[61]) );
  CFD2QXL \acc_reg[62]  ( .D(n420), .CP(clk), .CD(n1315), .Q(acc[62]) );
  CFD2QXL \h0_stg1_reg[0]  ( .D(n612), .CP(clk), .CD(n1339), .Q(h0_stg1[0]) );
  CFD2QXL \out1_stg1_reg[59]  ( .D(n945), .CP(clk), .CD(n1329), .Q(
        out1_stg1[59]) );
  CFD2QXL \out1_stg1_reg[58]  ( .D(n943), .CP(clk), .CD(n1330), .Q(
        out1_stg1[58]) );
  CFD2QXL \out1_stg1_reg[57]  ( .D(n941), .CP(clk), .CD(n1330), .Q(
        out1_stg1[57]) );
  CFD2QXL \out1_stg1_reg[56]  ( .D(n939), .CP(clk), .CD(n1330), .Q(
        out1_stg1[56]) );
  CFD2QXL \out1_stg1_reg[55]  ( .D(n937), .CP(clk), .CD(n1330), .Q(
        out1_stg1[55]) );
  CFD2QXL \out1_stg1_reg[53]  ( .D(n935), .CP(clk), .CD(n1330), .Q(
        out1_stg1[53]) );
  CFD2QXL \out1_stg1_reg[52]  ( .D(n933), .CP(clk), .CD(n1330), .Q(
        out1_stg1[52]) );
  CFD2QXL \out1_stg1_reg[51]  ( .D(n931), .CP(clk), .CD(n1331), .Q(
        out1_stg1[51]) );
  CFD2QXL \out1_stg1_reg[50]  ( .D(n929), .CP(clk), .CD(n1331), .Q(
        out1_stg1[50]) );
  CFD2QXL \out1_stg1_reg[49]  ( .D(n927), .CP(clk), .CD(n1331), .Q(
        out1_stg1[49]) );
  CFD2QXL \out1_stg1_reg[48]  ( .D(n925), .CP(clk), .CD(n1331), .Q(
        out1_stg1[48]) );
  CFD2QXL \out1_stg1_reg[47]  ( .D(n923), .CP(clk), .CD(n1307), .Q(
        out1_stg1[47]) );
  CFD2QXL \out1_stg1_reg[46]  ( .D(n921), .CP(clk), .CD(n1307), .Q(
        out1_stg1[46]) );
  CFD2QXL \out1_stg1_reg[45]  ( .D(n919), .CP(clk), .CD(n1307), .Q(
        out1_stg1[45]) );
  CFD2QXL \out1_stg1_reg[44]  ( .D(n917), .CP(clk), .CD(n1307), .Q(
        out1_stg1[44]) );
  CFD2QXL \out1_stg1_reg[43]  ( .D(n915), .CP(clk), .CD(n1308), .Q(
        out1_stg1[43]) );
  CFD2QXL \out1_stg1_reg[42]  ( .D(n913), .CP(clk), .CD(n1308), .Q(
        out1_stg1[42]) );
  CFD2QXL \out1_stg1_reg[41]  ( .D(n911), .CP(clk), .CD(n1308), .Q(
        out1_stg1[41]) );
  CFD2QXL \out1_stg1_reg[40]  ( .D(n909), .CP(clk), .CD(n1308), .Q(
        out1_stg1[40]) );
  CFD2QXL \out1_stg1_reg[39]  ( .D(n907), .CP(clk), .CD(n1308), .Q(
        out1_stg1[39]) );
  CFD2QXL \out1_stg1_reg[38]  ( .D(n905), .CP(clk), .CD(n1308), .Q(
        out1_stg1[38]) );
  CFD2QXL \out1_stg1_reg[37]  ( .D(n903), .CP(clk), .CD(n1309), .Q(
        out1_stg1[37]) );
  CFD2QXL \out1_stg1_reg[36]  ( .D(n901), .CP(clk), .CD(n1309), .Q(
        out1_stg1[36]) );
  CFD2QXL \out1_stg1_reg[35]  ( .D(n899), .CP(clk), .CD(n1309), .Q(
        out1_stg1[35]) );
  CFD2QXL \out1_stg1_reg[34]  ( .D(n897), .CP(clk), .CD(n1309), .Q(
        out1_stg1[34]) );
  CFD2QXL \out1_stg1_reg[33]  ( .D(n895), .CP(clk), .CD(n1309), .Q(
        out1_stg1[33]) );
  CFD2QXL \out1_stg1_reg[32]  ( .D(n893), .CP(clk), .CD(n1309), .Q(
        out1_stg1[32]) );
  CFD2QXL \out1_stg1_reg[31]  ( .D(n891), .CP(clk), .CD(n1309), .Q(
        out1_stg1[31]) );
  CFD2QXL \out1_stg1_reg[30]  ( .D(n889), .CP(clk), .CD(n1310), .Q(
        out1_stg1[30]) );
  CFD2QXL \out1_stg1_reg[29]  ( .D(n887), .CP(clk), .CD(n1310), .Q(
        out1_stg1[29]) );
  CFD2QXL \out1_stg1_reg[28]  ( .D(n885), .CP(clk), .CD(n1310), .Q(
        out1_stg1[28]) );
  CFD2QXL \out1_stg1_reg[27]  ( .D(n883), .CP(clk), .CD(n1310), .Q(
        out1_stg1[27]) );
  CFD2QXL \out1_stg1_reg[26]  ( .D(n881), .CP(clk), .CD(n1310), .Q(
        out1_stg1[26]) );
  CFD2QXL \out1_stg1_reg[25]  ( .D(n879), .CP(clk), .CD(n1310), .Q(
        out1_stg1[25]) );
  CFD2QXL \out1_stg1_reg[24]  ( .D(n877), .CP(clk), .CD(n1311), .Q(
        out1_stg1[24]) );
  CFD2QXL \out1_stg1_reg[23]  ( .D(n875), .CP(clk), .CD(n1311), .Q(
        out1_stg1[23]) );
  CFD2QXL \out1_stg1_reg[22]  ( .D(n873), .CP(clk), .CD(n1311), .Q(
        out1_stg1[22]) );
  CFD2QXL \out1_stg1_reg[21]  ( .D(n871), .CP(clk), .CD(n1311), .Q(
        out1_stg1[21]) );
  CFD2QXL \out1_stg1_reg[20]  ( .D(n869), .CP(clk), .CD(n1311), .Q(
        out1_stg1[20]) );
  CFD2QXL \out1_stg1_reg[19]  ( .D(n867), .CP(clk), .CD(n1311), .Q(
        out1_stg1[19]) );
  CFD2QXL \out1_stg1_reg[18]  ( .D(n865), .CP(clk), .CD(n1311), .Q(
        out1_stg1[18]) );
  CFD2QXL \out1_stg1_reg[17]  ( .D(n863), .CP(clk), .CD(n1312), .Q(
        out1_stg1[17]) );
  CFD2QXL \out1_stg1_reg[16]  ( .D(n861), .CP(clk), .CD(n1312), .Q(
        out1_stg1[16]) );
  CFD2QXL \out1_stg1_reg[15]  ( .D(n859), .CP(clk), .CD(n1312), .Q(
        out1_stg1[15]) );
  CFD2QXL \out1_stg1_reg[14]  ( .D(n857), .CP(clk), .CD(n1312), .Q(
        out1_stg1[14]) );
  CFD2QXL \out1_stg1_reg[13]  ( .D(n855), .CP(clk), .CD(n1312), .Q(
        out1_stg1[13]) );
  CFD2QXL \out1_stg1_reg[12]  ( .D(n853), .CP(clk), .CD(n1312), .Q(
        out1_stg1[12]) );
  CFD2QXL \out1_stg1_reg[11]  ( .D(n851), .CP(clk), .CD(n1313), .Q(
        out1_stg1[11]) );
  CFD2QXL \out1_stg1_reg[10]  ( .D(n849), .CP(clk), .CD(n1313), .Q(
        out1_stg1[10]) );
  CFD2QXL \out1_stg1_reg[9]  ( .D(n847), .CP(clk), .CD(n1313), .Q(out1_stg1[9]) );
  CFD2QXL \out1_stg1_reg[8]  ( .D(n845), .CP(clk), .CD(n1313), .Q(out1_stg1[8]) );
  CFD2QXL \out1_stg1_reg[7]  ( .D(n843), .CP(clk), .CD(n1313), .Q(out1_stg1[7]) );
  CFD2QXL \out1_stg1_reg[6]  ( .D(n841), .CP(clk), .CD(n1313), .Q(out1_stg1[6]) );
  CFD2QXL \out1_stg1_reg[5]  ( .D(n839), .CP(clk), .CD(n1314), .Q(out1_stg1[5]) );
  CFD2QXL \out1_stg1_reg[4]  ( .D(n837), .CP(clk), .CD(n1314), .Q(out1_stg1[4]) );
  CFD2QXL \out1_stg1_reg[3]  ( .D(n835), .CP(clk), .CD(n1314), .Q(out1_stg1[3]) );
  CFD2QXL \out1_stg1_reg[2]  ( .D(n833), .CP(clk), .CD(n1314), .Q(out1_stg1[2]) );
  CFD2QXL \out1_stg1_reg[1]  ( .D(n831), .CP(clk), .CD(n1314), .Q(out1_stg1[1]) );
  CFD2QXL \out1_stg1_reg[0]  ( .D(n829), .CP(clk), .CD(n1314), .Q(out1_stg1[0]) );
  CFD2QXL \out0_stg2_reg[0]  ( .D(n754), .CP(clk), .CD(n1338), .Q(out0_stg2[0]) );
  CFD2QXL \out0_stg2_reg[1]  ( .D(n753), .CP(clk), .CD(n1338), .Q(out0_stg2[1]) );
  CFD2QXL \out0_stg2_reg[2]  ( .D(n752), .CP(clk), .CD(n1338), .Q(out0_stg2[2]) );
  CFD2QXL \out0_stg2_reg[3]  ( .D(n751), .CP(clk), .CD(n1343), .Q(out0_stg2[3]) );
  CFD2QXL \out0_stg2_reg[4]  ( .D(n750), .CP(clk), .CD(n1337), .Q(out0_stg2[4]) );
  CFD2QXL \out0_stg2_reg[5]  ( .D(n749), .CP(clk), .CD(n1337), .Q(out0_stg2[5]) );
  CFD2QXL \out0_stg2_reg[6]  ( .D(n748), .CP(clk), .CD(n1336), .Q(out0_stg2[6]) );
  CFD2QXL \out0_stg2_reg[7]  ( .D(n747), .CP(clk), .CD(n1336), .Q(out0_stg2[7]) );
  CFD2QXL \out0_stg2_reg[8]  ( .D(n746), .CP(clk), .CD(n1335), .Q(out0_stg2[8]) );
  CFD2QXL \out0_stg2_reg[9]  ( .D(n745), .CP(clk), .CD(n1335), .Q(out0_stg2[9]) );
  CFD2QXL \out0_stg2_reg[10]  ( .D(n744), .CP(clk), .CD(n1335), .Q(
        out0_stg2[10]) );
  CFD2QXL \out0_stg2_reg[11]  ( .D(n743), .CP(clk), .CD(n1334), .Q(
        out0_stg2[11]) );
  CFD2QXL \out0_stg2_reg[12]  ( .D(n742), .CP(clk), .CD(n1334), .Q(
        out0_stg2[12]) );
  CFD2QXL \out0_stg2_reg[13]  ( .D(n741), .CP(clk), .CD(n1333), .Q(
        out0_stg2[13]) );
  CFD2QXL \out0_stg2_reg[14]  ( .D(n740), .CP(clk), .CD(n1333), .Q(
        out0_stg2[14]) );
  CFD2QXL \out0_stg2_reg[15]  ( .D(n739), .CP(clk), .CD(n1333), .Q(
        out0_stg2[15]) );
  CFD2QXL \out0_stg2_reg[16]  ( .D(n738), .CP(clk), .CD(n1332), .Q(
        out0_stg2[16]) );
  CFD2QXL \out0_stg2_reg[17]  ( .D(n737), .CP(clk), .CD(n1332), .Q(
        out0_stg2[17]) );
  CFD2QXL \out0_stg2_reg[18]  ( .D(n736), .CP(clk), .CD(n1332), .Q(
        out0_stg2[18]) );
  CFD2QXL \out0_stg2_reg[19]  ( .D(n735), .CP(clk), .CD(n1337), .Q(
        out0_stg2[19]) );
  CFD2QXL \out0_stg2_reg[20]  ( .D(n734), .CP(clk), .CD(n1355), .Q(
        out0_stg2[20]) );
  CFD2QXL \out0_stg2_reg[21]  ( .D(n733), .CP(clk), .CD(n1355), .Q(
        out0_stg2[21]) );
  CFD2QXL \out0_stg2_reg[22]  ( .D(n732), .CP(clk), .CD(n1355), .Q(
        out0_stg2[22]) );
  CFD2QXL \out0_stg2_reg[23]  ( .D(n731), .CP(clk), .CD(n1354), .Q(
        out0_stg2[23]) );
  CFD2QXL \out0_stg2_reg[24]  ( .D(n730), .CP(clk), .CD(n1354), .Q(
        out0_stg2[24]) );
  CFD2QXL \out0_stg2_reg[25]  ( .D(n729), .CP(clk), .CD(n1353), .Q(
        out0_stg2[25]) );
  CFD2QXL \out0_stg2_reg[26]  ( .D(n728), .CP(clk), .CD(n1353), .Q(
        out0_stg2[26]) );
  CFD2QXL \out0_stg2_reg[27]  ( .D(n727), .CP(clk), .CD(n1353), .Q(
        out0_stg2[27]) );
  CFD2QXL \out0_stg2_reg[28]  ( .D(n726), .CP(clk), .CD(n1352), .Q(
        out0_stg2[28]) );
  CFD2QXL \out0_stg2_reg[29]  ( .D(n725), .CP(clk), .CD(n1352), .Q(
        out0_stg2[29]) );
  CFD2QXL \out0_stg2_reg[30]  ( .D(n724), .CP(clk), .CD(n1352), .Q(
        out0_stg2[30]) );
  CFD2QXL \out0_stg2_reg[31]  ( .D(n723), .CP(clk), .CD(n1351), .Q(
        out0_stg2[31]) );
  CFD2QXL \out0_stg2_reg[32]  ( .D(n722), .CP(clk), .CD(n1351), .Q(
        out0_stg2[32]) );
  CFD2QXL \out0_stg2_reg[33]  ( .D(n721), .CP(clk), .CD(n1350), .Q(
        out0_stg2[33]) );
  CFD2QXL \out0_stg2_reg[34]  ( .D(n720), .CP(clk), .CD(n1350), .Q(
        out0_stg2[34]) );
  CFD2QXL \out0_stg2_reg[35]  ( .D(n719), .CP(clk), .CD(n1350), .Q(
        out0_stg2[35]) );
  CFD2QXL \out0_stg2_reg[36]  ( .D(n718), .CP(clk), .CD(n1349), .Q(
        out0_stg2[36]) );
  CFD2QXL \out0_stg2_reg[37]  ( .D(n717), .CP(clk), .CD(n1349), .Q(
        out0_stg2[37]) );
  CFD2QXL \out0_stg2_reg[38]  ( .D(n716), .CP(clk), .CD(n1348), .Q(
        out0_stg2[38]) );
  CFD2QXL \out0_stg2_reg[39]  ( .D(n715), .CP(clk), .CD(n1348), .Q(
        out0_stg2[39]) );
  CFD2QXL \out0_stg2_reg[40]  ( .D(n714), .CP(clk), .CD(n1348), .Q(
        out0_stg2[40]) );
  CFD2QXL \out0_stg2_reg[41]  ( .D(n713), .CP(clk), .CD(n1347), .Q(
        out0_stg2[41]) );
  CFD2QXL \out0_stg2_reg[42]  ( .D(n712), .CP(clk), .CD(n1347), .Q(
        out0_stg2[42]) );
  CFD2QXL \out0_stg2_reg[43]  ( .D(n711), .CP(clk), .CD(n1346), .Q(
        out0_stg2[43]) );
  CFD2QXL \out0_stg2_reg[44]  ( .D(n710), .CP(clk), .CD(n1346), .Q(
        out0_stg2[44]) );
  CFD2QXL \out0_stg2_reg[45]  ( .D(n709), .CP(clk), .CD(n1346), .Q(
        out0_stg2[45]) );
  CFD2QXL \out0_stg2_reg[46]  ( .D(n708), .CP(clk), .CD(n1345), .Q(
        out0_stg2[46]) );
  CFD2QXL \out0_stg2_reg[47]  ( .D(n707), .CP(clk), .CD(n1345), .Q(
        out0_stg2[47]) );
  CFD2QXL \out0_stg2_reg[48]  ( .D(n706), .CP(clk), .CD(n1345), .Q(
        out0_stg2[48]) );
  CFD2QXL \out0_stg2_reg[49]  ( .D(n705), .CP(clk), .CD(n1344), .Q(
        out0_stg2[49]) );
  CFD2QXL \out0_stg2_reg[50]  ( .D(n704), .CP(clk), .CD(n1344), .Q(
        out0_stg2[50]) );
  CFD2QXL \out0_stg2_reg[51]  ( .D(n703), .CP(clk), .CD(n1319), .Q(
        out0_stg2[51]) );
  CFD2QXL \out0_stg2_reg[52]  ( .D(n702), .CP(clk), .CD(n1319), .Q(
        out0_stg2[52]) );
  CFD2QXL \out0_stg2_reg[53]  ( .D(n701), .CP(clk), .CD(n1318), .Q(
        out0_stg2[53]) );
  CFD2QXL \out0_stg2_reg[54]  ( .D(n700), .CP(clk), .CD(n1318), .Q(
        out0_stg2[54]) );
  CFD2QXL \out0_stg2_reg[55]  ( .D(n699), .CP(clk), .CD(n1317), .Q(
        out0_stg2[55]) );
  CFD2QXL \out0_stg2_reg[56]  ( .D(n698), .CP(clk), .CD(n1317), .Q(
        out0_stg2[56]) );
  CFD2QXL \out0_stg2_reg[57]  ( .D(n697), .CP(clk), .CD(n1317), .Q(
        out0_stg2[57]) );
  CFD2QXL \out0_stg2_reg[58]  ( .D(n696), .CP(clk), .CD(n1316), .Q(
        out0_stg2[58]) );
  CFD2QXL \out0_stg2_reg[59]  ( .D(n695), .CP(clk), .CD(n1316), .Q(
        out0_stg2[59]) );
  CFD2QXL \out0_stg2_reg[60]  ( .D(n694), .CP(clk), .CD(n1316), .Q(
        out0_stg2[60]) );
  CFD2QXL \out0_stg2_reg[61]  ( .D(n693), .CP(clk), .CD(n1315), .Q(
        out0_stg2[61]) );
  CFD2QXL \out0_stg2_reg[62]  ( .D(n692), .CP(clk), .CD(n1315), .Q(
        out0_stg2[62]) );
  CFD2QXL \out1_stg2_reg[0]  ( .D(n545), .CP(clk), .CD(n1339), .Q(out1_stg2[0]) );
  CFD2QXL \out1_stg2_reg[1]  ( .D(n543), .CP(clk), .CD(n1338), .Q(out1_stg2[1]) );
  CFD2QXL \out1_stg2_reg[2]  ( .D(n541), .CP(clk), .CD(n1338), .Q(out1_stg2[2]) );
  CFD2QXL \out1_stg2_reg[3]  ( .D(n539), .CP(clk), .CD(n1337), .Q(out1_stg2[3]) );
  CFD2QXL \out1_stg2_reg[4]  ( .D(n537), .CP(clk), .CD(n1337), .Q(out1_stg2[4]) );
  CFD2QXL \out1_stg2_reg[5]  ( .D(n535), .CP(clk), .CD(n1337), .Q(out1_stg2[5]) );
  CFD2QXL \out1_stg2_reg[6]  ( .D(n533), .CP(clk), .CD(n1336), .Q(out1_stg2[6]) );
  CFD2QXL \out1_stg2_reg[7]  ( .D(n531), .CP(clk), .CD(n1336), .Q(out1_stg2[7]) );
  CFD2QXL \out1_stg2_reg[8]  ( .D(n529), .CP(clk), .CD(n1335), .Q(out1_stg2[8]) );
  CFD2QXL \out1_stg2_reg[9]  ( .D(n527), .CP(clk), .CD(n1335), .Q(out1_stg2[9]) );
  CFD2QXL \out1_stg2_reg[16]  ( .D(n513), .CP(clk), .CD(n1332), .Q(
        out1_stg2[16]) );
  CFD2QXL \acc_reg[0]  ( .D(n544), .CP(clk), .CD(n1339), .Q(acc[0]) );
  CFD2QXL \acc_reg[1]  ( .D(n542), .CP(clk), .CD(n1338), .Q(acc[1]) );
  CFD2QXL \acc_reg[2]  ( .D(n540), .CP(clk), .CD(n1338), .Q(acc[2]) );
  CFD2QXL \acc_reg[3]  ( .D(n538), .CP(clk), .CD(n1337), .Q(acc[3]) );
  CFD2QXL \acc_reg[4]  ( .D(n536), .CP(clk), .CD(n1337), .Q(acc[4]) );
  CFD2QXL \acc_reg[5]  ( .D(n534), .CP(clk), .CD(n1337), .Q(acc[5]) );
  CFD2QXL \acc_reg[6]  ( .D(n532), .CP(clk), .CD(n1336), .Q(acc[6]) );
  CFD2QXL \acc_reg[7]  ( .D(n530), .CP(clk), .CD(n1336), .Q(acc[7]) );
  CFD2QXL \acc_reg[8]  ( .D(n528), .CP(clk), .CD(n1336), .Q(acc[8]) );
  CFD2QXL \acc_reg[9]  ( .D(n526), .CP(clk), .CD(n1335), .Q(acc[9]) );
  CFD2QXL \acc_reg[10]  ( .D(n524), .CP(clk), .CD(n1335), .Q(acc[10]) );
  CFD2QXL \acc_reg[11]  ( .D(n522), .CP(clk), .CD(n1334), .Q(acc[11]) );
  CFD2QXL \acc_reg[12]  ( .D(n520), .CP(clk), .CD(n1334), .Q(acc[12]) );
  CFD2QXL \acc_reg[13]  ( .D(n518), .CP(clk), .CD(n1334), .Q(acc[13]) );
  CFD2QXL \acc_reg[14]  ( .D(n516), .CP(clk), .CD(n1333), .Q(acc[14]) );
  CFD2QXL \acc_reg[15]  ( .D(n514), .CP(clk), .CD(n1333), .Q(acc[15]) );
  CFD2QXL \acc_reg[16]  ( .D(n512), .CP(clk), .CD(n1332), .Q(acc[16]) );
  CFD2QXL \acc_reg[17]  ( .D(n510), .CP(clk), .CD(n1332), .Q(acc[17]) );
  CFD2QXL \acc_reg[18]  ( .D(n508), .CP(clk), .CD(n1332), .Q(acc[18]) );
  CFD2QXL \acc_reg[19]  ( .D(n506), .CP(clk), .CD(n1331), .Q(acc[19]) );
  CFD2QXL \acc_reg[20]  ( .D(n504), .CP(clk), .CD(n1356), .Q(acc[20]) );
  CFD2QXL \acc_reg[21]  ( .D(n502), .CP(clk), .CD(n1355), .Q(acc[21]) );
  CFD2QXL \acc_reg[22]  ( .D(n500), .CP(clk), .CD(n1355), .Q(acc[22]) );
  CFD2QXL \acc_reg[23]  ( .D(n498), .CP(clk), .CD(n1354), .Q(acc[23]) );
  CFD2QXL \acc_reg[24]  ( .D(n496), .CP(clk), .CD(n1354), .Q(acc[24]) );
  CFD2QXL \acc_reg[25]  ( .D(n494), .CP(clk), .CD(n1354), .Q(acc[25]) );
  CFD2QXL \acc_reg[26]  ( .D(n492), .CP(clk), .CD(n1353), .Q(acc[26]) );
  CFD2QXL \acc_reg[27]  ( .D(n490), .CP(clk), .CD(n1353), .Q(acc[27]) );
  CFD2QXL \acc_reg[28]  ( .D(n488), .CP(clk), .CD(n1352), .Q(acc[28]) );
  CFD2QXL \acc_reg[29]  ( .D(n486), .CP(clk), .CD(n1352), .Q(acc[29]) );
  CFD2QXL \acc_reg[30]  ( .D(n484), .CP(clk), .CD(n1352), .Q(acc[30]) );
  CFD2QXL \acc_reg[31]  ( .D(n482), .CP(clk), .CD(n1351), .Q(acc[31]) );
  CFD2QXL \out2_stg2_reg[56]  ( .D(n554), .CP(clk), .CD(n1324), .Q(
        out2_stg2[56]) );
  CFD2QXL \out2_stg2_reg[1]  ( .D(n609), .CP(clk), .CD(n1329), .Q(out2_stg2[1]) );
  CFD2QXL \out2_stg2_reg[3]  ( .D(n607), .CP(clk), .CD(n1328), .Q(out2_stg2[3]) );
  CFD2QXL \out2_stg2_reg[9]  ( .D(n601), .CP(clk), .CD(n1328), .Q(out2_stg2[9]) );
  CFD2QXL \out2_stg2_reg[11]  ( .D(n599), .CP(clk), .CD(n1328), .Q(
        out2_stg2[11]) );
  CFD2QXL \out2_stg2_reg[13]  ( .D(n597), .CP(clk), .CD(n1328), .Q(
        out2_stg2[13]) );
  CFD2QXL \out2_stg2_reg[15]  ( .D(n595), .CP(clk), .CD(n1327), .Q(
        out2_stg2[15]) );
  CFD2QXL \out2_stg2_reg[33]  ( .D(n577), .CP(clk), .CD(n1326), .Q(
        out2_stg2[33]) );
  CFD2QXL \out2_stg2_reg[35]  ( .D(n575), .CP(clk), .CD(n1326), .Q(
        out2_stg2[35]) );
  CFD2QXL \out2_stg2_reg[37]  ( .D(n573), .CP(clk), .CD(n1326), .Q(
        out2_stg2[37]) );
  CFD2QXL \out2_stg2_reg[39]  ( .D(n571), .CP(clk), .CD(n1326), .Q(
        out2_stg2[39]) );
  CFD2QXL \out2_stg2_reg[41]  ( .D(n569), .CP(clk), .CD(n1325), .Q(
        out2_stg2[41]) );
  CFD2QXL \out2_stg2_reg[43]  ( .D(n567), .CP(clk), .CD(n1325), .Q(
        out2_stg2[43]) );
  CFD2QXL \out2_stg2_reg[45]  ( .D(n565), .CP(clk), .CD(n1325), .Q(
        out2_stg2[45]) );
  CFD2QXL \out2_stg2_reg[47]  ( .D(n563), .CP(clk), .CD(n1325), .Q(
        out2_stg2[47]) );
  CFD2QXL \out2_stg2_reg[49]  ( .D(n561), .CP(clk), .CD(n1325), .Q(
        out2_stg2[49]) );
  CFD2QXL \out2_stg2_reg[51]  ( .D(n559), .CP(clk), .CD(n1325), .Q(
        out2_stg2[51]) );
  CFD2QXL \out2_stg2_reg[53]  ( .D(n557), .CP(clk), .CD(n1324), .Q(
        out2_stg2[53]) );
  CFD2QXL \out2_stg2_reg[55]  ( .D(n555), .CP(clk), .CD(n1324), .Q(
        out2_stg2[55]) );
  CFD2QXL \out2_stg2_reg[2]  ( .D(n608), .CP(clk), .CD(n1328), .Q(out2_stg2[2]) );
  CFD2QXL \out2_stg2_reg[4]  ( .D(n606), .CP(clk), .CD(n1328), .Q(out2_stg2[4]) );
  CFD2QXL \out2_stg2_reg[6]  ( .D(n604), .CP(clk), .CD(n1328), .Q(out2_stg2[6]) );
  CFD2QXL \out2_stg2_reg[8]  ( .D(n602), .CP(clk), .CD(n1328), .Q(out2_stg2[8]) );
  CFD2QXL \out2_stg2_reg[10]  ( .D(n600), .CP(clk), .CD(n1328), .Q(
        out2_stg2[10]) );
  CFD2QXL \out2_stg2_reg[12]  ( .D(n598), .CP(clk), .CD(n1328), .Q(
        out2_stg2[12]) );
  CFD2QXL \out2_stg2_reg[14]  ( .D(n596), .CP(clk), .CD(n1328), .Q(
        out2_stg2[14]) );
  CFD2QXL \out2_stg2_reg[16]  ( .D(n594), .CP(clk), .CD(n1327), .Q(
        out2_stg2[16]) );
  CFD2QXL \out2_stg2_reg[18]  ( .D(n592), .CP(clk), .CD(n1327), .Q(
        out2_stg2[18]) );
  CFD2QXL \out2_stg2_reg[20]  ( .D(n590), .CP(clk), .CD(n1327), .Q(
        out2_stg2[20]) );
  CFD2QXL \out2_stg2_reg[22]  ( .D(n588), .CP(clk), .CD(n1327), .Q(
        out2_stg2[22]) );
  CFD2QXL \out2_stg2_reg[24]  ( .D(n586), .CP(clk), .CD(n1327), .Q(
        out2_stg2[24]) );
  CFD2QXL \out2_stg2_reg[26]  ( .D(n584), .CP(clk), .CD(n1327), .Q(
        out2_stg2[26]) );
  CFD2QXL \out2_stg2_reg[28]  ( .D(n582), .CP(clk), .CD(n1326), .Q(
        out2_stg2[28]) );
  CFD2QXL \out2_stg2_reg[30]  ( .D(n580), .CP(clk), .CD(n1326), .Q(
        out2_stg2[30]) );
  CFD2QXL \out2_stg2_reg[32]  ( .D(n578), .CP(clk), .CD(n1326), .Q(
        out2_stg2[32]) );
  CFD2QXL \out2_stg2_reg[34]  ( .D(n576), .CP(clk), .CD(n1326), .Q(
        out2_stg2[34]) );
  CFD2QXL \out2_stg2_reg[36]  ( .D(n574), .CP(clk), .CD(n1326), .Q(
        out2_stg2[36]) );
  CFD2QXL \out2_stg2_reg[38]  ( .D(n572), .CP(clk), .CD(n1326), .Q(
        out2_stg2[38]) );
  CFD2QXL \out2_stg2_reg[40]  ( .D(n570), .CP(clk), .CD(n1326), .Q(
        out2_stg2[40]) );
  CFD2QXL \out2_stg2_reg[42]  ( .D(n568), .CP(clk), .CD(n1325), .Q(
        out2_stg2[42]) );
  CFD2QXL \out2_stg2_reg[44]  ( .D(n566), .CP(clk), .CD(n1325), .Q(
        out2_stg2[44]) );
  CFD2QXL \out2_stg2_reg[46]  ( .D(n564), .CP(clk), .CD(n1325), .Q(
        out2_stg2[46]) );
  CFD2QXL \out2_stg2_reg[48]  ( .D(n562), .CP(clk), .CD(n1325), .Q(
        out2_stg2[48]) );
  CFD2QXL \out2_stg2_reg[50]  ( .D(n560), .CP(clk), .CD(n1325), .Q(
        out2_stg2[50]) );
  CFD2QXL \out2_stg2_reg[52]  ( .D(n558), .CP(clk), .CD(n1325), .Q(
        out2_stg2[52]) );
  CFD2QXL \out2_stg2_reg[54]  ( .D(n556), .CP(clk), .CD(n1324), .Q(
        out2_stg2[54]) );
  CFD2QXL \out2_stg2_reg[0]  ( .D(n828), .CP(clk), .CD(n1329), .Q(out2_stg2[0]) );
  CFD2QXL \out2_stg2_reg[5]  ( .D(n605), .CP(clk), .CD(n1328), .Q(out2_stg2[5]) );
  CFD2QXL \out2_stg2_reg[7]  ( .D(n603), .CP(clk), .CD(n1328), .Q(out2_stg2[7]) );
  CFD2QXL \out2_stg2_reg[17]  ( .D(n593), .CP(clk), .CD(n1327), .Q(
        out2_stg2[17]) );
  CFD2QXL \out2_stg2_reg[19]  ( .D(n591), .CP(clk), .CD(n1327), .Q(
        out2_stg2[19]) );
  CFD2QXL \out2_stg2_reg[21]  ( .D(n589), .CP(clk), .CD(n1327), .Q(
        out2_stg2[21]) );
  CFD2QXL \out2_stg2_reg[23]  ( .D(n587), .CP(clk), .CD(n1327), .Q(
        out2_stg2[23]) );
  CFD2QXL \out2_stg2_reg[25]  ( .D(n585), .CP(clk), .CD(n1327), .Q(
        out2_stg2[25]) );
  CFD2QXL \out2_stg2_reg[27]  ( .D(n583), .CP(clk), .CD(n1327), .Q(
        out2_stg2[27]) );
  CFD2QXL \out2_stg2_reg[29]  ( .D(n581), .CP(clk), .CD(n1326), .Q(
        out2_stg2[29]) );
  CFD2QXL \out2_stg2_reg[31]  ( .D(n579), .CP(clk), .CD(n1326), .Q(
        out2_stg2[31]) );
  CFD2QXL _pushout_reg ( .D(n808), .CP(clk), .CD(n1340), .Q(pushout) );
  CFD2QXL \out0_stg0_reg[63]  ( .D(N78), .CP(clk), .CD(n1323), .Q(
        out0_stg0[63]) );
  CFD2QXL \out0_stg0_reg[41]  ( .D(N56), .CP(clk), .CD(n1347), .Q(
        out0_stg0[41]) );
  CFD2QXL \out0_stg0_reg[40]  ( .D(N55), .CP(clk), .CD(n1347), .Q(
        out0_stg0[40]) );
  CFD2QXL \out0_stg0_reg[39]  ( .D(N54), .CP(clk), .CD(n1348), .Q(
        out0_stg0[39]) );
  CFD2QXL \out0_stg0_reg[38]  ( .D(N53), .CP(clk), .CD(n1348), .Q(
        out0_stg0[38]) );
  CFD2QXL \out0_stg0_reg[37]  ( .D(N52), .CP(clk), .CD(n1349), .Q(
        out0_stg0[37]) );
  CFD2QXL \out0_stg0_reg[36]  ( .D(N51), .CP(clk), .CD(n1349), .Q(
        out0_stg0[36]) );
  CFD2QXL \out0_stg0_reg[35]  ( .D(N50), .CP(clk), .CD(n1349), .Q(
        out0_stg0[35]) );
  CFD2QXL \out0_stg0_reg[34]  ( .D(N49), .CP(clk), .CD(n1350), .Q(
        out0_stg0[34]) );
  CFD2QXL \out0_stg0_reg[33]  ( .D(N48), .CP(clk), .CD(n1350), .Q(
        out0_stg0[33]) );
  CFD2QXL \out0_stg0_reg[32]  ( .D(N47), .CP(clk), .CD(n1351), .Q(
        out0_stg0[32]) );
  CFD2QXL \out0_stg0_reg[31]  ( .D(N46), .CP(clk), .CD(n1351), .Q(
        out0_stg0[31]) );
  CFD2QXL \out0_stg0_reg[30]  ( .D(N45), .CP(clk), .CD(n1351), .Q(
        out0_stg0[30]) );
  CFD2QXL \out0_stg0_reg[29]  ( .D(N44), .CP(clk), .CD(n1352), .Q(
        out0_stg0[29]) );
  CFD2QXL \out0_stg0_reg[28]  ( .D(N43), .CP(clk), .CD(n1352), .Q(
        out0_stg0[28]) );
  CFD2QXL \out0_stg0_reg[27]  ( .D(N42), .CP(clk), .CD(n1353), .Q(
        out0_stg0[27]) );
  CFD2QXL \out0_stg0_reg[26]  ( .D(N41), .CP(clk), .CD(n1353), .Q(
        out0_stg0[26]) );
  CFD2QXL \out0_stg0_reg[25]  ( .D(N40), .CP(clk), .CD(n1353), .Q(
        out0_stg0[25]) );
  CFD2QXL \out0_stg0_reg[24]  ( .D(N39), .CP(clk), .CD(n1354), .Q(
        out0_stg0[24]) );
  CFD2QXL \out0_stg0_reg[23]  ( .D(N38), .CP(clk), .CD(n1354), .Q(
        out0_stg0[23]) );
  CFD2QXL \out0_stg0_reg[22]  ( .D(N37), .CP(clk), .CD(n1354), .Q(
        out0_stg0[22]) );
  CFD2QXL \out0_stg0_reg[21]  ( .D(N36), .CP(clk), .CD(n1355), .Q(
        out0_stg0[21]) );
  CFD2QXL \out0_stg0_reg[20]  ( .D(N35), .CP(clk), .CD(n1355), .Q(
        out0_stg0[20]) );
  CFD2QXL \out0_stg0_reg[19]  ( .D(N34), .CP(clk), .CD(n1356), .Q(
        out0_stg0[19]) );
  CFD2QXL \out0_stg0_reg[18]  ( .D(N33), .CP(clk), .CD(n1331), .Q(
        out0_stg0[18]) );
  CFD2QXL \out0_stg0_reg[17]  ( .D(N32), .CP(clk), .CD(n1332), .Q(
        out0_stg0[17]) );
  CFD2QXL \out0_stg0_reg[16]  ( .D(N31), .CP(clk), .CD(n1332), .Q(
        out0_stg0[16]) );
  CFD2QXL \out0_stg0_reg[14]  ( .D(N29), .CP(clk), .CD(n1333), .Q(
        out0_stg0[14]) );
  CFD2QXL \out0_stg0_reg[9]  ( .D(N24), .CP(clk), .CD(n1335), .Q(out0_stg0[9])
         );
  CFD2QXL \out0_stg0_reg[8]  ( .D(N23), .CP(clk), .CD(n1335), .Q(out0_stg0[8])
         );
  CFD2QXL \out0_stg0_reg[7]  ( .D(N22), .CP(clk), .CD(n1336), .Q(out0_stg0[7])
         );
  CFD2QXL \out0_stg0_reg[6]  ( .D(N21), .CP(clk), .CD(n1336), .Q(out0_stg0[6])
         );
  CFD2QXL \out0_stg0_reg[5]  ( .D(N20), .CP(clk), .CD(n1336), .Q(out0_stg0[5])
         );
  CFD2QXL \out0_stg0_reg[4]  ( .D(N19), .CP(clk), .CD(n1337), .Q(out0_stg0[4])
         );
  CFD2QXL \out0_stg0_reg[3]  ( .D(N18), .CP(clk), .CD(n1337), .Q(out0_stg0[3])
         );
  CFD2QXL \out0_stg0_reg[2]  ( .D(N17), .CP(clk), .CD(n1338), .Q(out0_stg0[2])
         );
  CFD2QXL \out0_stg0_reg[1]  ( .D(N16), .CP(clk), .CD(n1338), .Q(out0_stg0[1])
         );
  CFD2QXL \out0_stg0_reg[0]  ( .D(N15), .CP(clk), .CD(n1338), .Q(out0_stg0[0])
         );
  CFD2QXL \out1_stg0_reg[63]  ( .D(N78), .CP(clk), .CD(n1329), .Q(
        out1_stg0[63]) );
  CFD2QXL \out1_stg0_reg[41]  ( .D(N56), .CP(clk), .CD(n1308), .Q(
        out1_stg0[41]) );
  CFD2QXL \out1_stg0_reg[40]  ( .D(N55), .CP(clk), .CD(n1308), .Q(
        out1_stg0[40]) );
  CFD2QXL \out1_stg0_reg[39]  ( .D(N54), .CP(clk), .CD(n1308), .Q(
        out1_stg0[39]) );
  CFD2QXL \out1_stg0_reg[38]  ( .D(N53), .CP(clk), .CD(n1308), .Q(
        out1_stg0[38]) );
  CFD2QXL \out1_stg0_reg[37]  ( .D(N52), .CP(clk), .CD(n1308), .Q(
        out1_stg0[37]) );
  CFD2QXL \out1_stg0_reg[36]  ( .D(N51), .CP(clk), .CD(n1309), .Q(
        out1_stg0[36]) );
  CFD2QXL \out1_stg0_reg[35]  ( .D(N50), .CP(clk), .CD(n1309), .Q(
        out1_stg0[35]) );
  CFD2QXL \out1_stg0_reg[34]  ( .D(N49), .CP(clk), .CD(n1309), .Q(
        out1_stg0[34]) );
  CFD2QXL \out1_stg0_reg[33]  ( .D(N48), .CP(clk), .CD(n1309), .Q(
        out1_stg0[33]) );
  CFD2QXL \out1_stg0_reg[32]  ( .D(N47), .CP(clk), .CD(n1309), .Q(
        out1_stg0[32]) );
  CFD2QXL \out1_stg0_reg[31]  ( .D(N46), .CP(clk), .CD(n1309), .Q(
        out1_stg0[31]) );
  CFD2QXL \out1_stg0_reg[30]  ( .D(N45), .CP(clk), .CD(n1310), .Q(
        out1_stg0[30]) );
  CFD2QXL \out1_stg0_reg[29]  ( .D(N44), .CP(clk), .CD(n1310), .Q(
        out1_stg0[29]) );
  CFD2QXL \out1_stg0_reg[28]  ( .D(N43), .CP(clk), .CD(n1310), .Q(
        out1_stg0[28]) );
  CFD2QXL \out1_stg0_reg[27]  ( .D(N42), .CP(clk), .CD(n1310), .Q(
        out1_stg0[27]) );
  CFD2QXL \out1_stg0_reg[26]  ( .D(N41), .CP(clk), .CD(n1310), .Q(
        out1_stg0[26]) );
  CFD2QXL \out1_stg0_reg[25]  ( .D(N40), .CP(clk), .CD(n1310), .Q(
        out1_stg0[25]) );
  CFD2QXL \out1_stg0_reg[24]  ( .D(N39), .CP(clk), .CD(n1310), .Q(
        out1_stg0[24]) );
  CFD2QXL \out1_stg0_reg[23]  ( .D(N38), .CP(clk), .CD(n1311), .Q(
        out1_stg0[23]) );
  CFD2QXL \out1_stg0_reg[22]  ( .D(N37), .CP(clk), .CD(n1311), .Q(
        out1_stg0[22]) );
  CFD2QXL \out1_stg0_reg[21]  ( .D(N36), .CP(clk), .CD(n1311), .Q(
        out1_stg0[21]) );
  CFD2QXL \out1_stg0_reg[20]  ( .D(N35), .CP(clk), .CD(n1311), .Q(
        out1_stg0[20]) );
  CFD2QXL \out1_stg0_reg[19]  ( .D(N34), .CP(clk), .CD(n1311), .Q(
        out1_stg0[19]) );
  CFD2QXL \out1_stg0_reg[18]  ( .D(N33), .CP(clk), .CD(n1311), .Q(
        out1_stg0[18]) );
  CFD2QXL \out1_stg0_reg[17]  ( .D(N32), .CP(clk), .CD(n1312), .Q(
        out1_stg0[17]) );
  CFD2QXL \out1_stg0_reg[16]  ( .D(N31), .CP(clk), .CD(n1312), .Q(
        out1_stg0[16]) );
  CFD2QXL \out1_stg0_reg[14]  ( .D(N29), .CP(clk), .CD(n1312), .Q(
        out1_stg0[14]) );
  CFD2QXL \out1_stg0_reg[9]  ( .D(N24), .CP(clk), .CD(n1313), .Q(out1_stg0[9])
         );
  CFD2QXL \out1_stg0_reg[8]  ( .D(N23), .CP(clk), .CD(n1313), .Q(out1_stg0[8])
         );
  CFD2QXL \out1_stg0_reg[7]  ( .D(N22), .CP(clk), .CD(n1313), .Q(out1_stg0[7])
         );
  CFD2QXL \out1_stg0_reg[6]  ( .D(N21), .CP(clk), .CD(n1313), .Q(out1_stg0[6])
         );
  CFD2QXL \out1_stg0_reg[5]  ( .D(N20), .CP(clk), .CD(n1313), .Q(out1_stg0[5])
         );
  CFD2QXL \out1_stg0_reg[4]  ( .D(N19), .CP(clk), .CD(n1314), .Q(out1_stg0[4])
         );
  CFD2QXL \out1_stg0_reg[3]  ( .D(N18), .CP(clk), .CD(n1314), .Q(out1_stg0[3])
         );
  CFD2QXL \out1_stg0_reg[2]  ( .D(N17), .CP(clk), .CD(n1314), .Q(out1_stg0[2])
         );
  CFD2QXL \out1_stg0_reg[1]  ( .D(N16), .CP(clk), .CD(n1314), .Q(out1_stg0[1])
         );
  CFD2QXL \out1_stg0_reg[0]  ( .D(N15), .CP(clk), .CD(n1314), .Q(out1_stg0[0])
         );
  CFD2QXL \cmd0_stg0_reg[1]  ( .D(n1118), .CP(clk), .CD(n1340), .Q(
        cmd0_stg0[1]) );
  CFD2QXL \cmd0_stg1_reg[1]  ( .D(n1110), .CP(clk), .CD(n1340), .Q(
        cmd0_stg1[1]) );
  CFD2QXL \cmd0_stg0_reg[0]  ( .D(n1120), .CP(clk), .CD(n1340), .Q(
        cmd0_stg0[0]) );
  CFD2QXL \cmd0_stg1_reg[0]  ( .D(n1112), .CP(clk), .CD(n1340), .Q(
        cmd0_stg1[0]) );
  CFD2QXL push0_stg0_reg ( .D(n1122), .CP(clk), .CD(n1340), .Q(push0_stg0) );
  CFD2QXL push0_stg1_reg ( .D(n1114), .CP(clk), .CD(n1340), .Q(push0_stg1) );
  CFD1QXL cmd2_en_stg2_reg ( .D(n690), .CP(clk), .Q(cmd2_en_stg2) );
  CFD2QX1 \q0_reg[21]  ( .D(n1108), .CP(clk), .CD(n1307), .Q(q0[21]) );
  CFD2QX2 \q0_reg[31]  ( .D(n1098), .CP(clk), .CD(n1331), .Q(q0[31]) );
  CFD2QXL cmd1_en_stg2_d_reg ( .D(n1293), .CP(clk), .CD(n1314), .Q(
        cmd1_en_stg2_d) );
  CFD2QXL cmd0_en_stg2_d_reg ( .D(n1255), .CP(clk), .CD(n1315), .Q(
        cmd0_en_stg2_d) );
  CFD2QX2 \h0_reg[1]  ( .D(n617), .CP(clk), .CD(n1323), .Q(h0[1]) );
  CFD2QX1 \h0_reg[5]  ( .D(n629), .CP(clk), .CD(n1323), .Q(h0[5]) );
  CFD2QX1 \h0_reg[6]  ( .D(n632), .CP(clk), .CD(n1323), .Q(h0[6]) );
  CFD2QX1 \h0_reg[12]  ( .D(n638), .CP(clk), .CD(n1322), .Q(h0[12]) );
  CFD2QX2 \h0_reg[3]  ( .D(n623), .CP(clk), .CD(n1323), .Q(h0[3]) );
  CFD2QX1 \h0_reg[10]  ( .D(n636), .CP(clk), .CD(n1323), .Q(h0[10]) );
  CFD2QX2 \h0_reg[8]  ( .D(n816), .CP(clk), .CD(n1323), .Q(h0[8]) );
  CFD2QX1 \h0_reg[2]  ( .D(n620), .CP(clk), .CD(n1323), .Q(h0[2]) );
  CFD2QX2 \h0_reg[18]  ( .D(n813), .CP(clk), .CD(n1322), .Q(h0[18]) );
  CFD2QX2 \h0_reg[9]  ( .D(n814), .CP(clk), .CD(n1323), .Q(h0[9]) );
  CFD2QX1 \h0_reg[29]  ( .D(n819), .CP(clk), .CD(n1321), .Q(h0[29]) );
  CFD2QX1 \h0_reg[20]  ( .D(n821), .CP(clk), .CD(n1322), .Q(h0[20]) );
  CFD2QX2 \h0_reg[21]  ( .D(n822), .CP(clk), .CD(n1322), .Q(h0[21]) );
  CFD2QX2 \h0_reg[22]  ( .D(n820), .CP(clk), .CD(n1322), .Q(h0[22]) );
  CFD2QX1 \h0_reg[13]  ( .D(n817), .CP(clk), .CD(n1322), .Q(h0[13]) );
  CFD2QX1 \h0_reg[11]  ( .D(n823), .CP(clk), .CD(n1322), .Q(h0[11]) );
  CFD2QX1 \h0_reg[7]  ( .D(n633), .CP(clk), .CD(n1323), .Q(h0[7]) );
  CFD2QX1 \h0_reg[26]  ( .D(n652), .CP(clk), .CD(n1321), .Q(h0[26]) );
  CFD2QX1 \h0_reg[27]  ( .D(n824), .CP(clk), .CD(n1321), .Q(h0[27]) );
  CFD2QX1 \h0_reg[25]  ( .D(n825), .CP(clk), .CD(n1321), .Q(h0[25]) );
  CFD2QX1 \h0_reg[28]  ( .D(n654), .CP(clk), .CD(n1321), .Q(h0[28]) );
  CFD2QX1 \h0_reg[14]  ( .D(n818), .CP(clk), .CD(n1322), .Q(h0[14]) );
  CFD2QX1 \h0_reg[19]  ( .D(n826), .CP(clk), .CD(n1322), .Q(h0[19]) );
  CFD2QX2 \q0_reg[14]  ( .D(n672), .CP(clk), .CD(n1320), .Q(q0[14]) );
  CFD2QX1 \q0_reg[23]  ( .D(n809), .CP(clk), .CD(n1307), .Q(q0[23]) );
  CFD2QX1 \q0_reg[9]  ( .D(n810), .CP(clk), .CD(n1320), .Q(q0[9]) );
  CFD2QX1 \q0_reg[3]  ( .D(n661), .CP(clk), .CD(n1321), .Q(q0[3]) );
  CFD2QX1 \h0_reg[15]  ( .D(n641), .CP(clk), .CD(n1322), .Q(h0[15]) );
  CFD2QX4 \q0_reg[6]  ( .D(n664), .CP(clk), .CD(n1320), .Q(q0[6]) );
  CFD2QX1 \q0_reg[5]  ( .D(n663), .CP(clk), .CD(n1321), .Q(q0[5]) );
  CFD2QX1 \h0_reg[16]  ( .D(n812), .CP(clk), .CD(n1322), .Q(h0[16]) );
  CFD2QX1 \h0_reg[23]  ( .D(n811), .CP(clk), .CD(n1322), .Q(h0[23]) );
  CFD2QX1 \h0_reg[30]  ( .D(n827), .CP(clk), .CD(n1321), .Q(h0[30]) );
  CFD2QX1 \h0_reg[24]  ( .D(n1124), .CP(clk), .CD(n1321), .Q(h0[24]) );
  CFD2QX1 \q0_reg[11]  ( .D(n669), .CP(clk), .CD(n1320), .Q(q0[11]) );
  CFD2QX1 \h0_reg[31]  ( .D(n1125), .CP(clk), .CD(n1321), .Q(h0[31]) );
  CFD2QX2 \q0_reg[29]  ( .D(n687), .CP(clk), .CD(n1307), .Q(q0[29]) );
  CFD2QX1 \q0_reg[25]  ( .D(n1117), .CP(clk), .CD(n1319), .Q(q0[25]) );
  CFD2QX4 \q0_reg[4]  ( .D(n662), .CP(clk), .CD(n1321), .Q(q0[4]) );
  CFD2QX4 \q0_reg[28]  ( .D(n686), .CP(clk), .CD(n1325), .Q(q0[28]) );
  CFD2QX4 \q0_reg[24]  ( .D(n682), .CP(clk), .CD(n1319), .Q(q0[24]) );
  CFD1XL cmd0_en_stg2_reg ( .D(n755), .CP(clk), .Q(cmd0_en_stg2), .QN(n1226)
         );
  CFD2XL push0_stg2_reg ( .D(n1102), .CP(clk), .CD(n1973), .Q(push0_stg2), 
        .QN(n1972) );
  CFD2XL \out1_stg2_reg[14]  ( .D(n517), .CP(clk), .CD(n1973), .Q(
        out1_stg2[14]), .QN(n1703) );
  CFD2XL \out1_stg2_reg[12]  ( .D(n521), .CP(clk), .CD(n1973), .Q(
        out1_stg2[12]), .QN(n1711) );
  CFD2XL \out1_stg2_reg[10]  ( .D(n525), .CP(clk), .CD(n1973), .Q(
        out1_stg2[10]), .QN(n1719) );
  CFD2XL \out1_stg0_reg[10]  ( .D(N25), .CP(clk), .CD(n1973), .Q(out1_stg0[10]) );
  CFD2XL \out0_stg0_reg[10]  ( .D(N25), .CP(clk), .CD(n1973), .Q(out0_stg0[10]) );
  CFD2XL \out1_stg2_reg[31]  ( .D(n483), .CP(clk), .CD(n1973), .Q(
        out1_stg2[31]), .QN(n1635) );
  CFD2XL \out1_stg2_reg[30]  ( .D(n485), .CP(clk), .CD(n1973), .Q(
        out1_stg2[30]), .QN(n1639) );
  CFD2XL \out1_stg2_reg[29]  ( .D(n487), .CP(clk), .CD(n1973), .Q(
        out1_stg2[29]), .QN(n1643) );
  CFD2XL \out1_stg2_reg[28]  ( .D(n489), .CP(clk), .CD(n1973), .Q(
        out1_stg2[28]), .QN(n1647) );
  CFD2XL \out1_stg2_reg[27]  ( .D(n491), .CP(clk), .CD(n1973), .Q(
        out1_stg2[27]), .QN(n1651) );
  CFD2XL \out1_stg2_reg[26]  ( .D(n493), .CP(clk), .CD(n1973), .Q(
        out1_stg2[26]), .QN(n1655) );
  CFD2XL \out1_stg2_reg[25]  ( .D(n495), .CP(clk), .CD(n1973), .Q(
        out1_stg2[25]), .QN(n1659) );
  CFD2XL \out1_stg2_reg[24]  ( .D(n497), .CP(clk), .CD(n1973), .Q(
        out1_stg2[24]), .QN(n1663) );
  CFD2XL \out1_stg2_reg[22]  ( .D(n501), .CP(clk), .CD(n1973), .Q(
        out1_stg2[22]), .QN(n1671) );
  CFD2XL \out1_stg2_reg[21]  ( .D(n503), .CP(clk), .CD(n1973), .Q(
        out1_stg2[21]), .QN(n1675) );
  CFD2XL \out1_stg2_reg[20]  ( .D(n505), .CP(clk), .CD(n1973), .Q(
        out1_stg2[20]), .QN(n1679) );
  CFD2XL \out1_stg2_reg[19]  ( .D(n507), .CP(clk), .CD(n1973), .Q(
        out1_stg2[19]), .QN(n1683) );
  CFD2XL \out1_stg2_reg[18]  ( .D(n509), .CP(clk), .CD(n1973), .Q(
        out1_stg2[18]), .QN(n1687) );
  CFD2XL \out1_stg2_reg[17]  ( .D(n511), .CP(clk), .CD(n1973), .Q(
        out1_stg2[17]), .QN(n1691) );
  CFD2XL \out1_stg2_reg[23]  ( .D(n499), .CP(clk), .CD(n1973), .Q(
        out1_stg2[23]), .QN(n1667) );
  CFD2XL \out1_stg0_reg[11]  ( .D(N26), .CP(clk), .CD(n1973), .Q(out1_stg0[11]) );
  CFD2XL \out0_stg0_reg[11]  ( .D(N26), .CP(clk), .CD(n1973), .Q(out0_stg0[11]) );
  CFD2XL \out1_stg2_reg[32]  ( .D(n481), .CP(clk), .CD(n1973), .Q(
        out1_stg2[32]), .QN(n1631) );
  CFD2XL \out1_stg2_reg[15]  ( .D(n515), .CP(clk), .CD(n1973), .Q(
        out1_stg2[15]), .QN(n1699) );
  CFD2XL \out1_stg2_reg[13]  ( .D(n519), .CP(clk), .CD(n1973), .Q(
        out1_stg2[13]), .QN(n1707) );
  CFD2XL \out1_stg2_reg[11]  ( .D(n523), .CP(clk), .CD(n1973), .Q(
        out1_stg2[11]), .QN(n1715) );
  CFD2XL \out1_stg0_reg[13]  ( .D(N28), .CP(clk), .CD(n1973), .Q(out1_stg0[13]) );
  CFD2XL \out0_stg0_reg[13]  ( .D(N28), .CP(clk), .CD(n1973), .Q(out0_stg0[13]) );
  CFD2XL \out1_stg0_reg[15]  ( .D(N30), .CP(clk), .CD(n1973), .Q(out1_stg0[15]) );
  CFD2XL \out0_stg0_reg[15]  ( .D(N30), .CP(clk), .CD(n1973), .Q(out0_stg0[15]) );
  CFD2XL \out1_stg0_reg[12]  ( .D(N27), .CP(clk), .CD(n1973), .Q(out1_stg0[12]) );
  CFD2XL \out0_stg0_reg[12]  ( .D(N27), .CP(clk), .CD(n1973), .Q(out0_stg0[12]) );
  CFD2XL \out1_stg2_reg[63]  ( .D(n419), .CP(clk), .CD(n1973), .Q(
        out1_stg2[63]), .QN(n1505) );
  CFD2XL \out1_stg2_reg[62]  ( .D(n421), .CP(clk), .CD(n1973), .Q(
        out1_stg2[62]), .QN(n1511) );
  CFD2XL \out1_stg2_reg[61]  ( .D(n423), .CP(clk), .CD(n1973), .Q(
        out1_stg2[61]), .QN(n1515) );
  CFD2XL \out1_stg2_reg[60]  ( .D(n425), .CP(clk), .CD(n1973), .Q(
        out1_stg2[60]), .QN(n1519) );
  CFD2XL \out1_stg2_reg[59]  ( .D(n427), .CP(clk), .CD(n1973), .Q(
        out1_stg2[59]), .QN(n1523) );
  CFD2XL \out1_stg2_reg[58]  ( .D(n429), .CP(clk), .CD(n1973), .Q(
        out1_stg2[58]), .QN(n1527) );
  CFD2XL \out1_stg2_reg[57]  ( .D(n431), .CP(clk), .CD(n1973), .Q(
        out1_stg2[57]), .QN(n1531) );
  CFD2XL \out1_stg2_reg[56]  ( .D(n433), .CP(clk), .CD(n1973), .Q(
        out1_stg2[56]), .QN(n1535) );
  CFD2XL \out1_stg2_reg[55]  ( .D(n435), .CP(clk), .CD(n1973), .Q(
        out1_stg2[55]), .QN(n1539) );
  CFD2XL \out1_stg2_reg[54]  ( .D(n437), .CP(clk), .CD(n1973), .Q(
        out1_stg2[54]), .QN(n1543) );
  CFD2XL \out1_stg2_reg[53]  ( .D(n439), .CP(clk), .CD(n1973), .Q(
        out1_stg2[53]), .QN(n1547) );
  CFD2XL \out1_stg2_reg[52]  ( .D(n441), .CP(clk), .CD(n1973), .Q(
        out1_stg2[52]), .QN(n1551) );
  CFD2XL \out1_stg2_reg[51]  ( .D(n443), .CP(clk), .CD(n1973), .Q(
        out1_stg2[51]), .QN(n1555) );
  CFD2XL \out1_stg2_reg[50]  ( .D(n445), .CP(clk), .CD(n1973), .Q(
        out1_stg2[50]), .QN(n1559) );
  CFD2XL \out1_stg2_reg[49]  ( .D(n447), .CP(clk), .CD(n1973), .Q(
        out1_stg2[49]), .QN(n1563) );
  CFD2XL \out1_stg2_reg[48]  ( .D(n449), .CP(clk), .CD(n1973), .Q(
        out1_stg2[48]), .QN(n1567) );
  CFD2XL \out1_stg2_reg[47]  ( .D(n451), .CP(clk), .CD(n1973), .Q(
        out1_stg2[47]), .QN(n1571) );
  CFD2XL \out1_stg2_reg[46]  ( .D(n453), .CP(clk), .CD(n1973), .Q(
        out1_stg2[46]), .QN(n1575) );
  CFD2XL \out1_stg2_reg[45]  ( .D(n455), .CP(clk), .CD(n1973), .Q(
        out1_stg2[45]), .QN(n1579) );
  CFD2XL \out1_stg2_reg[44]  ( .D(n457), .CP(clk), .CD(n1973), .Q(
        out1_stg2[44]), .QN(n1583) );
  CFD2XL \out1_stg2_reg[43]  ( .D(n459), .CP(clk), .CD(n1973), .Q(
        out1_stg2[43]), .QN(n1587) );
  CFD2XL \out1_stg2_reg[42]  ( .D(n461), .CP(clk), .CD(n1973), .Q(
        out1_stg2[42]), .QN(n1591) );
  CFD2XL \out1_stg2_reg[41]  ( .D(n463), .CP(clk), .CD(n1973), .Q(
        out1_stg2[41]), .QN(n1595) );
  CFD2XL \out1_stg2_reg[40]  ( .D(n465), .CP(clk), .CD(n1973), .Q(
        out1_stg2[40]), .QN(n1599) );
  CFD2XL \out1_stg2_reg[39]  ( .D(n467), .CP(clk), .CD(n1973), .Q(
        out1_stg2[39]), .QN(n1603) );
  CFD2XL \out1_stg2_reg[38]  ( .D(n469), .CP(clk), .CD(n1973), .Q(
        out1_stg2[38]), .QN(n1607) );
  CFD2XL \out1_stg2_reg[37]  ( .D(n471), .CP(clk), .CD(n1973), .Q(
        out1_stg2[37]), .QN(n1611) );
  CFD2XL \out1_stg2_reg[36]  ( .D(n473), .CP(clk), .CD(n1973), .Q(
        out1_stg2[36]), .QN(n1615) );
  CFD2XL \out1_stg2_reg[35]  ( .D(n475), .CP(clk), .CD(n1973), .Q(
        out1_stg2[35]), .QN(n1619) );
  CFD2XL \out1_stg2_reg[34]  ( .D(n477), .CP(clk), .CD(n1973), .Q(
        out1_stg2[34]), .QN(n1623) );
  CFD2XL \out1_stg2_reg[33]  ( .D(n479), .CP(clk), .CD(n1973), .Q(
        out1_stg2[33]), .QN(n1627) );
  CFD1QXL roundit_reg ( .D(n611), .CP(clk), .Q(roundit) );
  CFD1QXL cmd1_en_stg2_reg ( .D(n756), .CP(clk), .Q(cmd1_en_stg2) );
  CFD2QX1 \q0_reg[18]  ( .D(n676), .CP(clk), .CD(n1320), .Q(q0[18]) );
  CFD2QX1 \q0_reg[26]  ( .D(n1101), .CP(clk), .CD(n1319), .Q(q0[26]) );
  CFD2QX1 \q0_reg[12]  ( .D(n1100), .CP(clk), .CD(n1320), .Q(q0[12]) );
  CFD2QX1 \q0_reg[8]  ( .D(n1099), .CP(clk), .CD(n1320), .Q(q0[8]) );
  CFD2QX1 \h0_reg[0]  ( .D(n614), .CP(clk), .CD(n1323), .Q(h0[0]) );
  CFD2QX1 \q0_reg[22]  ( .D(n1109), .CP(clk), .CD(n1319), .Q(q0[22]) );
  CFD2QX1 \h0_reg[4]  ( .D(n626), .CP(clk), .CD(n1323), .Q(h0[4]) );
  CFD2QX1 \h0_reg[17]  ( .D(n815), .CP(clk), .CD(n1322), .Q(h0[17]) );
  CFD2QX1 \q0_reg[16]  ( .D(n674), .CP(clk), .CD(n1320), .Q(q0[16]) );
  CFD2QX2 \q0_reg[17]  ( .D(n1104), .CP(clk), .CD(n1320), .Q(q0[17]) );
  CFD2QX1 \q0_reg[7]  ( .D(n665), .CP(clk), .CD(n1320), .Q(q0[7]) );
  CFD2QX1 \q0_reg[10]  ( .D(n792), .CP(clk), .CD(n1320), .Q(q0[10]) );
  CFD2QX1 \q0_reg[1]  ( .D(n659), .CP(clk), .CD(n1307), .Q(q0[1]) );
  CNIVX1 U921 ( .A(n658), .Z(n790) );
  CNIVX1 U922 ( .A(n660), .Z(n791) );
  CNIVX1 U923 ( .A(n668), .Z(n792) );
  CDLY1XL U924 ( .A(q0[23]), .Z(n793) );
  CDLY1XL U925 ( .A(n804), .Z(n794) );
  CDLY1XL U926 ( .A(q0[3]), .Z(n795) );
  CDLY1XL U927 ( .A(q0[9]), .Z(n796) );
  CNIVX3 U928 ( .A(n801), .Z(n1212) );
  CIVXL U929 ( .A(cmd1_en_stg2), .Z(n1268) );
  CIVXL U930 ( .A(cmd1_en_stg2), .Z(n1266) );
  CIVXL U931 ( .A(cmd1_en_stg2), .Z(n1265) );
  CIVX2 U932 ( .A(n797), .Z(n1378) );
  CIVDX1 U933 ( .A(cmd2_en_stg2), .Z0(n797), .Z1(n798) );
  CIVX2 U934 ( .A(n1436), .Z(n1300) );
  CAN3X1 U935 ( .A(cmd0[1]), .B(n1976), .C(push0), .Z(n799) );
  CIVXL U936 ( .A(n1267), .Z(n1289) );
  CIVXL U937 ( .A(n1267), .Z(n1288) );
  CAN4X1 U938 ( .A(n1917), .B(push0_stg2), .C(n1916), .D(n1915), .Z(n800) );
  CAN3XL U939 ( .A(cmd1_en_stg2_d), .B(n1379), .C(n1767), .Z(n801) );
  CNIVX1 U940 ( .A(n1972), .Z(n802) );
  CDLY1XL U941 ( .A(q0[25]), .Z(n803) );
  CNIVX4 U942 ( .A(q0[18]), .Z(n804) );
  CIVXL U943 ( .A(q0[17]), .Z(n805) );
  CIVX2 U944 ( .A(n805), .Z(n806) );
  CDLY1XL U945 ( .A(q0[21]), .Z(n807) );
  CNIVX1 U946 ( .A(_pushout_d), .Z(n808) );
  CNIVX1 U947 ( .A(n681), .Z(n809) );
  CNIVX1 U948 ( .A(n667), .Z(n810) );
  CNIVX1 U949 ( .A(n649), .Z(n811) );
  CNIVX1 U950 ( .A(n642), .Z(n812) );
  CNIVX1 U951 ( .A(n644), .Z(n813) );
  CNIVX1 U952 ( .A(n635), .Z(n814) );
  CNIVX1 U953 ( .A(n643), .Z(n815) );
  CNIVX1 U954 ( .A(n634), .Z(n816) );
  CMX2XL U955 ( .A0(h0[8]), .A1(h[8]), .S(n1384), .Z(n634) );
  CNIVX1 U956 ( .A(n639), .Z(n817) );
  CNIVX1 U957 ( .A(n640), .Z(n818) );
  CNIVX1 U958 ( .A(n655), .Z(n819) );
  CNIVX1 U959 ( .A(n648), .Z(n820) );
  CNIVX1 U960 ( .A(n646), .Z(n821) );
  CNIVX1 U961 ( .A(n647), .Z(n822) );
  CNIVX1 U962 ( .A(n637), .Z(n823) );
  CNIVX1 U963 ( .A(n653), .Z(n824) );
  CNIVX1 U964 ( .A(n651), .Z(n825) );
  CNIVX1 U965 ( .A(n645), .Z(n826) );
  CNIVX1 U966 ( .A(n656), .Z(n827) );
  CNIVX1 U967 ( .A(n610), .Z(n828) );
  CIVX3 U968 ( .A(out2_stg2[30]), .Z(n1440) );
  CIVX3 U969 ( .A(out2_stg2[28]), .Z(n1444) );
  CIVX3 U970 ( .A(out2_stg2[26]), .Z(n1448) );
  CIVX3 U971 ( .A(out2_stg2[24]), .Z(n1452) );
  CIVX3 U972 ( .A(out2_stg2[22]), .Z(n1456) );
  CIVX3 U973 ( .A(out2_stg2[20]), .Z(n1460) );
  CIVX3 U974 ( .A(out2_stg2[18]), .Z(n1464) );
  CIVX3 U975 ( .A(out2_stg2[16]), .Z(n1468) );
  CIVX3 U976 ( .A(out2_stg2[14]), .Z(n1472) );
  CIVX3 U977 ( .A(out2_stg2[12]), .Z(n1476) );
  CIVX3 U978 ( .A(out2_stg2[10]), .Z(n1480) );
  CIVX3 U979 ( .A(out2_stg2[8]), .Z(n1484) );
  CIVX3 U980 ( .A(out2_stg2[6]), .Z(n1488) );
  CIVX3 U981 ( .A(out2_stg2[4]), .Z(n1492) );
  CIVX3 U982 ( .A(out2_stg2[2]), .Z(n1496) );
  CIVX3 U983 ( .A(out2_stg2[15]), .Z(n1470) );
  CIVX3 U984 ( .A(out2_stg2[13]), .Z(n1474) );
  CIVX3 U985 ( .A(out2_stg2[11]), .Z(n1478) );
  CIVX3 U986 ( .A(out2_stg2[9]), .Z(n1482) );
  CIVX3 U987 ( .A(out2_stg2[3]), .Z(n1494) );
  CIVX3 U988 ( .A(out2_stg2[1]), .Z(n1498) );
  CMX2X2 U989 ( .A0(out0_stg2[62]), .A1(out0_stg1[62]), .S(n1232), .Z(n692) );
  CMX2X2 U990 ( .A0(out0_stg2[61]), .A1(out0_stg1[61]), .S(n1233), .Z(n693) );
  CMX2X2 U991 ( .A0(out0_stg2[60]), .A1(out0_stg1[60]), .S(n1234), .Z(n694) );
  CMX2X2 U992 ( .A0(out0_stg2[59]), .A1(out0_stg1[59]), .S(n1235), .Z(n695) );
  CMX2X2 U993 ( .A0(out0_stg2[58]), .A1(out0_stg1[58]), .S(n1236), .Z(n696) );
  CMX2X2 U994 ( .A0(out0_stg2[57]), .A1(out0_stg1[57]), .S(n1237), .Z(n697) );
  CMX2X2 U995 ( .A0(out0_stg2[56]), .A1(out0_stg1[56]), .S(n1238), .Z(n698) );
  CMX2X2 U996 ( .A0(out0_stg2[55]), .A1(out0_stg1[55]), .S(n1239), .Z(n699) );
  CMX2X2 U997 ( .A0(out0_stg2[54]), .A1(out0_stg1[54]), .S(n1240), .Z(n700) );
  CMX2X2 U998 ( .A0(out0_stg2[53]), .A1(out0_stg1[53]), .S(n1241), .Z(n701) );
  CMX2X2 U999 ( .A0(out0_stg2[52]), .A1(out0_stg1[52]), .S(n1242), .Z(n702) );
  CMX2X2 U1000 ( .A0(out0_stg2[51]), .A1(out0_stg1[51]), .S(n1243), .Z(n703)
         );
  CMX2X2 U1001 ( .A0(out0_stg2[50]), .A1(out0_stg1[50]), .S(n1244), .Z(n704)
         );
  CMX2X2 U1002 ( .A0(out0_stg2[49]), .A1(out0_stg1[49]), .S(n1245), .Z(n705)
         );
  CMX2X2 U1003 ( .A0(out0_stg2[48]), .A1(out0_stg1[48]), .S(n1246), .Z(n706)
         );
  CMX2X2 U1004 ( .A0(out0_stg2[47]), .A1(out0_stg1[47]), .S(n1247), .Z(n707)
         );
  CMX2X2 U1005 ( .A0(out0_stg2[46]), .A1(out0_stg1[46]), .S(n1248), .Z(n708)
         );
  CMX2X2 U1006 ( .A0(out0_stg2[45]), .A1(out0_stg1[45]), .S(n1249), .Z(n709)
         );
  CMX2X2 U1007 ( .A0(out0_stg2[44]), .A1(out0_stg1[44]), .S(n1250), .Z(n710)
         );
  CMX2X2 U1008 ( .A0(out0_stg2[43]), .A1(out0_stg1[43]), .S(n1251), .Z(n711)
         );
  CMX2X2 U1009 ( .A0(out0_stg2[42]), .A1(out0_stg1[42]), .S(n1252), .Z(n712)
         );
  CMX2X2 U1010 ( .A0(out0_stg2[41]), .A1(out0_stg1[41]), .S(n1253), .Z(n713)
         );
  CMX2X2 U1011 ( .A0(out0_stg2[40]), .A1(out0_stg1[40]), .S(n1254), .Z(n714)
         );
  CMX2X2 U1012 ( .A0(out0_stg2[39]), .A1(out0_stg1[39]), .S(n1255), .Z(n715)
         );
  CMX2X2 U1013 ( .A0(out0_stg2[38]), .A1(out0_stg1[38]), .S(n1256), .Z(n716)
         );
  CMX2X2 U1014 ( .A0(out0_stg2[37]), .A1(out0_stg1[37]), .S(n1257), .Z(n717)
         );
  CMX2X2 U1015 ( .A0(out0_stg2[36]), .A1(out0_stg1[36]), .S(n1258), .Z(n718)
         );
  CMX2X2 U1016 ( .A0(out0_stg2[35]), .A1(out0_stg1[35]), .S(n1259), .Z(n719)
         );
  CMX2X2 U1017 ( .A0(out0_stg2[34]), .A1(out0_stg1[34]), .S(n1257), .Z(n720)
         );
  CMX2X2 U1018 ( .A0(out0_stg2[33]), .A1(out0_stg1[33]), .S(n1258), .Z(n721)
         );
  CMX2X2 U1019 ( .A0(out0_stg2[32]), .A1(out0_stg1[32]), .S(n1259), .Z(n722)
         );
  CMX2X2 U1020 ( .A0(out0_stg2[31]), .A1(out0_stg1[31]), .S(n1262), .Z(n723)
         );
  CMX2X2 U1021 ( .A0(out0_stg2[30]), .A1(out0_stg1[30]), .S(n1254), .Z(n724)
         );
  CMX2X2 U1022 ( .A0(out0_stg2[29]), .A1(out0_stg1[29]), .S(n1256), .Z(n725)
         );
  CMX2X2 U1023 ( .A0(out0_stg2[28]), .A1(out0_stg1[28]), .S(n1261), .Z(n726)
         );
  CMX2X2 U1024 ( .A0(out0_stg2[27]), .A1(out0_stg1[27]), .S(n1260), .Z(n727)
         );
  CMX2X2 U1025 ( .A0(out0_stg2[26]), .A1(out0_stg1[26]), .S(n1260), .Z(n728)
         );
  CMX2X2 U1026 ( .A0(out0_stg2[25]), .A1(out0_stg1[25]), .S(n1261), .Z(n729)
         );
  CMX2X2 U1027 ( .A0(out0_stg2[24]), .A1(out0_stg1[24]), .S(n1262), .Z(n730)
         );
  CMX2X2 U1028 ( .A0(out0_stg2[23]), .A1(out0_stg1[23]), .S(n1233), .Z(n731)
         );
  CMX2X2 U1029 ( .A0(out0_stg2[22]), .A1(out0_stg1[22]), .S(n1231), .Z(n732)
         );
  CMX2X2 U1030 ( .A0(out0_stg2[21]), .A1(out0_stg1[21]), .S(n1232), .Z(n733)
         );
  CMX2X2 U1031 ( .A0(out0_stg2[20]), .A1(out0_stg1[20]), .S(n1233), .Z(n734)
         );
  CMX2X2 U1032 ( .A0(out0_stg2[19]), .A1(out0_stg1[19]), .S(n1234), .Z(n735)
         );
  CMX2X2 U1033 ( .A0(out0_stg2[18]), .A1(out0_stg1[18]), .S(n1235), .Z(n736)
         );
  CMX2X2 U1034 ( .A0(out0_stg2[17]), .A1(out0_stg1[17]), .S(n1236), .Z(n737)
         );
  CMX2X2 U1035 ( .A0(out0_stg2[16]), .A1(out0_stg1[16]), .S(n1237), .Z(n738)
         );
  CMX2X2 U1036 ( .A0(out0_stg2[15]), .A1(out0_stg1[15]), .S(n1238), .Z(n739)
         );
  CMX2X2 U1037 ( .A0(out0_stg2[14]), .A1(out0_stg1[14]), .S(n1239), .Z(n740)
         );
  CMX2X2 U1038 ( .A0(out0_stg2[13]), .A1(out0_stg1[13]), .S(n1240), .Z(n741)
         );
  CMX2X2 U1039 ( .A0(out0_stg2[12]), .A1(out0_stg1[12]), .S(n1241), .Z(n742)
         );
  CMX2X2 U1040 ( .A0(out0_stg2[11]), .A1(out0_stg1[11]), .S(n1242), .Z(n743)
         );
  CMX2X2 U1041 ( .A0(out0_stg2[10]), .A1(out0_stg1[10]), .S(n1243), .Z(n744)
         );
  CMX2X2 U1042 ( .A0(out0_stg2[9]), .A1(out0_stg1[9]), .S(n1244), .Z(n745) );
  CMX2X2 U1043 ( .A0(out0_stg2[8]), .A1(out0_stg1[8]), .S(n1245), .Z(n746) );
  CMX2X2 U1044 ( .A0(out0_stg2[7]), .A1(out0_stg1[7]), .S(n1246), .Z(n747) );
  CMX2X2 U1045 ( .A0(out0_stg2[6]), .A1(out0_stg1[6]), .S(n1247), .Z(n748) );
  CMX2X2 U1046 ( .A0(out0_stg2[5]), .A1(out0_stg1[5]), .S(n1248), .Z(n749) );
  CMX2X2 U1047 ( .A0(out0_stg2[4]), .A1(out0_stg1[4]), .S(n1249), .Z(n750) );
  CMX2X2 U1048 ( .A0(out0_stg2[3]), .A1(out0_stg1[3]), .S(n1250), .Z(n751) );
  CMX2X2 U1049 ( .A0(out0_stg2[2]), .A1(out0_stg1[2]), .S(n1251), .Z(n752) );
  CMX2X2 U1050 ( .A0(out0_stg2[1]), .A1(out0_stg1[1]), .S(n1252), .Z(n753) );
  CMX2X2 U1051 ( .A0(out0_stg2[0]), .A1(out0_stg1[0]), .S(n1253), .Z(n754) );
  CIVDX1 U1052 ( .A(out1_stg0[0]), .Z1(n830) );
  CNIVX1 U1053 ( .A(n830), .Z(n829) );
  CIVDX1 U1054 ( .A(out1_stg0[1]), .Z1(n832) );
  CNIVX1 U1055 ( .A(n832), .Z(n831) );
  CIVDX1 U1056 ( .A(out1_stg0[2]), .Z1(n834) );
  CNIVX1 U1057 ( .A(n834), .Z(n833) );
  CIVDX1 U1058 ( .A(out1_stg0[3]), .Z1(n836) );
  CNIVX1 U1059 ( .A(n836), .Z(n835) );
  CIVDX1 U1060 ( .A(out1_stg0[4]), .Z1(n838) );
  CNIVX1 U1061 ( .A(n838), .Z(n837) );
  CIVDX1 U1062 ( .A(out1_stg0[5]), .Z1(n840) );
  CNIVX1 U1063 ( .A(n840), .Z(n839) );
  CIVDX1 U1064 ( .A(out1_stg0[6]), .Z1(n842) );
  CNIVX1 U1065 ( .A(n842), .Z(n841) );
  CIVDX1 U1066 ( .A(out1_stg0[7]), .Z1(n844) );
  CNIVX1 U1067 ( .A(n844), .Z(n843) );
  CIVDX1 U1068 ( .A(out1_stg0[8]), .Z1(n846) );
  CNIVX1 U1069 ( .A(n846), .Z(n845) );
  CIVDX1 U1070 ( .A(out1_stg0[9]), .Z1(n848) );
  CNIVX1 U1071 ( .A(n848), .Z(n847) );
  CIVDX1 U1072 ( .A(out1_stg0[10]), .Z1(n850) );
  CNIVX1 U1073 ( .A(n850), .Z(n849) );
  CIVDX1 U1074 ( .A(out1_stg0[11]), .Z1(n852) );
  CNIVX1 U1075 ( .A(n852), .Z(n851) );
  CIVDX1 U1076 ( .A(out1_stg0[12]), .Z1(n854) );
  CNIVX1 U1077 ( .A(n854), .Z(n853) );
  CIVDX1 U1078 ( .A(out1_stg0[13]), .Z1(n856) );
  CNIVX1 U1079 ( .A(n856), .Z(n855) );
  CIVDX1 U1080 ( .A(out1_stg0[14]), .Z1(n858) );
  CNIVX1 U1081 ( .A(n858), .Z(n857) );
  CIVDX1 U1082 ( .A(out1_stg0[15]), .Z1(n860) );
  CNIVX1 U1083 ( .A(n860), .Z(n859) );
  CIVDX1 U1084 ( .A(out1_stg0[16]), .Z1(n862) );
  CNIVX1 U1085 ( .A(n862), .Z(n861) );
  CIVDX1 U1086 ( .A(out1_stg0[17]), .Z1(n864) );
  CNIVX1 U1087 ( .A(n864), .Z(n863) );
  CIVDX1 U1088 ( .A(out1_stg0[18]), .Z1(n866) );
  CNIVX1 U1089 ( .A(n866), .Z(n865) );
  CIVDX1 U1090 ( .A(out1_stg0[19]), .Z1(n868) );
  CNIVX1 U1091 ( .A(n868), .Z(n867) );
  CIVDX1 U1092 ( .A(out1_stg0[20]), .Z1(n870) );
  CNIVX1 U1093 ( .A(n870), .Z(n869) );
  CIVDX1 U1094 ( .A(out1_stg0[21]), .Z1(n872) );
  CNIVX1 U1095 ( .A(n872), .Z(n871) );
  CIVDX1 U1096 ( .A(out1_stg0[22]), .Z1(n874) );
  CNIVX1 U1097 ( .A(n874), .Z(n873) );
  CIVDX1 U1098 ( .A(out1_stg0[23]), .Z1(n876) );
  CNIVX1 U1099 ( .A(n876), .Z(n875) );
  CIVDX1 U1100 ( .A(out1_stg0[24]), .Z1(n878) );
  CNIVX1 U1101 ( .A(n878), .Z(n877) );
  CIVDX1 U1102 ( .A(out1_stg0[25]), .Z1(n880) );
  CNIVX1 U1103 ( .A(n880), .Z(n879) );
  CIVDX1 U1104 ( .A(out1_stg0[26]), .Z1(n882) );
  CNIVX1 U1105 ( .A(n882), .Z(n881) );
  CIVDX1 U1106 ( .A(out1_stg0[27]), .Z1(n884) );
  CNIVX1 U1107 ( .A(n884), .Z(n883) );
  CIVDX1 U1108 ( .A(out1_stg0[28]), .Z1(n886) );
  CNIVX1 U1109 ( .A(n886), .Z(n885) );
  CIVDX1 U1110 ( .A(out1_stg0[29]), .Z1(n888) );
  CNIVX1 U1111 ( .A(n888), .Z(n887) );
  CIVDX1 U1112 ( .A(out1_stg0[30]), .Z1(n890) );
  CNIVX1 U1113 ( .A(n890), .Z(n889) );
  CIVDX1 U1114 ( .A(out1_stg0[31]), .Z1(n892) );
  CNIVX1 U1115 ( .A(n892), .Z(n891) );
  CIVDX1 U1116 ( .A(out1_stg0[32]), .Z1(n894) );
  CNIVX1 U1117 ( .A(n894), .Z(n893) );
  CIVDX1 U1118 ( .A(out1_stg0[33]), .Z1(n896) );
  CNIVX1 U1119 ( .A(n896), .Z(n895) );
  CIVDX1 U1120 ( .A(out1_stg0[34]), .Z1(n898) );
  CNIVX1 U1121 ( .A(n898), .Z(n897) );
  CIVDX1 U1122 ( .A(out1_stg0[35]), .Z1(n900) );
  CNIVX1 U1123 ( .A(n900), .Z(n899) );
  CIVDX1 U1124 ( .A(out1_stg0[36]), .Z1(n902) );
  CNIVX1 U1125 ( .A(n902), .Z(n901) );
  CIVDX1 U1126 ( .A(out1_stg0[37]), .Z1(n904) );
  CNIVX1 U1127 ( .A(n904), .Z(n903) );
  CIVDX1 U1128 ( .A(out1_stg0[38]), .Z1(n906) );
  CNIVX1 U1129 ( .A(n906), .Z(n905) );
  CIVDX1 U1130 ( .A(out1_stg0[39]), .Z1(n908) );
  CNIVX1 U1131 ( .A(n908), .Z(n907) );
  CIVDX1 U1132 ( .A(out1_stg0[40]), .Z1(n910) );
  CNIVX1 U1133 ( .A(n910), .Z(n909) );
  CIVDX1 U1134 ( .A(out1_stg0[41]), .Z1(n912) );
  CNIVX1 U1135 ( .A(n912), .Z(n911) );
  CIVDX1 U1136 ( .A(out1_stg0[42]), .Z1(n914) );
  CNIVX1 U1137 ( .A(n914), .Z(n913) );
  CIVDX1 U1138 ( .A(out1_stg0[43]), .Z1(n916) );
  CNIVX1 U1139 ( .A(n916), .Z(n915) );
  CIVDX1 U1140 ( .A(out1_stg0[44]), .Z1(n918) );
  CNIVX1 U1141 ( .A(n918), .Z(n917) );
  CIVDX1 U1142 ( .A(out1_stg0[45]), .Z1(n920) );
  CNIVX1 U1143 ( .A(n920), .Z(n919) );
  CIVDX1 U1144 ( .A(out1_stg0[46]), .Z1(n922) );
  CNIVX1 U1145 ( .A(n922), .Z(n921) );
  CIVDX1 U1146 ( .A(out1_stg0[47]), .Z1(n924) );
  CNIVX1 U1147 ( .A(n924), .Z(n923) );
  CIVDX1 U1148 ( .A(out1_stg0[48]), .Z1(n926) );
  CNIVX1 U1149 ( .A(n926), .Z(n925) );
  CIVDX1 U1150 ( .A(out1_stg0[49]), .Z1(n928) );
  CNIVX1 U1151 ( .A(n928), .Z(n927) );
  CIVDX1 U1152 ( .A(out1_stg0[50]), .Z1(n930) );
  CNIVX1 U1153 ( .A(n930), .Z(n929) );
  CIVDX1 U1154 ( .A(out1_stg0[51]), .Z1(n932) );
  CNIVX1 U1155 ( .A(n932), .Z(n931) );
  CIVDX1 U1156 ( .A(out1_stg0[52]), .Z1(n934) );
  CNIVX1 U1157 ( .A(n934), .Z(n933) );
  CIVDX1 U1158 ( .A(out1_stg0[53]), .Z1(n936) );
  CNIVX1 U1159 ( .A(n936), .Z(n935) );
  CIVDX1 U1160 ( .A(out1_stg0[55]), .Z1(n938) );
  CNIVX1 U1161 ( .A(n938), .Z(n937) );
  CIVDX1 U1162 ( .A(out1_stg0[56]), .Z1(n940) );
  CNIVX1 U1163 ( .A(n940), .Z(n939) );
  CIVDX1 U1164 ( .A(out1_stg0[57]), .Z1(n942) );
  CNIVX1 U1165 ( .A(n942), .Z(n941) );
  CIVDX1 U1166 ( .A(out1_stg0[58]), .Z1(n944) );
  CNIVX1 U1167 ( .A(n944), .Z(n943) );
  CIVDX1 U1168 ( .A(out1_stg0[59]), .Z1(n946) );
  CNIVX1 U1169 ( .A(n946), .Z(n945) );
  CIVDX1 U1170 ( .A(cmd0_stg1[1]), .Z1(n948) );
  CNIVX1 U1171 ( .A(n948), .Z(n947) );
  CIVDX1 U1172 ( .A(cmd0_stg1[0]), .Z1(n950) );
  CNIVX1 U1173 ( .A(n950), .Z(n949) );
  CMX2X2 U1174 ( .A0(out0_stg2[63]), .A1(out0_stg1[63]), .S(n1231), .Z(n691)
         );
  CIVDX1 U1175 ( .A(out1_stg0[54]), .Z1(n952) );
  CNIVX1 U1176 ( .A(n952), .Z(n951) );
  CIVDX1 U1177 ( .A(out1_stg0[60]), .Z1(n954) );
  CNIVX1 U1178 ( .A(n954), .Z(n953) );
  CIVDX1 U1179 ( .A(out1_stg0[61]), .Z1(n956) );
  CNIVX1 U1180 ( .A(n956), .Z(n955) );
  CIVDX1 U1181 ( .A(out1_stg0[62]), .Z1(n958) );
  CNIVX1 U1182 ( .A(n958), .Z(n957) );
  CIVDX1 U1183 ( .A(out1_stg0[63]), .Z1(n960) );
  CNIVX1 U1184 ( .A(n960), .Z(n959) );
  CNIVX1 U1185 ( .A(n613), .Z(n961) );
  CNIVX1 U1186 ( .A(n616), .Z(n962) );
  CNIVX1 U1187 ( .A(n619), .Z(n963) );
  CNIVX1 U1188 ( .A(n622), .Z(n964) );
  CNIVX1 U1189 ( .A(h0[3]), .Z(n965) );
  CNIVX1 U1190 ( .A(n625), .Z(n966) );
  CNIVX1 U1191 ( .A(n628), .Z(n967) );
  CNIVX1 U1192 ( .A(n631), .Z(n968) );
  CNIVX1 U1193 ( .A(h0[6]), .Z(n969) );
  CMX2X2 U1194 ( .A0(z[0]), .A1(acc[0]), .S(n800), .Z(n758) );
  CMX2X2 U1195 ( .A0(z[1]), .A1(acc[1]), .S(n800), .Z(n759) );
  CMXI2X2 U1196 ( .A0(n1919), .A1(n1918), .S(n800), .Z(n760) );
  CMX2X2 U1197 ( .A0(z[3]), .A1(acc[3]), .S(n800), .Z(n761) );
  CMXI2X2 U1198 ( .A0(n1921), .A1(n1920), .S(n800), .Z(n762) );
  CMXI2X2 U1199 ( .A0(n1923), .A1(n1922), .S(n800), .Z(n763) );
  CMXI2X2 U1200 ( .A0(n1925), .A1(n1924), .S(n800), .Z(n764) );
  CMXI2X2 U1201 ( .A0(n1927), .A1(n1926), .S(n800), .Z(n765) );
  CMXI2X2 U1202 ( .A0(n1929), .A1(n1928), .S(n800), .Z(n766) );
  CMX2X2 U1203 ( .A0(z[9]), .A1(acc[9]), .S(n800), .Z(n767) );
  CMXI2X2 U1204 ( .A0(n1931), .A1(n1930), .S(n800), .Z(n768) );
  CMX2X2 U1205 ( .A0(z[11]), .A1(acc[11]), .S(n800), .Z(n769) );
  CMXI2X2 U1206 ( .A0(n1933), .A1(n1932), .S(n800), .Z(n770) );
  CMXI2X2 U1207 ( .A0(n1935), .A1(n1934), .S(n800), .Z(n771) );
  CMXI2X2 U1208 ( .A0(n1937), .A1(n1936), .S(n800), .Z(n772) );
  CMXI2X2 U1209 ( .A0(n1939), .A1(n1938), .S(n800), .Z(n773) );
  CMXI2X2 U1210 ( .A0(n1941), .A1(n1940), .S(n800), .Z(n774) );
  CMXI2X2 U1211 ( .A0(n1943), .A1(n1942), .S(n800), .Z(n775) );
  CMXI2X2 U1212 ( .A0(n1945), .A1(n1944), .S(n800), .Z(n776) );
  CMXI2X2 U1213 ( .A0(n1947), .A1(n1946), .S(n800), .Z(n777) );
  CMXI2X2 U1214 ( .A0(n1949), .A1(n1948), .S(n800), .Z(n778) );
  CMXI2X2 U1215 ( .A0(n1951), .A1(n1950), .S(n800), .Z(n779) );
  CMXI2X2 U1216 ( .A0(n1953), .A1(n1952), .S(n800), .Z(n780) );
  CMXI2X2 U1217 ( .A0(n1955), .A1(n1954), .S(n800), .Z(n781) );
  CMXI2X2 U1218 ( .A0(n1957), .A1(n1956), .S(n800), .Z(n782) );
  CMXI2X2 U1219 ( .A0(n1959), .A1(n1958), .S(n800), .Z(n783) );
  CMXI2X2 U1220 ( .A0(n1961), .A1(n1960), .S(n800), .Z(n784) );
  CMXI2X2 U1221 ( .A0(n1963), .A1(n1962), .S(n800), .Z(n785) );
  CMXI2X2 U1222 ( .A0(n1965), .A1(n1964), .S(n800), .Z(n786) );
  CMXI2X2 U1223 ( .A0(n1967), .A1(n1966), .S(n800), .Z(n787) );
  CMXI2X2 U1224 ( .A0(n1969), .A1(n1968), .S(n800), .Z(n788) );
  CMXI2X2 U1225 ( .A0(n1971), .A1(n1970), .S(n800), .Z(n789) );
  CIVDX1 U1226 ( .A(out0_stg0[0]), .Z1(n971) );
  CNIVX1 U1227 ( .A(n971), .Z(n970) );
  CIVDX1 U1228 ( .A(out0_stg0[1]), .Z1(n973) );
  CNIVX1 U1229 ( .A(n973), .Z(n972) );
  CIVDX1 U1230 ( .A(out0_stg0[2]), .Z1(n975) );
  CNIVX1 U1231 ( .A(n975), .Z(n974) );
  CIVDX1 U1232 ( .A(out0_stg0[3]), .Z1(n977) );
  CNIVX1 U1233 ( .A(n977), .Z(n976) );
  CIVDX1 U1234 ( .A(out0_stg0[4]), .Z1(n979) );
  CNIVX1 U1235 ( .A(n979), .Z(n978) );
  CIVDX1 U1236 ( .A(out0_stg0[5]), .Z1(n981) );
  CNIVX1 U1237 ( .A(n981), .Z(n980) );
  CIVDX1 U1238 ( .A(out0_stg0[6]), .Z1(n983) );
  CNIVX1 U1239 ( .A(n983), .Z(n982) );
  CIVDX1 U1240 ( .A(out0_stg0[7]), .Z1(n985) );
  CNIVX1 U1241 ( .A(n985), .Z(n984) );
  CIVDX1 U1242 ( .A(out0_stg0[8]), .Z1(n987) );
  CNIVX1 U1243 ( .A(n987), .Z(n986) );
  CIVDX1 U1244 ( .A(out0_stg0[9]), .Z1(n989) );
  CNIVX1 U1245 ( .A(n989), .Z(n988) );
  CIVDX1 U1246 ( .A(out0_stg0[10]), .Z1(n991) );
  CNIVX1 U1247 ( .A(n991), .Z(n990) );
  CIVDX1 U1248 ( .A(out0_stg0[11]), .Z1(n993) );
  CNIVX1 U1249 ( .A(n993), .Z(n992) );
  CIVDX1 U1250 ( .A(out0_stg0[12]), .Z1(n995) );
  CNIVX1 U1251 ( .A(n995), .Z(n994) );
  CIVDX1 U1252 ( .A(out0_stg0[13]), .Z1(n997) );
  CNIVX1 U1253 ( .A(n997), .Z(n996) );
  CIVDX1 U1254 ( .A(out0_stg0[14]), .Z1(n999) );
  CNIVX1 U1255 ( .A(n999), .Z(n998) );
  CIVDX1 U1256 ( .A(out0_stg0[15]), .Z1(n1001) );
  CNIVX1 U1257 ( .A(n1001), .Z(n1000) );
  CIVDX1 U1258 ( .A(out0_stg0[16]), .Z1(n1003) );
  CNIVX1 U1259 ( .A(n1003), .Z(n1002) );
  CIVDX1 U1260 ( .A(out0_stg0[17]), .Z1(n1005) );
  CNIVX1 U1261 ( .A(n1005), .Z(n1004) );
  CIVDX1 U1262 ( .A(out0_stg0[18]), .Z1(n1007) );
  CNIVX1 U1263 ( .A(n1007), .Z(n1006) );
  CIVDX1 U1264 ( .A(out0_stg0[19]), .Z1(n1009) );
  CNIVX1 U1265 ( .A(n1009), .Z(n1008) );
  CIVDX1 U1266 ( .A(out0_stg0[20]), .Z1(n1011) );
  CNIVX1 U1267 ( .A(n1011), .Z(n1010) );
  CIVDX1 U1268 ( .A(out0_stg0[21]), .Z1(n1013) );
  CNIVX1 U1269 ( .A(n1013), .Z(n1012) );
  CIVDX1 U1270 ( .A(out0_stg0[22]), .Z1(n1015) );
  CNIVX1 U1271 ( .A(n1015), .Z(n1014) );
  CIVDX1 U1272 ( .A(out0_stg0[23]), .Z1(n1017) );
  CNIVX1 U1273 ( .A(n1017), .Z(n1016) );
  CIVDX1 U1274 ( .A(out0_stg0[24]), .Z1(n1019) );
  CNIVX1 U1275 ( .A(n1019), .Z(n1018) );
  CIVDX1 U1276 ( .A(out0_stg0[25]), .Z1(n1021) );
  CNIVX1 U1277 ( .A(n1021), .Z(n1020) );
  CIVDX1 U1278 ( .A(out0_stg0[26]), .Z1(n1023) );
  CNIVX1 U1279 ( .A(n1023), .Z(n1022) );
  CIVDX1 U1280 ( .A(out0_stg0[27]), .Z1(n1025) );
  CNIVX1 U1281 ( .A(n1025), .Z(n1024) );
  CIVDX1 U1282 ( .A(out0_stg0[28]), .Z1(n1027) );
  CNIVX1 U1283 ( .A(n1027), .Z(n1026) );
  CIVDX1 U1284 ( .A(out0_stg0[29]), .Z1(n1029) );
  CNIVX1 U1285 ( .A(n1029), .Z(n1028) );
  CIVDX1 U1286 ( .A(out0_stg0[30]), .Z1(n1031) );
  CNIVX1 U1287 ( .A(n1031), .Z(n1030) );
  CIVDX1 U1288 ( .A(out0_stg0[31]), .Z1(n1033) );
  CNIVX1 U1289 ( .A(n1033), .Z(n1032) );
  CIVDX1 U1290 ( .A(out0_stg0[32]), .Z1(n1035) );
  CNIVX1 U1291 ( .A(n1035), .Z(n1034) );
  CIVDX1 U1292 ( .A(out0_stg0[33]), .Z1(n1037) );
  CNIVX1 U1293 ( .A(n1037), .Z(n1036) );
  CIVDX1 U1294 ( .A(out0_stg0[34]), .Z1(n1039) );
  CNIVX1 U1295 ( .A(n1039), .Z(n1038) );
  CIVDX1 U1296 ( .A(out0_stg0[35]), .Z1(n1041) );
  CNIVX1 U1297 ( .A(n1041), .Z(n1040) );
  CIVDX1 U1298 ( .A(out0_stg0[36]), .Z1(n1043) );
  CNIVX1 U1299 ( .A(n1043), .Z(n1042) );
  CIVDX1 U1300 ( .A(out0_stg0[37]), .Z1(n1045) );
  CNIVX1 U1301 ( .A(n1045), .Z(n1044) );
  CIVDX1 U1302 ( .A(out0_stg0[38]), .Z1(n1047) );
  CNIVX1 U1303 ( .A(n1047), .Z(n1046) );
  CIVDX1 U1304 ( .A(out0_stg0[39]), .Z1(n1049) );
  CNIVX1 U1305 ( .A(n1049), .Z(n1048) );
  CIVDX1 U1306 ( .A(out0_stg0[40]), .Z1(n1051) );
  CNIVX1 U1307 ( .A(n1051), .Z(n1050) );
  CIVDX1 U1308 ( .A(out0_stg0[41]), .Z1(n1053) );
  CNIVX1 U1309 ( .A(n1053), .Z(n1052) );
  CIVDX1 U1310 ( .A(out0_stg0[42]), .Z1(n1055) );
  CNIVX1 U1311 ( .A(n1055), .Z(n1054) );
  CIVDX1 U1312 ( .A(out0_stg0[43]), .Z1(n1057) );
  CNIVX1 U1313 ( .A(n1057), .Z(n1056) );
  CIVDX1 U1314 ( .A(out0_stg0[44]), .Z1(n1059) );
  CNIVX1 U1315 ( .A(n1059), .Z(n1058) );
  CIVDX1 U1316 ( .A(out0_stg0[45]), .Z1(n1061) );
  CNIVX1 U1317 ( .A(n1061), .Z(n1060) );
  CIVDX1 U1318 ( .A(out0_stg0[46]), .Z1(n1063) );
  CNIVX1 U1319 ( .A(n1063), .Z(n1062) );
  CIVDX1 U1320 ( .A(out0_stg0[47]), .Z1(n1065) );
  CNIVX1 U1321 ( .A(n1065), .Z(n1064) );
  CIVDX1 U1322 ( .A(out0_stg0[48]), .Z1(n1067) );
  CNIVX1 U1323 ( .A(n1067), .Z(n1066) );
  CIVDX1 U1324 ( .A(out0_stg0[49]), .Z1(n1069) );
  CNIVX1 U1325 ( .A(n1069), .Z(n1068) );
  CIVDX1 U1326 ( .A(out0_stg0[50]), .Z1(n1071) );
  CNIVX1 U1327 ( .A(n1071), .Z(n1070) );
  CIVDX1 U1328 ( .A(out0_stg0[51]), .Z1(n1073) );
  CNIVX1 U1329 ( .A(n1073), .Z(n1072) );
  CIVDX1 U1330 ( .A(out0_stg0[52]), .Z1(n1075) );
  CNIVX1 U1331 ( .A(n1075), .Z(n1074) );
  CIVDX1 U1332 ( .A(out0_stg0[53]), .Z1(n1077) );
  CNIVX1 U1333 ( .A(n1077), .Z(n1076) );
  CIVDX1 U1334 ( .A(out0_stg0[54]), .Z1(n1079) );
  CNIVX1 U1335 ( .A(n1079), .Z(n1078) );
  CIVDX1 U1336 ( .A(out0_stg0[55]), .Z1(n1081) );
  CNIVX1 U1337 ( .A(n1081), .Z(n1080) );
  CIVDX1 U1338 ( .A(out0_stg0[56]), .Z1(n1083) );
  CNIVX1 U1339 ( .A(n1083), .Z(n1082) );
  CIVDX1 U1340 ( .A(out0_stg0[57]), .Z1(n1085) );
  CNIVX1 U1341 ( .A(n1085), .Z(n1084) );
  CIVDX1 U1342 ( .A(out0_stg0[58]), .Z1(n1087) );
  CNIVX1 U1343 ( .A(n1087), .Z(n1086) );
  CIVDX1 U1344 ( .A(out0_stg0[59]), .Z1(n1089) );
  CNIVX1 U1345 ( .A(n1089), .Z(n1088) );
  CIVDX1 U1346 ( .A(out0_stg0[60]), .Z1(n1091) );
  CNIVX1 U1347 ( .A(n1091), .Z(n1090) );
  CIVDX1 U1348 ( .A(out0_stg0[61]), .Z1(n1093) );
  CNIVX1 U1349 ( .A(n1093), .Z(n1092) );
  CIVDX1 U1350 ( .A(out0_stg0[62]), .Z1(n1095) );
  CNIVX1 U1351 ( .A(n1095), .Z(n1094) );
  CIVDX1 U1352 ( .A(out0_stg0[63]), .Z1(n1097) );
  CNIVX1 U1353 ( .A(n1097), .Z(n1096) );
  CNIVX1 U1354 ( .A(n689), .Z(n1098) );
  CNIVX1 U1355 ( .A(n666), .Z(n1099) );
  CNIVX1 U1356 ( .A(n670), .Z(n1100) );
  CNIVX1 U1357 ( .A(n684), .Z(n1101) );
  CMX2XL U1358 ( .A0(q0[26]), .A1(q[26]), .S(n1380), .Z(n684) );
  CIVDX1 U1359 ( .A(push0_stg1), .Z1(n1103) );
  CNIVX1 U1360 ( .A(n1103), .Z(n1102) );
  CNIVX1 U1361 ( .A(n675), .Z(n1104) );
  CNIVX1 U1362 ( .A(h0[5]), .Z(n1105) );
  CNIVX1 U1363 ( .A(h0[1]), .Z(n1106) );
  CNIVX1 U1364 ( .A(h0[0]), .Z(n1107) );
  CNIVX1 U1365 ( .A(n679), .Z(n1108) );
  CNIVX1 U1366 ( .A(n680), .Z(n1109) );
  CMX2XL U1367 ( .A0(q0[22]), .A1(q[22]), .S(n1380), .Z(n680) );
  CIVDX1 U1368 ( .A(cmd0_stg0[1]), .Z1(n1111) );
  CNIVX1 U1369 ( .A(n1111), .Z(n1110) );
  CIVDX1 U1370 ( .A(cmd0_stg0[0]), .Z1(n1113) );
  CNIVX1 U1371 ( .A(n1113), .Z(n1112) );
  CIVDX1 U1372 ( .A(push0_stg0), .Z1(n1115) );
  CNIVX1 U1373 ( .A(n1115), .Z(n1114) );
  CNIVX1 U1374 ( .A(h0[4]), .Z(n1116) );
  CNIVX1 U1375 ( .A(n683), .Z(n1117) );
  CNIVX1 U1376 ( .A(n1119), .Z(n1118) );
  CNIVX1 U1377 ( .A(cmd0[1]), .Z(n1119) );
  CNIVX1 U1378 ( .A(n1121), .Z(n1120) );
  CNIVX1 U1379 ( .A(cmd0[0]), .Z(n1121) );
  CNIVX1 U1380 ( .A(n1123), .Z(n1122) );
  CNIVX1 U1381 ( .A(push0), .Z(n1123) );
  CNIVX1 U1382 ( .A(n650), .Z(n1124) );
  CNIVX1 U1383 ( .A(n657), .Z(n1125) );
  CIVX3 U1384 ( .A(rst), .Z(n1973) );
  CMX2XL U1385 ( .A0(n806), .A1(q[17]), .S(n1381), .Z(n675) );
  CMX2XL U1386 ( .A0(n794), .A1(q[18]), .S(n1381), .Z(n676) );
  CIVX3 U1387 ( .A(q0[16]), .Z(n1126) );
  CIVX8 U1388 ( .A(n1126), .Z(n1127) );
  CDLY1XL U1389 ( .A(q0[19]), .Z(n1128) );
  CDLY1XL U1390 ( .A(q0[29]), .Z(n1129) );
  CMX2XL U1391 ( .A0(n1127), .A1(q[16]), .S(n1381), .Z(n674) );
  CDLY1XL U1392 ( .A(q0[7]), .Z(n1130) );
  CDLY1XL U1393 ( .A(q0[13]), .Z(n1131) );
  CMX2XL U1394 ( .A0(h0[30]), .A1(h[30]), .S(n1382), .Z(n656) );
  CDLY1XL U1395 ( .A(h0[15]), .Z(n1132) );
  CDLY1XL U1396 ( .A(q0[1]), .Z(n1133) );
  CDLY1XL U1397 ( .A(q0[5]), .Z(n1134) );
  CDLY1XL U1398 ( .A(q0[11]), .Z(n1135) );
  CDLY1XL U1399 ( .A(q0[14]), .Z(n1208) );
  CMX2XL U1400 ( .A0(h0[14]), .A1(h[14]), .S(n1384), .Z(n640) );
  CIVXL U1401 ( .A(n795), .Z(n1136) );
  CIVX2 U1402 ( .A(n1136), .Z(n1137) );
  CDLY1XL U1403 ( .A(h0[28]), .Z(n1138) );
  CMX2XL U1404 ( .A0(h0[25]), .A1(h[25]), .S(n1383), .Z(n651) );
  CMX2XL U1405 ( .A0(q0[31]), .A1(q[31]), .S(n1380), .Z(n689) );
  CDLY1XL U1406 ( .A(q0[6]), .Z(n1139) );
  CDLY1XL U1407 ( .A(h0[26]), .Z(n1140) );
  CMX2XL U1408 ( .A0(q0[8]), .A1(q[8]), .S(n1381), .Z(n666) );
  CMX2XL U1409 ( .A0(n1139), .A1(q[6]), .S(n1382), .Z(n664) );
  CDLY1XL U1410 ( .A(h0[7]), .Z(n1141) );
  CMX2XL U1411 ( .A0(h0[11]), .A1(h[11]), .S(n1384), .Z(n637) );
  CMX2XL U1412 ( .A0(h0[13]), .A1(h[13]), .S(n1384), .Z(n639) );
  CMX2XL U1413 ( .A0(n803), .A1(q[25]), .S(n1380), .Z(n683) );
  CDLY1XL U1414 ( .A(q0[27]), .Z(n1209) );
  CMX2XL U1415 ( .A0(h0[22]), .A1(h[22]), .S(n1383), .Z(n648) );
  CMX2XL U1416 ( .A0(h0[21]), .A1(h[21]), .S(n1383), .Z(n647) );
  CMX2XL U1417 ( .A0(n796), .A1(q[9]), .S(n1381), .Z(n667) );
  CDLY1XL U1418 ( .A(q0[15]), .Z(n1142) );
  CMX2XL U1419 ( .A0(n1135), .A1(q[11]), .S(n1381), .Z(n669) );
  CMX2XL U1420 ( .A0(h0[9]), .A1(h[9]), .S(n1384), .Z(n635) );
  CMX2XL U1421 ( .A0(h0[18]), .A1(h[18]), .S(n1383), .Z(n644) );
  CMX2XL U1422 ( .A0(h0[17]), .A1(h[17]), .S(n1383), .Z(n643) );
  CDLY1XL U1423 ( .A(h0[2]), .Z(n1143) );
  CDLY1XL U1424 ( .A(h0[10]), .Z(n1144) );
  CDLY1XL U1425 ( .A(h0[12]), .Z(n1145) );
  CMX2XL U1426 ( .A0(n1106), .A1(h[1]), .S(n1385), .Z(n617) );
  CIVXL U1427 ( .A(n1106), .Z(n1911) );
  CANR2XL U1428 ( .A(n1759), .B(acc[24]), .C(n1758), .D(out0_stg2[24]), .Z(
        n1662) );
  CNR2XL U1429 ( .A(n2223), .B(n1219), .Z(n2264) );
  CND2X1 U1430 ( .A(n2179), .B(n1376), .Z(n2244) );
  CND2X1 U1431 ( .A(n2120), .B(n1376), .Z(n2183) );
  CMXI2XL U1432 ( .A0(n1900), .A1(n1204), .S(n1357), .Z(n2130) );
  CIVXL U1433 ( .A(n1899), .Z(n1900) );
  CANR2XL U1434 ( .A(n1759), .B(acc[63]), .C(n1758), .D(out0_stg2[63]), .Z(
        n1504) );
  CANR2XL U1435 ( .A(n1759), .B(acc[20]), .C(n1758), .D(out0_stg2[20]), .Z(
        n1678) );
  CANR2XL U1436 ( .A(acc[1]), .B(n1894), .C(out1_stg2[1]), .D(n1212), .Z(n1772) );
  CANR2XL U1437 ( .A(acc[2]), .B(n1894), .C(out1_stg2[2]), .D(n1212), .Z(n1774) );
  CANR2XL U1438 ( .A(acc[55]), .B(n1894), .C(out1_stg2[55]), .D(n1212), .Z(
        n1884) );
  CANR2XL U1439 ( .A(acc[52]), .B(n1894), .C(out1_stg2[52]), .D(n1212), .Z(
        n1874) );
  CANR2XL U1440 ( .A(acc[53]), .B(n1894), .C(out1_stg2[53]), .D(n1212), .Z(
        n1876) );
  CANR2XL U1441 ( .A(acc[54]), .B(n1894), .C(out1_stg2[54]), .D(n1212), .Z(
        n1878) );
  CANR2XL U1442 ( .A(acc[49]), .B(n1894), .C(out1_stg2[49]), .D(n1212), .Z(
        n1868) );
  CANR2XL U1443 ( .A(acc[50]), .B(n1894), .C(out1_stg2[50]), .D(n1212), .Z(
        n1870) );
  CANR2XL U1444 ( .A(acc[51]), .B(n1894), .C(out1_stg2[51]), .D(n1212), .Z(
        n1872) );
  CANR2XL U1445 ( .A(acc[48]), .B(n1894), .C(out1_stg2[48]), .D(n1212), .Z(
        n1866) );
  CANR2XL U1446 ( .A(acc[56]), .B(n1894), .C(out1_stg2[56]), .D(n1212), .Z(
        n1886) );
  CANR2XL U1447 ( .A(acc[47]), .B(n1894), .C(out1_stg2[47]), .D(n1212), .Z(
        n1864) );
  CANR2XL U1448 ( .A(acc[46]), .B(n1894), .C(out1_stg2[46]), .D(n1212), .Z(
        n1862) );
  CANR2XL U1449 ( .A(acc[45]), .B(n1894), .C(out1_stg2[45]), .D(n1212), .Z(
        n1860) );
  CANR2XL U1450 ( .A(acc[44]), .B(n1894), .C(out1_stg2[44]), .D(n1212), .Z(
        n1858) );
  CANR2XL U1451 ( .A(acc[41]), .B(n1894), .C(out1_stg2[41]), .D(n1212), .Z(
        n1852) );
  CANR2XL U1452 ( .A(acc[43]), .B(n1894), .C(out1_stg2[43]), .D(n1212), .Z(
        n1856) );
  CANR2XL U1453 ( .A(acc[42]), .B(n1894), .C(out1_stg2[42]), .D(n1212), .Z(
        n1854) );
  CANR2XL U1454 ( .A(acc[40]), .B(n1894), .C(out1_stg2[40]), .D(n1212), .Z(
        n1850) );
  CANR2XL U1455 ( .A(acc[39]), .B(n1894), .C(out1_stg2[39]), .D(n1212), .Z(
        n1848) );
  CANR2XL U1456 ( .A(acc[38]), .B(n1894), .C(out1_stg2[38]), .D(n1212), .Z(
        n1846) );
  CANR2XL U1457 ( .A(acc[37]), .B(n1894), .C(out1_stg2[37]), .D(n1212), .Z(
        n1844) );
  CANR2XL U1458 ( .A(acc[36]), .B(n1894), .C(out1_stg2[36]), .D(n1212), .Z(
        n1842) );
  CANR2XL U1459 ( .A(acc[35]), .B(n1894), .C(out1_stg2[35]), .D(n1212), .Z(
        n1840) );
  CANR2XL U1460 ( .A(acc[34]), .B(n1894), .C(out1_stg2[34]), .D(n1212), .Z(
        n1838) );
  CANR2XL U1461 ( .A(acc[33]), .B(n1894), .C(out1_stg2[33]), .D(n1212), .Z(
        n1836) );
  CANR2XL U1462 ( .A(acc[32]), .B(n1894), .C(out1_stg2[32]), .D(n1212), .Z(
        n1834) );
  CANR2XL U1463 ( .A(acc[31]), .B(n1894), .C(out1_stg2[31]), .D(n1212), .Z(
        n1832) );
  CANR2XL U1464 ( .A(acc[30]), .B(n1894), .C(out1_stg2[30]), .D(n1212), .Z(
        n1830) );
  CANR2XL U1465 ( .A(acc[29]), .B(n1894), .C(out1_stg2[29]), .D(n1212), .Z(
        n1828) );
  CANR2XL U1466 ( .A(acc[28]), .B(n1894), .C(out1_stg2[28]), .D(n1212), .Z(
        n1826) );
  CANR2XL U1467 ( .A(acc[27]), .B(n1894), .C(out1_stg2[27]), .D(n1212), .Z(
        n1824) );
  CANR2XL U1468 ( .A(acc[26]), .B(n1894), .C(out1_stg2[26]), .D(n1212), .Z(
        n1822) );
  CANR2XL U1469 ( .A(acc[25]), .B(n1894), .C(out1_stg2[25]), .D(n1212), .Z(
        n1820) );
  CANR2XL U1470 ( .A(acc[24]), .B(n1894), .C(out1_stg2[24]), .D(n1212), .Z(
        n1818) );
  CANR2XL U1471 ( .A(acc[23]), .B(n1894), .C(out1_stg2[23]), .D(n1212), .Z(
        n1816) );
  CANR2XL U1472 ( .A(acc[22]), .B(n1894), .C(out1_stg2[22]), .D(n1212), .Z(
        n1814) );
  CANR2XL U1473 ( .A(acc[21]), .B(n1894), .C(out1_stg2[21]), .D(n1212), .Z(
        n1812) );
  CANR2XL U1474 ( .A(acc[20]), .B(n1894), .C(out1_stg2[20]), .D(n1212), .Z(
        n1810) );
  CANR2XL U1475 ( .A(acc[19]), .B(n1894), .C(out1_stg2[19]), .D(n1212), .Z(
        n1808) );
  CANR2XL U1476 ( .A(acc[18]), .B(n1894), .C(out1_stg2[18]), .D(n1212), .Z(
        n1806) );
  CANR2XL U1477 ( .A(acc[17]), .B(n1894), .C(out1_stg2[17]), .D(n1212), .Z(
        n1804) );
  CANR2XL U1478 ( .A(acc[16]), .B(n1894), .C(out1_stg2[16]), .D(n1212), .Z(
        n1802) );
  CANR2XL U1479 ( .A(acc[15]), .B(n1894), .C(out1_stg2[15]), .D(n1212), .Z(
        n1800) );
  CANR2XL U1480 ( .A(acc[14]), .B(n1894), .C(out1_stg2[14]), .D(n1212), .Z(
        n1798) );
  CANR2XL U1481 ( .A(acc[13]), .B(n1894), .C(out1_stg2[13]), .D(n1212), .Z(
        n1796) );
  CANR2XL U1482 ( .A(acc[12]), .B(n1894), .C(out1_stg2[12]), .D(n1212), .Z(
        n1794) );
  CANR2XL U1483 ( .A(acc[11]), .B(n1894), .C(out1_stg2[11]), .D(n1212), .Z(
        n1792) );
  CANR2XL U1484 ( .A(acc[10]), .B(n1894), .C(out1_stg2[10]), .D(n1212), .Z(
        n1790) );
  CANR2XL U1485 ( .A(acc[9]), .B(n1894), .C(out1_stg2[9]), .D(n1212), .Z(n1788) );
  CANR2XL U1486 ( .A(acc[8]), .B(n1894), .C(out1_stg2[8]), .D(n1212), .Z(n1786) );
  CANR2XL U1487 ( .A(acc[7]), .B(n1894), .C(out1_stg2[7]), .D(n1212), .Z(n1784) );
  CANR2XL U1488 ( .A(acc[6]), .B(n1894), .C(out1_stg2[6]), .D(n1212), .Z(n1782) );
  CANR2XL U1489 ( .A(acc[5]), .B(n1894), .C(out1_stg2[5]), .D(n1212), .Z(n1780) );
  CANR2XL U1490 ( .A(acc[4]), .B(n1894), .C(out1_stg2[4]), .D(n1212), .Z(n1778) );
  CANR2XL U1491 ( .A(acc[3]), .B(n1894), .C(out1_stg2[3]), .D(n1212), .Z(n1776) );
  CANR2XL U1492 ( .A(n1759), .B(acc[18]), .C(n1758), .D(out0_stg2[18]), .Z(
        n1686) );
  CANR2XL U1493 ( .A(n1759), .B(acc[2]), .C(n1758), .D(out0_stg2[2]), .Z(n1750) );
  CANR2XL U1494 ( .A(n1759), .B(acc[11]), .C(n1758), .D(out0_stg2[11]), .Z(
        n1714) );
  CANR2XL U1495 ( .A(n1759), .B(acc[10]), .C(n1758), .D(out0_stg2[10]), .Z(
        n1718) );
  CANR2XL U1496 ( .A(n1759), .B(acc[23]), .C(n1758), .D(out0_stg2[23]), .Z(
        n1666) );
  CANR2XL U1497 ( .A(n1759), .B(acc[17]), .C(n1758), .D(out0_stg2[17]), .Z(
        n1690) );
  CANR2XL U1498 ( .A(n1759), .B(acc[25]), .C(n1758), .D(out0_stg2[25]), .Z(
        n1658) );
  CANR2XL U1499 ( .A(n1759), .B(acc[8]), .C(n1758), .D(out0_stg2[8]), .Z(n1726) );
  CANR2XL U1500 ( .A(n1759), .B(acc[19]), .C(n1758), .D(out0_stg2[19]), .Z(
        n1682) );
  CANR2XL U1501 ( .A(n1759), .B(acc[22]), .C(n1758), .D(out0_stg2[22]), .Z(
        n1670) );
  CANR2XL U1502 ( .A(n1759), .B(acc[6]), .C(n1758), .D(out0_stg2[6]), .Z(n1734) );
  CANR2XL U1503 ( .A(n1759), .B(acc[26]), .C(n1758), .D(out0_stg2[26]), .Z(
        n1654) );
  CANR2XL U1504 ( .A(n1759), .B(acc[28]), .C(n1758), .D(out0_stg2[28]), .Z(
        n1646) );
  CANR2XL U1505 ( .A(n1759), .B(acc[16]), .C(n1758), .D(out0_stg2[16]), .Z(
        n1694) );
  CANR2XL U1506 ( .A(n1759), .B(acc[27]), .C(n1758), .D(out0_stg2[27]), .Z(
        n1650) );
  CANR2XL U1507 ( .A(n1759), .B(acc[29]), .C(n1758), .D(out0_stg2[29]), .Z(
        n1642) );
  CANR2XL U1508 ( .A(n1759), .B(acc[4]), .C(n1758), .D(out0_stg2[4]), .Z(n1742) );
  CANR2XL U1509 ( .A(n1759), .B(acc[3]), .C(n1758), .D(out0_stg2[3]), .Z(n1746) );
  CANR2XL U1510 ( .A(n1759), .B(acc[14]), .C(n1758), .D(out0_stg2[14]), .Z(
        n1702) );
  CANR2XL U1511 ( .A(n1759), .B(acc[15]), .C(n1758), .D(out0_stg2[15]), .Z(
        n1698) );
  CANR2XL U1512 ( .A(n1759), .B(acc[7]), .C(n1758), .D(out0_stg2[7]), .Z(n1730) );
  CANR2XL U1513 ( .A(n1759), .B(acc[35]), .C(n1758), .D(out0_stg2[35]), .Z(
        n1618) );
  CANR2XL U1514 ( .A(n1759), .B(acc[13]), .C(n1758), .D(out0_stg2[13]), .Z(
        n1706) );
  CANR2XL U1515 ( .A(n1759), .B(acc[41]), .C(n1758), .D(out0_stg2[41]), .Z(
        n1594) );
  CANR2XL U1516 ( .A(n1759), .B(acc[21]), .C(n1758), .D(out0_stg2[21]), .Z(
        n1674) );
  CANR2XL U1517 ( .A(n1759), .B(acc[5]), .C(n1758), .D(out0_stg2[5]), .Z(n1738) );
  CANR2XL U1518 ( .A(n1759), .B(acc[30]), .C(n1758), .D(out0_stg2[30]), .Z(
        n1638) );
  CANR2XL U1519 ( .A(n1759), .B(acc[12]), .C(n1758), .D(out0_stg2[12]), .Z(
        n1710) );
  CANR2XL U1520 ( .A(n1759), .B(acc[31]), .C(n1758), .D(out0_stg2[31]), .Z(
        n1634) );
  CANR2XL U1521 ( .A(n1759), .B(acc[49]), .C(n1758), .D(out0_stg2[49]), .Z(
        n1562) );
  CANR2XL U1522 ( .A(n1759), .B(acc[33]), .C(n1758), .D(out0_stg2[33]), .Z(
        n1626) );
  CANR2XL U1523 ( .A(n1759), .B(acc[40]), .C(n1758), .D(out0_stg2[40]), .Z(
        n1598) );
  CANR2XL U1524 ( .A(n1759), .B(acc[34]), .C(n1758), .D(out0_stg2[34]), .Z(
        n1622) );
  CANR2XL U1525 ( .A(n1759), .B(acc[42]), .C(n1758), .D(out0_stg2[42]), .Z(
        n1590) );
  CANR2XL U1526 ( .A(n1759), .B(acc[43]), .C(n1758), .D(out0_stg2[43]), .Z(
        n1586) );
  CANR2XL U1527 ( .A(n1759), .B(acc[58]), .C(n1758), .D(out0_stg2[58]), .Z(
        n1526) );
  CANR2XL U1528 ( .A(n1759), .B(acc[57]), .C(n1758), .D(out0_stg2[57]), .Z(
        n1530) );
  CANR2XL U1529 ( .A(n1759), .B(acc[50]), .C(n1758), .D(out0_stg2[50]), .Z(
        n1558) );
  CANR2XL U1530 ( .A(n1759), .B(acc[48]), .C(n1758), .D(out0_stg2[48]), .Z(
        n1566) );
  CANR2XL U1531 ( .A(n1759), .B(acc[51]), .C(n1758), .D(out0_stg2[51]), .Z(
        n1554) );
  CANR2XL U1532 ( .A(n1759), .B(acc[56]), .C(n1758), .D(out0_stg2[56]), .Z(
        n1534) );
  CANR2XL U1533 ( .A(n1759), .B(acc[52]), .C(n1758), .D(out0_stg2[52]), .Z(
        n1550) );
  CANR2XL U1534 ( .A(n1759), .B(acc[32]), .C(n1758), .D(out0_stg2[32]), .Z(
        n1630) );
  CANR2XL U1535 ( .A(n1759), .B(acc[59]), .C(n1758), .D(out0_stg2[59]), .Z(
        n1522) );
  CANR2XL U1536 ( .A(n1759), .B(acc[44]), .C(n1758), .D(out0_stg2[44]), .Z(
        n1582) );
  CANR2XL U1537 ( .A(n1759), .B(acc[45]), .C(n1758), .D(out0_stg2[45]), .Z(
        n1578) );
  CANR2XL U1538 ( .A(n1759), .B(acc[53]), .C(n1758), .D(out0_stg2[53]), .Z(
        n1546) );
  CANR2XL U1539 ( .A(n1759), .B(acc[47]), .C(n1758), .D(out0_stg2[47]), .Z(
        n1570) );
  CANR2XL U1540 ( .A(n1759), .B(acc[38]), .C(n1758), .D(out0_stg2[38]), .Z(
        n1606) );
  CANR2XL U1541 ( .A(n1759), .B(acc[39]), .C(n1758), .D(out0_stg2[39]), .Z(
        n1602) );
  CANR2XL U1542 ( .A(n1759), .B(acc[36]), .C(n1758), .D(out0_stg2[36]), .Z(
        n1614) );
  CANR2XL U1543 ( .A(n1759), .B(acc[55]), .C(n1758), .D(out0_stg2[55]), .Z(
        n1538) );
  CANR2XL U1544 ( .A(n1759), .B(acc[54]), .C(n1758), .D(out0_stg2[54]), .Z(
        n1542) );
  CANR2XL U1545 ( .A(n1759), .B(acc[46]), .C(n1758), .D(out0_stg2[46]), .Z(
        n1574) );
  CANR2XL U1546 ( .A(acc[63]), .B(n1894), .C(out1_stg2[63]), .D(n1212), .Z(
        n1768) );
  CANR2XL U1547 ( .A(n1759), .B(acc[37]), .C(n1758), .D(out0_stg2[37]), .Z(
        n1610) );
  CANR2XL U1548 ( .A(n1759), .B(acc[60]), .C(n1758), .D(out0_stg2[60]), .Z(
        n1518) );
  CANR2XL U1549 ( .A(n1759), .B(acc[61]), .C(n1758), .D(out0_stg2[61]), .Z(
        n1514) );
  CANR2XL U1550 ( .A(acc[62]), .B(n1894), .C(out1_stg2[62]), .D(n1212), .Z(
        n1892) );
  CANR2XL U1551 ( .A(acc[0]), .B(n1894), .C(out1_stg2[0]), .D(n1212), .Z(n1770) );
  CANR2XL U1552 ( .A(acc[61]), .B(n1894), .C(out1_stg2[61]), .D(n1212), .Z(
        n1895) );
  CANR2XL U1553 ( .A(acc[60]), .B(n1894), .C(out1_stg2[60]), .D(n1212), .Z(
        n1888) );
  CANR2XL U1554 ( .A(acc[58]), .B(n1894), .C(out1_stg2[58]), .D(n1212), .Z(
        n1880) );
  CANR2XL U1555 ( .A(acc[59]), .B(n1894), .C(out1_stg2[59]), .D(n1212), .Z(
        n1890) );
  CANR2XL U1556 ( .A(n1759), .B(acc[62]), .C(n1758), .D(out0_stg2[62]), .Z(
        n1510) );
  CANR2XL U1557 ( .A(n2217), .B(n1146), .C(n2218), .D(n1300), .Z(n1437) );
  CANR2XL U1558 ( .A(n1206), .B(out0_stg2[11]), .C(N429), .D(n1205), .Z(n1713)
         );
  CANR2XL U1559 ( .A(n1206), .B(out0_stg2[9]), .C(N427), .D(n1205), .Z(n1721)
         );
  CANR2XL U1560 ( .A(n1206), .B(out0_stg2[3]), .C(N421), .D(n1205), .Z(n1745)
         );
  CANR2XL U1561 ( .A(n1206), .B(out0_stg2[1]), .C(N419), .D(n1205), .Z(n1753)
         );
  CANR2XL U1562 ( .A(n1207), .B(out1_stg2[0]), .C(acc[0]), .D(n802), .Z(n1756)
         );
  CANR2XL U1563 ( .A(n1206), .B(out0_stg2[0]), .C(N418), .D(n1205), .Z(n1757)
         );
  CMXI2XL U1564 ( .A0(n1991), .A1(n2284), .S(n1225), .Z(n1147) );
  CND2XL U1565 ( .A(n1378), .B(n1356), .Z(n1148) );
  CIVX1 U1566 ( .A(n2270), .Z(n1979) );
  CIVXL U1567 ( .A(n2269), .Z(n1978) );
  CNIVX1 U1568 ( .A(n1436), .Z(n1211) );
  CNIVX1 U1569 ( .A(n1436), .Z(n1210) );
  CIVX4 U1570 ( .A(n1501), .Z(n1762) );
  CIVX4 U1571 ( .A(n1502), .Z(n1759) );
  CIVX2 U1572 ( .A(n1370), .Z(n1366) );
  CIVX2 U1573 ( .A(n1370), .Z(n1365) );
  CIVX2 U1574 ( .A(n1370), .Z(n1367) );
  CIVX2 U1575 ( .A(n1370), .Z(n1368) );
  CIVX2 U1576 ( .A(n1363), .Z(n1357) );
  CIVX2 U1577 ( .A(n1363), .Z(n1359) );
  CIVX2 U1578 ( .A(n1363), .Z(n1360) );
  CIVX2 U1579 ( .A(n1363), .Z(n1361) );
  CIVX2 U1580 ( .A(n1363), .Z(n1358) );
  CNR2X1 U1581 ( .A(n2096), .B(n1213), .Z(n2165) );
  CNR2XL U1582 ( .A(n2113), .B(n1215), .Z(n2151) );
  CNR2XL U1583 ( .A(n2081), .B(n1214), .Z(n2158) );
  CNR2X1 U1584 ( .A(n2037), .B(n1216), .Z(n2172) );
  CNR2IX1 U1585 ( .B(acc_cmd2[63]), .A(n1357), .Z(n2019) );
  CNR2X1 U1586 ( .A(n2215), .B(n1221), .Z(n2283) );
  CNR2X1 U1587 ( .A(n2244), .B(n1219), .Z(n2269) );
  CNR2X1 U1588 ( .A(n2183), .B(n1218), .Z(n2270) );
  CNR2XL U1589 ( .A(n2137), .B(n1219), .Z(n2253) );
  CNR2X1 U1590 ( .A(n2191), .B(n1218), .Z(n2280) );
  CNR2X1 U1591 ( .A(n2187), .B(n1222), .Z(n2271) );
  CNR2XL U1592 ( .A(n2206), .B(n1218), .Z(n2262) );
  CNR2X1 U1593 ( .A(n2221), .B(n1223), .Z(n2263) );
  CNR2XL U1594 ( .A(n2242), .B(n1220), .Z(n2268) );
  CNR2XL U1595 ( .A(n2229), .B(n1221), .Z(n2267) );
  CNR2XL U1596 ( .A(n2227), .B(n1222), .Z(n2266) );
  CNR2XL U1597 ( .A(n2225), .B(n1223), .Z(n2265) );
  CNR2X1 U1598 ( .A(n2195), .B(n1223), .Z(n2281) );
  CNR2X1 U1599 ( .A(n2211), .B(n1222), .Z(n2282) );
  CND3XL U1600 ( .A(n1379), .B(n1765), .C(n1767), .Z(n1766) );
  CNR2X1 U1601 ( .A(n2100), .B(n1220), .Z(n2217) );
  CNIVX1 U1602 ( .A(n1897), .Z(n1304) );
  CNIVX1 U1603 ( .A(n1897), .Z(n1303) );
  CNIVX1 U1604 ( .A(n1897), .Z(n1302) );
  CNIVX1 U1605 ( .A(n1897), .Z(n1305) );
  CNIVX1 U1606 ( .A(n1897), .Z(n1301) );
  CIVX2 U1607 ( .A(n1370), .Z(n1364) );
  CNIVX1 U1608 ( .A(n1897), .Z(n1306) );
  CND2XL U1609 ( .A(n2065), .B(n1370), .Z(n2096) );
  CND2X1 U1610 ( .A(n2165), .B(n1376), .Z(n2215) );
  CND2X1 U1611 ( .A(n2127), .B(n1376), .Z(n2187) );
  CND2X1 U1612 ( .A(n2144), .B(n1376), .Z(n2191) );
  CND2XL U1613 ( .A(n2151), .B(n1376), .Z(n2195) );
  CND2XL U1614 ( .A(n2158), .B(n1376), .Z(n2211) );
  CND2X1 U1615 ( .A(n2019), .B(n1370), .Z(n2037) );
  CND2X1 U1616 ( .A(n2172), .B(n1376), .Z(n2100) );
  CND3XL U1617 ( .A(n1378), .B(n1435), .C(n1386), .Z(n1436) );
  CAN3X2 U1618 ( .A(n1224), .B(n1378), .C(n1435), .Z(n1146) );
  CIVX2 U1619 ( .A(n1376), .Z(n1374) );
  CIVX2 U1620 ( .A(n1376), .Z(n1372) );
  CIVX2 U1621 ( .A(n1376), .Z(n1373) );
  CNR3XL U1622 ( .A(n802), .B(n1974), .C(n1975), .Z(_pushout_d) );
  CIVX2 U1623 ( .A(n1376), .Z(n1375) );
  CIVX2 U1624 ( .A(n1376), .Z(n1371) );
  CNIVX1 U1625 ( .A(n1973), .Z(n1342) );
  CNIVX1 U1626 ( .A(n1973), .Z(n1326) );
  CNIVX1 U1627 ( .A(n1973), .Z(n1327) );
  CNIVX1 U1628 ( .A(n1973), .Z(n1328) );
  CNIVX1 U1629 ( .A(n1973), .Z(n1341) );
  CNIVX1 U1630 ( .A(n1973), .Z(n1322) );
  CNIVX1 U1631 ( .A(n1973), .Z(n1325) );
  CNIVX1 U1632 ( .A(n1973), .Z(n1343) );
  CNIVX1 U1633 ( .A(n1973), .Z(n1339) );
  CNIVX1 U1634 ( .A(n1973), .Z(n1324) );
  CNIVX1 U1635 ( .A(n1973), .Z(n1340) );
  CNIVX1 U1636 ( .A(n1973), .Z(n1314) );
  CNIVX1 U1637 ( .A(n1973), .Z(n1312) );
  CNIVX1 U1638 ( .A(n1973), .Z(n1311) );
  CNIVX1 U1639 ( .A(n1973), .Z(n1310) );
  CNIVX1 U1640 ( .A(n1973), .Z(n1309) );
  CNIVX1 U1641 ( .A(n1973), .Z(n1338) );
  CNIVX1 U1642 ( .A(n1973), .Z(n1337) );
  CNIVX1 U1643 ( .A(n1973), .Z(n1336) );
  CNIVX1 U1644 ( .A(n1973), .Z(n1335) );
  CNIVX1 U1645 ( .A(n1973), .Z(n1334) );
  CNIVX1 U1646 ( .A(n1973), .Z(n1333) );
  CNIVX1 U1647 ( .A(n1973), .Z(n1332) );
  CNIVX1 U1648 ( .A(n1973), .Z(n1355) );
  CNIVX1 U1649 ( .A(n1973), .Z(n1354) );
  CNIVX1 U1650 ( .A(n1973), .Z(n1353) );
  CNIVX1 U1651 ( .A(n1973), .Z(n1352) );
  CNIVX1 U1652 ( .A(n1973), .Z(n1351) );
  CNIVX1 U1653 ( .A(n1973), .Z(n1350) );
  CNIVX1 U1654 ( .A(n1973), .Z(n1349) );
  CNIVX1 U1655 ( .A(n1973), .Z(n1348) );
  CNIVX1 U1656 ( .A(n1973), .Z(n1323) );
  CNIVX1 U1657 ( .A(n1973), .Z(n1321) );
  CNIVX1 U1658 ( .A(n1973), .Z(n1320) );
  CNIVX1 U1659 ( .A(n1973), .Z(n1313) );
  CNIVX1 U1660 ( .A(n1973), .Z(n1347) );
  CNIVX1 U1661 ( .A(n1973), .Z(n1319) );
  CNIVX1 U1662 ( .A(n1973), .Z(n1308) );
  CNIVX1 U1663 ( .A(n1973), .Z(n1345) );
  CNIVX1 U1664 ( .A(n1973), .Z(n1316) );
  CNIVX1 U1665 ( .A(n1973), .Z(n1346) );
  CNIVX1 U1666 ( .A(n1973), .Z(n1344) );
  CNIVX1 U1667 ( .A(n1973), .Z(n1318) );
  CNIVX1 U1668 ( .A(n1973), .Z(n1317) );
  CNIVX1 U1669 ( .A(n1973), .Z(n1315) );
  CNIVX1 U1670 ( .A(n1973), .Z(n1307) );
  CNIVX1 U1671 ( .A(n1973), .Z(n1331) );
  CNIVX1 U1672 ( .A(n1973), .Z(n1329) );
  CNIVX1 U1673 ( .A(n1973), .Z(n1330) );
  CNIVX1 U1674 ( .A(n1973), .Z(n1356) );
  COND1XL U1675 ( .A(n1762), .B(n1571), .C(n1570), .Z(acc_cmd1[47]) );
  COND1XL U1676 ( .A(n1762), .B(n1567), .C(n1566), .Z(acc_cmd1[48]) );
  COND1XL U1677 ( .A(n1762), .B(n1667), .C(n1666), .Z(acc_cmd1[23]) );
  COND1XL U1678 ( .A(n1762), .B(n1679), .C(n1678), .Z(acc_cmd1[20]) );
  COND1XL U1679 ( .A(n1762), .B(n1583), .C(n1582), .Z(acc_cmd1[44]) );
  COND1XL U1680 ( .A(n1762), .B(n1647), .C(n1646), .Z(acc_cmd1[28]) );
  COND1XL U1681 ( .A(n1762), .B(n1671), .C(n1670), .Z(acc_cmd1[22]) );
  COND1XL U1682 ( .A(n1762), .B(n1551), .C(n1550), .Z(acc_cmd1[52]) );
  COND1XL U1683 ( .A(n1762), .B(n1655), .C(n1654), .Z(acc_cmd1[26]) );
  COND1XL U1684 ( .A(n1762), .B(n1663), .C(n1662), .Z(acc_cmd1[24]) );
  COND1XL U1685 ( .A(n1762), .B(n1563), .C(n1562), .Z(acc_cmd1[49]) );
  COND1XL U1686 ( .A(n1762), .B(n1559), .C(n1558), .Z(acc_cmd1[50]) );
  COND1XL U1687 ( .A(n1762), .B(n1695), .C(n1694), .Z(acc_cmd1[16]) );
  COND1XL U1688 ( .A(n1762), .B(n1643), .C(n1642), .Z(acc_cmd1[29]) );
  COND1XL U1689 ( .A(n1762), .B(n1675), .C(n1674), .Z(acc_cmd1[21]) );
  COND1XL U1690 ( .A(n1762), .B(n1547), .C(n1546), .Z(acc_cmd1[53]) );
  COND1XL U1691 ( .A(n1762), .B(n1751), .C(n1750), .Z(acc_cmd1[2]) );
  COND1XL U1692 ( .A(n1762), .B(n1635), .C(n1634), .Z(acc_cmd1[31]) );
  COND1XL U1693 ( .A(n1762), .B(n1543), .C(n1542), .Z(acc_cmd1[54]) );
  COND1XL U1694 ( .A(n1762), .B(n1703), .C(n1702), .Z(acc_cmd1[14]) );
  COND1XL U1695 ( .A(n1762), .B(n1711), .C(n1710), .Z(acc_cmd1[12]) );
  COND1XL U1696 ( .A(n1762), .B(n1761), .C(n1760), .Z(acc_cmd1[0]) );
  COND1XL U1697 ( .A(n1762), .B(n1555), .C(n1554), .Z(acc_cmd1[51]) );
  COND1XL U1698 ( .A(n1762), .B(n1535), .C(n1534), .Z(acc_cmd1[56]) );
  COND1XL U1699 ( .A(n1762), .B(n1743), .C(n1742), .Z(acc_cmd1[4]) );
  COND1XL U1700 ( .A(n1762), .B(n1539), .C(n1538), .Z(acc_cmd1[55]) );
  COND1XL U1701 ( .A(n1762), .B(n1527), .C(n1526), .Z(acc_cmd1[58]) );
  COND1XL U1702 ( .A(n1762), .B(n1531), .C(n1530), .Z(acc_cmd1[57]) );
  COND1XL U1703 ( .A(n1762), .B(n1523), .C(n1522), .Z(acc_cmd1[59]) );
  COND1XL U1704 ( .A(n1762), .B(n1515), .C(n1514), .Z(acc_cmd1[61]) );
  COND1XL U1705 ( .A(n1762), .B(n1519), .C(n1518), .Z(acc_cmd1[60]) );
  COND1XL U1706 ( .A(n1762), .B(n1511), .C(n1510), .Z(acc_cmd1[62]) );
  COND1XL U1707 ( .A(n1762), .B(n1505), .C(n1504), .Z(acc_cmd1[63]) );
  CIVX4 U1708 ( .A(n1503), .Z(n1758) );
  COND1XL U1709 ( .A(n1305), .B(n1883), .C(n1882), .Z(acc_cmd2[57]) );
  COND1XL U1710 ( .A(n1301), .B(n1771), .C(n1770), .Z(n1899) );
  COND1XL U1711 ( .A(n1762), .B(n1623), .C(n1622), .Z(acc_cmd1[34]) );
  COND1XL U1712 ( .A(n1762), .B(n1575), .C(n1574), .Z(acc_cmd1[46]) );
  COND1XL U1713 ( .A(n1762), .B(n1591), .C(n1590), .Z(acc_cmd1[42]) );
  COND1XL U1714 ( .A(n1762), .B(n1687), .C(n1686), .Z(acc_cmd1[18]) );
  COND1XL U1715 ( .A(n1762), .B(n1595), .C(n1594), .Z(acc_cmd1[41]) );
  COND1XL U1716 ( .A(n1762), .B(n1579), .C(n1578), .Z(acc_cmd1[45]) );
  COND1XL U1717 ( .A(n1762), .B(n1659), .C(n1658), .Z(acc_cmd1[25]) );
  COND1XL U1718 ( .A(n1762), .B(n1607), .C(n1606), .Z(acc_cmd1[38]) );
  COND1XL U1719 ( .A(n1762), .B(n1691), .C(n1690), .Z(acc_cmd1[17]) );
  COND1XL U1720 ( .A(n1762), .B(n1715), .C(n1714), .Z(acc_cmd1[11]) );
  COND1XL U1721 ( .A(n1762), .B(n1619), .C(n1618), .Z(acc_cmd1[35]) );
  COND1XL U1722 ( .A(n1762), .B(n1599), .C(n1598), .Z(acc_cmd1[40]) );
  COND1XL U1723 ( .A(n1762), .B(n1627), .C(n1626), .Z(acc_cmd1[33]) );
  COND1XL U1724 ( .A(n1762), .B(n1587), .C(n1586), .Z(acc_cmd1[43]) );
  COND1XL U1725 ( .A(n1762), .B(n1683), .C(n1682), .Z(acc_cmd1[19]) );
  COND1XL U1726 ( .A(n1762), .B(n1603), .C(n1602), .Z(acc_cmd1[39]) );
  COND1XL U1727 ( .A(n1762), .B(n1615), .C(n1614), .Z(acc_cmd1[36]) );
  COND1XL U1728 ( .A(n1762), .B(n1719), .C(n1718), .Z(acc_cmd1[10]) );
  COND1XL U1729 ( .A(n1762), .B(n1639), .C(n1638), .Z(acc_cmd1[30]) );
  COND1XL U1730 ( .A(n1762), .B(n1699), .C(n1698), .Z(acc_cmd1[15]) );
  COND1XL U1731 ( .A(n1762), .B(n1651), .C(n1650), .Z(acc_cmd1[27]) );
  COND1XL U1732 ( .A(n1762), .B(n1723), .C(n1722), .Z(acc_cmd1[9]) );
  COND1XL U1733 ( .A(n1762), .B(n1707), .C(n1706), .Z(acc_cmd1[13]) );
  COND1XL U1734 ( .A(n1762), .B(n1611), .C(n1610), .Z(acc_cmd1[37]) );
  COND1XL U1735 ( .A(n1762), .B(n1735), .C(n1734), .Z(acc_cmd1[6]) );
  COND1XL U1736 ( .A(n1762), .B(n1731), .C(n1730), .Z(acc_cmd1[7]) );
  COND1XL U1737 ( .A(n1762), .B(n1727), .C(n1726), .Z(acc_cmd1[8]) );
  COND1XL U1738 ( .A(n1762), .B(n1739), .C(n1738), .Z(acc_cmd1[5]) );
  COND1XL U1739 ( .A(n1762), .B(n1631), .C(n1630), .Z(acc_cmd1[32]) );
  COND1XL U1740 ( .A(n1762), .B(n1747), .C(n1746), .Z(acc_cmd1[3]) );
  COND1XL U1741 ( .A(n1762), .B(n1755), .C(n1754), .Z(acc_cmd1[1]) );
  COND1XL U1742 ( .A(n1301), .B(n1769), .C(n1768), .Z(acc_cmd2[63]) );
  COND1XL U1743 ( .A(n1306), .B(n1893), .C(n1892), .Z(acc_cmd2[62]) );
  COND1XL U1744 ( .A(n1306), .B(n1889), .C(n1888), .Z(acc_cmd2[60]) );
  COND1XL U1745 ( .A(n1306), .B(n1896), .C(n1895), .Z(acc_cmd2[61]) );
  COND1XL U1746 ( .A(n1306), .B(n1891), .C(n1890), .Z(acc_cmd2[59]) );
  COND1XL U1747 ( .A(n1305), .B(n1881), .C(n1880), .Z(acc_cmd2[58]) );
  CMX2X1 U1748 ( .A0(n1147), .A1(roundit), .S(n1148), .Z(n611) );
  COND1XL U1749 ( .A(n1378), .B(n1446), .C(n1445), .Z(n583) );
  COND1XL U1750 ( .A(n1378), .B(n1448), .C(n1447), .Z(n584) );
  COND1XL U1751 ( .A(n1378), .B(n1450), .C(n1449), .Z(n585) );
  COND1XL U1752 ( .A(n1379), .B(n1500), .C(n1499), .Z(n610) );
  COND1XL U1753 ( .A(n1379), .B(n1498), .C(n1497), .Z(n609) );
  COND1XL U1754 ( .A(n1379), .B(n1494), .C(n1493), .Z(n607) );
  COND1XL U1755 ( .A(n1379), .B(n1496), .C(n1495), .Z(n608) );
  COND1XL U1756 ( .A(n1378), .B(n1438), .C(n1437), .Z(n579) );
  COND1XL U1757 ( .A(n1379), .B(n1486), .C(n1485), .Z(n603) );
  COND1XL U1758 ( .A(n1379), .B(n1488), .C(n1487), .Z(n604) );
  COND1XL U1759 ( .A(n1379), .B(n1490), .C(n1489), .Z(n605) );
  COND1XL U1760 ( .A(n1379), .B(n1492), .C(n1491), .Z(n606) );
  COND1XL U1761 ( .A(n1378), .B(n1440), .C(n1439), .Z(n580) );
  COND1XL U1762 ( .A(n1378), .B(n1442), .C(n1441), .Z(n581) );
  COND1XL U1763 ( .A(n1378), .B(n1444), .C(n1443), .Z(n582) );
  COND1XL U1764 ( .A(n1379), .B(n1468), .C(n1467), .Z(n594) );
  COND1XL U1765 ( .A(n1379), .B(n1466), .C(n1465), .Z(n593) );
  COND1XL U1766 ( .A(n1379), .B(n1484), .C(n1483), .Z(n602) );
  COND1XL U1767 ( .A(n1379), .B(n1470), .C(n1469), .Z(n595) );
  COND1XL U1768 ( .A(n1379), .B(n1472), .C(n1471), .Z(n596) );
  COND1XL U1769 ( .A(n1379), .B(n1474), .C(n1473), .Z(n597) );
  COND1XL U1770 ( .A(n1379), .B(n1476), .C(n1475), .Z(n598) );
  COND1XL U1771 ( .A(n1379), .B(n1482), .C(n1481), .Z(n601) );
  COND1XL U1772 ( .A(n1378), .B(n1462), .C(n1461), .Z(n591) );
  COND1XL U1773 ( .A(n1379), .B(n1464), .C(n1463), .Z(n592) );
  COND1XL U1774 ( .A(n1379), .B(n1478), .C(n1477), .Z(n599) );
  COND1XL U1775 ( .A(n1379), .B(n1480), .C(n1479), .Z(n600) );
  COND1XL U1776 ( .A(n1378), .B(n1454), .C(n1453), .Z(n587) );
  COND1XL U1777 ( .A(n1378), .B(n1456), .C(n1455), .Z(n588) );
  COND1XL U1778 ( .A(n1378), .B(n1458), .C(n1457), .Z(n589) );
  COND1XL U1779 ( .A(n1378), .B(n1460), .C(n1459), .Z(n590) );
  COND1XL U1780 ( .A(n1378), .B(n1452), .C(n1451), .Z(n586) );
  CNIVX1 U1781 ( .A(pushin), .Z(n1385) );
  CNR2X1 U1782 ( .A(n1225), .B(n2284), .Z(N406) );
  CNR3XL U1783 ( .A(n1984), .B(n1225), .C(n1224), .Z(N405) );
  CNR3XL U1784 ( .A(n1978), .B(n1225), .C(n1224), .Z(N399) );
  CNR3XL U1785 ( .A(n1979), .B(n1225), .C(n1224), .Z(N400) );
  CNR3XL U1786 ( .A(n1981), .B(n1225), .C(n1224), .Z(N402) );
  CNR3XL U1787 ( .A(n1980), .B(n1225), .C(n1224), .Z(N401) );
  CNR3XL U1788 ( .A(n1982), .B(n1225), .C(n1224), .Z(N403) );
  CNR3XL U1789 ( .A(n1983), .B(n1225), .C(n1224), .Z(N404) );
  COAN1X1 U1790 ( .A(n1305), .B(n1887), .C(n1886), .Z(n1149) );
  COAN1X1 U1791 ( .A(n1305), .B(n1885), .C(n1884), .Z(n1150) );
  COAN1X1 U1792 ( .A(n1305), .B(n1873), .C(n1872), .Z(n1151) );
  COAN1X1 U1793 ( .A(n1305), .B(n1875), .C(n1874), .Z(n1152) );
  COAN1X1 U1794 ( .A(n1305), .B(n1877), .C(n1876), .Z(n1153) );
  COAN1X1 U1795 ( .A(n1305), .B(n1879), .C(n1878), .Z(n1154) );
  COAN1X1 U1796 ( .A(n1305), .B(n1865), .C(n1864), .Z(n1155) );
  COAN1X1 U1797 ( .A(n1305), .B(n1867), .C(n1866), .Z(n1156) );
  COAN1X1 U1798 ( .A(n1305), .B(n1869), .C(n1868), .Z(n1157) );
  COAN1X1 U1799 ( .A(n1305), .B(n1871), .C(n1870), .Z(n1158) );
  COAN1X1 U1800 ( .A(n1304), .B(n1849), .C(n1848), .Z(n1159) );
  COAN1X1 U1801 ( .A(n1304), .B(n1847), .C(n1846), .Z(n1160) );
  COAN1X1 U1802 ( .A(n1304), .B(n1845), .C(n1844), .Z(n1161) );
  COAN1X1 U1803 ( .A(n1304), .B(n1843), .C(n1842), .Z(n1162) );
  COAN1X1 U1804 ( .A(n1304), .B(n1841), .C(n1840), .Z(n1163) );
  COAN1X1 U1805 ( .A(n1303), .B(n1839), .C(n1838), .Z(n1164) );
  COAN1X1 U1806 ( .A(n1303), .B(n1837), .C(n1836), .Z(n1165) );
  COAN1X1 U1807 ( .A(n1303), .B(n1835), .C(n1834), .Z(n1166) );
  COAN1X1 U1808 ( .A(n1304), .B(n1863), .C(n1862), .Z(n1167) );
  COAN1X1 U1809 ( .A(n1304), .B(n1861), .C(n1860), .Z(n1168) );
  COAN1X1 U1810 ( .A(n1304), .B(n1859), .C(n1858), .Z(n1169) );
  COAN1X1 U1811 ( .A(n1304), .B(n1853), .C(n1852), .Z(n1170) );
  COAN1X1 U1812 ( .A(n1304), .B(n1851), .C(n1850), .Z(n1171) );
  COAN1X1 U1813 ( .A(n1304), .B(n1857), .C(n1856), .Z(n1172) );
  COAN1X1 U1814 ( .A(n1304), .B(n1855), .C(n1854), .Z(n1173) );
  COAN1X1 U1815 ( .A(n1303), .B(n1833), .C(n1832), .Z(n1174) );
  COAN1X1 U1816 ( .A(n1303), .B(n1831), .C(n1830), .Z(n1175) );
  COAN1X1 U1817 ( .A(n1303), .B(n1829), .C(n1828), .Z(n1176) );
  COAN1X1 U1818 ( .A(n1303), .B(n1827), .C(n1826), .Z(n1177) );
  COAN1X1 U1819 ( .A(n1303), .B(n1825), .C(n1824), .Z(n1178) );
  COAN1X1 U1820 ( .A(n1303), .B(n1823), .C(n1822), .Z(n1179) );
  COAN1X1 U1821 ( .A(n1303), .B(n1821), .C(n1820), .Z(n1180) );
  COAN1X1 U1822 ( .A(n1303), .B(n1819), .C(n1818), .Z(n1181) );
  COAN1X1 U1823 ( .A(n1303), .B(n1817), .C(n1816), .Z(n1182) );
  COAN1X1 U1824 ( .A(n1302), .B(n1815), .C(n1814), .Z(n1183) );
  COAN1X1 U1825 ( .A(n1302), .B(n1813), .C(n1812), .Z(n1184) );
  COAN1X1 U1826 ( .A(n1302), .B(n1811), .C(n1810), .Z(n1185) );
  COAN1X1 U1827 ( .A(n1302), .B(n1809), .C(n1808), .Z(n1186) );
  COAN1X1 U1828 ( .A(n1302), .B(n1807), .C(n1806), .Z(n1187) );
  COAN1X1 U1829 ( .A(n1302), .B(n1805), .C(n1804), .Z(n1188) );
  COAN1X1 U1830 ( .A(n1302), .B(n1803), .C(n1802), .Z(n1189) );
  COAN1X1 U1831 ( .A(n1302), .B(n1801), .C(n1800), .Z(n1190) );
  COAN1X1 U1832 ( .A(n1302), .B(n1799), .C(n1798), .Z(n1191) );
  COAN1X1 U1833 ( .A(n1302), .B(n1797), .C(n1796), .Z(n1192) );
  COAN1X1 U1834 ( .A(n1302), .B(n1795), .C(n1794), .Z(n1193) );
  COAN1X1 U1835 ( .A(n1302), .B(n1793), .C(n1792), .Z(n1194) );
  COAN1X1 U1836 ( .A(n1301), .B(n1791), .C(n1790), .Z(n1195) );
  COAN1X1 U1837 ( .A(n1301), .B(n1789), .C(n1788), .Z(n1196) );
  COAN1X1 U1838 ( .A(n1301), .B(n1787), .C(n1786), .Z(n1197) );
  COAN1X1 U1839 ( .A(n1301), .B(n1785), .C(n1784), .Z(n1198) );
  COAN1X1 U1840 ( .A(n1301), .B(n1783), .C(n1782), .Z(n1199) );
  COAN1X1 U1841 ( .A(n1301), .B(n1781), .C(n1780), .Z(n1200) );
  COAN1X1 U1842 ( .A(n1301), .B(n1779), .C(n1778), .Z(n1201) );
  COAN1X1 U1843 ( .A(n1301), .B(n1777), .C(n1776), .Z(n1202) );
  COAN1X1 U1844 ( .A(n1301), .B(n1775), .C(n1774), .Z(n1203) );
  COAN1X1 U1845 ( .A(n1301), .B(n1773), .C(n1772), .Z(n1204) );
  CAN2X1 U1846 ( .A(n1506), .B(push0_stg2), .Z(n1205) );
  CAN2X1 U1847 ( .A(n12), .B(push0_stg2), .Z(n1206) );
  CAN2X1 U1848 ( .A(n1507), .B(push0_stg2), .Z(n1207) );
  CNIVX1 U1849 ( .A(h0_stg1[2]), .Z(n1213) );
  CNIVX1 U1850 ( .A(h0_stg1[2]), .Z(n1216) );
  CNIVX1 U1851 ( .A(h0_stg1[2]), .Z(n1215) );
  CNIVX1 U1852 ( .A(h0_stg1[2]), .Z(n1214) );
  CNIVX1 U1853 ( .A(h0_stg1[2]), .Z(n1217) );
  CNIVX1 U1854 ( .A(h0_stg1[4]), .Z(n1223) );
  CNIVX1 U1855 ( .A(h0_stg1[4]), .Z(n1222) );
  CNIVX1 U1856 ( .A(h0_stg1[4]), .Z(n1219) );
  CNIVX1 U1857 ( .A(h0_stg1[4]), .Z(n1221) );
  CNIVX1 U1858 ( .A(h0_stg1[4]), .Z(n1220) );
  CNIVX1 U1859 ( .A(h0_stg1[4]), .Z(n1218) );
  CNIVX1 U1860 ( .A(pushin), .Z(n1384) );
  CNIVX1 U1861 ( .A(pushin), .Z(n1383) );
  CNIVX1 U1862 ( .A(pushin), .Z(n1381) );
  CNIVX1 U1863 ( .A(pushin), .Z(n1382) );
  CNIVX1 U1864 ( .A(pushin), .Z(n1380) );
  CNR2X1 U1865 ( .A(cmd0_stg2[0]), .B(cmd0_stg2[1]), .Z(n12) );
  CNIVX1 U1866 ( .A(h0_stg1[5]), .Z(n1224) );
  CNIVX1 U1867 ( .A(h0_stg1[6]), .Z(n1225) );
  CIVXL U1868 ( .A(cmd1_en_stg2), .Z(n1263) );
  CNR3XL U1869 ( .A(n1977), .B(n1119), .C(n1121), .Z(cmd0_en_stg0) );
  CNR3XL U1870 ( .A(n1976), .B(n1119), .C(n1977), .Z(cmd1_en_stg0) );
  CMX2XL U1871 ( .A0(n1128), .A1(q[19]), .S(n1381), .Z(n677) );
  CMX2XL U1872 ( .A0(n1134), .A1(q[5]), .S(n1382), .Z(n663) );
  CMX2XL U1873 ( .A0(n1142), .A1(q[15]), .S(n1381), .Z(n673) );
  CMX2XL U1874 ( .A0(n1137), .A1(q[3]), .S(n1382), .Z(n661) );
  CMX2XL U1875 ( .A0(n793), .A1(q[23]), .S(n1380), .Z(n681) );
  CMX2XL U1876 ( .A0(n1130), .A1(q[7]), .S(n1382), .Z(n665) );
  CMX2XL U1877 ( .A0(n807), .A1(q[21]), .S(n1380), .Z(n679) );
  CMX2XL U1878 ( .A0(n1129), .A1(q[29]), .S(n1380), .Z(n687) );
  CMX2XL U1879 ( .A0(n1209), .A1(q[27]), .S(n1380), .Z(n685) );
  CMX2XL U1880 ( .A0(n1133), .A1(q[1]), .S(n1382), .Z(n659) );
  CMX2XL U1881 ( .A0(n1131), .A1(q[13]), .S(n1381), .Z(n671) );
  CIVX2 U1882 ( .A(n797), .Z(n1379) );
  CIVX1 U1883 ( .A(cmd0_en_stg2), .Z(n1227) );
  CIVX1 U1884 ( .A(cmd0_en_stg2), .Z(n1228) );
  CIVX1 U1885 ( .A(cmd0_en_stg2), .Z(n1229) );
  CIVX1 U1886 ( .A(cmd0_en_stg2), .Z(n1230) );
  CIVXL U1887 ( .A(n1226), .Z(n1231) );
  CIVXL U1888 ( .A(n1226), .Z(n1232) );
  CIVXL U1889 ( .A(n1226), .Z(n1233) );
  CIVXL U1890 ( .A(n1226), .Z(n1234) );
  CIVX1 U1891 ( .A(n1227), .Z(n1235) );
  CIVX1 U1892 ( .A(n1227), .Z(n1236) );
  CIVX1 U1893 ( .A(n1227), .Z(n1237) );
  CIVX1 U1894 ( .A(n1227), .Z(n1238) );
  CIVX1 U1895 ( .A(n1227), .Z(n1239) );
  CIVX1 U1896 ( .A(n1228), .Z(n1240) );
  CIVX1 U1897 ( .A(n1228), .Z(n1241) );
  CIVX1 U1898 ( .A(n1228), .Z(n1242) );
  CIVX1 U1899 ( .A(n1228), .Z(n1243) );
  CIVX1 U1900 ( .A(n1228), .Z(n1244) );
  CIVX1 U1901 ( .A(n1229), .Z(n1245) );
  CIVX1 U1902 ( .A(n1229), .Z(n1246) );
  CIVX1 U1903 ( .A(n1229), .Z(n1247) );
  CIVX1 U1904 ( .A(n1229), .Z(n1248) );
  CIVX1 U1905 ( .A(n1229), .Z(n1249) );
  CIVX1 U1906 ( .A(n1230), .Z(n1250) );
  CIVX1 U1907 ( .A(n1230), .Z(n1251) );
  CIVX1 U1908 ( .A(n1230), .Z(n1252) );
  CIVX1 U1909 ( .A(n1230), .Z(n1253) );
  CIVX1 U1910 ( .A(n1230), .Z(n1254) );
  CIVXL U1911 ( .A(n1226), .Z(n1255) );
  CIVX1 U1912 ( .A(n1230), .Z(n1256) );
  CIVX1 U1913 ( .A(n1226), .Z(n1257) );
  CIVX1 U1914 ( .A(n1226), .Z(n1258) );
  CIVX1 U1915 ( .A(n1226), .Z(n1259) );
  CIVXL U1916 ( .A(n1226), .Z(n1260) );
  CIVXL U1917 ( .A(n1226), .Z(n1261) );
  CIVXL U1918 ( .A(n1226), .Z(n1262) );
  CIVX1 U1919 ( .A(cmd1_en_stg2), .Z(n1264) );
  CIVX1 U1920 ( .A(cmd1_en_stg2), .Z(n1267) );
  CIVXL U1921 ( .A(n1263), .Z(n1269) );
  CIVXL U1922 ( .A(n1263), .Z(n1270) );
  CIVXL U1923 ( .A(n1263), .Z(n1271) );
  CIVXL U1924 ( .A(n1263), .Z(n1272) );
  CIVX1 U1925 ( .A(n1264), .Z(n1273) );
  CIVX1 U1926 ( .A(n1264), .Z(n1274) );
  CIVX1 U1927 ( .A(n1264), .Z(n1275) );
  CIVX1 U1928 ( .A(n1264), .Z(n1276) );
  CIVX1 U1929 ( .A(n1264), .Z(n1277) );
  CIVX1 U1930 ( .A(n1265), .Z(n1278) );
  CIVX1 U1931 ( .A(n1265), .Z(n1279) );
  CIVX1 U1932 ( .A(n1265), .Z(n1280) );
  CIVX1 U1933 ( .A(n1265), .Z(n1281) );
  CIVX1 U1934 ( .A(n1265), .Z(n1282) );
  CIVX1 U1935 ( .A(n1266), .Z(n1283) );
  CIVX1 U1936 ( .A(n1266), .Z(n1284) );
  CIVX1 U1937 ( .A(n1266), .Z(n1285) );
  CIVX1 U1938 ( .A(n1266), .Z(n1286) );
  CIVX1 U1939 ( .A(n1266), .Z(n1287) );
  CIVXL U1940 ( .A(n1267), .Z(n1290) );
  CIVX1 U1941 ( .A(n1268), .Z(n1291) );
  CIVX1 U1942 ( .A(n1268), .Z(n1292) );
  CIVXL U1943 ( .A(n1268), .Z(n1293) );
  CIVX1 U1944 ( .A(n1268), .Z(n1294) );
  CIVX1 U1945 ( .A(n1268), .Z(n1295) );
  CIVX1 U1946 ( .A(n1266), .Z(n1296) );
  CIVX1 U1947 ( .A(n1268), .Z(n1297) );
  CIVXL U1948 ( .A(n1265), .Z(n1298) );
  CIVXL U1949 ( .A(n1264), .Z(n1299) );
  CIVXL U1950 ( .A(n1363), .Z(n1362) );
  CIVX1 U1951 ( .A(h0_stg1[0]), .Z(n1363) );
  CIVXL U1952 ( .A(n1370), .Z(n1369) );
  CIVX2 U1953 ( .A(h0_stg1[1]), .Z(n1370) );
  CIVX2 U1954 ( .A(h0_stg1[3]), .Z(n1376) );
  CIVXL U1955 ( .A(n1107), .Z(n1377) );
  CMX2X1 U1956 ( .A0(q0[30]), .A1(q[30]), .S(n1380), .Z(n688) );
  CMX2X1 U1957 ( .A0(q0[28]), .A1(q[28]), .S(n1380), .Z(n686) );
  CMX2X1 U1958 ( .A0(q0[24]), .A1(q[24]), .S(n1380), .Z(n682) );
  CMX2X1 U1959 ( .A0(q0[20]), .A1(q[20]), .S(n1380), .Z(n678) );
  CMX2X1 U1960 ( .A0(n1208), .A1(q[14]), .S(n1381), .Z(n672) );
  CMX2X1 U1961 ( .A0(q0[12]), .A1(q[12]), .S(n1381), .Z(n670) );
  CMX2X1 U1962 ( .A0(q0[10]), .A1(q[10]), .S(n1381), .Z(n668) );
  CMX2X1 U1963 ( .A0(q0[4]), .A1(q[4]), .S(n1382), .Z(n662) );
  CMX2X1 U1964 ( .A0(q0[2]), .A1(q[2]), .S(n1382), .Z(n660) );
  CMX2X1 U1965 ( .A0(q0[0]), .A1(q[0]), .S(n1382), .Z(n658) );
  CMX2X1 U1966 ( .A0(h0[31]), .A1(h[31]), .S(n1382), .Z(n657) );
  CMX2X1 U1967 ( .A0(h0[29]), .A1(h[29]), .S(n1382), .Z(n655) );
  CMX2X1 U1968 ( .A0(n1138), .A1(h[28]), .S(n1382), .Z(n654) );
  CMX2X1 U1969 ( .A0(h0[27]), .A1(h[27]), .S(n1383), .Z(n653) );
  CMX2X1 U1970 ( .A0(n1140), .A1(h[26]), .S(n1383), .Z(n652) );
  CMX2X1 U1971 ( .A0(h0[24]), .A1(h[24]), .S(n1383), .Z(n650) );
  CMX2X1 U1972 ( .A0(h0[23]), .A1(h[23]), .S(n1383), .Z(n649) );
  CMX2X1 U1973 ( .A0(h0[20]), .A1(h[20]), .S(n1383), .Z(n646) );
  CMX2X1 U1974 ( .A0(h0[19]), .A1(h[19]), .S(n1383), .Z(n645) );
  CMX2X1 U1975 ( .A0(h0[16]), .A1(h[16]), .S(n1383), .Z(n642) );
  CMX2X1 U1976 ( .A0(n1132), .A1(h[15]), .S(n1384), .Z(n641) );
  CMX2X1 U1977 ( .A0(n1145), .A1(h[12]), .S(n1384), .Z(n638) );
  CMX2X1 U1978 ( .A0(n1144), .A1(h[10]), .S(n1384), .Z(n636) );
  CMX2X1 U1979 ( .A0(n1141), .A1(h[7]), .S(n1384), .Z(n633) );
  CMX2X1 U1980 ( .A0(n969), .A1(h[6]), .S(n1384), .Z(n632) );
  CMX2X1 U1981 ( .A0(n1105), .A1(h[5]), .S(n1384), .Z(n629) );
  CMX2X1 U1982 ( .A0(n1116), .A1(h[4]), .S(n1384), .Z(n626) );
  CMX2X1 U1983 ( .A0(n965), .A1(h[3]), .S(n1385), .Z(n623) );
  CMX2X1 U1984 ( .A0(n1143), .A1(h[2]), .S(n1385), .Z(n620) );
  CMX2X1 U1985 ( .A0(n1107), .A1(h[0]), .S(n1385), .Z(n614) );
  CMX2X1 U1986 ( .A0(cmd0_en_stg1), .A1(n1234), .S(rst), .Z(n755) );
  CMXI2X1 U1987 ( .A0(n1985), .A1(n797), .S(rst), .Z(n690) );
  CMX2X1 U1988 ( .A0(out2_stg2[63]), .A1(N406), .S(n798), .Z(n547) );
  CMX2X1 U1989 ( .A0(out2_stg2[62]), .A1(N405), .S(n798), .Z(n548) );
  CMX2X1 U1990 ( .A0(out2_stg2[61]), .A1(N404), .S(n798), .Z(n549) );
  CMX2X1 U1991 ( .A0(out2_stg2[60]), .A1(N403), .S(n798), .Z(n550) );
  CMX2X1 U1992 ( .A0(out2_stg2[59]), .A1(N402), .S(n798), .Z(n551) );
  CMX2X1 U1993 ( .A0(out2_stg2[58]), .A1(N401), .S(n798), .Z(n552) );
  CMX2X1 U1994 ( .A0(out2_stg2[57]), .A1(N400), .S(n798), .Z(n553) );
  CMX2X1 U1995 ( .A0(out2_stg2[56]), .A1(N399), .S(n798), .Z(n554) );
  CIVX2 U1996 ( .A(n1225), .Z(n1435) );
  CIVX2 U1997 ( .A(n1224), .Z(n1386) );
  CIVX2 U1998 ( .A(n2268), .Z(n1388) );
  CIVX2 U1999 ( .A(out2_stg2[55]), .Z(n1387) );
  COND2X1 U2000 ( .A(n1210), .B(n1388), .C(n798), .D(n1387), .Z(n555) );
  CIVX2 U2001 ( .A(n2267), .Z(n1390) );
  CIVX2 U2002 ( .A(out2_stg2[54]), .Z(n1389) );
  COND2X1 U2003 ( .A(n1210), .B(n1390), .C(n798), .D(n1389), .Z(n556) );
  CIVX2 U2004 ( .A(n2266), .Z(n1392) );
  CIVX2 U2005 ( .A(out2_stg2[53]), .Z(n1391) );
  COND2X1 U2006 ( .A(n1211), .B(n1392), .C(n798), .D(n1391), .Z(n557) );
  CIVX2 U2007 ( .A(n2265), .Z(n1394) );
  CIVX2 U2008 ( .A(out2_stg2[52]), .Z(n1393) );
  COND2X1 U2009 ( .A(n1211), .B(n1394), .C(n798), .D(n1393), .Z(n558) );
  CIVX2 U2010 ( .A(n2264), .Z(n1396) );
  CIVX2 U2011 ( .A(out2_stg2[51]), .Z(n1395) );
  COND2X1 U2012 ( .A(n1210), .B(n1396), .C(n798), .D(n1395), .Z(n559) );
  CIVX2 U2013 ( .A(n2263), .Z(n1398) );
  CIVX2 U2014 ( .A(out2_stg2[50]), .Z(n1397) );
  COND2X1 U2015 ( .A(n1210), .B(n1398), .C(n798), .D(n1397), .Z(n560) );
  CIVX2 U2016 ( .A(n2262), .Z(n1400) );
  CIVX2 U2017 ( .A(out2_stg2[49]), .Z(n1399) );
  COND2X1 U2018 ( .A(n1211), .B(n1400), .C(n1378), .D(n1399), .Z(n561) );
  CIVX2 U2019 ( .A(n2253), .Z(n1402) );
  CIVX2 U2020 ( .A(out2_stg2[48]), .Z(n1401) );
  COND2X1 U2021 ( .A(n1211), .B(n1402), .C(n1378), .D(n1401), .Z(n562) );
  CIVX2 U2022 ( .A(n2252), .Z(n1404) );
  CIVX2 U2023 ( .A(out2_stg2[47]), .Z(n1403) );
  COND2X1 U2024 ( .A(n1210), .B(n1404), .C(n1378), .D(n1403), .Z(n563) );
  CIVX2 U2025 ( .A(n2251), .Z(n1406) );
  CIVX2 U2026 ( .A(out2_stg2[46]), .Z(n1405) );
  COND2X1 U2027 ( .A(n1210), .B(n1406), .C(n1378), .D(n1405), .Z(n564) );
  CIVX2 U2028 ( .A(n2250), .Z(n1408) );
  CIVX2 U2029 ( .A(out2_stg2[45]), .Z(n1407) );
  COND2X1 U2030 ( .A(n1211), .B(n1408), .C(n1378), .D(n1407), .Z(n565) );
  CIVX2 U2031 ( .A(n2249), .Z(n1410) );
  CIVX2 U2032 ( .A(out2_stg2[44]), .Z(n1409) );
  COND2X1 U2033 ( .A(n1211), .B(n1410), .C(n1378), .D(n1409), .Z(n566) );
  CIVX2 U2034 ( .A(n2248), .Z(n1412) );
  CIVX2 U2035 ( .A(out2_stg2[43]), .Z(n1411) );
  COND2X1 U2036 ( .A(n1210), .B(n1412), .C(n1378), .D(n1411), .Z(n567) );
  CIVX2 U2037 ( .A(n2247), .Z(n1414) );
  CIVX2 U2038 ( .A(out2_stg2[42]), .Z(n1413) );
  COND2X1 U2039 ( .A(n1210), .B(n1414), .C(n1378), .D(n1413), .Z(n568) );
  CIVX2 U2040 ( .A(n2246), .Z(n1416) );
  CIVX2 U2041 ( .A(out2_stg2[41]), .Z(n1415) );
  COND2X1 U2042 ( .A(n1211), .B(n1416), .C(n1378), .D(n1415), .Z(n569) );
  CIVX2 U2043 ( .A(n2311), .Z(n1418) );
  CIVX2 U2044 ( .A(out2_stg2[40]), .Z(n1417) );
  COND2X1 U2045 ( .A(n1211), .B(n1418), .C(n1378), .D(n1417), .Z(n570) );
  CIVX2 U2046 ( .A(n2305), .Z(n1420) );
  CIVX2 U2047 ( .A(out2_stg2[39]), .Z(n1419) );
  COND2X1 U2048 ( .A(n1210), .B(n1420), .C(n1378), .D(n1419), .Z(n571) );
  CIVX2 U2049 ( .A(n2299), .Z(n1422) );
  CIVX2 U2050 ( .A(out2_stg2[38]), .Z(n1421) );
  COND2X1 U2051 ( .A(n1210), .B(n1422), .C(n1378), .D(n1421), .Z(n572) );
  CIVX2 U2052 ( .A(n2291), .Z(n1424) );
  CIVX2 U2053 ( .A(out2_stg2[37]), .Z(n1423) );
  COND2X1 U2054 ( .A(n1211), .B(n1424), .C(n1378), .D(n1423), .Z(n573) );
  CIVX2 U2055 ( .A(n2278), .Z(n1426) );
  CIVX2 U2056 ( .A(out2_stg2[36]), .Z(n1425) );
  COND2X1 U2057 ( .A(n1211), .B(n1426), .C(n1378), .D(n1425), .Z(n574) );
  CIVX2 U2058 ( .A(n2260), .Z(n1428) );
  CIVX2 U2059 ( .A(out2_stg2[35]), .Z(n1427) );
  COND2X1 U2060 ( .A(n1210), .B(n1428), .C(n1378), .D(n1427), .Z(n575) );
  CIVX2 U2061 ( .A(n2240), .Z(n1430) );
  CIVX2 U2062 ( .A(out2_stg2[34]), .Z(n1429) );
  COND2X1 U2063 ( .A(n1210), .B(n1430), .C(n1378), .D(n1429), .Z(n576) );
  CIVX2 U2064 ( .A(n2220), .Z(n1432) );
  CIVX2 U2065 ( .A(out2_stg2[33]), .Z(n1431) );
  COND2X1 U2066 ( .A(n1211), .B(n1432), .C(n1378), .D(n1431), .Z(n577) );
  CIVX2 U2067 ( .A(n2219), .Z(n1434) );
  CIVX2 U2068 ( .A(out2_stg2[32]), .Z(n1433) );
  COND2X1 U2069 ( .A(n1434), .B(n1211), .C(n1378), .D(n1433), .Z(n578) );
  CIVX2 U2070 ( .A(out2_stg2[31]), .Z(n1438) );
  CANR2X1 U2071 ( .A(n2283), .B(n1146), .C(n2216), .D(n1300), .Z(n1439) );
  CIVX2 U2072 ( .A(out2_stg2[29]), .Z(n1442) );
  CANR2X1 U2073 ( .A(n2282), .B(n1146), .C(n2212), .D(n1300), .Z(n1441) );
  CANR2X1 U2074 ( .A(n2281), .B(n1146), .C(n2196), .D(n1300), .Z(n1443) );
  CIVX2 U2075 ( .A(out2_stg2[27]), .Z(n1446) );
  CANR2X1 U2076 ( .A(n2280), .B(n1146), .C(n2192), .D(n1300), .Z(n1445) );
  CANR2X1 U2077 ( .A(n2271), .B(n1146), .C(n2188), .D(n1300), .Z(n1447) );
  CIVX2 U2078 ( .A(out2_stg2[25]), .Z(n1450) );
  CANR2X1 U2079 ( .A(n2270), .B(n1146), .C(n2184), .D(n1300), .Z(n1449) );
  CANR2X1 U2080 ( .A(n2269), .B(n1146), .C(n2180), .D(n1300), .Z(n1451) );
  CIVX2 U2081 ( .A(out2_stg2[23]), .Z(n1454) );
  CANR2X1 U2082 ( .A(n2268), .B(n1146), .C(n2174), .D(n1300), .Z(n1453) );
  CANR2X1 U2083 ( .A(n2267), .B(n1146), .C(n2167), .D(n1300), .Z(n1455) );
  CIVX2 U2084 ( .A(out2_stg2[21]), .Z(n1458) );
  CANR2X1 U2085 ( .A(n2266), .B(n1146), .C(n2160), .D(n1300), .Z(n1457) );
  CANR2X1 U2086 ( .A(n2265), .B(n1146), .C(n2153), .D(n1300), .Z(n1459) );
  CIVX2 U2087 ( .A(out2_stg2[19]), .Z(n1462) );
  CANR2X1 U2088 ( .A(n2264), .B(n1146), .C(n2146), .D(n1300), .Z(n1461) );
  CANR2X1 U2089 ( .A(n2263), .B(n1146), .C(n2129), .D(n1300), .Z(n1463) );
  CIVX2 U2090 ( .A(out2_stg2[17]), .Z(n1466) );
  CANR2X1 U2091 ( .A(n2262), .B(n1146), .C(n2122), .D(n1300), .Z(n1465) );
  CANR2X1 U2092 ( .A(n2253), .B(n1146), .C(n2115), .D(n1300), .Z(n1467) );
  CANR2X1 U2093 ( .A(n2252), .B(n1146), .C(n2102), .D(n1300), .Z(n1469) );
  CANR2X1 U2094 ( .A(n2251), .B(n1146), .C(n2097), .D(n1300), .Z(n1471) );
  CANR2X1 U2095 ( .A(n2250), .B(n1146), .C(n2082), .D(n1300), .Z(n1473) );
  CANR2X1 U2096 ( .A(n2249), .B(n1146), .C(n2067), .D(n1300), .Z(n1475) );
  CANR2X1 U2097 ( .A(n2248), .B(n1146), .C(n2039), .D(n1300), .Z(n1477) );
  CANR2X1 U2098 ( .A(n2247), .B(n1146), .C(n2023), .D(n1300), .Z(n1479) );
  CANR2X1 U2099 ( .A(n2246), .B(n1146), .C(n2021), .D(n1300), .Z(n1481) );
  CANR2X1 U2100 ( .A(n2311), .B(n1146), .C(n2312), .D(n1300), .Z(n1483) );
  CIVX2 U2101 ( .A(out2_stg2[7]), .Z(n1486) );
  CANR2X1 U2102 ( .A(n2305), .B(n1146), .C(n2306), .D(n1300), .Z(n1485) );
  CANR2X1 U2103 ( .A(n2299), .B(n1146), .C(n2300), .D(n1300), .Z(n1487) );
  CIVX2 U2104 ( .A(out2_stg2[5]), .Z(n1490) );
  CANR2X1 U2105 ( .A(n2291), .B(n1146), .C(n2292), .D(n1300), .Z(n1489) );
  CANR2X1 U2106 ( .A(n2278), .B(n1146), .C(n2279), .D(n1300), .Z(n1491) );
  CANR2X1 U2107 ( .A(n2260), .B(n1146), .C(n2261), .D(n1300), .Z(n1493) );
  CANR2X1 U2108 ( .A(n2240), .B(n1146), .C(n2241), .D(n1300), .Z(n1495) );
  CANR2X1 U2109 ( .A(n2220), .B(n1146), .C(n2208), .D(n1300), .Z(n1497) );
  CIVX2 U2110 ( .A(out2_stg2[0]), .Z(n1500) );
  CANR2X1 U2111 ( .A(n2219), .B(n1146), .C(n2139), .D(n1300), .Z(n1499) );
  CMX2X1 U2112 ( .A0(cmd1_en_stg1), .A1(n1297), .S(rst), .Z(n756) );
  CIVX2 U2113 ( .A(cmd1_en_stg2_d), .Z(n1765) );
  CND2X1 U2114 ( .A(n1290), .B(n1765), .Z(n1501) );
  CIVX2 U2115 ( .A(cmd0_en_stg2_d), .Z(n1767) );
  CND2X1 U2116 ( .A(n1762), .B(n1767), .Z(n1502) );
  CND2X1 U2117 ( .A(n1762), .B(cmd0_en_stg2_d), .Z(n1503) );
  CMX2X1 U2118 ( .A0(out1_stg2[62]), .A1(N271), .S(n1269), .Z(n421) );
  CIVX2 U2119 ( .A(cmd0_stg2[0]), .Z(n1975) );
  CND2X1 U2120 ( .A(cmd0_stg2[1]), .B(n1975), .Z(n1917) );
  CIVX2 U2121 ( .A(n1917), .Z(n1506) );
  CANR2X1 U2122 ( .A(n1206), .B(out0_stg2[62]), .C(N480), .D(n1205), .Z(n1509)
         );
  CIVX2 U2123 ( .A(cmd0_stg2[1]), .Z(n1974) );
  CND2X1 U2124 ( .A(cmd0_stg2[0]), .B(n1974), .Z(n1916) );
  CIVX2 U2125 ( .A(n1916), .Z(n1507) );
  CANR2X1 U2126 ( .A(n1207), .B(out1_stg2[62]), .C(acc[62]), .D(n802), .Z(
        n1508) );
  CND2X1 U2127 ( .A(n1509), .B(n1508), .Z(n420) );
  CMX2X1 U2128 ( .A0(out1_stg2[61]), .A1(N270), .S(n1270), .Z(n423) );
  CANR2X1 U2129 ( .A(n1206), .B(out0_stg2[61]), .C(N479), .D(n1205), .Z(n1513)
         );
  CANR2X1 U2130 ( .A(n1207), .B(out1_stg2[61]), .C(acc[61]), .D(n802), .Z(
        n1512) );
  CND2X1 U2131 ( .A(n1513), .B(n1512), .Z(n422) );
  CMX2X1 U2132 ( .A0(out1_stg2[60]), .A1(N269), .S(n1271), .Z(n425) );
  CANR2X1 U2133 ( .A(n1206), .B(out0_stg2[60]), .C(N478), .D(n1205), .Z(n1517)
         );
  CANR2X1 U2134 ( .A(n1207), .B(out1_stg2[60]), .C(acc[60]), .D(n802), .Z(
        n1516) );
  CND2X1 U2135 ( .A(n1517), .B(n1516), .Z(n424) );
  CMX2X1 U2136 ( .A0(out1_stg2[59]), .A1(N268), .S(n1272), .Z(n427) );
  CANR2X1 U2137 ( .A(n1206), .B(out0_stg2[59]), .C(N477), .D(n1205), .Z(n1521)
         );
  CANR2X1 U2138 ( .A(n1207), .B(out1_stg2[59]), .C(acc[59]), .D(n802), .Z(
        n1520) );
  CND2X1 U2139 ( .A(n1521), .B(n1520), .Z(n426) );
  CMX2X1 U2140 ( .A0(out1_stg2[58]), .A1(N267), .S(n1273), .Z(n429) );
  CANR2X1 U2141 ( .A(n1206), .B(out0_stg2[58]), .C(N476), .D(n1205), .Z(n1525)
         );
  CANR2X1 U2142 ( .A(n1207), .B(out1_stg2[58]), .C(acc[58]), .D(n802), .Z(
        n1524) );
  CND2X1 U2143 ( .A(n1525), .B(n1524), .Z(n428) );
  CMX2X1 U2144 ( .A0(out1_stg2[57]), .A1(N266), .S(n1274), .Z(n431) );
  CANR2X1 U2145 ( .A(n1206), .B(out0_stg2[57]), .C(N475), .D(n1205), .Z(n1529)
         );
  CANR2X1 U2146 ( .A(n1207), .B(out1_stg2[57]), .C(acc[57]), .D(n802), .Z(
        n1528) );
  CND2X1 U2147 ( .A(n1529), .B(n1528), .Z(n430) );
  CMX2X1 U2148 ( .A0(out1_stg2[56]), .A1(N265), .S(n1275), .Z(n433) );
  CANR2X1 U2149 ( .A(n1206), .B(out0_stg2[56]), .C(N474), .D(n1205), .Z(n1533)
         );
  CANR2X1 U2150 ( .A(n1207), .B(out1_stg2[56]), .C(acc[56]), .D(n802), .Z(
        n1532) );
  CND2X1 U2151 ( .A(n1533), .B(n1532), .Z(n432) );
  CMX2X1 U2152 ( .A0(out1_stg2[55]), .A1(N264), .S(n1276), .Z(n435) );
  CANR2X1 U2153 ( .A(n1206), .B(out0_stg2[55]), .C(N473), .D(n1205), .Z(n1537)
         );
  CANR2X1 U2154 ( .A(n1207), .B(out1_stg2[55]), .C(acc[55]), .D(n802), .Z(
        n1536) );
  CND2X1 U2155 ( .A(n1537), .B(n1536), .Z(n434) );
  CMX2X1 U2156 ( .A0(out1_stg2[54]), .A1(N263), .S(n1277), .Z(n437) );
  CANR2X1 U2157 ( .A(n1206), .B(out0_stg2[54]), .C(N472), .D(n1205), .Z(n1541)
         );
  CANR2X1 U2158 ( .A(n1207), .B(out1_stg2[54]), .C(acc[54]), .D(n802), .Z(
        n1540) );
  CND2X1 U2159 ( .A(n1541), .B(n1540), .Z(n436) );
  CMX2X1 U2160 ( .A0(out1_stg2[53]), .A1(N262), .S(n1278), .Z(n439) );
  CANR2X1 U2161 ( .A(n1206), .B(out0_stg2[53]), .C(N471), .D(n1205), .Z(n1545)
         );
  CANR2X1 U2162 ( .A(n1207), .B(out1_stg2[53]), .C(acc[53]), .D(n802), .Z(
        n1544) );
  CND2X1 U2163 ( .A(n1545), .B(n1544), .Z(n438) );
  CMX2X1 U2164 ( .A0(out1_stg2[52]), .A1(N261), .S(n1279), .Z(n441) );
  CANR2X1 U2165 ( .A(n1206), .B(out0_stg2[52]), .C(N470), .D(n1205), .Z(n1549)
         );
  CANR2X1 U2166 ( .A(n1207), .B(out1_stg2[52]), .C(acc[52]), .D(n802), .Z(
        n1548) );
  CND2X1 U2167 ( .A(n1549), .B(n1548), .Z(n440) );
  CMX2X1 U2168 ( .A0(out1_stg2[51]), .A1(N260), .S(n1280), .Z(n443) );
  CANR2X1 U2169 ( .A(n1206), .B(out0_stg2[51]), .C(N469), .D(n1205), .Z(n1553)
         );
  CANR2X1 U2170 ( .A(n1207), .B(out1_stg2[51]), .C(acc[51]), .D(n802), .Z(
        n1552) );
  CND2X1 U2171 ( .A(n1553), .B(n1552), .Z(n442) );
  CMX2X1 U2172 ( .A0(out1_stg2[50]), .A1(N259), .S(n1281), .Z(n445) );
  CANR2X1 U2173 ( .A(n1206), .B(out0_stg2[50]), .C(N468), .D(n1205), .Z(n1557)
         );
  CANR2X1 U2174 ( .A(n1207), .B(out1_stg2[50]), .C(acc[50]), .D(n802), .Z(
        n1556) );
  CND2X1 U2175 ( .A(n1557), .B(n1556), .Z(n444) );
  CMX2X1 U2176 ( .A0(out1_stg2[49]), .A1(N258), .S(n1282), .Z(n447) );
  CANR2X1 U2177 ( .A(n1206), .B(out0_stg2[49]), .C(N467), .D(n1205), .Z(n1561)
         );
  CANR2X1 U2178 ( .A(n1207), .B(out1_stg2[49]), .C(acc[49]), .D(n802), .Z(
        n1560) );
  CND2X1 U2179 ( .A(n1561), .B(n1560), .Z(n446) );
  CMX2X1 U2180 ( .A0(out1_stg2[48]), .A1(N257), .S(n1283), .Z(n449) );
  CANR2X1 U2181 ( .A(n1206), .B(out0_stg2[48]), .C(N466), .D(n1205), .Z(n1565)
         );
  CANR2X1 U2182 ( .A(n1207), .B(out1_stg2[48]), .C(acc[48]), .D(n802), .Z(
        n1564) );
  CND2X1 U2183 ( .A(n1565), .B(n1564), .Z(n448) );
  CMX2X1 U2184 ( .A0(out1_stg2[47]), .A1(N256), .S(n1284), .Z(n451) );
  CANR2X1 U2185 ( .A(n1206), .B(out0_stg2[47]), .C(N465), .D(n1205), .Z(n1569)
         );
  CANR2X1 U2186 ( .A(n1207), .B(out1_stg2[47]), .C(acc[47]), .D(n802), .Z(
        n1568) );
  CND2X1 U2187 ( .A(n1569), .B(n1568), .Z(n450) );
  CMX2X1 U2188 ( .A0(out1_stg2[46]), .A1(N255), .S(n1285), .Z(n453) );
  CANR2X1 U2189 ( .A(n1206), .B(out0_stg2[46]), .C(N464), .D(n1205), .Z(n1573)
         );
  CANR2X1 U2190 ( .A(n1207), .B(out1_stg2[46]), .C(acc[46]), .D(n802), .Z(
        n1572) );
  CND2X1 U2191 ( .A(n1573), .B(n1572), .Z(n452) );
  CMX2X1 U2192 ( .A0(out1_stg2[45]), .A1(N254), .S(n1286), .Z(n455) );
  CANR2X1 U2193 ( .A(n1206), .B(out0_stg2[45]), .C(N463), .D(n1205), .Z(n1577)
         );
  CANR2X1 U2194 ( .A(n1207), .B(out1_stg2[45]), .C(acc[45]), .D(n802), .Z(
        n1576) );
  CND2X1 U2195 ( .A(n1577), .B(n1576), .Z(n454) );
  CMX2X1 U2196 ( .A0(out1_stg2[44]), .A1(N253), .S(n1287), .Z(n457) );
  CANR2X1 U2197 ( .A(n1206), .B(out0_stg2[44]), .C(N462), .D(n1205), .Z(n1581)
         );
  CANR2X1 U2198 ( .A(n1207), .B(out1_stg2[44]), .C(acc[44]), .D(n802), .Z(
        n1580) );
  CND2X1 U2199 ( .A(n1581), .B(n1580), .Z(n456) );
  CMX2X1 U2200 ( .A0(out1_stg2[43]), .A1(N252), .S(n1295), .Z(n459) );
  CANR2X1 U2201 ( .A(n1206), .B(out0_stg2[43]), .C(N461), .D(n1205), .Z(n1585)
         );
  CANR2X1 U2202 ( .A(n1207), .B(out1_stg2[43]), .C(acc[43]), .D(n802), .Z(
        n1584) );
  CND2X1 U2203 ( .A(n1585), .B(n1584), .Z(n458) );
  CMX2X1 U2204 ( .A0(out1_stg2[42]), .A1(N251), .S(n1288), .Z(n461) );
  CANR2X1 U2205 ( .A(n1206), .B(out0_stg2[42]), .C(N460), .D(n1205), .Z(n1589)
         );
  CANR2X1 U2206 ( .A(n1207), .B(out1_stg2[42]), .C(acc[42]), .D(n802), .Z(
        n1588) );
  CND2X1 U2207 ( .A(n1589), .B(n1588), .Z(n460) );
  CMX2X1 U2208 ( .A0(out1_stg2[41]), .A1(N250), .S(n1289), .Z(n463) );
  CANR2X1 U2209 ( .A(n1206), .B(out0_stg2[41]), .C(N459), .D(n1205), .Z(n1593)
         );
  CANR2X1 U2210 ( .A(n1207), .B(out1_stg2[41]), .C(acc[41]), .D(n802), .Z(
        n1592) );
  CND2X1 U2211 ( .A(n1593), .B(n1592), .Z(n462) );
  CMX2X1 U2212 ( .A0(out1_stg2[40]), .A1(N249), .S(n1289), .Z(n465) );
  CANR2X1 U2213 ( .A(n1206), .B(out0_stg2[40]), .C(N458), .D(n1205), .Z(n1597)
         );
  CANR2X1 U2214 ( .A(n1207), .B(out1_stg2[40]), .C(acc[40]), .D(n802), .Z(
        n1596) );
  CND2X1 U2215 ( .A(n1597), .B(n1596), .Z(n464) );
  CMX2X1 U2216 ( .A0(out1_stg2[39]), .A1(N248), .S(n1290), .Z(n467) );
  CANR2X1 U2217 ( .A(n1206), .B(out0_stg2[39]), .C(N457), .D(n1205), .Z(n1601)
         );
  CANR2X1 U2218 ( .A(n1207), .B(out1_stg2[39]), .C(acc[39]), .D(n802), .Z(
        n1600) );
  CND2X1 U2219 ( .A(n1601), .B(n1600), .Z(n466) );
  CMX2X1 U2220 ( .A0(out1_stg2[38]), .A1(N247), .S(n1291), .Z(n469) );
  CANR2X1 U2221 ( .A(n1206), .B(out0_stg2[38]), .C(N456), .D(n1205), .Z(n1605)
         );
  CANR2X1 U2222 ( .A(n1207), .B(out1_stg2[38]), .C(acc[38]), .D(n802), .Z(
        n1604) );
  CND2X1 U2223 ( .A(n1605), .B(n1604), .Z(n468) );
  CMX2X1 U2224 ( .A0(out1_stg2[37]), .A1(N246), .S(n1292), .Z(n471) );
  CANR2X1 U2225 ( .A(n1206), .B(out0_stg2[37]), .C(N455), .D(n1205), .Z(n1609)
         );
  CANR2X1 U2226 ( .A(n1207), .B(out1_stg2[37]), .C(acc[37]), .D(n802), .Z(
        n1608) );
  CND2X1 U2227 ( .A(n1609), .B(n1608), .Z(n470) );
  CMX2X1 U2228 ( .A0(out1_stg2[36]), .A1(N245), .S(n1293), .Z(n473) );
  CANR2X1 U2229 ( .A(n1206), .B(out0_stg2[36]), .C(N454), .D(n1205), .Z(n1613)
         );
  CANR2X1 U2230 ( .A(n1207), .B(out1_stg2[36]), .C(acc[36]), .D(n802), .Z(
        n1612) );
  CND2X1 U2231 ( .A(n1613), .B(n1612), .Z(n472) );
  CMX2X1 U2232 ( .A0(out1_stg2[35]), .A1(N244), .S(n1294), .Z(n475) );
  CANR2X1 U2233 ( .A(n1206), .B(out0_stg2[35]), .C(N453), .D(n1205), .Z(n1617)
         );
  CANR2X1 U2234 ( .A(n1207), .B(out1_stg2[35]), .C(acc[35]), .D(n802), .Z(
        n1616) );
  CND2X1 U2235 ( .A(n1617), .B(n1616), .Z(n474) );
  CMX2X1 U2236 ( .A0(out1_stg2[34]), .A1(N243), .S(n1295), .Z(n477) );
  CANR2X1 U2237 ( .A(n1206), .B(out0_stg2[34]), .C(N452), .D(n1205), .Z(n1621)
         );
  CANR2X1 U2238 ( .A(n1207), .B(out1_stg2[34]), .C(acc[34]), .D(n802), .Z(
        n1620) );
  CND2X1 U2239 ( .A(n1621), .B(n1620), .Z(n476) );
  CMX2X1 U2240 ( .A0(out1_stg2[33]), .A1(N242), .S(n1295), .Z(n479) );
  CANR2X1 U2241 ( .A(n1206), .B(out0_stg2[33]), .C(N451), .D(n1205), .Z(n1625)
         );
  CANR2X1 U2242 ( .A(n1207), .B(out1_stg2[33]), .C(acc[33]), .D(n802), .Z(
        n1624) );
  CND2X1 U2243 ( .A(n1625), .B(n1624), .Z(n478) );
  CMX2X1 U2244 ( .A0(out1_stg2[32]), .A1(N241), .S(n1296), .Z(n481) );
  CANR2X1 U2245 ( .A(n1206), .B(out0_stg2[32]), .C(N450), .D(n1205), .Z(n1629)
         );
  CANR2X1 U2246 ( .A(n1207), .B(out1_stg2[32]), .C(acc[32]), .D(n802), .Z(
        n1628) );
  CND2X1 U2247 ( .A(n1629), .B(n1628), .Z(n480) );
  CMX2X1 U2248 ( .A0(out1_stg2[31]), .A1(N240), .S(n1297), .Z(n483) );
  CANR2X1 U2249 ( .A(n1206), .B(out0_stg2[31]), .C(N449), .D(n1205), .Z(n1633)
         );
  CANR2X1 U2250 ( .A(n1207), .B(out1_stg2[31]), .C(acc[31]), .D(n802), .Z(
        n1632) );
  CND2X1 U2251 ( .A(n1633), .B(n1632), .Z(n482) );
  CMX2X1 U2252 ( .A0(out1_stg2[30]), .A1(N239), .S(n1292), .Z(n485) );
  CANR2X1 U2253 ( .A(n1206), .B(out0_stg2[30]), .C(N448), .D(n1205), .Z(n1637)
         );
  CANR2X1 U2254 ( .A(n1207), .B(out1_stg2[30]), .C(acc[30]), .D(n802), .Z(
        n1636) );
  CND2X1 U2255 ( .A(n1637), .B(n1636), .Z(n484) );
  CMX2X1 U2256 ( .A0(out1_stg2[29]), .A1(N238), .S(n1294), .Z(n487) );
  CANR2X1 U2257 ( .A(n1206), .B(out0_stg2[29]), .C(N447), .D(n1205), .Z(n1641)
         );
  CANR2X1 U2258 ( .A(n1207), .B(out1_stg2[29]), .C(acc[29]), .D(n802), .Z(
        n1640) );
  CND2X1 U2259 ( .A(n1641), .B(n1640), .Z(n486) );
  CMX2X1 U2260 ( .A0(out1_stg2[28]), .A1(N237), .S(n1291), .Z(n489) );
  CANR2X1 U2261 ( .A(n1206), .B(out0_stg2[28]), .C(N446), .D(n1205), .Z(n1645)
         );
  CANR2X1 U2262 ( .A(n1207), .B(out1_stg2[28]), .C(acc[28]), .D(n802), .Z(
        n1644) );
  CND2X1 U2263 ( .A(n1645), .B(n1644), .Z(n488) );
  CMX2X1 U2264 ( .A0(out1_stg2[27]), .A1(N236), .S(n1296), .Z(n491) );
  CANR2X1 U2265 ( .A(n1206), .B(out0_stg2[27]), .C(N445), .D(n1205), .Z(n1649)
         );
  CANR2X1 U2266 ( .A(n1207), .B(out1_stg2[27]), .C(acc[27]), .D(n802), .Z(
        n1648) );
  CND2X1 U2267 ( .A(n1649), .B(n1648), .Z(n490) );
  CMX2X1 U2268 ( .A0(out1_stg2[26]), .A1(N235), .S(n1297), .Z(n493) );
  CANR2X1 U2269 ( .A(n1206), .B(out0_stg2[26]), .C(N444), .D(n1205), .Z(n1653)
         );
  CANR2X1 U2270 ( .A(n1207), .B(out1_stg2[26]), .C(acc[26]), .D(n802), .Z(
        n1652) );
  CND2X1 U2271 ( .A(n1653), .B(n1652), .Z(n492) );
  CMX2X1 U2272 ( .A0(out1_stg2[25]), .A1(N234), .S(n1298), .Z(n495) );
  CANR2X1 U2273 ( .A(n1206), .B(out0_stg2[25]), .C(N443), .D(n1205), .Z(n1657)
         );
  CANR2X1 U2274 ( .A(n1207), .B(out1_stg2[25]), .C(acc[25]), .D(n802), .Z(
        n1656) );
  CND2X1 U2275 ( .A(n1657), .B(n1656), .Z(n494) );
  CMX2X1 U2276 ( .A0(out1_stg2[24]), .A1(N233), .S(n1299), .Z(n497) );
  CANR2X1 U2277 ( .A(n1206), .B(out0_stg2[24]), .C(N442), .D(n1205), .Z(n1661)
         );
  CANR2X1 U2278 ( .A(n1207), .B(out1_stg2[24]), .C(acc[24]), .D(n802), .Z(
        n1660) );
  CND2X1 U2279 ( .A(n1661), .B(n1660), .Z(n496) );
  CMX2X1 U2280 ( .A0(out1_stg2[23]), .A1(N232), .S(n1274), .Z(n499) );
  CANR2X1 U2281 ( .A(n1206), .B(out0_stg2[23]), .C(N441), .D(n1205), .Z(n1665)
         );
  CANR2X1 U2282 ( .A(n1207), .B(out1_stg2[23]), .C(acc[23]), .D(n802), .Z(
        n1664) );
  CND2X1 U2283 ( .A(n1665), .B(n1664), .Z(n498) );
  CMX2X1 U2284 ( .A0(out1_stg2[22]), .A1(N231), .S(n1296), .Z(n501) );
  CANR2X1 U2285 ( .A(n1206), .B(out0_stg2[22]), .C(N440), .D(n1205), .Z(n1669)
         );
  CANR2X1 U2286 ( .A(n1207), .B(out1_stg2[22]), .C(acc[22]), .D(n802), .Z(
        n1668) );
  CND2X1 U2287 ( .A(n1669), .B(n1668), .Z(n500) );
  CMX2X1 U2288 ( .A0(out1_stg2[21]), .A1(N230), .S(n1269), .Z(n503) );
  CANR2X1 U2289 ( .A(n1206), .B(out0_stg2[21]), .C(N439), .D(n1205), .Z(n1673)
         );
  CANR2X1 U2290 ( .A(n1207), .B(out1_stg2[21]), .C(acc[21]), .D(n802), .Z(
        n1672) );
  CND2X1 U2291 ( .A(n1673), .B(n1672), .Z(n502) );
  CMX2X1 U2292 ( .A0(out1_stg2[20]), .A1(N229), .S(n1270), .Z(n505) );
  CANR2X1 U2293 ( .A(n1206), .B(out0_stg2[20]), .C(N438), .D(n1205), .Z(n1677)
         );
  CANR2X1 U2294 ( .A(n1207), .B(out1_stg2[20]), .C(acc[20]), .D(n802), .Z(
        n1676) );
  CND2X1 U2295 ( .A(n1677), .B(n1676), .Z(n504) );
  CMX2X1 U2296 ( .A0(out1_stg2[19]), .A1(N228), .S(n1271), .Z(n507) );
  CANR2X1 U2297 ( .A(n1206), .B(out0_stg2[19]), .C(N437), .D(n1205), .Z(n1681)
         );
  CANR2X1 U2298 ( .A(n1207), .B(out1_stg2[19]), .C(acc[19]), .D(n802), .Z(
        n1680) );
  CND2X1 U2299 ( .A(n1681), .B(n1680), .Z(n506) );
  CMX2X1 U2300 ( .A0(out1_stg2[18]), .A1(N227), .S(n1272), .Z(n509) );
  CANR2X1 U2301 ( .A(n1206), .B(out0_stg2[18]), .C(N436), .D(n1205), .Z(n1685)
         );
  CANR2X1 U2302 ( .A(n1207), .B(out1_stg2[18]), .C(acc[18]), .D(n802), .Z(
        n1684) );
  CND2X1 U2303 ( .A(n1685), .B(n1684), .Z(n508) );
  CMX2X1 U2304 ( .A0(out1_stg2[17]), .A1(N226), .S(n1273), .Z(n511) );
  CANR2X1 U2305 ( .A(n1206), .B(out0_stg2[17]), .C(N435), .D(n1205), .Z(n1689)
         );
  CANR2X1 U2306 ( .A(n1207), .B(out1_stg2[17]), .C(acc[17]), .D(n802), .Z(
        n1688) );
  CND2X1 U2307 ( .A(n1689), .B(n1688), .Z(n510) );
  CMX2X1 U2308 ( .A0(out1_stg2[16]), .A1(N225), .S(n1274), .Z(n513) );
  CANR2X1 U2309 ( .A(n1206), .B(out0_stg2[16]), .C(N434), .D(n1205), .Z(n1693)
         );
  CANR2X1 U2310 ( .A(n1207), .B(out1_stg2[16]), .C(acc[16]), .D(n802), .Z(
        n1692) );
  CND2X1 U2311 ( .A(n1693), .B(n1692), .Z(n512) );
  CIVX2 U2312 ( .A(out1_stg2[16]), .Z(n1695) );
  CMX2X1 U2313 ( .A0(out1_stg2[15]), .A1(N224), .S(n1275), .Z(n515) );
  CANR2X1 U2314 ( .A(n1206), .B(out0_stg2[15]), .C(N433), .D(n1205), .Z(n1697)
         );
  CANR2X1 U2315 ( .A(n1207), .B(out1_stg2[15]), .C(acc[15]), .D(n802), .Z(
        n1696) );
  CND2X1 U2316 ( .A(n1697), .B(n1696), .Z(n514) );
  CMX2X1 U2317 ( .A0(out1_stg2[14]), .A1(N223), .S(n1276), .Z(n517) );
  CANR2X1 U2318 ( .A(n1206), .B(out0_stg2[14]), .C(N432), .D(n1205), .Z(n1701)
         );
  CANR2X1 U2319 ( .A(n1207), .B(out1_stg2[14]), .C(acc[14]), .D(n802), .Z(
        n1700) );
  CND2X1 U2320 ( .A(n1701), .B(n1700), .Z(n516) );
  CMX2X1 U2321 ( .A0(out1_stg2[13]), .A1(N222), .S(n1277), .Z(n519) );
  CANR2X1 U2322 ( .A(n1206), .B(out0_stg2[13]), .C(N431), .D(n1205), .Z(n1705)
         );
  CANR2X1 U2323 ( .A(n1207), .B(out1_stg2[13]), .C(acc[13]), .D(n802), .Z(
        n1704) );
  CND2X1 U2324 ( .A(n1705), .B(n1704), .Z(n518) );
  CMX2X1 U2325 ( .A0(out1_stg2[12]), .A1(N221), .S(n1278), .Z(n521) );
  CANR2X1 U2326 ( .A(n1206), .B(out0_stg2[12]), .C(N430), .D(n1205), .Z(n1709)
         );
  CANR2X1 U2327 ( .A(n1207), .B(out1_stg2[12]), .C(acc[12]), .D(n802), .Z(
        n1708) );
  CND2X1 U2328 ( .A(n1709), .B(n1708), .Z(n520) );
  CMX2X1 U2329 ( .A0(out1_stg2[11]), .A1(N220), .S(n1279), .Z(n523) );
  CANR2X1 U2330 ( .A(n1207), .B(out1_stg2[11]), .C(acc[11]), .D(n802), .Z(
        n1712) );
  CND2X1 U2331 ( .A(n1713), .B(n1712), .Z(n522) );
  CMX2X1 U2332 ( .A0(out1_stg2[10]), .A1(N219), .S(n1280), .Z(n525) );
  CANR2X1 U2333 ( .A(n1206), .B(out0_stg2[10]), .C(N428), .D(n1205), .Z(n1717)
         );
  CANR2X1 U2334 ( .A(n1207), .B(out1_stg2[10]), .C(acc[10]), .D(n802), .Z(
        n1716) );
  CND2X1 U2335 ( .A(n1717), .B(n1716), .Z(n524) );
  CMX2X1 U2336 ( .A0(out1_stg2[9]), .A1(N218), .S(n1281), .Z(n527) );
  CANR2X1 U2337 ( .A(n1207), .B(out1_stg2[9]), .C(acc[9]), .D(n802), .Z(n1720)
         );
  CND2X1 U2338 ( .A(n1721), .B(n1720), .Z(n526) );
  CIVX2 U2339 ( .A(out1_stg2[9]), .Z(n1723) );
  CANR2X1 U2340 ( .A(n1759), .B(acc[9]), .C(n1758), .D(out0_stg2[9]), .Z(n1722) );
  CMX2X1 U2341 ( .A0(out1_stg2[8]), .A1(N217), .S(n1282), .Z(n529) );
  CANR2X1 U2342 ( .A(n1206), .B(out0_stg2[8]), .C(N426), .D(n1205), .Z(n1725)
         );
  CANR2X1 U2343 ( .A(n1207), .B(out1_stg2[8]), .C(acc[8]), .D(n802), .Z(n1724)
         );
  CND2X1 U2344 ( .A(n1725), .B(n1724), .Z(n528) );
  CIVX2 U2345 ( .A(out1_stg2[8]), .Z(n1727) );
  CMX2X1 U2346 ( .A0(out1_stg2[7]), .A1(N216), .S(n1283), .Z(n531) );
  CANR2X1 U2347 ( .A(n1206), .B(out0_stg2[7]), .C(N425), .D(n1205), .Z(n1729)
         );
  CANR2X1 U2348 ( .A(n1207), .B(out1_stg2[7]), .C(acc[7]), .D(n802), .Z(n1728)
         );
  CND2X1 U2349 ( .A(n1729), .B(n1728), .Z(n530) );
  CIVX2 U2350 ( .A(out1_stg2[7]), .Z(n1731) );
  CMX2X1 U2351 ( .A0(out1_stg2[6]), .A1(N215), .S(n1284), .Z(n533) );
  CANR2X1 U2352 ( .A(n1206), .B(out0_stg2[6]), .C(N424), .D(n1205), .Z(n1733)
         );
  CANR2X1 U2353 ( .A(n1207), .B(out1_stg2[6]), .C(acc[6]), .D(n802), .Z(n1732)
         );
  CND2X1 U2354 ( .A(n1733), .B(n1732), .Z(n532) );
  CIVX2 U2355 ( .A(out1_stg2[6]), .Z(n1735) );
  CMX2X1 U2356 ( .A0(out1_stg2[5]), .A1(N214), .S(n1285), .Z(n535) );
  CANR2X1 U2357 ( .A(n1206), .B(out0_stg2[5]), .C(N423), .D(n1205), .Z(n1737)
         );
  CANR2X1 U2358 ( .A(n1207), .B(out1_stg2[5]), .C(acc[5]), .D(n802), .Z(n1736)
         );
  CND2X1 U2359 ( .A(n1737), .B(n1736), .Z(n534) );
  CIVX2 U2360 ( .A(out1_stg2[5]), .Z(n1739) );
  CMX2X1 U2361 ( .A0(out1_stg2[4]), .A1(N213), .S(n1286), .Z(n537) );
  CANR2X1 U2362 ( .A(n1206), .B(out0_stg2[4]), .C(N422), .D(n1205), .Z(n1741)
         );
  CANR2X1 U2363 ( .A(n1207), .B(out1_stg2[4]), .C(acc[4]), .D(n802), .Z(n1740)
         );
  CND2X1 U2364 ( .A(n1741), .B(n1740), .Z(n536) );
  CIVX2 U2365 ( .A(out1_stg2[4]), .Z(n1743) );
  CMX2X1 U2366 ( .A0(out1_stg2[3]), .A1(N212), .S(n1287), .Z(n539) );
  CANR2X1 U2367 ( .A(n1207), .B(out1_stg2[3]), .C(acc[3]), .D(n802), .Z(n1744)
         );
  CND2X1 U2368 ( .A(n1745), .B(n1744), .Z(n538) );
  CIVX2 U2369 ( .A(out1_stg2[3]), .Z(n1747) );
  CMX2X1 U2370 ( .A0(out1_stg2[2]), .A1(N211), .S(n1297), .Z(n541) );
  CANR2X1 U2371 ( .A(n1206), .B(out0_stg2[2]), .C(N420), .D(n1205), .Z(n1749)
         );
  CANR2X1 U2372 ( .A(n1207), .B(out1_stg2[2]), .C(acc[2]), .D(n802), .Z(n1748)
         );
  CND2X1 U2373 ( .A(n1749), .B(n1748), .Z(n540) );
  CIVX2 U2374 ( .A(out1_stg2[2]), .Z(n1751) );
  CMX2X1 U2375 ( .A0(out1_stg2[1]), .A1(N210), .S(n1288), .Z(n543) );
  CANR2X1 U2376 ( .A(n1207), .B(out1_stg2[1]), .C(acc[1]), .D(n802), .Z(n1752)
         );
  CND2X1 U2377 ( .A(n1753), .B(n1752), .Z(n542) );
  CIVX2 U2378 ( .A(out1_stg2[1]), .Z(n1755) );
  CANR2X1 U2379 ( .A(n1759), .B(acc[1]), .C(n1758), .D(out0_stg2[1]), .Z(n1754) );
  CMX2X1 U2380 ( .A0(out1_stg2[0]), .A1(N209), .S(n1289), .Z(n545) );
  CND2X1 U2381 ( .A(n1757), .B(n1756), .Z(n544) );
  CIVX2 U2382 ( .A(out1_stg2[0]), .Z(n1761) );
  CANR2X1 U2383 ( .A(n1759), .B(acc[0]), .C(n1758), .D(out0_stg2[0]), .Z(n1760) );
  CMX2X1 U2384 ( .A0(out1_stg2[63]), .A1(N272), .S(n1288), .Z(n419) );
  CANR2X1 U2385 ( .A(n1206), .B(out0_stg2[63]), .C(N481), .D(n1205), .Z(n1764)
         );
  CANR2X1 U2386 ( .A(n1207), .B(out1_stg2[63]), .C(acc[63]), .D(n802), .Z(
        n1763) );
  CND2X1 U2387 ( .A(n1764), .B(n1763), .Z(n546) );
  CND2X1 U2388 ( .A(cmd0_en_stg2_d), .B(n798), .Z(n1897) );
  CIVX2 U2389 ( .A(out0_stg2[63]), .Z(n1769) );
  CIVX2 U2390 ( .A(n1766), .Z(n1894) );
  CIVX2 U2391 ( .A(out0_stg2[0]), .Z(n1771) );
  CAN2X1 U2392 ( .A(n1899), .B(n1362), .Z(n1986) );
  CIVX2 U2393 ( .A(out0_stg2[1]), .Z(n1773) );
  CIVX2 U2394 ( .A(out0_stg2[2]), .Z(n1775) );
  CMXI2X1 U2395 ( .A0(n1204), .A1(n1203), .S(n1362), .Z(n2198) );
  CIVX2 U2396 ( .A(out0_stg2[3]), .Z(n1777) );
  CIVX2 U2397 ( .A(out0_stg2[4]), .Z(n1779) );
  CMXI2X1 U2398 ( .A0(n1202), .A1(n1201), .S(n1362), .Z(n2197) );
  CIVX2 U2399 ( .A(out0_stg2[5]), .Z(n1781) );
  CIVX2 U2400 ( .A(out0_stg2[6]), .Z(n1783) );
  CMXI2X1 U2401 ( .A0(n1200), .A1(n1199), .S(n1362), .Z(n2200) );
  CIVX2 U2402 ( .A(out0_stg2[7]), .Z(n1785) );
  CIVX2 U2403 ( .A(out0_stg2[8]), .Z(n1787) );
  CMXI2X1 U2404 ( .A0(n1198), .A1(n1197), .S(n1361), .Z(n2199) );
  CIVX2 U2405 ( .A(out0_stg2[9]), .Z(n1789) );
  CIVX2 U2406 ( .A(out0_stg2[10]), .Z(n1791) );
  CMXI2X1 U2407 ( .A0(n1196), .A1(n1195), .S(n1361), .Z(n1993) );
  CIVX2 U2408 ( .A(out0_stg2[11]), .Z(n1793) );
  CIVX2 U2409 ( .A(out0_stg2[12]), .Z(n1795) );
  CMXI2X1 U2410 ( .A0(n1194), .A1(n1193), .S(n1361), .Z(n1992) );
  CIVX2 U2411 ( .A(out0_stg2[13]), .Z(n1797) );
  CIVX2 U2412 ( .A(out0_stg2[14]), .Z(n1799) );
  CMXI2X1 U2413 ( .A0(n1192), .A1(n1191), .S(n1361), .Z(n1995) );
  CIVX2 U2414 ( .A(out0_stg2[15]), .Z(n1801) );
  CIVX2 U2415 ( .A(out0_stg2[16]), .Z(n1803) );
  CMXI2X1 U2416 ( .A0(n1190), .A1(n1189), .S(n1361), .Z(n1994) );
  CIVX2 U2417 ( .A(out0_stg2[17]), .Z(n1805) );
  CIVX2 U2418 ( .A(out0_stg2[18]), .Z(n1807) );
  CMXI2X1 U2419 ( .A0(n1188), .A1(n1187), .S(n1361), .Z(n1997) );
  CIVX2 U2420 ( .A(out0_stg2[19]), .Z(n1809) );
  CIVX2 U2421 ( .A(out0_stg2[20]), .Z(n1811) );
  CMXI2X1 U2422 ( .A0(n1186), .A1(n1185), .S(n1361), .Z(n1996) );
  CIVX2 U2423 ( .A(out0_stg2[21]), .Z(n1813) );
  CIVX2 U2424 ( .A(out0_stg2[22]), .Z(n1815) );
  CMXI2X1 U2425 ( .A0(n1184), .A1(n1183), .S(n1361), .Z(n1999) );
  CIVX2 U2426 ( .A(out0_stg2[23]), .Z(n1817) );
  CIVX2 U2427 ( .A(out0_stg2[24]), .Z(n1819) );
  CMXI2X1 U2428 ( .A0(n1182), .A1(n1181), .S(n1361), .Z(n1998) );
  CIVX2 U2429 ( .A(out0_stg2[25]), .Z(n1821) );
  CIVX2 U2430 ( .A(out0_stg2[26]), .Z(n1823) );
  CMXI2X1 U2431 ( .A0(n1180), .A1(n1179), .S(n1361), .Z(n2001) );
  CIVX2 U2432 ( .A(out0_stg2[27]), .Z(n1825) );
  CIVX2 U2433 ( .A(out0_stg2[28]), .Z(n1827) );
  CMXI2X1 U2434 ( .A0(n1178), .A1(n1177), .S(n1361), .Z(n2000) );
  CIVX2 U2435 ( .A(out0_stg2[29]), .Z(n1829) );
  CIVX2 U2436 ( .A(out0_stg2[30]), .Z(n1831) );
  CMXI2X1 U2437 ( .A0(n1176), .A1(n1175), .S(n1360), .Z(n2003) );
  CIVX2 U2438 ( .A(out0_stg2[31]), .Z(n1833) );
  CIVX2 U2439 ( .A(out0_stg2[32]), .Z(n1835) );
  CMXI2X1 U2440 ( .A0(n1174), .A1(n1166), .S(n1360), .Z(n2002) );
  CIVX2 U2441 ( .A(out0_stg2[33]), .Z(n1837) );
  CIVX2 U2442 ( .A(out0_stg2[34]), .Z(n1839) );
  CMXI2X1 U2443 ( .A0(n1165), .A1(n1164), .S(n1360), .Z(n2005) );
  CIVX2 U2444 ( .A(out0_stg2[35]), .Z(n1841) );
  CIVX2 U2445 ( .A(out0_stg2[36]), .Z(n1843) );
  CMXI2X1 U2446 ( .A0(n1163), .A1(n1162), .S(n1360), .Z(n2004) );
  CIVX2 U2447 ( .A(out0_stg2[37]), .Z(n1845) );
  CIVX2 U2448 ( .A(out0_stg2[38]), .Z(n1847) );
  CMXI2X1 U2449 ( .A0(n1161), .A1(n1160), .S(n1360), .Z(n2007) );
  CIVX2 U2450 ( .A(out0_stg2[39]), .Z(n1849) );
  CIVX2 U2451 ( .A(out0_stg2[40]), .Z(n1851) );
  CMXI2X1 U2452 ( .A0(n1159), .A1(n1171), .S(n1360), .Z(n2006) );
  CIVX2 U2453 ( .A(out0_stg2[41]), .Z(n1853) );
  CIVX2 U2454 ( .A(out0_stg2[42]), .Z(n1855) );
  CMXI2X1 U2455 ( .A0(n1170), .A1(n1173), .S(n1360), .Z(n2010) );
  CIVX2 U2456 ( .A(out0_stg2[43]), .Z(n1857) );
  CIVX2 U2457 ( .A(out0_stg2[44]), .Z(n1859) );
  CMXI2X1 U2458 ( .A0(n1172), .A1(n1169), .S(n1360), .Z(n2009) );
  CIVX2 U2459 ( .A(out0_stg2[45]), .Z(n1861) );
  CIVX2 U2460 ( .A(out0_stg2[46]), .Z(n1863) );
  CMXI2X1 U2461 ( .A0(n1168), .A1(n1167), .S(n1360), .Z(n2012) );
  CIVX2 U2462 ( .A(out0_stg2[47]), .Z(n1865) );
  CIVX2 U2463 ( .A(out0_stg2[48]), .Z(n1867) );
  CMXI2X1 U2464 ( .A0(n1155), .A1(n1156), .S(n1360), .Z(n2011) );
  CIVX2 U2465 ( .A(out0_stg2[49]), .Z(n1869) );
  CIVX2 U2466 ( .A(out0_stg2[50]), .Z(n1871) );
  CMXI2X1 U2467 ( .A0(n1157), .A1(n1158), .S(n1360), .Z(n2014) );
  CIVX2 U2468 ( .A(out0_stg2[51]), .Z(n1873) );
  CIVX2 U2469 ( .A(out0_stg2[52]), .Z(n1875) );
  CMXI2X1 U2470 ( .A0(n1151), .A1(n1152), .S(n1359), .Z(n2013) );
  CIVX2 U2471 ( .A(out0_stg2[53]), .Z(n1877) );
  CIVX2 U2472 ( .A(out0_stg2[54]), .Z(n1879) );
  CMXI2X1 U2473 ( .A0(n1153), .A1(n1154), .S(n1359), .Z(n2016) );
  CIVX2 U2474 ( .A(out0_stg2[58]), .Z(n1881) );
  CIVX2 U2475 ( .A(out0_stg2[57]), .Z(n1883) );
  CANR2X1 U2476 ( .A(acc[57]), .B(n1894), .C(out1_stg2[57]), .D(n1212), .Z(
        n1882) );
  CIVX2 U2477 ( .A(out0_stg2[55]), .Z(n1885) );
  CIVX2 U2478 ( .A(out0_stg2[56]), .Z(n1887) );
  CMXI2X1 U2479 ( .A0(n1150), .A1(n1149), .S(n1359), .Z(n2015) );
  CIVX2 U2480 ( .A(out0_stg2[60]), .Z(n1889) );
  CIVX2 U2481 ( .A(out0_stg2[59]), .Z(n1891) );
  CIVX2 U2482 ( .A(out0_stg2[62]), .Z(n1893) );
  CIVX2 U2483 ( .A(out0_stg2[61]), .Z(n1896) );
  CMXI2X1 U2484 ( .A0(n1195), .A1(n1194), .S(n1359), .Z(n2132) );
  CMXI2X1 U2485 ( .A0(n1193), .A1(n1192), .S(n1359), .Z(n2041) );
  CMXI2X1 U2486 ( .A0(n1191), .A1(n1190), .S(n1359), .Z(n2040) );
  CMXI2X1 U2487 ( .A0(n1189), .A1(n1188), .S(n1359), .Z(n2043) );
  CMXI2X1 U2488 ( .A0(n1187), .A1(n1186), .S(n1359), .Z(n2042) );
  CMXI2X1 U2489 ( .A0(n1185), .A1(n1184), .S(n1359), .Z(n2045) );
  CMXI2X1 U2490 ( .A0(n1183), .A1(n1182), .S(n1359), .Z(n2044) );
  CMXI2X1 U2491 ( .A0(n1181), .A1(n1180), .S(n1358), .Z(n2047) );
  CMXI2X1 U2492 ( .A0(n1179), .A1(n1178), .S(n1358), .Z(n2046) );
  CMXI2X1 U2493 ( .A0(n1177), .A1(n1176), .S(n1358), .Z(n2049) );
  CMXI2X1 U2494 ( .A0(n1175), .A1(n1174), .S(n1358), .Z(n2048) );
  CMXI2X1 U2495 ( .A0(n1166), .A1(n1165), .S(n1358), .Z(n2051) );
  CMXI2X1 U2496 ( .A0(n1164), .A1(n1163), .S(n1358), .Z(n2050) );
  CMXI2X1 U2497 ( .A0(n1162), .A1(n1161), .S(n1358), .Z(n2053) );
  CMXI2X1 U2498 ( .A0(n1160), .A1(n1159), .S(n1358), .Z(n2052) );
  CMXI2X1 U2499 ( .A0(n1171), .A1(n1170), .S(n1358), .Z(n2055) );
  CMXI2X1 U2500 ( .A0(n1173), .A1(n1172), .S(n1359), .Z(n2054) );
  CMXI2X1 U2501 ( .A0(n1169), .A1(n1168), .S(n1358), .Z(n2058) );
  CMXI2X1 U2502 ( .A0(n1167), .A1(n1155), .S(n1358), .Z(n2057) );
  CMXI2X1 U2503 ( .A0(n1156), .A1(n1157), .S(n1357), .Z(n2060) );
  CMXI2X1 U2504 ( .A0(n1158), .A1(n1151), .S(n1357), .Z(n2059) );
  CMXI2X1 U2505 ( .A0(n1152), .A1(n1153), .S(n1357), .Z(n2062) );
  CMXI2X1 U2506 ( .A0(n1154), .A1(n1150), .S(n1357), .Z(n2061) );
  CIVX2 U2507 ( .A(acc_cmd2[57]), .Z(n1898) );
  CMXI2X1 U2508 ( .A0(n1149), .A1(n1898), .S(n1357), .Z(n2064) );
  CMXI2X1 U2509 ( .A0(n1203), .A1(n1202), .S(n1357), .Z(n2232) );
  CMXI2X1 U2510 ( .A0(n1201), .A1(n1200), .S(n1357), .Z(n2231) );
  CMXI2X1 U2511 ( .A0(n1199), .A1(n1198), .S(n1357), .Z(n2234) );
  CMXI2X1 U2512 ( .A0(n1197), .A1(n1196), .S(n1357), .Z(n2233) );
  CIVX2 U2513 ( .A(h0_stg0[6]), .Z(n1902) );
  CIVX2 U2514 ( .A(n799), .Z(n1913) );
  CIVX2 U2515 ( .A(n969), .Z(n1901) );
  COND2X1 U2516 ( .A(n799), .B(n1902), .C(n1913), .D(n1901), .Z(n631) );
  CIVX2 U2517 ( .A(h0_stg0[5]), .Z(n1904) );
  CIVX2 U2518 ( .A(n1105), .Z(n1903) );
  COND2X1 U2519 ( .A(n799), .B(n1904), .C(n1913), .D(n1903), .Z(n628) );
  CIVX2 U2520 ( .A(h0_stg0[4]), .Z(n1906) );
  CIVX2 U2521 ( .A(n1116), .Z(n1905) );
  COND2X1 U2522 ( .A(n799), .B(n1906), .C(n1913), .D(n1905), .Z(n625) );
  CIVX2 U2523 ( .A(h0_stg0[3]), .Z(n1908) );
  CIVX2 U2524 ( .A(n965), .Z(n1907) );
  COND2X1 U2525 ( .A(n799), .B(n1908), .C(n1913), .D(n1907), .Z(n622) );
  CIVX2 U2526 ( .A(h0_stg0[2]), .Z(n1910) );
  CIVX2 U2527 ( .A(n1143), .Z(n1909) );
  COND2X1 U2528 ( .A(n799), .B(n1910), .C(n1913), .D(n1909), .Z(n619) );
  CIVX2 U2529 ( .A(h0_stg0[1]), .Z(n1912) );
  COND2X1 U2530 ( .A(n799), .B(n1912), .C(n1913), .D(n1911), .Z(n616) );
  CIVX2 U2531 ( .A(h0_stg0[0]), .Z(n1914) );
  COND2X1 U2532 ( .A(n799), .B(n1914), .C(n1377), .D(n1913), .Z(n613) );
  CIVX2 U2533 ( .A(n12), .Z(n1915) );
  CIVX2 U2534 ( .A(z[2]), .Z(n1919) );
  CIVX2 U2535 ( .A(acc[2]), .Z(n1918) );
  CIVX2 U2536 ( .A(z[4]), .Z(n1921) );
  CIVX2 U2537 ( .A(acc[4]), .Z(n1920) );
  CIVX2 U2538 ( .A(z[5]), .Z(n1923) );
  CIVX2 U2539 ( .A(acc[5]), .Z(n1922) );
  CIVX2 U2540 ( .A(z[6]), .Z(n1925) );
  CIVX2 U2541 ( .A(acc[6]), .Z(n1924) );
  CIVX2 U2542 ( .A(z[7]), .Z(n1927) );
  CIVX2 U2543 ( .A(acc[7]), .Z(n1926) );
  CIVX2 U2544 ( .A(z[8]), .Z(n1929) );
  CIVX2 U2545 ( .A(acc[8]), .Z(n1928) );
  CIVX2 U2546 ( .A(z[10]), .Z(n1931) );
  CIVX2 U2547 ( .A(acc[10]), .Z(n1930) );
  CIVX2 U2548 ( .A(z[12]), .Z(n1933) );
  CIVX2 U2549 ( .A(acc[12]), .Z(n1932) );
  CIVX2 U2550 ( .A(z[13]), .Z(n1935) );
  CIVX2 U2551 ( .A(acc[13]), .Z(n1934) );
  CIVX2 U2552 ( .A(z[14]), .Z(n1937) );
  CIVX2 U2553 ( .A(acc[14]), .Z(n1936) );
  CIVX2 U2554 ( .A(z[15]), .Z(n1939) );
  CIVX2 U2555 ( .A(acc[15]), .Z(n1938) );
  CIVX2 U2556 ( .A(z[16]), .Z(n1941) );
  CIVX2 U2557 ( .A(acc[16]), .Z(n1940) );
  CIVX2 U2558 ( .A(z[17]), .Z(n1943) );
  CIVX2 U2559 ( .A(acc[17]), .Z(n1942) );
  CIVX2 U2560 ( .A(z[18]), .Z(n1945) );
  CIVX2 U2561 ( .A(acc[18]), .Z(n1944) );
  CIVX2 U2562 ( .A(z[19]), .Z(n1947) );
  CIVX2 U2563 ( .A(acc[19]), .Z(n1946) );
  CIVX2 U2564 ( .A(z[20]), .Z(n1949) );
  CIVX2 U2565 ( .A(acc[20]), .Z(n1948) );
  CIVX2 U2566 ( .A(z[21]), .Z(n1951) );
  CIVX2 U2567 ( .A(acc[21]), .Z(n1950) );
  CIVX2 U2568 ( .A(z[22]), .Z(n1953) );
  CIVX2 U2569 ( .A(acc[22]), .Z(n1952) );
  CIVX2 U2570 ( .A(z[23]), .Z(n1955) );
  CIVX2 U2571 ( .A(acc[23]), .Z(n1954) );
  CIVX2 U2572 ( .A(z[24]), .Z(n1957) );
  CIVX2 U2573 ( .A(acc[24]), .Z(n1956) );
  CIVX2 U2574 ( .A(z[25]), .Z(n1959) );
  CIVX2 U2575 ( .A(acc[25]), .Z(n1958) );
  CIVX2 U2576 ( .A(z[26]), .Z(n1961) );
  CIVX2 U2577 ( .A(acc[26]), .Z(n1960) );
  CIVX2 U2578 ( .A(z[27]), .Z(n1963) );
  CIVX2 U2579 ( .A(acc[27]), .Z(n1962) );
  CIVX2 U2580 ( .A(z[28]), .Z(n1965) );
  CIVX2 U2581 ( .A(acc[28]), .Z(n1964) );
  CIVX2 U2582 ( .A(z[29]), .Z(n1967) );
  CIVX2 U2583 ( .A(acc[29]), .Z(n1966) );
  CIVX2 U2584 ( .A(z[30]), .Z(n1969) );
  CIVX2 U2585 ( .A(acc[30]), .Z(n1968) );
  CIVX2 U2586 ( .A(z[31]), .Z(n1971) );
  CIVX2 U2587 ( .A(acc[31]), .Z(n1970) );
  CIVX2 U2588 ( .A(n1120), .Z(n1976) );
  CIVX2 U2589 ( .A(n1122), .Z(n1977) );
  CIVX2 U2590 ( .A(n2271), .Z(n1980) );
  CIVX2 U2591 ( .A(n2280), .Z(n1981) );
  CIVX2 U2592 ( .A(n2281), .Z(n1982) );
  CIVX2 U2593 ( .A(n2282), .Z(n1983) );
  CIVX2 U2594 ( .A(n2283), .Z(n1984) );
  CIVX2 U2595 ( .A(cmd2_en_stg1), .Z(n1985) );
  CMXI2X1 U2596 ( .A0(n1986), .A1(n2198), .S(n1364), .Z(n1987) );
  CMXI2X1 U2597 ( .A0(n2197), .A1(n2200), .S(n1364), .Z(n2255) );
  CMXI2X1 U2598 ( .A0(n1987), .A1(n2255), .S(n1216), .Z(n1988) );
  CMXI2X1 U2599 ( .A0(n2199), .A1(n1993), .S(n1364), .Z(n2254) );
  CMXI2X1 U2600 ( .A0(n1992), .A1(n1995), .S(n1364), .Z(n2025) );
  CMXI2X1 U2601 ( .A0(n2254), .A1(n2025), .S(n1217), .Z(n2302) );
  CMXI2X1 U2602 ( .A0(n1988), .A1(n2302), .S(n1371), .Z(n1989) );
  CMXI2X1 U2603 ( .A0(n1994), .A1(n1997), .S(n1364), .Z(n2024) );
  CMXI2X1 U2604 ( .A0(n1996), .A1(n1999), .S(n1364), .Z(n2027) );
  CMXI2X1 U2605 ( .A0(n2024), .A1(n2027), .S(n1213), .Z(n2301) );
  CMXI2X1 U2606 ( .A0(n1998), .A1(n2001), .S(n1364), .Z(n2026) );
  CMXI2X1 U2607 ( .A0(n2000), .A1(n2003), .S(n1364), .Z(n2029) );
  CMXI2X1 U2608 ( .A0(n2026), .A1(n2029), .S(n1214), .Z(n2169) );
  CMXI2X1 U2609 ( .A0(n2301), .A1(n2169), .S(n1371), .Z(n2099) );
  CMXI2X1 U2610 ( .A0(n1989), .A1(n2099), .S(n1221), .Z(n1990) );
  CMXI2X1 U2611 ( .A0(n2002), .A1(n2005), .S(n1364), .Z(n2028) );
  CMXI2X1 U2612 ( .A0(n2004), .A1(n2007), .S(n1364), .Z(n2031) );
  CMXI2X1 U2613 ( .A0(n2028), .A1(n2031), .S(n1214), .Z(n2168) );
  CMXI2X1 U2614 ( .A0(n2006), .A1(n2010), .S(n1364), .Z(n2030) );
  CMXI2X1 U2615 ( .A0(n2009), .A1(n2012), .S(n1364), .Z(n2034) );
  CMXI2X1 U2616 ( .A0(n2030), .A1(n2034), .S(n1217), .Z(n2171) );
  CMXI2X1 U2617 ( .A0(n2168), .A1(n2171), .S(n1371), .Z(n2098) );
  CMXI2X1 U2618 ( .A0(n2011), .A1(n2014), .S(n1365), .Z(n2033) );
  CMXI2X1 U2619 ( .A0(n2013), .A1(n2016), .S(n1365), .Z(n2036) );
  CMXI2X1 U2620 ( .A0(n2033), .A1(n2036), .S(n1215), .Z(n2170) );
  CMX2X1 U2621 ( .A0(acc_cmd2[58]), .A1(acc_cmd2[57]), .S(n1363), .Z(n2018) );
  CMXI2X1 U2622 ( .A0(n2015), .A1(n2018), .S(n1365), .Z(n2035) );
  CMX2X1 U2623 ( .A0(acc_cmd2[60]), .A1(acc_cmd2[59]), .S(n1363), .Z(n2017) );
  CMX2X1 U2624 ( .A0(acc_cmd2[62]), .A1(acc_cmd2[61]), .S(n1363), .Z(n2020) );
  CMXI2X1 U2625 ( .A0(n2017), .A1(n2020), .S(n1365), .Z(n2038) );
  CMXI2X1 U2626 ( .A0(n2035), .A1(n2038), .S(n1216), .Z(n2173) );
  CMXI2X1 U2627 ( .A0(n2170), .A1(n2173), .S(n1371), .Z(n2101) );
  CMXI2X1 U2628 ( .A0(n2098), .A1(n2101), .S(n1219), .Z(n2218) );
  CMXI2X1 U2629 ( .A0(n1990), .A1(n2218), .S(n1224), .Z(n1991) );
  CND2IX1 U2630 ( .B(n1224), .A(n2217), .Z(n2284) );
  CMXI2X1 U2631 ( .A0(n1993), .A1(n1992), .S(n1365), .Z(n2285) );
  CMXI2X1 U2632 ( .A0(n1995), .A1(n1994), .S(n1365), .Z(n2069) );
  CMXI2X1 U2633 ( .A0(n2285), .A1(n2069), .S(n1217), .Z(n2202) );
  CMXI2X1 U2634 ( .A0(n1997), .A1(n1996), .S(n1365), .Z(n2068) );
  CMXI2X1 U2635 ( .A0(n1999), .A1(n1998), .S(n1365), .Z(n2071) );
  CMXI2X1 U2636 ( .A0(n2068), .A1(n2071), .S(n1215), .Z(n2117) );
  CMXI2X1 U2637 ( .A0(n2202), .A1(n2117), .S(n1371), .Z(n2008) );
  CMXI2X1 U2638 ( .A0(n2001), .A1(n2000), .S(n1365), .Z(n2070) );
  CMXI2X1 U2639 ( .A0(n2003), .A1(n2002), .S(n1365), .Z(n2073) );
  CMXI2X1 U2640 ( .A0(n2070), .A1(n2073), .S(n1213), .Z(n2116) );
  CMXI2X1 U2641 ( .A0(n2005), .A1(n2004), .S(n1365), .Z(n2072) );
  CMXI2X1 U2642 ( .A0(n2007), .A1(n2006), .S(n1365), .Z(n2075) );
  CMXI2X1 U2643 ( .A0(n2072), .A1(n2075), .S(n1213), .Z(n2119) );
  CMXI2X1 U2644 ( .A0(n2116), .A1(n2119), .S(n1371), .Z(n2182) );
  CMXI2X1 U2645 ( .A0(n2008), .A1(n2182), .S(n1220), .Z(n2021) );
  CMXI2X1 U2646 ( .A0(n2010), .A1(n2009), .S(n1366), .Z(n2074) );
  CMXI2X1 U2647 ( .A0(n2012), .A1(n2011), .S(n1366), .Z(n2078) );
  CMXI2X1 U2648 ( .A0(n2074), .A1(n2078), .S(n1214), .Z(n2118) );
  CMXI2X1 U2649 ( .A0(n2014), .A1(n2013), .S(n1366), .Z(n2077) );
  CMXI2X1 U2650 ( .A0(n2016), .A1(n2015), .S(n1366), .Z(n2080) );
  CMXI2X1 U2651 ( .A0(n2077), .A1(n2080), .S(n1215), .Z(n2121) );
  CMXI2X1 U2652 ( .A0(n2118), .A1(n2121), .S(n1371), .Z(n2181) );
  CMXI2X1 U2653 ( .A0(n2018), .A1(n2017), .S(n1366), .Z(n2079) );
  CMXI2X1 U2654 ( .A0(n2020), .A1(n2019), .S(n1366), .Z(n2081) );
  CMXI2X1 U2655 ( .A0(n2079), .A1(n2081), .S(n1216), .Z(n2120) );
  CMXI2X1 U2656 ( .A0(n2181), .A1(n2183), .S(n1221), .Z(n2246) );
  CMXI2X1 U2657 ( .A0(n2132), .A1(n2041), .S(n1366), .Z(n2293) );
  CMXI2X1 U2658 ( .A0(n2040), .A1(n2043), .S(n1366), .Z(n2084) );
  CMXI2X1 U2659 ( .A0(n2293), .A1(n2084), .S(n1214), .Z(n2236) );
  CMXI2X1 U2660 ( .A0(n2042), .A1(n2045), .S(n1366), .Z(n2083) );
  CMXI2X1 U2661 ( .A0(n2044), .A1(n2047), .S(n1366), .Z(n2086) );
  CMXI2X1 U2662 ( .A0(n2083), .A1(n2086), .S(n1216), .Z(n2124) );
  CMXI2X1 U2663 ( .A0(n2236), .A1(n2124), .S(n1371), .Z(n2022) );
  CMXI2X1 U2664 ( .A0(n2046), .A1(n2049), .S(n1366), .Z(n2085) );
  CMXI2X1 U2665 ( .A0(n2048), .A1(n2051), .S(n1366), .Z(n2088) );
  CMXI2X1 U2666 ( .A0(n2085), .A1(n2088), .S(n1217), .Z(n2123) );
  CMXI2X1 U2667 ( .A0(n2050), .A1(n2053), .S(n1367), .Z(n2087) );
  CMXI2X1 U2668 ( .A0(n2052), .A1(n2055), .S(n1367), .Z(n2090) );
  CMXI2X1 U2669 ( .A0(n2087), .A1(n2090), .S(n1213), .Z(n2126) );
  CMXI2X1 U2670 ( .A0(n2123), .A1(n2126), .S(n1371), .Z(n2186) );
  CMXI2X1 U2671 ( .A0(n2022), .A1(n2186), .S(n1222), .Z(n2023) );
  CMXI2X1 U2672 ( .A0(n2054), .A1(n2058), .S(n1367), .Z(n2089) );
  CMXI2X1 U2673 ( .A0(n2057), .A1(n2060), .S(n1367), .Z(n2093) );
  CMXI2X1 U2674 ( .A0(n2089), .A1(n2093), .S(n1217), .Z(n2125) );
  CMXI2X1 U2675 ( .A0(n2059), .A1(n2062), .S(n1367), .Z(n2092) );
  CMXI2X1 U2676 ( .A0(n2061), .A1(n2064), .S(n1367), .Z(n2095) );
  CMXI2X1 U2677 ( .A0(n2092), .A1(n2095), .S(n1215), .Z(n2128) );
  CMXI2X1 U2678 ( .A0(n2125), .A1(n2128), .S(n1371), .Z(n2185) );
  CMX2X1 U2679 ( .A0(acc_cmd2[59]), .A1(acc_cmd2[58]), .S(n1363), .Z(n2063) );
  CMX2X1 U2680 ( .A0(acc_cmd2[61]), .A1(acc_cmd2[60]), .S(n1363), .Z(n2066) );
  CMXI2X1 U2681 ( .A0(n2063), .A1(n2066), .S(n1367), .Z(n2094) );
  CMX2X1 U2682 ( .A0(acc_cmd2[63]), .A1(acc_cmd2[62]), .S(n1363), .Z(n2065) );
  CMXI2X1 U2683 ( .A0(n2094), .A1(n2096), .S(n1214), .Z(n2127) );
  CMXI2X1 U2684 ( .A0(n2185), .A1(n2187), .S(n1220), .Z(n2247) );
  CMXI2X1 U2685 ( .A0(n2025), .A1(n2024), .S(n1215), .Z(n2256) );
  CMXI2X1 U2686 ( .A0(n2027), .A1(n2026), .S(n1216), .Z(n2141) );
  CMXI2X1 U2687 ( .A0(n2256), .A1(n2141), .S(n1371), .Z(n2032) );
  CMXI2X1 U2688 ( .A0(n2029), .A1(n2028), .S(n1213), .Z(n2140) );
  CMXI2X1 U2689 ( .A0(n2031), .A1(n2030), .S(n1216), .Z(n2143) );
  CMXI2X1 U2690 ( .A0(n2140), .A1(n2143), .S(n1371), .Z(n2190) );
  CMXI2X1 U2691 ( .A0(n2032), .A1(n2190), .S(n1222), .Z(n2039) );
  CMXI2X1 U2692 ( .A0(n2034), .A1(n2033), .S(n1217), .Z(n2142) );
  CMXI2X1 U2693 ( .A0(n2036), .A1(n2035), .S(n1213), .Z(n2145) );
  CMXI2X1 U2694 ( .A0(n2142), .A1(n2145), .S(n1372), .Z(n2189) );
  CMXI2X1 U2695 ( .A0(n2038), .A1(n2037), .S(n1214), .Z(n2144) );
  CMXI2X1 U2696 ( .A0(n2189), .A1(n2191), .S(n1223), .Z(n2248) );
  CMXI2X1 U2697 ( .A0(n2041), .A1(n2040), .S(n1367), .Z(n2133) );
  CMXI2X1 U2698 ( .A0(n2043), .A1(n2042), .S(n1367), .Z(n2104) );
  CMXI2X1 U2699 ( .A0(n2133), .A1(n2104), .S(n1214), .Z(n2274) );
  CMXI2X1 U2700 ( .A0(n2045), .A1(n2044), .S(n1367), .Z(n2103) );
  CMXI2X1 U2701 ( .A0(n2047), .A1(n2046), .S(n1367), .Z(n2106) );
  CMXI2X1 U2702 ( .A0(n2103), .A1(n2106), .S(n1217), .Z(n2148) );
  CMXI2X1 U2703 ( .A0(n2274), .A1(n2148), .S(n1372), .Z(n2056) );
  CMXI2X1 U2704 ( .A0(n2049), .A1(n2048), .S(n1367), .Z(n2105) );
  CMXI2X1 U2705 ( .A0(n2051), .A1(n2050), .S(n1368), .Z(n2108) );
  CMXI2X1 U2706 ( .A0(n2105), .A1(n2108), .S(n1215), .Z(n2147) );
  CMXI2X1 U2707 ( .A0(n2053), .A1(n2052), .S(n1368), .Z(n2107) );
  CMXI2X1 U2708 ( .A0(n2055), .A1(n2054), .S(n1368), .Z(n2110) );
  CMXI2X1 U2709 ( .A0(n2107), .A1(n2110), .S(n1216), .Z(n2150) );
  CMXI2X1 U2710 ( .A0(n2147), .A1(n2150), .S(n1372), .Z(n2194) );
  CMXI2X1 U2711 ( .A0(n2056), .A1(n2194), .S(n1218), .Z(n2067) );
  CMXI2X1 U2712 ( .A0(n2058), .A1(n2057), .S(n1368), .Z(n2109) );
  CMXI2X1 U2713 ( .A0(n2060), .A1(n2059), .S(n1368), .Z(n2112) );
  CMXI2X1 U2714 ( .A0(n2109), .A1(n2112), .S(n1217), .Z(n2149) );
  CMXI2X1 U2715 ( .A0(n2062), .A1(n2061), .S(n1368), .Z(n2111) );
  CMXI2X1 U2716 ( .A0(n2064), .A1(n2063), .S(n1368), .Z(n2114) );
  CMXI2X1 U2717 ( .A0(n2111), .A1(n2114), .S(n1215), .Z(n2152) );
  CMXI2X1 U2718 ( .A0(n2149), .A1(n2152), .S(n1372), .Z(n2193) );
  CMXI2X1 U2719 ( .A0(n2066), .A1(n2065), .S(n1368), .Z(n2113) );
  CMXI2X1 U2720 ( .A0(n2193), .A1(n2195), .S(n1219), .Z(n2249) );
  CMXI2X1 U2721 ( .A0(n2069), .A1(n2068), .S(n1213), .Z(n2287) );
  CMXI2X1 U2722 ( .A0(n2071), .A1(n2070), .S(n1213), .Z(n2155) );
  CMXI2X1 U2723 ( .A0(n2287), .A1(n2155), .S(n1372), .Z(n2076) );
  CMXI2X1 U2724 ( .A0(n2073), .A1(n2072), .S(n1214), .Z(n2154) );
  CMXI2X1 U2725 ( .A0(n2075), .A1(n2074), .S(n1215), .Z(n2157) );
  CMXI2X1 U2726 ( .A0(n2154), .A1(n2157), .S(n1372), .Z(n2210) );
  CMXI2X1 U2727 ( .A0(n2076), .A1(n2210), .S(n1220), .Z(n2082) );
  CMXI2X1 U2728 ( .A0(n2078), .A1(n2077), .S(n1216), .Z(n2156) );
  CMXI2X1 U2729 ( .A0(n2080), .A1(n2079), .S(n1214), .Z(n2159) );
  CMXI2X1 U2730 ( .A0(n2156), .A1(n2159), .S(n1372), .Z(n2209) );
  CMXI2X1 U2731 ( .A0(n2209), .A1(n2211), .S(n1221), .Z(n2250) );
  CMXI2X1 U2732 ( .A0(n2084), .A1(n2083), .S(n1216), .Z(n2295) );
  CMXI2X1 U2733 ( .A0(n2086), .A1(n2085), .S(n1217), .Z(n2162) );
  CMXI2X1 U2734 ( .A0(n2295), .A1(n2162), .S(n1372), .Z(n2091) );
  CMXI2X1 U2735 ( .A0(n2088), .A1(n2087), .S(n1213), .Z(n2161) );
  CMXI2X1 U2736 ( .A0(n2090), .A1(n2089), .S(n1217), .Z(n2164) );
  CMXI2X1 U2737 ( .A0(n2161), .A1(n2164), .S(n1372), .Z(n2214) );
  CMXI2X1 U2738 ( .A0(n2091), .A1(n2214), .S(n1223), .Z(n2097) );
  CMXI2X1 U2739 ( .A0(n2093), .A1(n2092), .S(n1215), .Z(n2163) );
  CMXI2X1 U2740 ( .A0(n2095), .A1(n2094), .S(n1214), .Z(n2166) );
  CMXI2X1 U2741 ( .A0(n2163), .A1(n2166), .S(n1372), .Z(n2213) );
  CMXI2X1 U2742 ( .A0(n2213), .A1(n2215), .S(n1221), .Z(n2251) );
  CMXI2X1 U2743 ( .A0(n2099), .A1(n2098), .S(n1222), .Z(n2102) );
  CMXI2X1 U2744 ( .A0(n2101), .A1(n2100), .S(n1223), .Z(n2252) );
  CMXI2X1 U2745 ( .A0(n2104), .A1(n2103), .S(n1215), .Z(n2307) );
  CMXI2X1 U2746 ( .A0(n2106), .A1(n2105), .S(n1216), .Z(n2176) );
  CMXI2X1 U2747 ( .A0(n2307), .A1(n2176), .S(n1372), .Z(n2135) );
  CMXI2X1 U2748 ( .A0(n2108), .A1(n2107), .S(n1213), .Z(n2175) );
  CMXI2X1 U2749 ( .A0(n2110), .A1(n2109), .S(n1216), .Z(n2178) );
  CMXI2X1 U2750 ( .A0(n2175), .A1(n2178), .S(n1372), .Z(n2138) );
  CMXI2X1 U2751 ( .A0(n2135), .A1(n2138), .S(n1218), .Z(n2115) );
  CMXI2X1 U2752 ( .A0(n2112), .A1(n2111), .S(n1217), .Z(n2177) );
  CMXI2X1 U2753 ( .A0(n2114), .A1(n2113), .S(n1213), .Z(n2179) );
  CMXI2X1 U2754 ( .A0(n2177), .A1(n2179), .S(n1373), .Z(n2137) );
  CMXI2X1 U2755 ( .A0(n2117), .A1(n2116), .S(n1373), .Z(n2204) );
  CMXI2X1 U2756 ( .A0(n2119), .A1(n2118), .S(n1373), .Z(n2207) );
  CMXI2X1 U2757 ( .A0(n2204), .A1(n2207), .S(n1222), .Z(n2122) );
  CMXI2X1 U2758 ( .A0(n2121), .A1(n2120), .S(n1373), .Z(n2206) );
  CMXI2X1 U2759 ( .A0(n2124), .A1(n2123), .S(n1373), .Z(n2238) );
  CMXI2X1 U2760 ( .A0(n2126), .A1(n2125), .S(n1373), .Z(n2222) );
  CMXI2X1 U2761 ( .A0(n2238), .A1(n2222), .S(n1218), .Z(n2129) );
  CMXI2X1 U2762 ( .A0(n2128), .A1(n2127), .S(n1373), .Z(n2221) );
  CMXI2X1 U2763 ( .A0(n2130), .A1(n2232), .S(n1368), .Z(n2131) );
  CMXI2X1 U2764 ( .A0(n2231), .A1(n2234), .S(n1368), .Z(n2273) );
  CMXI2X1 U2765 ( .A0(n2131), .A1(n2273), .S(n1214), .Z(n2134) );
  CMXI2X1 U2766 ( .A0(n2233), .A1(n2132), .S(n1368), .Z(n2272) );
  CMXI2X1 U2767 ( .A0(n2272), .A1(n2133), .S(n1214), .Z(n2308) );
  CMXI2X1 U2768 ( .A0(n2134), .A1(n2308), .S(n1373), .Z(n2136) );
  CMXI2X1 U2769 ( .A0(n2136), .A1(n2135), .S(n1219), .Z(n2139) );
  CMXI2X1 U2770 ( .A0(n2138), .A1(n2137), .S(n1220), .Z(n2219) );
  CMXI2X1 U2771 ( .A0(n2141), .A1(n2140), .S(n1373), .Z(n2258) );
  CMXI2X1 U2772 ( .A0(n2143), .A1(n2142), .S(n1373), .Z(n2224) );
  CMXI2X1 U2773 ( .A0(n2258), .A1(n2224), .S(n1221), .Z(n2146) );
  CMXI2X1 U2774 ( .A0(n2145), .A1(n2144), .S(n1373), .Z(n2223) );
  CMXI2X1 U2775 ( .A0(n2148), .A1(n2147), .S(n1373), .Z(n2276) );
  CMXI2X1 U2776 ( .A0(n2150), .A1(n2149), .S(n1374), .Z(n2226) );
  CMXI2X1 U2777 ( .A0(n2276), .A1(n2226), .S(n1222), .Z(n2153) );
  CMXI2X1 U2778 ( .A0(n2152), .A1(n2151), .S(n1374), .Z(n2225) );
  CMXI2X1 U2779 ( .A0(n2155), .A1(n2154), .S(n1374), .Z(n2289) );
  CMXI2X1 U2780 ( .A0(n2157), .A1(n2156), .S(n1374), .Z(n2228) );
  CMXI2X1 U2781 ( .A0(n2289), .A1(n2228), .S(n1223), .Z(n2160) );
  CMXI2X1 U2782 ( .A0(n2159), .A1(n2158), .S(n1374), .Z(n2227) );
  CMXI2X1 U2783 ( .A0(n2162), .A1(n2161), .S(n1374), .Z(n2297) );
  CMXI2X1 U2784 ( .A0(n2164), .A1(n2163), .S(n1374), .Z(n2230) );
  CMXI2X1 U2785 ( .A0(n2297), .A1(n2230), .S(n1219), .Z(n2167) );
  CMXI2X1 U2786 ( .A0(n2166), .A1(n2165), .S(n1374), .Z(n2229) );
  CMXI2X1 U2787 ( .A0(n2169), .A1(n2168), .S(n1374), .Z(n2303) );
  CMXI2X1 U2788 ( .A0(n2171), .A1(n2170), .S(n1374), .Z(n2243) );
  CMXI2X1 U2789 ( .A0(n2303), .A1(n2243), .S(n1223), .Z(n2174) );
  CMXI2X1 U2790 ( .A0(n2173), .A1(n2172), .S(n1374), .Z(n2242) );
  CMXI2X1 U2791 ( .A0(n2176), .A1(n2175), .S(n1374), .Z(n2309) );
  CMXI2X1 U2792 ( .A0(n2178), .A1(n2177), .S(n1375), .Z(n2245) );
  CMXI2X1 U2793 ( .A0(n2309), .A1(n2245), .S(n1218), .Z(n2180) );
  CMXI2X1 U2794 ( .A0(n2182), .A1(n2181), .S(n1219), .Z(n2184) );
  CMXI2X1 U2795 ( .A0(n2186), .A1(n2185), .S(n1220), .Z(n2188) );
  CMXI2X1 U2796 ( .A0(n2190), .A1(n2189), .S(n1218), .Z(n2192) );
  CMXI2X1 U2797 ( .A0(n2194), .A1(n2193), .S(n1220), .Z(n2196) );
  CMXI2X1 U2798 ( .A0(n2198), .A1(n2197), .S(n1368), .Z(n2201) );
  CMXI2X1 U2799 ( .A0(n2200), .A1(n2199), .S(n1369), .Z(n2286) );
  CMXI2X1 U2800 ( .A0(n2201), .A1(n2286), .S(n1217), .Z(n2203) );
  CMXI2X1 U2801 ( .A0(n2203), .A1(n2202), .S(n1375), .Z(n2205) );
  CMXI2X1 U2802 ( .A0(n2205), .A1(n2204), .S(n1221), .Z(n2208) );
  CMXI2X1 U2803 ( .A0(n2207), .A1(n2206), .S(n1222), .Z(n2220) );
  CMXI2X1 U2804 ( .A0(n2210), .A1(n2209), .S(n1223), .Z(n2212) );
  CMXI2X1 U2805 ( .A0(n2214), .A1(n2213), .S(n1218), .Z(n2216) );
  CMXI2X1 U2806 ( .A0(n2222), .A1(n2221), .S(n1219), .Z(n2240) );
  CMXI2X1 U2807 ( .A0(n2224), .A1(n2223), .S(n1221), .Z(n2260) );
  CMXI2X1 U2808 ( .A0(n2226), .A1(n2225), .S(n1219), .Z(n2278) );
  CMXI2X1 U2809 ( .A0(n2228), .A1(n2227), .S(n1220), .Z(n2291) );
  CMXI2X1 U2810 ( .A0(n2230), .A1(n2229), .S(n1221), .Z(n2299) );
  CMXI2X1 U2811 ( .A0(n2232), .A1(n2231), .S(n1369), .Z(n2235) );
  CMXI2X1 U2812 ( .A0(n2234), .A1(n2233), .S(n1369), .Z(n2294) );
  CMXI2X1 U2813 ( .A0(n2235), .A1(n2294), .S(n1215), .Z(n2237) );
  CMXI2X1 U2814 ( .A0(n2237), .A1(n2236), .S(n1375), .Z(n2239) );
  CMXI2X1 U2815 ( .A0(n2239), .A1(n2238), .S(n1222), .Z(n2241) );
  CMXI2X1 U2816 ( .A0(n2243), .A1(n2242), .S(n1220), .Z(n2305) );
  CMXI2X1 U2817 ( .A0(n2245), .A1(n2244), .S(n1222), .Z(n2311) );
  CMXI2X1 U2818 ( .A0(n2255), .A1(n2254), .S(n1216), .Z(n2257) );
  CMXI2X1 U2819 ( .A0(n2257), .A1(n2256), .S(n1375), .Z(n2259) );
  CMXI2X1 U2820 ( .A0(n2259), .A1(n2258), .S(n1223), .Z(n2261) );
  CMXI2X1 U2821 ( .A0(n2273), .A1(n2272), .S(n1217), .Z(n2275) );
  CMXI2X1 U2822 ( .A0(n2275), .A1(n2274), .S(n1375), .Z(n2277) );
  CMXI2X1 U2823 ( .A0(n2277), .A1(n2276), .S(n1218), .Z(n2279) );
  CMXI2X1 U2824 ( .A0(n2286), .A1(n2285), .S(n1215), .Z(n2288) );
  CMXI2X1 U2825 ( .A0(n2288), .A1(n2287), .S(n1375), .Z(n2290) );
  CMXI2X1 U2826 ( .A0(n2290), .A1(n2289), .S(n1219), .Z(n2292) );
  CMXI2X1 U2827 ( .A0(n2294), .A1(n2293), .S(n1213), .Z(n2296) );
  CMXI2X1 U2828 ( .A0(n2296), .A1(n2295), .S(n1375), .Z(n2298) );
  CMXI2X1 U2829 ( .A0(n2298), .A1(n2297), .S(n1220), .Z(n2300) );
  CMXI2X1 U2830 ( .A0(n2302), .A1(n2301), .S(n1375), .Z(n2304) );
  CMXI2X1 U2831 ( .A0(n2304), .A1(n2303), .S(n1221), .Z(n2306) );
  CMXI2X1 U2832 ( .A0(n2308), .A1(n2307), .S(n1375), .Z(n2310) );
  CMXI2X1 U2833 ( .A0(n2310), .A1(n2309), .S(n1223), .Z(n2312) );
endmodule

