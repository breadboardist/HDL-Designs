
module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push0, cmd0_en_0, cmd1_en_0, cmd2_en_0, cmd0_en_1, cmd1_en_1, push0_0,
         cmd0_en_2_d, cmd1_en_2_d, push0_2, push0_1, cmd2_en_1, cmd2_en_2,
         cmd0_en_2, cmd1_en_2, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         roundit, n851, n852, n853, n854, n855, n859, n862, n863, n864, n865,
         n866, n867, n868, n870, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n885, n889, n891, n892, n897, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n916, n917, n919, n920, n921, n922, n923, n924, n925,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n938, n940,
         n946, n949, n950, n952, n957, n959, n961, n973, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1057,
         n1116, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022;
  wire   [1:0] cmd0;
  wire   [1:0] cmd0_0;
  wire   [1:0] cmd0_2;
  wire   [1:0] cmd0_1;
  wire   [63:0] out0_2;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] acc;
  wire   [63:0] out1_2;
  wire   [63:0] out1_0;
  wire   [63:0] out1_1;
  wire   [63:0] out2_2;
  wire   [6:0] h0_1;
  wire   [6:0] h0_0;

  CFD2QX1 cmd0_en_2_d_reg ( .D(cmd0_en_2), .CP(clk), .CD(n7935), .Q(
        cmd0_en_2_d) );
  CFD2QX1 cmd1_en_2_d_reg ( .D(n8022), .CP(clk), .CD(n7935), .Q(cmd1_en_2_d)
         );
  CFD2QX1 \out0_2_reg[1]  ( .D(n1183), .CP(clk), .CD(n7935), .Q(out0_2[1]) );
  CFD2QX1 \out0_2_reg[2]  ( .D(n1182), .CP(clk), .CD(n7935), .Q(out0_2[2]) );
  CFD2QX1 \out0_2_reg[3]  ( .D(n1181), .CP(clk), .CD(n7935), .Q(out0_2[3]) );
  CFD2QX1 \out0_2_reg[4]  ( .D(n1180), .CP(clk), .CD(n7935), .Q(out0_2[4]) );
  CFD2QX1 \out0_2_reg[5]  ( .D(n1179), .CP(clk), .CD(n7935), .Q(out0_2[5]) );
  CFD2QX1 \out0_2_reg[6]  ( .D(n1178), .CP(clk), .CD(n7935), .Q(out0_2[6]) );
  CFD2QX1 \out0_2_reg[7]  ( .D(n1177), .CP(clk), .CD(n7935), .Q(out0_2[7]) );
  CFD2QX1 \out0_2_reg[8]  ( .D(n1176), .CP(clk), .CD(n7935), .Q(out0_2[8]) );
  CFD2QX1 \out0_2_reg[9]  ( .D(n1175), .CP(clk), .CD(n7935), .Q(out0_2[9]) );
  CFD2QX1 \out0_2_reg[10]  ( .D(n1174), .CP(clk), .CD(n7935), .Q(out0_2[10])
         );
  CFD2QX1 \out0_2_reg[11]  ( .D(n1173), .CP(clk), .CD(n7935), .Q(out0_2[11])
         );
  CFD2QX1 \out0_2_reg[12]  ( .D(n1172), .CP(clk), .CD(n7935), .Q(out0_2[12])
         );
  CFD2QX1 \out0_2_reg[13]  ( .D(n1171), .CP(clk), .CD(n7935), .Q(out0_2[13])
         );
  CFD2QX1 \out0_2_reg[14]  ( .D(n1170), .CP(clk), .CD(n7935), .Q(out0_2[14])
         );
  CFD2QX1 \out0_2_reg[15]  ( .D(n1169), .CP(clk), .CD(n7935), .Q(out0_2[15])
         );
  CFD2QX1 \out0_2_reg[19]  ( .D(n1165), .CP(clk), .CD(n7935), .Q(out0_2[19])
         );
  CFD2QX1 \out0_2_reg[22]  ( .D(n1162), .CP(clk), .CD(n7935), .Q(out0_2[22])
         );
  CFD2QX1 \out0_2_reg[23]  ( .D(n1161), .CP(clk), .CD(n7935), .Q(out0_2[23])
         );
  CFD2QX1 \out0_2_reg[24]  ( .D(n1160), .CP(clk), .CD(n7935), .Q(out0_2[24])
         );
  CFD2QX1 \out0_2_reg[25]  ( .D(n1159), .CP(clk), .CD(n7935), .Q(out0_2[25])
         );
  CFD2QX1 \out0_2_reg[26]  ( .D(n1158), .CP(clk), .CD(n7935), .Q(out0_2[26])
         );
  CFD2QX1 \out0_2_reg[27]  ( .D(n1157), .CP(clk), .CD(n7935), .Q(out0_2[27])
         );
  CFD2QX1 \out0_2_reg[31]  ( .D(n1153), .CP(clk), .CD(n7935), .Q(out0_2[31])
         );
  CFD2QX1 \out0_2_reg[35]  ( .D(n1149), .CP(clk), .CD(n7935), .Q(out0_2[35])
         );
  CFD2QX1 \out0_2_reg[40]  ( .D(n1144), .CP(clk), .CD(n7935), .Q(out0_2[40])
         );
  CFD2QX1 \out0_2_reg[41]  ( .D(n1143), .CP(clk), .CD(n7935), .Q(out0_2[41])
         );
  CFD2QX1 \out0_2_reg[43]  ( .D(n1141), .CP(clk), .CD(n7935), .Q(out0_2[43])
         );
  CFD2QX1 \out0_2_reg[47]  ( .D(n1137), .CP(clk), .CD(n7935), .Q(out0_2[47])
         );
  CFD2QX1 \out1_2_reg[0]  ( .D(n7934), .CP(clk), .CD(n7935), .Q(out1_2[0]) );
  CFD2QX1 \out1_2_reg[1]  ( .D(n7933), .CP(clk), .CD(n7935), .Q(out1_2[1]) );
  CFD2QX1 \out1_2_reg[2]  ( .D(n7932), .CP(clk), .CD(n7935), .Q(out1_2[2]) );
  CFD2QX1 \out1_2_reg[4]  ( .D(n1116), .CP(clk), .CD(n7935), .Q(out1_2[4]) );
  CFD2QX1 \acc_reg[24]  ( .D(n1017), .CP(clk), .CD(n7935), .Q(acc[24]) );
  CFD2QX1 \acc_reg[4]  ( .D(n997), .CP(clk), .CD(n7935), .Q(acc[4]) );
  CFD2QX1 \q0_reg[16]  ( .D(n1316), .CP(clk), .CD(n7935), .Q(q0[16]) );
  CFD2QX1 \h0_reg[9]  ( .D(n938), .CP(clk), .CD(n7935), .Q(h0[9]) );
  CFD2QX1 \h0_reg[6]  ( .D(n935), .CP(clk), .CD(n7935), .Q(h0[6]) );
  CFD2QX1 \h0_1_reg[1]  ( .D(n1291), .CP(clk), .CD(n7935), .Q(h0_1[1]) );
  CFD2QX1 \h0_1_reg[0]  ( .D(n1290), .CP(clk), .CD(n7935), .Q(h0_1[0]) );
  CFD2QXL \out1_0_reg[46]  ( .D(N61), .CP(clk), .CD(n7935), .Q(out1_0[46]) );
  CFD2QXL \out1_0_reg[47]  ( .D(N62), .CP(clk), .CD(n7935), .Q(out1_0[47]) );
  CFD2QXL \out1_0_reg[49]  ( .D(N64), .CP(clk), .CD(n7935), .Q(out1_0[49]) );
  CFD2QXL \out1_0_reg[57]  ( .D(N72), .CP(clk), .CD(n7935), .Q(out1_0[57]) );
  CFD2QXL \out1_0_reg[35]  ( .D(N50), .CP(clk), .CD(n7935), .Q(out1_0[35]) );
  CFD2QXL \out2_2_reg[3]  ( .D(n3199), .CP(clk), .CD(n7935), .Q(out2_2[3]) );
  CFD2QXL \out2_2_reg[4]  ( .D(n3188), .CP(clk), .CD(n7935), .Q(out2_2[4]) );
  CFD2QXL \out2_2_reg[9]  ( .D(n3142), .CP(clk), .CD(n7935), .Q(out2_2[9]) );
  CFD2QXL \out2_2_reg[12]  ( .D(n3135), .CP(clk), .CD(n7935), .Q(out2_2[12])
         );
  CFD2QXL \out2_2_reg[14]  ( .D(n1448), .CP(clk), .CD(n7935), .Q(out2_2[14])
         );
  CFD2QXL \out2_2_reg[21]  ( .D(n3094), .CP(clk), .CD(n7935), .Q(out2_2[21])
         );
  CFD2QXL \out1_0_reg[63]  ( .D(N78), .CP(clk), .CD(n7935), .Q(out1_0[63]) );
  CFD2QXL \out1_0_reg[40]  ( .D(N55), .CP(clk), .CD(n7935), .Q(out1_0[40]) );
  CFD2QXL \out1_0_reg[39]  ( .D(N54), .CP(clk), .CD(n7935), .Q(out1_0[39]) );
  CFD2QXL \out1_0_reg[38]  ( .D(N53), .CP(clk), .CD(n7935), .Q(out1_0[38]) );
  CFD2QXL \out1_0_reg[37]  ( .D(N52), .CP(clk), .CD(n7935), .Q(out1_0[37]) );
  CFD2QXL \out1_0_reg[36]  ( .D(N51), .CP(clk), .CD(n7935), .Q(out1_0[36]) );
  CFD2QXL \out1_0_reg[34]  ( .D(N49), .CP(clk), .CD(n7935), .Q(out1_0[34]) );
  CFD2QXL \out1_0_reg[33]  ( .D(N48), .CP(clk), .CD(n7935), .Q(out1_0[33]) );
  CFD2QXL \out1_0_reg[32]  ( .D(N47), .CP(clk), .CD(n7935), .Q(out1_0[32]) );
  CFD2QXL \out1_0_reg[31]  ( .D(N46), .CP(clk), .CD(n7935), .Q(out1_0[31]) );
  CFD2QXL \out1_0_reg[30]  ( .D(N45), .CP(clk), .CD(n7935), .Q(out1_0[30]) );
  CFD2QXL \out1_0_reg[29]  ( .D(N44), .CP(clk), .CD(n7935), .Q(out1_0[29]) );
  CFD2QXL \out1_0_reg[28]  ( .D(N43), .CP(clk), .CD(n7935), .Q(out1_0[28]) );
  CFD2QXL \out1_0_reg[27]  ( .D(N42), .CP(clk), .CD(n7935), .Q(out1_0[27]) );
  CFD2QXL \out1_0_reg[26]  ( .D(N41), .CP(clk), .CD(n7935), .Q(out1_0[26]) );
  CFD2QXL \out1_0_reg[24]  ( .D(N39), .CP(clk), .CD(n7935), .Q(out1_0[24]) );
  CFD2QXL \out1_0_reg[23]  ( .D(N38), .CP(clk), .CD(n7935), .Q(out1_0[23]) );
  CFD2QXL \out1_0_reg[22]  ( .D(N37), .CP(clk), .CD(n7935), .Q(out1_0[22]) );
  CFD2QXL \out1_0_reg[21]  ( .D(N36), .CP(clk), .CD(n7935), .Q(out1_0[21]) );
  CFD2QXL \out1_0_reg[20]  ( .D(N35), .CP(clk), .CD(n7935), .Q(out1_0[20]) );
  CFD2QXL \out1_0_reg[19]  ( .D(N34), .CP(clk), .CD(n7935), .Q(out1_0[19]) );
  CFD2QXL \out1_0_reg[18]  ( .D(N33), .CP(clk), .CD(n7935), .Q(out1_0[18]) );
  CFD2QXL \out1_0_reg[17]  ( .D(N32), .CP(clk), .CD(n7935), .Q(out1_0[17]) );
  CFD2QXL \out1_0_reg[16]  ( .D(N31), .CP(clk), .CD(n7935), .Q(out1_0[16]) );
  CFD2QXL \out1_0_reg[15]  ( .D(N30), .CP(clk), .CD(n7935), .Q(out1_0[15]) );
  CFD2QXL \out1_0_reg[14]  ( .D(N29), .CP(clk), .CD(n7935), .Q(out1_0[14]) );
  CFD2QXL \out1_0_reg[13]  ( .D(N28), .CP(clk), .CD(n7935), .Q(out1_0[13]) );
  CFD2QXL \out1_0_reg[12]  ( .D(N27), .CP(clk), .CD(n7935), .Q(out1_0[12]) );
  CFD2QXL \out1_0_reg[11]  ( .D(N26), .CP(clk), .CD(n7935), .Q(out1_0[11]) );
  CFD2QXL \out1_0_reg[10]  ( .D(N25), .CP(clk), .CD(n7935), .Q(out1_0[10]) );
  CFD2QXL \out1_0_reg[9]  ( .D(N24), .CP(clk), .CD(n7935), .Q(out1_0[9]) );
  CFD2QXL \out1_0_reg[8]  ( .D(N23), .CP(clk), .CD(n7935), .Q(out1_0[8]) );
  CFD2QXL \out1_0_reg[7]  ( .D(N22), .CP(clk), .CD(n7935), .Q(out1_0[7]) );
  CFD2QXL \out1_0_reg[6]  ( .D(N21), .CP(clk), .CD(n7935), .Q(out1_0[6]) );
  CFD2QXL \out1_0_reg[52]  ( .D(N67), .CP(clk), .CD(n7935), .Q(out1_0[52]) );
  CFD2QXL \out1_0_reg[54]  ( .D(N69), .CP(clk), .CD(n7935), .Q(out1_0[54]) );
  CFD2QXL \out1_0_reg[58]  ( .D(N73), .CP(clk), .CD(n7935), .Q(out1_0[58]) );
  CFD2QXL \out1_0_reg[62]  ( .D(N77), .CP(clk), .CD(n7935), .Q(out1_0[62]) );
  CFD2QXL \out2_2_reg[5]  ( .D(n2892), .CP(clk), .CD(n7935), .Q(out2_2[5]) );
  CFD2QXL \out2_2_reg[7]  ( .D(n855), .CP(clk), .CD(n7935), .Q(out2_2[7]) );
  CFD1QXL roundit_reg ( .D(n2940), .CP(clk), .Q(roundit) );
  CFD2QXL \out2_2_reg[28]  ( .D(n1431), .CP(clk), .CD(n7935), .Q(out2_2[28])
         );
  CFD2QXL \out2_2_reg[27]  ( .D(n1433), .CP(clk), .CD(n7935), .Q(out2_2[27])
         );
  CFD2QXL \out2_2_reg[11]  ( .D(n1434), .CP(clk), .CD(n7935), .Q(out2_2[11])
         );
  CFD2QXL \out2_2_reg[24]  ( .D(n3023), .CP(clk), .CD(n7935), .Q(out2_2[24])
         );
  CFD2QXL \out2_2_reg[8]  ( .D(n3158), .CP(clk), .CD(n7935), .Q(out2_2[8]) );
  CFD2QXL \acc_reg[25]  ( .D(n1018), .CP(clk), .CD(n7935), .Q(acc[25]) );
  CFD2QXL \acc_reg[23]  ( .D(n1016), .CP(clk), .CD(n7935), .Q(acc[23]) );
  CFD2QXL \acc_reg[22]  ( .D(n1015), .CP(clk), .CD(n7935), .Q(acc[22]) );
  CFD2QXL \acc_reg[21]  ( .D(n1289), .CP(clk), .CD(n7935), .Q(acc[21]) );
  CFD2QXL \acc_reg[20]  ( .D(n1283), .CP(clk), .CD(n7935), .Q(acc[20]) );
  CFD2QXL \acc_reg[19]  ( .D(n1012), .CP(clk), .CD(n7935), .Q(acc[19]) );
  CFD2QXL \acc_reg[18]  ( .D(n1011), .CP(clk), .CD(n7935), .Q(acc[18]) );
  CFD2QXL \acc_reg[15]  ( .D(n1008), .CP(clk), .CD(n7935), .Q(acc[15]) );
  CFD2QXL \acc_reg[13]  ( .D(n1006), .CP(clk), .CD(n7935), .Q(acc[13]) );
  CFD2QXL \acc_reg[7]  ( .D(n1000), .CP(clk), .CD(n7935), .Q(acc[7]) );
  CFD2QXL \acc_reg[6]  ( .D(n999), .CP(clk), .CD(n7935), .Q(acc[6]) );
  CFD2QXL \acc_reg[5]  ( .D(n998), .CP(clk), .CD(n7935), .Q(acc[5]) );
  CFD2QXL \acc_reg[3]  ( .D(n996), .CP(clk), .CD(n7935), .Q(acc[3]) );
  CFD2QXL \out2_2_reg[0]  ( .D(n892), .CP(clk), .CD(n7935), .Q(out2_2[0]) );
  CFD2QXL \out1_2_reg[8]  ( .D(n7927), .CP(clk), .CD(n7935), .Q(out1_2[8]) );
  CFD2QXL \out1_2_reg[9]  ( .D(n7926), .CP(clk), .CD(n7935), .Q(out1_2[9]) );
  CFD2QXL \out1_2_reg[10]  ( .D(n7925), .CP(clk), .CD(n7935), .Q(out1_2[10])
         );
  CFD2QXL \out2_2_reg[22]  ( .D(n1393), .CP(clk), .CD(n7935), .Q(out2_2[22])
         );
  CFD2QXL \out2_2_reg[6]  ( .D(n3052), .CP(clk), .CD(n7935), .Q(out2_2[6]) );
  CFD2QXL \out2_2_reg[19]  ( .D(n1390), .CP(clk), .CD(n7935), .Q(out2_2[19])
         );
  CFD2QXL \out2_2_reg[1]  ( .D(n865), .CP(clk), .CD(n7935), .Q(out2_2[1]) );
  CFD2QXL \out2_2_reg[30]  ( .D(n1288), .CP(clk), .CD(n7935), .Q(out2_2[30])
         );
  CFD2QXL \out2_2_reg[26]  ( .D(n2856), .CP(clk), .CD(n7935), .Q(out2_2[26])
         );
  CFD2QXL \out2_2_reg[18]  ( .D(n2850), .CP(clk), .CD(n7935), .Q(out2_2[18])
         );
  CFD2QXL \out2_2_reg[10]  ( .D(n2837), .CP(clk), .CD(n7935), .Q(out2_2[10])
         );
  CFD2QXL \acc_reg[63]  ( .D(n1274), .CP(clk), .CD(n7935), .Q(acc[63]) );
  CFD2QXL \acc_reg[48]  ( .D(n1280), .CP(clk), .CD(n7935), .Q(acc[48]) );
  CFD2QXL \acc_reg[47]  ( .D(n1040), .CP(clk), .CD(n7935), .Q(acc[47]) );
  CFD2QXL \acc_reg[46]  ( .D(n1344), .CP(clk), .CD(n7935), .Q(acc[46]) );
  CFD2QXL \acc_reg[43]  ( .D(n1036), .CP(clk), .CD(n7935), .Q(acc[43]) );
  CFD2QXL \acc_reg[41]  ( .D(n1034), .CP(clk), .CD(n7935), .Q(acc[41]) );
  CFD2QXL \acc_reg[40]  ( .D(n1033), .CP(clk), .CD(n7935), .Q(acc[40]) );
  CFD2QXL \acc_reg[34]  ( .D(n1343), .CP(clk), .CD(n7935), .Q(acc[34]) );
  CFD2QXL \out2_2_reg[2]  ( .D(n885), .CP(clk), .CD(n7935), .Q(out2_2[2]) );
  CFD2QXL \out0_2_reg[54]  ( .D(n1130), .CP(clk), .CD(n7935), .Q(out0_2[54])
         );
  CFD2QXL \out0_2_reg[58]  ( .D(n1126), .CP(clk), .CD(n7935), .Q(out0_2[58])
         );
  CFD2QXL \out1_2_reg[3]  ( .D(n7931), .CP(clk), .CD(n7935), .Q(out1_2[3]) );
  CFD2QXL \out1_2_reg[14]  ( .D(n7921), .CP(clk), .CD(n7935), .Q(out1_2[14])
         );
  CFD2QXL \acc_reg[14]  ( .D(n1007), .CP(clk), .CD(n7935), .Q(acc[14]) );
  CFD2QXL \acc_reg[31]  ( .D(n1024), .CP(clk), .CD(n7935), .Q(acc[31]) );
  CFD2QXL \acc_reg[30]  ( .D(n1286), .CP(clk), .CD(n7935), .Q(acc[30]) );
  CFD2QXL \acc_reg[29]  ( .D(n1285), .CP(clk), .CD(n7935), .Q(acc[29]) );
  CFD2QXL \acc_reg[27]  ( .D(n1020), .CP(clk), .CD(n7935), .Q(acc[27]) );
  CFD2QXL \acc_reg[26]  ( .D(n1019), .CP(clk), .CD(n7935), .Q(acc[26]) );
  CFD2QXL \out1_2_reg[5]  ( .D(n7930), .CP(clk), .CD(n7935), .Q(out1_2[5]) );
  CFD2QXL \out1_2_reg[6]  ( .D(n7929), .CP(clk), .CD(n7935), .Q(out1_2[6]) );
  CFD2QXL \out1_2_reg[7]  ( .D(n7928), .CP(clk), .CD(n7935), .Q(out1_2[7]) );
  CFD2QXL \out1_2_reg[11]  ( .D(n7924), .CP(clk), .CD(n7935), .Q(out1_2[11])
         );
  CFD2QXL \out1_2_reg[12]  ( .D(n7923), .CP(clk), .CD(n7935), .Q(out1_2[12])
         );
  CFD2QXL \out1_2_reg[13]  ( .D(n7922), .CP(clk), .CD(n7935), .Q(out1_2[13])
         );
  CFD2QXL \out1_2_reg[15]  ( .D(n7920), .CP(clk), .CD(n7935), .Q(out1_2[15])
         );
  CFD2QXL \out1_2_reg[16]  ( .D(n7919), .CP(clk), .CD(n7935), .Q(out1_2[16])
         );
  CFD2QXL \out1_2_reg[17]  ( .D(n7918), .CP(clk), .CD(n7935), .Q(out1_2[17])
         );
  CFD2QXL \out1_2_reg[18]  ( .D(n7917), .CP(clk), .CD(n7935), .Q(out1_2[18])
         );
  CFD2QXL \out1_2_reg[19]  ( .D(n7916), .CP(clk), .CD(n7935), .Q(out1_2[19])
         );
  CFD2QXL \out1_2_reg[20]  ( .D(n7915), .CP(clk), .CD(n7935), .Q(out1_2[20])
         );
  CFD2QXL \out1_2_reg[21]  ( .D(n7914), .CP(clk), .CD(n7935), .Q(out1_2[21])
         );
  CFD2QXL \out1_2_reg[22]  ( .D(n7913), .CP(clk), .CD(n7935), .Q(out1_2[22])
         );
  CFD2QXL \out1_2_reg[23]  ( .D(n7912), .CP(clk), .CD(n7935), .Q(out1_2[23])
         );
  CFD2QXL \out1_2_reg[24]  ( .D(n7911), .CP(clk), .CD(n7935), .Q(out1_2[24])
         );
  CFD2QXL \out1_2_reg[25]  ( .D(n7910), .CP(clk), .CD(n7935), .Q(out1_2[25])
         );
  CFD2QXL \out1_2_reg[26]  ( .D(n7909), .CP(clk), .CD(n7935), .Q(out1_2[26])
         );
  CFD2QXL \out1_2_reg[27]  ( .D(n7908), .CP(clk), .CD(n7935), .Q(out1_2[27])
         );
  CFD2QXL \out1_2_reg[28]  ( .D(n7907), .CP(clk), .CD(n7935), .Q(out1_2[28])
         );
  CFD2QXL \out1_2_reg[29]  ( .D(n7906), .CP(clk), .CD(n7935), .Q(out1_2[29])
         );
  CFD2QXL \out1_2_reg[30]  ( .D(n7905), .CP(clk), .CD(n7935), .Q(out1_2[30])
         );
  CFD2QXL \out1_2_reg[31]  ( .D(n7904), .CP(clk), .CD(n7935), .Q(out1_2[31])
         );
  CFD2QXL \out1_2_reg[32]  ( .D(n7903), .CP(clk), .CD(n7935), .Q(out1_2[32])
         );
  CFD2QXL \out1_2_reg[33]  ( .D(n7902), .CP(clk), .CD(n7935), .Q(out1_2[33])
         );
  CFD2QXL \out1_2_reg[34]  ( .D(n7901), .CP(clk), .CD(n7935), .Q(out1_2[34])
         );
  CFD2QXL \out1_2_reg[35]  ( .D(n7900), .CP(clk), .CD(n7935), .Q(out1_2[35])
         );
  CFD2QXL \out1_2_reg[36]  ( .D(n7899), .CP(clk), .CD(n7935), .Q(out1_2[36])
         );
  CFD2QXL \out1_2_reg[37]  ( .D(n7898), .CP(clk), .CD(n7935), .Q(out1_2[37])
         );
  CFD2QXL \out1_2_reg[38]  ( .D(n7897), .CP(clk), .CD(n7935), .Q(out1_2[38])
         );
  CFD2QXL \out1_2_reg[39]  ( .D(n7896), .CP(clk), .CD(n7935), .Q(out1_2[39])
         );
  CFD2QXL \out1_2_reg[40]  ( .D(n7895), .CP(clk), .CD(n7935), .Q(out1_2[40])
         );
  CFD2QXL \out1_2_reg[41]  ( .D(n7894), .CP(clk), .CD(n7935), .Q(out1_2[41])
         );
  CFD2QXL \out1_2_reg[42]  ( .D(n7893), .CP(clk), .CD(n7935), .Q(out1_2[42])
         );
  CFD2QXL \out1_2_reg[43]  ( .D(n7892), .CP(clk), .CD(n7935), .Q(out1_2[43])
         );
  CFD2QXL \out1_2_reg[44]  ( .D(n7891), .CP(clk), .CD(n7935), .Q(out1_2[44])
         );
  CFD2QXL \out1_2_reg[45]  ( .D(n7890), .CP(clk), .CD(n7935), .Q(out1_2[45])
         );
  CFD2QXL \out1_2_reg[46]  ( .D(n7889), .CP(clk), .CD(n7935), .Q(out1_2[46])
         );
  CFD2QXL \out1_2_reg[47]  ( .D(n7888), .CP(clk), .CD(n7935), .Q(out1_2[47])
         );
  CFD2QXL \out1_2_reg[48]  ( .D(n7887), .CP(clk), .CD(n7935), .Q(out1_2[48])
         );
  CFD2QXL \out1_2_reg[49]  ( .D(n7886), .CP(clk), .CD(n7935), .Q(out1_2[49])
         );
  CFD2QXL \out1_2_reg[50]  ( .D(n7885), .CP(clk), .CD(n7935), .Q(out1_2[50])
         );
  CFD2QXL \out1_2_reg[51]  ( .D(n7884), .CP(clk), .CD(n7935), .Q(out1_2[51])
         );
  CFD2QXL \out1_2_reg[52]  ( .D(n7883), .CP(clk), .CD(n7935), .Q(out1_2[52])
         );
  CFD2QXL \out1_2_reg[53]  ( .D(n7882), .CP(clk), .CD(n7935), .Q(out1_2[53])
         );
  CFD2QXL \out1_2_reg[54]  ( .D(n7881), .CP(clk), .CD(n7935), .Q(out1_2[54])
         );
  CFD2QXL \out1_2_reg[55]  ( .D(n7880), .CP(clk), .CD(n7935), .Q(out1_2[55])
         );
  CFD2QXL \out1_2_reg[56]  ( .D(n7879), .CP(clk), .CD(n7935), .Q(out1_2[56])
         );
  CFD2QXL \out1_2_reg[57]  ( .D(n7878), .CP(clk), .CD(n7935), .Q(out1_2[57])
         );
  CFD2QXL \out1_2_reg[58]  ( .D(n7877), .CP(clk), .CD(n7935), .Q(out1_2[58])
         );
  CFD2QXL \out1_2_reg[59]  ( .D(n7876), .CP(clk), .CD(n7935), .Q(out1_2[59])
         );
  CFD2QXL \out1_2_reg[60]  ( .D(n7875), .CP(clk), .CD(n7935), .Q(out1_2[60])
         );
  CFD2QXL \out1_2_reg[61]  ( .D(n7874), .CP(clk), .CD(n7935), .Q(out1_2[61])
         );
  CFD2QXL \out1_2_reg[62]  ( .D(n7873), .CP(clk), .CD(n7935), .Q(out1_2[62])
         );
  CFD2QXL \out1_2_reg[63]  ( .D(n1057), .CP(clk), .CD(n7935), .Q(out1_2[63])
         );
  CFD2XL \out1_0_reg[41]  ( .D(N56), .CP(clk), .CD(n7935), .Q(out1_0[41]) );
  CFD2XL \out1_0_reg[43]  ( .D(N58), .CP(clk), .CD(n7935), .Q(out1_0[43]) );
  CFD2XL \out1_0_reg[42]  ( .D(N57), .CP(clk), .CD(n7935), .Q(out1_0[42]) );
  CFD2XL \out1_0_reg[45]  ( .D(N60), .CP(clk), .CD(n7935), .Q(out1_0[45]) );
  CFD2XL \out1_0_reg[48]  ( .D(N63), .CP(clk), .CD(n7935), .Q(out1_0[48]) );
  CFD2XL \out1_0_reg[50]  ( .D(N65), .CP(clk), .CD(n7935), .Q(out1_0[50]) );
  CFD2XL \out1_0_reg[51]  ( .D(N66), .CP(clk), .CD(n7935), .Q(out1_0[51]) );
  CFD2XL \out1_0_reg[53]  ( .D(N68), .CP(clk), .CD(n7935), .Q(out1_0[53]) );
  CFD2XL \out1_0_reg[55]  ( .D(N70), .CP(clk), .CD(n7935), .Q(out1_0[55]) );
  CFD2XL \out1_0_reg[59]  ( .D(N74), .CP(clk), .CD(n7935), .Q(out1_0[59]) );
  CFD2XL \out1_0_reg[61]  ( .D(N76), .CP(clk), .CD(n7935), .Q(out1_0[61]) );
  CFD2XL \out1_0_reg[44]  ( .D(N59), .CP(clk), .CD(n7935), .Q(out1_0[44]) );
  CFD4X2 \q0_reg[5]  ( .D(n1432), .CP(clk), .SD(n7935), .Q(n7863), .QN(q0[5])
         );
  CFD4X2 \q0_reg[13]  ( .D(n2627), .CP(clk), .SD(n7935), .Q(n7864), .QN(q0[13]) );
  CFD4X1 \q0_reg[31]  ( .D(n2681), .CP(clk), .SD(n7935), .Q(n7870), .QN(q0[31]) );
  CFD4X2 \q0_reg[29]  ( .D(n2679), .CP(clk), .SD(n7935), .Q(n7853), .QN(q0[29]) );
  CFD2XL \out1_0_reg[60]  ( .D(N75), .CP(clk), .CD(n7935), .Q(out1_0[60]) );
  CFD2XL \out1_0_reg[56]  ( .D(N71), .CP(clk), .CD(n7935), .Q(out1_0[56]) );
  CFD4X2 \q0_reg[10]  ( .D(n1473), .CP(clk), .SD(n7935), .Q(n7868), .QN(q0[10]) );
  CFD4X2 \q0_reg[11]  ( .D(n2678), .CP(clk), .SD(n7935), .Q(n7872), .QN(q0[11]) );
  CFD4X2 \q0_reg[1]  ( .D(n2669), .CP(clk), .SD(n7935), .Q(n2624), .QN(q0[1])
         );
  CFD4X2 \q0_reg[19]  ( .D(n2677), .CP(clk), .SD(n7935), .Q(n2658), .QN(q0[19]) );
  CFD4X2 \q0_reg[27]  ( .D(n2626), .CP(clk), .SD(n7935), .Q(n7851), .QN(q0[27]) );
  CFD4X2 \q0_reg[7]  ( .D(n2668), .CP(clk), .SD(n7935), .Q(n2582), .QN(q0[7])
         );
  CFD4X2 \q0_reg[30]  ( .D(n7856), .CP(clk), .SD(n7935), .QN(q0[30]) );
  CFD4X2 \q0_reg[15]  ( .D(n2676), .CP(clk), .SD(n7935), .Q(n7861), .QN(q0[15]) );
  CFD4X2 \q0_reg[2]  ( .D(n7855), .CP(clk), .SD(n7935), .QN(q0[2]) );
  CFD4X2 \q0_reg[3]  ( .D(n2667), .CP(clk), .SD(n7935), .Q(n7862), .QN(q0[3])
         );
  CFD4X1 \q0_reg[24]  ( .D(n2680), .CP(clk), .SD(n7935), .Q(n7871), .QN(q0[24]) );
  CFD4X2 \q0_reg[21]  ( .D(n2675), .CP(clk), .SD(n7935), .Q(n7866), .QN(q0[21]) );
  CFD4X2 \q0_reg[26]  ( .D(n1294), .CP(clk), .SD(n7935), .QN(q0[26]) );
  CFD4X2 \q0_reg[9]  ( .D(n2665), .CP(clk), .SD(n7935), .Q(n7858), .QN(q0[9])
         );
  CFD2QX2 \q0_reg[12]  ( .D(n973), .CP(clk), .CD(n7935), .Q(q0[12]) );
  CFD2QX2 \q0_reg[8]  ( .D(n1439), .CP(clk), .CD(n7935), .Q(q0[8]) );
  CFD4X2 \q0_reg[17]  ( .D(n2674), .CP(clk), .SD(n7935), .Q(n7865), .QN(n7860)
         );
  CFD4X2 \q0_reg[14]  ( .D(n2664), .CP(clk), .SD(n7935), .Q(n7859), .QN(q0[14]) );
  CFD2QX2 \q0_reg[18]  ( .D(n1354), .CP(clk), .CD(n7935), .Q(q0[18]) );
  CFD4X2 \q0_reg[25]  ( .D(n2673), .CP(clk), .SD(n7935), .Q(n7867), .QN(q0[25]) );
  CFD4X2 \q0_reg[23]  ( .D(n2672), .CP(clk), .SD(n7935), .Q(n7869), .QN(q0[23]) );
  CFD2XL push0_2_reg ( .D(n1482), .CP(clk), .CD(n7935), .Q(push0_2), .QN(n8004) );
  CFD2XL \cmd0_2_reg[1]  ( .D(n1490), .CP(clk), .CD(n7935), .Q(cmd0_2[1]) );
  CFD2XL \cmd0_2_reg[0]  ( .D(n1306), .CP(clk), .CD(n7935), .Q(cmd0_2[0]), 
        .QN(n7937) );
  CFD2XL push0_1_reg ( .D(n1492), .CP(clk), .CD(n7935), .Q(push0_1) );
  CFD2XL \out1_1_reg[63]  ( .D(n1494), .CP(clk), .CD(n7935), .Q(out1_1[63]) );
  CFD2XL \out1_1_reg[62]  ( .D(n1302), .CP(clk), .CD(n7935), .Q(out1_1[62]) );
  CFD2XL \out1_1_reg[58]  ( .D(n1500), .CP(clk), .CD(n7935), .Q(out1_1[58]) );
  CFD2XL \out1_1_reg[57]  ( .D(n1504), .CP(clk), .CD(n7935), .Q(out1_1[57]) );
  CFD2XL \out1_1_reg[54]  ( .D(n1498), .CP(clk), .CD(n7935), .Q(out1_1[54]) );
  CFD2XL \out1_1_reg[52]  ( .D(n1506), .CP(clk), .CD(n7935), .Q(out1_1[52]) );
  CFD2XL \out1_1_reg[49]  ( .D(n1480), .CP(clk), .CD(n7935), .Q(out1_1[49]) );
  CFD2XL \out1_1_reg[47]  ( .D(n1502), .CP(clk), .CD(n7935), .Q(out1_1[47]) );
  CFD2XL \out1_1_reg[46]  ( .D(n1304), .CP(clk), .CD(n7935), .Q(out1_1[46]) );
  CFD2XL \out1_1_reg[40]  ( .D(n1268), .CP(clk), .CD(n7935), .Q(out1_1[40]) );
  CFD2XL \out1_1_reg[39]  ( .D(n1325), .CP(clk), .CD(n7935), .Q(out1_1[39]) );
  CFD2XL \out1_1_reg[38]  ( .D(n1295), .CP(clk), .CD(n7935), .Q(out1_1[38]) );
  CFD2XL \out1_1_reg[37]  ( .D(n1312), .CP(clk), .CD(n7935), .Q(out1_1[37]) );
  CFD2XL \out1_1_reg[36]  ( .D(n1317), .CP(clk), .CD(n7935), .Q(out1_1[36]) );
  CFD2XL \out1_1_reg[35]  ( .D(n1350), .CP(clk), .CD(n7935), .Q(out1_1[35]) );
  CFD2XL \out1_1_reg[34]  ( .D(n1348), .CP(clk), .CD(n7935), .Q(out1_1[34]) );
  CFD2XL \out1_1_reg[33]  ( .D(n1319), .CP(clk), .CD(n7935), .Q(out1_1[33]) );
  CFD2XL \out1_1_reg[32]  ( .D(n1451), .CP(clk), .CD(n7935), .Q(out1_1[32]) );
  CFD2XL \out1_1_reg[31]  ( .D(n1308), .CP(clk), .CD(n7935), .Q(out1_1[31]) );
  CFD2XL \out1_1_reg[30]  ( .D(n1533), .CP(clk), .CD(n7935), .Q(out1_1[30]) );
  CFD2XL \out1_1_reg[29]  ( .D(n1321), .CP(clk), .CD(n7935), .Q(out1_1[29]) );
  CFD2XL \out1_1_reg[28]  ( .D(n1300), .CP(clk), .CD(n7935), .Q(out1_1[28]) );
  CFD2XL \out1_1_reg[27]  ( .D(n1526), .CP(clk), .CD(n7935), .Q(out1_1[27]) );
  CFD2XL \out1_1_reg[26]  ( .D(n1467), .CP(clk), .CD(n7935), .Q(out1_1[26]) );
  CFD2XL \out1_1_reg[25]  ( .D(n1471), .CP(clk), .CD(n7935), .Q(out1_1[25]) );
  CFD2XL \out1_1_reg[24]  ( .D(n1275), .CP(clk), .CD(n7935), .Q(out1_1[24]) );
  CFD2XL \out1_1_reg[23]  ( .D(n1528), .CP(clk), .CD(n7935), .Q(out1_1[23]) );
  CFD2XL \out1_1_reg[22]  ( .D(n1496), .CP(clk), .CD(n7935), .Q(out1_1[22]) );
  CFD2XL \out1_1_reg[21]  ( .D(n1531), .CP(clk), .CD(n7935), .Q(out1_1[21]) );
  CFD2XL \out1_1_reg[20]  ( .D(n1461), .CP(clk), .CD(n7935), .Q(out1_1[20]) );
  CFD2XL \out1_1_reg[19]  ( .D(n1346), .CP(clk), .CD(n7935), .Q(out1_1[19]) );
  CFD2XL \out1_1_reg[18]  ( .D(n1352), .CP(clk), .CD(n7935), .Q(out1_1[18]) );
  CFD2XL \out1_1_reg[17]  ( .D(n1453), .CP(clk), .CD(n7935), .Q(out1_1[17]) );
  CFD2XL \out1_1_reg[16]  ( .D(n1469), .CP(clk), .CD(n7935), .Q(out1_1[16]) );
  CFD2XL \out1_1_reg[15]  ( .D(n1359), .CP(clk), .CD(n7935), .Q(out1_1[15]) );
  CFD2XL \out1_1_reg[14]  ( .D(n1355), .CP(clk), .CD(n7935), .Q(out1_1[14]) );
  CFD2XL \out1_1_reg[13]  ( .D(n1329), .CP(clk), .CD(n7935), .Q(out1_1[13]) );
  CFD2XL \out1_1_reg[12]  ( .D(n1465), .CP(clk), .CD(n7935), .Q(out1_1[12]) );
  CFD2XL \out1_1_reg[11]  ( .D(n1436), .CP(clk), .CD(n7935), .Q(out1_1[11]) );
  CFD2XL \out1_1_reg[10]  ( .D(n1444), .CP(clk), .CD(n7935), .Q(out1_1[10]) );
  CFD2XL \out1_1_reg[9]  ( .D(n1457), .CP(clk), .CD(n7935), .Q(out1_1[9]) );
  CFD2XL \out1_1_reg[8]  ( .D(n1459), .CP(clk), .CD(n7935), .Q(out1_1[8]) );
  CFD2XL \out1_1_reg[7]  ( .D(n1378), .CP(clk), .CD(n7935), .Q(out1_1[7]) );
  CFD2XL \out1_1_reg[6]  ( .D(n1455), .CP(clk), .CD(n7935), .Q(out1_1[6]) );
  CFD2XL \out1_1_reg[5]  ( .D(n1463), .CP(clk), .CD(n7935), .Q(out1_1[5]) );
  CFD2XL \out1_1_reg[4]  ( .D(n1476), .CP(clk), .CD(n7935), .Q(out1_1[4]) );
  CFD2XL \out1_1_reg[3]  ( .D(n1474), .CP(clk), .CD(n7935), .Q(out1_1[3]) );
  CFD2XL \out1_1_reg[2]  ( .D(n1478), .CP(clk), .CD(n7935), .Q(out1_1[2]) );
  CFD2XL \out1_1_reg[1]  ( .D(n1310), .CP(clk), .CD(n7935), .Q(out1_1[1]) );
  CFD2XL \out1_1_reg[0]  ( .D(n1484), .CP(clk), .CD(n7935), .Q(out1_1[0]) );
  CFD2XL \cmd0_1_reg[1]  ( .D(n1298), .CP(clk), .CD(n7935), .Q(cmd0_1[1]) );
  CFD2XL \cmd0_1_reg[0]  ( .D(n1314), .CP(clk), .CD(n7935), .Q(cmd0_1[0]) );
  CFD2XL \out1_1_reg[61]  ( .D(n1323), .CP(clk), .CD(n7935), .Q(out1_1[61]) );
  CFD2XL \out1_1_reg[60]  ( .D(n1380), .CP(clk), .CD(n7935), .Q(out1_1[60]) );
  CFD2XL \out1_1_reg[59]  ( .D(n1520), .CP(clk), .CD(n7935), .Q(out1_1[59]) );
  CFD2XL \out1_1_reg[56]  ( .D(n1524), .CP(clk), .CD(n7935), .Q(out1_1[56]) );
  CFD2XL \out1_1_reg[55]  ( .D(n1514), .CP(clk), .CD(n7935), .Q(out1_1[55]) );
  CFD2XL \out1_1_reg[53]  ( .D(n1522), .CP(clk), .CD(n7935), .Q(out1_1[53]) );
  CFD2XL \out1_1_reg[51]  ( .D(n1518), .CP(clk), .CD(n7935), .Q(out1_1[51]) );
  CFD2XL \out1_1_reg[50]  ( .D(n1512), .CP(clk), .CD(n7935), .Q(out1_1[50]) );
  CFD2XL \out1_1_reg[48]  ( .D(n1516), .CP(clk), .CD(n7935), .Q(out1_1[48]) );
  CFD2XL \out1_1_reg[45]  ( .D(n1508), .CP(clk), .CD(n7935), .Q(out1_1[45]) );
  CFD2XL \out1_1_reg[44]  ( .D(n1510), .CP(clk), .CD(n7935), .Q(out1_1[44]) );
  CFD2XL \out1_1_reg[43]  ( .D(n1357), .CP(clk), .CD(n7935), .Q(out1_1[43]) );
  CFD2XL \out1_1_reg[42]  ( .D(n1327), .CP(clk), .CD(n7935), .Q(out1_1[42]) );
  CFD2XL \out1_1_reg[41]  ( .D(n1486), .CP(clk), .CD(n7935), .Q(out1_1[41]) );
  CFD2XL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n7935), .Q(cmd0[1]) );
  CFD2XL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n7935), .Q(cmd0[0]) );
  CFD2XL push0_0_reg ( .D(n1488), .CP(clk), .CD(n7935), .Q(push0_0) );
  CFD2XL \cmd0_0_reg[1]  ( .D(n1442), .CP(clk), .CD(n7935), .Q(cmd0_0[1]) );
  CFD2XL \out0_2_reg[33]  ( .D(n1151), .CP(clk), .CD(n7935), .Q(out0_2[33]) );
  CFD2XL \out0_2_reg[32]  ( .D(n1152), .CP(clk), .CD(n7935), .Q(out0_2[32]), 
        .QN(n2683) );
  CFD2XL \out1_0_reg[0]  ( .D(n1297), .CP(clk), .CD(n7935), .Q(out1_0[0]) );
  CFD2XL \cmd0_0_reg[0]  ( .D(n1281), .CP(clk), .CD(n7935), .Q(cmd0_0[0]) );
  CFD2XL push0_reg ( .D(pushin), .CP(clk), .CD(n7935), .Q(push0) );
  CFD2XL cmd0_en_1_reg ( .D(cmd0_en_0), .CP(clk), .CD(n7935), .Q(cmd0_en_1) );
  CFD2XL cmd1_en_1_reg ( .D(cmd1_en_0), .CP(clk), .CD(n7935), .Q(cmd1_en_1) );
  CFD2XL cmd2_en_1_reg ( .D(cmd2_en_0), .CP(clk), .CD(n7935), .Q(cmd2_en_1), 
        .QN(n7936) );
  CFD2XL _pushout_reg ( .D(n8021), .CP(clk), .CD(n7935), .Q(pushout) );
  CFD2XL \h0_1_reg[2]  ( .D(n921), .CP(clk), .CD(n7935), .Q(h0_1[2]), .QN(
        n8012) );
  CFD2XL \h0_1_reg[3]  ( .D(n924), .CP(clk), .CD(n7935), .Q(h0_1[3]), .QN(
        n8013) );
  CFD2XL \dout_reg[24]  ( .D(n1213), .CP(clk), .CD(n7935), .Q(z[24]) );
  CFD2XL \dout_reg[17]  ( .D(n1424), .CP(clk), .CD(n7935), .Q(z[17]) );
  CFD2XL \dout_reg[16]  ( .D(n1423), .CP(clk), .CD(n7935), .Q(z[16]) );
  CFD2XL \dout_reg[12]  ( .D(n1201), .CP(clk), .CD(n7935), .Q(z[12]) );
  CFD2XL \dout_reg[11]  ( .D(n1200), .CP(clk), .CD(n7935), .Q(z[11]) );
  CFD2XL \dout_reg[10]  ( .D(n1199), .CP(clk), .CD(n7935), .Q(z[10]) );
  CFD2XL \dout_reg[9]  ( .D(n1198), .CP(clk), .CD(n7935), .Q(z[9]) );
  CFD2XL \dout_reg[8]  ( .D(n1197), .CP(clk), .CD(n7935), .Q(z[8]) );
  CFD2XL \dout_reg[2]  ( .D(n1419), .CP(clk), .CD(n7935), .Q(z[2]) );
  CFD2XL \dout_reg[1]  ( .D(n1190), .CP(clk), .CD(n7935), .Q(z[1]) );
  CFD2XL \dout_reg[0]  ( .D(n1189), .CP(clk), .CD(n7935), .Q(z[0]) );
  CFD2XL \h0_0_reg[5]  ( .D(n931), .CP(clk), .CD(n7935), .Q(h0_0[5]) );
  CFD2XL \h0_0_reg[1]  ( .D(n1418), .CP(clk), .CD(n7935), .Q(h0_0[1]) );
  CFD2XL \dout_reg[31]  ( .D(n1417), .CP(clk), .CD(n7935), .Q(z[31]) );
  CFD2XL \dout_reg[30]  ( .D(n1416), .CP(clk), .CD(n7935), .Q(z[30]) );
  CFD2XL \dout_reg[29]  ( .D(n1415), .CP(clk), .CD(n7935), .Q(z[29]) );
  CFD2XL \dout_reg[28]  ( .D(n1414), .CP(clk), .CD(n7935), .Q(z[28]) );
  CFD2XL \dout_reg[27]  ( .D(n1413), .CP(clk), .CD(n7935), .Q(z[27]) );
  CFD2XL \dout_reg[26]  ( .D(n1412), .CP(clk), .CD(n7935), .Q(z[26]) );
  CFD2XL \dout_reg[25]  ( .D(n1411), .CP(clk), .CD(n7935), .Q(z[25]) );
  CFD2XL \dout_reg[23]  ( .D(n1410), .CP(clk), .CD(n7935), .Q(z[23]) );
  CFD2XL \dout_reg[22]  ( .D(n1409), .CP(clk), .CD(n7935), .Q(z[22]) );
  CFD2XL \dout_reg[21]  ( .D(n1408), .CP(clk), .CD(n7935), .Q(z[21]) );
  CFD2XL \dout_reg[20]  ( .D(n1407), .CP(clk), .CD(n7935), .Q(z[20]) );
  CFD2XL \dout_reg[19]  ( .D(n1406), .CP(clk), .CD(n7935), .Q(z[19]) );
  CFD2XL \dout_reg[18]  ( .D(n1405), .CP(clk), .CD(n7935), .Q(z[18]) );
  CFD2XL \dout_reg[15]  ( .D(n1404), .CP(clk), .CD(n7935), .Q(z[15]) );
  CFD2XL \dout_reg[14]  ( .D(n1403), .CP(clk), .CD(n7935), .Q(z[14]) );
  CFD2XL \dout_reg[13]  ( .D(n1402), .CP(clk), .CD(n7935), .Q(z[13]) );
  CFD2XL \dout_reg[7]  ( .D(n1401), .CP(clk), .CD(n7935), .Q(z[7]) );
  CFD2XL \dout_reg[6]  ( .D(n1400), .CP(clk), .CD(n7935), .Q(z[6]) );
  CFD2XL \dout_reg[5]  ( .D(n1399), .CP(clk), .CD(n7935), .Q(z[5]) );
  CFD2XL \dout_reg[4]  ( .D(n1193), .CP(clk), .CD(n7935), .Q(z[4]) );
  CFD2XL \dout_reg[3]  ( .D(n1397), .CP(clk), .CD(n7935), .Q(z[3]) );
  CFD2XL \h0_1_reg[6]  ( .D(n933), .CP(clk), .CD(n7935), .Q(h0_1[6]), .QN(
        n8019) );
  CFD2XL \h0_1_reg[5]  ( .D(n930), .CP(clk), .CD(n7935), .Q(h0_1[5]), .QN(
        n8016) );
  CFD2XL \h0_1_reg[4]  ( .D(n927), .CP(clk), .CD(n7935), .Q(h0_1[4]), .QN(
        n8020) );
  CFD2XL \h0_0_reg[6]  ( .D(n934), .CP(clk), .CD(n7935), .Q(h0_0[6]) );
  CFD2XL \h0_0_reg[4]  ( .D(n928), .CP(clk), .CD(n7935), .Q(h0_0[4]) );
  CFD2XL \h0_0_reg[3]  ( .D(n1428), .CP(clk), .CD(n7935), .Q(h0_0[3]) );
  CFD2XL \h0_0_reg[2]  ( .D(n1337), .CP(clk), .CD(n7935), .Q(h0_0[2]) );
  CFD2XL \h0_0_reg[0]  ( .D(n1336), .CP(clk), .CD(n7935), .Q(h0_0[0]) );
  CFD2XL \out1_0_reg[1]  ( .D(N16), .CP(clk), .CD(n7935), .Q(out1_0[1]) );
  CFD2XL \out0_2_reg[63]  ( .D(n1121), .CP(clk), .CD(n7935), .Q(out0_2[63]), 
        .QN(n8011) );
  CFD2XL \out0_2_reg[62]  ( .D(n1122), .CP(clk), .CD(n7935), .Q(out0_2[62]), 
        .QN(n7938) );
  CFD2XL \out0_2_reg[61]  ( .D(n1123), .CP(clk), .CD(n7935), .Q(out0_2[61]), 
        .QN(n7940) );
  CFD2XL \out0_2_reg[60]  ( .D(n1124), .CP(clk), .CD(n7935), .Q(out0_2[60]), 
        .QN(n7943) );
  CFD2XL \out0_2_reg[55]  ( .D(n1129), .CP(clk), .CD(n7935), .Q(out0_2[55]), 
        .QN(n2648) );
  CFD2XL \out0_2_reg[53]  ( .D(n1131), .CP(clk), .CD(n7935), .Q(out0_2[53]), 
        .QN(n2640) );
  CFD2XL \out0_2_reg[52]  ( .D(n1132), .CP(clk), .CD(n7935), .Q(out0_2[52]), 
        .QN(n2635) );
  CFD2XL \out1_0_reg[2]  ( .D(N17), .CP(clk), .CD(n7935), .Q(out1_0[2]) );
  CFD2XL \out2_2_reg[63]  ( .D(n882), .CP(clk), .CD(n7935), .Q(out2_2[63]) );
  CFD2XL \out2_2_reg[61]  ( .D(n881), .CP(clk), .CD(n7935), .Q(out2_2[61]) );
  CFD2XL \out2_2_reg[56]  ( .D(n911), .CP(clk), .CD(n7935), .Q(out2_2[56]), 
        .QN(n7951) );
  CFD2XL \out1_0_reg[4]  ( .D(N19), .CP(clk), .CD(n7935), .Q(out1_0[4]) );
  CFD2XL \out2_2_reg[57]  ( .D(n877), .CP(clk), .CD(n7935), .Q(out2_2[57]), 
        .QN(n7949) );
  CFD2XL \acc_reg[39]  ( .D(n1032), .CP(clk), .CD(n7935), .Q(acc[39]), .QN(
        n7980) );
  CFD2XL \acc_reg[35]  ( .D(n1028), .CP(clk), .CD(n7935), .Q(acc[35]), .QN(
        n7988) );
  CFD2XL \acc_reg[51]  ( .D(n1044), .CP(clk), .CD(n7935), .Q(acc[51]), .QN(
        n7962) );
  CFD2XL \out1_0_reg[3]  ( .D(N18), .CP(clk), .CD(n7935), .Q(out1_0[3]) );
  CFD2XL \out2_2_reg[53]  ( .D(n879), .CP(clk), .CD(n7935), .Q(out2_2[53]), 
        .QN(n7957) );
  CFD2XL \acc_reg[49]  ( .D(n1042), .CP(clk), .CD(n7935), .Q(acc[49]), .QN(
        n7966) );
  CFD2XL \acc_reg[37]  ( .D(n1030), .CP(clk), .CD(n7935), .Q(acc[37]), .QN(
        n7984) );
  CFD2XL \acc_reg[53]  ( .D(n1293), .CP(clk), .CD(n7935), .Q(acc[53]), .QN(
        n7958) );
  CFD2XL \acc_reg[55]  ( .D(n1270), .CP(clk), .CD(n7935), .Q(acc[55]), .QN(
        n7954) );
  CFD2XL \out2_2_reg[45]  ( .D(n873), .CP(clk), .CD(n7935), .Q(out2_2[45]), 
        .QN(n7970) );
  CFD2XL \out2_2_reg[52]  ( .D(n908), .CP(clk), .CD(n7935), .Q(out2_2[52]), 
        .QN(n7959) );
  CFD2XL \out2_2_reg[37]  ( .D(n870), .CP(clk), .CD(n7935), .Q(out2_2[37]), 
        .QN(n7983) );
  CFD2XL \out2_2_reg[62]  ( .D(n1426), .CP(clk), .CD(n7935), .Q(out2_2[62]) );
  CFD2XL \out2_2_reg[47]  ( .D(n874), .CP(clk), .CD(n7935), .Q(out2_2[47]), 
        .QN(n7968) );
  CFD2XL \acc_reg[44]  ( .D(n1384), .CP(clk), .CD(n7935), .Q(acc[44]), .QN(
        n7973) );
  CFD2XL \acc_reg[36]  ( .D(n1029), .CP(clk), .CD(n7935), .Q(acc[36]), .QN(
        n7986) );
  CFD2XL \out2_2_reg[41]  ( .D(n862), .CP(clk), .CD(n7935), .Q(out2_2[41]), 
        .QN(n7977) );
  CFD2XL \acc_reg[61]  ( .D(n1054), .CP(clk), .CD(n7935), .Q(acc[61]), .QN(
        n7941) );
  CFD2XL \acc_reg[59]  ( .D(n1052), .CP(clk), .CD(n7935), .Q(acc[59]), .QN(
        n7946) );
  CFD2XL \acc_reg[57]  ( .D(n1050), .CP(clk), .CD(n7935), .Q(acc[57]), .QN(
        n7950) );
  CFD2XL \acc_reg[52]  ( .D(n1045), .CP(clk), .CD(n7935), .Q(acc[52]), .QN(
        n7960) );
  CFD2XL \out2_2_reg[59]  ( .D(n880), .CP(clk), .CD(n7935), .QN(n7945) );
  CFD2XL \out2_2_reg[60]  ( .D(n913), .CP(clk), .CD(n7935), .QN(n7942) );
  CFD2XL \acc_reg[62]  ( .D(n1331), .CP(clk), .CD(n7935), .Q(acc[62]), .QN(
        n7939) );
  CFD2XL \acc_reg[50]  ( .D(n1332), .CP(clk), .CD(n7935), .Q(acc[50]), .QN(
        n7964) );
  CFD2XL \acc_reg[42]  ( .D(n1035), .CP(clk), .CD(n7935), .Q(acc[42]), .QN(
        n7976) );
  CFD2XL \acc_reg[38]  ( .D(n1031), .CP(clk), .CD(n7935), .Q(acc[38]), .QN(
        n7982) );
  CFD2XL \acc_reg[56]  ( .D(n1049), .CP(clk), .CD(n7935), .Q(acc[56]), .QN(
        n7952) );
  CFD2XL \out2_2_reg[46]  ( .D(n906), .CP(clk), .CD(n7935), .Q(out2_2[46]), 
        .QN(n7969) );
  CFD2XL \acc_reg[60]  ( .D(n1427), .CP(clk), .CD(n7935), .Q(acc[60]), .QN(
        n7944) );
  CFD2XL \out2_2_reg[31]  ( .D(n851), .CP(clk), .CD(n7935), .Q(out2_2[31]), 
        .QN(n7994) );
  CFD2XL \out2_2_reg[49]  ( .D(n878), .CP(clk), .CD(n7935), .Q(out2_2[49]), 
        .QN(n7965) );
  CFD2XL \out2_2_reg[42]  ( .D(n904), .CP(clk), .CD(n7935), .Q(out2_2[42]), 
        .QN(n7975) );
  CFD2XL \out2_2_reg[38]  ( .D(n902), .CP(clk), .CD(n7935), .Q(out2_2[38]), 
        .QN(n7981) );
  CFD2XL \acc_reg[33]  ( .D(n1026), .CP(clk), .CD(n7935), .Q(acc[33]), .QN(
        n7991) );
  CFD2XL \out2_2_reg[58]  ( .D(n912), .CP(clk), .CD(n7935), .Q(out2_2[58]), 
        .QN(n7947) );
  CFD2XL \out2_2_reg[50]  ( .D(n905), .CP(clk), .CD(n7935), .Q(out2_2[50]), 
        .QN(n7963) );
  CFD2XL \out2_2_reg[48]  ( .D(n909), .CP(clk), .CD(n7935), .Q(out2_2[48]), 
        .QN(n7967) );
  CFD2XL \acc_reg[32]  ( .D(n1025), .CP(clk), .CD(n7935), .Q(acc[32]), .QN(
        n7993) );
  CFD2XL \out2_2_reg[34]  ( .D(n897), .CP(clk), .CD(n7935), .Q(out2_2[34]), 
        .QN(n7989) );
  CFD2XL \out2_2_reg[55]  ( .D(n875), .CP(clk), .CD(n7935), .Q(out2_2[55]), 
        .QN(n7953) );
  CFD2XL \out2_2_reg[39]  ( .D(n854), .CP(clk), .CD(n7935), .Q(out2_2[39]), 
        .QN(n7979) );
  CFD2XL \out2_2_reg[35]  ( .D(n859), .CP(clk), .CD(n7935), .Q(out2_2[35]), 
        .QN(n7987) );
  CFD2XL \out2_2_reg[32]  ( .D(n901), .CP(clk), .CD(n7935), .Q(out2_2[32]), 
        .QN(n7992) );
  CFD2XL \out2_2_reg[33]  ( .D(n866), .CP(clk), .CD(n7935), .Q(out2_2[33]), 
        .QN(n7990) );
  CFD2XL \out2_2_reg[36]  ( .D(n900), .CP(clk), .CD(n7935), .Q(out2_2[36]), 
        .QN(n7985) );
  CFD2XL \out1_0_reg[5]  ( .D(N20), .CP(clk), .CD(n7935), .Q(out1_0[5]) );
  CFD2XL \out2_2_reg[23]  ( .D(n853), .CP(clk), .CD(n7935), .Q(out2_2[23]), 
        .QN(n7998) );
  CFD2XL \out2_2_reg[20]  ( .D(n889), .CP(clk), .CD(n7935), .Q(out2_2[20]), 
        .QN(n7999) );
  CFD2XL \acc_reg[54]  ( .D(n1047), .CP(clk), .CD(n7935), .Q(acc[54]), .QN(
        n7956) );
  CFD2XL \out2_2_reg[29]  ( .D(n1292), .CP(clk), .CD(n7935), .Q(out2_2[29]), 
        .QN(n7995) );
  CFD2XL \out2_2_reg[51]  ( .D(n1383), .CP(clk), .CD(n7935), .Q(out2_2[51]), 
        .QN(n7961) );
  CFD2XL \out2_2_reg[15]  ( .D(n852), .CP(clk), .CD(n7935), .Q(out2_2[15]), 
        .QN(n8002) );
  CFD2XL \acc_reg[58]  ( .D(n1382), .CP(clk), .CD(n7935), .Q(acc[58]), .QN(
        n7948) );
  CFD2XL \out2_2_reg[54]  ( .D(n910), .CP(clk), .CD(n7935), .Q(out2_2[54]), 
        .QN(n7955) );
  CFD2XL \out2_2_reg[17]  ( .D(n864), .CP(clk), .CD(n7935), .Q(out2_2[17]), 
        .QN(n8000) );
  CFD2XL \out2_2_reg[16]  ( .D(n891), .CP(clk), .CD(n7935), .Q(out2_2[16]), 
        .QN(n8001) );
  CFD2XL \out2_2_reg[40]  ( .D(n903), .CP(clk), .CD(n7935), .Q(out2_2[40]), 
        .QN(n7978) );
  CFD2XL \out2_2_reg[44]  ( .D(n907), .CP(clk), .CD(n7935), .Q(out2_2[44]), 
        .QN(n7972) );
  CFD2XL \out2_2_reg[43]  ( .D(n1340), .CP(clk), .CD(n7935), .Q(out2_2[43]), 
        .QN(n7974) );
  CFD2XL \out2_2_reg[13]  ( .D(n867), .CP(clk), .CD(n7935), .Q(out2_2[13]), 
        .QN(n8003) );
  CFD2XL \out2_2_reg[25]  ( .D(n1362), .CP(clk), .CD(n7935), .Q(out2_2[25]), 
        .QN(n7997) );
  CFD4XL \acc_reg[45]  ( .D(n1365), .CP(clk), .SD(n7935), .Q(n7971), .QN(
        acc[45]) );
  CFD2X1 \acc_reg[28]  ( .D(n1370), .CP(clk), .CD(n7935), .Q(acc[28]), .QN(
        n7996) );
  CFD3QX1 cmd2_en_2_reg ( .D(n1186), .CP(clk), .CD(1'b1), .SD(1'b1), .Q(
        cmd2_en_2) );
  CFD2XL \out1_0_reg[25]  ( .D(N40), .CP(clk), .CD(n7935), .Q(out1_0[25]) );
  CFD4X1 \q0_reg[4]  ( .D(n7857), .CP(clk), .SD(n7935), .Q(n7852), .QN(q0[4])
         );
  CFD4X2 \q0_reg[22]  ( .D(n7848), .CP(clk), .SD(n7935), .QN(q0[22]) );
  CFD2X1 \out0_2_reg[51]  ( .D(n1435), .CP(clk), .CD(n7935), .Q(out0_2[51]), 
        .QN(n2650) );
  CFD2X1 \out0_2_reg[49]  ( .D(n1446), .CP(clk), .CD(n7935), .Q(out0_2[49]), 
        .QN(n2639) );
  CFD2X1 \out0_2_reg[50]  ( .D(n1447), .CP(clk), .CD(n7935), .Q(out0_2[50]), 
        .QN(n2634) );
  CFD2X1 \out0_2_reg[56]  ( .D(n1394), .CP(clk), .CD(n7935), .Q(out0_2[56]), 
        .QN(n2641) );
  CFD2X1 \out0_2_reg[36]  ( .D(n1395), .CP(clk), .CD(n7935), .Q(out0_2[36]), 
        .QN(n2644) );
  CFD2X1 \out0_2_reg[57]  ( .D(n1396), .CP(clk), .CD(n7935), .Q(out0_2[57]), 
        .QN(n2636) );
  CFD2X1 \out0_2_reg[46]  ( .D(n1449), .CP(clk), .CD(n7935), .Q(out0_2[46]), 
        .QN(n2632) );
  CFD2X1 \out0_2_reg[48]  ( .D(n1391), .CP(clk), .CD(n7935), .Q(out0_2[48]), 
        .QN(n2633) );
  CFD2X1 \out0_2_reg[42]  ( .D(n1341), .CP(clk), .CD(n7935), .Q(out0_2[42]), 
        .QN(n2631) );
  CFD2X1 \out0_2_reg[59]  ( .D(n1386), .CP(clk), .CD(n7935), .Q(out0_2[59]), 
        .QN(n2637) );
  CFD2X1 \out0_2_reg[39]  ( .D(n1338), .CP(clk), .CD(n7935), .Q(out0_2[39]), 
        .QN(n2638) );
  CFD2X1 \out0_2_reg[37]  ( .D(n1441), .CP(clk), .CD(n7935), .Q(out0_2[37]), 
        .QN(n2649) );
  CFD2X1 \out0_2_reg[38]  ( .D(n1438), .CP(clk), .CD(n7935), .Q(out0_2[38]), 
        .QN(n2643) );
  CFD2X1 \out0_2_reg[34]  ( .D(n1342), .CP(clk), .CD(n7935), .Q(out0_2[34]), 
        .QN(n2642) );
  CFD2X1 \out0_2_reg[44]  ( .D(n1339), .CP(clk), .CD(n7935), .Q(out0_2[44]), 
        .QN(n2645) );
  CFD2X1 \out0_2_reg[16]  ( .D(n1279), .CP(clk), .CD(n7935), .Q(out0_2[16]), 
        .QN(n2653) );
  CFD2X1 \out0_2_reg[17]  ( .D(n1440), .CP(clk), .CD(n7935), .Q(out0_2[17]), 
        .QN(n2654) );
  CFD2X1 \out0_2_reg[18]  ( .D(n1530), .CP(clk), .CD(n7935), .Q(out0_2[18]), 
        .QN(n2652) );
  CFD2X1 \out0_2_reg[28]  ( .D(n1278), .CP(clk), .CD(n7935), .Q(out0_2[28]), 
        .QN(n2646) );
  CFD2X1 \out0_2_reg[29]  ( .D(n1389), .CP(clk), .CD(n7935), .Q(out0_2[29]), 
        .QN(n2655) );
  CFD2X1 \out0_2_reg[30]  ( .D(n1450), .CP(clk), .CD(n7935), .Q(out0_2[30]), 
        .QN(n2647) );
  CFD2X1 \out0_2_reg[21]  ( .D(n1364), .CP(clk), .CD(n7935), .Q(out0_2[21]), 
        .QN(n2651) );
  CFD2X1 \out0_2_reg[20]  ( .D(n1363), .CP(clk), .CD(n7935), .Q(out0_2[20]), 
        .QN(n2630) );
  CFD2X1 \out0_2_reg[0]  ( .D(n1184), .CP(clk), .CD(n7935), .Q(out0_2[0]), 
        .QN(n2684) );
  CFD2QX4 \h0_reg[5]  ( .D(n932), .CP(clk), .CD(n7935), .Q(h0[5]) );
  CFD2QX4 \h0_reg[1]  ( .D(n920), .CP(clk), .CD(n7935), .Q(h0[1]) );
  CFD2X1 \acc_reg[0]  ( .D(n1272), .CP(clk), .CD(n7935), .Q(acc[0]), .QN(n8010) );
  CFD2X1 \acc_reg[2]  ( .D(n1282), .CP(clk), .CD(n7935), .Q(acc[2]), .QN(n8008) );
  CFD2X1 \acc_reg[8]  ( .D(n1001), .CP(clk), .CD(n7935), .Q(acc[8]), .QN(n8007) );
  CFD2X1 \acc_reg[9]  ( .D(n1002), .CP(clk), .CD(n7935), .Q(acc[9]), .QN(n8006) );
  CFD2X1 \acc_reg[17]  ( .D(n1010), .CP(clk), .CD(n7935), .Q(acc[17]), .QN(
        n8014) );
  CFD2X1 \acc_reg[16]  ( .D(n1009), .CP(clk), .CD(n7935), .Q(acc[16]), .QN(
        n8015) );
  CFD2X1 \acc_reg[12]  ( .D(n1005), .CP(clk), .CD(n7935), .Q(acc[12]), .QN(
        n8017) );
  CFD2X1 \acc_reg[11]  ( .D(n1004), .CP(clk), .CD(n7935), .Q(acc[11]), .QN(
        n8018) );
  CFD2X1 \acc_reg[10]  ( .D(n1003), .CP(clk), .CD(n7935), .Q(acc[10]), .QN(
        n8005) );
  CFD2X1 \acc_reg[1]  ( .D(n1334), .CP(clk), .CD(n7935), .Q(acc[1]), .QN(n8009) );
  CFD1QXL cmd1_en_2_reg ( .D(n1187), .CP(clk), .Q(cmd1_en_2) );
  CFD2X1 \out0_2_reg[45]  ( .D(n1333), .CP(clk), .CD(n7935), .Q(out0_2[45]), 
        .QN(n2629) );
  CFD2QX4 \h0_reg[17]  ( .D(n946), .CP(clk), .CD(n7935), .Q(h0[17]) );
  CFD2QX4 \h0_reg[20]  ( .D(n949), .CP(clk), .CD(n7935), .Q(h0[20]) );
  CFD2QX4 \h0_reg[23]  ( .D(n952), .CP(clk), .CD(n7935), .Q(h0[23]) );
  CFD4X4 \h0_reg[12]  ( .D(n7854), .CP(clk), .SD(n7935), .QN(h0[12]) );
  CFD1QX1 cmd0_en_2_reg ( .D(n1188), .CP(clk), .Q(cmd0_en_2) );
  CFD2QX4 \h0_reg[24]  ( .D(n2905), .CP(clk), .CD(n7935), .Q(h0[24]) );
  CFD2QX4 \h0_reg[2]  ( .D(n923), .CP(clk), .CD(n7935), .Q(h0[2]) );
  CFD2QX4 \h0_reg[3]  ( .D(n2893), .CP(clk), .CD(n7935), .Q(h0[3]) );
  CFD2QX4 \h0_reg[18]  ( .D(n2902), .CP(clk), .CD(n7935), .Q(h0[18]) );
  CFD2QX4 \h0_reg[27]  ( .D(n2908), .CP(clk), .CD(n7935), .Q(h0[27]) );
  CFD2QX4 \h0_reg[22]  ( .D(n2904), .CP(clk), .CD(n7935), .Q(h0[22]) );
  CFD2QX4 \h0_reg[29]  ( .D(n2909), .CP(clk), .CD(n7935), .Q(h0[29]) );
  CFD2QX4 \h0_reg[28]  ( .D(n957), .CP(clk), .CD(n7935), .Q(h0[28]) );
  CFD2QX4 \h0_reg[10]  ( .D(n2896), .CP(clk), .CD(n7935), .Q(h0[10]) );
  CFD2QX4 \h0_reg[31]  ( .D(n2910), .CP(clk), .CD(n7935), .Q(h0[31]) );
  CFD2QX4 \h0_reg[11]  ( .D(n940), .CP(clk), .CD(n7935), .Q(h0[11]) );
  CFD2QX4 \h0_reg[30]  ( .D(n959), .CP(clk), .CD(n7935), .Q(h0[30]) );
  CFD2QX4 \h0_reg[8]  ( .D(n2895), .CP(clk), .CD(n7935), .Q(h0[8]) );
  CFD2QX4 \h0_reg[19]  ( .D(n2903), .CP(clk), .CD(n7935), .Q(h0[19]) );
  CFD2QX4 \h0_reg[25]  ( .D(n2906), .CP(clk), .CD(n7935), .Q(h0[25]) );
  CFD2QX4 \h0_reg[26]  ( .D(n2907), .CP(clk), .CD(n7935), .Q(h0[26]) );
  CFD2QX4 \h0_reg[15]  ( .D(n2900), .CP(clk), .CD(n7935), .Q(h0[15]) );
  CFD2QX4 \h0_reg[16]  ( .D(n2901), .CP(clk), .CD(n7935), .Q(h0[16]) );
  CFD2QX4 \h0_reg[13]  ( .D(n2898), .CP(clk), .CD(n7935), .Q(h0[13]) );
  CFD2QX4 \h0_reg[7]  ( .D(n2894), .CP(clk), .CD(n7935), .Q(h0[7]) );
  CFD2QX4 \h0_reg[14]  ( .D(n2899), .CP(clk), .CD(n7935), .Q(h0[14]) );
  CFD2QX2 \q0_reg[0]  ( .D(n1277), .CP(clk), .CD(n7935), .Q(q0[0]) );
  CFD2QX1 \h0_reg[4]  ( .D(n929), .CP(clk), .CD(n7935), .Q(h0[4]) );
  CFD2QX2 \q0_reg[28]  ( .D(n2943), .CP(clk), .CD(n7935), .Q(q0[28]) );
  CFD2X1 \q0_reg[20]  ( .D(n1271), .CP(clk), .CD(n7935), .Q(n2464), .QN(n2465)
         );
  CFD2QX2 \q0_reg[6]  ( .D(n1273), .CP(clk), .CD(n7935), .Q(q0[6]) );
  CFD2QX1 \h0_reg[21]  ( .D(n950), .CP(clk), .CD(n7935), .Q(h0[21]) );
  CFD2QX2 \h0_reg[0]  ( .D(n917), .CP(clk), .CD(n7935), .Q(h0[0]) );
  CND2X1 U1292 ( .A(n1266), .B(n5340), .Z(n1568) );
  CNIVXL U1293 ( .A(n6110), .Z(n1222) );
  CND2X2 U1294 ( .A(n5003), .B(n5004), .Z(n5602) );
  CND2X2 U1295 ( .A(n1223), .B(n2459), .Z(n6277) );
  CND2X2 U1296 ( .A(n2458), .B(n2457), .Z(n1223) );
  CND2X2 U1297 ( .A(n5939), .B(n1224), .Z(n6049) );
  COND1X2 U1298 ( .A(n5938), .B(n5937), .C(n5936), .Z(n1224) );
  CNR2X2 U1299 ( .A(n5985), .B(n6293), .Z(n5869) );
  COND1X2 U1300 ( .A(n1225), .B(n5600), .C(n5599), .Z(n5676) );
  CNR2X2 U1301 ( .A(n5597), .B(n1584), .Z(n1225) );
  CIVX1 U1302 ( .A(q0[11]), .Z(n2606) );
  CND2X1 U1303 ( .A(n2450), .B(n6169), .Z(n2505) );
  CENX2 U1304 ( .A(n6149), .B(n5935), .Z(n6169) );
  CENX2 U1305 ( .A(n6417), .B(h0[23]), .Z(n2283) );
  CENX2 U1306 ( .A(n5978), .B(n5865), .Z(n5945) );
  CNR2X2 U1307 ( .A(n7003), .B(n7018), .Z(n7035) );
  CNR2X2 U1308 ( .A(n6272), .B(n6271), .Z(n7003) );
  CND2X1 U1309 ( .A(n2407), .B(n6277), .Z(n6263) );
  CENX1 U1310 ( .A(n6220), .B(n6171), .Z(n2407) );
  CNIVXL U1311 ( .A(n7205), .Z(n1226) );
  CND2IX2 U1312 ( .B(n2294), .A(n2657), .Z(n4965) );
  CND2X4 U1313 ( .A(n4965), .B(n4964), .Z(n5223) );
  CENX2 U1314 ( .A(n5209), .B(n2466), .Z(n5210) );
  CND2X2 U1315 ( .A(n1230), .B(n1227), .Z(n2466) );
  CND2X2 U1316 ( .A(n1229), .B(n1228), .Z(n1227) );
  CIVX2 U1317 ( .A(n6702), .Z(n1228) );
  CIVX2 U1318 ( .A(n4946), .Z(n1229) );
  CND2IX1 U1319 ( .B(n6703), .A(n1231), .Z(n1230) );
  CIVX2 U1320 ( .A(n5096), .Z(n1231) );
  CNR2X2 U1321 ( .A(n5378), .B(n5379), .Z(n5381) );
  CNIVX4 U1322 ( .A(n6703), .Z(n6473) );
  CNIVX1 U1323 ( .A(n6530), .Z(n6474) );
  CNIVX1 U1324 ( .A(h0[3]), .Z(n1232) );
  CENX1 U1325 ( .A(q0[3]), .B(q0[4]), .Z(n3350) );
  COND2X2 U1326 ( .A(n2571), .B(n4996), .C(n2488), .D(n5578), .Z(n5591) );
  CNR2X2 U1327 ( .A(n5592), .B(n5591), .Z(n5590) );
  CENX2 U1328 ( .A(n1233), .B(n2345), .Z(n5365) );
  CENX2 U1329 ( .A(n4977), .B(n4976), .Z(n1233) );
  CENX2 U1330 ( .A(n4880), .B(n4879), .Z(n4743) );
  COND2X2 U1331 ( .A(n6703), .B(n4756), .C(n2515), .D(n4796), .Z(n4880) );
  CIVX2 U1332 ( .A(n2560), .Z(n2569) );
  CND2X2 U1333 ( .A(n1235), .B(n1234), .Z(n6874) );
  CND2X2 U1334 ( .A(n1237), .B(n6853), .Z(n1234) );
  COND1X2 U1335 ( .A(n6853), .B(n1237), .C(n6852), .Z(n1235) );
  CENX1 U1336 ( .A(n1237), .B(n1236), .Z(n6833) );
  CENX1 U1337 ( .A(n6853), .B(n6852), .Z(n1236) );
  CENX1 U1338 ( .A(n6849), .B(n6801), .Z(n1237) );
  COND1X2 U1339 ( .A(n5476), .B(n5475), .C(n5474), .Z(n5478) );
  COND2X2 U1340 ( .A(n6405), .B(n2294), .C(n7114), .D(n6470), .Z(n6516) );
  CNIVX4 U1341 ( .A(n4432), .Z(n1238) );
  COND2X2 U1342 ( .A(n7203), .B(n4736), .C(n4715), .D(n7217), .Z(n4751) );
  COND1X2 U1343 ( .A(n6331), .B(n6332), .C(n6330), .Z(n6334) );
  CND2X1 U1344 ( .A(n4981), .B(n5363), .Z(n4982) );
  CENX2 U1345 ( .A(n2098), .B(n4908), .Z(n5363) );
  CIVX4 U1346 ( .A(n6972), .Z(n4662) );
  CIVXL U1347 ( .A(n7011), .Z(n7490) );
  COAN1X1 U1348 ( .A(n7011), .B(n5504), .C(n7496), .Z(n5513) );
  CND2X1 U1349 ( .A(n1240), .B(n1239), .Z(n5806) );
  CND2XL U1350 ( .A(n5721), .B(n5722), .Z(n1239) );
  COND1XL U1351 ( .A(n5722), .B(n5721), .C(n5720), .Z(n1240) );
  CENX2 U1352 ( .A(n1241), .B(n5721), .Z(n5683) );
  CENX2 U1353 ( .A(n5722), .B(n5720), .Z(n1241) );
  CENX1 U1354 ( .A(n6647), .B(h0[18]), .Z(n5565) );
  CENX1 U1355 ( .A(n5637), .B(n5638), .Z(n5041) );
  COND1X2 U1356 ( .A(n5037), .B(n5038), .C(n5036), .Z(n5638) );
  CND2X1 U1357 ( .A(n2307), .B(n1913), .Z(n1914) );
  CENX1 U1358 ( .A(n6810), .B(n1242), .Z(n6815) );
  CENX2 U1359 ( .A(n6812), .B(n6811), .Z(n1242) );
  CND2X2 U1360 ( .A(n1245), .B(n1243), .Z(n2536) );
  CIVX2 U1361 ( .A(n5838), .Z(n1243) );
  CND2X2 U1362 ( .A(n1244), .B(n5753), .Z(n5838) );
  COND1X2 U1363 ( .A(n5751), .B(n5752), .C(n5750), .Z(n1244) );
  CIVX2 U1364 ( .A(n5840), .Z(n1245) );
  CIVX2 U1365 ( .A(n1246), .Z(n2661) );
  COND1X2 U1366 ( .A(n7433), .B(n7235), .C(n1247), .Z(n1246) );
  CANR1X2 U1367 ( .A(n7234), .B(n1249), .C(n1248), .Z(n1247) );
  COND1X2 U1368 ( .A(n7233), .B(n7449), .C(n7232), .Z(n1248) );
  CND2X2 U1369 ( .A(n7166), .B(n7165), .Z(n7449) );
  CIVX2 U1370 ( .A(n7263), .Z(n7234) );
  CND2X2 U1371 ( .A(n7162), .B(n7161), .Z(n7263) );
  CND2X2 U1372 ( .A(n7264), .B(n1249), .Z(n7235) );
  CNR2IX2 U1373 ( .B(n1250), .A(n7191), .Z(n1249) );
  CNR2X2 U1374 ( .A(n7165), .B(n7166), .Z(n7191) );
  CIVX2 U1375 ( .A(n7233), .Z(n1250) );
  CNR2X2 U1376 ( .A(n7187), .B(n7186), .Z(n7233) );
  CND2X2 U1377 ( .A(n1252), .B(n1251), .Z(n7264) );
  CIVX2 U1378 ( .A(n7162), .Z(n1251) );
  CIVX2 U1379 ( .A(n7130), .Z(n1252) );
  CND2X2 U1380 ( .A(n7157), .B(n7156), .Z(n7433) );
  CENXL U1381 ( .A(n7494), .B(n1253), .Z(N39) );
  CAN2XL U1382 ( .A(n2297), .B(n6381), .Z(n1253) );
  CENXL U1383 ( .A(n4657), .B(n2255), .Z(N36) );
  COND2X1 U1384 ( .A(n3493), .B(n7537), .C(n3492), .D(n5160), .Z(n3508) );
  CND2X1 U1385 ( .A(n3496), .B(n3495), .Z(n1593) );
  CND2X1 U1386 ( .A(n4638), .B(n4637), .Z(n7528) );
  CENX1 U1387 ( .A(n3802), .B(n3430), .Z(n3747) );
  COND1X1 U1388 ( .A(n3801), .B(n3802), .C(n3800), .Z(n3804) );
  COND1X1 U1389 ( .A(n3533), .B(n3535), .C(n3532), .Z(n3421) );
  CENX1 U1390 ( .A(n3533), .B(n3532), .Z(n3534) );
  CENXL U1391 ( .A(n7475), .B(n1254), .Z(N47) );
  CAN2XL U1392 ( .A(n5079), .B(n7309), .Z(n1254) );
  CND2X1 U1393 ( .A(n4464), .B(n4465), .Z(n4405) );
  CND2X4 U1394 ( .A(n4402), .B(n4401), .Z(n4465) );
  CANR1X1 U1395 ( .A(n7151), .B(n2438), .C(n7149), .Z(n2541) );
  CND2X1 U1396 ( .A(n2403), .B(n6474), .Z(n6475) );
  COND1X1 U1397 ( .A(n6530), .B(n2403), .C(n6531), .Z(n6476) );
  CIVX8 U1398 ( .A(n3615), .Z(n6118) );
  CENX1 U1399 ( .A(n3458), .B(n3457), .Z(n3472) );
  CANR5CX1 U1400 ( .A(n2033), .B(n3560), .C(n3559), .Z(n1970) );
  CENX1 U1401 ( .A(n3597), .B(n3596), .Z(n3599) );
  COND1XL U1402 ( .A(n3468), .B(n3467), .C(n3466), .Z(n1255) );
  CENX1 U1403 ( .A(n3551), .B(n3536), .Z(n3739) );
  CND2X1 U1404 ( .A(n3431), .B(n3433), .Z(n3374) );
  CENX1 U1405 ( .A(n3608), .B(n2656), .Z(n3609) );
  CND2X1 U1406 ( .A(n3608), .B(n2656), .Z(n3582) );
  COND1X1 U1407 ( .A(n3574), .B(n3572), .C(n3573), .Z(n3516) );
  CENX2 U1408 ( .A(n5372), .B(n1256), .Z(n5382) );
  CEOX2 U1409 ( .A(n5370), .B(n5371), .Z(n1256) );
  CND2IX2 U1410 ( .B(n4818), .A(n4820), .Z(n4821) );
  COND1X2 U1411 ( .A(n2559), .B(n5389), .C(n5387), .Z(n5391) );
  COND1X1 U1412 ( .A(n5528), .B(n5527), .C(n5526), .Z(n1257) );
  COND1X1 U1413 ( .A(n5528), .B(n5527), .C(n5526), .Z(n2404) );
  CIVXL U1414 ( .A(n5061), .Z(n5058) );
  CND2X1 U1415 ( .A(n5945), .B(n5946), .Z(n5948) );
  CENX1 U1416 ( .A(n2363), .B(n5330), .Z(n1258) );
  COND1XL U1417 ( .A(n6983), .B(n6984), .C(n6982), .Z(n6986) );
  COND2X2 U1418 ( .A(n4538), .B(n2295), .C(n7114), .D(n5169), .Z(n5299) );
  CAOR1XL U1419 ( .A(n7218), .B(n1226), .C(n7216), .Z(n7225) );
  CENXL U1420 ( .A(n6118), .B(h0[1]), .Z(n3614) );
  CENXL U1421 ( .A(n5793), .B(h0[1]), .Z(n3680) );
  CENX1 U1422 ( .A(n6769), .B(h0[19]), .Z(n6145) );
  COND2XL U1423 ( .A(n7853), .B(n7126), .C(n7124), .D(n4678), .Z(n1259) );
  CIVXL U1424 ( .A(n5512), .Z(n1260) );
  CNR2XL U1425 ( .A(n6280), .B(n2286), .Z(n1261) );
  CMXI2XL U1426 ( .A0(n5923), .A1(q[7]), .S(n7682), .Z(n2668) );
  CENX2 U1427 ( .A(q0[1]), .B(q0[2]), .Z(n4492) );
  CIVX2 U1428 ( .A(n5574), .Z(n5575) );
  CIVDX4 U1429 ( .A(q0[19]), .Z0(n4390), .Z1(n6769) );
  CNIVXL U1430 ( .A(n6211), .Z(n1262) );
  CENX2 U1431 ( .A(n2583), .B(h0[20]), .Z(n4958) );
  CNIVX1 U1432 ( .A(n4751), .Z(n2468) );
  CENX2 U1433 ( .A(n6769), .B(h0[7]), .Z(n5097) );
  CENX1 U1434 ( .A(n6415), .B(n6509), .Z(n6535) );
  COND1X2 U1435 ( .A(n6414), .B(n2396), .C(n6413), .Z(n6509) );
  COND1X1 U1436 ( .A(n6632), .B(n6633), .C(n6631), .Z(n6635) );
  CND3X1 U1437 ( .A(n2371), .B(n2372), .C(n2373), .Z(n6632) );
  CENX2 U1438 ( .A(h0[8]), .B(n7092), .Z(n4774) );
  COND1X2 U1439 ( .A(n5807), .B(n5806), .C(n5805), .Z(n5809) );
  CIVX2 U1440 ( .A(n4962), .Z(n1263) );
  COND2X1 U1441 ( .A(n7126), .B(n5756), .C(n2433), .D(n5798), .Z(n1264) );
  CENX1 U1442 ( .A(n6570), .B(n6533), .Z(n1265) );
  CENX1 U1443 ( .A(n6570), .B(n6533), .Z(n6908) );
  CENX2 U1444 ( .A(n6417), .B(h0[20]), .Z(n4661) );
  CND2X4 U1445 ( .A(n6065), .B(n6064), .Z(n6135) );
  CEO3X2 U1446 ( .A(n4751), .B(n4750), .C(n4749), .Z(n4912) );
  CND2X2 U1447 ( .A(n5389), .B(n2559), .Z(n5390) );
  COND1X2 U1448 ( .A(n5083), .B(n5081), .C(n5080), .Z(n4842) );
  CENX2 U1449 ( .A(n5856), .B(n5757), .Z(n5880) );
  CND2XL U1450 ( .A(n6046), .B(n6045), .Z(n6047) );
  COND2XL U1451 ( .A(n6870), .B(n5167), .C(n6829), .D(n5166), .Z(n1266) );
  CND2X2 U1452 ( .A(n7290), .B(n7318), .Z(n7267) );
  CFA1X2 U1453 ( .A(n6167), .B(n6166), .CI(n6165), .CO(n6219), .S(n6134) );
  COND2XL U1454 ( .A(n6974), .B(n5634), .C(n5692), .D(n6972), .Z(n1267) );
  CND2XL U1455 ( .A(n4824), .B(n4818), .Z(n4706) );
  CIVX8 U1456 ( .A(n7867), .Z(n7134) );
  CNIVX3 U1457 ( .A(out1_0[40]), .Z(n1269) );
  CNIVX1 U1458 ( .A(n1269), .Z(n1268) );
  COND3X2 U1459 ( .A(n2652), .B(n2685), .C(n2239), .D(n2242), .Z(n1011) );
  CNIVX1 U1460 ( .A(n1048), .Z(n1270) );
  CNIVX1 U1461 ( .A(n2897), .Z(n1271) );
  CNIVX1 U1462 ( .A(n993), .Z(n1272) );
  CNIVX1 U1463 ( .A(n2941), .Z(n1273) );
  CNIVX1 U1464 ( .A(n2725), .Z(n1274) );
  CNIVX3 U1465 ( .A(out1_0[24]), .Z(n1276) );
  CNIVX1 U1466 ( .A(n1276), .Z(n1275) );
  CNIVX1 U1467 ( .A(n961), .Z(n1277) );
  COND3X2 U1468 ( .A(n2685), .B(n2014), .C(n2015), .D(n2017), .Z(n998) );
  COND3X2 U1469 ( .A(n2685), .B(n2226), .C(n2227), .D(n2230), .Z(n999) );
  COND3X2 U1470 ( .A(n2685), .B(n2231), .C(n2232), .D(n2234), .Z(n1000) );
  COND3X2 U1471 ( .A(n2685), .B(n2235), .C(n2236), .D(n2238), .Z(n1006) );
  COND3X2 U1472 ( .A(n2685), .B(n2079), .C(n2080), .D(n2082), .Z(n1008) );
  CNIVX1 U1473 ( .A(n1156), .Z(n1278) );
  CNIVX1 U1474 ( .A(n1168), .Z(n1279) );
  CNIVX1 U1475 ( .A(n1041), .Z(n1280) );
  CNIVX1 U1476 ( .A(n1335), .Z(n1281) );
  COND3X2 U1477 ( .A(n2685), .B(n1900), .C(n1901), .D(n1903), .Z(n996) );
  CNIVX1 U1478 ( .A(n995), .Z(n1282) );
  CNIVX1 U1479 ( .A(n1013), .Z(n1283) );
  CMXI2X2 U1480 ( .A0(n1284), .A1(q[22]), .S(n7682), .Z(n7848) );
  CNIVX1 U1481 ( .A(q0[22]), .Z(n1284) );
  CNIVX2 U1482 ( .A(n1022), .Z(n1285) );
  CNIVX1 U1483 ( .A(n1287), .Z(n1286) );
  CNIVXL U1484 ( .A(n1023), .Z(n1287) );
  CNIVX1 U1485 ( .A(n2862), .Z(n1288) );
  CNIVX2 U1486 ( .A(n1014), .Z(n1289) );
  CNIVX1 U1487 ( .A(n2863), .Z(n1290) );
  CNIVX1 U1488 ( .A(n2864), .Z(n1291) );
  CNIVX1 U1489 ( .A(n868), .Z(n1292) );
  COND3X2 U1490 ( .A(n2685), .B(n2191), .C(n2192), .D(n2195), .Z(n1047) );
  CNIVX1 U1491 ( .A(n1046), .Z(n1293) );
  CNIVX1 U1492 ( .A(n2666), .Z(n1294) );
  CNIVX3 U1493 ( .A(out1_0[38]), .Z(n1296) );
  CNIVX1 U1494 ( .A(n1296), .Z(n1295) );
  CNIVX1 U1495 ( .A(N15), .Z(n1297) );
  CNR2IXL U1496 ( .B(n7538), .A(n7537), .Z(N15) );
  CNIVX3 U1497 ( .A(cmd0_0[1]), .Z(n1299) );
  CNIVX1 U1498 ( .A(n1299), .Z(n1298) );
  CNIVX3 U1499 ( .A(out1_0[28]), .Z(n1301) );
  CNIVX1 U1500 ( .A(n1301), .Z(n1300) );
  CNIVX3 U1501 ( .A(out1_0[62]), .Z(n1303) );
  CNIVX1 U1502 ( .A(n1303), .Z(n1302) );
  CNIVX3 U1503 ( .A(out1_0[46]), .Z(n1305) );
  CNIVX1 U1504 ( .A(n1305), .Z(n1304) );
  CNIVX3 U1505 ( .A(cmd0_1[0]), .Z(n1307) );
  CNIVX1 U1506 ( .A(n1307), .Z(n1306) );
  CNIVX3 U1507 ( .A(out1_0[31]), .Z(n1309) );
  CNIVX1 U1508 ( .A(n1309), .Z(n1308) );
  CNIVX3 U1509 ( .A(out1_0[1]), .Z(n1311) );
  CNIVX1 U1510 ( .A(n1311), .Z(n1310) );
  CNIVX3 U1511 ( .A(out1_0[37]), .Z(n1313) );
  CNIVX1 U1512 ( .A(n1313), .Z(n1312) );
  CNIVX3 U1513 ( .A(cmd0_0[0]), .Z(n1315) );
  CNIVX1 U1514 ( .A(n1315), .Z(n1314) );
  CNIVX1 U1515 ( .A(n2942), .Z(n1316) );
  CNIVX3 U1516 ( .A(out1_0[36]), .Z(n1318) );
  CNIVX1 U1517 ( .A(n1318), .Z(n1317) );
  CNIVX3 U1518 ( .A(out1_0[33]), .Z(n1320) );
  CNIVX1 U1519 ( .A(n1320), .Z(n1319) );
  CNIVX3 U1520 ( .A(out1_0[29]), .Z(n1322) );
  CNIVX1 U1521 ( .A(n1322), .Z(n1321) );
  CNIVX3 U1522 ( .A(out1_0[61]), .Z(n1324) );
  CNIVX1 U1523 ( .A(n1324), .Z(n1323) );
  CNIVX3 U1524 ( .A(out1_0[39]), .Z(n1326) );
  CNIVX1 U1525 ( .A(n1326), .Z(n1325) );
  CNIVX3 U1526 ( .A(out1_0[42]), .Z(n1328) );
  CNIVX1 U1527 ( .A(n1328), .Z(n1327) );
  CNIVX3 U1528 ( .A(out1_0[13]), .Z(n1330) );
  CNIVX1 U1529 ( .A(n1330), .Z(n1329) );
  CNIVX1 U1530 ( .A(n1055), .Z(n1331) );
  CNIVX2 U1531 ( .A(n1043), .Z(n1332) );
  CMXI2XL U1532 ( .A0(h0[12]), .A1(h[12]), .S(pushin), .Z(n7854) );
  CNIVX1 U1533 ( .A(n1139), .Z(n1333) );
  CNIVX1 U1534 ( .A(n994), .Z(n1334) );
  CNIVX1 U1535 ( .A(cmd0[0]), .Z(n1335) );
  CNIVX1 U1536 ( .A(n916), .Z(n1336) );
  CNIVX1 U1537 ( .A(n922), .Z(n1337) );
  CNIVX1 U1538 ( .A(n1145), .Z(n1338) );
  CNIVX1 U1539 ( .A(n1140), .Z(n1339) );
  CNIVX1 U1540 ( .A(n872), .Z(n1340) );
  CNIVX1 U1541 ( .A(n1142), .Z(n1341) );
  CNIVX1 U1542 ( .A(n1150), .Z(n1342) );
  CNIVX1 U1543 ( .A(n1027), .Z(n1343) );
  COND3X2 U1544 ( .A(n2654), .B(n2685), .C(n3325), .D(n3324), .Z(n1010) );
  CNIVX1 U1545 ( .A(n1345), .Z(n1344) );
  CNIVXL U1546 ( .A(n1039), .Z(n1345) );
  COND3XL U1547 ( .A(n2685), .B(n2632), .C(n3241), .D(n3240), .Z(n1039) );
  CNIVX3 U1548 ( .A(out1_0[19]), .Z(n1347) );
  CNIVX1 U1549 ( .A(n1347), .Z(n1346) );
  CNIVX3 U1550 ( .A(out1_0[34]), .Z(n1349) );
  CNIVX1 U1551 ( .A(n1349), .Z(n1348) );
  CNIVX3 U1552 ( .A(out1_0[35]), .Z(n1351) );
  CNIVX1 U1553 ( .A(n1351), .Z(n1350) );
  CNIVX3 U1554 ( .A(out1_0[18]), .Z(n1353) );
  CNIVX1 U1555 ( .A(n1353), .Z(n1352) );
  CNIVX1 U1556 ( .A(n2946), .Z(n1354) );
  CNIVX3 U1557 ( .A(out1_0[14]), .Z(n1356) );
  CNIVX1 U1558 ( .A(n1356), .Z(n1355) );
  CNIVX3 U1559 ( .A(out1_0[43]), .Z(n1358) );
  CNIVX1 U1560 ( .A(n1358), .Z(n1357) );
  CNIVX3 U1561 ( .A(out1_0[15]), .Z(n1360) );
  CNIVX1 U1562 ( .A(n1360), .Z(n1359) );
  CMX2X1 U1563 ( .A0(n1361), .A1(n2264), .S(n7846), .Z(n7932) );
  CNIVX1 U1564 ( .A(out1_2[2]), .Z(n1361) );
  CNIVX1 U1565 ( .A(n863), .Z(n1362) );
  COND11X1 U1566 ( .A(n7734), .B(n7733), .C(n7732), .D(n7731), .Z(n863) );
  CNIVX1 U1567 ( .A(n1164), .Z(n1363) );
  CNIVX1 U1568 ( .A(n1163), .Z(n1364) );
  CNIVX1 U1569 ( .A(n7850), .Z(n1365) );
  CNIVX1 U1570 ( .A(n4385), .Z(n1366) );
  CNIVX1 U1571 ( .A(n4386), .Z(n1367) );
  CNIVX1 U1572 ( .A(n4387), .Z(n1368) );
  CNIVX1 U1573 ( .A(n7679), .Z(n1369) );
  CNIVX1 U1574 ( .A(n1021), .Z(n1370) );
  CNIVX1 U1575 ( .A(n4369), .Z(n1371) );
  CAOR2X2 U1576 ( .A(out2_2[61]), .B(n7751), .C(n7696), .D(n7738), .Z(n881) );
  CNIVX1 U1577 ( .A(n4370), .Z(n1372) );
  CNIVX1 U1578 ( .A(n4371), .Z(n1373) );
  CNIVX1 U1579 ( .A(n4374), .Z(n1374) );
  COND3X2 U1580 ( .A(n2685), .B(n2638), .C(n3278), .D(n3277), .Z(n1032) );
  CNIVX1 U1581 ( .A(n4388), .Z(n1375) );
  COND3X2 U1582 ( .A(n2685), .B(n2650), .C(n4352), .D(n4351), .Z(n1044) );
  CNIVX1 U1583 ( .A(n4381), .Z(n1376) );
  CNIVX1 U1584 ( .A(n4372), .Z(n1377) );
  CNIVX3 U1585 ( .A(out1_0[7]), .Z(n1379) );
  CNIVX1 U1586 ( .A(n1379), .Z(n1378) );
  CNIVX3 U1587 ( .A(out1_0[60]), .Z(n1381) );
  CNIVX1 U1588 ( .A(n1381), .Z(n1380) );
  COND3X2 U1589 ( .A(n2685), .B(n2643), .C(n4297), .D(n4296), .Z(n1031) );
  CNIVX1 U1590 ( .A(n1051), .Z(n1382) );
  COND3X2 U1591 ( .A(n2685), .B(n2631), .C(n3236), .D(n3235), .Z(n1035) );
  CNIVX1 U1592 ( .A(n876), .Z(n1383) );
  COND3X2 U1593 ( .A(n2685), .B(n2649), .C(n4347), .D(n4346), .Z(n1030) );
  COND3X2 U1594 ( .A(n2685), .B(n2639), .C(n3289), .D(n3288), .Z(n1042) );
  COND3X2 U1595 ( .A(n2685), .B(n2635), .C(n3257), .D(n3256), .Z(n1045) );
  COND3X2 U1596 ( .A(n2685), .B(n2636), .C(n3261), .D(n3260), .Z(n1050) );
  COND3X2 U1597 ( .A(n2685), .B(n2637), .C(n3265), .D(n3264), .Z(n1052) );
  COND3X2 U1598 ( .A(n7940), .B(n2685), .C(n2106), .D(n2107), .Z(n1054) );
  COND3X2 U1599 ( .A(n2685), .B(n2644), .C(n4302), .D(n4301), .Z(n1029) );
  CNIVX1 U1600 ( .A(n1385), .Z(n1384) );
  CNIVX1 U1601 ( .A(n1037), .Z(n1385) );
  CNIVX1 U1602 ( .A(n1125), .Z(n1386) );
  COND3X2 U1603 ( .A(n2685), .B(n2683), .C(n1996), .D(n1999), .Z(n1025) );
  CNIVX1 U1604 ( .A(n4368), .Z(n1387) );
  CNIVX1 U1605 ( .A(n4373), .Z(n1388) );
  CMXI2X1 U1606 ( .A0(n7751), .A1(n7936), .S(n7935), .Z(n1186) );
  CNIVX1 U1607 ( .A(n1155), .Z(n1389) );
  CNIVX1 U1608 ( .A(n3033), .Z(n1390) );
  CNIVX1 U1609 ( .A(n1136), .Z(n1391) );
  CMXI2X2 U1610 ( .A0(n1392), .A1(q[4]), .S(n7682), .Z(n7857) );
  CNIVX1 U1611 ( .A(q0[4]), .Z(n1392) );
  CNIVX1 U1612 ( .A(n3059), .Z(n1393) );
  CNIVX1 U1613 ( .A(n1128), .Z(n1394) );
  CNIVX1 U1614 ( .A(n1148), .Z(n1395) );
  CNIVX1 U1615 ( .A(n1127), .Z(n1396) );
  CNIVX1 U1616 ( .A(n1192), .Z(n1397) );
  CMX2X2 U1617 ( .A0(n1398), .A1(z[4]), .S(n7681), .Z(n1193) );
  CNIVX1 U1618 ( .A(acc[4]), .Z(n1398) );
  CNIVX1 U1619 ( .A(n1194), .Z(n1399) );
  CNIVX1 U1620 ( .A(n1195), .Z(n1400) );
  CNIVX1 U1621 ( .A(n1196), .Z(n1401) );
  CNIVX1 U1622 ( .A(n1202), .Z(n1402) );
  CNIVX1 U1623 ( .A(n1203), .Z(n1403) );
  CNIVX1 U1624 ( .A(n1204), .Z(n1404) );
  CNIVX1 U1625 ( .A(n1207), .Z(n1405) );
  CNIVX1 U1626 ( .A(n1208), .Z(n1406) );
  CNIVX1 U1627 ( .A(n1209), .Z(n1407) );
  CNIVX1 U1628 ( .A(n1210), .Z(n1408) );
  CNIVX1 U1629 ( .A(n1211), .Z(n1409) );
  CNIVX1 U1630 ( .A(n1212), .Z(n1410) );
  CNIVX1 U1631 ( .A(n1214), .Z(n1411) );
  CNIVX1 U1632 ( .A(n1215), .Z(n1412) );
  CNIVX1 U1633 ( .A(n1216), .Z(n1413) );
  CNIVX1 U1634 ( .A(n1217), .Z(n1414) );
  CNIVX1 U1635 ( .A(n1218), .Z(n1415) );
  CNIVX1 U1636 ( .A(n1219), .Z(n1416) );
  CNIVX1 U1637 ( .A(n1220), .Z(n1417) );
  CNIVX1 U1638 ( .A(n919), .Z(n1418) );
  CMX2X4 U1639 ( .A0(acc[0]), .A1(z[0]), .S(n7681), .Z(n1189) );
  CMX2X4 U1640 ( .A0(acc[1]), .A1(z[1]), .S(n7681), .Z(n1190) );
  CNIVX1 U1641 ( .A(n1191), .Z(n1419) );
  CMX2X4 U1642 ( .A0(acc[2]), .A1(z[2]), .S(n7681), .Z(n1191) );
  CNIVX1 U1643 ( .A(acc[9]), .Z(n1420) );
  CMX2X4 U1644 ( .A0(n1420), .A1(z[9]), .S(n7681), .Z(n1198) );
  CNIVX1 U1645 ( .A(acc[11]), .Z(n1421) );
  CMX2X4 U1646 ( .A0(n1421), .A1(z[11]), .S(n7681), .Z(n1200) );
  CNIVX1 U1647 ( .A(acc[12]), .Z(n1422) );
  CMX2XL U1648 ( .A0(acc[16]), .A1(z[16]), .S(n7681), .Z(n1205) );
  CNIVX1 U1649 ( .A(n1205), .Z(n1423) );
  CNIVX1 U1650 ( .A(n1206), .Z(n1424) );
  CMX2X4 U1651 ( .A0(acc[17]), .A1(z[17]), .S(n7681), .Z(n1206) );
  CNIVX1 U1652 ( .A(acc[24]), .Z(n1425) );
  CNIVX1 U1653 ( .A(n914), .Z(n1426) );
  CNIVX1 U1654 ( .A(n1053), .Z(n1427) );
  COND3X2 U1655 ( .A(n2685), .B(n2641), .C(n4285), .D(n4284), .Z(n1049) );
  CNIVX1 U1656 ( .A(n925), .Z(n1428) );
  CNIVX1 U1657 ( .A(acc[8]), .Z(n1429) );
  COND3X2 U1658 ( .A(n2653), .B(n2685), .C(n1880), .D(n1883), .Z(n1009) );
  CNIVX1 U1659 ( .A(acc[10]), .Z(n1430) );
  CNIVX1 U1660 ( .A(n3071), .Z(n1431) );
  CNIVX3 U1661 ( .A(n2628), .Z(n1432) );
  CNIVX1 U1662 ( .A(n3076), .Z(n1433) );
  CNIVX1 U1663 ( .A(n3089), .Z(n1434) );
  CNIVX1 U1664 ( .A(n1133), .Z(n1435) );
  CNIVX3 U1665 ( .A(out1_0[11]), .Z(n1437) );
  CNIVX1 U1666 ( .A(n1437), .Z(n1436) );
  CNIVX1 U1667 ( .A(n1146), .Z(n1438) );
  CNIVX1 U1668 ( .A(n3090), .Z(n1439) );
  CNIVX1 U1669 ( .A(n1167), .Z(n1440) );
  CNIVX1 U1670 ( .A(n1147), .Z(n1441) );
  CNIVX1 U1671 ( .A(n1443), .Z(n1442) );
  CNIVX1 U1672 ( .A(cmd0[1]), .Z(n1443) );
  CNIVX3 U1673 ( .A(out1_0[10]), .Z(n1445) );
  CNIVX1 U1674 ( .A(n1445), .Z(n1444) );
  CIVXL U1675 ( .A(out2_2[21]), .Z(n4279) );
  CNIVX1 U1676 ( .A(n1135), .Z(n1446) );
  CNIVX1 U1677 ( .A(n1134), .Z(n1447) );
  CNIVX1 U1678 ( .A(n3117), .Z(n1448) );
  CNIVX1 U1679 ( .A(n1138), .Z(n1449) );
  CIVXL U1680 ( .A(out2_2[9]), .Z(n3333) );
  CNIVX1 U1681 ( .A(n1154), .Z(n1450) );
  CNIVX3 U1682 ( .A(out1_0[32]), .Z(n1452) );
  CNIVX1 U1683 ( .A(n1452), .Z(n1451) );
  CNIVX3 U1684 ( .A(out1_0[17]), .Z(n1454) );
  CNIVX1 U1685 ( .A(n1454), .Z(n1453) );
  CNIVX3 U1686 ( .A(out1_0[6]), .Z(n1456) );
  CNIVX1 U1687 ( .A(n1456), .Z(n1455) );
  CNIVX3 U1688 ( .A(out1_0[9]), .Z(n1458) );
  CNIVX1 U1689 ( .A(n1458), .Z(n1457) );
  CNIVX3 U1690 ( .A(out1_0[8]), .Z(n1460) );
  CNIVX1 U1691 ( .A(n1460), .Z(n1459) );
  CNIVX3 U1692 ( .A(out1_0[20]), .Z(n1462) );
  CNIVX1 U1693 ( .A(n1462), .Z(n1461) );
  CNIVX3 U1694 ( .A(out1_0[5]), .Z(n1464) );
  CNIVX1 U1695 ( .A(n1464), .Z(n1463) );
  CNIVX3 U1696 ( .A(out1_0[12]), .Z(n1466) );
  CNIVX1 U1697 ( .A(n1466), .Z(n1465) );
  CNIVX3 U1698 ( .A(out1_0[26]), .Z(n1468) );
  CNIVX1 U1699 ( .A(n1468), .Z(n1467) );
  CNIVX3 U1700 ( .A(out1_0[16]), .Z(n1470) );
  CNIVX1 U1701 ( .A(n1470), .Z(n1469) );
  CNIVX3 U1702 ( .A(out1_0[25]), .Z(n1472) );
  CNIVX1 U1703 ( .A(n1472), .Z(n1471) );
  CNIVXL U1704 ( .A(n2682), .Z(n1473) );
  CNIVX3 U1705 ( .A(out1_0[3]), .Z(n1475) );
  CNIVX1 U1706 ( .A(n1475), .Z(n1474) );
  CNIVX3 U1707 ( .A(out1_0[4]), .Z(n1477) );
  CNIVX1 U1708 ( .A(n1477), .Z(n1476) );
  CNIVX3 U1709 ( .A(out1_0[2]), .Z(n1479) );
  CNIVX1 U1710 ( .A(n1479), .Z(n1478) );
  CNIVX3 U1711 ( .A(out1_0[49]), .Z(n1481) );
  CNIVX1 U1712 ( .A(n1481), .Z(n1480) );
  CNIVX3 U1713 ( .A(push0_1), .Z(n1483) );
  CNIVX1 U1714 ( .A(n1483), .Z(n1482) );
  CNIVX3 U1715 ( .A(out1_0[0]), .Z(n1485) );
  CNIVX1 U1716 ( .A(n1485), .Z(n1484) );
  CNIVX3 U1717 ( .A(out1_0[41]), .Z(n1487) );
  CNIVX1 U1718 ( .A(n1487), .Z(n1486) );
  CNIVX1 U1719 ( .A(n1489), .Z(n1488) );
  CNIVX1 U1720 ( .A(push0), .Z(n1489) );
  CNIVX3 U1721 ( .A(cmd0_1[1]), .Z(n1491) );
  CNIVX1 U1722 ( .A(n1491), .Z(n1490) );
  CNIVX3 U1723 ( .A(push0_0), .Z(n1493) );
  CNIVX1 U1724 ( .A(n1493), .Z(n1492) );
  CNIVX3 U1725 ( .A(out1_0[63]), .Z(n1495) );
  CNIVX1 U1726 ( .A(n1495), .Z(n1494) );
  CNIVX3 U1727 ( .A(out1_0[22]), .Z(n1497) );
  CNIVX1 U1728 ( .A(n1497), .Z(n1496) );
  CNIVX3 U1729 ( .A(out1_0[54]), .Z(n1499) );
  CNIVX1 U1730 ( .A(n1499), .Z(n1498) );
  CNIVX3 U1731 ( .A(out1_0[58]), .Z(n1501) );
  CNIVX1 U1732 ( .A(n1501), .Z(n1500) );
  CNIVX3 U1733 ( .A(out1_0[47]), .Z(n1503) );
  CNIVX1 U1734 ( .A(n1503), .Z(n1502) );
  CNIVX3 U1735 ( .A(out1_0[57]), .Z(n1505) );
  CNIVX1 U1736 ( .A(n1505), .Z(n1504) );
  CMXI2X2 U1737 ( .A0(n4367), .A1(q[24]), .S(n7682), .Z(n2680) );
  CNIVX3 U1738 ( .A(out1_0[52]), .Z(n1507) );
  CNIVX1 U1739 ( .A(n1507), .Z(n1506) );
  CNIVX3 U1740 ( .A(out1_0[45]), .Z(n1509) );
  CNIVX1 U1741 ( .A(n1509), .Z(n1508) );
  CNIVX3 U1742 ( .A(out1_0[44]), .Z(n1511) );
  CNIVX1 U1743 ( .A(n1511), .Z(n1510) );
  CNIVX3 U1744 ( .A(out1_0[50]), .Z(n1513) );
  CNIVX1 U1745 ( .A(n1513), .Z(n1512) );
  CNIVX3 U1746 ( .A(out1_0[55]), .Z(n1515) );
  CNIVX1 U1747 ( .A(n1515), .Z(n1514) );
  CNIVX3 U1748 ( .A(out1_0[48]), .Z(n1517) );
  CNIVX1 U1749 ( .A(n1517), .Z(n1516) );
  CNIVX3 U1750 ( .A(out1_0[51]), .Z(n1519) );
  CNIVX1 U1751 ( .A(n1519), .Z(n1518) );
  CNIVX3 U1752 ( .A(out1_0[59]), .Z(n1521) );
  CNIVX1 U1753 ( .A(n1521), .Z(n1520) );
  CNIVX3 U1754 ( .A(out1_0[53]), .Z(n1523) );
  CNIVX1 U1755 ( .A(n1523), .Z(n1522) );
  CNIVX3 U1756 ( .A(out1_0[56]), .Z(n1525) );
  CNIVX1 U1757 ( .A(n1525), .Z(n1524) );
  CNIVX3 U1758 ( .A(out1_0[27]), .Z(n1527) );
  CNIVX1 U1759 ( .A(n1527), .Z(n1526) );
  CNIVX3 U1760 ( .A(out1_0[23]), .Z(n1529) );
  CNIVX1 U1761 ( .A(n1529), .Z(n1528) );
  CNIVX1 U1762 ( .A(n1166), .Z(n1530) );
  CNIVX3 U1763 ( .A(out1_0[21]), .Z(n1532) );
  CNIVX1 U1764 ( .A(n1532), .Z(n1531) );
  CNIVX3 U1765 ( .A(out1_0[30]), .Z(n1534) );
  CNIVX1 U1766 ( .A(n1534), .Z(n1533) );
  CNIVX4 U1767 ( .A(n6576), .Z(n6527) );
  CND2X1 U1768 ( .A(n5092), .B(n5091), .Z(n1537) );
  CND2X1 U1769 ( .A(n1535), .B(n1536), .Z(n1538) );
  CND2X2 U1770 ( .A(n1537), .B(n1538), .Z(n5093) );
  CIVXL U1771 ( .A(n5092), .Z(n1535) );
  CIVX2 U1772 ( .A(n5091), .Z(n1536) );
  CENX2 U1773 ( .A(n1594), .B(n3487), .Z(n1599) );
  CND2XL U1774 ( .A(n2308), .B(n6267), .Z(n1539) );
  CENX1 U1775 ( .A(n1540), .B(n5432), .Z(n5442) );
  CENX1 U1776 ( .A(n5433), .B(n5434), .Z(n1540) );
  CND2X1 U1777 ( .A(n5289), .B(n5290), .Z(n1543) );
  CND2X2 U1778 ( .A(n1541), .B(n1542), .Z(n1544) );
  CND2X2 U1779 ( .A(n1543), .B(n1544), .Z(n5518) );
  CIVXL U1780 ( .A(n5290), .Z(n1541) );
  CIVX2 U1781 ( .A(n5289), .Z(n1542) );
  COR2XL U1782 ( .A(n5984), .B(n6210), .Z(n6099) );
  COND1XL U1783 ( .A(n6827), .B(n6969), .C(n6826), .Z(n6890) );
  CND2X4 U1784 ( .A(n4717), .B(n4716), .Z(n4897) );
  CNIVX4 U1785 ( .A(n3796), .Z(n1545) );
  CND2X2 U1786 ( .A(n5436), .B(n5435), .Z(n5465) );
  COAN1X2 U1787 ( .A(n7858), .B(n3353), .C(n3351), .Z(n1588) );
  CIVXL U1788 ( .A(n7039), .Z(n7030) );
  CNIVX1 U1789 ( .A(n6197), .Z(n2439) );
  CAN2XL U1790 ( .A(n2308), .B(n6267), .Z(n1546) );
  CENX1 U1791 ( .A(q0[24]), .B(q0[23]), .Z(n1547) );
  CIVX2 U1792 ( .A(n4659), .Z(n1548) );
  CIVX3 U1793 ( .A(n7171), .Z(n1549) );
  CIVX2 U1794 ( .A(n4658), .Z(n4659) );
  CIVXL U1795 ( .A(n4683), .Z(n4658) );
  CIVX4 U1796 ( .A(n4683), .Z(n4684) );
  CND2X2 U1797 ( .A(n6281), .B(n6280), .Z(n7047) );
  CIVXL U1798 ( .A(n1546), .Z(n1550) );
  CENX1 U1799 ( .A(n5090), .B(n5089), .Z(n5248) );
  CENXL U1800 ( .A(n5088), .B(n5087), .Z(n5089) );
  CNIVX1 U1801 ( .A(n2658), .Z(n1551) );
  CND2X1 U1802 ( .A(q0[15]), .B(q0[16]), .Z(n1554) );
  CND2X2 U1803 ( .A(n1552), .B(n1553), .Z(n1555) );
  CND2X4 U1804 ( .A(n1554), .B(n1555), .Z(n4670) );
  CIVX2 U1805 ( .A(q0[15]), .Z(n1552) );
  CIVX2 U1806 ( .A(q0[16]), .Z(n1553) );
  CNIVX16 U1807 ( .A(n4670), .Z(n6765) );
  CND2IX2 U1808 ( .B(n4763), .A(n4662), .Z(n4667) );
  CENX2 U1809 ( .A(n5932), .B(n6185), .Z(n4763) );
  COND1X1 U1810 ( .A(n4703), .B(n4705), .C(n4702), .Z(n4674) );
  CNIVX4 U1811 ( .A(n3459), .Z(n1556) );
  CNIVX4 U1812 ( .A(n3459), .Z(n1557) );
  CNIVX1 U1813 ( .A(n3459), .Z(n6525) );
  CEO3X1 U1814 ( .A(n6720), .B(n6721), .C(n6722), .Z(n6743) );
  CND2XL U1815 ( .A(n6720), .B(n6722), .Z(n1558) );
  CND2X1 U1816 ( .A(n6720), .B(n6721), .Z(n1559) );
  CND2X1 U1817 ( .A(n6722), .B(n6721), .Z(n1560) );
  CND3X2 U1818 ( .A(n1558), .B(n1559), .C(n1560), .Z(n6777) );
  CANR1XL U1819 ( .A(n6961), .B(n7415), .C(n6960), .Z(n1561) );
  CANR1XL U1820 ( .A(n6961), .B(n7415), .C(n6960), .Z(n1562) );
  COND1X1 U1821 ( .A(n6778), .B(n6777), .C(n6776), .Z(n6780) );
  CENX2 U1822 ( .A(n6723), .B(n6777), .Z(n6811) );
  CANR1X1 U1823 ( .A(n6961), .B(n7415), .C(n6960), .Z(n6962) );
  CNR2X4 U1824 ( .A(n1587), .B(n5468), .Z(n5503) );
  CND2X1 U1825 ( .A(n2464), .B(n2658), .Z(n2590) );
  COND1XL U1826 ( .A(n7051), .B(n6963), .C(n1561), .Z(n1563) );
  CND2X1 U1827 ( .A(n6952), .B(n6951), .Z(n7340) );
  CEN3X2 U1828 ( .A(n5327), .B(n5326), .C(n5325), .Z(n2347) );
  CND2X1 U1829 ( .A(n6083), .B(n6067), .Z(n6068) );
  CND2X1 U1830 ( .A(n5480), .B(n5479), .Z(n1566) );
  CND2X2 U1831 ( .A(n1564), .B(n1565), .Z(n1567) );
  CND2X2 U1832 ( .A(n1566), .B(n1567), .Z(n5481) );
  CIVX2 U1833 ( .A(n5480), .Z(n1564) );
  CIVX2 U1834 ( .A(n5479), .Z(n1565) );
  CEO3X2 U1835 ( .A(n5341), .B(n5339), .C(n5340), .Z(n5424) );
  CND2XL U1836 ( .A(n1266), .B(n5339), .Z(n1569) );
  CND2X1 U1837 ( .A(n5340), .B(n5339), .Z(n1570) );
  CND3X1 U1838 ( .A(n1568), .B(n1569), .C(n1570), .Z(n5320) );
  CIVXL U1839 ( .A(n2442), .Z(n2443) );
  CENX2 U1840 ( .A(n5413), .B(n5412), .Z(n5454) );
  CENXL U1841 ( .A(n2454), .B(h0[25]), .Z(n6492) );
  CND2X2 U1842 ( .A(n2604), .B(n2605), .Z(n1571) );
  CND2X1 U1843 ( .A(n2604), .B(n2605), .Z(n5603) );
  CND2X1 U1844 ( .A(n5651), .B(n5673), .Z(n1574) );
  CND2X2 U1845 ( .A(n1572), .B(n1573), .Z(n1575) );
  CND2X2 U1846 ( .A(n1574), .B(n1575), .Z(n5775) );
  CIVX2 U1847 ( .A(n5651), .Z(n1572) );
  CIVXL U1848 ( .A(n5673), .Z(n1573) );
  CIVX3 U1849 ( .A(n5775), .Z(n5661) );
  COND1XL U1850 ( .A(n7527), .B(n7525), .C(n7528), .Z(n1576) );
  CNIVXL U1851 ( .A(n5666), .Z(n1577) );
  CND2X1 U1852 ( .A(n5631), .B(n5752), .Z(n1580) );
  CND2X2 U1853 ( .A(n1578), .B(n1579), .Z(n1581) );
  CND2X2 U1854 ( .A(n1580), .B(n1581), .Z(n5671) );
  CIVX2 U1855 ( .A(n5631), .Z(n1578) );
  CIVX2 U1856 ( .A(n5752), .Z(n1579) );
  COND2X4 U1857 ( .A(n7171), .B(n6669), .C(n6774), .D(n6641), .Z(n6678) );
  CNIVX4 U1858 ( .A(n3382), .Z(n1582) );
  CNIVX2 U1859 ( .A(n3382), .Z(n6766) );
  CENX1 U1860 ( .A(n6179), .B(n6180), .Z(n6147) );
  CENX1 U1861 ( .A(n6181), .B(n6147), .Z(n6224) );
  COND1X1 U1862 ( .A(n6224), .B(n6225), .C(n6223), .Z(n6227) );
  CMX2XL U1863 ( .A0(h0[17]), .A1(h[17]), .S(n7682), .Z(n946) );
  CIVXL U1864 ( .A(n4397), .Z(n1583) );
  CEO3X2 U1865 ( .A(n5623), .B(n4993), .C(n5621), .Z(n1584) );
  CIVXL U1866 ( .A(n6525), .Z(n1585) );
  CIVX2 U1867 ( .A(n1585), .Z(n1586) );
  CNR2X2 U1868 ( .A(n5511), .B(n5467), .Z(n1587) );
  CIVX4 U1869 ( .A(n2582), .Z(n2583) );
  CND2XL U1870 ( .A(n6088), .B(n6090), .Z(n6091) );
  CENX2 U1871 ( .A(n6217), .B(n6219), .Z(n6171) );
  CND2X1 U1872 ( .A(n5237), .B(n5235), .Z(n4938) );
  CND2X1 U1873 ( .A(n4498), .B(n4497), .Z(n4541) );
  COND1XL U1874 ( .A(n4508), .B(n4505), .C(n4506), .Z(n4498) );
  CND2X1 U1875 ( .A(n6624), .B(n6623), .Z(n6625) );
  CENX1 U1876 ( .A(n6672), .B(n6671), .Z(n6621) );
  CND2XL U1877 ( .A(n6902), .B(n6903), .Z(n6609) );
  CENX1 U1878 ( .A(n7173), .B(h0[3]), .Z(n5755) );
  CND2X2 U1879 ( .A(n2379), .B(n2380), .Z(n6358) );
  COR2XL U1880 ( .A(n7114), .B(n6301), .Z(n2380) );
  COND2X1 U1881 ( .A(n6701), .B(n6146), .C(n6765), .D(n6188), .Z(n6180) );
  COND1X1 U1882 ( .A(n6142), .B(n6141), .C(n6140), .Z(n6143) );
  CNIVX1 U1883 ( .A(n5277), .Z(n5131) );
  CNIVX2 U1884 ( .A(n5237), .Z(n5238) );
  CFA1X1 U1885 ( .A(n4874), .B(n4873), .CI(n4872), .CO(n4815), .S(n5085) );
  CENX1 U1886 ( .A(n5613), .B(n5612), .Z(n5071) );
  CND3X1 U1887 ( .A(n2474), .B(n2475), .C(n2476), .Z(n5559) );
  CENX1 U1888 ( .A(h0[27]), .B(n6970), .Z(n6866) );
  CND2X1 U1889 ( .A(n6986), .B(n6985), .Z(n7072) );
  CND2XL U1890 ( .A(n6984), .B(n6983), .Z(n6985) );
  CND2X1 U1891 ( .A(n3648), .B(n3650), .Z(n3635) );
  CND2X1 U1892 ( .A(n3751), .B(n3750), .Z(n3752) );
  COND1X1 U1893 ( .A(n3751), .B(n3750), .C(n3749), .Z(n3753) );
  CENX1 U1894 ( .A(n4567), .B(n4566), .Z(n4568) );
  CIVX2 U1895 ( .A(n2299), .Z(n2300) );
  CND2X1 U1896 ( .A(n6690), .B(n6689), .Z(n6691) );
  CND2X1 U1897 ( .A(n6549), .B(n6548), .Z(n6658) );
  COND1X1 U1898 ( .A(n3588), .B(n3591), .C(n3589), .Z(n3571) );
  CENX1 U1899 ( .A(n3427), .B(n2031), .Z(n3438) );
  CND2X1 U1900 ( .A(n4552), .B(n4550), .Z(n4468) );
  COND1X1 U1901 ( .A(n4550), .B(n4552), .C(n4549), .Z(n4469) );
  CIVX2 U1902 ( .A(n5259), .Z(n5222) );
  CND2X1 U1903 ( .A(n6447), .B(n6446), .Z(n6448) );
  CND2X1 U1904 ( .A(n6899), .B(n6901), .Z(n6611) );
  COND1X1 U1905 ( .A(n5946), .B(n5945), .C(n5944), .Z(n5949) );
  CND2X1 U1906 ( .A(n5938), .B(n5937), .Z(n5939) );
  CNIVX1 U1907 ( .A(n5424), .Z(n5345) );
  COND2X1 U1908 ( .A(n7228), .B(n5755), .C(n5818), .D(n2381), .Z(n5857) );
  CND2XL U1909 ( .A(n6501), .B(n6500), .Z(n6502) );
  COND1X1 U1910 ( .A(n6504), .B(n6505), .C(n6528), .Z(n6507) );
  CND2X1 U1911 ( .A(n6505), .B(n6504), .Z(n6506) );
  CND2X1 U1912 ( .A(n7009), .B(n7010), .Z(n7011) );
  CENX1 U1913 ( .A(n5801), .B(n5800), .Z(n5803) );
  COND2X1 U1914 ( .A(n2449), .B(n3391), .C(n1557), .D(n3402), .Z(n3359) );
  CND2XL U1915 ( .A(n3762), .B(n3761), .Z(n3763) );
  CENX1 U1916 ( .A(n5106), .B(h0[20]), .Z(n4495) );
  COND2X1 U1917 ( .A(n6703), .B(n5995), .C(n2514), .D(n5994), .Z(n6017) );
  COND1X1 U1918 ( .A(n6239), .B(n6238), .C(n6237), .Z(n6242) );
  COND1X1 U1919 ( .A(n6126), .B(n6127), .C(n6125), .Z(n6129) );
  CND2X1 U1920 ( .A(n6127), .B(n6126), .Z(n6128) );
  CNIVX1 U1921 ( .A(n5622), .Z(n4993) );
  COND2X1 U1922 ( .A(n6972), .B(n6868), .C(n6824), .D(n6974), .Z(n6889) );
  COND2X1 U1923 ( .A(n6640), .B(n7065), .C(n2477), .D(n6676), .Z(n6680) );
  COND2X1 U1924 ( .A(n7205), .B(n6642), .C(n7203), .D(n6708), .Z(n6679) );
  COND1XL U1925 ( .A(n6879), .B(n6878), .C(n6877), .Z(n6881) );
  CNIVX2 U1926 ( .A(n4861), .Z(n3674) );
  CENX1 U1927 ( .A(n5701), .B(h0[7]), .Z(n3512) );
  COND2X1 U1928 ( .A(n6522), .B(n3500), .C(n6293), .D(n3450), .Z(n3494) );
  CENX1 U1929 ( .A(h0[11]), .B(n5566), .Z(n3490) );
  CENX1 U1930 ( .A(n3766), .B(n3767), .Z(n3358) );
  CENX1 U1931 ( .A(n4472), .B(n4404), .Z(n4466) );
  CNIVX1 U1932 ( .A(n5327), .Z(n5198) );
  CNIVX1 U1933 ( .A(n5293), .Z(n5206) );
  CND2X1 U1934 ( .A(n5084), .B(n5086), .Z(n4875) );
  COND1X1 U1935 ( .A(n5086), .B(n5084), .C(n5085), .Z(n4876) );
  CND2X1 U1936 ( .A(n4898), .B(n4897), .Z(n4899) );
  COND1X1 U1937 ( .A(n6012), .B(n6013), .C(n6011), .Z(n6015) );
  CND2X1 U1938 ( .A(n6034), .B(n6033), .Z(n6035) );
  CND2X1 U1939 ( .A(n6354), .B(n6353), .Z(n6355) );
  COND1X1 U1940 ( .A(n6342), .B(n6343), .C(n6341), .Z(n6345) );
  CND2X1 U1941 ( .A(n6343), .B(n6342), .Z(n6344) );
  CND2X1 U1942 ( .A(n6350), .B(n6349), .Z(n6432) );
  CND2XL U1943 ( .A(n6244), .B(n6246), .Z(n6247) );
  COND1X1 U1944 ( .A(n6246), .B(n6244), .C(n6245), .Z(n6248) );
  COND1X1 U1945 ( .A(n6180), .B(n6181), .C(n6179), .Z(n6183) );
  CND3X1 U1946 ( .A(n6054), .B(n6056), .C(n6055), .Z(n6061) );
  CND2X2 U1947 ( .A(n5594), .B(n5593), .Z(n5736) );
  CND2IX1 U1948 ( .B(n5590), .A(n5589), .Z(n5594) );
  CND3X1 U1949 ( .A(n2517), .B(n2518), .C(n2519), .Z(n5737) );
  CND2X1 U1950 ( .A(n5586), .B(n5585), .Z(n5587) );
  COND1X1 U1951 ( .A(n5585), .B(n5586), .C(n5584), .Z(n5588) );
  CIVX2 U1952 ( .A(n5106), .Z(n2510) );
  CENX1 U1953 ( .A(n5932), .B(h0[8]), .Z(n4688) );
  CENX1 U1954 ( .A(n6699), .B(h0[23]), .Z(n6300) );
  CEOX1 U1955 ( .A(h0[13]), .B(n7851), .Z(n6309) );
  CND2XL U1956 ( .A(n6598), .B(n6597), .Z(n6599) );
  COND1X1 U1957 ( .A(n6427), .B(n6428), .C(n6426), .Z(n6430) );
  CND2X1 U1958 ( .A(n6394), .B(n6393), .Z(n6395) );
  COND1X1 U1959 ( .A(n6393), .B(n6394), .C(n6392), .Z(n6396) );
  CNIVX1 U1960 ( .A(n7217), .Z(n7123) );
  COND1X1 U1961 ( .A(n4559), .B(n4560), .C(n4558), .Z(n4562) );
  COND1X1 U1962 ( .A(n4594), .B(n4595), .C(n4593), .Z(n4597) );
  CND2X1 U1963 ( .A(n4595), .B(n4594), .Z(n4596) );
  CND3X1 U1964 ( .A(n2354), .B(n2355), .C(n2356), .Z(n5448) );
  CND2X1 U1965 ( .A(n4585), .B(n4583), .Z(n4462) );
  CND2X1 U1966 ( .A(n5131), .B(n5280), .Z(n5132) );
  COND1X1 U1967 ( .A(n5280), .B(n5131), .C(n5278), .Z(n5133) );
  CNIVX2 U1968 ( .A(n5012), .Z(n4908) );
  CNIVX1 U1969 ( .A(n6085), .Z(n6067) );
  CNIVX1 U1970 ( .A(n6136), .Z(n6137) );
  CND2X1 U1971 ( .A(n7391), .B(n7395), .Z(n6959) );
  CND2XL U1972 ( .A(n5788), .B(n5787), .Z(n5789) );
  COND1X1 U1973 ( .A(n5560), .B(n5561), .C(n5559), .Z(n5563) );
  COND1X1 U1974 ( .A(n7145), .B(n7146), .C(n7144), .Z(n7148) );
  CND2XL U1975 ( .A(n7146), .B(n7145), .Z(n7147) );
  CND2X1 U1976 ( .A(n6792), .B(n6791), .Z(n6832) );
  COND2X1 U1977 ( .A(n7217), .B(n6823), .C(n7203), .D(n6891), .Z(n6862) );
  COND1X1 U1978 ( .A(n6725), .B(n6726), .C(n6724), .Z(n6728) );
  CND2XL U1979 ( .A(n6726), .B(n6725), .Z(n6727) );
  CIVX4 U1980 ( .A(n4783), .Z(n4732) );
  CNIVX2 U1981 ( .A(n4786), .Z(n4792) );
  CENX1 U1982 ( .A(n7173), .B(h0[1]), .Z(n5039) );
  CENX1 U1983 ( .A(n7173), .B(h0[2]), .Z(n5700) );
  CENX1 U1984 ( .A(n2660), .B(h0[19]), .Z(n5709) );
  CNIVX1 U1985 ( .A(n7051), .Z(n7052) );
  CND2X1 U1986 ( .A(n7260), .B(n7264), .Z(n7164) );
  CNIVX1 U1987 ( .A(n6992), .Z(n6993) );
  CNIVX1 U1988 ( .A(n6658), .Z(n6659) );
  COND2X1 U1989 ( .A(n7119), .B(n7118), .C(n7171), .D(n7135), .Z(n7144) );
  COND1X1 U1990 ( .A(n7097), .B(n7098), .C(n7096), .Z(n7100) );
  CFA1X1 U1991 ( .A(n7069), .B(n7068), .CI(n7067), .CO(n7098), .S(n7076) );
  CENX1 U1992 ( .A(n7097), .B(n7096), .Z(n7070) );
  CND2XL U1993 ( .A(n7072), .B(n7071), .Z(n2325) );
  CND2XL U1994 ( .A(n7073), .B(n7072), .Z(n2323) );
  COND1X1 U1995 ( .A(n3650), .B(n3648), .C(n3649), .Z(n1861) );
  CND2XL U1996 ( .A(n3440), .B(n3437), .Z(n3428) );
  COND1X1 U1997 ( .A(n3440), .B(n3437), .C(n3438), .Z(n3429) );
  CND2X1 U1998 ( .A(n3523), .B(n3524), .Z(n3466) );
  CNR2X1 U1999 ( .A(n3523), .B(n3524), .Z(n3468) );
  CND2X1 U2000 ( .A(n4619), .B(n4618), .Z(n4620) );
  COND1X1 U2001 ( .A(n4618), .B(n4619), .C(n4617), .Z(n4621) );
  CND2X1 U2002 ( .A(n4589), .B(n4587), .Z(n4570) );
  COND1X1 U2003 ( .A(n4587), .B(n4589), .C(n4586), .Z(n4571) );
  CND2XL U2004 ( .A(n5244), .B(n5243), .Z(n5240) );
  COND1X1 U2005 ( .A(n5243), .B(n5244), .C(n5245), .Z(n5241) );
  CNIVX1 U2006 ( .A(n5388), .Z(n2559) );
  CNIVX1 U2007 ( .A(n5361), .Z(n4981) );
  CND2XL U2008 ( .A(n6070), .B(n6008), .Z(n6009) );
  CND2X1 U2009 ( .A(n6332), .B(n6331), .Z(n6333) );
  CND2XL U2010 ( .A(n6784), .B(n6783), .Z(n6785) );
  CNR2X1 U2011 ( .A(n6784), .B(n6783), .Z(n6787) );
  CND2X1 U2012 ( .A(n6734), .B(n6733), .Z(n6735) );
  COND1X1 U2013 ( .A(n6733), .B(n6734), .C(n6732), .Z(n6736) );
  CENX1 U2014 ( .A(n6783), .B(n6784), .Z(n6758) );
  CENX1 U2015 ( .A(n6690), .B(n6630), .Z(n6712) );
  CND2X1 U2016 ( .A(n6685), .B(n6684), .Z(n6686) );
  COND1X1 U2017 ( .A(n6684), .B(n6685), .C(n6683), .Z(n6687) );
  CENX1 U2018 ( .A(n5106), .B(h0[28]), .Z(n4710) );
  CND2X1 U2019 ( .A(n4940), .B(n4942), .Z(n4700) );
  COND1X1 U2020 ( .A(n4940), .B(n4942), .C(n4939), .Z(n4701) );
  CNR2X1 U2021 ( .A(n6701), .B(n5704), .Z(n5705) );
  CND2X1 U2022 ( .A(n5487), .B(n5486), .Z(n5498) );
  CND2X1 U2023 ( .A(n6894), .B(n6893), .Z(n6895) );
  COND1X1 U2024 ( .A(n3625), .B(n3626), .C(n3624), .Z(n3622) );
  CND2X1 U2025 ( .A(n3626), .B(n3625), .Z(n3621) );
  CENX1 U2026 ( .A(n3599), .B(n3598), .Z(n3733) );
  CND2X1 U2027 ( .A(n3591), .B(n3588), .Z(n3570) );
  CANR1X1 U2028 ( .A(n6387), .B(n6386), .C(n3727), .Z(n3728) );
  CND2XL U2029 ( .A(n3598), .B(n3597), .Z(n3521) );
  COND1X1 U2030 ( .A(n3597), .B(n3598), .C(n3596), .Z(n3522) );
  CND2X1 U2031 ( .A(n3551), .B(n3550), .Z(n3552) );
  COND1X1 U2032 ( .A(n3551), .B(n3550), .C(n3549), .Z(n3553) );
  CND2X1 U2033 ( .A(n6089), .B(n6088), .Z(n6092) );
  CND2X1 U2034 ( .A(n8012), .B(n8013), .Z(n7553) );
  CIVX2 U2035 ( .A(n7763), .Z(n3169) );
  CIVX2 U2036 ( .A(n7770), .Z(n3172) );
  CIVX2 U2037 ( .A(n7553), .Z(n7582) );
  CNR2X1 U2038 ( .A(n7425), .B(n7236), .Z(n7315) );
  COND2X1 U2039 ( .A(n5911), .B(n4949), .C(n5912), .D(n4854), .Z(n5130) );
  CND2X1 U2040 ( .A(n5941), .B(n5940), .Z(n5942) );
  COND1X1 U2041 ( .A(n5941), .B(n5940), .C(n5918), .Z(n5943) );
  CND2X1 U2042 ( .A(n5025), .B(n5024), .Z(n5026) );
  COND1X1 U2043 ( .A(n5024), .B(n5025), .C(n5023), .Z(n5027) );
  CND2X1 U2044 ( .A(q0[3]), .B(n2532), .Z(n2534) );
  CENX1 U2045 ( .A(n6699), .B(h0[12]), .Z(n4699) );
  CENX1 U2046 ( .A(n5188), .B(n5187), .Z(n5189) );
  CND2XL U2047 ( .A(n4963), .B(n2657), .Z(n5214) );
  CND2XL U2048 ( .A(n2658), .B(n4419), .Z(n4420) );
  CND2X1 U2049 ( .A(n7724), .B(n8020), .Z(n7722) );
  CIVX2 U2050 ( .A(n7722), .Z(n7738) );
  CND3X1 U2051 ( .A(cmd0_2[1]), .B(cmd0_2[0]), .C(push0_2), .Z(n7681) );
  CDLY1XL U2052 ( .A(q0[14]), .Z(n3211) );
  CIVX2 U2053 ( .A(n7432), .Z(n7192) );
  CNIVX1 U2054 ( .A(n7374), .Z(n7384) );
  CIVX2 U2055 ( .A(n7758), .Z(n7747) );
  CIVX2 U2056 ( .A(n7744), .Z(n7755) );
  CIVX2 U2057 ( .A(n7766), .Z(n3173) );
  COR2X1 U2058 ( .A(n3724), .B(n3723), .Z(n6389) );
  CNR2X1 U2059 ( .A(n3731), .B(n3730), .Z(n7503) );
  CND2X1 U2060 ( .A(n8020), .B(n8016), .Z(n7729) );
  CNR2X1 U2061 ( .A(h0_1[5]), .B(h0_1[6]), .Z(n7724) );
  COND1XL U2062 ( .A(n5125), .B(n5127), .C(n5124), .Z(n4849) );
  CNIVX4 U2063 ( .A(h0[9]), .Z(n5927) );
  CND2X1 U2064 ( .A(n5762), .B(n5761), .Z(n5879) );
  CIVDX2 U2065 ( .A(q0[27]), .Z0(n4851), .Z1(n7062) );
  CNIVX8 U2066 ( .A(h0[0]), .Z(n7539) );
  CENX1 U2067 ( .A(n7092), .B(h0[2]), .Z(n5212) );
  CND2X1 U2068 ( .A(n5345), .B(n5426), .Z(n5346) );
  CND2X1 U2069 ( .A(n5858), .B(n5857), .Z(n5859) );
  CNR2X1 U2070 ( .A(n5867), .B(n6522), .Z(n5868) );
  CND2X1 U2071 ( .A(n6503), .B(n6502), .Z(n6602) );
  CMX2X2 U2072 ( .A0(h0_1[4]), .A1(h0_0[4]), .S(cmd2_en_1), .Z(n927) );
  CMX2X1 U2073 ( .A0(h0_1[5]), .A1(h0_0[5]), .S(cmd2_en_1), .Z(n930) );
  CMX2X2 U2074 ( .A0(h0_1[6]), .A1(h0_0[6]), .S(cmd2_en_1), .Z(n933) );
  CAN2XL U2075 ( .A(n5396), .B(n5393), .Z(n4647) );
  COND1XL U2076 ( .A(n7495), .B(n7494), .C(n7493), .Z(n7499) );
  CANR1XL U2077 ( .A(n7492), .B(n7491), .C(n7490), .Z(n7493) );
  CIVX2 U2078 ( .A(n5932), .Z(n2315) );
  COND2X1 U2079 ( .A(n5171), .B(n5695), .C(n4886), .D(n5170), .Z(n5339) );
  COND1X1 U2080 ( .A(n5952), .B(n5951), .C(n5950), .Z(n6168) );
  CENX1 U2081 ( .A(n7092), .B(n2513), .Z(n4961) );
  COND1X1 U2082 ( .A(n5203), .B(n5201), .C(n5202), .Z(n4936) );
  CND2XL U2083 ( .A(n5201), .B(n5203), .Z(n4935) );
  CENX1 U2084 ( .A(h0[14]), .B(n6417), .Z(n5294) );
  CENX1 U2085 ( .A(h0[31]), .B(n5923), .Z(n6115) );
  COND1X1 U2086 ( .A(n6588), .B(n6586), .C(n6587), .Z(n6549) );
  CND2X1 U2087 ( .A(n6586), .B(n6588), .Z(n6548) );
  COND1X1 U2088 ( .A(n6789), .B(n6790), .C(n6788), .Z(n6792) );
  CND2X1 U2089 ( .A(n6790), .B(n6789), .Z(n6791) );
  CND2X1 U2090 ( .A(n5224), .B(n5225), .Z(n4966) );
  CENX1 U2091 ( .A(n4922), .B(n7539), .Z(n1589) );
  COND2XL U2092 ( .A(n2572), .B(n1589), .C(n2489), .D(n3614), .Z(n1590) );
  CND2XL U2093 ( .A(n6191), .B(n4399), .Z(n1591) );
  COND2X1 U2094 ( .A(n7858), .B(n2573), .C(n2491), .D(n1591), .Z(n1592) );
  CEOX1 U2095 ( .A(n1590), .B(n1592), .Z(n3649) );
  CAN2X1 U2096 ( .A(n1590), .B(n1592), .Z(n3629) );
  CAN2X2 U2097 ( .A(n3451), .B(n1593), .Z(n1594) );
  CNR2XL U2098 ( .A(n5695), .B(n3454), .Z(n1595) );
  CNR2XL U2099 ( .A(n5696), .B(n3444), .Z(n1596) );
  CNR2X2 U2100 ( .A(n1595), .B(n1596), .Z(n1597) );
  CIVX2 U2101 ( .A(n3487), .Z(n1598) );
  CANR5CX4 U2102 ( .A(n1594), .B(n1597), .C(n1598), .Z(n3524) );
  CENX2 U2103 ( .A(n1597), .B(n1599), .Z(n3529) );
  CANR2XL U2104 ( .A(n2979), .B(n3173), .C(n3169), .D(n2980), .Z(n1600) );
  CANR2XL U2105 ( .A(n2995), .B(n2978), .C(n3172), .D(n2977), .Z(n1601) );
  CND2X1 U2106 ( .A(n1600), .B(n1601), .Z(n3160) );
  COND1XL U2107 ( .A(n4127), .B(n4096), .C(n4097), .Z(n1602) );
  CANR1XL U2108 ( .A(n3983), .B(n4130), .C(n1602), .Z(n4100) );
  COND1XL U2109 ( .A(n7667), .B(n4006), .C(n4007), .Z(n1603) );
  CANR1XL U2110 ( .A(n3954), .B(n7669), .C(n1603), .Z(n4027) );
  CANR2X1 U2111 ( .A(n4260), .B(n7747), .C(n7755), .D(n4246), .Z(n1604) );
  CANR2X1 U2112 ( .A(n4245), .B(n7582), .C(n7762), .D(n4261), .Z(n1605) );
  CND2X1 U2113 ( .A(n1604), .B(n1605), .Z(n4240) );
  CANR2XL U2114 ( .A(n2995), .B(n3132), .C(n3098), .D(n3172), .Z(n1606) );
  CANR2XL U2115 ( .A(n3099), .B(n3173), .C(n3130), .D(n3169), .Z(n1607) );
  CND2X1 U2116 ( .A(n1606), .B(n1607), .Z(n7557) );
  COND1XL U2117 ( .A(n7541), .B(n7675), .C(n7771), .Z(n1608) );
  COND1XL U2118 ( .A(n7729), .B(n7542), .C(n1608), .Z(n1609) );
  CND2XL U2119 ( .A(out2_2[29]), .B(n7751), .Z(n1610) );
  COND4CX1 U2120 ( .A(n7698), .B(n7543), .C(n1609), .D(n1610), .Z(n868) );
  CNR2IXL U2121 ( .B(n7804), .A(n7803), .Z(n1611) );
  CANR1XL U2122 ( .A(n7807), .B(n7806), .C(n7805), .Z(n1612) );
  CENX1 U2123 ( .A(n1611), .B(n1612), .Z(n1613) );
  CMX2XL U2124 ( .A0(out1_2[18]), .A1(n1613), .S(n8022), .Z(n7917) );
  COND1XL U2125 ( .A(n7487), .B(n7494), .C(n7008), .Z(n1614) );
  CND2XL U2126 ( .A(n7011), .B(n7492), .Z(n1615) );
  CENXL U2127 ( .A(n1615), .B(n1614), .Z(N41) );
  CNR2XL U2128 ( .A(n3691), .B(n5696), .Z(n1616) );
  CNR2XL U2129 ( .A(n3699), .B(n5695), .Z(n1617) );
  CNR2X1 U2130 ( .A(n1616), .B(n1617), .Z(n3705) );
  CND2X1 U2131 ( .A(acc[54]), .B(n2758), .Z(n1618) );
  CANR2XL U2132 ( .A(n2737), .B(out1_2[54]), .C(n2928), .D(out0_2[54]), .Z(
        n1619) );
  CND2X1 U2133 ( .A(n1618), .B(n1619), .Z(n2984) );
  CND2X1 U2134 ( .A(out2_2[10]), .B(out2_2[9]), .Z(n1620) );
  CNR2X1 U2135 ( .A(n3312), .B(n1620), .Z(n2734) );
  CANR2XL U2136 ( .A(n7552), .B(n2995), .C(n3172), .D(n3174), .Z(n1621) );
  COND1XL U2137 ( .A(n3145), .B(n7766), .C(n1621), .Z(n1622) );
  CANR1XL U2138 ( .A(n3171), .B(n3169), .C(n1622), .Z(n7743) );
  CNR2IXL U2139 ( .B(n4058), .A(n4059), .Z(n1623) );
  CNR2XL U2140 ( .A(n7816), .B(n4057), .Z(n1624) );
  CND2XL U2141 ( .A(n1624), .B(n7817), .Z(n1625) );
  COND1XL U2142 ( .A(n4057), .B(n7824), .C(n4060), .Z(n1626) );
  CANR1XL U2143 ( .A(n1624), .B(n7827), .C(n1626), .Z(n1627) );
  COND1XL U2144 ( .A(n7830), .B(n1625), .C(n1627), .Z(n1628) );
  CNR2XL U2145 ( .A(n1625), .B(n7818), .Z(n1629) );
  CANR1XL U2146 ( .A(n3949), .B(n1629), .C(n1628), .Z(n1630) );
  CENX1 U2147 ( .A(n1623), .B(n1630), .Z(n1631) );
  CMX2XL U2148 ( .A0(out1_2[61]), .A1(n1631), .S(n7846), .Z(n7874) );
  CND2XL U2149 ( .A(n4212), .B(n4211), .Z(n1632) );
  CENX1 U2150 ( .A(n7806), .B(n1632), .Z(n1633) );
  CMX2XL U2151 ( .A0(out1_2[16]), .A1(n1633), .S(n8022), .Z(n7919) );
  CNR2X1 U2152 ( .A(n7693), .B(n7727), .Z(n1634) );
  COND2X1 U2153 ( .A(n7729), .B(n3116), .C(n7724), .D(n7692), .Z(n1635) );
  CND2XL U2154 ( .A(out2_2[30]), .B(n7751), .Z(n1636) );
  COND11X1 U2155 ( .A(n3075), .B(n1634), .C(n1635), .D(n1636), .Z(n2862) );
  CND2X1 U2156 ( .A(acc[49]), .B(n2758), .Z(n1637) );
  CANR2XL U2157 ( .A(n2737), .B(out1_2[49]), .C(n2928), .D(out0_2[49]), .Z(
        n1638) );
  CND2X1 U2158 ( .A(n1637), .B(n1638), .Z(n2969) );
  CND2X1 U2159 ( .A(acc[53]), .B(n2758), .Z(n1639) );
  CANR2XL U2160 ( .A(n2737), .B(out1_2[53]), .C(n2928), .D(out0_2[53]), .Z(
        n1640) );
  CND2X1 U2161 ( .A(n1639), .B(n1640), .Z(n2983) );
  CNR2IX1 U2162 ( .B(n4291), .A(n4292), .Z(n4298) );
  CANR2XL U2163 ( .A(n3018), .B(n2995), .C(n3019), .D(n3169), .Z(n1641) );
  CANR2XL U2164 ( .A(n2989), .B(n3173), .C(n2988), .D(n3172), .Z(n1642) );
  CND2X1 U2165 ( .A(n1641), .B(n1642), .Z(n3039) );
  CANR2XL U2166 ( .A(n2984), .B(n2995), .C(n3173), .D(n2980), .Z(n1643) );
  CANR2XL U2167 ( .A(n3169), .B(n2982), .C(n3172), .D(n2978), .Z(n1644) );
  CND2X1 U2168 ( .A(n1643), .B(n1644), .Z(n3035) );
  CANR2XL U2169 ( .A(n2974), .B(n3173), .C(n2973), .D(n3169), .Z(n1645) );
  CANR2XL U2170 ( .A(n2975), .B(n2995), .C(n2976), .D(n3172), .Z(n1646) );
  CND2X1 U2171 ( .A(n1645), .B(n1646), .Z(n3161) );
  CNR2IXL U2172 ( .B(n4009), .A(n4008), .Z(n1647) );
  CNR2IXL U2173 ( .B(n4119), .A(n4115), .Z(n1648) );
  CND2XL U2174 ( .A(n1648), .B(n7817), .Z(n1649) );
  CIVXL U2175 ( .A(n4118), .Z(n1650) );
  COND1XL U2176 ( .A(n4115), .B(n1650), .C(n4116), .Z(n1651) );
  CANR1XL U2177 ( .A(n1648), .B(n7827), .C(n1651), .Z(n1652) );
  COND1XL U2178 ( .A(n7830), .B(n1649), .C(n1652), .Z(n1653) );
  CNR2XL U2179 ( .A(n1649), .B(n7818), .Z(n1654) );
  CANR1XL U2180 ( .A(n3949), .B(n1654), .C(n1653), .Z(n1655) );
  CENX1 U2181 ( .A(n1647), .B(n1655), .Z(n1656) );
  CMX2XL U2182 ( .A0(out1_2[59]), .A1(n1656), .S(n7846), .Z(n7876) );
  CIVXL U2183 ( .A(n4228), .Z(n1657) );
  CIVXL U2184 ( .A(n7792), .Z(n1658) );
  CNR2IXL U2185 ( .B(n4226), .A(n4230), .Z(n1659) );
  COND4CXL U2186 ( .A(n4227), .B(n1658), .C(n4231), .D(n1659), .Z(n1660) );
  COND3XL U2187 ( .A(n4230), .B(n1657), .C(n4229), .D(n1660), .Z(n1661) );
  CND2IXL U2188 ( .B(n4232), .A(n4233), .Z(n1662) );
  CENX1 U2189 ( .A(n1661), .B(n1662), .Z(n1663) );
  CMX2XL U2190 ( .A0(out1_2[15]), .A1(n1663), .S(cmd1_en_2), .Z(n7920) );
  COND2XL U2191 ( .A(n7770), .B(n7765), .C(n7766), .D(n7748), .Z(n1664) );
  COND2X1 U2192 ( .A(n7763), .B(n7769), .C(n7764), .D(n2663), .Z(n1665) );
  CANR4CX1 U2193 ( .A(n1664), .B(n1665), .C(n7772), .D(n7771), .Z(n1666) );
  CIVX1 U2194 ( .A(n7743), .Z(n1667) );
  COND2XL U2195 ( .A(n2662), .B(n7745), .C(n7744), .D(n1667), .Z(n1668) );
  COND4CXL U2196 ( .A(n7746), .B(n7747), .C(n1668), .D(n8020), .Z(n1669) );
  COND3X1 U2197 ( .A(n8020), .B(n7750), .C(n1666), .D(n1669), .Z(n1670) );
  CANR2X1 U2198 ( .A(n7751), .B(out2_2[1]), .C(n7778), .D(n7752), .Z(n1671) );
  CND2X1 U2199 ( .A(n7780), .B(n7753), .Z(n1672) );
  CND3XL U2200 ( .A(n1672), .B(n1671), .C(n1670), .Z(n865) );
  CANR5CXL U2201 ( .A(n1699), .B(n1698), .C(n1697), .Z(n1673) );
  CIVX2 U2202 ( .A(n1673), .Z(n3610) );
  CND2X1 U2203 ( .A(acc[56]), .B(n2758), .Z(n1674) );
  CANR2XL U2204 ( .A(n2737), .B(out1_2[56]), .C(n2928), .D(out0_2[56]), .Z(
        n1675) );
  CND2X1 U2205 ( .A(n1674), .B(n1675), .Z(n2978) );
  CENXL U2206 ( .A(n1817), .B(n1818), .Z(n1676) );
  CENXL U2207 ( .A(n3690), .B(n1676), .Z(n3709) );
  CNR2IXL U2208 ( .B(n3270), .A(n3285), .Z(n4316) );
  CANR2XL U2209 ( .A(n3173), .B(n3009), .C(n3169), .D(n3008), .Z(n1677) );
  CANR2XL U2210 ( .A(n2995), .B(n3011), .C(n3172), .D(n3010), .Z(n1678) );
  CND2XL U2211 ( .A(n1677), .B(n1678), .Z(n3164) );
  CANR2XL U2212 ( .A(n2983), .B(n3169), .C(n3172), .D(n2984), .Z(n1679) );
  CANR2XL U2213 ( .A(n3173), .B(n2982), .C(n2995), .D(n2981), .Z(n1680) );
  CND2X1 U2214 ( .A(n1679), .B(n1680), .Z(n3159) );
  CANR2X1 U2215 ( .A(n3173), .B(n2967), .C(n2969), .D(n3172), .Z(n1681) );
  CANR2XL U2216 ( .A(n2997), .B(n2995), .C(n2968), .D(n3169), .Z(n1682) );
  CND2X1 U2217 ( .A(n1681), .B(n1682), .Z(n4262) );
  CANR2XL U2218 ( .A(n2737), .B(out1_2[4]), .C(n2928), .D(out0_2[4]), .Z(n1683) );
  COND1XL U2219 ( .A(n2670), .B(n2961), .C(n1683), .Z(n7748) );
  CNR2IXL U2220 ( .B(n4144), .A(n4143), .Z(n1684) );
  CND2XL U2221 ( .A(n4146), .B(n7817), .Z(n1685) );
  CNR2XL U2222 ( .A(n1685), .B(n7818), .Z(n1686) );
  CND2XL U2223 ( .A(n4146), .B(n7827), .Z(n1687) );
  COND3XL U2224 ( .A(n7830), .B(n1685), .C(n4145), .D(n1687), .Z(n1688) );
  CANR1XL U2225 ( .A(n3949), .B(n1686), .C(n1688), .Z(n1689) );
  CENX1 U2226 ( .A(n1684), .B(n1689), .Z(n1690) );
  CMX2XL U2227 ( .A0(out1_2[57]), .A1(n1690), .S(n7846), .Z(n7878) );
  COND2XL U2228 ( .A(n7556), .B(n3189), .C(n4254), .D(n3113), .Z(n1691) );
  COND1XL U2229 ( .A(n3175), .B(n7557), .C(n8019), .Z(n1692) );
  CANR3X1 U2230 ( .A(n4249), .B(n7559), .C(n1691), .D(n1692), .Z(n1693) );
  CND3XL U2231 ( .A(n3054), .B(n3053), .C(n7543), .Z(n1694) );
  COND3X1 U2232 ( .A(n7739), .B(n4266), .C(n1693), .D(n1694), .Z(n1695) );
  CND2X1 U2233 ( .A(n7751), .B(out2_2[6]), .Z(n1696) );
  COND4CX1 U2234 ( .A(n4272), .B(n7741), .C(n1695), .D(n1696), .Z(n3052) );
  COND2XL U2235 ( .A(n5695), .B(n3616), .C(n4886), .D(n3585), .Z(n1697) );
  COND2X1 U2236 ( .A(n5912), .B(n3584), .C(n4443), .D(n3617), .Z(n1698) );
  COND2XL U2237 ( .A(n2569), .B(n3614), .C(n2490), .D(n3583), .Z(n1699) );
  CENX1 U2238 ( .A(n1697), .B(n1698), .Z(n1700) );
  CENX1 U2239 ( .A(n1699), .B(n1700), .Z(n3636) );
  CND2X1 U2240 ( .A(acc[51]), .B(n2758), .Z(n1701) );
  CANR2XL U2241 ( .A(n2737), .B(out1_2[51]), .C(n2928), .D(out0_2[51]), .Z(
        n1702) );
  CND2X1 U2242 ( .A(n1701), .B(n1702), .Z(n2970) );
  CND2X1 U2243 ( .A(acc[60]), .B(n2758), .Z(n1703) );
  CANR2XL U2244 ( .A(n2737), .B(out1_2[60]), .C(n2928), .D(out0_2[60]), .Z(
        n1704) );
  CND2X1 U2245 ( .A(n1703), .B(n1704), .Z(n2975) );
  CIVX1 U2246 ( .A(n2708), .Z(n1705) );
  CNR3X1 U2247 ( .A(n4292), .B(n3225), .C(n1705), .Z(n3279) );
  CANR2XL U2248 ( .A(n3173), .B(n3100), .C(n3099), .D(n3172), .Z(n1706) );
  CANR2XL U2249 ( .A(n3130), .B(n2995), .C(n3098), .D(n3169), .Z(n1707) );
  CND2X1 U2250 ( .A(n1706), .B(n1707), .Z(n3078) );
  CANR2X1 U2251 ( .A(n2987), .B(n2995), .C(n3169), .D(n2994), .Z(n1708) );
  CANR2X1 U2252 ( .A(n2993), .B(n3173), .C(n3172), .D(n2996), .Z(n1709) );
  CND2X1 U2253 ( .A(n1708), .B(n1709), .Z(n4260) );
  CND2IX1 U2254 ( .B(h0_1[1]), .A(h0_1[0]), .Z(n7763) );
  CIVXL U2255 ( .A(n7830), .Z(n1710) );
  CANR1XL U2256 ( .A(n7817), .B(n1710), .C(n7827), .Z(n1711) );
  CND2XL U2257 ( .A(n7817), .B(n3949), .Z(n1712) );
  COND1XL U2258 ( .A(n7818), .B(n1712), .C(n1711), .Z(n1713) );
  CND2XL U2259 ( .A(n4146), .B(n4145), .Z(n1714) );
  CENX1 U2260 ( .A(n1713), .B(n1714), .Z(n1715) );
  CMX2XL U2261 ( .A0(out1_2[56]), .A1(n1715), .S(n7846), .Z(n7879) );
  CIVXL U2262 ( .A(n7792), .Z(n1716) );
  COND4CXL U2263 ( .A(n4227), .B(n1716), .C(n4231), .D(n4219), .Z(n1717) );
  CND2XL U2264 ( .A(n4218), .B(n1717), .Z(n1718) );
  CND2IXL U2265 ( .B(n4214), .A(n4215), .Z(n1719) );
  CENX1 U2266 ( .A(n1718), .B(n1719), .Z(n1720) );
  CMX2XL U2267 ( .A0(out1_2[13]), .A1(n1720), .S(cmd1_en_2), .Z(n7922) );
  CANR5CXL U2268 ( .A(n6677), .B(n1798), .C(n1799), .Z(n1721) );
  CIVX1 U2269 ( .A(n1721), .Z(n6724) );
  CND2X1 U2270 ( .A(acc[50]), .B(n2758), .Z(n1722) );
  CANR2XL U2271 ( .A(n2737), .B(out1_2[50]), .C(n2928), .D(out0_2[50]), .Z(
        n1723) );
  CND2X1 U2272 ( .A(n1722), .B(n1723), .Z(n2967) );
  CND2X1 U2273 ( .A(acc[42]), .B(n2758), .Z(n1724) );
  CANR2XL U2274 ( .A(n2737), .B(out1_2[42]), .C(n2928), .D(out0_2[42]), .Z(
        n1725) );
  CND2X1 U2275 ( .A(n1724), .B(n1725), .Z(n2990) );
  CND2X1 U2276 ( .A(acc[61]), .B(n2758), .Z(n1726) );
  CANR2XL U2277 ( .A(n2737), .B(out1_2[61]), .C(n2928), .D(out0_2[61]), .Z(
        n1727) );
  CND2X1 U2278 ( .A(n1726), .B(n1727), .Z(n2973) );
  CND2XL U2279 ( .A(n5566), .B(n4399), .Z(n1728) );
  COND2XL U2280 ( .A(n7862), .B(n5695), .C(n5696), .D(n1728), .Z(n3700) );
  CANR2XL U2281 ( .A(n3173), .B(n2975), .C(n2977), .D(n3169), .Z(n1729) );
  CANR2XL U2282 ( .A(n3172), .B(n2979), .C(n2980), .D(n2995), .Z(n1730) );
  CND2X1 U2283 ( .A(n1729), .B(n1730), .Z(n3122) );
  CANR2X1 U2284 ( .A(n3009), .B(n2995), .C(n3169), .D(n3003), .Z(n1731) );
  CANR2X1 U2285 ( .A(n3005), .B(n3173), .C(n3172), .D(n3004), .Z(n1732) );
  CND2X1 U2286 ( .A(n1731), .B(n1732), .Z(n4245) );
  CANR2X1 U2287 ( .A(n2970), .B(n2995), .C(n3169), .D(n2981), .Z(n1733) );
  CANR2X1 U2288 ( .A(n2984), .B(n3173), .C(n3172), .D(n2983), .Z(n1734) );
  CND2X1 U2289 ( .A(n1733), .B(n1734), .Z(n4263) );
  CAOR2XL U2290 ( .A(out0_2[1]), .B(n2928), .C(n2737), .D(out1_2[1]), .Z(n1735) );
  CANR1XL U2291 ( .A(n2758), .B(acc[1]), .C(n1735), .Z(n7749) );
  CANR2XL U2292 ( .A(n2995), .B(n3013), .C(n3172), .D(n3012), .Z(n1736) );
  CANR2XL U2293 ( .A(n3169), .B(n3015), .C(n3173), .D(n3014), .Z(n1737) );
  CND2XL U2294 ( .A(n1736), .B(n1737), .Z(n3162) );
  CND2IXL U2295 ( .B(n7228), .A(n6978), .Z(n1738) );
  CND2IXL U2296 ( .B(n2382), .A(n6976), .Z(n1739) );
  CND2X2 U2297 ( .A(n1738), .B(n1739), .Z(n7081) );
  CENXL U2298 ( .A(n5566), .B(n7539), .Z(n1740) );
  COND2XL U2299 ( .A(n4886), .B(n3699), .C(n5695), .D(n1740), .Z(n1770) );
  CIVX1 U2300 ( .A(n2719), .Z(n1741) );
  CND4X1 U2301 ( .A(out2_2[54]), .B(out2_2[53]), .C(n2717), .D(n1741), .Z(
        n2726) );
  CNR2IX1 U2302 ( .B(n3242), .A(n4292), .Z(n3248) );
  CANR5CXL U2303 ( .A(n1817), .B(n1818), .C(n3690), .Z(n1742) );
  CIVXL U2304 ( .A(n1742), .Z(n3710) );
  CANR5CXL U2305 ( .A(n3606), .B(n3603), .C(n3604), .Z(n1743) );
  CIVX1 U2306 ( .A(n1743), .Z(n3730) );
  CANR2XL U2307 ( .A(n2990), .B(n2995), .C(n3173), .D(n2996), .Z(n1744) );
  CANR2XL U2308 ( .A(n3169), .B(n2987), .C(n3172), .D(n2994), .Z(n1745) );
  CND2X1 U2309 ( .A(n1744), .B(n1745), .Z(n3038) );
  CANR2XL U2310 ( .A(n2995), .B(n3012), .C(n3008), .D(n3173), .Z(n1746) );
  CANR2XL U2311 ( .A(n3172), .B(n3011), .C(n3014), .D(n3169), .Z(n1747) );
  CND2X1 U2312 ( .A(n1746), .B(n1747), .Z(n3114) );
  CNR2IXL U2313 ( .B(n4136), .A(n4135), .Z(n1748) );
  CNR2IXL U2314 ( .B(n4137), .A(n4141), .Z(n1749) );
  CND2XL U2315 ( .A(n4138), .B(n1749), .Z(n1750) );
  CNR2XL U2316 ( .A(n1750), .B(n7818), .Z(n1751) );
  CIVXL U2317 ( .A(n4139), .Z(n1752) );
  COND1XL U2318 ( .A(n4141), .B(n1752), .C(n4140), .Z(n1753) );
  CANR1XL U2319 ( .A(n1749), .B(n4142), .C(n1753), .Z(n1754) );
  COND1XL U2320 ( .A(n7830), .B(n1750), .C(n1754), .Z(n1755) );
  CANR1XL U2321 ( .A(n3949), .B(n1751), .C(n1755), .Z(n1756) );
  CENX1 U2322 ( .A(n1748), .B(n1756), .Z(n1757) );
  CMX2XL U2323 ( .A0(out1_2[55]), .A1(n1757), .S(n7846), .Z(n7880) );
  COND1XL U2324 ( .A(n4217), .B(n7792), .C(n4216), .Z(n1758) );
  CND2XL U2325 ( .A(n4219), .B(n4218), .Z(n1759) );
  CENX1 U2326 ( .A(n1758), .B(n1759), .Z(n1760) );
  CMX2XL U2327 ( .A0(out1_2[12]), .A1(n1760), .S(cmd1_en_2), .Z(n7923) );
  CANR11XL U2328 ( .A(n3154), .B(n3155), .C(n3074), .D(n3075), .Z(n1761) );
  COND1XL U2329 ( .A(n7727), .B(n3152), .C(n1761), .Z(n1762) );
  CND2X1 U2330 ( .A(n7751), .B(out2_2[24]), .Z(n1763) );
  COND4CXL U2331 ( .A(n7771), .B(n7685), .C(n1762), .D(n1763), .Z(n3023) );
  CANR5CXL U2332 ( .A(n1851), .B(n1852), .C(n6975), .Z(n1764) );
  CIVX1 U2333 ( .A(n1764), .Z(n7067) );
  CNR2XL U2334 ( .A(n7537), .B(n3634), .Z(n1765) );
  CNR2XL U2335 ( .A(n5160), .B(n3659), .Z(n1766) );
  CNR2X1 U2336 ( .A(n1765), .B(n1766), .Z(n1807) );
  CND2X1 U2337 ( .A(acc[44]), .B(n2758), .Z(n1767) );
  CANR2XL U2338 ( .A(n2737), .B(out1_2[44]), .C(n2928), .D(out0_2[44]), .Z(
        n1768) );
  CND2X1 U2339 ( .A(n1767), .B(n1768), .Z(n2994) );
  COND2XL U2340 ( .A(n7537), .B(n3697), .C(n5160), .D(n3698), .Z(n1769) );
  CEOXL U2341 ( .A(n1769), .B(n1770), .Z(n3701) );
  CAN2XL U2342 ( .A(n1769), .B(n1770), .Z(n3706) );
  CNR2IX1 U2343 ( .B(n3213), .A(n3321), .Z(n3295) );
  CENX1 U2344 ( .A(n3684), .B(n3683), .Z(n1771) );
  CENX1 U2345 ( .A(n3685), .B(n1771), .Z(n3711) );
  CND2XL U2346 ( .A(n2995), .B(n2973), .Z(n1772) );
  CANR2XL U2347 ( .A(n2974), .B(n3172), .C(n2976), .D(n3169), .Z(n1773) );
  CND2X1 U2348 ( .A(n1772), .B(n1773), .Z(n3118) );
  CND2IX1 U2349 ( .B(n3312), .A(n3339), .Z(n3332) );
  CND2IX1 U2350 ( .B(n2729), .A(n4281), .Z(n3258) );
  COND1XL U2351 ( .A(n4221), .B(n4224), .C(n4225), .Z(n1774) );
  CANR1XL U2352 ( .A(n3909), .B(n4222), .C(n1774), .Z(n4216) );
  CNR2XL U2353 ( .A(n3145), .B(n2663), .Z(n1775) );
  COND2XL U2354 ( .A(n3143), .B(n7763), .C(n7770), .D(n3144), .Z(n1776) );
  CANR3XL U2355 ( .A(n3146), .B(n3173), .C(n1775), .D(n1776), .Z(n7761) );
  CNR2IXL U2356 ( .B(n4112), .A(n4111), .Z(n1777) );
  CND2XL U2357 ( .A(n4114), .B(n4138), .Z(n1778) );
  CNR2XL U2358 ( .A(n1778), .B(n7818), .Z(n1779) );
  CND2XL U2359 ( .A(n4114), .B(n4142), .Z(n1780) );
  COND3XL U2360 ( .A(n7830), .B(n1778), .C(n4113), .D(n1780), .Z(n1781) );
  CANR1XL U2361 ( .A(n3949), .B(n1779), .C(n1781), .Z(n1782) );
  CENX1 U2362 ( .A(n1777), .B(n1782), .Z(n1783) );
  CMX2XL U2363 ( .A0(out1_2[53]), .A1(n1783), .S(n7846), .Z(n7882) );
  CNR2IXL U2364 ( .B(n4235), .A(n4234), .Z(n1784) );
  CIVXL U2365 ( .A(n7785), .Z(n1785) );
  CIVXL U2366 ( .A(n7787), .Z(n1786) );
  COND1XL U2367 ( .A(n7785), .B(n1786), .C(n7786), .Z(n1787) );
  CANR11XL U2368 ( .A(n7788), .B(n7789), .C(n1785), .D(n1787), .Z(n1788) );
  CENX1 U2369 ( .A(n1784), .B(n1788), .Z(n1789) );
  CMX2XL U2370 ( .A0(out1_2[7]), .A1(n1789), .S(n8022), .Z(n7928) );
  CND2XL U2371 ( .A(n3082), .B(n3074), .Z(n1790) );
  COND2X1 U2372 ( .A(n3084), .B(n1790), .C(n7727), .D(n3085), .Z(n1791) );
  CANR3X1 U2373 ( .A(n7684), .B(n7771), .C(n3075), .D(n1791), .Z(n1792) );
  CAOR1X1 U2374 ( .A(out2_2[27]), .B(n7751), .C(n1792), .Z(n3076) );
  CANR5CXL U2375 ( .A(n6889), .B(n6890), .C(n6888), .Z(n1793) );
  CIVXL U2376 ( .A(n1793), .Z(n6988) );
  COND2X1 U2377 ( .A(n7537), .B(n4393), .C(n5160), .D(n3778), .Z(n1794) );
  COND2XL U2378 ( .A(n6114), .B(n3777), .C(n3368), .D(n4515), .Z(n1795) );
  CENX1 U2379 ( .A(n4458), .B(n1794), .Z(n1796) );
  CENX1 U2380 ( .A(n1795), .B(n1796), .Z(n4560) );
  CANR5CXL U2381 ( .A(n4458), .B(n1794), .C(n1795), .Z(n1797) );
  CIVXL U2382 ( .A(n1797), .Z(n4591) );
  COND2X1 U2383 ( .A(n6703), .B(n6648), .C(n2514), .D(n6704), .Z(n1798) );
  COND2X1 U2384 ( .A(n2294), .B(n6649), .C(n7114), .D(n6670), .Z(n1799) );
  CENX1 U2385 ( .A(n6677), .B(n1798), .Z(n1800) );
  CENX1 U2386 ( .A(n1799), .B(n1800), .Z(n6693) );
  CIVX2 U2387 ( .A(n6604), .Z(n1801) );
  CND2XL U2388 ( .A(n6607), .B(n6606), .Z(n1802) );
  COND1X4 U2389 ( .A(n1801), .B(n6605), .C(n1802), .Z(n6904) );
  CENXL U2390 ( .A(n1963), .B(n1962), .Z(n1803) );
  CENXL U2391 ( .A(n7059), .B(n1803), .Z(n7068) );
  COND2X1 U2392 ( .A(n6523), .B(n3517), .C(n6211), .D(n3518), .Z(n1804) );
  CND2XL U2393 ( .A(n6417), .B(n4399), .Z(n1805) );
  COND2X1 U2394 ( .A(n6211), .B(n2606), .C(n6523), .D(n1805), .Z(n1806) );
  CEOX1 U2395 ( .A(n1804), .B(n1806), .Z(n3607) );
  CAN2X2 U2396 ( .A(n1804), .B(n1806), .Z(n3593) );
  CND2IXL U2397 ( .B(n2488), .A(n7539), .Z(n1808) );
  CIVXL U2398 ( .A(n3665), .Z(n1809) );
  CANR5CX1 U2399 ( .A(n1807), .B(n1808), .C(n1809), .Z(n3648) );
  CENXL U2400 ( .A(n1807), .B(n3665), .Z(n1810) );
  CENX1 U2401 ( .A(n1808), .B(n1810), .Z(n3666) );
  CND2XL U2402 ( .A(acc[48]), .B(n2758), .Z(n1811) );
  CANR2XL U2403 ( .A(n2737), .B(out1_2[48]), .C(n2928), .D(out0_2[48]), .Z(
        n1812) );
  CND2X1 U2404 ( .A(n1811), .B(n1812), .Z(n2968) );
  CND2XL U2405 ( .A(acc[52]), .B(n2758), .Z(n1813) );
  CANR2XL U2406 ( .A(n2737), .B(out1_2[52]), .C(n2928), .D(out0_2[52]), .Z(
        n1814) );
  CND2X1 U2407 ( .A(n1813), .B(n1814), .Z(n2981) );
  CND2XL U2408 ( .A(acc[57]), .B(n2758), .Z(n1815) );
  CANR2XL U2409 ( .A(n2737), .B(out1_2[57]), .C(n2928), .D(out0_2[57]), .Z(
        n1816) );
  CND2X1 U2410 ( .A(n1815), .B(n1816), .Z(n2980) );
  COND2XL U2411 ( .A(n5696), .B(n3689), .C(n5695), .D(n3691), .Z(n1817) );
  COND2XL U2412 ( .A(n7537), .B(n3686), .C(n5160), .D(n3693), .Z(n1818) );
  CANR2XL U2413 ( .A(n3017), .B(n3173), .C(n3002), .D(n3169), .Z(n1819) );
  CANR2XL U2414 ( .A(n3005), .B(n2995), .C(n3020), .D(n3172), .Z(n1820) );
  CND2XL U2415 ( .A(n1819), .B(n1820), .Z(n3051) );
  CANR2XL U2416 ( .A(n2983), .B(n2995), .C(n3169), .D(n2984), .Z(n1821) );
  CANR2XL U2417 ( .A(n3173), .B(n2978), .C(n3172), .D(n2982), .Z(n1822) );
  CND2X1 U2418 ( .A(n1821), .B(n1822), .Z(n3136) );
  CANR2X1 U2419 ( .A(n2973), .B(n3172), .C(n2976), .D(n3173), .Z(n1823) );
  CANR2X1 U2420 ( .A(n2975), .B(n3169), .C(n2979), .D(n2995), .Z(n1824) );
  CND2X1 U2421 ( .A(n1823), .B(n1824), .Z(n3065) );
  CND2IX1 U2422 ( .B(n3268), .A(n3269), .Z(n3285) );
  CND2IX1 U2423 ( .B(n2719), .A(n3253), .Z(n3290) );
  COND1XL U2424 ( .A(n4199), .B(n4195), .C(n4196), .Z(n1825) );
  CANR1XL U2425 ( .A(n4183), .B(n3929), .C(n1825), .Z(n1826) );
  COND1XL U2426 ( .A(n3930), .B(n4177), .C(n1826), .Z(n7569) );
  CND2IX1 U2427 ( .B(n2735), .A(n3313), .Z(n3218) );
  CANR2X1 U2428 ( .A(n7755), .B(n7584), .C(n7583), .D(n7762), .Z(n1827) );
  CANR2XL U2429 ( .A(n7582), .B(n7580), .C(n7577), .D(n7747), .Z(n1828) );
  CND2XL U2430 ( .A(n1827), .B(n1828), .Z(n3091) );
  CANR2XL U2431 ( .A(n3172), .B(n3132), .C(n3131), .D(n2995), .Z(n1829) );
  CANR2XL U2432 ( .A(n3130), .B(n3173), .C(n3129), .D(n3169), .Z(n1830) );
  CND2X1 U2433 ( .A(n1829), .B(n1830), .Z(n7759) );
  CIVXL U2434 ( .A(n3311), .Z(n1831) );
  CANR2XL U2435 ( .A(n4363), .B(out1_2[10]), .C(n1430), .D(n4350), .Z(n1832)
         );
  CNR2X1 U2436 ( .A(n3332), .B(n3333), .Z(n1833) );
  CEOX1 U2437 ( .A(n1833), .B(out2_2[10]), .Z(n1834) );
  CND2X1 U2438 ( .A(n4344), .B(n1834), .Z(n1835) );
  COND3XL U2439 ( .A(n2685), .B(n1831), .C(n1832), .D(n1835), .Z(n1003) );
  CND2X1 U2440 ( .A(cmd0[1]), .B(push0), .Z(n1836) );
  CNR2X1 U2441 ( .A(cmd0[0]), .B(n1836), .Z(cmd2_en_0) );
  CNR2IXL U2442 ( .B(n4097), .A(n4096), .Z(n1837) );
  CND2XL U2443 ( .A(n4128), .B(n4129), .Z(n1838) );
  CNR2XL U2444 ( .A(n1838), .B(n7818), .Z(n1839) );
  CND2XL U2445 ( .A(n4128), .B(n4130), .Z(n1840) );
  COND3XL U2446 ( .A(n7830), .B(n1838), .C(n4127), .D(n1840), .Z(n1841) );
  CANR1XL U2447 ( .A(n3949), .B(n1839), .C(n1841), .Z(n1842) );
  CENX1 U2448 ( .A(n1837), .B(n1842), .Z(n1843) );
  CMX2XL U2449 ( .A0(out1_2[51]), .A1(n1843), .S(n7846), .Z(n7884) );
  CNR2IXL U2450 ( .B(n7786), .A(n7785), .Z(n1844) );
  CANR1XL U2451 ( .A(n7789), .B(n7788), .C(n7787), .Z(n1845) );
  CENX1 U2452 ( .A(n1844), .B(n1845), .Z(n1846) );
  CMX2XL U2453 ( .A0(out1_2[6]), .A1(n1846), .S(n8022), .Z(n7929) );
  CNR2XL U2454 ( .A(n3134), .B(n7727), .Z(n1847) );
  CANR3X1 U2455 ( .A(n7683), .B(n7771), .C(n1847), .D(n3075), .Z(n1848) );
  COND1XL U2456 ( .A(n7729), .B(n3133), .C(n1848), .Z(n1849) );
  COND1XL U2457 ( .A(n2865), .B(n4310), .C(n1849), .Z(n3071) );
  CND2XL U2458 ( .A(n6380), .B(n6378), .Z(n1850) );
  CENX1 U2459 ( .A(n6379), .B(n1850), .Z(N30) );
  COND2X1 U2460 ( .A(n2433), .B(n6980), .C(n2282), .D(n6867), .Z(n1851) );
  COND2XL U2461 ( .A(n7228), .B(n6865), .C(n2381), .D(n6977), .Z(n1852) );
  CENX1 U2462 ( .A(n6975), .B(n1851), .Z(n1853) );
  CENX1 U2463 ( .A(n1852), .B(n1853), .Z(n6982) );
  COND2X1 U2464 ( .A(n6293), .B(n3500), .C(n3501), .D(n6211), .Z(n1854) );
  COND2X1 U2465 ( .A(n5912), .B(n3497), .C(n5911), .D(n3511), .Z(n1855) );
  CENX1 U2466 ( .A(n3520), .B(n1854), .Z(n1856) );
  CENX1 U2467 ( .A(n1855), .B(n1856), .Z(n3559) );
  CANR5CX1 U2468 ( .A(n3520), .B(n1854), .C(n1855), .Z(n1857) );
  CIVX1 U2469 ( .A(n1857), .Z(n3503) );
  CENXL U2470 ( .A(n2026), .B(n4557), .Z(n1858) );
  CENX1 U2471 ( .A(n2025), .B(n1858), .Z(n4612) );
  CND2X1 U2472 ( .A(n6902), .B(n6903), .Z(n1859) );
  CND2X2 U2473 ( .A(n2303), .B(n1859), .Z(n1860) );
  CENX2 U2474 ( .A(n6904), .B(n1860), .Z(n6916) );
  CND2X2 U2475 ( .A(n1861), .B(n3635), .Z(n3637) );
  CND2XL U2476 ( .A(acc[47]), .B(n2758), .Z(n1862) );
  CANR2XL U2477 ( .A(n2737), .B(out1_2[47]), .C(n2928), .D(out0_2[47]), .Z(
        n1863) );
  CND2X1 U2478 ( .A(n1862), .B(n1863), .Z(n2997) );
  CND2XL U2479 ( .A(acc[59]), .B(n2758), .Z(n1864) );
  CANR2XL U2480 ( .A(n2737), .B(out1_2[59]), .C(n2928), .D(out0_2[59]), .Z(
        n1865) );
  CND2X1 U2481 ( .A(n1864), .B(n1865), .Z(n2979) );
  CMXI2XL U2482 ( .A0(n2976), .A1(n2974), .S(h0_1[0]), .Z(n1866) );
  COR2X1 U2483 ( .A(h0_1[1]), .B(n1866), .Z(n3037) );
  CANR2X1 U2484 ( .A(n3018), .B(n3173), .C(n3172), .D(n3017), .Z(n1867) );
  CANR2X1 U2485 ( .A(n3002), .B(n2995), .C(n3169), .D(n3020), .Z(n1868) );
  CND2X1 U2486 ( .A(n1867), .B(n1868), .Z(n4246) );
  CANR2X1 U2487 ( .A(n2982), .B(n2995), .C(n3169), .D(n2978), .Z(n1869) );
  CANR2X1 U2488 ( .A(n2977), .B(n3173), .C(n3172), .D(n2980), .Z(n1870) );
  CND2X1 U2489 ( .A(n1869), .B(n1870), .Z(n3066) );
  CND2X1 U2490 ( .A(n7536), .B(n7535), .Z(n1871) );
  CND2X2 U2491 ( .A(n1871), .B(n7534), .Z(n4278) );
  COND1XL U2492 ( .A(n4116), .B(n4008), .C(n4009), .Z(n1872) );
  CANR1XL U2493 ( .A(n3996), .B(n4118), .C(n1872), .Z(n7824) );
  COND1XL U2494 ( .A(n7804), .B(n7793), .C(n7794), .Z(n1873) );
  CANR1XL U2495 ( .A(n7805), .B(n3924), .C(n1873), .Z(n4177) );
  CND2IX1 U2496 ( .B(n2945), .A(n4353), .Z(n4286) );
  CENX1 U2497 ( .A(n3548), .B(n3547), .Z(n1874) );
  CND2X1 U2498 ( .A(n1874), .B(n3740), .Z(n6373) );
  CIVXL U2499 ( .A(n4383), .Z(n1875) );
  CANR2XL U2500 ( .A(n4363), .B(out1_2[12]), .C(n1422), .D(n4350), .Z(n1876)
         );
  CNR2X1 U2501 ( .A(n3319), .B(n3318), .Z(n1877) );
  CENX1 U2502 ( .A(n3320), .B(n1877), .Z(n1878) );
  CND2X1 U2503 ( .A(n4344), .B(n1878), .Z(n1879) );
  COND3XL U2504 ( .A(n2685), .B(n1875), .C(n1876), .D(n1879), .Z(n1005) );
  CANR2XL U2505 ( .A(n4363), .B(out1_2[16]), .C(acc[16]), .D(n4350), .Z(n1880)
         );
  CNR2X1 U2506 ( .A(n3321), .B(n8002), .Z(n1881) );
  CENX1 U2507 ( .A(n8001), .B(n1881), .Z(n1882) );
  CND2X1 U2508 ( .A(n4344), .B(n1882), .Z(n1883) );
  CIVX1 U2509 ( .A(n3340), .Z(n1884) );
  CANR2XL U2510 ( .A(n4363), .B(n1361), .C(acc[2]), .D(n4350), .Z(n1885) );
  CNR2X1 U2511 ( .A(n4364), .B(n3341), .Z(n1886) );
  CEOX1 U2512 ( .A(n1886), .B(out2_2[2]), .Z(n1887) );
  CND2X1 U2513 ( .A(n4344), .B(n1887), .Z(n1888) );
  COND3XL U2514 ( .A(n2685), .B(n1884), .C(n1885), .D(n1888), .Z(n995) );
  CIVXL U2515 ( .A(n7830), .Z(n1889) );
  CANR1XL U2516 ( .A(n4129), .B(n1889), .C(n4130), .Z(n1890) );
  CND2X1 U2517 ( .A(n3949), .B(n4129), .Z(n1891) );
  COND1XL U2518 ( .A(n7818), .B(n1891), .C(n1890), .Z(n1892) );
  CND2XL U2519 ( .A(n4128), .B(n4127), .Z(n1893) );
  CENX1 U2520 ( .A(n1892), .B(n1893), .Z(n1894) );
  CMX2XL U2521 ( .A0(out1_2[50]), .A1(n1894), .S(n7846), .Z(n7885) );
  CND2XL U2522 ( .A(n4223), .B(n4220), .Z(n1895) );
  CND2XL U2523 ( .A(n4223), .B(n4222), .Z(n1896) );
  COND3X1 U2524 ( .A(n7792), .B(n1895), .C(n4221), .D(n1896), .Z(n1897) );
  CND2IXL U2525 ( .B(n4224), .A(n4225), .Z(n1898) );
  CENX1 U2526 ( .A(n1897), .B(n1898), .Z(n1899) );
  CMX2XL U2527 ( .A0(out1_2[11]), .A1(n1899), .S(cmd1_en_2), .Z(n7924) );
  CIVXL U2528 ( .A(n4379), .Z(n1900) );
  CANR2XL U2529 ( .A(n4363), .B(out1_2[3]), .C(acc[3]), .D(n4350), .Z(n1901)
         );
  CEOX1 U2530 ( .A(n3198), .B(n2944), .Z(n1902) );
  CND2X1 U2531 ( .A(n4344), .B(n1902), .Z(n1903) );
  CIVX2 U2532 ( .A(n7746), .Z(n1904) );
  COND2XL U2533 ( .A(n4254), .B(n7581), .C(n3175), .D(n1904), .Z(n1905) );
  COND1XL U2534 ( .A(n3148), .B(n7745), .C(n8019), .Z(n1906) );
  CANR3XL U2535 ( .A(n4251), .B(n7743), .C(n1905), .D(n1906), .Z(n1907) );
  COND1XL U2536 ( .A(n4266), .B(n7688), .C(n1907), .Z(n1908) );
  COND2XL U2537 ( .A(n3091), .B(n7727), .C(n4267), .D(n7689), .Z(n1909) );
  COND2XL U2538 ( .A(n2865), .B(n2891), .C(n1908), .D(n1909), .Z(n2892) );
  CND2XL U2539 ( .A(n6380), .B(n6379), .Z(n1910) );
  CND2XL U2540 ( .A(n1910), .B(n6378), .Z(n1911) );
  CND2XL U2541 ( .A(n3743), .B(n6377), .Z(n1912) );
  CENX1 U2542 ( .A(n1911), .B(n1912), .Z(N31) );
  CND2XL U2543 ( .A(n6890), .B(n6888), .Z(n1913) );
  CENX1 U2544 ( .A(n6889), .B(n1914), .Z(n6882) );
  COND2X1 U2545 ( .A(n7228), .B(n6553), .C(n2382), .D(n6645), .Z(n1915) );
  COND2X1 U2546 ( .A(n2433), .B(n6650), .C(n2282), .D(n6462), .Z(n1916) );
  CENX1 U2547 ( .A(n6620), .B(n1915), .Z(n1917) );
  CENX1 U2548 ( .A(n1916), .B(n1917), .Z(n6623) );
  CANR5CX1 U2549 ( .A(n6620), .B(n1915), .C(n1916), .Z(n1918) );
  CIVX2 U2550 ( .A(n1918), .Z(n6671) );
  COND2XL U2551 ( .A(n4959), .B(n3579), .C(n4957), .D(n3565), .Z(n1919) );
  COND2XL U2552 ( .A(n5695), .B(n3585), .C(n4886), .D(n3564), .Z(n1920) );
  CANR5CXL U2553 ( .A(n3607), .B(n1919), .C(n1920), .Z(n1921) );
  CIVX1 U2554 ( .A(n1921), .Z(n3591) );
  CENX1 U2555 ( .A(n3607), .B(n1919), .Z(n1922) );
  CENX2 U2556 ( .A(n1920), .B(n1922), .Z(n3625) );
  CND2XL U2557 ( .A(acc[43]), .B(n2758), .Z(n1923) );
  CANR2XL U2558 ( .A(n2737), .B(out1_2[43]), .C(n2928), .D(out0_2[43]), .Z(
        n1924) );
  CND2X1 U2559 ( .A(n1923), .B(n1924), .Z(n2987) );
  CANR5CX1 U2560 ( .A(n1976), .B(n1975), .C(n6401), .Z(n1925) );
  CIVX2 U2561 ( .A(n1925), .Z(n6499) );
  CANR5CX1 U2562 ( .A(n3685), .B(n3684), .C(n3683), .Z(n1926) );
  CIVX2 U2563 ( .A(n1926), .Z(n3712) );
  CANR5CXL U2564 ( .A(n3678), .B(n3677), .C(n3676), .Z(n1927) );
  CIVXL U2565 ( .A(n1927), .Z(n3715) );
  CIVX1 U2566 ( .A(n3694), .Z(n1928) );
  CANR1X2 U2567 ( .A(n3696), .B(n3695), .C(n1928), .Z(n4360) );
  CND2IX1 U2568 ( .B(n3231), .A(n3232), .Z(n4328) );
  CND2IX1 U2569 ( .B(n3294), .A(n3295), .Z(n4280) );
  CND2XL U2570 ( .A(n7755), .B(n3122), .Z(n1929) );
  CANR2X1 U2571 ( .A(n3136), .B(n7582), .C(n3118), .D(n2859), .Z(n1930) );
  CND2X1 U2572 ( .A(n1929), .B(n1930), .Z(n7689) );
  CANR2X1 U2573 ( .A(n3181), .B(n7582), .C(n7755), .D(n3182), .Z(n1931) );
  CANR2X1 U2574 ( .A(n3160), .B(n7747), .C(n2859), .D(n3159), .Z(n1932) );
  CND2X1 U2575 ( .A(n1931), .B(n1932), .Z(n3134) );
  CNR2XL U2576 ( .A(n3145), .B(n7763), .Z(n1933) );
  COND2XL U2577 ( .A(n3143), .B(n7770), .C(n7766), .D(n3144), .Z(n1934) );
  CANR3X1 U2578 ( .A(n3174), .B(n2995), .C(n1933), .D(n1934), .Z(n4252) );
  CANR2X1 U2579 ( .A(n4363), .B(out1_2[60]), .C(acc[60]), .D(n8004), .Z(n1935)
         );
  CNR2X1 U2580 ( .A(n4318), .B(n7945), .Z(n1936) );
  CENX1 U2581 ( .A(n7942), .B(n1936), .Z(n1937) );
  CND2X1 U2582 ( .A(n4344), .B(n1937), .Z(n1938) );
  COND3X1 U2583 ( .A(n2685), .B(n7943), .C(n1935), .D(n1938), .Z(n1053) );
  CNR2IXL U2584 ( .B(n4132), .A(n4131), .Z(n1939) );
  CNR2XL U2585 ( .A(n7818), .B(n4134), .Z(n1940) );
  COND1XL U2586 ( .A(n4134), .B(n7830), .C(n4133), .Z(n1941) );
  CANR1XL U2587 ( .A(n3949), .B(n1940), .C(n1941), .Z(n1942) );
  CENX1 U2588 ( .A(n1939), .B(n1942), .Z(n1943) );
  CMX2XL U2589 ( .A0(out1_2[49]), .A1(n1943), .S(n7846), .Z(n7886) );
  CND2X1 U2590 ( .A(n4239), .B(n7788), .Z(n1944) );
  CND2XL U2591 ( .A(n1944), .B(n4238), .Z(n1945) );
  CND2IXL U2592 ( .B(n4236), .A(n4237), .Z(n1946) );
  CENX1 U2593 ( .A(n1945), .B(n1946), .Z(n1947) );
  CMX2XL U2594 ( .A0(out1_2[5]), .A1(n1947), .S(n8022), .Z(n7930) );
  CND2XL U2595 ( .A(n6375), .B(n6379), .Z(n1948) );
  COND3X1 U2596 ( .A(n6376), .B(n6378), .C(n6377), .D(n1948), .Z(n1949) );
  CND2XL U2597 ( .A(n6373), .B(n6374), .Z(n1950) );
  CENX1 U2598 ( .A(n1949), .B(n1950), .Z(N32) );
  COND1XL U2599 ( .A(n3148), .B(n3113), .C(n8019), .Z(n1951) );
  COND2XL U2600 ( .A(n7557), .B(n3189), .C(n4254), .D(n3114), .Z(n1952) );
  CANR3XL U2601 ( .A(n3115), .B(n4257), .C(n1951), .D(n1952), .Z(n1953) );
  COND1XL U2602 ( .A(n7727), .B(n3116), .C(n1953), .Z(n1954) );
  COND2X1 U2603 ( .A(n4266), .B(n7693), .C(n4267), .D(n7692), .Z(n1955) );
  COND2XL U2604 ( .A(n2865), .B(n3219), .C(n1954), .D(n1955), .Z(n3117) );
  CANR5CXL U2605 ( .A(n6434), .B(n6435), .C(n6436), .Z(n1956) );
  CIVX1 U2606 ( .A(n1956), .Z(n6596) );
  COND2X1 U2607 ( .A(n6293), .B(n3349), .C(n6418), .D(n3386), .Z(n1957) );
  COND2X1 U2608 ( .A(n6703), .B(n3388), .C(n2514), .D(n3356), .Z(n1958) );
  CENX1 U2609 ( .A(n3359), .B(n1957), .Z(n1959) );
  CENX1 U2610 ( .A(n1958), .B(n1959), .Z(n3433) );
  CANR5CXL U2611 ( .A(n3359), .B(n1957), .C(n1958), .Z(n1960) );
  CIVX1 U2612 ( .A(n1960), .Z(n3782) );
  CANR5CX1 U2613 ( .A(n2049), .B(n2048), .C(n6539), .Z(n1961) );
  CIVX2 U2614 ( .A(n1961), .Z(n6624) );
  COND2X1 U2615 ( .A(n6969), .B(n6968), .C(n7171), .D(n7053), .Z(n1962) );
  COND2X1 U2616 ( .A(n2293), .B(n6971), .C(n7114), .D(n7066), .Z(n1963) );
  CANR5CX1 U2617 ( .A(n7059), .B(n1962), .C(n1963), .Z(n1964) );
  CIVX1 U2618 ( .A(n1964), .Z(n7086) );
  CANR5CXL U2619 ( .A(n2086), .B(n2088), .C(n4563), .Z(n1965) );
  CIVX1 U2620 ( .A(n1965), .Z(n4610) );
  CND2X1 U2621 ( .A(n6880), .B(n6881), .Z(n1966) );
  CND2X2 U2622 ( .A(n6885), .B(n6886), .Z(n1967) );
  CENX2 U2623 ( .A(n1966), .B(n1967), .Z(n1968) );
  CENX2 U2624 ( .A(n6990), .B(n1968), .Z(n6991) );
  CANR5CXL U2625 ( .A(n6990), .B(n1966), .C(n1967), .Z(n1969) );
  CIVX1 U2626 ( .A(n1969), .Z(n7074) );
  CIVX1 U2627 ( .A(n1970), .Z(n3596) );
  CND2X1 U2628 ( .A(acc[38]), .B(n2671), .Z(n1971) );
  CANR2XL U2629 ( .A(n2737), .B(out1_2[38]), .C(n2928), .D(out0_2[38]), .Z(
        n1972) );
  CND2X1 U2630 ( .A(n1971), .B(n1972), .Z(n3018) );
  CND2X1 U2631 ( .A(acc[45]), .B(n2758), .Z(n1973) );
  CANR2XL U2632 ( .A(n2737), .B(out1_2[45]), .C(n2928), .D(out0_2[45]), .Z(
        n1974) );
  CND2X1 U2633 ( .A(n1973), .B(n1974), .Z(n2996) );
  COND2X1 U2634 ( .A(n6701), .B(n6300), .C(n6765), .D(n6410), .Z(n1975) );
  COND2X1 U2635 ( .A(n6974), .B(n6302), .C(n6972), .D(n6416), .Z(n1976) );
  CENX1 U2636 ( .A(n6401), .B(n1976), .Z(n1977) );
  CENX1 U2637 ( .A(n1975), .B(n1977), .Z(n6393) );
  CIVXL U2638 ( .A(n3702), .Z(n1978) );
  CNR2XL U2639 ( .A(n3702), .B(n3692), .Z(n1979) );
  COND2X1 U2640 ( .A(n3705), .B(n1979), .C(n3703), .D(n1978), .Z(n3708) );
  CENXL U2641 ( .A(n3663), .B(n3662), .Z(n1980) );
  CENX1 U2642 ( .A(n3664), .B(n1980), .Z(n1981) );
  CENX1 U2643 ( .A(n3666), .B(n3667), .Z(n1982) );
  CENX1 U2644 ( .A(n1981), .B(n1982), .Z(n3716) );
  CANR5CXL U2645 ( .A(n3666), .B(n3667), .C(n1981), .Z(n1983) );
  CIVXL U2646 ( .A(n1983), .Z(n3717) );
  CANR5CX1 U2647 ( .A(n3638), .B(n3636), .C(n3637), .Z(n1984) );
  CIVX2 U2648 ( .A(n1984), .Z(n3723) );
  CANR2X1 U2649 ( .A(n3019), .B(n2995), .C(n3169), .D(n2988), .Z(n1985) );
  CANR2X1 U2650 ( .A(n2990), .B(n3173), .C(n3172), .D(n2989), .Z(n1986) );
  CND2X1 U2651 ( .A(n1985), .B(n1986), .Z(n4261) );
  CND2IX1 U2652 ( .B(n3300), .A(n3326), .Z(n4317) );
  CAOR2XL U2653 ( .A(n7582), .B(n3122), .C(n7755), .D(n3118), .Z(n7725) );
  CIVXL U2654 ( .A(n3338), .Z(n1987) );
  CANR2XL U2655 ( .A(n4363), .B(out1_2[8]), .C(n1429), .D(n4350), .Z(n1988) );
  CND2X1 U2656 ( .A(n3339), .B(out2_2[7]), .Z(n1989) );
  CENX1 U2657 ( .A(out2_2[8]), .B(n1989), .Z(n1990) );
  CND2X1 U2658 ( .A(n4344), .B(n1990), .Z(n1991) );
  COND3XL U2659 ( .A(n2685), .B(n1987), .C(n1988), .D(n1991), .Z(n1001) );
  CANR2X1 U2660 ( .A(n4363), .B(n4362), .C(acc[0]), .D(n4350), .Z(n1992) );
  COND3X1 U2661 ( .A(out2_2[0]), .B(roundit), .C(n4344), .D(n4364), .Z(n1993)
         );
  COND3XL U2662 ( .A(n2684), .B(n2685), .C(n1992), .D(n1993), .Z(n993) );
  CND2XL U2663 ( .A(n3085), .B(n7738), .Z(n1994) );
  CND2XL U2664 ( .A(out2_2[43]), .B(n7751), .Z(n1995) );
  COND3X1 U2665 ( .A(n7684), .B(n7742), .C(n1994), .D(n1995), .Z(n872) );
  CANR2XL U2666 ( .A(n4363), .B(out1_2[32]), .C(acc[32]), .D(n4350), .Z(n1996)
         );
  CND2X1 U2667 ( .A(n4353), .B(out2_2[31]), .Z(n1997) );
  CEOX1 U2668 ( .A(n7992), .B(n1997), .Z(n1998) );
  CND2X1 U2669 ( .A(n4344), .B(n1998), .Z(n1999) );
  CNR2IXL U2670 ( .B(n4021), .A(n4020), .Z(n2000) );
  CNR2IXL U2671 ( .B(n4078), .A(n4072), .Z(n2001) );
  CND2XL U2672 ( .A(n4075), .B(n2001), .Z(n2002) );
  CIVXL U2673 ( .A(n4076), .Z(n2003) );
  COND1XL U2674 ( .A(n4072), .B(n2003), .C(n4073), .Z(n2004) );
  CANR1XL U2675 ( .A(n2001), .B(n4077), .C(n2004), .Z(n2005) );
  COND1XL U2676 ( .A(n7659), .B(n2002), .C(n2005), .Z(n2006) );
  CNR2XL U2677 ( .A(n2002), .B(n7656), .Z(n2007) );
  CANR1XL U2678 ( .A(n3949), .B(n2007), .C(n2006), .Z(n2008) );
  CENX1 U2679 ( .A(n2000), .B(n2008), .Z(n2009) );
  CMX2XL U2680 ( .A0(out1_2[47]), .A1(n2009), .S(n7846), .Z(n7888) );
  CIVXL U2681 ( .A(n7792), .Z(n2010) );
  CANR1XL U2682 ( .A(n4220), .B(n2010), .C(n4222), .Z(n2011) );
  CND2XL U2683 ( .A(n4223), .B(n4221), .Z(n2012) );
  CEOXL U2684 ( .A(n2011), .B(n2012), .Z(n2013) );
  CMX2XL U2685 ( .A0(out1_2[10]), .A1(n2013), .S(n8022), .Z(n7925) );
  CIVXL U2686 ( .A(n4377), .Z(n2014) );
  CANR2XL U2687 ( .A(n4363), .B(out1_2[5]), .C(acc[5]), .D(n4350), .Z(n2015)
         );
  CENX1 U2688 ( .A(n2732), .B(n2891), .Z(n2016) );
  CND2X1 U2689 ( .A(n2016), .B(n4344), .Z(n2017) );
  CND2XL U2690 ( .A(n6384), .B(n6383), .Z(n2018) );
  CEOXL U2691 ( .A(n2432), .B(n2018), .Z(N33) );
  COND2XL U2692 ( .A(n7727), .B(n3133), .C(n3134), .D(n4266), .Z(n2019) );
  CANR1XL U2693 ( .A(n3168), .B(n4249), .C(n2019), .Z(n2020) );
  COND2XL U2694 ( .A(n3162), .B(n4254), .C(n3163), .D(n3175), .Z(n2021) );
  CANR3X1 U2695 ( .A(n4272), .B(n7683), .C(h0_1[6]), .D(n2021), .Z(n2022) );
  COND3XL U2696 ( .A(n7759), .B(n3189), .C(n2020), .D(n2022), .Z(n2023) );
  COND1XL U2697 ( .A(n2865), .B(n3320), .C(n2023), .Z(n3135) );
  CENXL U2698 ( .A(n6314), .B(n6312), .Z(n2024) );
  CENX1 U2699 ( .A(n6313), .B(n2024), .Z(n6346) );
  CANR5CX1 U2700 ( .A(n3613), .B(n3611), .C(n3612), .Z(n2656) );
  CNR2IX2 U2701 ( .B(n4517), .A(n4516), .Z(n2025) );
  COND2XL U2702 ( .A(n2489), .B(n4519), .C(n2571), .D(n4518), .Z(n2026) );
  CANR5CXL U2703 ( .A(n4557), .B(n2025), .C(n2026), .Z(n2027) );
  CIVX1 U2704 ( .A(n2027), .Z(n4556) );
  CND2X1 U2705 ( .A(n6607), .B(n6606), .Z(n2028) );
  CND2X2 U2706 ( .A(n2395), .B(n2028), .Z(n2029) );
  CENX2 U2707 ( .A(n6604), .B(n2029), .Z(n6919) );
  CENXL U2708 ( .A(n2091), .B(n2089), .Z(n2030) );
  CENX1 U2709 ( .A(n2090), .B(n2030), .Z(n3685) );
  CENX1 U2710 ( .A(n3426), .B(n3425), .Z(n2031) );
  CND2XL U2711 ( .A(n3595), .B(n3592), .Z(n2032) );
  CND2X1 U2712 ( .A(n2032), .B(n3519), .Z(n2033) );
  CENX1 U2713 ( .A(n3559), .B(n3560), .Z(n2034) );
  CENX1 U2714 ( .A(n2033), .B(n2034), .Z(n3601) );
  CND2X1 U2715 ( .A(n5244), .B(n5243), .Z(n2035) );
  CND2X2 U2716 ( .A(n2338), .B(n2035), .Z(n2036) );
  CENX2 U2717 ( .A(n5245), .B(n2036), .Z(n5290) );
  CND2X1 U2718 ( .A(acc[46]), .B(n2758), .Z(n2037) );
  CANR2XL U2719 ( .A(n2737), .B(out1_2[46]), .C(n2928), .D(out0_2[46]), .Z(
        n2038) );
  CND2X1 U2720 ( .A(n2037), .B(n2038), .Z(n2993) );
  CND2X1 U2721 ( .A(acc[55]), .B(n2758), .Z(n2039) );
  CANR2XL U2722 ( .A(n2737), .B(out1_2[55]), .C(n2928), .D(out0_2[55]), .Z(
        n2040) );
  CND2X1 U2723 ( .A(n2039), .B(n2040), .Z(n2982) );
  CENX1 U2724 ( .A(n7075), .B(n7076), .Z(n2041) );
  CENX1 U2725 ( .A(n7074), .B(n2041), .Z(n7000) );
  CENX1 U2726 ( .A(n3657), .B(n3656), .Z(n2042) );
  CENX1 U2727 ( .A(n3658), .B(n2042), .Z(n3718) );
  CANR2XL U2728 ( .A(n2983), .B(n3173), .C(n3169), .D(n2970), .Z(n2043) );
  CANR2XL U2729 ( .A(n3172), .B(n2981), .C(n2995), .D(n2967), .Z(n2044) );
  CND2X1 U2730 ( .A(n2043), .B(n2044), .Z(n3040) );
  CIVX1 U2731 ( .A(n4276), .Z(n2045) );
  CANR1X2 U2732 ( .A(n4278), .B(n4277), .C(n2045), .Z(n7524) );
  CANR2XL U2733 ( .A(n2995), .B(n3099), .C(n3097), .D(n3172), .Z(n2046) );
  CANR2XL U2734 ( .A(n3104), .B(n3173), .C(n3100), .D(n3169), .Z(n2047) );
  CND2X1 U2735 ( .A(n2046), .B(n2047), .Z(n7581) );
  COND2X1 U2736 ( .A(n7205), .B(n6497), .C(n7203), .D(n6461), .Z(n2048) );
  COND2X1 U2737 ( .A(n1582), .B(n6479), .C(n6765), .D(n6487), .Z(n2049) );
  CENX1 U2738 ( .A(n6539), .B(n2049), .Z(n2050) );
  CENX1 U2739 ( .A(n2048), .B(n2050), .Z(n6552) );
  CENX1 U2740 ( .A(n2173), .B(n4745), .Z(n2051) );
  CENX1 U2741 ( .A(n2172), .B(n2051), .Z(n4914) );
  CANR2X1 U2742 ( .A(out1_2[62]), .B(n4363), .C(n4344), .D(n3267), .Z(n2052)
         );
  CND2X1 U2743 ( .A(n8004), .B(acc[62]), .Z(n2053) );
  COND3X1 U2744 ( .A(n2685), .B(n7938), .C(n2052), .D(n2053), .Z(n1055) );
  CNR2IXL U2745 ( .B(n4031), .A(n4030), .Z(n2054) );
  CND2XL U2746 ( .A(n4033), .B(n4075), .Z(n2055) );
  CNR2XL U2747 ( .A(n2055), .B(n7656), .Z(n2056) );
  CND2XL U2748 ( .A(n4033), .B(n4077), .Z(n2057) );
  COND3XL U2749 ( .A(n7659), .B(n2055), .C(n4032), .D(n2057), .Z(n2058) );
  CANR1XL U2750 ( .A(n3949), .B(n2056), .C(n2058), .Z(n2059) );
  CENX1 U2751 ( .A(n2054), .B(n2059), .Z(n2060) );
  CMX2XL U2752 ( .A0(out1_2[45]), .A1(n2060), .S(n7846), .Z(n7890) );
  CNR2IXL U2753 ( .B(n4025), .A(n4024), .Z(n2061) );
  CNR2XL U2754 ( .A(n4039), .B(n4037), .Z(n2062) );
  COND1XL U2755 ( .A(n4037), .B(n4040), .C(n4038), .Z(n2063) );
  CANR1XL U2756 ( .A(n3949), .B(n2062), .C(n2063), .Z(n2064) );
  CENX1 U2757 ( .A(n2061), .B(n2064), .Z(n2065) );
  CMX2XL U2758 ( .A0(out1_2[39]), .A1(n2065), .S(n7846), .Z(n7896) );
  CNR2IXL U2759 ( .B(n4166), .A(n4165), .Z(n2066) );
  CNR2XL U2760 ( .A(n7635), .B(n7566), .Z(n2067) );
  COND1XL U2761 ( .A(n7566), .B(n7638), .C(n7567), .Z(n2068) );
  CANR1XL U2762 ( .A(n7806), .B(n2067), .C(n2068), .Z(n2069) );
  CENX1 U2763 ( .A(n2066), .B(n2069), .Z(n2070) );
  CMX2XL U2764 ( .A0(out1_2[25]), .A1(n2070), .S(n7846), .Z(n7910) );
  CIVXL U2765 ( .A(n1373), .Z(n2071) );
  CANR2XL U2766 ( .A(n4363), .B(out1_2[26]), .C(acc[26]), .D(n4350), .Z(n2072)
         );
  CNR2X1 U2767 ( .A(n4317), .B(n7997), .Z(n2073) );
  CEOX1 U2768 ( .A(n2073), .B(out2_2[26]), .Z(n2074) );
  CND2X1 U2769 ( .A(n4344), .B(n2074), .Z(n2075) );
  COND3X1 U2770 ( .A(n2685), .B(n2071), .C(n2072), .D(n2075), .Z(n1019) );
  COND1XL U2771 ( .A(n7790), .B(n7792), .C(n7791), .Z(n2076) );
  CND2IXL U2772 ( .B(n4208), .A(n4209), .Z(n2077) );
  CENX1 U2773 ( .A(n2076), .B(n2077), .Z(n2078) );
  CMX2XL U2774 ( .A0(out1_2[9]), .A1(n2078), .S(n8022), .Z(n7926) );
  CIVXL U2775 ( .A(n4380), .Z(n2079) );
  CANR2XL U2776 ( .A(n4363), .B(out1_2[15]), .C(acc[15]), .D(n4350), .Z(n2080)
         );
  CEOX1 U2777 ( .A(n8002), .B(n3321), .Z(n2081) );
  CND2X1 U2778 ( .A(n4344), .B(n2081), .Z(n2082) );
  COND1XL U2779 ( .A(n2432), .B(n4624), .C(n6384), .Z(n2083) );
  CND2XL U2780 ( .A(n4634), .B(n4635), .Z(n2084) );
  CENX1 U2781 ( .A(n2083), .B(n2084), .Z(N34) );
  CENX1 U2782 ( .A(n6021), .B(n6023), .Z(n2085) );
  CENX2 U2783 ( .A(n6005), .B(n2085), .Z(n6013) );
  CND2IXL U2784 ( .B(n5112), .A(n6525), .Z(n6577) );
  CND2X2 U2785 ( .A(n3763), .B(n3764), .Z(n2086) );
  CENX2 U2786 ( .A(n4563), .B(n2086), .Z(n2087) );
  CND2X1 U2787 ( .A(n3768), .B(n3769), .Z(n2088) );
  CENX2 U2788 ( .A(n2087), .B(n2088), .Z(n4618) );
  CNR2IX1 U2789 ( .B(n7539), .A(n4957), .Z(n2089) );
  COND2X1 U2790 ( .A(n7537), .B(n3675), .C(n5160), .D(n3686), .Z(n2090) );
  COND2XL U2791 ( .A(n5695), .B(n3689), .C(n4886), .D(n3673), .Z(n2091) );
  CANR5CXL U2792 ( .A(n2089), .B(n2090), .C(n2091), .Z(n2092) );
  CIVXL U2793 ( .A(n2092), .Z(n3676) );
  CENX1 U2794 ( .A(n3630), .B(n3629), .Z(n2093) );
  CENX1 U2795 ( .A(n3628), .B(n2093), .Z(n3638) );
  CENX1 U2796 ( .A(n3496), .B(n3495), .Z(n2094) );
  CENX1 U2797 ( .A(n3494), .B(n2094), .Z(n2095) );
  CENX1 U2798 ( .A(n3503), .B(n3504), .Z(n2096) );
  CENX1 U2799 ( .A(n2095), .B(n2096), .Z(n3597) );
  CANR5CX1 U2800 ( .A(n3503), .B(n3504), .C(n2095), .Z(n2097) );
  CIVX2 U2801 ( .A(n2097), .Z(n3527) );
  CENX2 U2802 ( .A(n5013), .B(n5014), .Z(n2098) );
  CND2X1 U2803 ( .A(acc[35]), .B(n2671), .Z(n2099) );
  CANR2XL U2804 ( .A(n2737), .B(out1_2[35]), .C(n2928), .D(out0_2[35]), .Z(
        n2100) );
  CND2X1 U2805 ( .A(n2099), .B(n2100), .Z(n3002) );
  CAN2XL U2806 ( .A(n7417), .B(n7422), .Z(n7344) );
  COND1X1 U2807 ( .A(n6398), .B(n6399), .C(n6397), .Z(n2101) );
  CND2X2 U2808 ( .A(n2101), .B(n6400), .Z(n6501) );
  CND2X2 U2809 ( .A(n7379), .B(n7385), .Z(n2102) );
  CNR2X2 U2810 ( .A(n7164), .B(n2102), .Z(n7131) );
  COND1XL U2811 ( .A(n5342), .B(n5344), .C(n2342), .Z(n2103) );
  CND2X1 U2812 ( .A(n2103), .B(n2444), .Z(n5329) );
  COND2X1 U2813 ( .A(n6969), .B(n5863), .C(n5989), .D(n7171), .Z(n5977) );
  COR2X1 U2814 ( .A(n3709), .B(n3708), .Z(n4277) );
  CIVXL U2815 ( .A(n3631), .Z(n2104) );
  COND1XL U2816 ( .A(n7539), .B(n2104), .C(n5160), .Z(n6370) );
  CND2IX1 U2817 ( .B(n4315), .A(n4316), .Z(n4319) );
  CND2IX1 U2818 ( .B(n2706), .A(n3279), .Z(n3237) );
  CND2IX1 U2819 ( .B(h0_1[0]), .A(h0_1[1]), .Z(n7770) );
  CENX1 U2820 ( .A(n4865), .B(n4864), .Z(n2105) );
  CENX1 U2821 ( .A(n4863), .B(n2105), .Z(n4917) );
  CANR2XL U2822 ( .A(out1_2[61]), .B(n4363), .C(n4344), .D(n2716), .Z(n2106)
         );
  CND2X1 U2823 ( .A(n8004), .B(acc[61]), .Z(n2107) );
  CND2XL U2824 ( .A(n7535), .B(n7534), .Z(n2108) );
  CENX1 U2825 ( .A(n7536), .B(n2108), .Z(N19) );
  CNR2IXL U2826 ( .B(n4035), .A(n4034), .Z(n2109) );
  CND2XL U2827 ( .A(n7654), .B(n7655), .Z(n2110) );
  CND2XL U2828 ( .A(n7654), .B(n7657), .Z(n2111) );
  COND3XL U2829 ( .A(n7659), .B(n2110), .C(n7653), .D(n2111), .Z(n2112) );
  CNR2XL U2830 ( .A(n2110), .B(n7656), .Z(n2113) );
  CANR1XL U2831 ( .A(n3949), .B(n2113), .C(n2112), .Z(n2114) );
  CENX1 U2832 ( .A(n2109), .B(n2114), .Z(n2115) );
  CMX2XL U2833 ( .A0(out1_2[43]), .A1(n2115), .S(n7846), .Z(n7892) );
  CIVX2 U2834 ( .A(n3949), .Z(n2116) );
  COND1XL U2835 ( .A(n4039), .B(n2116), .C(n4040), .Z(n2117) );
  CND2IXL U2836 ( .B(n4037), .A(n4038), .Z(n2118) );
  CENX1 U2837 ( .A(n2117), .B(n2118), .Z(n2119) );
  CMX2X1 U2838 ( .A0(out1_2[38]), .A1(n2119), .S(n7846), .Z(n7897) );
  CNR2IXL U2839 ( .B(n4005), .A(n4004), .Z(n2120) );
  CNR2XL U2840 ( .A(n4026), .B(n4041), .Z(n2121) );
  COND1XL U2841 ( .A(n4041), .B(n4027), .C(n4042), .Z(n2122) );
  CANR1XL U2842 ( .A(n3949), .B(n2121), .C(n2122), .Z(n2123) );
  CENX1 U2843 ( .A(n2120), .B(n2123), .Z(n2124) );
  CMX2XL U2844 ( .A0(out1_2[37]), .A1(n2124), .S(n7846), .Z(n7898) );
  CND2XL U2845 ( .A(n4192), .B(n3949), .Z(n2125) );
  CND2X1 U2846 ( .A(n2125), .B(n4191), .Z(n2126) );
  CND2IXL U2847 ( .B(n4107), .A(n4108), .Z(n2127) );
  CENX1 U2848 ( .A(n2126), .B(n2127), .Z(n2128) );
  CMX2XL U2849 ( .A0(out1_2[33]), .A1(n2128), .S(n7846), .Z(n7902) );
  CNR2IXL U2850 ( .B(n4164), .A(n4163), .Z(n2129) );
  CNR2XL U2851 ( .A(n4176), .B(n4173), .Z(n2130) );
  COND1XL U2852 ( .A(n4173), .B(n4177), .C(n4174), .Z(n2131) );
  CANR1XL U2853 ( .A(n7806), .B(n2130), .C(n2131), .Z(n2132) );
  CENX1 U2854 ( .A(n2129), .B(n2132), .Z(n2133) );
  CMX2XL U2855 ( .A0(out1_2[21]), .A1(n2133), .S(n7846), .Z(n7914) );
  CANR1XL U2856 ( .A(n4231), .B(n4226), .C(n4228), .Z(n2134) );
  CND2XL U2857 ( .A(n4226), .B(n4227), .Z(n2135) );
  COND1XL U2858 ( .A(n7792), .B(n2135), .C(n2134), .Z(n2136) );
  CND2IXL U2859 ( .B(n4230), .A(n4229), .Z(n2137) );
  CENX1 U2860 ( .A(n2136), .B(n2137), .Z(n2138) );
  CMX2XL U2861 ( .A0(out1_2[14]), .A1(n2138), .S(cmd1_en_2), .Z(n7921) );
  COND1XL U2862 ( .A(n7840), .B(n7839), .C(n7838), .Z(n2139) );
  CND2IXL U2863 ( .B(n7841), .A(n7842), .Z(n2140) );
  CENX1 U2864 ( .A(n2139), .B(n2140), .Z(n2141) );
  CMX2XL U2865 ( .A0(out1_2[3]), .A1(n2141), .S(n7846), .Z(n7931) );
  CNR2IXL U2866 ( .B(n7531), .A(n7533), .Z(n2142) );
  CENX1 U2867 ( .A(n7532), .B(n2142), .Z(N24) );
  CNR2IXL U2868 ( .B(n7504), .A(n7503), .Z(n2143) );
  CENX1 U2869 ( .A(n7505), .B(n2143), .Z(N28) );
  COND2XL U2870 ( .A(n7745), .B(n3189), .C(n3175), .D(n7581), .Z(n2144) );
  COND1XL U2871 ( .A(n4254), .B(n7580), .C(n8019), .Z(n2145) );
  CANR3XL U2872 ( .A(n4249), .B(n7746), .C(n2144), .D(n2145), .Z(n2146) );
  COND1XL U2873 ( .A(n4267), .B(n7725), .C(n2146), .Z(n2147) );
  COND2X1 U2874 ( .A(n7727), .B(n7730), .C(n4266), .D(n7728), .Z(n2148) );
  COND2XL U2875 ( .A(n2865), .B(n3333), .C(n2147), .D(n2148), .Z(n3142) );
  CIVX1 U2876 ( .A(n4378), .Z(n2149) );
  CANR2XL U2877 ( .A(n4350), .B(n1398), .C(n2947), .D(n4363), .Z(n2150) );
  CNR2X1 U2878 ( .A(n2944), .B(n3198), .Z(n2151) );
  CENX1 U2879 ( .A(n3187), .B(n2151), .Z(n2152) );
  CND2X1 U2880 ( .A(n4344), .B(n2152), .Z(n2153) );
  COND3XL U2881 ( .A(n2685), .B(n2149), .C(n2150), .D(n2153), .Z(n997) );
  CNR2IXL U2882 ( .B(n7844), .A(n7843), .Z(n2154) );
  CENX1 U2883 ( .A(n2154), .B(n7845), .Z(n2155) );
  CMX2X1 U2884 ( .A0(n7847), .A1(n2155), .S(n7846), .Z(n7933) );
  COND1X1 U2885 ( .A(n6357), .B(n6359), .C(n6358), .Z(n2156) );
  CND2X2 U2886 ( .A(n2156), .B(n2378), .Z(n6439) );
  CENX1 U2887 ( .A(n6392), .B(n6394), .Z(n2157) );
  CENX1 U2888 ( .A(n6393), .B(n2157), .Z(n6428) );
  CENX1 U2889 ( .A(n5737), .B(n5735), .Z(n2158) );
  CENX2 U2890 ( .A(n5595), .B(n2158), .Z(n5677) );
  CANR5CX1 U2891 ( .A(n6816), .B(n6817), .C(n6815), .Z(n2159) );
  CIVX2 U2892 ( .A(n2159), .Z(n6951) );
  CNR2XL U2893 ( .A(n2381), .B(n5906), .Z(n2160) );
  CNR2X1 U2894 ( .A(n5818), .B(n7228), .Z(n2161) );
  CNR2X2 U2895 ( .A(n2160), .B(n2161), .Z(n5918) );
  CND2XL U2896 ( .A(n6940), .B(n6941), .Z(n2162) );
  COND1X1 U2897 ( .A(n7327), .B(n2391), .C(n2162), .Z(n7438) );
  CANR2XL U2898 ( .A(n2969), .B(n3173), .C(n3172), .D(n2968), .Z(n2163) );
  CANR2XL U2899 ( .A(n2995), .B(n2993), .C(n3169), .D(n2997), .Z(n2164) );
  CND2X1 U2900 ( .A(n2163), .B(n2164), .Z(n3041) );
  CND2X1 U2901 ( .A(acc[27]), .B(n2671), .Z(n2165) );
  CANR2XL U2902 ( .A(n2737), .B(out1_2[27]), .C(n2928), .D(out0_2[27]), .Z(
        n2166) );
  CND2X1 U2903 ( .A(n2165), .B(n2166), .Z(n3014) );
  CENX2 U2904 ( .A(n5224), .B(n5223), .Z(n2167) );
  CENX2 U2905 ( .A(n5226), .B(n2167), .Z(n5270) );
  CND2IX1 U2906 ( .B(n4293), .A(n4298), .Z(n4343) );
  CANR2XL U2907 ( .A(n4262), .B(n7582), .C(n7755), .D(n4263), .Z(n2168) );
  CANR2XL U2908 ( .A(n2859), .B(n3066), .C(n7747), .D(n3065), .Z(n2169) );
  CND2XL U2909 ( .A(n2168), .B(n2169), .Z(n7699) );
  CANR2XL U2910 ( .A(n3160), .B(n7755), .C(n3161), .D(n2859), .Z(n2170) );
  CND2XL U2911 ( .A(n7582), .B(n3159), .Z(n2171) );
  CND2X1 U2912 ( .A(n2171), .B(n2170), .Z(n7712) );
  COND2X1 U2913 ( .A(n7537), .B(n4735), .C(n5160), .D(n4710), .Z(n2172) );
  COND2X1 U2914 ( .A(n1556), .B(n4740), .C(n6576), .D(n4708), .Z(n2173) );
  CANR5CX1 U2915 ( .A(n4745), .B(n2173), .C(n2172), .Z(n2174) );
  CIVX2 U2916 ( .A(n2174), .Z(n4896) );
  CENX2 U2917 ( .A(n7871), .B(n6411), .Z(n2175) );
  CND2X4 U2918 ( .A(n2175), .B(n1547), .Z(n6969) );
  CAN2X2 U2919 ( .A(n4968), .B(n4969), .Z(n4921) );
  CENX1 U2920 ( .A(q0[5]), .B(n7852), .Z(n2176) );
  CENX1 U2921 ( .A(q0[4]), .B(q0[3]), .Z(n2177) );
  CND2X4 U2922 ( .A(n2176), .B(n2177), .Z(n5911) );
  COND1X1 U2923 ( .A(n5874), .B(n5873), .C(n5875), .Z(n2178) );
  CND2X2 U2924 ( .A(n2178), .B(n5876), .Z(n5946) );
  COND2X1 U2925 ( .A(n2433), .B(n6496), .C(n2282), .D(n6420), .Z(n2179) );
  COND2X1 U2926 ( .A(n6523), .B(n6521), .C(n6419), .D(n6418), .Z(n2180) );
  CENXL U2927 ( .A(n6513), .B(n2179), .Z(n2181) );
  CENX1 U2928 ( .A(n2180), .B(n2181), .Z(n6534) );
  CANR5CXL U2929 ( .A(n6513), .B(n2179), .C(n2180), .Z(n2182) );
  CIVX1 U2930 ( .A(n2182), .Z(n6540) );
  CANR2XL U2931 ( .A(n4363), .B(out1_2[45]), .C(acc[45]), .D(n4350), .Z(n2183)
         );
  COND1XL U2932 ( .A(n2685), .B(n2629), .C(n2183), .Z(n2184) );
  CEOX1 U2933 ( .A(n7970), .B(n3237), .Z(n2185) );
  CANR1XL U2934 ( .A(n4344), .B(n2185), .C(n2184), .Z(n7850) );
  CIVXL U2935 ( .A(out0_2[58]), .Z(n2186) );
  CANR2XL U2936 ( .A(n4363), .B(out1_2[58]), .C(acc[58]), .D(n4350), .Z(n2187)
         );
  CNR2X1 U2937 ( .A(n3258), .B(n7949), .Z(n2188) );
  CENX1 U2938 ( .A(n7947), .B(n2188), .Z(n2189) );
  CND2X1 U2939 ( .A(n4344), .B(n2189), .Z(n2190) );
  COND3X1 U2940 ( .A(n2685), .B(n2186), .C(n2187), .D(n2190), .Z(n1051) );
  CIVXL U2941 ( .A(out0_2[54]), .Z(n2191) );
  CANR2XL U2942 ( .A(n4363), .B(out1_2[54]), .C(acc[54]), .D(n4350), .Z(n2192)
         );
  CNR2X1 U2943 ( .A(n3290), .B(n7957), .Z(n2193) );
  CENX1 U2944 ( .A(n7955), .B(n2193), .Z(n2194) );
  CND2X1 U2945 ( .A(n4344), .B(n2194), .Z(n2195) );
  CND2XL U2946 ( .A(n4277), .B(n4276), .Z(n2196) );
  CENX1 U2947 ( .A(n4278), .B(n2196), .Z(N20) );
  CIVX1 U2948 ( .A(n2965), .Z(n2197) );
  CANR2XL U2949 ( .A(n4363), .B(out1_2[33]), .C(acc[33]), .D(n4350), .Z(n2198)
         );
  CEOX1 U2950 ( .A(n7990), .B(n4286), .Z(n2199) );
  CND2X1 U2951 ( .A(n4344), .B(n2199), .Z(n2200) );
  COND3X1 U2952 ( .A(n2685), .B(n2197), .C(n2198), .D(n2200), .Z(n1026) );
  CNR2IXL U2953 ( .B(n4359), .A(n4358), .Z(n2201) );
  CENX1 U2954 ( .A(n4360), .B(n2201), .Z(N18) );
  CNR2IXL U2955 ( .B(n4046), .A(n4045), .Z(n2202) );
  COND1XL U2956 ( .A(n7645), .B(n7659), .C(n7646), .Z(n2203) );
  CNR2XL U2957 ( .A(n7656), .B(n7645), .Z(n2204) );
  CANR1XL U2958 ( .A(n3949), .B(n2204), .C(n2203), .Z(n2205) );
  CENX1 U2959 ( .A(n2202), .B(n2205), .Z(n2206) );
  CMX2XL U2960 ( .A0(out1_2[41]), .A1(n2206), .S(n7846), .Z(n7894) );
  CNR2IXL U2961 ( .B(n4042), .A(n4041), .Z(n2207) );
  CANR1XL U2962 ( .A(n4044), .B(n3949), .C(n4043), .Z(n2208) );
  CENX1 U2963 ( .A(n2207), .B(n2208), .Z(n2209) );
  CMX2XL U2964 ( .A0(out1_2[36]), .A1(n2209), .S(n7846), .Z(n7899) );
  CNR2IXL U2965 ( .B(n4007), .A(n4006), .Z(n2210) );
  CIVXL U2966 ( .A(n7666), .Z(n2211) );
  CIVXL U2967 ( .A(n7669), .Z(n2212) );
  COND1XL U2968 ( .A(n7666), .B(n2212), .C(n7667), .Z(n2213) );
  CANR11X1 U2969 ( .A(n3949), .B(n7670), .C(n2211), .D(n2213), .Z(n2214) );
  CENX1 U2970 ( .A(n2210), .B(n2214), .Z(n2215) );
  CMX2XL U2971 ( .A0(out1_2[35]), .A1(n2215), .S(n7846), .Z(n7900) );
  CND2XL U2972 ( .A(n4212), .B(n7806), .Z(n2216) );
  CND2X1 U2973 ( .A(n2216), .B(n4211), .Z(n2217) );
  CND2IXL U2974 ( .B(n4160), .A(n4161), .Z(n2218) );
  CENX1 U2975 ( .A(n2217), .B(n2218), .Z(n2219) );
  CMX2XL U2976 ( .A0(out1_2[17]), .A1(n2219), .S(n7846), .Z(n7918) );
  CANR2XL U2977 ( .A(n4363), .B(out1_2[30]), .C(acc[30]), .D(n4350), .Z(n2220)
         );
  CNR2X1 U2978 ( .A(n4319), .B(n7995), .Z(n2221) );
  CEOX1 U2979 ( .A(n2221), .B(out2_2[30]), .Z(n2222) );
  CND2X1 U2980 ( .A(n4344), .B(n2222), .Z(n2223) );
  COND3X1 U2981 ( .A(n2685), .B(n2647), .C(n2220), .D(n2223), .Z(n1023) );
  CNR2IXL U2982 ( .B(n7791), .A(n7790), .Z(n2224) );
  CENX1 U2983 ( .A(n2224), .B(n7792), .Z(n2225) );
  CMX2XL U2984 ( .A0(out1_2[8]), .A1(n2225), .S(n8022), .Z(n7927) );
  CIVXL U2985 ( .A(n4376), .Z(n2226) );
  CANR2XL U2986 ( .A(n4363), .B(out1_2[6]), .C(acc[6]), .D(n4350), .Z(n2227)
         );
  CND2X1 U2987 ( .A(n2732), .B(out2_2[5]), .Z(n2228) );
  CENX1 U2988 ( .A(out2_2[6]), .B(n2228), .Z(n2229) );
  CND2X1 U2989 ( .A(n4344), .B(n2229), .Z(n2230) );
  CIVXL U2990 ( .A(n4375), .Z(n2231) );
  CANR2XL U2991 ( .A(n4363), .B(out1_2[7]), .C(acc[7]), .D(n4350), .Z(n2232)
         );
  CENX1 U2992 ( .A(n3339), .B(n4270), .Z(n2233) );
  CND2X1 U2993 ( .A(n2233), .B(n4344), .Z(n2234) );
  CIVXL U2994 ( .A(n4382), .Z(n2235) );
  CANR2XL U2995 ( .A(n4363), .B(out1_2[13]), .C(acc[13]), .D(n4350), .Z(n2236)
         );
  CEOX1 U2996 ( .A(n8003), .B(n3218), .Z(n2237) );
  CND2X1 U2997 ( .A(n4344), .B(n2237), .Z(n2238) );
  CANR2XL U2998 ( .A(n4363), .B(out1_2[18]), .C(acc[18]), .D(n4350), .Z(n2239)
         );
  CND2X1 U2999 ( .A(n3322), .B(out2_2[17]), .Z(n2240) );
  CENX1 U3000 ( .A(out2_2[18]), .B(n2240), .Z(n2241) );
  CND2X1 U3001 ( .A(n4344), .B(n2241), .Z(n2242) );
  CIVXL U3002 ( .A(n1387), .Z(n2243) );
  CANR2XL U3003 ( .A(n4363), .B(out1_2[22]), .C(acc[22]), .D(n4350), .Z(n2244)
         );
  CNR2X1 U3004 ( .A(n4280), .B(n4279), .Z(n2245) );
  CEOX1 U3005 ( .A(n2245), .B(out2_2[22]), .Z(n2246) );
  CND2X1 U3006 ( .A(n4344), .B(n2246), .Z(n2247) );
  COND3X1 U3007 ( .A(n2685), .B(n2243), .C(n2244), .D(n2247), .Z(n1015) );
  COND1XL U3008 ( .A(n7533), .B(n7532), .C(n7531), .Z(n2248) );
  CND2IXL U3009 ( .B(n7529), .A(n7530), .Z(n2249) );
  CENX1 U3010 ( .A(n2248), .B(n2249), .Z(N25) );
  CND2XL U3011 ( .A(n6389), .B(n4087), .Z(n2250) );
  CENX1 U3012 ( .A(n6388), .B(n2250), .Z(N26) );
  COND1XL U3013 ( .A(n7503), .B(n7505), .C(n7504), .Z(n2251) );
  CND2IXL U3014 ( .B(n7501), .A(n7502), .Z(n2252) );
  CENX1 U3015 ( .A(n2251), .B(n2252), .Z(N29) );
  COND1XL U3016 ( .A(n7526), .B(n2432), .C(n7525), .Z(n2253) );
  CND2IXL U3017 ( .B(n7527), .A(n7528), .Z(n2254) );
  CENX1 U3018 ( .A(n2253), .B(n2254), .Z(N35) );
  CND2XL U3019 ( .A(n4656), .B(n4655), .Z(n2255) );
  CIVX1 U3020 ( .A(n3284), .Z(n2256) );
  CANR2XL U3021 ( .A(n4363), .B(out1_2[24]), .C(n1425), .D(n4350), .Z(n2257)
         );
  CND2X1 U3022 ( .A(n3326), .B(out2_2[23]), .Z(n2258) );
  CENX1 U3023 ( .A(out2_2[24]), .B(n2258), .Z(n2259) );
  CND2X1 U3024 ( .A(n4344), .B(n2259), .Z(n2260) );
  COND3XL U3025 ( .A(n2685), .B(n2256), .C(n2257), .D(n2260), .Z(n1017) );
  CND2XL U3026 ( .A(n4239), .B(n4238), .Z(n2261) );
  CENX1 U3027 ( .A(n7788), .B(n2261), .Z(n2262) );
  CMX2X1 U3028 ( .A0(n2947), .A1(n2262), .S(n7846), .Z(n1116) );
  CNR2IXL U3029 ( .B(n7838), .A(n7840), .Z(n2263) );
  CENX1 U3030 ( .A(n2263), .B(n7839), .Z(n2264) );
  CIVXL U3031 ( .A(n4362), .Z(n2265) );
  COND1XL U3032 ( .A(n2964), .B(out1_1[0]), .C(n7845), .Z(n2266) );
  CMXI2X1 U3033 ( .A0(n2265), .A1(n2266), .S(n7846), .Z(n7934) );
  CENX1 U3034 ( .A(n6028), .B(n6027), .Z(n2267) );
  CENX1 U3035 ( .A(n6026), .B(n2267), .Z(n6012) );
  CND2IX1 U3036 ( .B(n5803), .A(n5804), .Z(n6055) );
  COND2X1 U3037 ( .A(n6701), .B(n6644), .C(n6700), .D(n6765), .Z(n6698) );
  CENX1 U3038 ( .A(n5211), .B(n2448), .Z(n2268) );
  CND2X1 U3039 ( .A(n2268), .B(n5267), .Z(n5227) );
  CEOX1 U3040 ( .A(n5559), .B(n5560), .Z(n2593) );
  CENX1 U3041 ( .A(n6251), .B(n6253), .Z(n2269) );
  CENX1 U3042 ( .A(n6250), .B(n2269), .Z(n6259) );
  CENX1 U3043 ( .A(n5682), .B(n5684), .Z(n2270) );
  CENX1 U3044 ( .A(n2343), .B(n2270), .Z(n5679) );
  CAOR1X1 U3045 ( .A(n2569), .B(n2491), .C(n6292), .Z(n6447) );
  CENX1 U3046 ( .A(n6427), .B(n6426), .Z(n2271) );
  CENX1 U3047 ( .A(n6428), .B(n2271), .Z(n6454) );
  CENX1 U3048 ( .A(n6839), .B(n6838), .Z(n2272) );
  CENX1 U3049 ( .A(n6781), .B(n2272), .Z(n6856) );
  COND2X1 U3050 ( .A(n7228), .B(n5039), .C(n2382), .D(n5700), .Z(n2273) );
  CENX1 U3051 ( .A(n5618), .B(n2273), .Z(n5637) );
  CANR2X1 U3052 ( .A(n7808), .B(out0_2[11]), .C(out1_2[11]), .D(n3902), .Z(
        n2274) );
  COND1XL U3053 ( .A(n8018), .B(n7810), .C(n2274), .Z(n3908) );
  CENX1 U3054 ( .A(n3677), .B(n3676), .Z(n2275) );
  CENX1 U3055 ( .A(n3678), .B(n2275), .Z(n3713) );
  COND2X1 U3056 ( .A(n2294), .B(n6470), .C(n7114), .D(n6471), .Z(n2403) );
  CND2X1 U3057 ( .A(n6803), .B(n6804), .Z(n6806) );
  CND2IX1 U3058 ( .B(n3247), .A(n3248), .Z(n3286) );
  CND4X1 U3059 ( .A(n7450), .B(n7132), .C(n7373), .D(n7131), .Z(n7169) );
  CIVX1 U3060 ( .A(n7384), .Z(n2276) );
  CANR1XL U3061 ( .A(n7375), .B(n7385), .C(n2276), .Z(n7376) );
  CAN3X1 U3062 ( .A(n5949), .B(n5948), .C(n5947), .Z(n5951) );
  COAN1X1 U3063 ( .A(n6371), .B(n6370), .C(n6372), .Z(N16) );
  CIVXL U3064 ( .A(n6706), .Z(n2277) );
  CNIVXL U3065 ( .A(h0[21]), .Z(n2278) );
  CNIVX4 U3066 ( .A(h0[21]), .Z(n2279) );
  CNIVX4 U3067 ( .A(h0[21]), .Z(n2280) );
  CENX1 U3068 ( .A(n5734), .B(n5733), .Z(n2281) );
  CNIVX1 U3069 ( .A(n5806), .Z(n5734) );
  CND2X2 U3070 ( .A(n4676), .B(n2555), .Z(n2282) );
  CND2X2 U3071 ( .A(n4676), .B(n2555), .Z(n7126) );
  COND2X1 U3072 ( .A(n2564), .B(n5765), .C(n2487), .D(n5796), .Z(n5844) );
  CENX1 U3073 ( .A(n6417), .B(h0[23]), .Z(n5708) );
  CANR1XL U3074 ( .A(n4641), .B(n4640), .C(n1576), .Z(n2284) );
  CENXL U3075 ( .A(n5203), .B(n5202), .Z(n2285) );
  CENX1 U3076 ( .A(n5203), .B(n5202), .Z(n5204) );
  CNIVX4 U3077 ( .A(n6969), .Z(n6774) );
  CENX1 U3078 ( .A(n6678), .B(n6679), .Z(n6643) );
  COND1X1 U3079 ( .A(n3729), .B(n4086), .C(n3728), .Z(n7500) );
  CND2X2 U3080 ( .A(n6368), .B(n6367), .Z(n7454) );
  CEO3X2 U3081 ( .A(n6454), .B(n6453), .C(n6455), .Z(n6368) );
  CND2X1 U3082 ( .A(n6565), .B(n6564), .Z(n6485) );
  CENX1 U3083 ( .A(n6565), .B(n6564), .Z(n6566) );
  CEO3X2 U3084 ( .A(n6288), .B(n6286), .C(n6289), .Z(n2286) );
  CND2X1 U3085 ( .A(n5645), .B(n5647), .Z(n2289) );
  CND2X2 U3086 ( .A(n2287), .B(n2288), .Z(n2290) );
  CND2X2 U3087 ( .A(n2289), .B(n2290), .Z(n5042) );
  CIVX2 U3088 ( .A(n5645), .Z(n2287) );
  CIVX2 U3089 ( .A(n5647), .Z(n2288) );
  CENXL U3090 ( .A(n5648), .B(n5042), .Z(n2291) );
  CENXL U3091 ( .A(n5648), .B(n5042), .Z(n2292) );
  CNIVX4 U3092 ( .A(n7113), .Z(n2293) );
  CNIVX4 U3093 ( .A(n7113), .Z(n2294) );
  CNIVX4 U3094 ( .A(n7113), .Z(n2295) );
  CENXL U3095 ( .A(n5648), .B(n5042), .Z(n2398) );
  CND2X2 U3096 ( .A(n4535), .B(n2374), .Z(n7113) );
  CND2X1 U3097 ( .A(n5165), .B(n5164), .Z(n2493) );
  CAN2X1 U3098 ( .A(n6291), .B(n6290), .Z(n2296) );
  CENX1 U3099 ( .A(n5257), .B(n5256), .Z(n5258) );
  CNR2XL U3100 ( .A(n5256), .B(n5257), .Z(n5221) );
  CND2XL U3101 ( .A(n5256), .B(n5257), .Z(n5220) );
  CNIVX4 U3102 ( .A(n5711), .Z(n6702) );
  CND2XL U3103 ( .A(n5737), .B(n5736), .Z(n5738) );
  CENX1 U3104 ( .A(h0[11]), .B(n6828), .Z(n4765) );
  CENX1 U3105 ( .A(n6460), .B(h0[11]), .Z(n5989) );
  CENXL U3106 ( .A(n5932), .B(h0[25]), .Z(n6676) );
  CNIVX1 U3107 ( .A(n7012), .Z(n2297) );
  CND2X1 U3108 ( .A(n6291), .B(n6290), .Z(n6367) );
  CEOX1 U3109 ( .A(n3478), .B(n3477), .Z(n3558) );
  CIVX2 U3110 ( .A(n2298), .Z(n3483) );
  CND2X1 U3111 ( .A(n3478), .B(n3477), .Z(n2298) );
  CENX1 U3112 ( .A(n3548), .B(n3547), .Z(n3741) );
  COND2X2 U3113 ( .A(n6770), .B(n4951), .C(n5097), .D(n6870), .Z(n5150) );
  COND1X1 U3114 ( .A(n5061), .B(n5060), .C(n5059), .Z(n5062) );
  CIVX2 U3115 ( .A(n6790), .Z(n2299) );
  CND2X1 U3116 ( .A(n4628), .B(n4626), .Z(n4622) );
  COND1X1 U3117 ( .A(n4626), .B(n4628), .C(n4625), .Z(n4623) );
  CNIVX1 U3118 ( .A(n5749), .Z(n5750) );
  CENX2 U3119 ( .A(n5288), .B(n5287), .Z(n5289) );
  CND2X1 U3120 ( .A(n4792), .B(n4791), .Z(n4793) );
  CENX1 U3121 ( .A(n5473), .B(n5472), .Z(n5492) );
  CND2XL U3122 ( .A(n5314), .B(n5313), .Z(n5315) );
  CENXL U3123 ( .A(n5312), .B(n5313), .Z(n4478) );
  CND2X2 U3124 ( .A(n2301), .B(n2302), .Z(n2303) );
  CIVX2 U3125 ( .A(n6903), .Z(n2301) );
  CIVX2 U3126 ( .A(n6902), .Z(n2302) );
  CNIVX1 U3127 ( .A(n6882), .Z(n2304) );
  CND2X1 U3128 ( .A(n2305), .B(n2306), .Z(n2307) );
  CIVXL U3129 ( .A(n6890), .Z(n2305) );
  CIVXL U3130 ( .A(n6888), .Z(n2306) );
  CND2X2 U3131 ( .A(n2552), .B(n2553), .Z(n2308) );
  CND2X1 U3132 ( .A(n6032), .B(n6033), .Z(n2311) );
  CND2X2 U3133 ( .A(n2309), .B(n2310), .Z(n2312) );
  CND2X2 U3134 ( .A(n2311), .B(n2312), .Z(n6037) );
  CIVX2 U3135 ( .A(n6032), .Z(n2309) );
  CIVX2 U3136 ( .A(n6033), .Z(n2310) );
  CND2X1 U3137 ( .A(n5094), .B(n5092), .Z(n4971) );
  CND2IXL U3138 ( .B(n7860), .A(q0[16]), .Z(n2600) );
  COND2X1 U3139 ( .A(n7252), .B(n7172), .C(n7253), .D(n7207), .Z(n7194) );
  CND2X1 U3140 ( .A(n4783), .B(n4782), .Z(n4784) );
  COND2XL U3141 ( .A(n7252), .B(n7223), .C(n7253), .D(n7251), .Z(n7250) );
  CAOR1XL U3142 ( .A(n7253), .B(n7252), .C(n7251), .Z(n7277) );
  COND2XL U3143 ( .A(n7252), .B(n7219), .C(n7253), .D(n7223), .Z(n7224) );
  COND2XL U3144 ( .A(n7252), .B(n7207), .C(n7253), .D(n7219), .Z(n7220) );
  CND2X1 U3145 ( .A(n7098), .B(n7097), .Z(n7099) );
  CENX1 U3146 ( .A(n7070), .B(n7098), .Z(n7102) );
  CIVXL U3147 ( .A(n6382), .Z(n7494) );
  CND2X1 U3148 ( .A(n3802), .B(n3801), .Z(n3803) );
  COND2X1 U3149 ( .A(n6765), .B(n3789), .C(n3401), .D(n1582), .Z(n3760) );
  CIVXL U3150 ( .A(n7489), .Z(n2313) );
  CIVXL U3151 ( .A(n2313), .Z(n2314) );
  CND2X1 U3152 ( .A(n5932), .B(n2512), .Z(n2317) );
  CND2X2 U3153 ( .A(n2315), .B(n2316), .Z(n2318) );
  CND2X2 U3154 ( .A(n2317), .B(n2318), .Z(n5219) );
  CIVX2 U3155 ( .A(n2512), .Z(n2316) );
  CND2XL U3156 ( .A(n4863), .B(n4864), .Z(n2319) );
  CND2X1 U3157 ( .A(n4863), .B(n4865), .Z(n2320) );
  CND2XL U3158 ( .A(n4864), .B(n4865), .Z(n2321) );
  CND3X1 U3159 ( .A(n2319), .B(n2320), .C(n2321), .Z(n4825) );
  COND1X1 U3160 ( .A(n4916), .B(n4917), .C(n4915), .Z(n4871) );
  CND2X4 U3161 ( .A(n7439), .B(n7443), .Z(n7337) );
  CND2XL U3162 ( .A(n6357), .B(n6359), .Z(n2378) );
  CND2X1 U3163 ( .A(n6348), .B(n6347), .Z(n6349) );
  CENXL U3164 ( .A(n7173), .B(h0[25]), .Z(n7174) );
  CENX2 U3165 ( .A(n6011), .B(n6013), .Z(n6006) );
  COND1X1 U3166 ( .A(n4825), .B(n4828), .C(n4826), .Z(n4693) );
  CND2X1 U3167 ( .A(n4828), .B(n4825), .Z(n4692) );
  COND1X1 U3168 ( .A(n5087), .B(n5090), .C(n5088), .Z(n4841) );
  CND2X1 U3169 ( .A(n5087), .B(n5090), .Z(n4840) );
  CEOX1 U3170 ( .A(n3463), .B(h0[1]), .Z(n3460) );
  CND2X1 U3171 ( .A(n6941), .B(n6940), .Z(n2322) );
  CND2X1 U3172 ( .A(n6941), .B(n6940), .Z(n7326) );
  CND2X1 U3173 ( .A(n5375), .B(n5374), .Z(n5376) );
  COND1X2 U3174 ( .A(n5374), .B(n5375), .C(n5373), .Z(n5377) );
  CEO3X2 U3175 ( .A(n7073), .B(n7072), .C(n7071), .Z(n7075) );
  CND2X1 U3176 ( .A(n7073), .B(n7071), .Z(n2324) );
  CND3X2 U3177 ( .A(n2323), .B(n2324), .C(n2325), .Z(n7101) );
  CND2XL U3178 ( .A(n7076), .B(n7074), .Z(n2326) );
  CND2X1 U3179 ( .A(n7076), .B(n7075), .Z(n2327) );
  CND2X1 U3180 ( .A(n7074), .B(n7075), .Z(n2328) );
  CND3X1 U3181 ( .A(n2326), .B(n2327), .C(n2328), .Z(n7153) );
  CNIVX2 U3182 ( .A(n7323), .Z(n7379) );
  CND2XL U3183 ( .A(n5812), .B(n2333), .Z(n2331) );
  CND2X1 U3184 ( .A(n2329), .B(n2330), .Z(n2332) );
  CND2X2 U3185 ( .A(n2331), .B(n2332), .Z(n5703) );
  CIVXL U3186 ( .A(n5812), .Z(n2329) );
  CIVXL U3187 ( .A(n5811), .Z(n2330) );
  COND2XL U3188 ( .A(n5911), .B(n5702), .C(n5912), .D(n5794), .Z(n2333) );
  COND2XL U3189 ( .A(n5911), .B(n5702), .C(n5912), .D(n5794), .Z(n2334) );
  COND2XL U3190 ( .A(n5911), .B(n5702), .C(n5912), .D(n5794), .Z(n5811) );
  CNR2X1 U3191 ( .A(n5520), .B(n5519), .Z(n2335) );
  CND2X2 U3192 ( .A(n2336), .B(n2337), .Z(n2338) );
  CIVX2 U3193 ( .A(n5244), .Z(n2336) );
  CIVX2 U3194 ( .A(n5243), .Z(n2337) );
  CNR2X1 U3195 ( .A(n5520), .B(n5519), .Z(n5553) );
  CND2X1 U3196 ( .A(n5286), .B(n5285), .Z(n5519) );
  CENX1 U3197 ( .A(n5843), .B(n5844), .Z(n5766) );
  CIVX2 U3198 ( .A(n5161), .Z(n5303) );
  CENX1 U3199 ( .A(n5932), .B(h0[7]), .Z(n4860) );
  CND2X1 U3200 ( .A(n4707), .B(n4706), .Z(n4909) );
  CND2X1 U3201 ( .A(n5961), .B(n5963), .Z(n5903) );
  CND2IX2 U3202 ( .B(n6418), .A(n5101), .Z(n5102) );
  CENX2 U3203 ( .A(n6232), .B(n6101), .Z(n6253) );
  CNIVX2 U3204 ( .A(n5464), .Z(n5507) );
  CENX1 U3205 ( .A(n5335), .B(n5334), .Z(n2339) );
  CIVX2 U3206 ( .A(q0[12]), .Z(n2340) );
  CIVX2 U3207 ( .A(n2340), .Z(n2341) );
  COND2XL U3208 ( .A(n2569), .B(n5193), .C(n2489), .D(n5192), .Z(n2342) );
  CANR1X1 U3209 ( .A(n7411), .B(n7406), .C(n7294), .Z(n7295) );
  COND1X1 U3210 ( .A(n7291), .B(n7290), .C(n2625), .Z(n7406) );
  CENX2 U3211 ( .A(n5389), .B(n5242), .Z(n5520) );
  CENX2 U3212 ( .A(n5373), .B(n5374), .Z(n5137) );
  CENX1 U3213 ( .A(h0[7]), .B(n6970), .Z(n4773) );
  CNIVX1 U3214 ( .A(n5683), .Z(n2343) );
  COND2X1 U3215 ( .A(n2565), .B(n3372), .C(n2488), .D(n3786), .Z(n3770) );
  CIVX2 U3216 ( .A(n4975), .Z(n2344) );
  CIVX3 U3217 ( .A(n2344), .Z(n2345) );
  CENX1 U3218 ( .A(n4815), .B(n4814), .Z(n4816) );
  COND1X1 U3219 ( .A(n4815), .B(n4817), .C(n4814), .Z(n4777) );
  CIVX8 U3220 ( .A(n2598), .Z(n6409) );
  CND2X1 U3221 ( .A(n2440), .B(n5848), .Z(n5851) );
  CANR11X2 U3222 ( .A(n3744), .B(n6374), .C(n3743), .D(n3742), .Z(n2346) );
  CANR11XL U3223 ( .A(n3744), .B(n6374), .C(n3743), .D(n3742), .Z(n3745) );
  COND1XL U3224 ( .A(n6023), .B(n6022), .C(n6021), .Z(n6025) );
  CND2XL U3225 ( .A(n6023), .B(n6022), .Z(n6024) );
  COND2X1 U3226 ( .A(n2294), .B(n6002), .C(n7114), .D(n6001), .Z(n6023) );
  CNR2X4 U3227 ( .A(n7028), .B(n2366), .Z(n6283) );
  CIVX12 U3228 ( .A(n7866), .Z(n5932) );
  CAOR1X1 U3229 ( .A(n2477), .B(n7065), .C(n7064), .Z(n7080) );
  CENX2 U3230 ( .A(n5439), .B(n5438), .Z(n5441) );
  CND2X2 U3231 ( .A(n5576), .B(n5575), .Z(n2348) );
  CND2X1 U3232 ( .A(n5576), .B(n5575), .Z(n2349) );
  CND2XL U3233 ( .A(n5576), .B(n5575), .Z(n5730) );
  CIVX2 U3234 ( .A(n5573), .Z(n5576) );
  CIVXL U3235 ( .A(n7313), .Z(n2350) );
  CIVXL U3236 ( .A(n2350), .Z(n2351) );
  CANR1X1 U3237 ( .A(n7353), .B(n7358), .C(n7155), .Z(n2352) );
  CEOX2 U3238 ( .A(n4433), .B(n4431), .Z(n2353) );
  CEOX2 U3239 ( .A(n2353), .B(n1238), .Z(n4550) );
  CND2XL U3240 ( .A(n4432), .B(n4431), .Z(n2354) );
  CND2X1 U3241 ( .A(n4432), .B(n4433), .Z(n2355) );
  CND2XL U3242 ( .A(n4431), .B(n4433), .Z(n2356) );
  COND1X1 U3243 ( .A(n4578), .B(n4581), .C(n4579), .Z(n4573) );
  CND2X1 U3244 ( .A(n5320), .B(n5174), .Z(n5175) );
  CNIVX1 U3245 ( .A(n6032), .Z(n6034) );
  CNIVX1 U3246 ( .A(n6591), .Z(n2357) );
  CENX1 U3247 ( .A(n5977), .B(n5976), .Z(n5865) );
  COND1X1 U3248 ( .A(n6893), .B(n6894), .C(n6892), .Z(n6896) );
  CIVX2 U3249 ( .A(n6169), .Z(n2503) );
  CENX1 U3250 ( .A(n6417), .B(h0[25]), .Z(n5985) );
  CIVX2 U3251 ( .A(n2611), .Z(n2358) );
  CANR1X1 U3252 ( .A(n2525), .B(n6928), .C(n2482), .Z(n2359) );
  CANR1X1 U3253 ( .A(n2525), .B(n6928), .C(n2482), .Z(n2623) );
  CEOX1 U3254 ( .A(h0[17]), .B(n2484), .Z(n4859) );
  CIVXL U3255 ( .A(n7319), .Z(n2360) );
  CND2IX2 U3256 ( .B(n7425), .A(n2361), .Z(n7275) );
  CNR2X2 U3257 ( .A(n7236), .B(n2360), .Z(n2361) );
  CENX1 U3258 ( .A(n2454), .B(h0[16]), .Z(n5866) );
  CNIVX1 U3259 ( .A(n5956), .Z(n2362) );
  CNIVX1 U3260 ( .A(n5331), .Z(n2363) );
  COND2XL U3261 ( .A(n2563), .B(n5192), .C(n2489), .D(n5111), .Z(n2364) );
  COND2XL U3262 ( .A(n2563), .B(n5192), .C(n2491), .D(n5111), .Z(n2365) );
  COND2X1 U3263 ( .A(n2563), .B(n5192), .C(n2491), .D(n5111), .Z(n5188) );
  CND2IX2 U3264 ( .B(n6703), .A(n5710), .Z(n5715) );
  CENXL U3265 ( .A(n5932), .B(h0[24]), .Z(n6640) );
  CENXL U3266 ( .A(n5932), .B(n7539), .Z(n4398) );
  CENXL U3267 ( .A(n5932), .B(h0[23]), .Z(n6584) );
  CENXL U3268 ( .A(n5932), .B(h0[18]), .Z(n6184) );
  CENXL U3269 ( .A(n5932), .B(h0[26]), .Z(n6746) );
  CENXL U3270 ( .A(n5932), .B(h0[22]), .Z(n6489) );
  CENXL U3271 ( .A(n5932), .B(n2279), .Z(n6481) );
  CENXL U3272 ( .A(n5932), .B(h0[27]), .Z(n6793) );
  CENXL U3273 ( .A(n5932), .B(h0[19]), .Z(n6302) );
  CENX1 U3274 ( .A(n5932), .B(h0[30]), .Z(n6973) );
  CENXL U3275 ( .A(n5932), .B(h0[20]), .Z(n6416) );
  CENXL U3276 ( .A(h0[31]), .B(n1583), .Z(n7064) );
  CNR2X2 U3277 ( .A(n6281), .B(n6280), .Z(n2366) );
  CANR1X1 U3278 ( .A(n7472), .B(n6270), .C(n6269), .Z(n2367) );
  CANR1X1 U3279 ( .A(n7472), .B(n6270), .C(n6269), .Z(n2368) );
  CENX2 U3280 ( .A(q0[10]), .B(q0[9]), .Z(n2369) );
  CANR1X1 U3281 ( .A(n7472), .B(n6270), .C(n6269), .Z(n7004) );
  CENX2 U3282 ( .A(q0[10]), .B(q0[9]), .Z(n3578) );
  CEOX2 U3283 ( .A(n6550), .B(n6552), .Z(n2370) );
  CEOX2 U3284 ( .A(n2370), .B(n6551), .Z(n6587) );
  CND2XL U3285 ( .A(n6551), .B(n6552), .Z(n2371) );
  CND2X1 U3286 ( .A(n6551), .B(n6550), .Z(n2372) );
  CND2XL U3287 ( .A(n6552), .B(n6550), .Z(n2373) );
  CENX1 U3288 ( .A(q0[22]), .B(q0[21]), .Z(n2374) );
  CND2XL U3289 ( .A(n6633), .B(n6632), .Z(n6634) );
  CENX1 U3290 ( .A(q0[21]), .B(q0[22]), .Z(n5168) );
  CANR1X1 U3291 ( .A(n7344), .B(n7343), .C(n7342), .Z(n7345) );
  COND2X1 U3292 ( .A(n5911), .B(n5181), .C(n5912), .D(n5095), .Z(n5255) );
  COND2X1 U3293 ( .A(n5911), .B(n4720), .C(n5912), .D(n4726), .Z(n4746) );
  CENX2 U3294 ( .A(n5270), .B(n5269), .Z(n2375) );
  CENXL U3295 ( .A(n5270), .B(n5269), .Z(n5403) );
  CND2X2 U3296 ( .A(n6925), .B(n6924), .Z(n2376) );
  CND2X1 U3297 ( .A(n4891), .B(n4890), .Z(n4892) );
  CND2IX1 U3298 ( .B(n5569), .A(n2412), .Z(n2414) );
  CND2X1 U3299 ( .A(n6778), .B(n6777), .Z(n6779) );
  CEOX1 U3300 ( .A(n7864), .B(h0[25]), .Z(n6100) );
  CEOX2 U3301 ( .A(n6359), .B(n6357), .Z(n2377) );
  CEOX2 U3302 ( .A(n2377), .B(n6358), .Z(n6347) );
  COR2X1 U3303 ( .A(n2294), .B(n6212), .Z(n2379) );
  CND2X2 U3304 ( .A(n6439), .B(n6438), .Z(n6440) );
  COND1X1 U3305 ( .A(n6348), .B(n6347), .C(n6346), .Z(n6350) );
  CND2XL U3306 ( .A(n6260), .B(n6259), .Z(n6261) );
  CNIVX4 U3307 ( .A(n4800), .Z(n2381) );
  CNIVX4 U3308 ( .A(n4800), .Z(n2382) );
  CNIVX2 U3309 ( .A(n4800), .Z(n7301) );
  CEO3X2 U3310 ( .A(n4912), .B(n4913), .C(n4914), .Z(n5138) );
  CND2XL U3311 ( .A(n4912), .B(n4914), .Z(n2383) );
  CND2X1 U3312 ( .A(n4912), .B(n4913), .Z(n2384) );
  CND2X1 U3313 ( .A(n4914), .B(n4913), .Z(n2385) );
  CND3X2 U3314 ( .A(n2383), .B(n2384), .C(n2385), .Z(n4976) );
  CND2X4 U3315 ( .A(n3643), .B(n3366), .Z(n3364) );
  CENX2 U3316 ( .A(n6103), .B(h0[1]), .Z(n4722) );
  COND1X1 U3317 ( .A(n5528), .B(n2399), .C(n5526), .Z(n2386) );
  COND1X1 U3318 ( .A(n5528), .B(n2399), .C(n5526), .Z(n6928) );
  CND2X1 U3319 ( .A(n6041), .B(n5982), .Z(n2389) );
  CND2X2 U3320 ( .A(n2387), .B(n2388), .Z(n2390) );
  CND2X2 U3321 ( .A(n2389), .B(n2390), .Z(n6007) );
  CIVX2 U3322 ( .A(n6041), .Z(n2387) );
  CIVX2 U3323 ( .A(n5982), .Z(n2388) );
  CND2X2 U3324 ( .A(n7374), .B(n7378), .Z(n6941) );
  CANR1X1 U3325 ( .A(n7457), .B(n6933), .C(n6932), .Z(n2391) );
  CANR1X1 U3326 ( .A(n7457), .B(n6933), .C(n6932), .Z(n2392) );
  CND2X2 U3327 ( .A(n2393), .B(n2394), .Z(n2395) );
  CIVX2 U3328 ( .A(n6607), .Z(n2393) );
  CIVX2 U3329 ( .A(n6606), .Z(n2394) );
  CANR1X1 U3330 ( .A(n7457), .B(n6933), .C(n6932), .Z(n7382) );
  COR2XL U3331 ( .A(n6114), .B(n4487), .Z(n4407) );
  CNIVX1 U3332 ( .A(n6969), .Z(n2396) );
  CNIVXL U3333 ( .A(n6969), .Z(n2397) );
  CNIVXL U3334 ( .A(n6969), .Z(n6307) );
  CNIVXL U3335 ( .A(n6969), .Z(n6468) );
  CNIVX1 U3336 ( .A(n6969), .Z(n7119) );
  COND1X1 U3337 ( .A(n6624), .B(n6623), .C(n6622), .Z(n6626) );
  CEOX2 U3338 ( .A(n2582), .B(h0[30]), .Z(n5924) );
  CENXL U3339 ( .A(n5648), .B(n5042), .Z(n5657) );
  CEO3X2 U3340 ( .A(n6983), .B(n6982), .C(n6984), .Z(n6994) );
  CND2X2 U3341 ( .A(n7407), .B(n7411), .Z(n7296) );
  COND2X2 U3342 ( .A(n7114), .B(n6772), .C(n6731), .D(n7095), .Z(n6803) );
  CANR1X1 U3343 ( .A(n5516), .B(n5515), .C(n5534), .Z(n2399) );
  CANR1X1 U3344 ( .A(n5516), .B(n5515), .C(n5534), .Z(n5527) );
  CND2X2 U3345 ( .A(n2602), .B(n2603), .Z(n2605) );
  COND1X1 U3346 ( .A(n6501), .B(n6500), .C(n6499), .Z(n6503) );
  COND1X2 U3347 ( .A(n5647), .B(n5648), .C(n5646), .Z(n5650) );
  CIVXL U3348 ( .A(n5583), .Z(n2400) );
  CIVXL U3349 ( .A(n2400), .Z(n2401) );
  CEO3X2 U3350 ( .A(n6501), .B(n6499), .C(n6500), .Z(n6606) );
  CND2X1 U3351 ( .A(n5561), .B(n5560), .Z(n5562) );
  CENX1 U3352 ( .A(n6460), .B(h0[18]), .Z(n6469) );
  COND1X1 U3353 ( .A(n7051), .B(n6963), .C(n6962), .Z(n2473) );
  COND1XL U3354 ( .A(n7051), .B(n7339), .C(n1562), .Z(n7149) );
  COND1X2 U3355 ( .A(n7236), .B(n7427), .C(n2661), .Z(n7313) );
  CEOX2 U3356 ( .A(n5677), .B(n5676), .Z(n2402) );
  CENX1 U3357 ( .A(n5677), .B(n5676), .Z(n5601) );
  CND2X1 U3358 ( .A(n6680), .B(n6679), .Z(n6681) );
  COND1X1 U3359 ( .A(n6679), .B(n6680), .C(n6678), .Z(n6682) );
  CND2X2 U3360 ( .A(n4682), .B(n4681), .Z(n5073) );
  CND2X2 U3361 ( .A(n2413), .B(n2414), .Z(n5682) );
  CENX1 U3362 ( .A(h0[10]), .B(n6828), .Z(n4718) );
  COND2X2 U3363 ( .A(n6701), .B(n4767), .C(n6765), .D(n5048), .Z(n5068) );
  COR2XL U3364 ( .A(n1557), .B(n6000), .Z(n5817) );
  CENX2 U3365 ( .A(n5701), .B(h0[26]), .Z(n4797) );
  COND1X2 U3366 ( .A(n6121), .B(n6122), .C(n6120), .Z(n6124) );
  COND1XL U3367 ( .A(n7476), .B(n7475), .C(n7474), .Z(n7477) );
  COND1XL U3368 ( .A(n7462), .B(n7475), .C(n7461), .Z(n7463) );
  COND1XL U3369 ( .A(n7475), .B(n7045), .C(n7044), .Z(n7050) );
  CANR1X1 U3370 ( .A(n6283), .B(n7038), .C(n6282), .Z(n2405) );
  CANR1X1 U3371 ( .A(n6283), .B(n7038), .C(n6282), .Z(n2406) );
  CANR1X1 U3372 ( .A(n6283), .B(n7038), .C(n6282), .Z(n6284) );
  CENXL U3373 ( .A(n6171), .B(n6220), .Z(n6275) );
  CENX2 U3374 ( .A(n4702), .B(n4703), .Z(n4704) );
  CND2X4 U3375 ( .A(n4667), .B(n4666), .Z(n4703) );
  CND2X1 U3376 ( .A(n5205), .B(n2285), .Z(n2410) );
  CND2X2 U3377 ( .A(n2409), .B(n2408), .Z(n2411) );
  CND2X2 U3378 ( .A(n2410), .B(n2411), .Z(n5292) );
  CIVX2 U3379 ( .A(n5205), .Z(n2408) );
  CIVX2 U3380 ( .A(n5204), .Z(n2409) );
  CNIVX1 U3381 ( .A(n5201), .Z(n5205) );
  CENX1 U3382 ( .A(n7134), .B(n7674), .Z(n4771) );
  CND2XL U3383 ( .A(n5568), .B(n5569), .Z(n2413) );
  CIVXL U3384 ( .A(n5568), .Z(n2412) );
  CENXL U3385 ( .A(n5741), .B(n5743), .Z(n5568) );
  CENX1 U3386 ( .A(n7134), .B(h0[26]), .Z(n6968) );
  COND1X2 U3387 ( .A(n4439), .B(n4441), .C(n4438), .Z(n4395) );
  CND2X1 U3388 ( .A(n5470), .B(n5469), .Z(n5430) );
  CNIVX1 U3389 ( .A(n5469), .Z(n5473) );
  CNIVX1 U3390 ( .A(n5246), .Z(n2415) );
  CND2X1 U3391 ( .A(n5365), .B(n5364), .Z(n2418) );
  CND2X2 U3392 ( .A(n2416), .B(n2417), .Z(n2419) );
  CND2X2 U3393 ( .A(n2418), .B(n2419), .Z(n5368) );
  CIVX2 U3394 ( .A(n5365), .Z(n2416) );
  CIVX2 U3395 ( .A(n5364), .Z(n2417) );
  CND2X2 U3396 ( .A(n3755), .B(n4421), .Z(n2420) );
  CND2X2 U3397 ( .A(n3755), .B(n4421), .Z(n6870) );
  CND2X1 U3398 ( .A(n7151), .B(n2438), .Z(n2421) );
  CIVXL U3399 ( .A(n1563), .Z(n2422) );
  CND2X2 U3400 ( .A(n2421), .B(n2422), .Z(n7314) );
  COND1X1 U3401 ( .A(n5180), .B(n5178), .C(n5177), .Z(n5123) );
  CENX1 U3402 ( .A(h0[25]), .B(n5104), .Z(n4846) );
  CND2X1 U3403 ( .A(n5485), .B(n5484), .Z(n5486) );
  COND1X1 U3404 ( .A(n5484), .B(n5485), .C(n5483), .Z(n5487) );
  CND2X1 U3405 ( .A(n6363), .B(n6214), .Z(n2425) );
  CND2X2 U3406 ( .A(n2423), .B(n2424), .Z(n2426) );
  CND2X2 U3407 ( .A(n2425), .B(n2426), .Z(n6288) );
  CIVXL U3408 ( .A(n6363), .Z(n2423) );
  CIVX2 U3409 ( .A(n6214), .Z(n2424) );
  CND2X1 U3410 ( .A(n6362), .B(n6360), .Z(n2429) );
  CND2X2 U3411 ( .A(n2427), .B(n2428), .Z(n2430) );
  CND2X2 U3412 ( .A(n2429), .B(n2430), .Z(n6214) );
  CIVX2 U3413 ( .A(n6362), .Z(n2427) );
  CIVX2 U3414 ( .A(n6360), .Z(n2428) );
  CNIVXL U3415 ( .A(n5462), .Z(n2455) );
  COND1X2 U3416 ( .A(n6883), .B(n6884), .C(n6882), .Z(n6886) );
  CNIVX1 U3417 ( .A(n5547), .Z(n2431) );
  COAN1XL U3418 ( .A(n3746), .B(n3808), .C(n3745), .Z(n2432) );
  CNIVX4 U3419 ( .A(n4675), .Z(n2433) );
  CNIVX2 U3420 ( .A(n4675), .Z(n7124) );
  CNIVX1 U3421 ( .A(n6857), .Z(n2434) );
  CNIVX2 U3422 ( .A(n7340), .Z(n7421) );
  CND2X1 U3423 ( .A(n4817), .B(n4815), .Z(n4776) );
  CIVXL U3424 ( .A(n4670), .Z(n2435) );
  CIVXL U3425 ( .A(n2435), .Z(n2436) );
  CNR2X2 U3426 ( .A(n7466), .B(n7465), .Z(n2446) );
  CEO3X2 U3427 ( .A(n6856), .B(n6855), .C(n2434), .Z(n6952) );
  CMX2XL U3428 ( .A0(n2280), .A1(h[21]), .S(n7682), .Z(n950) );
  CENX1 U3429 ( .A(n7134), .B(h0[2]), .Z(n4954) );
  CND2X1 U3430 ( .A(n6455), .B(n6454), .Z(n6456) );
  CNIVX2 U3431 ( .A(n5482), .Z(n2437) );
  CEO3X2 U3432 ( .A(n6893), .B(n6892), .C(n6894), .Z(n6954) );
  CND2X1 U3433 ( .A(n4581), .B(n4578), .Z(n4572) );
  CND2XL U3434 ( .A(n4508), .B(n4505), .Z(n4497) );
  CENXL U3435 ( .A(n4506), .B(n4505), .Z(n4507) );
  COND1X1 U3436 ( .A(n6942), .B(n2392), .C(n2322), .Z(n2438) );
  COND1X1 U3437 ( .A(n6942), .B(n7382), .C(n7326), .Z(n7150) );
  COND1X1 U3438 ( .A(n6438), .B(n6439), .C(n6437), .Z(n6441) );
  CND2X2 U3439 ( .A(n5715), .B(n5714), .Z(n2440) );
  CND2XL U3440 ( .A(n6065), .B(n6064), .Z(n2441) );
  CIVXL U3441 ( .A(h0[6]), .Z(n2442) );
  CEO3X2 U3442 ( .A(n5343), .B(n5344), .C(n5342), .Z(n5423) );
  CND2X1 U3443 ( .A(n5342), .B(n5344), .Z(n2444) );
  CND2X1 U3444 ( .A(n5476), .B(n5475), .Z(n5477) );
  CENXL U3445 ( .A(n6653), .B(n6493), .Z(n2445) );
  CENXL U3446 ( .A(n6653), .B(n6493), .Z(n6661) );
  CENX1 U3447 ( .A(n6652), .B(n6651), .Z(n6493) );
  CND2XL U3448 ( .A(n6158), .B(n6157), .Z(n6159) );
  COND1XL U3449 ( .A(n6157), .B(n6158), .C(n6156), .Z(n6160) );
  CND2X2 U3450 ( .A(n6768), .B(n6767), .Z(n6845) );
  CNR2X2 U3451 ( .A(n7466), .B(n7465), .Z(n6268) );
  CND2XL U3452 ( .A(n7497), .B(n1260), .Z(n7498) );
  CND2X1 U3453 ( .A(n4948), .B(n4947), .Z(n5231) );
  CND2X2 U3454 ( .A(n7469), .B(n6270), .Z(n7020) );
  CENX2 U3455 ( .A(h0[27]), .B(n2583), .Z(n5754) );
  COND1X2 U3456 ( .A(n6096), .B(n2396), .C(n6095), .Z(n6232) );
  CIVXL U3457 ( .A(n5793), .Z(n2447) );
  CND2IX1 U3458 ( .B(q0[16]), .A(n2599), .Z(n2601) );
  CNIVX1 U3459 ( .A(n5210), .Z(n2448) );
  CND2X4 U3460 ( .A(n3347), .B(n3346), .Z(n2449) );
  CND2IXL U3461 ( .B(n6663), .A(n6662), .Z(n6664) );
  COND1X1 U3462 ( .A(n5952), .B(n5951), .C(n5950), .Z(n2450) );
  COND1XL U3463 ( .A(n5952), .B(n5951), .C(n5950), .Z(n2451) );
  COND1X1 U3464 ( .A(n5332), .B(n5335), .C(n5333), .Z(n5266) );
  CNR2X2 U3465 ( .A(n5078), .B(n5077), .Z(n7310) );
  CIVXL U3466 ( .A(n5959), .Z(n2452) );
  CIVX2 U3467 ( .A(n2452), .Z(n2453) );
  CENX1 U3468 ( .A(n6061), .B(n5820), .Z(n5959) );
  CIVX2 U3469 ( .A(n1551), .Z(n2454) );
  CENX1 U3470 ( .A(n3569), .B(n3568), .Z(n3589) );
  CND2X1 U3471 ( .A(n3568), .B(n3567), .Z(n3479) );
  COND2X1 U3472 ( .A(n5580), .B(n6114), .C(n3368), .D(n5754), .Z(n5720) );
  CND2X1 U3473 ( .A(n3368), .B(n6114), .Z(n6117) );
  CND2X1 U3474 ( .A(n6761), .B(n6760), .Z(n6762) );
  COND1X1 U3475 ( .A(n6761), .B(n6760), .C(n6759), .Z(n6763) );
  CND2X1 U3476 ( .A(n4441), .B(n4439), .Z(n4394) );
  CND2XL U3477 ( .A(n5187), .B(n2364), .Z(n5120) );
  CENX1 U3478 ( .A(n6324), .B(n6326), .Z(n6195) );
  CIVXL U3479 ( .A(n6324), .Z(n6325) );
  CND2X1 U3480 ( .A(n6266), .B(n6265), .Z(n7307) );
  CNIVX2 U3481 ( .A(n5045), .Z(n4754) );
  CENX2 U3482 ( .A(n5044), .B(n5043), .Z(n4755) );
  CNIVX16 U3483 ( .A(n5168), .Z(n7114) );
  CND2X1 U3484 ( .A(n5956), .B(n5957), .Z(n2539) );
  CEOX1 U3485 ( .A(n2582), .B(h0[29]), .Z(n5910) );
  COND1X1 U3486 ( .A(n5480), .B(n5479), .C(n5482), .Z(n5457) );
  CND2X1 U3487 ( .A(n5479), .B(n5480), .Z(n5456) );
  CND2X1 U3488 ( .A(n6653), .B(n6652), .Z(n6654) );
  CIVX2 U3489 ( .A(n6187), .Z(n6444) );
  CND2X2 U3490 ( .A(n5522), .B(n5521), .Z(n5549) );
  CEOX1 U3491 ( .A(n7853), .B(h0[19]), .Z(n6795) );
  CND2X1 U3492 ( .A(n6884), .B(n6883), .Z(n6885) );
  CENX1 U3493 ( .A(n6647), .B(h0[10]), .Z(n5190) );
  CND2X2 U3494 ( .A(n6264), .B(n6263), .Z(n6280) );
  CIVX2 U3495 ( .A(n3759), .Z(n2456) );
  CENX1 U3496 ( .A(h0[28]), .B(n5104), .Z(n4887) );
  CND3XL U3497 ( .A(n7132), .B(n7131), .C(n7373), .Z(n7448) );
  CENX2 U3498 ( .A(n6531), .B(n6530), .Z(n6532) );
  CNR2X2 U3499 ( .A(n2308), .B(n6267), .Z(n7460) );
  CENX1 U3500 ( .A(h0[30]), .B(n2531), .Z(n5567) );
  CNIVX2 U3501 ( .A(n5140), .Z(n5141) );
  CND2X1 U3502 ( .A(n5140), .B(n5138), .Z(n4973) );
  CND2X1 U3503 ( .A(n6259), .B(n6130), .Z(n2459) );
  CIVXL U3504 ( .A(n6259), .Z(n2457) );
  CIVX2 U3505 ( .A(n6130), .Z(n2458) );
  CND2X1 U3506 ( .A(n6260), .B(n6258), .Z(n2462) );
  CND2X2 U3507 ( .A(n2460), .B(n2461), .Z(n2463) );
  CND2X2 U3508 ( .A(n2462), .B(n2463), .Z(n6130) );
  CIVX2 U3509 ( .A(n6258), .Z(n2460) );
  CIVX2 U3510 ( .A(n6260), .Z(n2461) );
  CNIVX4 U3511 ( .A(n6639), .Z(n2477) );
  CND2XL U3512 ( .A(n6314), .B(n6313), .Z(n6316) );
  COND1X1 U3513 ( .A(n6314), .B(n6313), .C(n6312), .Z(n6315) );
  COND1X1 U3514 ( .A(n6209), .B(n6969), .C(n6208), .Z(n6313) );
  CANR1X1 U3515 ( .A(n7271), .B(n7267), .C(n7241), .Z(n7242) );
  CEO3X2 U3516 ( .A(n4921), .B(n4920), .C(n4919), .Z(n5235) );
  CAOR1X1 U3517 ( .A(n6871), .B(n2420), .C(n6869), .Z(n6965) );
  CANR1X1 U3518 ( .A(n6929), .B(n2404), .C(n6927), .Z(n2467) );
  CANR1X1 U3519 ( .A(n6929), .B(n2404), .C(n6927), .Z(n7362) );
  CND2X1 U3520 ( .A(n5198), .B(n5325), .Z(n5199) );
  CND2X1 U3521 ( .A(n4631), .B(n4630), .Z(n4632) );
  COND1X1 U3522 ( .A(n4631), .B(n4630), .C(n4629), .Z(n4633) );
  CIVX3 U3523 ( .A(n4867), .Z(n7095) );
  COND2X1 U3524 ( .A(n6974), .B(n6481), .C(n6972), .D(n6489), .Z(n6518) );
  CND2X1 U3525 ( .A(n6857), .B(n6856), .Z(n6858) );
  CND2X2 U3526 ( .A(n5165), .B(n5164), .Z(n5321) );
  CENX1 U3527 ( .A(n7134), .B(h0[5]), .Z(n4772) );
  CND2X1 U3528 ( .A(n5368), .B(n5367), .Z(n2471) );
  CND2X2 U3529 ( .A(n2469), .B(n2470), .Z(n2472) );
  CND2X2 U3530 ( .A(n2471), .B(n2472), .Z(n5386) );
  CIVX2 U3531 ( .A(n5368), .Z(n2469) );
  CIVX2 U3532 ( .A(n5367), .Z(n2470) );
  CNR2X2 U3533 ( .A(n7020), .B(n6285), .Z(n2525) );
  CENX1 U3534 ( .A(n6491), .B(h0[10]), .Z(n4477) );
  COND2X2 U3535 ( .A(n2449), .B(n4389), .C(n1586), .D(n4477), .Z(n4414) );
  CENX2 U3536 ( .A(n5441), .B(n2339), .Z(n5489) );
  CEO3X2 U3537 ( .A(n6632), .B(n6633), .C(n6631), .Z(n6662) );
  CENX1 U3538 ( .A(n5329), .B(n5328), .Z(n5330) );
  CND2X1 U3539 ( .A(n6233), .B(n6232), .Z(n6234) );
  CEO3X2 U3540 ( .A(n5072), .B(n5074), .C(n5073), .Z(n5044) );
  CND2XL U3541 ( .A(n5072), .B(n5073), .Z(n2474) );
  CND2XL U3542 ( .A(n5072), .B(n5074), .Z(n2475) );
  CND2X1 U3543 ( .A(n5073), .B(n5074), .Z(n2476) );
  CND2X1 U3544 ( .A(n5432), .B(n5434), .Z(n2478) );
  CND2X1 U3545 ( .A(n5432), .B(n5433), .Z(n2479) );
  CND2X1 U3546 ( .A(n5434), .B(n5433), .Z(n2480) );
  CND3X2 U3547 ( .A(n2478), .B(n2479), .C(n2480), .Z(n5398) );
  CND2X1 U3548 ( .A(n5302), .B(n5301), .Z(n5434) );
  CNIVX4 U3549 ( .A(n6974), .Z(n7065) );
  CND2X1 U3550 ( .A(n5845), .B(n5844), .Z(n5846) );
  COND1X1 U3551 ( .A(n5844), .B(n5845), .C(n5843), .Z(n5847) );
  CENX1 U3552 ( .A(n5845), .B(n5766), .Z(n5878) );
  COND2XL U3553 ( .A(n2396), .B(n7078), .C(n7171), .D(n7118), .Z(n7109) );
  COND2XL U3554 ( .A(n6719), .B(n7053), .C(n7171), .D(n7078), .Z(n7088) );
  COND2X1 U3555 ( .A(n7171), .B(n5863), .C(n6969), .D(n5763), .Z(n5845) );
  CND2X1 U3556 ( .A(n6428), .B(n6427), .Z(n6429) );
  CND2X1 U3557 ( .A(n6921), .B(n6919), .Z(n6922) );
  COND1X2 U3558 ( .A(n6589), .B(n6591), .C(n6590), .Z(n6574) );
  COND1X1 U3559 ( .A(n6285), .B(n7004), .C(n6284), .Z(n2481) );
  COND1X1 U3560 ( .A(n6285), .B(n2367), .C(n2405), .Z(n2482) );
  COND1X1 U3561 ( .A(n6285), .B(n2368), .C(n2406), .Z(n6927) );
  CND2XL U3562 ( .A(n5462), .B(n5356), .Z(n5357) );
  CENXL U3563 ( .A(n6038), .B(n6037), .Z(n6039) );
  CENX2 U3564 ( .A(n2556), .B(n5082), .Z(n5373) );
  CNIVX1 U3565 ( .A(n5001), .Z(n2483) );
  CND2X2 U3566 ( .A(n2484), .B(n2485), .Z(n2486) );
  CND2X4 U3567 ( .A(n2486), .B(n3344), .Z(n3346) );
  CIVX2 U3568 ( .A(q0[11]), .Z(n2484) );
  CIVX2 U3569 ( .A(n7864), .Z(n2485) );
  CND2X1 U3570 ( .A(n6812), .B(n6811), .Z(n6813) );
  CEO3X2 U3571 ( .A(n6085), .B(n6083), .C(n6084), .Z(n6089) );
  CND2X1 U3572 ( .A(n5679), .B(n5601), .Z(n2621) );
  CNIVX4 U3573 ( .A(n4737), .Z(n2487) );
  CNIVX4 U3574 ( .A(n4737), .Z(n2488) );
  CNIVX4 U3575 ( .A(n4737), .Z(n2489) );
  CNIVX4 U3576 ( .A(n4737), .Z(n2490) );
  CNIVX4 U3577 ( .A(n4737), .Z(n2491) );
  CND2X1 U3578 ( .A(n7862), .B(q0[2]), .Z(n2533) );
  COR2XL U3579 ( .A(n2449), .B(n5815), .Z(n5816) );
  CND2XL U3580 ( .A(n5686), .B(n5685), .Z(n2492) );
  CNIVX1 U3581 ( .A(n5492), .Z(n5494) );
  CND2X1 U3582 ( .A(n6570), .B(n6569), .Z(n6571) );
  COR2XL U3583 ( .A(n2436), .B(n4766), .Z(n4671) );
  CND3XL U3584 ( .A(n5784), .B(n5783), .C(n5782), .Z(n5785) );
  CND2X1 U3585 ( .A(n5784), .B(n5783), .Z(n5788) );
  CND2X1 U3586 ( .A(n5053), .B(n5628), .Z(n2496) );
  CND2X2 U3587 ( .A(n2494), .B(n2495), .Z(n2497) );
  CND2X2 U3588 ( .A(n2497), .B(n2496), .Z(n5608) );
  CIVX2 U3589 ( .A(n5053), .Z(n2494) );
  CIVXL U3590 ( .A(n5628), .Z(n2495) );
  CND2XL U3591 ( .A(n5627), .B(n5626), .Z(n2500) );
  CND2X1 U3592 ( .A(n2498), .B(n2499), .Z(n2501) );
  CND2X2 U3593 ( .A(n2500), .B(n2501), .Z(n5053) );
  CIVXL U3594 ( .A(n5627), .Z(n2498) );
  CIVXL U3595 ( .A(n5626), .Z(n2499) );
  CND2X1 U3596 ( .A(n5686), .B(n5685), .Z(n5835) );
  CNIVX1 U3597 ( .A(n6173), .Z(n2502) );
  CND2X2 U3598 ( .A(n2503), .B(n2504), .Z(n2506) );
  CND2X2 U3599 ( .A(n2505), .B(n2506), .Z(n5953) );
  CIVX2 U3600 ( .A(n6168), .Z(n2504) );
  CENXL U3601 ( .A(n5591), .B(n5592), .Z(n4998) );
  CND2X1 U3602 ( .A(n5020), .B(n5019), .Z(n5021) );
  CND2X1 U3603 ( .A(n5030), .B(n5029), .Z(n5031) );
  COND1X1 U3604 ( .A(n5030), .B(n5029), .C(n5028), .Z(n5032) );
  CND2X1 U3605 ( .A(n3542), .B(n3541), .Z(n3543) );
  CENXL U3606 ( .A(n5560), .B(n5559), .Z(n2507) );
  CND2X1 U3607 ( .A(n5180), .B(n5178), .Z(n5122) );
  COND1X1 U3608 ( .A(n5290), .B(n5287), .C(n5288), .Z(n5286) );
  CND2X4 U3609 ( .A(n4794), .B(n4793), .Z(n5024) );
  CND2X4 U3610 ( .A(n4785), .B(n4784), .Z(n5023) );
  CND2X2 U3611 ( .A(n5829), .B(n5828), .Z(n2508) );
  CND2XL U3612 ( .A(n5829), .B(n5828), .Z(n6087) );
  CIVXL U3613 ( .A(n5079), .Z(n2509) );
  COND1X1 U3614 ( .A(n5328), .B(n5331), .C(n5329), .Z(n5197) );
  CNIVXL U3615 ( .A(h0[4]), .Z(n2511) );
  CNIVX4 U3616 ( .A(h0[4]), .Z(n2512) );
  CNIVX4 U3617 ( .A(h0[4]), .Z(n2513) );
  CNIVX4 U3618 ( .A(n5711), .Z(n2514) );
  CNIVX4 U3619 ( .A(n5711), .Z(n2515) );
  COND1X2 U3620 ( .A(n5507), .B(n5506), .C(n5505), .Z(n5466) );
  CENX1 U3621 ( .A(q0[30]), .B(q0[29]), .Z(n2516) );
  CIVDX2 U3622 ( .A(q0[29]), .Z0(n4679), .Z1(n7090) );
  CENX1 U3623 ( .A(q0[30]), .B(q0[29]), .Z(n4800) );
  CND2X1 U3624 ( .A(n5014), .B(n5013), .Z(n5015) );
  CND2X2 U3625 ( .A(n2341), .B(n3343), .Z(n3347) );
  CND2X1 U3626 ( .A(n3345), .B(q0[11]), .Z(n3343) );
  CENX1 U3627 ( .A(n2279), .B(n5104), .Z(n5171) );
  CENX1 U3628 ( .A(n6305), .B(h0[14]), .Z(n6209) );
  CENXL U3629 ( .A(n5932), .B(h0[3]), .Z(n5157) );
  COND2X1 U3630 ( .A(n5160), .B(n5159), .C(n7537), .D(n5158), .Z(n5305) );
  CENX1 U3631 ( .A(n6647), .B(h0[12]), .Z(n4946) );
  CNR2X2 U3632 ( .A(n3737), .B(n3736), .Z(n3809) );
  CENX1 U3633 ( .A(n6647), .B(h0[31]), .Z(n6704) );
  CENX1 U3634 ( .A(n6647), .B(n5927), .Z(n5191) );
  CENXL U3635 ( .A(n6647), .B(n7674), .Z(n4486) );
  CENX1 U3636 ( .A(n6647), .B(h0[8]), .Z(n4479) );
  CENXL U3637 ( .A(n7539), .B(n6647), .Z(n3361) );
  CENXL U3638 ( .A(n6647), .B(n2512), .Z(n3787) );
  CENXL U3639 ( .A(n6647), .B(h0[3]), .Z(n3356) );
  CND2X1 U3640 ( .A(n5081), .B(n5083), .Z(n4843) );
  CEO3X2 U3641 ( .A(n5583), .B(n5581), .C(n5582), .Z(n5609) );
  CND2XL U3642 ( .A(n2401), .B(n5582), .Z(n2517) );
  CND2XL U3643 ( .A(n2401), .B(n5581), .Z(n2518) );
  CND2X1 U3644 ( .A(n5582), .B(n5581), .Z(n2519) );
  CND2X1 U3645 ( .A(n5002), .B(n5001), .Z(n5003) );
  COND2X1 U3646 ( .A(n7126), .B(n5798), .C(n5907), .D(n7124), .Z(n5889) );
  COND1X1 U3647 ( .A(n5092), .B(n5094), .C(n5091), .Z(n4972) );
  CNIVX1 U3648 ( .A(n6286), .Z(n6287) );
  CNIVX2 U3649 ( .A(n2433), .Z(n7253) );
  CND2X1 U3650 ( .A(n6142), .B(n5931), .Z(n2522) );
  CND2X2 U3651 ( .A(n2520), .B(n2521), .Z(n2523) );
  CND2X2 U3652 ( .A(n2522), .B(n2523), .Z(n6148) );
  CIVXL U3653 ( .A(n6142), .Z(n2520) );
  CIVX2 U3654 ( .A(n5931), .Z(n2521) );
  COND2X1 U3655 ( .A(n6114), .B(n5924), .C(n3368), .D(n6115), .Z(n6142) );
  CDLY1XL U3656 ( .A(q0[28]), .Z(n2524) );
  CND2X1 U3657 ( .A(n5509), .B(n5508), .Z(n5510) );
  CNR2X1 U3658 ( .A(n7020), .B(n6285), .Z(n6929) );
  CENX1 U3659 ( .A(n5448), .B(n5449), .Z(n4430) );
  CND2X1 U3660 ( .A(n5450), .B(n5449), .Z(n5451) );
  CND2X1 U3661 ( .A(n5597), .B(n1584), .Z(n5599) );
  CND2XL U3662 ( .A(n5211), .B(n5209), .Z(n4947) );
  CENX1 U3663 ( .A(n5211), .B(n5210), .Z(n5268) );
  COR2XL U3664 ( .A(n7009), .B(n7010), .Z(n7492) );
  CND2X1 U3665 ( .A(n5506), .B(n5507), .Z(n5509) );
  COND1X1 U3666 ( .A(n5507), .B(n5506), .C(n5505), .Z(n5508) );
  CEO3X2 U3667 ( .A(n5492), .B(n5493), .C(n5495), .Z(n5499) );
  CND2X1 U3668 ( .A(n6066), .B(n6134), .Z(n2528) );
  CND2X2 U3669 ( .A(n2527), .B(n2526), .Z(n2529) );
  CND2X2 U3670 ( .A(n2528), .B(n2529), .Z(n6172) );
  CIVX2 U3671 ( .A(n6134), .Z(n2526) );
  CIVX2 U3672 ( .A(n6066), .Z(n2527) );
  CND2X1 U3673 ( .A(n5250), .B(n5252), .Z(n5153) );
  COND1X1 U3674 ( .A(n5250), .B(n5252), .C(n5249), .Z(n5154) );
  CIVXL U3675 ( .A(n7461), .Z(n2530) );
  CND2X2 U3676 ( .A(n2533), .B(n2534), .Z(n3371) );
  CIVX2 U3677 ( .A(n7862), .Z(n2531) );
  CIVX2 U3678 ( .A(q0[2]), .Z(n2532) );
  CND2IX1 U3679 ( .B(n5398), .A(n2347), .Z(n5350) );
  CND2X2 U3680 ( .A(n5457), .B(n5456), .Z(n5488) );
  CND2X1 U3681 ( .A(n5838), .B(n5840), .Z(n2535) );
  CND2X2 U3682 ( .A(n2535), .B(n2536), .Z(n5767) );
  CEO3X2 U3683 ( .A(n5955), .B(n5957), .C(n2362), .Z(n6084) );
  CND2XL U3684 ( .A(n5955), .B(n5956), .Z(n2537) );
  CND2XL U3685 ( .A(n5955), .B(n5957), .Z(n2538) );
  CND3X1 U3686 ( .A(n2537), .B(n2538), .C(n2539), .Z(n6072) );
  CNIVX1 U3687 ( .A(n6072), .Z(n6008) );
  CNR2X1 U3688 ( .A(n7503), .B(n7501), .Z(n3735) );
  CND2X1 U3689 ( .A(n5369), .B(n5371), .Z(n4877) );
  CNR2X2 U3690 ( .A(n7275), .B(n7291), .Z(n7407) );
  COND1X2 U3691 ( .A(n5613), .B(n5614), .C(n5612), .Z(n5616) );
  CENXL U3692 ( .A(n7134), .B(h0[22]), .Z(n6718) );
  CENXL U3693 ( .A(n7134), .B(h0[23]), .Z(n6773) );
  CENXL U3694 ( .A(n7134), .B(h0[24]), .Z(n6827) );
  CENXL U3695 ( .A(n7134), .B(h0[27]), .Z(n7053) );
  CENXL U3696 ( .A(n7134), .B(h0[28]), .Z(n7078) );
  CENXL U3697 ( .A(n7134), .B(h0[29]), .Z(n7118) );
  CENXL U3698 ( .A(n7134), .B(h0[30]), .Z(n7135) );
  CENXL U3699 ( .A(n7134), .B(h0[19]), .Z(n6583) );
  CND2X1 U3700 ( .A(n5416), .B(n5415), .Z(n5417) );
  CENX1 U3701 ( .A(n5416), .B(n5415), .Z(n4415) );
  COND1X1 U3702 ( .A(n6219), .B(n6218), .C(n6217), .Z(n6222) );
  CND2X1 U3703 ( .A(n6122), .B(n6121), .Z(n6123) );
  CNR2X2 U3704 ( .A(n5511), .B(n5467), .Z(n5504) );
  CENX1 U3705 ( .A(q0[14]), .B(q0[13]), .Z(n2540) );
  CENX1 U3706 ( .A(q0[14]), .B(q0[13]), .Z(n5711) );
  CANR1X1 U3707 ( .A(n7151), .B(n7150), .C(n2473), .Z(n7352) );
  CENX2 U3708 ( .A(n5179), .B(n5180), .Z(n5325) );
  CENX2 U3709 ( .A(n5178), .B(n5177), .Z(n5179) );
  CEO3X2 U3710 ( .A(n6883), .B(n6884), .C(n2304), .Z(n6893) );
  COND2X2 U3711 ( .A(n5578), .B(n2566), .C(n2490), .D(n5765), .Z(n5722) );
  CENXL U3712 ( .A(n6490), .B(h0[23]), .Z(n6000) );
  CND2IXL U3713 ( .B(n7538), .A(n6490), .Z(n3462) );
  CENXL U3714 ( .A(n6490), .B(h0[22]), .Z(n5815) );
  CENXL U3715 ( .A(n7539), .B(n6490), .Z(n3461) );
  CENX2 U3716 ( .A(n5801), .B(n5800), .Z(n5716) );
  COND1X1 U3717 ( .A(n6712), .B(n6713), .C(n6711), .Z(n6716) );
  CND2IXL U3718 ( .B(n4834), .A(n4833), .Z(n4690) );
  COND1X2 U3719 ( .A(n5444), .B(n5443), .C(n5442), .Z(n5436) );
  CENXL U3720 ( .A(n5034), .B(n5035), .Z(n4660) );
  CND2X1 U3721 ( .A(n5076), .B(n5075), .Z(n2544) );
  CND2X2 U3722 ( .A(n2542), .B(n2543), .Z(n2545) );
  CND2X2 U3723 ( .A(n2544), .B(n2545), .Z(n5078) );
  CIVX2 U3724 ( .A(n5076), .Z(n2542) );
  CIVX2 U3725 ( .A(n5075), .Z(n2543) );
  CIVX3 U3726 ( .A(n7864), .Z(n5888) );
  CND2X1 U3727 ( .A(n5268), .B(n5267), .Z(n2548) );
  CND2X2 U3728 ( .A(n2546), .B(n2547), .Z(n2549) );
  CND2X2 U3729 ( .A(n2548), .B(n2549), .Z(n5269) );
  CIVX2 U3730 ( .A(n5268), .Z(n2546) );
  CIVX2 U3731 ( .A(n5267), .Z(n2547) );
  COND1X2 U3732 ( .A(n5222), .B(n5221), .C(n5220), .Z(n5267) );
  CND2X1 U3733 ( .A(n5774), .B(n5885), .Z(n2552) );
  CND2X2 U3734 ( .A(n2551), .B(n2550), .Z(n2553) );
  CIVX2 U3735 ( .A(n5885), .Z(n2550) );
  CIVX2 U3736 ( .A(n5774), .Z(n2551) );
  CIVXL U3737 ( .A(n4760), .Z(n2554) );
  CENX1 U3738 ( .A(q0[27]), .B(q0[28]), .Z(n2555) );
  CENX1 U3739 ( .A(q0[28]), .B(q0[27]), .Z(n4675) );
  CIVX3 U3740 ( .A(n2433), .Z(n6797) );
  CNIVX2 U3741 ( .A(n6170), .Z(n5954) );
  CNIVX4 U3742 ( .A(q0[1]), .Z(n3580) );
  CIVX3 U3743 ( .A(n6576), .Z(n5112) );
  CNR2X1 U3744 ( .A(n5035), .B(n5034), .Z(n5038) );
  COND2X1 U3745 ( .A(n6418), .B(n4661), .C(n5984), .D(n5050), .Z(n5034) );
  CENX1 U3746 ( .A(n2510), .B(n4411), .Z(n4496) );
  CENX1 U3747 ( .A(n3447), .B(n2510), .Z(n3493) );
  CENX4 U3748 ( .A(n4732), .B(n4782), .Z(n4733) );
  CNIVX1 U3749 ( .A(n5083), .Z(n2556) );
  COR2XL U3750 ( .A(n6974), .B(n5692), .Z(n5694) );
  CENX4 U3751 ( .A(n4734), .B(n4733), .Z(n4903) );
  CIVXL U3752 ( .A(n2607), .Z(n2557) );
  COR2XL U3753 ( .A(n6273), .B(n6274), .Z(n2558) );
  CIVX3 U3754 ( .A(n3352), .Z(n2560) );
  CIVX2 U3755 ( .A(n3352), .Z(n2561) );
  CIVX2 U3756 ( .A(n2560), .Z(n2562) );
  CIVX2 U3757 ( .A(n2561), .Z(n2563) );
  CIVX1 U3758 ( .A(n2560), .Z(n2564) );
  CIVX1 U3759 ( .A(n2560), .Z(n2565) );
  CIVX1 U3760 ( .A(n2561), .Z(n2566) );
  CIVX1 U3761 ( .A(n2561), .Z(n2567) );
  CIVX1 U3762 ( .A(n1588), .Z(n2568) );
  CIVX1 U3763 ( .A(n1588), .Z(n2570) );
  CIVX1 U3764 ( .A(n1588), .Z(n2571) );
  CIVX1 U3765 ( .A(n1588), .Z(n2572) );
  CIVX1 U3766 ( .A(n2560), .Z(n2573) );
  CIVXL U3767 ( .A(n2560), .Z(n2574) );
  CIVXL U3768 ( .A(n1588), .Z(n2575) );
  CIVXL U3769 ( .A(n1588), .Z(n2576) );
  CIVXL U3770 ( .A(n1588), .Z(n2577) );
  CIVXL U3771 ( .A(n2560), .Z(n2578) );
  CIVXL U3772 ( .A(n2560), .Z(n2579) );
  CIVXL U3773 ( .A(n2560), .Z(n2580) );
  CIVX4 U3774 ( .A(q0[9]), .Z(n3615) );
  CIVX4 U3775 ( .A(n7858), .Z(n6191) );
  CIVXL U3776 ( .A(n7375), .Z(n2581) );
  CND2X1 U3777 ( .A(n5443), .B(n5444), .Z(n5435) );
  CIVX4 U3778 ( .A(n4685), .Z(n7218) );
  CND2X2 U3779 ( .A(n3379), .B(n4670), .Z(n2584) );
  CND2X1 U3780 ( .A(n5249), .B(n5250), .Z(n2587) );
  CND2X2 U3781 ( .A(n2585), .B(n2586), .Z(n2588) );
  CND2X2 U3782 ( .A(n2587), .B(n2588), .Z(n5251) );
  CIVX2 U3783 ( .A(n5250), .Z(n2585) );
  CIVX2 U3784 ( .A(n5249), .Z(n2586) );
  CND2X1 U3785 ( .A(n3379), .B(n4670), .Z(n3382) );
  CND2X2 U3786 ( .A(n2600), .B(n2601), .Z(n3379) );
  COND2X2 U3787 ( .A(n4798), .B(n5160), .C(n7537), .D(n5046), .Z(n5064) );
  CND2X2 U3788 ( .A(n2589), .B(n2465), .Z(n2591) );
  CND2X2 U3789 ( .A(n2591), .B(n2590), .Z(n4396) );
  CIVX2 U3790 ( .A(n4390), .Z(n2589) );
  CND2X1 U3791 ( .A(n2507), .B(n5561), .Z(n2594) );
  CND2X2 U3792 ( .A(n2592), .B(n2593), .Z(n2595) );
  CND2X2 U3793 ( .A(n2594), .B(n2595), .Z(n5655) );
  CIVXL U3794 ( .A(n5561), .Z(n2592) );
  CND2X1 U3795 ( .A(n4880), .B(n4881), .Z(n4882) );
  COND1X2 U3796 ( .A(n7021), .B(n7018), .C(n7019), .Z(n7038) );
  CNIVX2 U3797 ( .A(n5604), .Z(n5010) );
  CIVX8 U3798 ( .A(n4684), .Z(n7171) );
  CNR2IX2 U3799 ( .B(n7539), .A(n7171), .Z(n5306) );
  CND2IX2 U3800 ( .B(n7171), .A(n6825), .Z(n6826) );
  CND2IX2 U3801 ( .B(n7171), .A(n6094), .Z(n6095) );
  CEO3XL U3802 ( .A(n2398), .B(n5658), .C(n5655), .Z(n2596) );
  CENX1 U3803 ( .A(n5723), .B(n5724), .Z(n5635) );
  COND2X2 U3804 ( .A(n2562), .B(n5908), .C(n2491), .D(n5933), .Z(n5969) );
  COND1X2 U3805 ( .A(n5489), .B(n5490), .C(n5488), .Z(n5459) );
  CENX2 U3806 ( .A(n6417), .B(h0[24]), .Z(n5867) );
  CIVX2 U3807 ( .A(n2606), .Z(n2597) );
  CND2X1 U3808 ( .A(n5490), .B(n5489), .Z(n5458) );
  CIVX2 U3809 ( .A(n7860), .Z(n2598) );
  CIVX2 U3810 ( .A(n7865), .Z(n2599) );
  CND2X1 U3811 ( .A(n4999), .B(n5596), .Z(n2604) );
  CIVX2 U3812 ( .A(n4999), .Z(n2602) );
  CIVXL U3813 ( .A(n5596), .Z(n2603) );
  CENX1 U3814 ( .A(n5589), .B(n4998), .Z(n5596) );
  COAN1XL U3815 ( .A(n7021), .B(n7018), .C(n7019), .Z(n2607) );
  CND2X1 U3816 ( .A(n5773), .B(n5772), .Z(n2608) );
  CND2XL U3817 ( .A(n5660), .B(n5659), .Z(n2609) );
  CND2X2 U3818 ( .A(n5660), .B(n5659), .Z(n5777) );
  COND1X2 U3819 ( .A(n5549), .B(n5523), .C(n5542), .Z(n5524) );
  CND2X1 U3820 ( .A(n5671), .B(n5672), .Z(n2612) );
  CND2X2 U3821 ( .A(n2610), .B(n2611), .Z(n2613) );
  CND2X2 U3822 ( .A(n2612), .B(n2613), .Z(n5651) );
  CIVX2 U3823 ( .A(n5671), .Z(n2610) );
  CIVX2 U3824 ( .A(n5672), .Z(n2611) );
  COND1X1 U3825 ( .A(n6288), .B(n6289), .C(n6287), .Z(n6291) );
  CND2X2 U3826 ( .A(n7466), .B(n7465), .Z(n7468) );
  CND2X1 U3827 ( .A(n6089), .B(n6090), .Z(n6093) );
  CNIVX8 U3828 ( .A(n4687), .Z(n7203) );
  COND1X1 U3829 ( .A(n6169), .B(n6170), .C(n2451), .Z(n2614) );
  COND1X1 U3830 ( .A(n6169), .B(n6170), .C(n2450), .Z(n6216) );
  CIVX3 U3831 ( .A(n7862), .Z(n5104) );
  CMX2XL U3832 ( .A0(h0_0[1]), .A1(h0[1]), .S(cmd2_en_0), .Z(n919) );
  CENXL U3833 ( .A(n3210), .B(h0[1]), .Z(n3203) );
  CENX1 U3834 ( .A(n7092), .B(h0[1]), .Z(n5169) );
  CENX1 U3835 ( .A(n6460), .B(h0[1]), .Z(n4955) );
  CNR2X1 U3836 ( .A(n5518), .B(n5517), .Z(n5555) );
  CIVXL U3837 ( .A(n7036), .Z(n2615) );
  CIVX3 U3838 ( .A(q0[15]), .Z(n4366) );
  CMX2XL U3839 ( .A0(h0[11]), .A1(h[11]), .S(pushin), .Z(n940) );
  CND2X1 U3840 ( .A(n2502), .B(n6172), .Z(n6176) );
  CENX1 U3841 ( .A(n7092), .B(h0[11]), .Z(n5690) );
  CEOX2 U3842 ( .A(n5958), .B(n5960), .Z(n2616) );
  CEOX2 U3843 ( .A(n2616), .B(n2453), .Z(n6090) );
  CND2X1 U3844 ( .A(n5959), .B(n5958), .Z(n2617) );
  CND2X1 U3845 ( .A(n5959), .B(n5960), .Z(n2618) );
  CND2X1 U3846 ( .A(n5958), .B(n5960), .Z(n2619) );
  CND3X2 U3847 ( .A(n2617), .B(n2618), .C(n2619), .Z(n6070) );
  COND1X1 U3848 ( .A(n6008), .B(n6070), .C(n6071), .Z(n6010) );
  CND2X1 U3849 ( .A(n2620), .B(n2402), .Z(n2622) );
  CND2X2 U3850 ( .A(n2621), .B(n2622), .Z(n5769) );
  CIVXL U3851 ( .A(n5679), .Z(n2620) );
  COND1X1 U3852 ( .A(n5672), .B(n5673), .C(n5671), .Z(n5675) );
  CIVX8 U3853 ( .A(n7853), .Z(n6103) );
  CND2X4 U3854 ( .A(n3367), .B(n3366), .Z(n3368) );
  CIVX2 U3855 ( .A(n6293), .Z(n5099) );
  COAN1X1 U3856 ( .A(n7291), .B(n7318), .C(n7289), .Z(n2625) );
  CIVX4 U3857 ( .A(n7538), .Z(n4399) );
  COND2X1 U3858 ( .A(n2420), .B(n5866), .C(n6770), .D(n5992), .Z(n5899) );
  CNR2X2 U3859 ( .A(n8013), .B(h0_1[2]), .Z(n2859) );
  CIVX2 U3860 ( .A(n2663), .Z(n2995) );
  CNIVXL U3861 ( .A(cmd2_en_2), .Z(n2865) );
  CIVX2 U3862 ( .A(n2865), .Z(n7751) );
  CIVX4 U3863 ( .A(n2670), .Z(n2758) );
  CMXI2XL U3864 ( .A0(n7062), .A1(q[27]), .S(n7682), .Z(n2626) );
  CMXI2XL U3865 ( .A0(n6491), .A1(q[13]), .S(n7682), .Z(n2627) );
  CMXI2XL U3866 ( .A0(q0[5]), .A1(q[5]), .S(n7682), .Z(n2628) );
  CNIVXL U3867 ( .A(out0_2[52]), .Z(n7677) );
  CNIVXL U3868 ( .A(out0_2[53]), .Z(n7678) );
  CIVXL U3869 ( .A(n5711), .Z(n5712) );
  CEOX1 U3870 ( .A(n7092), .B(h0[3]), .Z(n2657) );
  CNIVX4 U3871 ( .A(n5911), .Z(n4443) );
  CIVX3 U3872 ( .A(n4534), .Z(n2659) );
  CIVX8 U3873 ( .A(n4366), .Z(n2660) );
  CIVXL U3874 ( .A(n5306), .Z(n5162) );
  CIVXL U3875 ( .A(n2737), .Z(n2927) );
  CNR2IX4 U3876 ( .B(cmd1_en_2_d), .A(n2736), .Z(n2737) );
  CAN2X4 U3877 ( .A(cmd0_en_2_d), .B(cmd2_en_2), .Z(n2928) );
  CNIVX2 U3878 ( .A(pushin), .Z(n7682) );
  CNIVX1 U3879 ( .A(n8004), .Z(n4350) );
  COND1X2 U3880 ( .A(n3948), .B(n4151), .C(n3947), .Z(n3949) );
  CIVX2 U3881 ( .A(n6376), .Z(n3743) );
  CAN2X1 U3882 ( .A(n2704), .B(cmd0_2[0]), .Z(n4363) );
  COR2X1 U3883 ( .A(h0_1[1]), .B(h0_1[0]), .Z(n2663) );
  CMXI2X1 U3884 ( .A0(n3211), .A1(q[14]), .S(n7682), .Z(n2664) );
  CMXI2XL U3885 ( .A0(n6118), .A1(q[9]), .S(n7682), .Z(n2665) );
  CMXI2XL U3886 ( .A0(n4686), .A1(q[26]), .S(n7682), .Z(n2666) );
  CMXI2XL U3887 ( .A0(n5566), .A1(q[3]), .S(n7682), .Z(n2667) );
  CMXI2XL U3888 ( .A0(n3210), .A1(q[1]), .S(n7682), .Z(n2669) );
  CIVDX2 U3889 ( .A(n2764), .Z0(n2670), .Z1(n2671) );
  CIVDX2 U3890 ( .A(cmd1_en_2_d), .Z0(n3883), .Z1(n3902) );
  CMXI2XL U3891 ( .A0(n2659), .A1(q[23]), .S(n7682), .Z(n2672) );
  CMXI2XL U3892 ( .A0(n6460), .A1(q[25]), .S(n7682), .Z(n2673) );
  CMXI2XL U3893 ( .A0(n6699), .A1(q[17]), .S(n7682), .Z(n2674) );
  CMXI2XL U3894 ( .A0(n5932), .A1(q[21]), .S(n7682), .Z(n2675) );
  CMXI2XL U3895 ( .A0(n2660), .A1(q[15]), .S(n7682), .Z(n2676) );
  CMXI2XL U3896 ( .A0(n2456), .A1(q[19]), .S(n7682), .Z(n2677) );
  CMXI2XL U3897 ( .A0(n2597), .A1(q[11]), .S(n7682), .Z(n2678) );
  CMXI2XL U3898 ( .A0(n7090), .A1(q[29]), .S(n7682), .Z(n2679) );
  CMXI2XL U3899 ( .A0(n7279), .A1(q[31]), .S(n7682), .Z(n2681) );
  CMX2XL U3900 ( .A0(n2464), .A1(q[20]), .S(n7682), .Z(n2897) );
  CMX2XL U3901 ( .A0(h0[7]), .A1(h[7]), .S(pushin), .Z(n2894) );
  CMX2XL U3902 ( .A0(h0[8]), .A1(h[8]), .S(pushin), .Z(n2895) );
  CMX2XL U3903 ( .A0(h0[10]), .A1(h[10]), .S(pushin), .Z(n2896) );
  CMX2XL U3904 ( .A0(h0[13]), .A1(h[13]), .S(pushin), .Z(n2898) );
  CMX2XL U3905 ( .A0(h0[14]), .A1(h[14]), .S(pushin), .Z(n2899) );
  CMX2XL U3906 ( .A0(h0[15]), .A1(h[15]), .S(pushin), .Z(n2900) );
  CMX2XL U3907 ( .A0(h0[16]), .A1(h[16]), .S(pushin), .Z(n2901) );
  CMX2XL U3908 ( .A0(h0[18]), .A1(h[18]), .S(pushin), .Z(n2902) );
  CMX2XL U3909 ( .A0(h0[19]), .A1(h[19]), .S(pushin), .Z(n2903) );
  CMX2XL U3910 ( .A0(h0[22]), .A1(h[22]), .S(pushin), .Z(n2904) );
  CMX2XL U3911 ( .A0(h0[24]), .A1(h[24]), .S(pushin), .Z(n2905) );
  CMX2XL U3912 ( .A0(h0[25]), .A1(h[25]), .S(pushin), .Z(n2906) );
  CMX2XL U3913 ( .A0(h0[26]), .A1(h[26]), .S(pushin), .Z(n2907) );
  CMX2XL U3914 ( .A0(h0[27]), .A1(h[27]), .S(pushin), .Z(n2908) );
  CMX2XL U3915 ( .A0(h0[29]), .A1(h[29]), .S(pushin), .Z(n2909) );
  CMX2XL U3916 ( .A0(h0[31]), .A1(h[31]), .S(n7682), .Z(n2910) );
  CMX2XL U3917 ( .A0(q0[6]), .A1(q[6]), .S(n7682), .Z(n2941) );
  CIVX8 U3918 ( .A(n3643), .Z(n5923) );
  CMXI2XL U3919 ( .A0(q0[10]), .A1(q[10]), .S(n7682), .Z(n2682) );
  COND11X1 U3920 ( .A(n3075), .B(n3032), .C(n3031), .D(n3030), .Z(n3033) );
  COND2X1 U3921 ( .A(n2865), .B(n4279), .C(n3093), .D(n3092), .Z(n3094) );
  CNIVX1 U3922 ( .A(cmd1_en_2), .Z(n7846) );
  CNIVXL U3923 ( .A(out0_2[32]), .Z(n2966) );
  CNIVXL U3924 ( .A(out0_2[0]), .Z(n4361) );
  CNIVXL U3925 ( .A(out0_2[55]), .Z(n4323) );
  CNR2X1 U3927 ( .A(n8004), .B(cmd0_2[1]), .Z(n2704) );
  CND2X1 U3928 ( .A(n2704), .B(n7937), .Z(n2685) );
  CND2X1 U3929 ( .A(out2_2[15]), .B(out2_2[16]), .Z(n3299) );
  CND2XL U3930 ( .A(out2_2[17]), .B(out2_2[18]), .Z(n2686) );
  CNR2X1 U3931 ( .A(n3299), .B(n2686), .Z(n3213) );
  CND2XL U3932 ( .A(out2_2[19]), .B(out2_2[20]), .Z(n3294) );
  CND2XL U3933 ( .A(out2_2[21]), .B(out2_2[22]), .Z(n2687) );
  CNR2X1 U3934 ( .A(n3294), .B(n2687), .Z(n2688) );
  CND2X1 U3935 ( .A(n3213), .B(n2688), .Z(n3268) );
  CND2XL U3936 ( .A(out2_2[23]), .B(out2_2[24]), .Z(n3300) );
  CND2XL U3937 ( .A(out2_2[25]), .B(out2_2[26]), .Z(n2689) );
  CNR2X1 U3938 ( .A(n3300), .B(n2689), .Z(n3270) );
  CND2XL U3939 ( .A(out2_2[27]), .B(out2_2[28]), .Z(n4315) );
  CND2XL U3940 ( .A(out2_2[29]), .B(out2_2[30]), .Z(n2690) );
  CNR2X1 U3941 ( .A(n4315), .B(n2690), .Z(n2691) );
  CND2X1 U3942 ( .A(n3270), .B(n2691), .Z(n2692) );
  CNR2X1 U3943 ( .A(n3268), .B(n2692), .Z(n2699) );
  CND2XL U3944 ( .A(out2_2[7]), .B(out2_2[8]), .Z(n3312) );
  CND2XL U3945 ( .A(out2_2[11]), .B(out2_2[12]), .Z(n2735) );
  CND2XL U3946 ( .A(out2_2[13]), .B(out2_2[14]), .Z(n2693) );
  CNR2X1 U3947 ( .A(n2735), .B(n2693), .Z(n2694) );
  CND2X1 U3948 ( .A(n2734), .B(n2694), .Z(n2698) );
  CND2XL U3949 ( .A(out2_2[3]), .B(out2_2[4]), .Z(n2731) );
  CND2XL U3950 ( .A(out2_2[5]), .B(out2_2[6]), .Z(n2695) );
  CNR2X1 U3951 ( .A(n2731), .B(n2695), .Z(n2697) );
  CND2XL U3952 ( .A(out2_2[1]), .B(out2_2[2]), .Z(n2696) );
  CND2X1 U3953 ( .A(out2_2[0]), .B(roundit), .Z(n4364) );
  CNR2X1 U3954 ( .A(n2696), .B(n4364), .Z(n2730) );
  CND2X1 U3955 ( .A(n2697), .B(n2730), .Z(n2733) );
  CNR2X2 U3956 ( .A(n2698), .B(n2733), .Z(n3269) );
  CND2X2 U3957 ( .A(n2699), .B(n3269), .Z(n4292) );
  CND2XL U3958 ( .A(out2_2[31]), .B(out2_2[32]), .Z(n2945) );
  CND2XL U3959 ( .A(out2_2[33]), .B(out2_2[34]), .Z(n2700) );
  CNR2X1 U3960 ( .A(n2945), .B(n2700), .Z(n4291) );
  CND2XL U3961 ( .A(out2_2[35]), .B(out2_2[36]), .Z(n4293) );
  CND2XL U3962 ( .A(out2_2[37]), .B(out2_2[38]), .Z(n2701) );
  CNR2X1 U3963 ( .A(n4293), .B(n2701), .Z(n2702) );
  CND2X1 U3964 ( .A(n4291), .B(n2702), .Z(n3225) );
  CND2XL U3965 ( .A(out2_2[39]), .B(out2_2[40]), .Z(n3231) );
  CND2XL U3966 ( .A(out2_2[41]), .B(out2_2[42]), .Z(n2703) );
  CNR2XL U3967 ( .A(n3231), .B(n2703), .Z(n2708) );
  CND2XL U3968 ( .A(out2_2[43]), .B(out2_2[44]), .Z(n2706) );
  CAN3X2 U3969 ( .A(n7937), .B(cmd0_2[1]), .C(push0_2), .Z(n4344) );
  CND2XL U3970 ( .A(out2_2[45]), .B(out2_2[46]), .Z(n2705) );
  CNR2XL U3971 ( .A(n2706), .B(n2705), .Z(n2707) );
  CND2XL U3972 ( .A(n2708), .B(n2707), .Z(n2709) );
  CNR2X1 U3973 ( .A(n3225), .B(n2709), .Z(n3242) );
  CND2XL U3974 ( .A(out2_2[47]), .B(out2_2[48]), .Z(n3247) );
  CND2XL U3975 ( .A(out2_2[49]), .B(out2_2[50]), .Z(n2710) );
  CNR2X1 U3976 ( .A(n3247), .B(n2710), .Z(n2717) );
  CND2XL U3977 ( .A(out2_2[51]), .B(out2_2[52]), .Z(n2719) );
  CND2XL U3978 ( .A(out2_2[55]), .B(out2_2[56]), .Z(n2729) );
  CND2XL U3979 ( .A(out2_2[57]), .B(out2_2[58]), .Z(n2711) );
  CNR2X1 U3980 ( .A(n2729), .B(n2711), .Z(n3262) );
  CNR2XL U3981 ( .A(n7945), .B(n7942), .Z(n2712) );
  CND2XL U3982 ( .A(n3262), .B(n2712), .Z(n2713) );
  CNR2XL U3983 ( .A(n2726), .B(n2713), .Z(n2714) );
  CND2XL U3984 ( .A(n3242), .B(n2714), .Z(n2715) );
  CNR2X1 U3985 ( .A(n2715), .B(n4292), .Z(n2720) );
  CND2XL U3986 ( .A(n3242), .B(n2717), .Z(n2718) );
  CNR2X1 U3987 ( .A(n2718), .B(n4292), .Z(n3253) );
  CHA1XL U3988 ( .A(out2_2[61]), .B(n2720), .CO(n3266), .S(n2716) );
  CEOXL U3989 ( .A(out2_2[63]), .B(n2721), .Z(n2722) );
  CND2XL U3990 ( .A(n2722), .B(n4344), .Z(n2724) );
  CANR2XL U3991 ( .A(n4363), .B(out1_2[63]), .C(acc[63]), .D(n4350), .Z(n2723)
         );
  COND3X1 U3992 ( .A(n8011), .B(n2685), .C(n2724), .D(n2723), .Z(n2725) );
  CIVXL U3993 ( .A(n2726), .Z(n2727) );
  CND2XL U3994 ( .A(n3242), .B(n2727), .Z(n2728) );
  CNR2X1 U3995 ( .A(n2728), .B(n4292), .Z(n4281) );
  CNIVX1 U3996 ( .A(out0_2[5]), .Z(n4377) );
  CIVXL U3997 ( .A(n2730), .Z(n2944) );
  CNR2XL U3998 ( .A(n2944), .B(n2731), .Z(n2732) );
  CIVXL U3999 ( .A(out2_2[5]), .Z(n2891) );
  CNIVX1 U4000 ( .A(out0_2[6]), .Z(n4376) );
  CNIVX1 U4001 ( .A(out0_2[7]), .Z(n4375) );
  CIVX1 U4002 ( .A(n2733), .Z(n3339) );
  CIVXL U4003 ( .A(out2_2[7]), .Z(n4270) );
  CNIVX1 U4004 ( .A(out0_2[13]), .Z(n4382) );
  CND2X1 U4005 ( .A(n3339), .B(n2734), .Z(n3319) );
  CIVX2 U4006 ( .A(n3319), .Z(n3313) );
  CNIVX1 U4007 ( .A(out0_2[15]), .Z(n4380) );
  CIVX1 U4008 ( .A(n3269), .Z(n3321) );
  CIVX1 U4009 ( .A(cmd0_en_2_d), .Z(n2948) );
  CND2X1 U4010 ( .A(n2948), .B(cmd2_en_2), .Z(n2736) );
  CNR2X1 U4011 ( .A(n2736), .B(cmd1_en_2_d), .Z(n2764) );
  CND2XL U4012 ( .A(n2764), .B(acc[62]), .Z(n2740) );
  CND2XL U4013 ( .A(n2737), .B(out1_2[62]), .Z(n2739) );
  CND2XL U4014 ( .A(n2928), .B(out0_2[62]), .Z(n2738) );
  CND3XL U4015 ( .A(n2740), .B(n2739), .C(n2738), .Z(n2976) );
  CND2X1 U4016 ( .A(h0_1[0]), .B(h0_1[1]), .Z(n7766) );
  CIVXL U4017 ( .A(n3065), .Z(n2748) );
  CND2X1 U4018 ( .A(n8013), .B(h0_1[2]), .Z(n7744) );
  CND2XL U4019 ( .A(n2671), .B(acc[58]), .Z(n2743) );
  CND2XL U4020 ( .A(n2737), .B(out1_2[58]), .Z(n2742) );
  CND2XL U4021 ( .A(n2928), .B(out0_2[58]), .Z(n2741) );
  CND3XL U4022 ( .A(n2743), .B(n2742), .C(n2741), .Z(n2977) );
  CND2X1 U4023 ( .A(n2758), .B(acc[63]), .Z(n2746) );
  CND2XL U4024 ( .A(n2737), .B(out1_2[63]), .Z(n2745) );
  CND2X1 U4025 ( .A(n2928), .B(out0_2[63]), .Z(n2744) );
  CND3X1 U4026 ( .A(n2746), .B(n2745), .C(n2744), .Z(n2974) );
  CND2X1 U4027 ( .A(n2974), .B(n2995), .Z(n2934) );
  CIVX1 U4028 ( .A(n2934), .Z(n3064) );
  CANR2XL U4029 ( .A(n3066), .B(n7582), .C(n3064), .D(n2859), .Z(n2747) );
  COND1XL U4030 ( .A(n2748), .B(n7744), .C(n2747), .Z(n7716) );
  CAOR2X2 U4031 ( .A(out2_2[55]), .B(n7751), .C(n7716), .D(n7738), .Z(n875) );
  CANR2XL U4032 ( .A(n2995), .B(n2969), .C(n3169), .D(n2967), .Z(n2750) );
  CANR2XL U4033 ( .A(n3173), .B(n2981), .C(n3172), .D(n2970), .Z(n2749) );
  CND2X1 U4034 ( .A(n2750), .B(n2749), .Z(n3137) );
  CANR2XL U4035 ( .A(n3137), .B(n7582), .C(n7755), .D(n3136), .Z(n2752) );
  CND2X1 U4036 ( .A(h0_1[3]), .B(h0_1[2]), .Z(n7758) );
  CANR2XL U4037 ( .A(n2859), .B(n3122), .C(n7747), .D(n3118), .Z(n2751) );
  CND2X1 U4038 ( .A(n2752), .B(n2751), .Z(n7752) );
  CAOR2X2 U4039 ( .A(out2_2[49]), .B(n7751), .C(n7752), .D(n7738), .Z(n878) );
  CND2XL U4040 ( .A(h0_1[5]), .B(h0_1[4]), .Z(n4267) );
  CIVX1 U4041 ( .A(n4267), .Z(n4272) );
  CND2XL U4042 ( .A(n2973), .B(n3173), .Z(n2756) );
  CND2XL U4043 ( .A(n2977), .B(n2995), .Z(n2755) );
  CND2XL U4044 ( .A(n2975), .B(n3172), .Z(n2754) );
  CND2XL U4045 ( .A(n2979), .B(n3169), .Z(n2753) );
  CND4X1 U4046 ( .A(n2756), .B(n2755), .C(n2754), .D(n2753), .Z(n3034) );
  CND2XL U4047 ( .A(n3034), .B(n8012), .Z(n2757) );
  COND1XL U4048 ( .A(n8012), .B(n3037), .C(n2757), .Z(n2841) );
  CND2XL U4049 ( .A(n2841), .B(n8013), .Z(n7737) );
  CANR2XL U4050 ( .A(n7582), .B(n3038), .C(n7755), .D(n3041), .Z(n2761) );
  CND2XL U4051 ( .A(n3040), .B(n2859), .Z(n2760) );
  CND2XL U4052 ( .A(n3035), .B(n7747), .Z(n2759) );
  CND3XL U4053 ( .A(n2761), .B(n2760), .C(n2759), .Z(n7735) );
  CNR2XL U4054 ( .A(n8016), .B(h0_1[4]), .Z(n2919) );
  CIVX1 U4055 ( .A(n2919), .Z(n4266) );
  CNR2X1 U4056 ( .A(n7553), .B(n7729), .Z(n4251) );
  CANR2X1 U4057 ( .A(n2737), .B(out1_2[12]), .C(n2928), .D(out0_2[12]), .Z(
        n2762) );
  COND1XL U4058 ( .A(n2670), .B(n8017), .C(n2762), .Z(n3131) );
  CAOR2XL U4059 ( .A(out0_2[10]), .B(n2928), .C(n2737), .D(out1_2[10]), .Z(
        n2763) );
  CANR1XL U4060 ( .A(n2758), .B(acc[10]), .C(n2763), .Z(n3144) );
  CNR2XL U4061 ( .A(n3144), .B(n2663), .Z(n2768) );
  CIVXL U4062 ( .A(acc[13]), .Z(n3899) );
  CANR2X1 U4063 ( .A(n2737), .B(out1_2[13]), .C(n2928), .D(out0_2[13]), .Z(
        n2765) );
  COND1XL U4064 ( .A(n2670), .B(n3899), .C(n2765), .Z(n3129) );
  CANR2X1 U4065 ( .A(n2737), .B(out1_2[11]), .C(n2928), .D(out0_2[11]), .Z(
        n2766) );
  COND1XL U4066 ( .A(n2670), .B(n8018), .C(n2766), .Z(n3146) );
  CAOR2XL U4067 ( .A(n3173), .B(n3129), .C(n3169), .D(n3146), .Z(n2767) );
  CANR3XL U4068 ( .A(n3172), .B(n3131), .C(n2768), .D(n2767), .Z(n7559) );
  CNR2X1 U4069 ( .A(n7729), .B(n7744), .Z(n4249) );
  CIVX1 U4070 ( .A(n4249), .Z(n3148) );
  CANR2X1 U4071 ( .A(n2737), .B(out1_2[17]), .C(n2928), .D(out0_2[17]), .Z(
        n2769) );
  COND1XL U4072 ( .A(n2670), .B(n8014), .C(n2769), .Z(n3099) );
  CIVXL U4073 ( .A(acc[15]), .Z(n3904) );
  CANR2X1 U4074 ( .A(n2737), .B(out1_2[15]), .C(n2928), .D(out0_2[15]), .Z(
        n2770) );
  COND1XL U4075 ( .A(n2670), .B(n3904), .C(n2770), .Z(n3130) );
  CIVXL U4076 ( .A(out1_2[14]), .Z(n2772) );
  CANR2XL U4077 ( .A(n2671), .B(acc[14]), .C(out0_2[14]), .D(n2928), .Z(n2771)
         );
  COND1XL U4078 ( .A(n2772), .B(n2927), .C(n2771), .Z(n3132) );
  CANR2X1 U4079 ( .A(n2737), .B(out1_2[16]), .C(n2928), .D(out0_2[16]), .Z(
        n2773) );
  COND1XL U4080 ( .A(n2670), .B(n8015), .C(n2773), .Z(n3098) );
  CIVXL U4081 ( .A(acc[24]), .Z(n3863) );
  CANR2XL U4082 ( .A(n2737), .B(out1_2[24]), .C(n2928), .D(out0_2[24]), .Z(
        n2774) );
  COND1XL U4083 ( .A(n2670), .B(n3863), .C(n2774), .Z(n3013) );
  CIVXL U4084 ( .A(acc[23]), .Z(n3861) );
  CANR2XL U4085 ( .A(n2737), .B(out1_2[23]), .C(n2928), .D(out0_2[23]), .Z(
        n2775) );
  COND1XL U4086 ( .A(n2670), .B(n3861), .C(n2775), .Z(n3103) );
  CANR2XL U4087 ( .A(n3172), .B(n3013), .C(n3169), .D(n3103), .Z(n2779) );
  CIVXL U4088 ( .A(acc[22]), .Z(n3859) );
  CANR2XL U4089 ( .A(n2737), .B(out1_2[22]), .C(out0_2[22]), .D(n2928), .Z(
        n2776) );
  COND1XL U4090 ( .A(n3859), .B(n2670), .C(n2776), .Z(n3106) );
  CIVXL U4091 ( .A(acc[25]), .Z(n3865) );
  CANR2XL U4092 ( .A(n2737), .B(out1_2[25]), .C(n2928), .D(out0_2[25]), .Z(
        n2777) );
  COND1XL U4093 ( .A(n2670), .B(n3865), .C(n2777), .Z(n3015) );
  CANR2XL U4094 ( .A(n2995), .B(n3106), .C(n3173), .D(n3015), .Z(n2778) );
  CAN2X1 U4095 ( .A(n2779), .B(n2778), .Z(n3115) );
  CIVXL U4096 ( .A(n3115), .Z(n2780) );
  CNR2X1 U4097 ( .A(n7729), .B(n7758), .Z(n3192) );
  CIVX2 U4098 ( .A(n3192), .Z(n4254) );
  COND2XL U4099 ( .A(n3148), .B(n7557), .C(n2780), .D(n4254), .Z(n2788) );
  CIVX2 U4100 ( .A(n7729), .Z(n3074) );
  CND2X1 U4101 ( .A(n7762), .B(n3074), .Z(n3175) );
  CIVXL U4102 ( .A(acc[18]), .Z(n3851) );
  CANR2XL U4103 ( .A(n2737), .B(out1_2[18]), .C(n2928), .D(out0_2[18]), .Z(
        n2781) );
  COND1XL U4104 ( .A(n2670), .B(n3851), .C(n2781), .Z(n3100) );
  CIVXL U4105 ( .A(acc[19]), .Z(n3853) );
  CANR2XL U4106 ( .A(n2737), .B(out1_2[19]), .C(n2928), .D(out0_2[19]), .Z(
        n2782) );
  COND1XL U4107 ( .A(n2670), .B(n3853), .C(n2782), .Z(n3097) );
  CANR2XL U4108 ( .A(n2995), .B(n3100), .C(n3169), .D(n3097), .Z(n2786) );
  CIVXL U4109 ( .A(acc[21]), .Z(n3857) );
  CANR2XL U4110 ( .A(n2737), .B(out1_2[21]), .C(n2928), .D(out0_2[21]), .Z(
        n2783) );
  COND1XL U4111 ( .A(n2670), .B(n3857), .C(n2783), .Z(n3105) );
  CIVXL U4112 ( .A(acc[20]), .Z(n3855) );
  CANR2XL U4113 ( .A(n2737), .B(out1_2[20]), .C(out0_2[20]), .D(n2928), .Z(
        n2784) );
  COND1XL U4114 ( .A(n3855), .B(n2670), .C(n2784), .Z(n3104) );
  CANR2XL U4115 ( .A(n3173), .B(n3105), .C(n3172), .D(n3104), .Z(n2785) );
  CND2X1 U4116 ( .A(n2786), .B(n2785), .Z(n3113) );
  COND1XL U4117 ( .A(n3175), .B(n3113), .C(n8019), .Z(n2787) );
  CANR3XL U4118 ( .A(n4251), .B(n7559), .C(n2788), .D(n2787), .Z(n2834) );
  CND2XL U4119 ( .A(n2671), .B(acc[29]), .Z(n2791) );
  CND2XL U4120 ( .A(n2737), .B(out1_2[29]), .Z(n2790) );
  CND2XL U4121 ( .A(n2928), .B(out0_2[29]), .Z(n2789) );
  CND3XL U4122 ( .A(n2791), .B(n2790), .C(n2789), .Z(n3008) );
  CND2XL U4123 ( .A(n2671), .B(acc[26]), .Z(n2794) );
  CND2XL U4124 ( .A(n2737), .B(out1_2[26]), .Z(n2793) );
  CND2XL U4125 ( .A(n2928), .B(out0_2[26]), .Z(n2792) );
  CND3XL U4126 ( .A(n2794), .B(n2793), .C(n2792), .Z(n3012) );
  CND2XL U4127 ( .A(n2671), .B(acc[28]), .Z(n2797) );
  CND2XL U4128 ( .A(n2737), .B(out1_2[28]), .Z(n2796) );
  CND2XL U4129 ( .A(n2928), .B(out0_2[28]), .Z(n2795) );
  CND3XL U4130 ( .A(n2797), .B(n2796), .C(n2795), .Z(n3011) );
  CND2XL U4131 ( .A(n2671), .B(acc[37]), .Z(n2800) );
  CND2XL U4132 ( .A(n2737), .B(out1_2[37]), .Z(n2799) );
  CND2XL U4133 ( .A(n2928), .B(out0_2[37]), .Z(n2798) );
  CND3XL U4134 ( .A(n2800), .B(n2799), .C(n2798), .Z(n3017) );
  CND2XL U4135 ( .A(n2671), .B(acc[34]), .Z(n2803) );
  CND2XL U4136 ( .A(n2737), .B(out1_2[34]), .Z(n2802) );
  CND2XL U4137 ( .A(n2928), .B(out0_2[34]), .Z(n2801) );
  CND3XL U4138 ( .A(n2803), .B(n2802), .C(n2801), .Z(n3005) );
  CND2XL U4139 ( .A(n2671), .B(acc[36]), .Z(n2806) );
  CND2XL U4140 ( .A(n2737), .B(out1_2[36]), .Z(n2805) );
  CND2XL U4141 ( .A(n2928), .B(out0_2[36]), .Z(n2804) );
  CND3XL U4142 ( .A(n2806), .B(n2805), .C(n2804), .Z(n3020) );
  CND2XL U4143 ( .A(n2671), .B(acc[31]), .Z(n2809) );
  CND2XL U4144 ( .A(n2737), .B(out1_2[31]), .Z(n2808) );
  CND2XL U4145 ( .A(n2928), .B(out0_2[31]), .Z(n2807) );
  CND3XL U4146 ( .A(n2809), .B(n2808), .C(n2807), .Z(n3009) );
  CND2XL U4147 ( .A(n3009), .B(n3169), .Z(n2822) );
  CND2XL U4148 ( .A(n2671), .B(acc[33]), .Z(n2812) );
  CND2XL U4149 ( .A(n2737), .B(out1_2[33]), .Z(n2811) );
  CND2XL U4150 ( .A(n2928), .B(out0_2[33]), .Z(n2810) );
  CND3XL U4151 ( .A(n2812), .B(n2811), .C(n2810), .Z(n3004) );
  CND2XL U4152 ( .A(n3004), .B(n3173), .Z(n2821) );
  CND2XL U4153 ( .A(n2671), .B(acc[30]), .Z(n2815) );
  CND2XL U4154 ( .A(n2737), .B(out1_2[30]), .Z(n2814) );
  CND2XL U4155 ( .A(n2928), .B(out0_2[30]), .Z(n2813) );
  CND3XL U4156 ( .A(n2815), .B(n2814), .C(n2813), .Z(n3010) );
  CND2XL U4157 ( .A(n3010), .B(n2995), .Z(n2820) );
  CND2XL U4158 ( .A(n2671), .B(acc[32]), .Z(n2818) );
  CND2XL U4159 ( .A(n2737), .B(out1_2[32]), .Z(n2817) );
  CND2XL U4160 ( .A(n2928), .B(out0_2[32]), .Z(n2816) );
  CND3XL U4161 ( .A(n2818), .B(n2817), .C(n2816), .Z(n3003) );
  CND2XL U4162 ( .A(n3003), .B(n3172), .Z(n2819) );
  CND4X1 U4163 ( .A(n2822), .B(n2821), .C(n2820), .D(n2819), .Z(n3048) );
  CAOR2XL U4164 ( .A(n2859), .B(n3051), .C(n7755), .D(n3048), .Z(n2823) );
  CANR1XL U4165 ( .A(n7582), .B(n3114), .C(n2823), .Z(n2852) );
  CNR2X1 U4166 ( .A(n8020), .B(h0_1[5]), .Z(n7543) );
  CND2XL U4167 ( .A(n2671), .B(acc[39]), .Z(n2826) );
  CND2XL U4168 ( .A(n2737), .B(out1_2[39]), .Z(n2825) );
  CND2XL U4169 ( .A(n2928), .B(out0_2[39]), .Z(n2824) );
  CND3XL U4170 ( .A(n2826), .B(n2825), .C(n2824), .Z(n3019) );
  CND2XL U4171 ( .A(n2671), .B(acc[41]), .Z(n2829) );
  CND2XL U4172 ( .A(n2737), .B(out1_2[41]), .Z(n2828) );
  CND2XL U4173 ( .A(n2928), .B(out0_2[41]), .Z(n2827) );
  CND3XL U4174 ( .A(n2829), .B(n2828), .C(n2827), .Z(n2989) );
  CND2XL U4175 ( .A(n2671), .B(acc[40]), .Z(n2832) );
  CND2XL U4176 ( .A(n2737), .B(out1_2[40]), .Z(n2831) );
  CND2XL U4177 ( .A(n2928), .B(out0_2[40]), .Z(n2830) );
  CND3XL U4178 ( .A(n2832), .B(n2831), .C(n2830), .Z(n2988) );
  CND2XL U4179 ( .A(n3039), .B(n7747), .Z(n2851) );
  CND3XL U4180 ( .A(n2852), .B(n7543), .C(n2851), .Z(n2833) );
  COND3XL U4181 ( .A(n7735), .B(n4266), .C(n2834), .D(n2833), .Z(n2836) );
  CND2XL U4182 ( .A(n7751), .B(out2_2[10]), .Z(n2835) );
  COND4CXL U4183 ( .A(n4272), .B(n7737), .C(n2836), .D(n2835), .Z(n2837) );
  CNIVXL U4184 ( .A(h0_1[3]), .Z(n7680) );
  CND2XL U4185 ( .A(n3035), .B(n7755), .Z(n2839) );
  CND2XL U4186 ( .A(n3040), .B(n7582), .Z(n2838) );
  CND2X1 U4187 ( .A(n2839), .B(n2838), .Z(n2840) );
  CANR1XL U4188 ( .A(n7680), .B(n2841), .C(n2840), .Z(n7723) );
  CIVX1 U4189 ( .A(n7724), .Z(n7771) );
  CIVX2 U4190 ( .A(n7543), .Z(n7727) );
  CANR2XL U4191 ( .A(n7582), .B(n3051), .C(n7755), .D(n3039), .Z(n2844) );
  CND2XL U4192 ( .A(n3041), .B(n7747), .Z(n2843) );
  CND2XL U4193 ( .A(n3038), .B(n2859), .Z(n2842) );
  CND3XL U4194 ( .A(n2844), .B(n2843), .C(n2842), .Z(n7720) );
  CND2XL U4195 ( .A(n3114), .B(n2859), .Z(n7550) );
  CIVXL U4196 ( .A(n3113), .Z(n2845) );
  COND2XL U4197 ( .A(n7553), .B(n2845), .C(n3115), .D(n7744), .Z(n2846) );
  CANR1XL U4198 ( .A(n7747), .B(n3048), .C(n2846), .Z(n7551) );
  CNR2X1 U4199 ( .A(h0_1[4]), .B(h0_1[6]), .Z(n7726) );
  CNR2X1 U4200 ( .A(n7724), .B(n7726), .Z(n3075) );
  CANR11XL U4201 ( .A(n3074), .B(n7550), .C(n7551), .D(n3075), .Z(n2847) );
  COND1XL U4202 ( .A(n7727), .B(n7720), .C(n2847), .Z(n2849) );
  CND2XL U4203 ( .A(n7751), .B(out2_2[18]), .Z(n2848) );
  COND4CXL U4204 ( .A(n7723), .B(n7771), .C(n2849), .D(n2848), .Z(n2850) );
  CNIVX1 U4205 ( .A(out0_2[3]), .Z(n4379) );
  CIVXL U4206 ( .A(out2_2[3]), .Z(n3198) );
  CND3XL U4207 ( .A(n2852), .B(n3074), .C(n2851), .Z(n2853) );
  CIVXL U4208 ( .A(n3075), .Z(n3055) );
  COND3XL U4209 ( .A(n7727), .B(n7735), .C(n2853), .D(n3055), .Z(n2855) );
  CND2XL U4210 ( .A(n7751), .B(out2_2[26]), .Z(n2854) );
  COND4CXL U4211 ( .A(n7771), .B(n7737), .C(n2855), .D(n2854), .Z(n2856) );
  CANR2XL U4212 ( .A(n2859), .B(n3035), .C(n7755), .D(n3040), .Z(n2858) );
  CANR2XL U4213 ( .A(n7582), .B(n3041), .C(n7747), .D(n3034), .Z(n2857) );
  CND2X1 U4214 ( .A(n2858), .B(n2857), .Z(n7693) );
  CNR2XL U4215 ( .A(n3037), .B(n7553), .Z(n7692) );
  CIVDX1 U4216 ( .A(n2859), .Z0(n2662), .Z1(n7762) );
  CANR2XL U4217 ( .A(n7747), .B(n3038), .C(n7762), .D(n3039), .Z(n2861) );
  CANR2XL U4218 ( .A(n7582), .B(n3048), .C(n7755), .D(n3051), .Z(n2860) );
  CND2XL U4219 ( .A(n2861), .B(n2860), .Z(n3116) );
  CAOR2X2 U4220 ( .A(out2_2[53]), .B(n7751), .C(n7689), .D(n7738), .Z(n879) );
  CMX2XL U4221 ( .A0(h0_1[0]), .A1(h0_0[0]), .S(cmd2_en_1), .Z(n2863) );
  CMX2XL U4222 ( .A0(h0_1[1]), .A1(h0_0[1]), .S(cmd2_en_1), .Z(n2864) );
  CANR2XL U4223 ( .A(n3173), .B(n2994), .C(n3172), .D(n2987), .Z(n2867) );
  CANR2XL U4224 ( .A(n2995), .B(n2989), .C(n3169), .D(n2990), .Z(n2866) );
  CND2X1 U4225 ( .A(n2867), .B(n2866), .Z(n7574) );
  CANR2XL U4226 ( .A(n7747), .B(n3137), .C(n7755), .D(n7574), .Z(n2873) );
  CANR2XL U4227 ( .A(n2995), .B(n3017), .C(n3173), .D(n2988), .Z(n2869) );
  CANR2XL U4228 ( .A(n3172), .B(n3019), .C(n3169), .D(n3018), .Z(n2868) );
  CND2X1 U4229 ( .A(n2869), .B(n2868), .Z(n7576) );
  CANR2XL U4230 ( .A(n2995), .B(n2996), .C(n3169), .D(n2993), .Z(n2871) );
  CANR2XL U4231 ( .A(n3173), .B(n2968), .C(n3172), .D(n2997), .Z(n2870) );
  CND2X1 U4232 ( .A(n2871), .B(n2870), .Z(n7575) );
  CANR2XL U4233 ( .A(n7582), .B(n7576), .C(n7762), .D(n7575), .Z(n2872) );
  CND2XL U4234 ( .A(n2873), .B(n2872), .Z(n7688) );
  CIVXL U4235 ( .A(acc[7]), .Z(n3885) );
  CANR2X1 U4236 ( .A(n2737), .B(out1_2[7]), .C(n2928), .D(out0_2[7]), .Z(n2874) );
  COND1XL U4237 ( .A(n2670), .B(n3885), .C(n2874), .Z(n3174) );
  CAOR2XL U4238 ( .A(out0_2[8]), .B(n2928), .C(n2737), .D(out1_2[8]), .Z(n2875) );
  CANR1XL U4239 ( .A(n2758), .B(acc[8]), .C(n2875), .Z(n3145) );
  CIVXL U4240 ( .A(acc[5]), .Z(n3879) );
  CANR2X1 U4241 ( .A(n2737), .B(out1_2[5]), .C(n2928), .D(out0_2[5]), .Z(n2876) );
  COND1XL U4242 ( .A(n2670), .B(n3879), .C(n2876), .Z(n7552) );
  CIVXL U4243 ( .A(acc[6]), .Z(n3882) );
  CANR2X1 U4244 ( .A(n2737), .B(out1_2[6]), .C(n2928), .D(out0_2[6]), .Z(n2877) );
  COND1XL U4245 ( .A(n2670), .B(n3882), .C(n2877), .Z(n3171) );
  CANR2XL U4246 ( .A(n3173), .B(n3098), .C(n3172), .D(n3130), .Z(n2879) );
  CANR2XL U4247 ( .A(n3169), .B(n3132), .C(n2995), .D(n3129), .Z(n2878) );
  CAN2X1 U4248 ( .A(n2879), .B(n2878), .Z(n7746) );
  CAOR2XL U4249 ( .A(out0_2[9]), .B(n2928), .C(n2737), .D(out1_2[9]), .Z(n2880) );
  CANR1XL U4250 ( .A(n2758), .B(acc[9]), .C(n2880), .Z(n3143) );
  CIVXL U4251 ( .A(n3143), .Z(n3045) );
  CND2XL U4252 ( .A(n3045), .B(n2995), .Z(n2882) );
  CANR2XL U4253 ( .A(n3173), .B(n3131), .C(n3172), .D(n3146), .Z(n2881) );
  COND3XL U4254 ( .A(n3144), .B(n7763), .C(n2882), .D(n2881), .Z(n7745) );
  CANR2XL U4255 ( .A(n3173), .B(n3013), .C(n3172), .D(n3103), .Z(n2884) );
  CANR2XL U4256 ( .A(n2995), .B(n3105), .C(n3169), .D(n3106), .Z(n2883) );
  CND2X1 U4257 ( .A(n2884), .B(n2883), .Z(n7580) );
  CANR2XL U4258 ( .A(n3173), .B(n3020), .C(n3172), .D(n3002), .Z(n2886) );
  CANR2XL U4259 ( .A(n2995), .B(n3004), .C(n3169), .D(n3005), .Z(n2885) );
  CND2X1 U4260 ( .A(n2886), .B(n2885), .Z(n7577) );
  CANR2XL U4261 ( .A(n3015), .B(n2995), .C(n3169), .D(n3012), .Z(n2888) );
  CANR2XL U4262 ( .A(n3173), .B(n3011), .C(n3172), .D(n3014), .Z(n2887) );
  CND2X1 U4263 ( .A(n2888), .B(n2887), .Z(n7584) );
  CANR2XL U4264 ( .A(n3173), .B(n3003), .C(n3172), .D(n3009), .Z(n2890) );
  CANR2XL U4265 ( .A(n2995), .B(n3008), .C(n3169), .D(n3010), .Z(n2889) );
  CND2X1 U4266 ( .A(n2890), .B(n2889), .Z(n7583) );
  CMX2XL U4267 ( .A0(n1232), .A1(h[3]), .S(pushin), .Z(n2893) );
  CANR2XL U4268 ( .A(n2995), .B(n3097), .C(n3169), .D(n3104), .Z(n2912) );
  CANR2XL U4269 ( .A(n3173), .B(n3106), .C(n3172), .D(n3105), .Z(n2911) );
  CND2X1 U4270 ( .A(n2912), .B(n2911), .Z(n4253) );
  CANR2XL U4271 ( .A(n7582), .B(n3078), .C(n7755), .D(n4253), .Z(n2918) );
  CANR2XL U4272 ( .A(n2995), .B(n3103), .C(n3169), .D(n3013), .Z(n2914) );
  CANR2XL U4273 ( .A(n3015), .B(n3172), .C(n3173), .D(n3012), .Z(n2913) );
  CND2X1 U4274 ( .A(n2914), .B(n2913), .Z(n4244) );
  CANR2XL U4275 ( .A(n3173), .B(n3010), .C(n3172), .D(n3008), .Z(n2916) );
  CANR2XL U4276 ( .A(n2995), .B(n3014), .C(n3169), .D(n3011), .Z(n2915) );
  CND2X1 U4277 ( .A(n2916), .B(n2915), .Z(n4243) );
  CANR2XL U4278 ( .A(n4244), .B(n2859), .C(n7747), .D(n4243), .Z(n2917) );
  CND2XL U4279 ( .A(n2918), .B(n2917), .Z(n4271) );
  CANR2XL U4280 ( .A(n4271), .B(n7543), .C(n2919), .D(n4240), .Z(n2937) );
  CANR2XL U4281 ( .A(n3173), .B(n3132), .C(n3172), .D(n3129), .Z(n2921) );
  CANR2XL U4282 ( .A(n2995), .B(n3146), .C(n3169), .D(n3131), .Z(n2920) );
  CND2X1 U4283 ( .A(n2921), .B(n2920), .Z(n3077) );
  CIVXL U4284 ( .A(acc[3]), .Z(n2955) );
  CANR2X1 U4285 ( .A(n2737), .B(out1_2[3]), .C(n2928), .D(out0_2[3]), .Z(n2922) );
  COND1XL U4286 ( .A(n2670), .B(n2955), .C(n2922), .Z(n7765) );
  CIVXL U4287 ( .A(acc[4]), .Z(n2961) );
  CANR2XL U4288 ( .A(n2995), .B(n7765), .C(n3169), .D(n7748), .Z(n2924) );
  CANR2XL U4289 ( .A(n3173), .B(n3171), .C(n3172), .D(n7552), .Z(n2923) );
  CND2XL U4290 ( .A(n2924), .B(n2923), .Z(n3190) );
  CANR2XL U4291 ( .A(n3192), .B(n3077), .C(n4249), .D(n3190), .Z(n2932) );
  CIVXL U4292 ( .A(out1_2[2]), .Z(n2926) );
  CANR2XL U4293 ( .A(n2671), .B(acc[2]), .C(n2928), .D(out0_2[2]), .Z(n2925)
         );
  COND1XL U4294 ( .A(n2927), .B(n2926), .C(n2925), .Z(n7769) );
  CAOR2XL U4295 ( .A(out0_2[0]), .B(n2928), .C(n2737), .D(out1_2[0]), .Z(n2929) );
  CANR1XL U4296 ( .A(n2758), .B(acc[0]), .C(n2929), .Z(n7767) );
  COND2XL U4297 ( .A(n7770), .B(n7749), .C(n7767), .D(n7763), .Z(n2930) );
  COND4CXL U4298 ( .A(n3173), .B(n7769), .C(n2930), .D(n4251), .Z(n2931) );
  COND3XL U4299 ( .A(n4252), .B(n3175), .C(n2932), .D(n2931), .Z(n2933) );
  CANR1XL U4300 ( .A(n4272), .B(n7699), .C(n2933), .Z(n2936) );
  CNR2X1 U4301 ( .A(n2934), .B(n7553), .Z(n7700) );
  CND3XL U4302 ( .A(n7700), .B(n3074), .C(h0_1[6]), .Z(n2935) );
  COND4CXL U4303 ( .A(n2937), .B(n2936), .C(h0_1[6]), .D(n2935), .Z(n2939) );
  CIVX12 U4304 ( .A(rst), .Z(n7935) );
  CND2X1 U4305 ( .A(n2865), .B(n7935), .Z(n2938) );
  CMX2XL U4306 ( .A0(n2939), .A1(roundit), .S(n2938), .Z(n2940) );
  CMX2XL U4307 ( .A0(q0[16]), .A1(q[16]), .S(n7682), .Z(n2942) );
  CMX2XL U4308 ( .A0(n2524), .A1(q[28]), .S(n7682), .Z(n2943) );
  CNIVX1 U4309 ( .A(out0_2[4]), .Z(n4378) );
  CIVXL U4310 ( .A(out2_2[4]), .Z(n3187) );
  CNIVX1 U4311 ( .A(out1_2[4]), .Z(n2947) );
  CIVX1 U4312 ( .A(n4292), .Z(n4353) );
  CNIVX1 U4313 ( .A(out0_2[33]), .Z(n2965) );
  CMX2XL U4314 ( .A0(q0[18]), .A1(q[18]), .S(n7682), .Z(n2946) );
  CND2X4 U4315 ( .A(n3883), .B(n2948), .Z(n7810) );
  CNR2IX2 U4316 ( .B(cmd0_en_2_d), .A(cmd1_en_2_d), .Z(n2950) );
  CNIVX4 U4317 ( .A(n2950), .Z(n4054) );
  CIVX1 U4318 ( .A(n3883), .Z(n4053) );
  CANR2XL U4319 ( .A(n4054), .B(out0_2[0]), .C(out1_2[0]), .D(n4053), .Z(n2949) );
  COND1XL U4320 ( .A(n8010), .B(n7810), .C(n2949), .Z(n2964) );
  CND2X1 U4321 ( .A(n2964), .B(out1_1[0]), .Z(n7845) );
  CNIVX4 U4322 ( .A(n2950), .Z(n7808) );
  CANR2XL U4323 ( .A(n7808), .B(out0_2[1]), .C(out1_2[1]), .D(n4053), .Z(n2951) );
  COND1XL U4324 ( .A(n8009), .B(n7810), .C(n2951), .Z(n2952) );
  CNR2XL U4325 ( .A(n2952), .B(out1_1[1]), .Z(n7843) );
  CND2X1 U4326 ( .A(n2952), .B(out1_1[1]), .Z(n7844) );
  COND1X1 U4327 ( .A(n7845), .B(n7843), .C(n7844), .Z(n2963) );
  CANR2XL U4328 ( .A(n4054), .B(out0_2[2]), .C(out1_2[2]), .D(n4053), .Z(n2953) );
  COND1XL U4329 ( .A(n8008), .B(n7810), .C(n2953), .Z(n2956) );
  CNR2XL U4330 ( .A(n2956), .B(out1_1[2]), .Z(n7840) );
  CANR2XL U4331 ( .A(n7808), .B(out0_2[3]), .C(out1_2[3]), .D(n4053), .Z(n2954) );
  COND1XL U4332 ( .A(n2955), .B(n7810), .C(n2954), .Z(n2957) );
  CNR2XL U4333 ( .A(n2957), .B(out1_1[3]), .Z(n7841) );
  CNR2XL U4334 ( .A(n7840), .B(n7841), .Z(n2959) );
  CND2XL U4335 ( .A(n2956), .B(out1_1[2]), .Z(n7838) );
  CND2XL U4336 ( .A(n2957), .B(out1_1[3]), .Z(n7842) );
  COND1XL U4337 ( .A(n7838), .B(n7841), .C(n7842), .Z(n2958) );
  CANR1X1 U4338 ( .A(n2963), .B(n2959), .C(n2958), .Z(n3892) );
  CIVX2 U4339 ( .A(n3892), .Z(n7788) );
  CANR2XL U4340 ( .A(n7808), .B(out0_2[4]), .C(out1_2[4]), .D(n4053), .Z(n2960) );
  COND1XL U4341 ( .A(n2961), .B(n7810), .C(n2960), .Z(n2962) );
  CNR2XL U4342 ( .A(n2962), .B(out1_1[4]), .Z(n3880) );
  CIVXL U4343 ( .A(n3880), .Z(n4239) );
  CND2X1 U4344 ( .A(n2962), .B(out1_1[4]), .Z(n4238) );
  CIVX1 U4345 ( .A(n2963), .Z(n7839) );
  CNIVX1 U4346 ( .A(out1_2[0]), .Z(n4362) );
  CMX2X1 U4347 ( .A0(n2965), .A1(out1_1[33]), .S(cmd0_en_2), .Z(n1151) );
  CMX2X1 U4348 ( .A0(n2966), .A1(out1_1[32]), .S(cmd0_en_2), .Z(n1152) );
  CNIVX1 U4349 ( .A(out0_2[24]), .Z(n3284) );
  CMX2X1 U4350 ( .A0(n3284), .A1(out1_1[24]), .S(cmd0_en_2), .Z(n1160) );
  CNIVX1 U4351 ( .A(out0_2[10]), .Z(n3311) );
  CMX2X1 U4352 ( .A0(n3311), .A1(out1_1[10]), .S(cmd0_en_2), .Z(n1174) );
  CNIVX1 U4353 ( .A(out0_2[9]), .Z(n3331) );
  CMX2X1 U4354 ( .A0(n3331), .A1(out1_1[9]), .S(cmd0_en_2), .Z(n1175) );
  CNIVX1 U4355 ( .A(out0_2[8]), .Z(n3338) );
  CMX2X1 U4356 ( .A0(n3338), .A1(out1_1[8]), .S(cmd0_en_2), .Z(n1176) );
  CNIVX1 U4357 ( .A(out0_2[2]), .Z(n3340) );
  CMX2X1 U4358 ( .A0(n3340), .A1(out1_1[2]), .S(cmd0_en_2), .Z(n1182) );
  CNIVX1 U4359 ( .A(out0_2[1]), .Z(n3205) );
  CMX2X1 U4360 ( .A0(n3205), .A1(out1_1[1]), .S(cmd0_en_2), .Z(n1183) );
  CMX2X1 U4361 ( .A0(n4361), .A1(out1_1[0]), .S(cmd0_en_2), .Z(n1184) );
  CMX2X1 U4362 ( .A0(h0_0[5]), .A1(h0[5]), .S(cmd2_en_0), .Z(n931) );
  CMX2X2 U4363 ( .A0(n1429), .A1(z[8]), .S(n7681), .Z(n1197) );
  CMX2X2 U4364 ( .A0(n1430), .A1(z[10]), .S(n7681), .Z(n1199) );
  CMX2X2 U4365 ( .A0(n1422), .A1(z[12]), .S(n7681), .Z(n1201) );
  CAOR2X2 U4366 ( .A(out2_2[57]), .B(n7751), .C(n7725), .D(n7738), .Z(n877) );
  CNIVX1 U4367 ( .A(cmd1_en_2), .Z(n8022) );
  CANR2XL U4368 ( .A(n2995), .B(n2968), .C(n3172), .D(n2967), .Z(n2972) );
  CANR2XL U4369 ( .A(n3173), .B(n2970), .C(n3169), .D(n2969), .Z(n2971) );
  CND2X1 U4370 ( .A(n2972), .B(n2971), .Z(n3182) );
  CANR2XL U4371 ( .A(n3182), .B(n7582), .C(n7747), .D(n3161), .Z(n2986) );
  CANR2XL U4372 ( .A(n2859), .B(n3160), .C(n7755), .D(n3159), .Z(n2985) );
  CND2X1 U4373 ( .A(n2986), .B(n2985), .Z(n7779) );
  CAOR2X2 U4374 ( .A(out2_2[48]), .B(n7751), .C(n7779), .D(n7738), .Z(n909) );
  CANR2X1 U4375 ( .A(n7582), .B(n3160), .C(n7755), .D(n3161), .Z(n7685) );
  CANR2XL U4376 ( .A(n2995), .B(n2988), .C(n3173), .D(n2987), .Z(n2992) );
  CANR2XL U4377 ( .A(n3172), .B(n2990), .C(n3169), .D(n2989), .Z(n2991) );
  CND2X1 U4378 ( .A(n2992), .B(n2991), .Z(n3179) );
  CANR2XL U4379 ( .A(n2995), .B(n2994), .C(n3172), .D(n2993), .Z(n2999) );
  CANR2XL U4380 ( .A(n3173), .B(n2997), .C(n3169), .D(n2996), .Z(n2998) );
  CND2X1 U4381 ( .A(n2999), .B(n2998), .Z(n3181) );
  CANR2XL U4382 ( .A(n7582), .B(n3179), .C(n7755), .D(n3181), .Z(n3001) );
  CANR2XL U4383 ( .A(n3182), .B(n2859), .C(n7747), .D(n3159), .Z(n3000) );
  CND2XL U4384 ( .A(n3001), .B(n3000), .Z(n3152) );
  CANR2XL U4385 ( .A(n2995), .B(n3003), .C(n3173), .D(n3002), .Z(n3007) );
  CANR2XL U4386 ( .A(n3172), .B(n3005), .C(n3169), .D(n3004), .Z(n3006) );
  CND2X1 U4387 ( .A(n3007), .B(n3006), .Z(n3165) );
  CAOR2XL U4388 ( .A(n7755), .B(n3164), .C(n3162), .D(n7582), .Z(n3016) );
  CANR1XL U4389 ( .A(n7762), .B(n3165), .C(n3016), .Z(n3155) );
  CANR2XL U4390 ( .A(n3172), .B(n3018), .C(n3169), .D(n3017), .Z(n3022) );
  CANR2XL U4391 ( .A(n2995), .B(n3020), .C(n3173), .D(n3019), .Z(n3021) );
  CND2X1 U4392 ( .A(n3022), .B(n3021), .Z(n3180) );
  CND2XL U4393 ( .A(n3180), .B(n7747), .Z(n3154) );
  CANR2XL U4394 ( .A(n4253), .B(n7582), .C(n7762), .D(n4243), .Z(n3025) );
  CANR2XL U4395 ( .A(n4244), .B(n7755), .C(n7747), .D(n4245), .Z(n3024) );
  CND2XL U4396 ( .A(n3025), .B(n3024), .Z(n3195) );
  CNR2XL U4397 ( .A(n3195), .B(n7729), .Z(n3032) );
  CANR2XL U4398 ( .A(n7582), .B(n4263), .C(n7755), .D(n3066), .Z(n3027) );
  CANR2XL U4399 ( .A(n3065), .B(n2859), .C(n7747), .D(n3064), .Z(n3026) );
  CND2X1 U4400 ( .A(n3027), .B(n3026), .Z(n7705) );
  CANR2XL U4401 ( .A(n7582), .B(n4246), .C(n7747), .D(n4262), .Z(n3029) );
  CANR2XL U4402 ( .A(n2859), .B(n4260), .C(n7755), .D(n4261), .Z(n3028) );
  CND2XL U4403 ( .A(n3029), .B(n3028), .Z(n7703) );
  COND2XL U4404 ( .A(n7724), .B(n7705), .C(n7727), .D(n7703), .Z(n3031) );
  CND2XL U4405 ( .A(n7751), .B(out2_2[19]), .Z(n3030) );
  CANR2XL U4406 ( .A(n7582), .B(n3035), .C(n7755), .D(n3034), .Z(n3036) );
  COAN1XL U4407 ( .A(n2662), .B(n3037), .C(n3036), .Z(n7741) );
  CANR2XL U4408 ( .A(n7582), .B(n3039), .C(n7755), .D(n3038), .Z(n3044) );
  CND2XL U4409 ( .A(n3040), .B(n7747), .Z(n3043) );
  CND2XL U4410 ( .A(n3041), .B(n2859), .Z(n3042) );
  CND3XL U4411 ( .A(n3044), .B(n3043), .C(n3042), .Z(n7739) );
  CANR2XL U4412 ( .A(n3045), .B(n3173), .C(n2995), .D(n3171), .Z(n3047) );
  CND2XL U4413 ( .A(n3174), .B(n3169), .Z(n3046) );
  COND3XL U4414 ( .A(n3145), .B(n7770), .C(n3047), .D(n3046), .Z(n7556) );
  CIVX1 U4415 ( .A(n4251), .Z(n3189) );
  CIVXL U4416 ( .A(n3048), .Z(n3049) );
  COND2XL U4417 ( .A(n3049), .B(n2662), .C(n3115), .D(n7553), .Z(n3050) );
  CANR1XL U4418 ( .A(n7755), .B(n3114), .C(n3050), .Z(n3054) );
  CND2XL U4419 ( .A(n3051), .B(n7747), .Z(n3053) );
  CND3XL U4420 ( .A(n3054), .B(n3074), .C(n3053), .Z(n3056) );
  COND3XL U4421 ( .A(n7727), .B(n7739), .C(n3056), .D(n3055), .Z(n3058) );
  CND2XL U4422 ( .A(out2_2[22]), .B(n7751), .Z(n3057) );
  COND4CXL U4423 ( .A(n7741), .B(n7771), .C(n3058), .D(n3057), .Z(n3059) );
  CND2X1 U4424 ( .A(n7724), .B(h0_1[4]), .Z(n7742) );
  CND2XL U4425 ( .A(n3152), .B(n7738), .Z(n3061) );
  CND2XL U4426 ( .A(out2_2[40]), .B(n7751), .Z(n3060) );
  COND3X2 U4427 ( .A(n7685), .B(n7742), .C(n3061), .D(n3060), .Z(n903) );
  CND2X1 U4428 ( .A(n3161), .B(n7582), .Z(n7683) );
  CND2XL U4429 ( .A(n3134), .B(n7738), .Z(n3063) );
  CND2XL U4430 ( .A(out2_2[44]), .B(n7751), .Z(n3062) );
  COND3X2 U4431 ( .A(n7683), .B(n7742), .C(n3063), .D(n3062), .Z(n907) );
  CANR2X1 U4432 ( .A(n3065), .B(n7582), .C(n7755), .D(n3064), .Z(n7684) );
  CANR2XL U4433 ( .A(n7582), .B(n4260), .C(n7747), .D(n3066), .Z(n3068) );
  CANR2XL U4434 ( .A(n2859), .B(n4263), .C(n7755), .D(n4262), .Z(n3067) );
  CND2XL U4435 ( .A(n3068), .B(n3067), .Z(n3085) );
  CMX2X2 U4436 ( .A0(n1425), .A1(z[24]), .S(n7681), .Z(n1213) );
  CIVXL U4437 ( .A(out2_2[28]), .Z(n4310) );
  CANR2XL U4438 ( .A(n7582), .B(n3164), .C(n7747), .D(n3179), .Z(n3070) );
  CANR2XL U4439 ( .A(n2859), .B(n3180), .C(n7755), .D(n3165), .Z(n3069) );
  CND2XL U4440 ( .A(n3070), .B(n3069), .Z(n3133) );
  CIVXL U4441 ( .A(n4246), .Z(n3073) );
  CANR2XL U4442 ( .A(n7582), .B(n4243), .C(n7755), .D(n4245), .Z(n3072) );
  COND1XL U4443 ( .A(n3073), .B(n2662), .C(n3072), .Z(n3084) );
  CND2XL U4444 ( .A(n4261), .B(n7747), .Z(n3082) );
  CIVX1 U4445 ( .A(n3077), .Z(n4250) );
  CIVX1 U4446 ( .A(n3078), .Z(n4256) );
  CANR2XL U4447 ( .A(n4251), .B(n4250), .C(n4249), .D(n4256), .Z(n3081) );
  CIVXL U4448 ( .A(n4244), .Z(n3079) );
  CANR1XL U4449 ( .A(n3192), .B(n3079), .C(h0_1[6]), .Z(n3080) );
  COND3XL U4450 ( .A(n3175), .B(n4253), .C(n3081), .D(n3080), .Z(n3087) );
  CND2XL U4451 ( .A(n3082), .B(n7543), .Z(n3083) );
  COND2XL U4452 ( .A(n4266), .B(n3085), .C(n3084), .D(n3083), .Z(n3086) );
  CANR3XL U4453 ( .A(n4272), .B(n7684), .C(n3087), .D(n3086), .Z(n3088) );
  CAOR1XL U4454 ( .A(out2_2[11]), .B(n7751), .C(n3088), .Z(n3089) );
  CMX2XL U4455 ( .A0(q0[8]), .A1(q[8]), .S(n7682), .Z(n3090) );
  COND2XL U4456 ( .A(n7727), .B(n7688), .C(n7729), .D(n3091), .Z(n3093) );
  CANR1XL U4457 ( .A(n7726), .B(n7689), .C(n7724), .Z(n3092) );
  CANR2XL U4458 ( .A(n2859), .B(n3179), .C(n7755), .D(n3180), .Z(n3096) );
  CANR2XL U4459 ( .A(n7582), .B(n3165), .C(n7747), .D(n3181), .Z(n3095) );
  CND2XL U4460 ( .A(n3096), .B(n3095), .Z(n7781) );
  CANR2XL U4461 ( .A(n2995), .B(n3098), .C(n3173), .D(n3097), .Z(n3102) );
  CANR2XL U4462 ( .A(n3172), .B(n3100), .C(n3169), .D(n3099), .Z(n3101) );
  CND2XL U4463 ( .A(n3102), .B(n3101), .Z(n3149) );
  CANR2XL U4464 ( .A(n3149), .B(n7582), .C(n7747), .D(n3164), .Z(n3110) );
  CANR2XL U4465 ( .A(n2995), .B(n3104), .C(n3173), .D(n3103), .Z(n3108) );
  CANR2XL U4466 ( .A(n3172), .B(n3106), .C(n3169), .D(n3105), .Z(n3107) );
  CND2X1 U4467 ( .A(n3108), .B(n3107), .Z(n3163) );
  CANR2XL U4468 ( .A(n3163), .B(n7755), .C(n7762), .D(n3162), .Z(n3109) );
  CND2XL U4469 ( .A(n3110), .B(n3109), .Z(n7777) );
  COND2XL U4470 ( .A(n7727), .B(n7781), .C(n7729), .D(n7777), .Z(n3112) );
  CANR1XL U4471 ( .A(n7726), .B(n7779), .C(n7724), .Z(n3111) );
  COND2X1 U4472 ( .A(n2865), .B(n8001), .C(n3112), .D(n3111), .Z(n891) );
  CIVX1 U4473 ( .A(out2_2[14]), .Z(n3219) );
  CIVXL U4474 ( .A(n3175), .Z(n4257) );
  CND2X1 U4475 ( .A(n3118), .B(n7582), .Z(n7675) );
  COND2XL U4476 ( .A(n3175), .B(n7580), .C(n3148), .D(n7581), .Z(n3119) );
  CANR1XL U4477 ( .A(n4272), .B(n7675), .C(n3119), .Z(n3121) );
  CANR1XL U4478 ( .A(n4251), .B(n7746), .C(h0_1[6]), .Z(n3120) );
  COND3XL U4479 ( .A(n4254), .B(n7584), .C(n3121), .D(n3120), .Z(n3128) );
  CANR2XL U4480 ( .A(n7575), .B(n7582), .C(n7747), .D(n3122), .Z(n3124) );
  CANR2XL U4481 ( .A(n3137), .B(n7755), .C(n2859), .D(n3136), .Z(n3123) );
  CND2XL U4482 ( .A(n3124), .B(n3123), .Z(n7540) );
  CANR2XL U4483 ( .A(n7747), .B(n7574), .C(n2859), .D(n7576), .Z(n3126) );
  CANR2XL U4484 ( .A(n7582), .B(n7583), .C(n7755), .D(n7577), .Z(n3125) );
  CND2XL U4485 ( .A(n3126), .B(n3125), .Z(n7542) );
  COND2XL U4486 ( .A(n4266), .B(n7540), .C(n7542), .D(n7727), .Z(n3127) );
  COND2X1 U4487 ( .A(n2865), .B(n8003), .C(n3128), .D(n3127), .Z(n867) );
  CIVXL U4488 ( .A(out2_2[12]), .Z(n3320) );
  CIVXL U4489 ( .A(n3149), .Z(n3168) );
  CANR2XL U4490 ( .A(n7582), .B(n7574), .C(n7755), .D(n7575), .Z(n3139) );
  CANR2XL U4491 ( .A(n3137), .B(n2859), .C(n7747), .D(n3136), .Z(n3138) );
  CND2X1 U4492 ( .A(n3139), .B(n3138), .Z(n7728) );
  CANR2XL U4493 ( .A(n7747), .B(n7576), .C(n7762), .D(n7577), .Z(n3141) );
  CANR2XL U4494 ( .A(n7582), .B(n7584), .C(n7755), .D(n7583), .Z(n3140) );
  CND2XL U4495 ( .A(n3141), .B(n3140), .Z(n7730) );
  CND2XL U4496 ( .A(n7761), .B(n4251), .Z(n3147) );
  COND3XL U4497 ( .A(n4254), .B(n3163), .C(n3147), .D(n8019), .Z(n3151) );
  COND2XL U4498 ( .A(n3175), .B(n3149), .C(n3148), .D(n7759), .Z(n3150) );
  CANR3XL U4499 ( .A(n4272), .B(n7685), .C(n3151), .D(n3150), .Z(n3157) );
  CNR2XL U4500 ( .A(n3152), .B(n4266), .Z(n3153) );
  CANR11XL U4501 ( .A(n3155), .B(n7543), .C(n3154), .D(n3153), .Z(n3156) );
  CAOR2XL U4502 ( .A(out2_2[8]), .B(n7751), .C(n3157), .D(n3156), .Z(n3158) );
  CAOR2X2 U4503 ( .A(out2_2[52]), .B(n7751), .C(n7712), .D(n7738), .Z(n908) );
  CANR2XL U4504 ( .A(n3163), .B(n7582), .C(n7755), .D(n3162), .Z(n3167) );
  CANR2XL U4505 ( .A(n7747), .B(n3165), .C(n7762), .D(n3164), .Z(n3166) );
  CND2XL U4506 ( .A(n3167), .B(n3166), .Z(n7544) );
  CANR2XL U4507 ( .A(n7761), .B(n4249), .C(n3192), .D(n3168), .Z(n3178) );
  CAOR2XL U4508 ( .A(n2995), .B(n7748), .C(n3169), .D(n7552), .Z(n3170) );
  CANR1XL U4509 ( .A(n3172), .B(n3171), .C(n3170), .Z(n7756) );
  CND2XL U4510 ( .A(n3174), .B(n3173), .Z(n7754) );
  COND1XL U4511 ( .A(n3175), .B(n7759), .C(n8019), .Z(n3176) );
  CANR11XL U4512 ( .A(n4251), .B(n7756), .C(n7754), .D(n3176), .Z(n3177) );
  COND3XL U4513 ( .A(n7727), .B(n7544), .C(n3178), .D(n3177), .Z(n3186) );
  CANR2XL U4514 ( .A(n7582), .B(n3180), .C(n7755), .D(n3179), .Z(n3184) );
  CANR2XL U4515 ( .A(n7747), .B(n3182), .C(n7762), .D(n3181), .Z(n3183) );
  CND2XL U4516 ( .A(n3184), .B(n3183), .Z(n7713) );
  COND2XL U4517 ( .A(n4267), .B(n7712), .C(n7713), .D(n4266), .Z(n3185) );
  COND2X1 U4518 ( .A(n2865), .B(n3187), .C(n3186), .D(n3185), .Z(n3188) );
  CANR2XL U4519 ( .A(n4252), .B(n4249), .C(n4257), .D(n4250), .Z(n3194) );
  CNR2XL U4520 ( .A(n3190), .B(n3189), .Z(n3191) );
  CANR3XL U4521 ( .A(n3192), .B(n4256), .C(n3191), .D(h0_1[6]), .Z(n3193) );
  COND3XL U4522 ( .A(n7727), .B(n3195), .C(n3194), .D(n3193), .Z(n3197) );
  COND2XL U4523 ( .A(n4267), .B(n7705), .C(n4266), .D(n7703), .Z(n3196) );
  COND2XL U4524 ( .A(n2865), .B(n3198), .C(n3197), .D(n3196), .Z(n3199) );
  CMX2XL U4525 ( .A0(q0[30]), .A1(q[30]), .S(n7682), .Z(n3200) );
  CIVX2 U4526 ( .A(n3200), .Z(n7856) );
  CIVX8 U4527 ( .A(q0[0]), .Z(n7537) );
  CND2X4 U4528 ( .A(n3580), .B(n7537), .Z(n5160) );
  CNIVX1 U4529 ( .A(n3580), .Z(n3210) );
  CENX1 U4530 ( .A(n3210), .B(h0[2]), .Z(n3698) );
  COND2X1 U4531 ( .A(n5160), .B(n3203), .C(n7537), .D(n3698), .Z(n3202) );
  CNIVX4 U4532 ( .A(n4492), .Z(n4886) );
  CNR2IX1 U4533 ( .B(n7539), .A(n4886), .Z(n3201) );
  COR2X1 U4534 ( .A(n3202), .B(n3201), .Z(n3695) );
  CND2X1 U4535 ( .A(n3202), .B(n3201), .Z(n3694) );
  CND2X1 U4536 ( .A(n3695), .B(n3694), .Z(n3204) );
  COND2XL U4537 ( .A(n5160), .B(n7539), .C(n7537), .D(n3203), .Z(n6371) );
  CIVX8 U4538 ( .A(n2624), .Z(n5106) );
  CNIVX4 U4539 ( .A(n5106), .Z(n3631) );
  CND2X1 U4540 ( .A(n6371), .B(n6370), .Z(n6372) );
  CIVX1 U4541 ( .A(n6372), .Z(n3696) );
  CENX1 U4542 ( .A(n3204), .B(n3696), .Z(N17) );
  CIVXL U4543 ( .A(n3205), .Z(n3209) );
  CIVXL U4544 ( .A(out2_2[1]), .Z(n3341) );
  CEOXL U4545 ( .A(n4364), .B(n3341), .Z(n3206) );
  CND2XL U4546 ( .A(n3206), .B(n4344), .Z(n3208) );
  CNIVX1 U4547 ( .A(out1_2[1]), .Z(n7847) );
  CANR2X1 U4548 ( .A(n4363), .B(n7847), .C(acc[1]), .D(n4350), .Z(n3207) );
  COND3XL U4549 ( .A(n3209), .B(n2685), .C(n3208), .D(n3207), .Z(n994) );
  CNIVX4 U4550 ( .A(n3345), .Z(n3463) );
  CIVX8 U4551 ( .A(n3463), .Z(n6491) );
  CIVX2 U4552 ( .A(n7858), .Z(n4922) );
  CMX2XL U4553 ( .A0(q0[2]), .A1(q[2]), .S(n7682), .Z(n3212) );
  CIVXL U4554 ( .A(n3212), .Z(n7855) );
  CIVX1 U4555 ( .A(n3295), .Z(n3305) );
  CIVXL U4556 ( .A(out2_2[19]), .Z(n3306) );
  CNR2X1 U4557 ( .A(n3305), .B(n3306), .Z(n3214) );
  CENX1 U4558 ( .A(n3214), .B(n7999), .Z(n3215) );
  CND2XL U4559 ( .A(n3215), .B(n4344), .Z(n3217) );
  CANR2XL U4560 ( .A(n4363), .B(out1_2[20]), .C(acc[20]), .D(n4350), .Z(n3216)
         );
  COND3XL U4561 ( .A(n2685), .B(n2630), .C(n3217), .D(n3216), .Z(n1013) );
  CNIVX1 U4562 ( .A(out0_2[14]), .Z(n4381) );
  CIVXL U4563 ( .A(n1376), .Z(n3224) );
  CNR2X1 U4564 ( .A(n3218), .B(n8003), .Z(n3220) );
  CENX1 U4565 ( .A(n3220), .B(n3219), .Z(n3221) );
  CND2XL U4566 ( .A(n3221), .B(n4344), .Z(n3223) );
  CANR2XL U4567 ( .A(n4363), .B(out1_2[14]), .C(acc[14]), .D(n4350), .Z(n3222)
         );
  COND3XL U4568 ( .A(n2685), .B(n3224), .C(n3223), .D(n3222), .Z(n1007) );
  CNIVX1 U4569 ( .A(out0_2[40]), .Z(n7679) );
  CIVXL U4570 ( .A(n1369), .Z(n3230) );
  CNR2X1 U4571 ( .A(n4292), .B(n3225), .Z(n3232) );
  CIVX1 U4572 ( .A(n3232), .Z(n3275) );
  CNR2X1 U4573 ( .A(n3275), .B(n7979), .Z(n3226) );
  CENX1 U4574 ( .A(n3226), .B(n7978), .Z(n3227) );
  CND2XL U4575 ( .A(n3227), .B(n4344), .Z(n3229) );
  CANR2XL U4576 ( .A(n4363), .B(out1_2[40]), .C(acc[40]), .D(n4350), .Z(n3228)
         );
  COND3XL U4577 ( .A(n2685), .B(n3230), .C(n3229), .D(n3228), .Z(n1033) );
  CNR2X1 U4578 ( .A(n4328), .B(n7977), .Z(n3233) );
  CENX1 U4579 ( .A(n3233), .B(n7975), .Z(n3234) );
  CND2XL U4580 ( .A(n3234), .B(n4344), .Z(n3236) );
  CANR2XL U4581 ( .A(n4363), .B(out1_2[42]), .C(acc[42]), .D(n4350), .Z(n3235)
         );
  CNR2X1 U4582 ( .A(n3237), .B(n7970), .Z(n3238) );
  CENX1 U4583 ( .A(n3238), .B(n7969), .Z(n3239) );
  CND2XL U4584 ( .A(n3239), .B(n4344), .Z(n3241) );
  CANR2XL U4585 ( .A(n4363), .B(out1_2[46]), .C(acc[46]), .D(n4350), .Z(n3240)
         );
  CIVX1 U4586 ( .A(n3248), .Z(n4338) );
  CNR2X1 U4587 ( .A(n4338), .B(n7968), .Z(n3243) );
  CENX1 U4588 ( .A(n3243), .B(n7967), .Z(n3244) );
  CND2XL U4589 ( .A(n3244), .B(n4344), .Z(n3246) );
  CANR2XL U4590 ( .A(n4363), .B(out1_2[48]), .C(acc[48]), .D(n4350), .Z(n3245)
         );
  COND3XL U4591 ( .A(n2685), .B(n2633), .C(n3246), .D(n3245), .Z(n1041) );
  CNR2X1 U4592 ( .A(n3286), .B(n7965), .Z(n3249) );
  CENX1 U4593 ( .A(n3249), .B(n7963), .Z(n3250) );
  CND2XL U4594 ( .A(n3250), .B(n4344), .Z(n3252) );
  CANR2XL U4595 ( .A(n4363), .B(out1_2[50]), .C(acc[50]), .D(n4350), .Z(n3251)
         );
  COND3XL U4596 ( .A(n2685), .B(n2634), .C(n3252), .D(n3251), .Z(n1043) );
  CIVX1 U4597 ( .A(n3253), .Z(n4348) );
  CNR2X1 U4598 ( .A(n4348), .B(n7961), .Z(n3254) );
  CENX1 U4599 ( .A(n3254), .B(n7959), .Z(n3255) );
  CND2XL U4600 ( .A(n3255), .B(n4344), .Z(n3257) );
  CANR2XL U4601 ( .A(n4363), .B(out1_2[52]), .C(acc[52]), .D(n4350), .Z(n3256)
         );
  CEOXL U4602 ( .A(n7949), .B(n3258), .Z(n3259) );
  CND2XL U4603 ( .A(n3259), .B(n4344), .Z(n3261) );
  CANR2XL U4604 ( .A(n4363), .B(out1_2[57]), .C(acc[57]), .D(n4350), .Z(n3260)
         );
  CND2X1 U4605 ( .A(n4281), .B(n3262), .Z(n4318) );
  CEOXL U4606 ( .A(n7945), .B(n4318), .Z(n3263) );
  CND2XL U4607 ( .A(n3263), .B(n4344), .Z(n3265) );
  CANR2XL U4608 ( .A(n4363), .B(out1_2[59]), .C(acc[59]), .D(n8004), .Z(n3264)
         );
  CHA1XL U4609 ( .A(out2_2[62]), .B(n3266), .CO(n2721), .S(n3267) );
  CNIVX1 U4610 ( .A(out0_2[27]), .Z(n4370) );
  CIVXL U4611 ( .A(n1372), .Z(n3274) );
  CIVXL U4612 ( .A(out2_2[27]), .Z(n4308) );
  CIVX1 U4613 ( .A(n4316), .Z(n4309) );
  CEOXL U4614 ( .A(n4308), .B(n4309), .Z(n3271) );
  CND2XL U4615 ( .A(n3271), .B(n4344), .Z(n3273) );
  CANR2XL U4616 ( .A(n4363), .B(out1_2[27]), .C(acc[27]), .D(n4350), .Z(n3272)
         );
  COND3XL U4617 ( .A(n3274), .B(n2685), .C(n3273), .D(n3272), .Z(n1020) );
  CEOXL U4618 ( .A(n7979), .B(n3275), .Z(n3276) );
  CND2XL U4619 ( .A(n3276), .B(n4344), .Z(n3278) );
  CANR2XL U4620 ( .A(n4363), .B(out1_2[39]), .C(acc[39]), .D(n4350), .Z(n3277)
         );
  CNIVX1 U4621 ( .A(out0_2[43]), .Z(n4386) );
  CIVXL U4622 ( .A(n1367), .Z(n3283) );
  CIVX1 U4623 ( .A(n3279), .Z(n4303) );
  CEOXL U4624 ( .A(n7974), .B(n4303), .Z(n3280) );
  CND2XL U4625 ( .A(n3280), .B(n4344), .Z(n3282) );
  CANR2XL U4626 ( .A(n4363), .B(out1_2[43]), .C(acc[43]), .D(n4350), .Z(n3281)
         );
  COND3XL U4627 ( .A(n2685), .B(n3283), .C(n3282), .D(n3281), .Z(n1036) );
  CIVX2 U4628 ( .A(n3285), .Z(n3326) );
  CEOXL U4629 ( .A(n7965), .B(n3286), .Z(n3287) );
  CND2XL U4630 ( .A(n3287), .B(n4344), .Z(n3289) );
  CANR2XL U4631 ( .A(n4363), .B(out1_2[49]), .C(acc[49]), .D(n4350), .Z(n3288)
         );
  CEOXL U4632 ( .A(n7957), .B(n3290), .Z(n3291) );
  CND2XL U4633 ( .A(n3291), .B(n4344), .Z(n3293) );
  CANR2XL U4634 ( .A(n4363), .B(out1_2[53]), .C(acc[53]), .D(n4350), .Z(n3292)
         );
  COND3XL U4635 ( .A(n2685), .B(n2640), .C(n3293), .D(n3292), .Z(n1046) );
  CEOXL U4636 ( .A(n4279), .B(n4280), .Z(n3296) );
  CND2XL U4637 ( .A(n3296), .B(n4344), .Z(n3298) );
  CANR2XL U4638 ( .A(n4363), .B(out1_2[21]), .C(acc[21]), .D(n4350), .Z(n3297)
         );
  COND3XL U4639 ( .A(n2651), .B(n2685), .C(n3298), .D(n3297), .Z(n1014) );
  CNR2X1 U4640 ( .A(n3321), .B(n3299), .Z(n3322) );
  CNIVX1 U4641 ( .A(out0_2[25]), .Z(n4372) );
  CIVXL U4642 ( .A(n1377), .Z(n3304) );
  CEOXL U4643 ( .A(n7997), .B(n4317), .Z(n3301) );
  CND2XL U4644 ( .A(n3301), .B(n4344), .Z(n3303) );
  CANR2XL U4645 ( .A(n4363), .B(out1_2[25]), .C(acc[25]), .D(n4350), .Z(n3302)
         );
  COND3XL U4646 ( .A(n3304), .B(n2685), .C(n3303), .D(n3302), .Z(n1018) );
  CNIVX1 U4647 ( .A(out0_2[19]), .Z(n4374) );
  CIVXL U4648 ( .A(n1374), .Z(n3310) );
  CEOXL U4649 ( .A(n3306), .B(n3305), .Z(n3307) );
  CND2XL U4650 ( .A(n3307), .B(n4344), .Z(n3309) );
  CANR2XL U4651 ( .A(n4363), .B(out1_2[19]), .C(acc[19]), .D(n4350), .Z(n3308)
         );
  COND3XL U4652 ( .A(n3310), .B(n2685), .C(n3309), .D(n3308), .Z(n1012) );
  CNIVX1 U4653 ( .A(out0_2[11]), .Z(n4384) );
  CIVXL U4654 ( .A(n4384), .Z(n3317) );
  CIVXL U4655 ( .A(out2_2[11]), .Z(n3318) );
  CENX1 U4656 ( .A(n3313), .B(n3318), .Z(n3314) );
  CND2XL U4657 ( .A(n3314), .B(n4344), .Z(n3316) );
  CANR2XL U4658 ( .A(n4363), .B(out1_2[11]), .C(n1421), .D(n4350), .Z(n3315)
         );
  COND3XL U4659 ( .A(n3317), .B(n2685), .C(n3316), .D(n3315), .Z(n1004) );
  CNIVX1 U4660 ( .A(out0_2[12]), .Z(n4383) );
  CENX1 U4661 ( .A(n3322), .B(n8000), .Z(n3323) );
  CND2XL U4662 ( .A(n3323), .B(n4344), .Z(n3325) );
  CANR2XL U4663 ( .A(n4363), .B(out1_2[17]), .C(acc[17]), .D(n4350), .Z(n3324)
         );
  CNIVX1 U4664 ( .A(out0_2[23]), .Z(n4373) );
  CIVXL U4665 ( .A(n1388), .Z(n3330) );
  CENX1 U4666 ( .A(n3326), .B(n7998), .Z(n3327) );
  CND2XL U4667 ( .A(n3327), .B(n4344), .Z(n3329) );
  CANR2XL U4668 ( .A(n4363), .B(out1_2[23]), .C(acc[23]), .D(n4350), .Z(n3328)
         );
  COND3XL U4669 ( .A(n3330), .B(n2685), .C(n3329), .D(n3328), .Z(n1016) );
  CIVXL U4670 ( .A(n3331), .Z(n3337) );
  CEOXL U4671 ( .A(n3333), .B(n3332), .Z(n3334) );
  CND2XL U4672 ( .A(n3334), .B(n4344), .Z(n3336) );
  CANR2XL U4673 ( .A(n4363), .B(out1_2[9]), .C(n1420), .D(n4350), .Z(n3335) );
  COND3XL U4674 ( .A(n3337), .B(n2685), .C(n3336), .D(n3335), .Z(n1002) );
  CMX2XL U4675 ( .A0(n5927), .A1(h[9]), .S(n7682), .Z(n938) );
  CIVX4 U4676 ( .A(n7863), .Z(n5701) );
  CDLY1XL U4677 ( .A(n2341), .Z(n3342) );
  CMX2XL U4678 ( .A0(n3342), .A1(q[12]), .S(n7682), .Z(n973) );
  CMX2XL U4679 ( .A0(h0[30]), .A1(h[30]), .S(n7682), .Z(n959) );
  CIVX2 U4680 ( .A(q0[13]), .Z(n3345) );
  CIVX2 U4681 ( .A(q0[12]), .Z(n3344) );
  CND2X4 U4682 ( .A(n3347), .B(n3346), .Z(n6576) );
  CENX1 U4683 ( .A(n6491), .B(n2512), .Z(n3391) );
  CENX2 U4684 ( .A(q0[11]), .B(q0[12]), .Z(n3459) );
  CENX1 U4685 ( .A(n5888), .B(h0[5]), .Z(n3402) );
  CENX2 U4686 ( .A(q0[15]), .B(n7859), .Z(n3348) );
  CND2X4 U4687 ( .A(n3348), .B(n2540), .Z(n6703) );
  CIVX8 U4688 ( .A(n7861), .Z(n6647) );
  CENX1 U4689 ( .A(n6647), .B(h0[2]), .Z(n3388) );
  CENX2 U4690 ( .A(q0[11]), .B(n7868), .Z(n3449) );
  CND2X2 U4691 ( .A(n3449), .B(n2369), .Z(n6418) );
  CIVX12 U4692 ( .A(n7872), .Z(n6417) );
  CNIVX4 U4693 ( .A(h0[6]), .Z(n7674) );
  CENX1 U4694 ( .A(n6417), .B(n7674), .Z(n3386) );
  CNIVX4 U4695 ( .A(n3578), .Z(n6293) );
  CENX1 U4696 ( .A(n6417), .B(h0[7]), .Z(n3349) );
  CND2X2 U4697 ( .A(n3578), .B(n3449), .Z(n6211) );
  CNIVX4 U4698 ( .A(n2369), .Z(n6523) );
  CENX1 U4699 ( .A(n6417), .B(h0[8]), .Z(n3775) );
  COND2X1 U4700 ( .A(n3349), .B(n6211), .C(n6523), .D(n3775), .Z(n3772) );
  CIVX4 U4701 ( .A(n7863), .Z(n5793) );
  CENX1 U4702 ( .A(h0[13]), .B(n5793), .Z(n3404) );
  CNIVX16 U4703 ( .A(n3350), .Z(n5912) );
  CENX1 U4704 ( .A(h0[14]), .B(n5793), .Z(n3774) );
  COND2X1 U4705 ( .A(n5911), .B(n3404), .C(n5912), .D(n3774), .Z(n3771) );
  CNR2X2 U4706 ( .A(q0[8]), .B(q0[7]), .Z(n3353) );
  CND2X2 U4707 ( .A(q0[8]), .B(q0[7]), .Z(n3354) );
  CND2X2 U4708 ( .A(n3354), .B(n7858), .Z(n3351) );
  COND1X2 U4709 ( .A(n3615), .B(n3353), .C(n3351), .Z(n3352) );
  CENX1 U4710 ( .A(n6118), .B(n5927), .Z(n3372) );
  CIVX2 U4711 ( .A(n3353), .Z(n3355) );
  CND2X2 U4712 ( .A(n3355), .B(n3354), .Z(n4737) );
  CENX1 U4713 ( .A(n6191), .B(h0[10]), .Z(n3786) );
  COND2X1 U4714 ( .A(n2515), .B(n3787), .C(n6473), .D(n3356), .Z(n3765) );
  CNIVX4 U4715 ( .A(h0[0]), .Z(n7538) );
  CIVX2 U4716 ( .A(q0[18]), .Z(n3357) );
  CND2X2 U4717 ( .A(n3357), .B(n7865), .Z(n3754) );
  CND2X2 U4718 ( .A(q0[18]), .B(n7860), .Z(n4419) );
  CND2X2 U4719 ( .A(n3754), .B(n4419), .Z(n6871) );
  CNIVX4 U4720 ( .A(n6871), .Z(n6770) );
  CNR2IX1 U4721 ( .B(n7538), .A(n6770), .Z(n3766) );
  CENX1 U4722 ( .A(n5106), .B(h0[17]), .Z(n3373) );
  CENX1 U4723 ( .A(n5106), .B(h0[18]), .Z(n3778) );
  COND2X2 U4724 ( .A(n5160), .B(n3373), .C(n7537), .D(n3778), .Z(n3767) );
  CENX1 U4725 ( .A(n3765), .B(n3358), .Z(n3781) );
  CEO3X2 U4726 ( .A(n3782), .B(n3780), .C(n3781), .Z(n3796) );
  CND2IX1 U4727 ( .B(n7539), .A(n6647), .Z(n3360) );
  COND2X1 U4728 ( .A(n7861), .B(n6703), .C(n3360), .D(n2514), .Z(n3446) );
  CENX1 U4729 ( .A(n6647), .B(h0[1]), .Z(n3389) );
  COND2X1 U4730 ( .A(n6703), .B(n3361), .C(n2514), .D(n3389), .Z(n3445) );
  CENX1 U4731 ( .A(n6191), .B(n7674), .Z(n3453) );
  CENX1 U4732 ( .A(n6191), .B(h0[7]), .Z(n3397) );
  COND2X1 U4733 ( .A(n2577), .B(n3453), .C(n2490), .D(n3397), .Z(n3457) );
  CENX1 U4734 ( .A(n5793), .B(h0[10]), .Z(n3465) );
  CENX1 U4735 ( .A(n5793), .B(h0[11]), .Z(n3394) );
  COND2X1 U4736 ( .A(n5911), .B(n3465), .C(n5912), .D(n3394), .Z(n3456) );
  CENX1 U4737 ( .A(n5106), .B(h0[14]), .Z(n3448) );
  CIVX4 U4738 ( .A(n2624), .Z(n4861) );
  CENX1 U4739 ( .A(n4861), .B(h0[15]), .Z(n3393) );
  COND2X1 U4740 ( .A(n5160), .B(n3448), .C(n7537), .D(n3393), .Z(n3455) );
  COND1X1 U4741 ( .A(n3457), .B(n3456), .C(n3455), .Z(n3363) );
  CND2X1 U4742 ( .A(n3457), .B(n3456), .Z(n3362) );
  CND2X2 U4743 ( .A(n3363), .B(n3362), .Z(n3442) );
  CENX1 U4744 ( .A(n6491), .B(h0[2]), .Z(n3452) );
  CENX1 U4745 ( .A(n6491), .B(h0[3]), .Z(n3390) );
  COND2X1 U4746 ( .A(n2449), .B(n3452), .C(n1557), .D(n3390), .Z(n3486) );
  CNR2X2 U4747 ( .A(q0[6]), .B(q0[5]), .Z(n3365) );
  CND2X2 U4748 ( .A(q0[6]), .B(q0[5]), .Z(n3366) );
  COND1X4 U4749 ( .A(n3643), .B(n3365), .C(n3364), .Z(n6114) );
  CENX1 U4750 ( .A(h0[8]), .B(n5923), .Z(n3464) );
  CIVX2 U4751 ( .A(n3365), .Z(n3367) );
  CENX1 U4752 ( .A(n5927), .B(n5923), .Z(n3395) );
  COND2X1 U4753 ( .A(n6114), .B(n3464), .C(n3368), .D(n3395), .Z(n3485) );
  CENX1 U4754 ( .A(n6417), .B(n2513), .Z(n3450) );
  CENX1 U4755 ( .A(n6417), .B(h0[5]), .Z(n3387) );
  COND2X1 U4756 ( .A(n6418), .B(n3450), .C(n6523), .D(n3387), .Z(n3484) );
  COND1X1 U4757 ( .A(n3443), .B(n3442), .C(n3441), .Z(n3370) );
  CND2X1 U4758 ( .A(n3442), .B(n3443), .Z(n3369) );
  CND2X2 U4759 ( .A(n3370), .B(n3369), .Z(n3431) );
  CENX1 U4760 ( .A(h0[14]), .B(n5104), .Z(n3385) );
  CND2X4 U4761 ( .A(n4492), .B(n3371), .Z(n5695) );
  CENX1 U4762 ( .A(h0[15]), .B(n2531), .Z(n3400) );
  COND2X1 U4763 ( .A(n3385), .B(n5695), .C(n4886), .D(n3400), .Z(n3378) );
  CENX1 U4764 ( .A(n6118), .B(h0[8]), .Z(n3396) );
  COND2X1 U4765 ( .A(n2562), .B(n3396), .C(n2488), .D(n3372), .Z(n3377) );
  CENX1 U4766 ( .A(n5106), .B(h0[16]), .Z(n3392) );
  COND2X1 U4767 ( .A(n5160), .B(n3392), .C(n7537), .D(n3373), .Z(n3376) );
  COND1X2 U4768 ( .A(n3433), .B(n3431), .C(n3432), .Z(n3375) );
  CND2X2 U4769 ( .A(n3375), .B(n3374), .Z(n3794) );
  CNIVX4 U4770 ( .A(n6114), .Z(n4959) );
  CENX1 U4771 ( .A(h0[11]), .B(n5923), .Z(n3408) );
  CNIVX4 U4772 ( .A(n3368), .Z(n4957) );
  CENX1 U4773 ( .A(n5923), .B(h0[12]), .Z(n3777) );
  COND2X1 U4774 ( .A(n4959), .B(n3408), .C(n4957), .D(n3777), .Z(n3792) );
  CFA1X1 U4775 ( .A(n3378), .B(n3377), .CI(n3376), .CO(n3791), .S(n3432) );
  CND2XL U4776 ( .A(n4399), .B(n6409), .Z(n3381) );
  CIVXL U4777 ( .A(n6409), .Z(n4365) );
  CIVX4 U4778 ( .A(n2584), .Z(n3788) );
  CND2IXL U4779 ( .B(n4365), .A(n3788), .Z(n3380) );
  COND1XL U4780 ( .A(n2436), .B(n3381), .C(n3380), .Z(n3407) );
  CENX1 U4781 ( .A(n6409), .B(h0[1]), .Z(n3401) );
  CNIVX4 U4782 ( .A(n7860), .Z(n6699) );
  CENX1 U4783 ( .A(n7538), .B(n6699), .Z(n3383) );
  COND2X2 U4784 ( .A(n6765), .B(n3401), .C(n3383), .D(n1582), .Z(n3406) );
  CENX2 U4785 ( .A(n3794), .B(n3795), .Z(n3384) );
  CENX2 U4786 ( .A(n1545), .B(n3384), .Z(n3802) );
  CENX1 U4787 ( .A(h0[13]), .B(n5566), .Z(n3444) );
  CNIVX4 U4788 ( .A(n4492), .Z(n5696) );
  COND2X1 U4789 ( .A(n5695), .B(n3444), .C(n5696), .D(n3385), .Z(n3413) );
  COND2X1 U4790 ( .A(n6211), .B(n3387), .C(n6293), .D(n3386), .Z(n3412) );
  COND2X1 U4791 ( .A(n6703), .B(n3389), .C(n2515), .D(n3388), .Z(n3411) );
  CNR2IX1 U4792 ( .B(n7539), .A(n6765), .Z(n3416) );
  COND2X1 U4793 ( .A(n1557), .B(n3391), .C(n3390), .D(n2449), .Z(n3415) );
  COND2X1 U4794 ( .A(n5160), .B(n3393), .C(n7537), .D(n3392), .Z(n3414) );
  CENX1 U4795 ( .A(h0[12]), .B(n5793), .Z(n3405) );
  COND2X1 U4796 ( .A(n5911), .B(n3394), .C(n5912), .D(n3405), .Z(n3419) );
  CENX1 U4797 ( .A(h0[10]), .B(n5923), .Z(n3409) );
  COND2X1 U4798 ( .A(n6114), .B(n3395), .C(n3368), .D(n3409), .Z(n3418) );
  COND2X1 U4799 ( .A(n2567), .B(n3397), .C(n2489), .D(n3396), .Z(n3417) );
  COND1X1 U4800 ( .A(n3425), .B(n3426), .C(n3427), .Z(n3399) );
  CND2X1 U4801 ( .A(n3425), .B(n3426), .Z(n3398) );
  CND2X2 U4802 ( .A(n3399), .B(n3398), .Z(n3751) );
  CENX1 U4803 ( .A(h0[16]), .B(n5566), .Z(n3773) );
  COND2X1 U4804 ( .A(n5695), .B(n3400), .C(n5696), .D(n3773), .Z(n3762) );
  CENX1 U4805 ( .A(n6409), .B(h0[2]), .Z(n3789) );
  CENX1 U4806 ( .A(n6491), .B(n7674), .Z(n3776) );
  COND2X1 U4807 ( .A(n2449), .B(n3402), .C(n1556), .D(n3776), .Z(n3761) );
  CENX1 U4808 ( .A(n3760), .B(n3761), .Z(n3403) );
  CENX2 U4809 ( .A(n3762), .B(n3403), .Z(n3750) );
  COND2X1 U4810 ( .A(n4443), .B(n3405), .C(n5912), .D(n3404), .Z(n3424) );
  CHA1X1 U4811 ( .A(n3407), .B(n3406), .CO(n3790), .S(n3423) );
  COND2X1 U4812 ( .A(n4959), .B(n3409), .C(n4957), .D(n3408), .Z(n3422) );
  CENX2 U4813 ( .A(n3750), .B(n3749), .Z(n3410) );
  CENX2 U4814 ( .A(n3751), .B(n3410), .Z(n3801) );
  CFA1X1 U4815 ( .A(n3413), .B(n3412), .CI(n3411), .CO(n3425), .S(n3533) );
  CFA1X1 U4816 ( .A(n3416), .B(n3415), .CI(n3414), .CO(n3426), .S(n3535) );
  CFA1X1 U4817 ( .A(n3419), .B(n3418), .CI(n3417), .CO(n3427), .S(n3532) );
  CND2X1 U4818 ( .A(n3535), .B(n3533), .Z(n3420) );
  CND2X2 U4819 ( .A(n3421), .B(n3420), .Z(n3440) );
  CFA1X1 U4820 ( .A(n3424), .B(n3423), .CI(n3422), .CO(n3749), .S(n3437) );
  CND2X2 U4821 ( .A(n3429), .B(n3428), .Z(n3800) );
  CENX2 U4822 ( .A(n3801), .B(n3800), .Z(n3430) );
  CIVX2 U4823 ( .A(n3431), .Z(n3436) );
  CENX1 U4824 ( .A(n3433), .B(n3432), .Z(n3434) );
  CIVX2 U4825 ( .A(n3434), .Z(n3435) );
  CENX2 U4826 ( .A(n3436), .B(n3435), .Z(n3546) );
  CENX2 U4827 ( .A(n3438), .B(n3437), .Z(n3439) );
  CENX2 U4828 ( .A(n3440), .B(n3439), .Z(n3547) );
  CEO3X2 U4829 ( .A(n3443), .B(n3442), .C(n3441), .Z(n3523) );
  CENX1 U4830 ( .A(h0[12]), .B(n5566), .Z(n3454) );
  CHA1X1 U4831 ( .A(n3446), .B(n3445), .CO(n3443), .S(n3487) );
  CNR2IX1 U4832 ( .B(n7539), .A(n2514), .Z(n3495) );
  CIVX2 U4833 ( .A(h0[13]), .Z(n3447) );
  COND2X2 U4834 ( .A(n7537), .B(n3448), .C(n3493), .D(n5160), .Z(n3496) );
  CND2X2 U4835 ( .A(n3449), .B(n2369), .Z(n6522) );
  CENX1 U4836 ( .A(n6417), .B(h0[3]), .Z(n3500) );
  CNIVX4 U4837 ( .A(n3578), .Z(n5984) );
  COND1X1 U4838 ( .A(n3495), .B(n3496), .C(n3494), .Z(n3451) );
  COND2X1 U4839 ( .A(n6527), .B(n3460), .C(n1586), .D(n3452), .Z(n3476) );
  CENX1 U4840 ( .A(n6118), .B(h0[5]), .Z(n3498) );
  COND2X1 U4841 ( .A(n2568), .B(n3498), .C(n2489), .D(n3453), .Z(n3475) );
  CNIVX4 U4842 ( .A(q0[3]), .Z(n5566) );
  COND2X1 U4843 ( .A(n5695), .B(n3490), .C(n5696), .D(n3454), .Z(n3474) );
  CENX1 U4844 ( .A(n3456), .B(n3455), .Z(n3458) );
  CIVX3 U4845 ( .A(n3345), .Z(n6490) );
  COND2X1 U4846 ( .A(n3461), .B(n2449), .C(n1557), .D(n3460), .Z(n3478) );
  COND2X1 U4847 ( .A(n2449), .B(n3463), .C(n3462), .D(n1556), .Z(n3477) );
  CIVDX3 U4848 ( .A(q0[7]), .Z0(n3643), .Z1(n5909) );
  CENX1 U4849 ( .A(n5909), .B(h0[7]), .Z(n3488) );
  COND2X1 U4850 ( .A(n4959), .B(n3488), .C(n4957), .D(n3464), .Z(n3482) );
  CENX1 U4851 ( .A(n5793), .B(n5927), .Z(n3497) );
  COND2X2 U4852 ( .A(n5912), .B(n3465), .C(n4443), .D(n3497), .Z(n3481) );
  CIVX2 U4853 ( .A(n3526), .Z(n3467) );
  COND1X2 U4854 ( .A(n3468), .B(n3467), .C(n3466), .Z(n3545) );
  COND1X1 U4855 ( .A(n3546), .B(n3547), .C(n1255), .Z(n3470) );
  CND2X1 U4856 ( .A(n3546), .B(n3547), .Z(n3469) );
  CND2X2 U4857 ( .A(n3470), .B(n3469), .Z(n3748) );
  CNR2X1 U4858 ( .A(n3747), .B(n3748), .Z(n4624) );
  CFA1X1 U4859 ( .A(n3473), .B(n3472), .CI(n3471), .CO(n3526), .S(n3541) );
  CFA1X1 U4860 ( .A(n3476), .B(n3475), .CI(n3474), .CO(n3473), .S(n3507) );
  CNIVX4 U4861 ( .A(h0[9]), .Z(n6185) );
  CENXL U4862 ( .A(n6185), .B(n5566), .Z(n3564) );
  CENXL U4863 ( .A(h0[10]), .B(n5104), .Z(n3491) );
  COND2X1 U4864 ( .A(n5695), .B(n3564), .C(n5696), .D(n3491), .Z(n3567) );
  CENX1 U4865 ( .A(n5923), .B(h0[5]), .Z(n3565) );
  CENX1 U4866 ( .A(n5923), .B(n7674), .Z(n3489) );
  COND2X2 U4867 ( .A(n4959), .B(n3565), .C(n4957), .D(n3489), .Z(n3568) );
  CENX1 U4868 ( .A(n6417), .B(h0[1]), .Z(n3517) );
  CENX1 U4869 ( .A(n6417), .B(h0[2]), .Z(n3501) );
  COND2X1 U4870 ( .A(n6211), .B(n3517), .C(n6293), .D(n3501), .Z(n3566) );
  COND1X2 U4871 ( .A(n3567), .B(n3568), .C(n3566), .Z(n3480) );
  CND2X2 U4872 ( .A(n3480), .B(n3479), .Z(n3557) );
  CNR2IX1 U4873 ( .B(n7538), .A(n1557), .Z(n3563) );
  CENX1 U4874 ( .A(n4861), .B(h0[11]), .Z(n3513) );
  CENX1 U4875 ( .A(n3580), .B(h0[12]), .Z(n3492) );
  COND2X1 U4876 ( .A(n5160), .B(n3513), .C(n7537), .D(n3492), .Z(n3562) );
  CENX1 U4877 ( .A(n6118), .B(h0[3]), .Z(n3514) );
  CENX1 U4878 ( .A(n4922), .B(n2513), .Z(n3499) );
  COND2X1 U4879 ( .A(n2575), .B(n3514), .C(n2488), .D(n3499), .Z(n3561) );
  CFA1X1 U4880 ( .A(n3483), .B(n3482), .CI(n3481), .CO(n3471), .S(n3505) );
  CENX2 U4881 ( .A(n3541), .B(n3542), .Z(n3502) );
  CFA1X1 U4882 ( .A(n3486), .B(n3485), .CI(n3484), .CO(n3441), .S(n3528) );
  COND2X1 U4883 ( .A(n6114), .B(n3489), .C(n3368), .D(n3488), .Z(n3510) );
  COND2X1 U4884 ( .A(n5695), .B(n3491), .C(n3490), .D(n4886), .Z(n3509) );
  CENX1 U4885 ( .A(n5793), .B(h0[8]), .Z(n3511) );
  COND2X1 U4886 ( .A(n2566), .B(n3499), .C(n2490), .D(n3498), .Z(n3520) );
  CEO3X2 U4887 ( .A(n3528), .B(n3529), .C(n3527), .Z(n3539) );
  CENX2 U4888 ( .A(n3502), .B(n3539), .Z(n3737) );
  CFA1X1 U4889 ( .A(n3507), .B(n3506), .CI(n3505), .CO(n3542), .S(n3598) );
  CFA1X1 U4890 ( .A(n3509), .B(n3510), .CI(n3508), .CO(n3504), .S(n3560) );
  COND2X1 U4891 ( .A(n4443), .B(n3512), .C(n5912), .D(n3511), .Z(n3592) );
  CENX1 U4892 ( .A(n5793), .B(n7674), .Z(n3584) );
  COND2X2 U4893 ( .A(n5911), .B(n3584), .C(n3512), .D(n5912), .Z(n3574) );
  CENX1 U4894 ( .A(n4861), .B(h0[10]), .Z(n3581) );
  COND2X1 U4895 ( .A(n5160), .B(n3581), .C(n7537), .D(n3513), .Z(n3572) );
  CENX1 U4896 ( .A(n6118), .B(h0[2]), .Z(n3583) );
  COND2X1 U4897 ( .A(n2579), .B(n3583), .C(n2490), .D(n3514), .Z(n3573) );
  CND2X2 U4898 ( .A(n3572), .B(n3574), .Z(n3515) );
  CND2X4 U4899 ( .A(n3516), .B(n3515), .Z(n3595) );
  CENX1 U4900 ( .A(n2597), .B(n7539), .Z(n3518) );
  COND1X2 U4901 ( .A(n3592), .B(n3595), .C(n3593), .Z(n3519) );
  CND2X2 U4902 ( .A(n3522), .B(n3521), .Z(n3736) );
  CENX2 U4903 ( .A(n3524), .B(n3523), .Z(n3525) );
  CENX2 U4904 ( .A(n3525), .B(n3526), .Z(n3551) );
  COND1X1 U4905 ( .A(n3528), .B(n3529), .C(n3527), .Z(n3531) );
  CND2X1 U4906 ( .A(n3529), .B(n3528), .Z(n3530) );
  CND2X2 U4907 ( .A(n3531), .B(n3530), .Z(n3549) );
  CENX2 U4908 ( .A(n3535), .B(n3534), .Z(n3550) );
  CENX2 U4909 ( .A(n3549), .B(n3550), .Z(n3536) );
  CIVX2 U4910 ( .A(n3542), .Z(n3538) );
  CIVX2 U4911 ( .A(n3541), .Z(n3537) );
  CND2X2 U4912 ( .A(n3538), .B(n3537), .Z(n3540) );
  CND2X2 U4913 ( .A(n3540), .B(n3539), .Z(n3544) );
  CND2X2 U4914 ( .A(n3544), .B(n3543), .Z(n3738) );
  CNR2X2 U4915 ( .A(n3739), .B(n3738), .Z(n6376) );
  CNR2X2 U4916 ( .A(n3809), .B(n6376), .Z(n6375) );
  CENX2 U4917 ( .A(n3546), .B(n3545), .Z(n3548) );
  CIVX2 U4918 ( .A(n3741), .Z(n3555) );
  CND2X2 U4919 ( .A(n3553), .B(n3552), .Z(n3740) );
  CIVX2 U4920 ( .A(n3740), .Z(n3554) );
  CND2X2 U4921 ( .A(n3555), .B(n3554), .Z(n6374) );
  CND2X2 U4922 ( .A(n6375), .B(n6374), .Z(n3746) );
  CFA1X1 U4923 ( .A(n3558), .B(n3557), .CI(n3556), .CO(n3506), .S(n3602) );
  CFA1X1 U4924 ( .A(n3563), .B(n3561), .CI(n3562), .CO(n3556), .S(n3588) );
  CENXL U4925 ( .A(h0[8]), .B(n5566), .Z(n3585) );
  CENX1 U4926 ( .A(n5923), .B(n2513), .Z(n3579) );
  CENX1 U4927 ( .A(n3567), .B(n3566), .Z(n3569) );
  CND2X2 U4928 ( .A(n3571), .B(n3570), .Z(n3600) );
  CNIVX1 U4929 ( .A(n3572), .Z(n3577) );
  CIVX2 U4930 ( .A(n3573), .Z(n3575) );
  CENX2 U4931 ( .A(n3575), .B(n3574), .Z(n3576) );
  CENX2 U4932 ( .A(n3577), .B(n3576), .Z(n3608) );
  CNR2IXL U4933 ( .B(n7539), .A(n2369), .Z(n3613) );
  CENX1 U4934 ( .A(n5923), .B(h0[3]), .Z(n3618) );
  COND2X1 U4935 ( .A(n3618), .B(n6114), .C(n3368), .D(n3579), .Z(n3611) );
  CENX1 U4936 ( .A(n3580), .B(n5927), .Z(n3633) );
  COND2X1 U4937 ( .A(n5160), .B(n3633), .C(n7537), .D(n3581), .Z(n3612) );
  CIVX2 U4938 ( .A(n3582), .Z(n3587) );
  CENX1 U4939 ( .A(n5793), .B(h0[5]), .Z(n3617) );
  CENXL U4940 ( .A(h0[7]), .B(n5566), .Z(n3616) );
  CIVX2 U4941 ( .A(n3610), .Z(n3586) );
  COND2X2 U4942 ( .A(n3608), .B(n2656), .C(n3587), .D(n3586), .Z(n3603) );
  CENX2 U4943 ( .A(n3589), .B(n3588), .Z(n3590) );
  CENX2 U4944 ( .A(n3591), .B(n3590), .Z(n3606) );
  CENX1 U4945 ( .A(n3593), .B(n3592), .Z(n3594) );
  CENX1 U4946 ( .A(n3595), .B(n3594), .Z(n3604) );
  CFA1X1 U4947 ( .A(n3602), .B(n3601), .CI(n3600), .CO(n3732), .S(n3731) );
  CNR2X2 U4948 ( .A(n3733), .B(n3732), .Z(n7501) );
  CENX2 U4949 ( .A(n3604), .B(n3603), .Z(n3605) );
  CENX2 U4950 ( .A(n3606), .B(n3605), .Z(n3726) );
  CENX2 U4951 ( .A(n3610), .B(n3609), .Z(n3626) );
  CEO3X2 U4952 ( .A(n3613), .B(n3612), .C(n3611), .Z(n3628) );
  CENXL U4953 ( .A(n5566), .B(n7674), .Z(n3640) );
  COND2X1 U4954 ( .A(n5695), .B(n3640), .C(n4886), .D(n3616), .Z(n3653) );
  CENX1 U4955 ( .A(n5793), .B(n2512), .Z(n3632) );
  COND2X1 U4956 ( .A(n4443), .B(n3632), .C(n5912), .D(n3617), .Z(n3652) );
  CENX1 U4957 ( .A(n5923), .B(h0[2]), .Z(n3644) );
  COND2X1 U4958 ( .A(n6114), .B(n3644), .C(n4957), .D(n3618), .Z(n3651) );
  COND1X1 U4959 ( .A(n3628), .B(n3629), .C(n3630), .Z(n3620) );
  CND2X1 U4960 ( .A(n3628), .B(n3629), .Z(n3619) );
  CND2X2 U4961 ( .A(n3620), .B(n3619), .Z(n3624) );
  CND2X2 U4962 ( .A(n3622), .B(n3621), .Z(n3725) );
  CNR2X1 U4963 ( .A(n3726), .B(n3725), .Z(n3623) );
  CIVX2 U4964 ( .A(n3623), .Z(n6386) );
  CENX2 U4965 ( .A(n3625), .B(n3624), .Z(n3627) );
  CENX2 U4966 ( .A(n3627), .B(n3626), .Z(n3724) );
  CENX1 U4967 ( .A(n3631), .B(h0[7]), .Z(n3659) );
  CENX1 U4968 ( .A(n3631), .B(h0[8]), .Z(n3634) );
  CENX1 U4969 ( .A(n5793), .B(n1232), .Z(n3661) );
  COND2X1 U4970 ( .A(n4443), .B(n3661), .C(n5912), .D(n3632), .Z(n3665) );
  COND2X1 U4971 ( .A(n5160), .B(n3634), .C(n7537), .D(n3633), .Z(n3650) );
  CND2X1 U4972 ( .A(n6386), .B(n6389), .Z(n3729) );
  CENX2 U4973 ( .A(n3637), .B(n3636), .Z(n3639) );
  CENX2 U4974 ( .A(n3639), .B(n3638), .Z(n3720) );
  CENXL U4975 ( .A(n5566), .B(h0[5]), .Z(n3660) );
  COND2X1 U4976 ( .A(n5695), .B(n3660), .C(n3640), .D(n5696), .Z(n3663) );
  CENX1 U4977 ( .A(n7539), .B(n5923), .Z(n3641) );
  CENX1 U4978 ( .A(n5923), .B(h0[1]), .Z(n3645) );
  COND2X1 U4979 ( .A(n4959), .B(n3641), .C(n3368), .D(n3645), .Z(n3669) );
  CND2IX1 U4980 ( .B(n7539), .A(n5923), .Z(n3642) );
  COND2X1 U4981 ( .A(n3643), .B(n6114), .C(n3642), .D(n3368), .Z(n3668) );
  COND2X1 U4982 ( .A(n4959), .B(n3645), .C(n4957), .D(n3644), .Z(n3662) );
  COND1X1 U4983 ( .A(n3663), .B(n3664), .C(n3662), .Z(n3647) );
  CND2X1 U4984 ( .A(n3664), .B(n3663), .Z(n3646) );
  CND2X2 U4985 ( .A(n3647), .B(n3646), .Z(n3657) );
  CEO3X1 U4986 ( .A(n3650), .B(n3649), .C(n3648), .Z(n3658) );
  CFA1X1 U4987 ( .A(n3653), .B(n3652), .CI(n3651), .CO(n3630), .S(n3656) );
  COND1X1 U4988 ( .A(n3657), .B(n3658), .C(n3656), .Z(n3655) );
  CND2X1 U4989 ( .A(n3658), .B(n3657), .Z(n3654) );
  CND2X1 U4990 ( .A(n3655), .B(n3654), .Z(n3719) );
  CNR2X2 U4991 ( .A(n3720), .B(n3719), .Z(n7529) );
  CENX1 U4992 ( .A(n3674), .B(n7674), .Z(n3675) );
  COND2X1 U4993 ( .A(n5160), .B(n3675), .C(n7537), .D(n3659), .Z(n3672) );
  CENXL U4994 ( .A(n5566), .B(n2512), .Z(n3673) );
  COND2X1 U4995 ( .A(n5695), .B(n3673), .C(n5696), .D(n3660), .Z(n3671) );
  CENX1 U4996 ( .A(n5793), .B(h0[2]), .Z(n3679) );
  COND2X1 U4997 ( .A(n4443), .B(n3679), .C(n5912), .D(n3661), .Z(n3670) );
  CNR2X1 U4998 ( .A(n3718), .B(n3717), .Z(n7533) );
  CNR2X1 U4999 ( .A(n7529), .B(n7533), .Z(n3722) );
  CHA1X1 U5000 ( .A(n3669), .B(n3668), .CO(n3664), .S(n3677) );
  CFA1X1 U5001 ( .A(n3672), .B(n3671), .CI(n3670), .CO(n3667), .S(n3678) );
  CENXL U5002 ( .A(n5566), .B(h0[3]), .Z(n3689) );
  CENX1 U5003 ( .A(n3674), .B(h0[5]), .Z(n3686) );
  CNR2X1 U5004 ( .A(n3716), .B(n3715), .Z(n7515) );
  COND2X1 U5005 ( .A(n4443), .B(n3680), .C(n5912), .D(n3679), .Z(n3684) );
  CENX1 U5006 ( .A(n5793), .B(n7539), .Z(n3681) );
  COND2X1 U5007 ( .A(n5911), .B(n3681), .C(n5912), .D(n3680), .Z(n3688) );
  CND2X1 U5008 ( .A(n4399), .B(n5793), .Z(n3682) );
  COND2X1 U5009 ( .A(n5911), .B(n2447), .C(n3682), .D(n5912), .Z(n3687) );
  COR2X1 U5010 ( .A(n3713), .B(n3712), .Z(n7507) );
  CENX1 U5011 ( .A(n4861), .B(n2513), .Z(n3693) );
  CHA1X1 U5012 ( .A(n3688), .B(n3687), .CO(n3683), .S(n3690) );
  CENXL U5013 ( .A(n5566), .B(h0[2]), .Z(n3691) );
  CNR2X1 U5014 ( .A(n3711), .B(n3710), .Z(n7520) );
  CENXL U5015 ( .A(n5566), .B(h0[1]), .Z(n3699) );
  CNR2IX1 U5016 ( .B(n7538), .A(n5912), .Z(n3692) );
  CIVX1 U5017 ( .A(n3692), .Z(n3703) );
  CENX1 U5018 ( .A(n4861), .B(n1232), .Z(n3697) );
  COND2X1 U5019 ( .A(n5160), .B(n3697), .C(n7537), .D(n3693), .Z(n3702) );
  CNR2X1 U5020 ( .A(n3701), .B(n3700), .Z(n4358) );
  CND2X1 U5021 ( .A(n3701), .B(n3700), .Z(n4359) );
  COND1X1 U5022 ( .A(n4360), .B(n4358), .C(n4359), .Z(n7536) );
  CENX1 U5023 ( .A(n3703), .B(n3702), .Z(n3704) );
  CENX1 U5024 ( .A(n3705), .B(n3704), .Z(n3707) );
  COR2X1 U5025 ( .A(n3707), .B(n3706), .Z(n7535) );
  CND2X1 U5026 ( .A(n3707), .B(n3706), .Z(n7534) );
  CND2X1 U5027 ( .A(n3709), .B(n3708), .Z(n4276) );
  CND2X1 U5028 ( .A(n3711), .B(n3710), .Z(n7521) );
  COND1X2 U5029 ( .A(n7520), .B(n7524), .C(n7521), .Z(n7508) );
  CND2X1 U5030 ( .A(n3713), .B(n3712), .Z(n7506) );
  CIVX1 U5031 ( .A(n7506), .Z(n3714) );
  CANR1X1 U5032 ( .A(n7507), .B(n7508), .C(n3714), .Z(n7519) );
  CND2X1 U5033 ( .A(n3716), .B(n3715), .Z(n7516) );
  COND1X1 U5034 ( .A(n7515), .B(n7519), .C(n7516), .Z(n7514) );
  CND2X1 U5035 ( .A(n3718), .B(n3717), .Z(n7531) );
  CND2X1 U5036 ( .A(n3720), .B(n3719), .Z(n7530) );
  COND1X1 U5037 ( .A(n7531), .B(n7529), .C(n7530), .Z(n3721) );
  CANR1X1 U5038 ( .A(n3722), .B(n7514), .C(n3721), .Z(n4086) );
  CND2X1 U5039 ( .A(n3724), .B(n3723), .Z(n4087) );
  CIVX2 U5040 ( .A(n4087), .Z(n6387) );
  CND2X1 U5041 ( .A(n3726), .B(n3725), .Z(n6385) );
  CIVX2 U5042 ( .A(n6385), .Z(n3727) );
  CND2X2 U5043 ( .A(n3731), .B(n3730), .Z(n7504) );
  CND2X2 U5044 ( .A(n3733), .B(n3732), .Z(n7502) );
  COND1X2 U5045 ( .A(n7504), .B(n7501), .C(n7502), .Z(n3734) );
  CANR1X2 U5046 ( .A(n3735), .B(n7500), .C(n3734), .Z(n3808) );
  CND2X2 U5047 ( .A(n3737), .B(n3736), .Z(n6378) );
  CND2X2 U5048 ( .A(n3739), .B(n3738), .Z(n6377) );
  CND2X2 U5049 ( .A(n6378), .B(n6377), .Z(n3744) );
  CIVX2 U5050 ( .A(n6373), .Z(n3742) );
  COND1X2 U5051 ( .A(n3746), .B(n3808), .C(n2346), .Z(n4640) );
  CND2X2 U5052 ( .A(n3748), .B(n3747), .Z(n6384) );
  CND2X2 U5053 ( .A(n3753), .B(n3752), .Z(n4619) );
  CND2X2 U5054 ( .A(n3759), .B(n4419), .Z(n3755) );
  CIVDX4 U5055 ( .A(n4390), .Z0(n6828), .Z1(n3759) );
  CND2X2 U5056 ( .A(n3754), .B(n6828), .Z(n4421) );
  CENX1 U5057 ( .A(n7539), .B(n2456), .Z(n3756) );
  CENXL U5058 ( .A(n6828), .B(h0[1]), .Z(n4437) );
  COND2X1 U5059 ( .A(n2420), .B(n3756), .C(n6770), .D(n4437), .Z(n3757) );
  CIVX2 U5060 ( .A(n3757), .Z(n4516) );
  CNIVX4 U5061 ( .A(n6871), .Z(n6829) );
  CND2IX1 U5062 ( .B(n7539), .A(n2456), .Z(n3758) );
  COND2X1 U5063 ( .A(n6870), .B(n3759), .C(n6829), .D(n3758), .Z(n4517) );
  CENX1 U5064 ( .A(n4516), .B(n4517), .Z(n4563) );
  COND1X1 U5065 ( .A(n3761), .B(n3762), .C(n3760), .Z(n3764) );
  COND1X1 U5066 ( .A(n3767), .B(n3766), .C(n3765), .Z(n3769) );
  CND2X1 U5067 ( .A(n3767), .B(n3766), .Z(n3768) );
  CFA1X1 U5068 ( .A(n3772), .B(n3771), .CI(n3770), .CO(n4559), .S(n3780) );
  CENX1 U5069 ( .A(h0[17]), .B(n5566), .Z(n4434) );
  COND2X1 U5070 ( .A(n5695), .B(n3773), .C(n4886), .D(n4434), .Z(n4461) );
  CENX1 U5071 ( .A(h0[15]), .B(n5793), .Z(n4442) );
  COND2X1 U5072 ( .A(n5911), .B(n3774), .C(n5912), .D(n4442), .Z(n4460) );
  CENX1 U5073 ( .A(n6417), .B(n5927), .Z(n4446) );
  COND2X1 U5074 ( .A(n6522), .B(n3775), .C(n6523), .D(n4446), .Z(n4459) );
  CENX1 U5075 ( .A(n6491), .B(h0[7]), .Z(n4445) );
  COND2X1 U5076 ( .A(n2449), .B(n3776), .C(n1556), .D(n4445), .Z(n4458) );
  CENX1 U5077 ( .A(n5923), .B(h0[13]), .Z(n4515) );
  CENX1 U5078 ( .A(n5106), .B(h0[19]), .Z(n4393) );
  CEO3X2 U5079 ( .A(n4559), .B(n4558), .C(n4560), .Z(n4617) );
  CENX2 U5080 ( .A(n4618), .B(n4617), .Z(n3779) );
  CENX2 U5081 ( .A(n4619), .B(n3779), .Z(n4630) );
  CIVX2 U5082 ( .A(n3780), .Z(n3785) );
  CNR2X1 U5083 ( .A(n3781), .B(n3782), .Z(n3784) );
  CND2X1 U5084 ( .A(n3782), .B(n3781), .Z(n3783) );
  COND1X2 U5085 ( .A(n3785), .B(n3784), .C(n3783), .Z(n4595) );
  CENX1 U5086 ( .A(n6118), .B(h0[11]), .Z(n4518) );
  COND2X1 U5087 ( .A(n2563), .B(n3786), .C(n2488), .D(n4518), .Z(n4457) );
  CENX1 U5088 ( .A(n6647), .B(h0[5]), .Z(n4435) );
  COND2X1 U5089 ( .A(n2277), .B(n3787), .C(n2514), .D(n4435), .Z(n4456) );
  CIVX8 U5090 ( .A(n3788), .Z(n6701) );
  CENX1 U5091 ( .A(n6409), .B(h0[3]), .Z(n4392) );
  COND2X1 U5092 ( .A(n6701), .B(n3789), .C(n6765), .D(n4392), .Z(n4455) );
  CFA1X1 U5093 ( .A(n3792), .B(n3791), .CI(n3790), .CO(n4593), .S(n3795) );
  CENX2 U5094 ( .A(n4594), .B(n4593), .Z(n3793) );
  CENX2 U5095 ( .A(n4595), .B(n3793), .Z(n4631) );
  COND1X2 U5096 ( .A(n3795), .B(n3796), .C(n3794), .Z(n3798) );
  CND2X2 U5097 ( .A(n3796), .B(n3795), .Z(n3797) );
  CND2X2 U5098 ( .A(n3798), .B(n3797), .Z(n4629) );
  CENX2 U5099 ( .A(n4631), .B(n4629), .Z(n3799) );
  CENX2 U5100 ( .A(n4630), .B(n3799), .Z(n3806) );
  CND2X2 U5101 ( .A(n3804), .B(n3803), .Z(n3805) );
  CND2X2 U5102 ( .A(n3805), .B(n3806), .Z(n4634) );
  CNR2X2 U5103 ( .A(n3806), .B(n3805), .Z(n3807) );
  CIVX3 U5104 ( .A(n3807), .Z(n4635) );
  CIVXL U5105 ( .A(n3808), .Z(n6379) );
  CIVX2 U5106 ( .A(n3809), .Z(n6380) );
  CANR2XL U5107 ( .A(n7808), .B(out0_2[61]), .C(out1_2[61]), .D(n4053), .Z(
        n3810) );
  COND1XL U5108 ( .A(n7941), .B(n7810), .C(n3810), .Z(n3811) );
  CNR2XL U5109 ( .A(n3811), .B(out1_1[61]), .Z(n4059) );
  CND2XL U5110 ( .A(n3811), .B(out1_1[61]), .Z(n4058) );
  CANR2XL U5111 ( .A(n7808), .B(out0_2[32]), .C(out1_2[32]), .D(n3902), .Z(
        n3812) );
  COND1XL U5112 ( .A(n7993), .B(n7810), .C(n3812), .Z(n3950) );
  CNR2X1 U5113 ( .A(n3950), .B(out1_1[32]), .Z(n4109) );
  CANR2XL U5114 ( .A(n7808), .B(out0_2[33]), .C(out1_2[33]), .D(n3902), .Z(
        n3813) );
  COND1XL U5115 ( .A(n7991), .B(n7810), .C(n3813), .Z(n3951) );
  CNR2X1 U5116 ( .A(n3951), .B(out1_1[33]), .Z(n4107) );
  CNR2X1 U5117 ( .A(n4109), .B(n4107), .Z(n7670) );
  CIVXL U5118 ( .A(acc[34]), .Z(n3815) );
  CANR2XL U5119 ( .A(n7808), .B(out0_2[34]), .C(out1_2[34]), .D(n3902), .Z(
        n3814) );
  COND1XL U5120 ( .A(n3815), .B(n7810), .C(n3814), .Z(n3952) );
  CNR2X1 U5121 ( .A(n3952), .B(out1_1[34]), .Z(n7666) );
  CANR2XL U5122 ( .A(n7808), .B(out0_2[35]), .C(out1_2[35]), .D(n3902), .Z(
        n3816) );
  COND1XL U5123 ( .A(n7988), .B(n7810), .C(n3816), .Z(n3953) );
  CNR2XL U5124 ( .A(n3953), .B(out1_1[35]), .Z(n4006) );
  CNR2X1 U5125 ( .A(n7666), .B(n4006), .Z(n3954) );
  CND2X1 U5126 ( .A(n7670), .B(n3954), .Z(n4026) );
  CANR2XL U5127 ( .A(n7808), .B(out0_2[36]), .C(out1_2[36]), .D(n3902), .Z(
        n3817) );
  COND1XL U5128 ( .A(n7986), .B(n7810), .C(n3817), .Z(n3955) );
  CNR2X1 U5129 ( .A(n3955), .B(out1_1[36]), .Z(n4041) );
  CANR2XL U5130 ( .A(n7808), .B(out0_2[37]), .C(out1_2[37]), .D(n3902), .Z(
        n3818) );
  COND1XL U5131 ( .A(n7984), .B(n7810), .C(n3818), .Z(n3956) );
  CNR2X1 U5132 ( .A(n3956), .B(out1_1[37]), .Z(n4004) );
  CNR2X1 U5133 ( .A(n4041), .B(n4004), .Z(n4029) );
  CANR2XL U5134 ( .A(n7808), .B(out0_2[38]), .C(out1_2[38]), .D(n3902), .Z(
        n3819) );
  COND1XL U5135 ( .A(n7982), .B(n7810), .C(n3819), .Z(n3957) );
  CNR2XL U5136 ( .A(n3957), .B(out1_1[38]), .Z(n4037) );
  CANR2XL U5137 ( .A(n7808), .B(out0_2[39]), .C(out1_2[39]), .D(n3902), .Z(
        n3820) );
  COND1XL U5138 ( .A(n7980), .B(n7810), .C(n3820), .Z(n3958) );
  CNR2XL U5139 ( .A(n3958), .B(out1_1[39]), .Z(n4024) );
  CNR2XL U5140 ( .A(n4037), .B(n4024), .Z(n3960) );
  CND2X1 U5141 ( .A(n4029), .B(n3960), .Z(n3962) );
  CNR2X1 U5142 ( .A(n4026), .B(n3962), .Z(n7649) );
  CIVXL U5143 ( .A(acc[40]), .Z(n3822) );
  CANR2XL U5144 ( .A(n4054), .B(out0_2[40]), .C(out1_2[40]), .D(n3868), .Z(
        n3821) );
  COND1XL U5145 ( .A(n3822), .B(n7810), .C(n3821), .Z(n3963) );
  CNR2X1 U5146 ( .A(n3963), .B(out1_1[40]), .Z(n7645) );
  CIVXL U5147 ( .A(acc[41]), .Z(n3824) );
  CANR2XL U5148 ( .A(n4054), .B(out0_2[41]), .C(out1_2[41]), .D(n3868), .Z(
        n3823) );
  COND1XL U5149 ( .A(n3824), .B(n7810), .C(n3823), .Z(n3964) );
  CNR2X1 U5150 ( .A(n3964), .B(out1_1[41]), .Z(n4045) );
  CNR2X1 U5151 ( .A(n7645), .B(n4045), .Z(n7655) );
  CANR2XL U5152 ( .A(n4054), .B(out0_2[42]), .C(out1_2[42]), .D(n3902), .Z(
        n3825) );
  COND1XL U5153 ( .A(n7976), .B(n7810), .C(n3825), .Z(n3965) );
  CNR2XL U5154 ( .A(n3965), .B(out1_1[42]), .Z(n4036) );
  CIVXL U5155 ( .A(acc[43]), .Z(n3827) );
  CANR2XL U5156 ( .A(n4054), .B(out0_2[43]), .C(out1_2[43]), .D(n3902), .Z(
        n3826) );
  COND1XL U5157 ( .A(n3827), .B(n7810), .C(n3826), .Z(n3966) );
  CNR2XL U5158 ( .A(n3966), .B(out1_1[43]), .Z(n4034) );
  CNR2XL U5159 ( .A(n4036), .B(n4034), .Z(n3968) );
  CND2X1 U5160 ( .A(n7655), .B(n3968), .Z(n4022) );
  CANR2XL U5161 ( .A(n4054), .B(out0_2[44]), .C(out1_2[44]), .D(n3902), .Z(
        n3828) );
  COND1XL U5162 ( .A(n7973), .B(n7810), .C(n3828), .Z(n3969) );
  CNR2X1 U5163 ( .A(n3969), .B(out1_1[44]), .Z(n3998) );
  CANR2XL U5164 ( .A(n4054), .B(out0_2[45]), .C(out1_2[45]), .D(n3902), .Z(
        n3829) );
  COND1XL U5165 ( .A(n7971), .B(n7810), .C(n3829), .Z(n3970) );
  CNR2X1 U5166 ( .A(n3970), .B(out1_1[45]), .Z(n4030) );
  CNR2X1 U5167 ( .A(n3998), .B(n4030), .Z(n4078) );
  CIVXL U5168 ( .A(acc[46]), .Z(n3831) );
  CANR2XL U5169 ( .A(n4054), .B(out0_2[46]), .C(out1_2[46]), .D(n3902), .Z(
        n3830) );
  COND1XL U5170 ( .A(n3831), .B(n7810), .C(n3830), .Z(n3971) );
  CNR2X1 U5171 ( .A(n3971), .B(out1_1[46]), .Z(n4072) );
  CIVXL U5172 ( .A(acc[47]), .Z(n3833) );
  CANR2XL U5173 ( .A(n4054), .B(out0_2[47]), .C(out1_2[47]), .D(n3902), .Z(
        n3832) );
  COND1XL U5174 ( .A(n3833), .B(n7810), .C(n3832), .Z(n3972) );
  CNR2XL U5175 ( .A(n3972), .B(out1_1[47]), .Z(n4020) );
  CNR2XL U5176 ( .A(n4072), .B(n4020), .Z(n3974) );
  CND2X1 U5177 ( .A(n4078), .B(n3974), .Z(n3976) );
  CNR2X1 U5178 ( .A(n4022), .B(n3976), .Z(n3978) );
  CND2X1 U5179 ( .A(n7649), .B(n3978), .Z(n7818) );
  CIVXL U5180 ( .A(acc[48]), .Z(n3835) );
  CANR2XL U5181 ( .A(n4054), .B(out0_2[48]), .C(out1_2[48]), .D(n3902), .Z(
        n3834) );
  COND1XL U5182 ( .A(n3835), .B(n7810), .C(n3834), .Z(n3979) );
  CNR2X1 U5183 ( .A(n3979), .B(out1_1[48]), .Z(n4134) );
  CANR2XL U5184 ( .A(n4054), .B(out0_2[49]), .C(out1_2[49]), .D(n3902), .Z(
        n3836) );
  COND1XL U5185 ( .A(n7966), .B(n7810), .C(n3836), .Z(n3980) );
  CNR2X1 U5186 ( .A(n3980), .B(out1_1[49]), .Z(n4131) );
  CNR2X1 U5187 ( .A(n4134), .B(n4131), .Z(n4129) );
  CANR2XL U5188 ( .A(n4054), .B(out0_2[50]), .C(out1_2[50]), .D(n3902), .Z(
        n3837) );
  COND1XL U5189 ( .A(n7964), .B(n7810), .C(n3837), .Z(n3981) );
  CNR2X1 U5190 ( .A(n3981), .B(out1_1[50]), .Z(n4098) );
  CANR2XL U5191 ( .A(n4054), .B(out0_2[51]), .C(out1_2[51]), .D(n3868), .Z(
        n3838) );
  COND1XL U5192 ( .A(n7962), .B(n7810), .C(n3838), .Z(n3982) );
  CNR2X1 U5193 ( .A(n3982), .B(out1_1[51]), .Z(n4096) );
  CNR2X1 U5194 ( .A(n4098), .B(n4096), .Z(n3983) );
  CND2X1 U5195 ( .A(n4129), .B(n3983), .Z(n4101) );
  CANR2XL U5196 ( .A(n7808), .B(out0_2[52]), .C(out1_2[52]), .D(n3902), .Z(
        n3839) );
  COND1XL U5197 ( .A(n7960), .B(n7810), .C(n3839), .Z(n3984) );
  CNR2X1 U5198 ( .A(n3984), .B(out1_1[52]), .Z(n4099) );
  CANR2XL U5199 ( .A(n4054), .B(out0_2[53]), .C(out1_2[53]), .D(n3902), .Z(
        n3840) );
  COND1XL U5200 ( .A(n7958), .B(n7810), .C(n3840), .Z(n3985) );
  CNR2X1 U5201 ( .A(n3985), .B(out1_1[53]), .Z(n4111) );
  CNR2X1 U5202 ( .A(n4099), .B(n4111), .Z(n4137) );
  CANR2XL U5203 ( .A(n4054), .B(out0_2[54]), .C(out1_2[54]), .D(n3868), .Z(
        n3841) );
  COND1XL U5204 ( .A(n7956), .B(n7810), .C(n3841), .Z(n3986) );
  CNR2XL U5205 ( .A(n3986), .B(out1_1[54]), .Z(n4141) );
  CANR2XL U5206 ( .A(n7808), .B(out0_2[55]), .C(out1_2[55]), .D(n3902), .Z(
        n3842) );
  COND1XL U5207 ( .A(n7954), .B(n7810), .C(n3842), .Z(n3987) );
  CNR2XL U5208 ( .A(n3987), .B(out1_1[55]), .Z(n4135) );
  CNR2XL U5209 ( .A(n4141), .B(n4135), .Z(n3989) );
  CND2X1 U5210 ( .A(n4137), .B(n3989), .Z(n3991) );
  CNR2X1 U5211 ( .A(n4101), .B(n3991), .Z(n7817) );
  CANR2XL U5212 ( .A(n4054), .B(out0_2[56]), .C(out1_2[56]), .D(n4053), .Z(
        n3843) );
  COND1XL U5213 ( .A(n7952), .B(n7810), .C(n3843), .Z(n3992) );
  CNR2X1 U5214 ( .A(n3992), .B(out1_1[56]), .Z(n4110) );
  CANR2XL U5215 ( .A(n7808), .B(out0_2[57]), .C(out1_2[57]), .D(n4053), .Z(
        n3844) );
  COND1XL U5216 ( .A(n7950), .B(n7810), .C(n3844), .Z(n3993) );
  CNR2X1 U5217 ( .A(n3993), .B(out1_1[57]), .Z(n4143) );
  CNR2X1 U5218 ( .A(n4110), .B(n4143), .Z(n4119) );
  CANR2XL U5219 ( .A(n4054), .B(out0_2[58]), .C(out1_2[58]), .D(n4053), .Z(
        n3845) );
  COND1XL U5220 ( .A(n7948), .B(n7810), .C(n3845), .Z(n3994) );
  CNR2X1 U5221 ( .A(n3994), .B(out1_1[58]), .Z(n4115) );
  CANR2XL U5222 ( .A(n7808), .B(out0_2[59]), .C(out1_2[59]), .D(n4053), .Z(
        n3846) );
  COND1XL U5223 ( .A(n7946), .B(n7810), .C(n3846), .Z(n3995) );
  CNR2X1 U5224 ( .A(n3995), .B(out1_1[59]), .Z(n4008) );
  CNR2X1 U5225 ( .A(n4115), .B(n4008), .Z(n3996) );
  CND2X1 U5226 ( .A(n4119), .B(n3996), .Z(n7816) );
  CANR2XL U5227 ( .A(n7808), .B(out0_2[60]), .C(out1_2[60]), .D(n4053), .Z(
        n3847) );
  COND1XL U5228 ( .A(n7944), .B(n7810), .C(n3847), .Z(n3997) );
  CNR2XL U5229 ( .A(n3997), .B(out1_1[60]), .Z(n4057) );
  CANR2XL U5230 ( .A(n7808), .B(out0_2[16]), .C(out1_2[16]), .D(n3902), .Z(
        n3848) );
  COND1XL U5231 ( .A(n8015), .B(n7810), .C(n3848), .Z(n3920) );
  CNR2XL U5232 ( .A(n3920), .B(out1_1[16]), .Z(n4162) );
  CANR2XL U5233 ( .A(n4054), .B(out0_2[17]), .C(out1_2[17]), .D(n3902), .Z(
        n3849) );
  COND1XL U5234 ( .A(n8014), .B(n7810), .C(n3849), .Z(n3921) );
  CNR2X1 U5235 ( .A(n3921), .B(out1_1[17]), .Z(n4160) );
  CNR2XL U5236 ( .A(n4162), .B(n4160), .Z(n7807) );
  CANR2XL U5237 ( .A(n7808), .B(out0_2[18]), .C(out1_2[18]), .D(n3902), .Z(
        n3850) );
  COND1XL U5238 ( .A(n3851), .B(n7810), .C(n3850), .Z(n3922) );
  CNR2X1 U5239 ( .A(n3922), .B(out1_1[18]), .Z(n7803) );
  CANR2XL U5240 ( .A(n4054), .B(out0_2[19]), .C(out1_2[19]), .D(n3902), .Z(
        n3852) );
  COND1XL U5241 ( .A(n3853), .B(n7810), .C(n3852), .Z(n3923) );
  CNR2XL U5242 ( .A(n3923), .B(out1_1[19]), .Z(n7793) );
  CNR2X1 U5243 ( .A(n7803), .B(n7793), .Z(n3924) );
  CND2X1 U5244 ( .A(n7807), .B(n3924), .Z(n4176) );
  CANR2XL U5245 ( .A(n7808), .B(out0_2[20]), .C(out1_2[20]), .D(n3902), .Z(
        n3854) );
  COND1XL U5246 ( .A(n3855), .B(n7810), .C(n3854), .Z(n3925) );
  CNR2X1 U5247 ( .A(n3925), .B(out1_1[20]), .Z(n4173) );
  CIVX1 U5248 ( .A(n3883), .Z(n3868) );
  CANR2XL U5249 ( .A(n7808), .B(out0_2[21]), .C(out1_2[21]), .D(n3868), .Z(
        n3856) );
  COND1XL U5250 ( .A(n3857), .B(n7810), .C(n3856), .Z(n3926) );
  CNR2X1 U5251 ( .A(n3926), .B(out1_1[21]), .Z(n4163) );
  CNR2X1 U5252 ( .A(n4173), .B(n4163), .Z(n4185) );
  CANR2XL U5253 ( .A(n4054), .B(out0_2[22]), .C(out1_2[22]), .D(n3868), .Z(
        n3858) );
  COND1XL U5254 ( .A(n3859), .B(n7810), .C(n3858), .Z(n3927) );
  CNR2XL U5255 ( .A(n3927), .B(out1_1[22]), .Z(n4201) );
  CANR2XL U5256 ( .A(n7808), .B(out0_2[23]), .C(out1_2[23]), .D(n3868), .Z(
        n3860) );
  COND1XL U5257 ( .A(n3861), .B(n7810), .C(n3860), .Z(n3928) );
  CNR2XL U5258 ( .A(n3928), .B(out1_1[23]), .Z(n4195) );
  CNR2XL U5259 ( .A(n4201), .B(n4195), .Z(n3929) );
  CND2X1 U5260 ( .A(n4185), .B(n3929), .Z(n3930) );
  CNR2X1 U5261 ( .A(n4176), .B(n3930), .Z(n7570) );
  CANR2XL U5262 ( .A(n4054), .B(out0_2[24]), .C(out1_2[24]), .D(n3868), .Z(
        n3862) );
  COND1XL U5263 ( .A(n3863), .B(n7810), .C(n3862), .Z(n3931) );
  CNR2X1 U5264 ( .A(n3931), .B(out1_1[24]), .Z(n7566) );
  CANR2XL U5265 ( .A(n4054), .B(out0_2[25]), .C(out1_2[25]), .D(n3868), .Z(
        n3864) );
  COND1XL U5266 ( .A(n3865), .B(n7810), .C(n3864), .Z(n3932) );
  CNR2X1 U5267 ( .A(n3932), .B(out1_1[25]), .Z(n4165) );
  CNR2X1 U5268 ( .A(n7566), .B(n4165), .Z(n7634) );
  CIVXL U5269 ( .A(acc[26]), .Z(n3867) );
  CANR2XL U5270 ( .A(n7808), .B(out0_2[26]), .C(out1_2[26]), .D(n3868), .Z(
        n3866) );
  COND1XL U5271 ( .A(n3867), .B(n7810), .C(n3866), .Z(n3933) );
  CNR2X1 U5272 ( .A(n3933), .B(out1_1[26]), .Z(n4150) );
  CIVXL U5273 ( .A(acc[27]), .Z(n3870) );
  CANR2XL U5274 ( .A(n4054), .B(out0_2[27]), .C(out1_2[27]), .D(n3868), .Z(
        n3869) );
  COND1XL U5275 ( .A(n3870), .B(n7810), .C(n3869), .Z(n3934) );
  CNR2X1 U5276 ( .A(n3934), .B(out1_1[27]), .Z(n4147) );
  CNR2X1 U5277 ( .A(n4150), .B(n4147), .Z(n3936) );
  CND2X1 U5278 ( .A(n7634), .B(n3936), .Z(n7592) );
  CANR2XL U5279 ( .A(n7808), .B(out0_2[28]), .C(out1_2[28]), .D(n3902), .Z(
        n3871) );
  COND1XL U5280 ( .A(n7996), .B(n7810), .C(n3871), .Z(n3937) );
  CNR2X1 U5281 ( .A(n3937), .B(out1_1[28]), .Z(n4167) );
  CIVXL U5282 ( .A(acc[29]), .Z(n3873) );
  CANR2XL U5283 ( .A(n7808), .B(out0_2[29]), .C(out1_2[29]), .D(n3868), .Z(
        n3872) );
  COND1XL U5284 ( .A(n3873), .B(n7810), .C(n3872), .Z(n3938) );
  CNR2X1 U5285 ( .A(n3938), .B(out1_1[29]), .Z(n7589) );
  CNR2X1 U5286 ( .A(n4167), .B(n7589), .Z(n7615) );
  CIVXL U5287 ( .A(acc[30]), .Z(n3875) );
  CANR2XL U5288 ( .A(n7808), .B(out0_2[30]), .C(out1_2[30]), .D(n3902), .Z(
        n3874) );
  COND1XL U5289 ( .A(n3875), .B(n7810), .C(n3874), .Z(n3939) );
  CNR2X1 U5290 ( .A(n3939), .B(out1_1[30]), .Z(n7621) );
  CIVXL U5291 ( .A(acc[31]), .Z(n3877) );
  CANR2XL U5292 ( .A(n7808), .B(out0_2[31]), .C(out1_2[31]), .D(n3902), .Z(
        n3876) );
  COND1XL U5293 ( .A(n3877), .B(n7810), .C(n3876), .Z(n3940) );
  CNR2XL U5294 ( .A(n3940), .B(out1_1[31]), .Z(n7612) );
  CNR2XL U5295 ( .A(n7621), .B(n7612), .Z(n3942) );
  CND2XL U5296 ( .A(n7615), .B(n3942), .Z(n3944) );
  CNR2X1 U5297 ( .A(n7592), .B(n3944), .Z(n3946) );
  CND2X1 U5298 ( .A(n7570), .B(n3946), .Z(n3948) );
  CANR2XL U5299 ( .A(n7808), .B(out0_2[5]), .C(out1_2[5]), .D(n4053), .Z(n3878) );
  COND1XL U5300 ( .A(n3879), .B(n7810), .C(n3878), .Z(n3886) );
  CNR2XL U5301 ( .A(n3886), .B(out1_1[5]), .Z(n4236) );
  CNR2XL U5302 ( .A(n3880), .B(n4236), .Z(n7789) );
  CANR2XL U5303 ( .A(n7808), .B(out0_2[6]), .C(out1_2[6]), .D(n4053), .Z(n3881) );
  COND1XL U5304 ( .A(n3882), .B(n7810), .C(n3881), .Z(n3887) );
  CNR2XL U5305 ( .A(n3887), .B(out1_1[6]), .Z(n7785) );
  CANR2XL U5306 ( .A(n7808), .B(out0_2[7]), .C(out1_2[7]), .D(n3868), .Z(n3884) );
  COND1XL U5307 ( .A(n3885), .B(n7810), .C(n3884), .Z(n3888) );
  CNR2XL U5308 ( .A(n3888), .B(out1_1[7]), .Z(n4234) );
  CNR2XL U5309 ( .A(n7785), .B(n4234), .Z(n3890) );
  CND2XL U5310 ( .A(n7789), .B(n3890), .Z(n3893) );
  CND2XL U5311 ( .A(n3886), .B(out1_1[5]), .Z(n4237) );
  COND1XL U5312 ( .A(n4238), .B(n4236), .C(n4237), .Z(n7787) );
  CND2XL U5313 ( .A(n3887), .B(out1_1[6]), .Z(n7786) );
  CND2XL U5314 ( .A(n3888), .B(out1_1[7]), .Z(n4235) );
  COND1XL U5315 ( .A(n7786), .B(n4234), .C(n4235), .Z(n3889) );
  CANR1XL U5316 ( .A(n7787), .B(n3890), .C(n3889), .Z(n3891) );
  COND1X1 U5317 ( .A(n3893), .B(n3892), .C(n3891), .Z(n4207) );
  CANR2XL U5318 ( .A(n7808), .B(out0_2[8]), .C(out1_2[8]), .D(n3868), .Z(n3894) );
  COND1XL U5319 ( .A(n8007), .B(n7810), .C(n3894), .Z(n3905) );
  CNR2X1 U5320 ( .A(n3905), .B(out1_1[8]), .Z(n7790) );
  CANR2XL U5321 ( .A(n7808), .B(out0_2[9]), .C(out1_2[9]), .D(n3868), .Z(n3895) );
  COND1XL U5322 ( .A(n8006), .B(n7810), .C(n3895), .Z(n3906) );
  CNR2X1 U5323 ( .A(n3906), .B(out1_1[9]), .Z(n4208) );
  CNR2X1 U5324 ( .A(n7790), .B(n4208), .Z(n4220) );
  CANR2XL U5325 ( .A(n7808), .B(out0_2[10]), .C(out1_2[10]), .D(n3902), .Z(
        n3896) );
  COND1XL U5326 ( .A(n8005), .B(n7810), .C(n3896), .Z(n3907) );
  CNR2X1 U5327 ( .A(n3907), .B(out1_1[10]), .Z(n4210) );
  CNR2XL U5328 ( .A(n3908), .B(out1_1[11]), .Z(n4224) );
  CNR2X1 U5329 ( .A(n4210), .B(n4224), .Z(n3909) );
  CND2X1 U5330 ( .A(n4220), .B(n3909), .Z(n4217) );
  CANR2XL U5331 ( .A(n7808), .B(out0_2[12]), .C(out1_2[12]), .D(n3902), .Z(
        n3897) );
  COND1XL U5332 ( .A(n8017), .B(n7810), .C(n3897), .Z(n3910) );
  CNR2X1 U5333 ( .A(n3910), .B(out1_1[12]), .Z(n4213) );
  CANR2XL U5334 ( .A(n7808), .B(out0_2[13]), .C(out1_2[13]), .D(n3902), .Z(
        n3898) );
  COND1XL U5335 ( .A(n3899), .B(n7810), .C(n3898), .Z(n3911) );
  CNR2X1 U5336 ( .A(n3911), .B(out1_1[13]), .Z(n4214) );
  CNR2X1 U5337 ( .A(n4213), .B(n4214), .Z(n4226) );
  CIVXL U5338 ( .A(acc[14]), .Z(n3901) );
  CANR2XL U5339 ( .A(n7808), .B(out0_2[14]), .C(out1_2[14]), .D(n3902), .Z(
        n3900) );
  COND1XL U5340 ( .A(n3901), .B(n7810), .C(n3900), .Z(n3912) );
  CNR2XL U5341 ( .A(n3912), .B(out1_1[14]), .Z(n4230) );
  CANR2XL U5342 ( .A(n7808), .B(out0_2[15]), .C(out1_2[15]), .D(n3902), .Z(
        n3903) );
  COND1XL U5343 ( .A(n3904), .B(n7810), .C(n3903), .Z(n3913) );
  CNR2XL U5344 ( .A(n3913), .B(out1_1[15]), .Z(n4232) );
  CNR2XL U5345 ( .A(n4230), .B(n4232), .Z(n3915) );
  CND2X1 U5346 ( .A(n4226), .B(n3915), .Z(n3917) );
  CNR2X1 U5347 ( .A(n4217), .B(n3917), .Z(n3919) );
  CND2X1 U5348 ( .A(n3905), .B(out1_1[8]), .Z(n7791) );
  CND2X1 U5349 ( .A(n3906), .B(out1_1[9]), .Z(n4209) );
  COND1X1 U5350 ( .A(n7791), .B(n4208), .C(n4209), .Z(n4222) );
  CND2X1 U5351 ( .A(n3907), .B(out1_1[10]), .Z(n4221) );
  CND2XL U5352 ( .A(n3908), .B(out1_1[11]), .Z(n4225) );
  CND2X1 U5353 ( .A(n3910), .B(out1_1[12]), .Z(n4218) );
  CND2XL U5354 ( .A(n3911), .B(out1_1[13]), .Z(n4215) );
  COND1XL U5355 ( .A(n4218), .B(n4214), .C(n4215), .Z(n4228) );
  CND2XL U5356 ( .A(n3912), .B(out1_1[14]), .Z(n4229) );
  CND2XL U5357 ( .A(n3913), .B(out1_1[15]), .Z(n4233) );
  COND1XL U5358 ( .A(n4229), .B(n4232), .C(n4233), .Z(n3914) );
  CANR1XL U5359 ( .A(n4228), .B(n3915), .C(n3914), .Z(n3916) );
  COND1X1 U5360 ( .A(n3917), .B(n4216), .C(n3916), .Z(n3918) );
  CANR1X1 U5361 ( .A(n4207), .B(n3919), .C(n3918), .Z(n4151) );
  CND2X1 U5362 ( .A(n3920), .B(out1_1[16]), .Z(n4211) );
  CND2XL U5363 ( .A(n3921), .B(out1_1[17]), .Z(n4161) );
  COND1X1 U5364 ( .A(n4211), .B(n4160), .C(n4161), .Z(n7805) );
  CND2XL U5365 ( .A(n3922), .B(out1_1[18]), .Z(n7804) );
  CND2XL U5366 ( .A(n3923), .B(out1_1[19]), .Z(n7794) );
  CND2XL U5367 ( .A(n3925), .B(out1_1[20]), .Z(n4174) );
  CND2XL U5368 ( .A(n3926), .B(out1_1[21]), .Z(n4164) );
  COND1XL U5369 ( .A(n4174), .B(n4163), .C(n4164), .Z(n4183) );
  CND2XL U5370 ( .A(n3927), .B(out1_1[22]), .Z(n4199) );
  CND2XL U5371 ( .A(n3928), .B(out1_1[23]), .Z(n4196) );
  CND2XL U5372 ( .A(n3931), .B(out1_1[24]), .Z(n7567) );
  CND2XL U5373 ( .A(n3932), .B(out1_1[25]), .Z(n4166) );
  COND1XL U5374 ( .A(n7567), .B(n4165), .C(n4166), .Z(n7636) );
  CND2XL U5375 ( .A(n3933), .B(out1_1[26]), .Z(n7632) );
  CND2XL U5376 ( .A(n3934), .B(out1_1[27]), .Z(n4148) );
  COND1XL U5377 ( .A(n7632), .B(n4147), .C(n4148), .Z(n3935) );
  CANR1XL U5378 ( .A(n7636), .B(n3936), .C(n3935), .Z(n7593) );
  CND2XL U5379 ( .A(n3937), .B(out1_1[28]), .Z(n7594) );
  CND2XL U5380 ( .A(n3938), .B(out1_1[29]), .Z(n7590) );
  COND1XL U5381 ( .A(n7594), .B(n7589), .C(n7590), .Z(n7618) );
  CND2XL U5382 ( .A(n3939), .B(out1_1[30]), .Z(n7619) );
  CND2XL U5383 ( .A(n3940), .B(out1_1[31]), .Z(n7613) );
  COND1XL U5384 ( .A(n7619), .B(n7612), .C(n7613), .Z(n3941) );
  CANR1XL U5385 ( .A(n7618), .B(n3942), .C(n3941), .Z(n3943) );
  COND1XL U5386 ( .A(n3944), .B(n7593), .C(n3943), .Z(n3945) );
  CANR1X1 U5387 ( .A(n7569), .B(n3946), .C(n3945), .Z(n3947) );
  CND2X1 U5388 ( .A(n3950), .B(out1_1[32]), .Z(n4191) );
  CND2XL U5389 ( .A(n3951), .B(out1_1[33]), .Z(n4108) );
  COND1X1 U5390 ( .A(n4191), .B(n4107), .C(n4108), .Z(n7669) );
  CND2XL U5391 ( .A(n3952), .B(out1_1[34]), .Z(n7667) );
  CND2XL U5392 ( .A(n3953), .B(out1_1[35]), .Z(n4007) );
  CND2XL U5393 ( .A(n3955), .B(out1_1[36]), .Z(n4042) );
  CND2XL U5394 ( .A(n3956), .B(out1_1[37]), .Z(n4005) );
  COND1XL U5395 ( .A(n4042), .B(n4004), .C(n4005), .Z(n4028) );
  CND2XL U5396 ( .A(n3957), .B(out1_1[38]), .Z(n4038) );
  CND2XL U5397 ( .A(n3958), .B(out1_1[39]), .Z(n4025) );
  COND1XL U5398 ( .A(n4038), .B(n4024), .C(n4025), .Z(n3959) );
  CANR1XL U5399 ( .A(n4028), .B(n3960), .C(n3959), .Z(n3961) );
  COND1X1 U5400 ( .A(n3962), .B(n4027), .C(n3961), .Z(n7648) );
  CND2XL U5401 ( .A(n3963), .B(out1_1[40]), .Z(n7646) );
  CND2XL U5402 ( .A(n3964), .B(out1_1[41]), .Z(n4046) );
  COND1XL U5403 ( .A(n7646), .B(n4045), .C(n4046), .Z(n7657) );
  CND2XL U5404 ( .A(n3965), .B(out1_1[42]), .Z(n7653) );
  CND2XL U5405 ( .A(n3966), .B(out1_1[43]), .Z(n4035) );
  COND1XL U5406 ( .A(n7653), .B(n4034), .C(n4035), .Z(n3967) );
  CANR1XL U5407 ( .A(n7657), .B(n3968), .C(n3967), .Z(n4023) );
  CND2XL U5408 ( .A(n3969), .B(out1_1[44]), .Z(n4032) );
  CND2XL U5409 ( .A(n3970), .B(out1_1[45]), .Z(n4031) );
  COND1XL U5410 ( .A(n4032), .B(n4030), .C(n4031), .Z(n4076) );
  CND2XL U5411 ( .A(n3971), .B(out1_1[46]), .Z(n4073) );
  CND2XL U5412 ( .A(n3972), .B(out1_1[47]), .Z(n4021) );
  COND1XL U5413 ( .A(n4073), .B(n4020), .C(n4021), .Z(n3973) );
  CANR1XL U5414 ( .A(n4076), .B(n3974), .C(n3973), .Z(n3975) );
  COND1X1 U5415 ( .A(n3976), .B(n4023), .C(n3975), .Z(n3977) );
  CANR1X2 U5416 ( .A(n7648), .B(n3978), .C(n3977), .Z(n7830) );
  CND2XL U5417 ( .A(n3979), .B(out1_1[48]), .Z(n4133) );
  CND2XL U5418 ( .A(n3980), .B(out1_1[49]), .Z(n4132) );
  COND1XL U5419 ( .A(n4133), .B(n4131), .C(n4132), .Z(n4130) );
  CND2XL U5420 ( .A(n3981), .B(out1_1[50]), .Z(n4127) );
  CND2XL U5421 ( .A(n3982), .B(out1_1[51]), .Z(n4097) );
  CND2XL U5422 ( .A(n3984), .B(out1_1[52]), .Z(n4113) );
  CND2XL U5423 ( .A(n3985), .B(out1_1[53]), .Z(n4112) );
  COND1XL U5424 ( .A(n4113), .B(n4111), .C(n4112), .Z(n4139) );
  CND2XL U5425 ( .A(n3986), .B(out1_1[54]), .Z(n4140) );
  CND2XL U5426 ( .A(n3987), .B(out1_1[55]), .Z(n4136) );
  COND1XL U5427 ( .A(n4140), .B(n4135), .C(n4136), .Z(n3988) );
  CANR1XL U5428 ( .A(n4139), .B(n3989), .C(n3988), .Z(n3990) );
  COND1X1 U5429 ( .A(n3991), .B(n4100), .C(n3990), .Z(n7827) );
  CND2X1 U5430 ( .A(n3992), .B(out1_1[56]), .Z(n4145) );
  CND2XL U5431 ( .A(n3993), .B(out1_1[57]), .Z(n4144) );
  COND1XL U5432 ( .A(n4145), .B(n4143), .C(n4144), .Z(n4118) );
  CND2XL U5433 ( .A(n3994), .B(out1_1[58]), .Z(n4116) );
  CND2XL U5434 ( .A(n3995), .B(out1_1[59]), .Z(n4009) );
  CND2XL U5435 ( .A(n3997), .B(out1_1[60]), .Z(n4060) );
  CIVX1 U5436 ( .A(n3998), .Z(n4033) );
  CND2XL U5437 ( .A(n4033), .B(n4032), .Z(n4002) );
  CIVX1 U5438 ( .A(n7649), .Z(n7656) );
  CNR2XL U5439 ( .A(n7656), .B(n4022), .Z(n4000) );
  CIVX1 U5440 ( .A(n7648), .Z(n7659) );
  COND1XL U5441 ( .A(n4022), .B(n7659), .C(n4023), .Z(n3999) );
  CANR1XL U5442 ( .A(n4000), .B(n3949), .C(n3999), .Z(n4001) );
  CEOXL U5443 ( .A(n4002), .B(n4001), .Z(n4003) );
  CMX2XL U5444 ( .A0(out1_2[44]), .A1(n4003), .S(n7846), .Z(n7891) );
  CIVXL U5445 ( .A(n4057), .Z(n4010) );
  CND2XL U5446 ( .A(n4010), .B(n4060), .Z(n4018) );
  CIVXL U5447 ( .A(n7816), .Z(n4012) );
  CND2XL U5448 ( .A(n7817), .B(n4012), .Z(n4014) );
  CNR2XL U5449 ( .A(n7818), .B(n4014), .Z(n4016) );
  CIVXL U5450 ( .A(n7824), .Z(n4011) );
  CANR1XL U5451 ( .A(n4012), .B(n7827), .C(n4011), .Z(n4013) );
  COND1XL U5452 ( .A(n4014), .B(n7830), .C(n4013), .Z(n4015) );
  CANR1XL U5453 ( .A(n4016), .B(n3949), .C(n4015), .Z(n4017) );
  CEOXL U5454 ( .A(n4018), .B(n4017), .Z(n4019) );
  CMX2XL U5455 ( .A0(out1_2[60]), .A1(n4019), .S(n8022), .Z(n7875) );
  CIVXL U5456 ( .A(n4022), .Z(n4075) );
  CIVXL U5457 ( .A(n4023), .Z(n4077) );
  CIVXL U5458 ( .A(n4026), .Z(n4044) );
  CND2XL U5459 ( .A(n4044), .B(n4029), .Z(n4039) );
  CIVXL U5460 ( .A(n4027), .Z(n4043) );
  CANR1XL U5461 ( .A(n4029), .B(n4043), .C(n4028), .Z(n4040) );
  CIVXL U5462 ( .A(n4036), .Z(n7654) );
  CIVXL U5463 ( .A(n4134), .Z(n4047) );
  CND2XL U5464 ( .A(n4047), .B(n4133), .Z(n4051) );
  CIVXL U5465 ( .A(n7818), .Z(n4049) );
  CIVXL U5466 ( .A(n7830), .Z(n4048) );
  CANR1XL U5467 ( .A(n4049), .B(n3949), .C(n4048), .Z(n4050) );
  CEOXL U5468 ( .A(n4051), .B(n4050), .Z(n4052) );
  CMX2XL U5469 ( .A0(out1_2[48]), .A1(n4052), .S(n8022), .Z(n7887) );
  CANR2XL U5470 ( .A(n4054), .B(out0_2[62]), .C(out1_2[62]), .D(n4053), .Z(
        n4055) );
  COND1XL U5471 ( .A(n7939), .B(n7810), .C(n4055), .Z(n4056) );
  COR2X1 U5472 ( .A(n4056), .B(out1_1[62]), .Z(n7822) );
  CND2XL U5473 ( .A(n4056), .B(out1_1[62]), .Z(n7819) );
  CND2XL U5474 ( .A(n7822), .B(n7819), .Z(n4070) );
  CNR2XL U5475 ( .A(n4057), .B(n4059), .Z(n7815) );
  CIVXL U5476 ( .A(n7815), .Z(n4062) );
  CNR2XL U5477 ( .A(n7816), .B(n4062), .Z(n4064) );
  CND2XL U5478 ( .A(n7817), .B(n4064), .Z(n4066) );
  CNR2XL U5479 ( .A(n7818), .B(n4066), .Z(n4068) );
  COND1XL U5480 ( .A(n4060), .B(n4059), .C(n4058), .Z(n7821) );
  CIVXL U5481 ( .A(n7821), .Z(n4061) );
  COND1XL U5482 ( .A(n4062), .B(n7824), .C(n4061), .Z(n4063) );
  CANR1XL U5483 ( .A(n4064), .B(n7827), .C(n4063), .Z(n4065) );
  COND1XL U5484 ( .A(n4066), .B(n7830), .C(n4065), .Z(n4067) );
  CANR1XL U5485 ( .A(n4068), .B(n3949), .C(n4067), .Z(n4069) );
  CEOXL U5486 ( .A(n4070), .B(n4069), .Z(n4071) );
  CMX2XL U5487 ( .A0(out1_2[62]), .A1(n4071), .S(n8022), .Z(n7873) );
  CIVXL U5488 ( .A(n4072), .Z(n4074) );
  CND2XL U5489 ( .A(n4074), .B(n4073), .Z(n4084) );
  CND2XL U5490 ( .A(n4075), .B(n4078), .Z(n4080) );
  CNR2XL U5491 ( .A(n7656), .B(n4080), .Z(n4082) );
  CANR1XL U5492 ( .A(n4078), .B(n4077), .C(n4076), .Z(n4079) );
  COND1XL U5493 ( .A(n4080), .B(n7659), .C(n4079), .Z(n4081) );
  CANR1XL U5494 ( .A(n4082), .B(n3949), .C(n4081), .Z(n4083) );
  CEOXL U5495 ( .A(n4084), .B(n4083), .Z(n4085) );
  CMX2XL U5496 ( .A0(out1_2[46]), .A1(n4085), .S(n8022), .Z(n7889) );
  CIVXL U5497 ( .A(n4086), .Z(n6388) );
  CIVXL U5498 ( .A(n4141), .Z(n4088) );
  CND2XL U5499 ( .A(n4088), .B(n4140), .Z(n4094) );
  CIVXL U5500 ( .A(n4101), .Z(n4138) );
  CND2XL U5501 ( .A(n4138), .B(n4137), .Z(n4090) );
  CNR2XL U5502 ( .A(n7818), .B(n4090), .Z(n4092) );
  CIVXL U5503 ( .A(n4100), .Z(n4142) );
  CANR1XL U5504 ( .A(n4137), .B(n4142), .C(n4139), .Z(n4089) );
  COND1XL U5505 ( .A(n4090), .B(n7830), .C(n4089), .Z(n4091) );
  CANR1XL U5506 ( .A(n4092), .B(n3949), .C(n4091), .Z(n4093) );
  CEOXL U5507 ( .A(n4094), .B(n4093), .Z(n4095) );
  CMX2XL U5508 ( .A0(out1_2[54]), .A1(n4095), .S(n8022), .Z(n7881) );
  CIVX1 U5509 ( .A(n4098), .Z(n4128) );
  CIVX1 U5510 ( .A(n4099), .Z(n4114) );
  CND2XL U5511 ( .A(n4114), .B(n4113), .Z(n4105) );
  CNR2XL U5512 ( .A(n7818), .B(n4101), .Z(n4103) );
  COND1XL U5513 ( .A(n4101), .B(n7830), .C(n4100), .Z(n4102) );
  CANR1XL U5514 ( .A(n4103), .B(n3949), .C(n4102), .Z(n4104) );
  CEOXL U5515 ( .A(n4105), .B(n4104), .Z(n4106) );
  CMX2XL U5516 ( .A0(out1_2[52]), .A1(n4106), .S(n8022), .Z(n7883) );
  CIVX1 U5517 ( .A(n4109), .Z(n4192) );
  CIVX1 U5518 ( .A(n4110), .Z(n4146) );
  CIVXL U5519 ( .A(n4115), .Z(n4117) );
  CND2XL U5520 ( .A(n4117), .B(n4116), .Z(n4125) );
  CND2XL U5521 ( .A(n7817), .B(n4119), .Z(n4121) );
  CNR2XL U5522 ( .A(n7818), .B(n4121), .Z(n4123) );
  CANR1XL U5523 ( .A(n4119), .B(n7827), .C(n4118), .Z(n4120) );
  COND1XL U5524 ( .A(n4121), .B(n7830), .C(n4120), .Z(n4122) );
  CANR1XL U5525 ( .A(n4123), .B(n3949), .C(n4122), .Z(n4124) );
  CEOXL U5526 ( .A(n4125), .B(n4124), .Z(n4126) );
  CMX2XL U5527 ( .A0(out1_2[58]), .A1(n4126), .S(n8022), .Z(n7877) );
  CIVXL U5528 ( .A(n4147), .Z(n4149) );
  CND2XL U5529 ( .A(n4149), .B(n4148), .Z(n4158) );
  CIVX1 U5530 ( .A(n7570), .Z(n7635) );
  CIVXL U5531 ( .A(n4150), .Z(n7633) );
  CND2XL U5532 ( .A(n7634), .B(n7633), .Z(n4154) );
  CNR2XL U5533 ( .A(n7635), .B(n4154), .Z(n4156) );
  CIVX2 U5534 ( .A(n4151), .Z(n7806) );
  CIVX1 U5535 ( .A(n7569), .Z(n7638) );
  CIVXL U5536 ( .A(n7632), .Z(n4152) );
  CANR1XL U5537 ( .A(n7633), .B(n7636), .C(n4152), .Z(n4153) );
  COND1XL U5538 ( .A(n4154), .B(n7638), .C(n4153), .Z(n4155) );
  CANR1XL U5539 ( .A(n4156), .B(n7806), .C(n4155), .Z(n4157) );
  CEOXL U5540 ( .A(n4158), .B(n4157), .Z(n4159) );
  CMX2XL U5541 ( .A0(out1_2[27]), .A1(n4159), .S(n7846), .Z(n7908) );
  CIVXL U5542 ( .A(n4162), .Z(n4212) );
  CIVXL U5543 ( .A(n4167), .Z(n7596) );
  CND2XL U5544 ( .A(n7596), .B(n7594), .Z(n4171) );
  CNR2XL U5545 ( .A(n7635), .B(n7592), .Z(n4169) );
  COND1XL U5546 ( .A(n7592), .B(n7638), .C(n7593), .Z(n4168) );
  CANR1XL U5547 ( .A(n4169), .B(n7806), .C(n4168), .Z(n4170) );
  CEOXL U5548 ( .A(n4171), .B(n4170), .Z(n4172) );
  CMX2XL U5549 ( .A0(out1_2[28]), .A1(n4172), .S(cmd1_en_2), .Z(n7907) );
  CIVXL U5550 ( .A(n4173), .Z(n4175) );
  CND2XL U5551 ( .A(n4175), .B(n4174), .Z(n4179) );
  CIVXL U5552 ( .A(n4176), .Z(n4182) );
  CIVXL U5553 ( .A(n4177), .Z(n4184) );
  CANR1XL U5554 ( .A(n4182), .B(n7806), .C(n4184), .Z(n4178) );
  CEOXL U5555 ( .A(n4179), .B(n4178), .Z(n4180) );
  CMX2XL U5556 ( .A0(out1_2[20]), .A1(n4180), .S(cmd1_en_2), .Z(n7915) );
  CIVXL U5557 ( .A(n4201), .Z(n4181) );
  CND2XL U5558 ( .A(n4181), .B(n4199), .Z(n4189) );
  CND2XL U5559 ( .A(n4182), .B(n4185), .Z(n4198) );
  CIVXL U5560 ( .A(n4198), .Z(n4187) );
  CANR1XL U5561 ( .A(n4185), .B(n4184), .C(n4183), .Z(n4200) );
  CIVXL U5562 ( .A(n4200), .Z(n4186) );
  CANR1XL U5563 ( .A(n4187), .B(n7806), .C(n4186), .Z(n4188) );
  CEOXL U5564 ( .A(n4189), .B(n4188), .Z(n4190) );
  CMX2XL U5565 ( .A0(out1_2[22]), .A1(n4190), .S(cmd1_en_2), .Z(n7913) );
  CND2X1 U5566 ( .A(n4192), .B(n4191), .Z(n4193) );
  CENX1 U5567 ( .A(n3949), .B(n4193), .Z(n4194) );
  CMX2XL U5568 ( .A0(out1_2[32]), .A1(n4194), .S(cmd1_en_2), .Z(n7903) );
  CIVXL U5569 ( .A(n4195), .Z(n4197) );
  CND2XL U5570 ( .A(n4197), .B(n4196), .Z(n4205) );
  CNR2XL U5571 ( .A(n4198), .B(n4201), .Z(n4203) );
  COND1XL U5572 ( .A(n4201), .B(n4200), .C(n4199), .Z(n4202) );
  CANR1XL U5573 ( .A(n4203), .B(n7806), .C(n4202), .Z(n4204) );
  CEOXL U5574 ( .A(n4205), .B(n4204), .Z(n4206) );
  CMX2XL U5575 ( .A0(out1_2[23]), .A1(n4206), .S(cmd1_en_2), .Z(n7912) );
  CIVX2 U5576 ( .A(n4207), .Z(n7792) );
  CIVXL U5577 ( .A(n4217), .Z(n4227) );
  CIVXL U5578 ( .A(n4216), .Z(n4231) );
  CIVX1 U5579 ( .A(n4210), .Z(n4223) );
  CIVX1 U5580 ( .A(n4213), .Z(n4219) );
  CIVX1 U5581 ( .A(n4240), .Z(n4275) );
  CIVXL U5582 ( .A(n7726), .Z(n7541) );
  CNR2X1 U5583 ( .A(n7541), .B(n8016), .Z(n7780) );
  CANR2XL U5584 ( .A(n7700), .B(n7780), .C(out2_2[31]), .D(n7751), .Z(n4242)
         );
  CIVX1 U5585 ( .A(n7742), .Z(n7704) );
  CND2XL U5586 ( .A(n7699), .B(n7704), .Z(n4241) );
  COND3XL U5587 ( .A(n4275), .B(n7722), .C(n4242), .D(n4241), .Z(n851) );
  CANR2XL U5588 ( .A(n4244), .B(n7582), .C(n7755), .D(n4243), .Z(n4248) );
  CANR2XL U5589 ( .A(n7747), .B(n4246), .C(n7762), .D(n4245), .Z(n4247) );
  CND2XL U5590 ( .A(n4248), .B(n4247), .Z(n7547) );
  CANR2XL U5591 ( .A(n4252), .B(n4251), .C(n4250), .D(n4249), .Z(n4259) );
  COND1XL U5592 ( .A(n4254), .B(n4253), .C(n8019), .Z(n4255) );
  CANR1XL U5593 ( .A(n4257), .B(n4256), .C(n4255), .Z(n4258) );
  COND3XL U5594 ( .A(n7727), .B(n7547), .C(n4259), .D(n4258), .Z(n4269) );
  CANR2XL U5595 ( .A(n7582), .B(n4261), .C(n7755), .D(n4260), .Z(n4265) );
  CANR2XL U5596 ( .A(n7747), .B(n4263), .C(n7762), .D(n4262), .Z(n4264) );
  CND2XL U5597 ( .A(n4265), .B(n4264), .Z(n7717) );
  COND2XL U5598 ( .A(n4267), .B(n7716), .C(n4266), .D(n7717), .Z(n4268) );
  COND2XL U5599 ( .A(n2865), .B(n4270), .C(n4269), .D(n4268), .Z(n855) );
  CANR2XL U5600 ( .A(n4271), .B(n7738), .C(n7780), .D(n7699), .Z(n4274) );
  CND2X1 U5601 ( .A(n4272), .B(n8019), .Z(n7565) );
  CIVX1 U5602 ( .A(n7565), .Z(n7778) );
  CANR2XL U5603 ( .A(n7700), .B(n7778), .C(out2_2[15]), .D(n7751), .Z(n4273)
         );
  COND3XL U5604 ( .A(n4275), .B(n7742), .C(n4274), .D(n4273), .Z(n852) );
  CNIVX1 U5605 ( .A(out0_2[22]), .Z(n4368) );
  CIVX1 U5606 ( .A(n4281), .Z(n4324) );
  CNR2X1 U5607 ( .A(n4324), .B(n7953), .Z(n4282) );
  CENX1 U5608 ( .A(n4282), .B(n7951), .Z(n4283) );
  CND2XL U5609 ( .A(n4283), .B(n4344), .Z(n4285) );
  CANR2XL U5610 ( .A(n4363), .B(out1_2[56]), .C(acc[56]), .D(n4350), .Z(n4284)
         );
  CNR2X1 U5611 ( .A(n4286), .B(n7990), .Z(n4287) );
  CENX1 U5612 ( .A(n4287), .B(n7989), .Z(n4288) );
  CND2XL U5613 ( .A(n4288), .B(n4344), .Z(n4290) );
  CANR2XL U5614 ( .A(n4363), .B(out1_2[34]), .C(acc[34]), .D(n4350), .Z(n4289)
         );
  COND3XL U5615 ( .A(n2685), .B(n2642), .C(n4290), .D(n4289), .Z(n1027) );
  CNR2X1 U5616 ( .A(n4343), .B(n7983), .Z(n4294) );
  CENX1 U5617 ( .A(n4294), .B(n7981), .Z(n4295) );
  CND2XL U5618 ( .A(n4295), .B(n4344), .Z(n4297) );
  CANR2XL U5619 ( .A(n4363), .B(out1_2[38]), .C(acc[38]), .D(n4350), .Z(n4296)
         );
  CIVX1 U5620 ( .A(n4298), .Z(n4333) );
  CNR2X1 U5621 ( .A(n4333), .B(n7987), .Z(n4299) );
  CENX1 U5622 ( .A(n4299), .B(n7985), .Z(n4300) );
  CND2XL U5623 ( .A(n4300), .B(n4344), .Z(n4302) );
  CANR2XL U5624 ( .A(n4363), .B(out1_2[36]), .C(acc[36]), .D(n4350), .Z(n4301)
         );
  CNR2X1 U5625 ( .A(n4303), .B(n7974), .Z(n4304) );
  CENX1 U5626 ( .A(n4304), .B(n7972), .Z(n4305) );
  CND2XL U5627 ( .A(n4305), .B(n4344), .Z(n4307) );
  CANR2XL U5628 ( .A(n4363), .B(out1_2[44]), .C(acc[44]), .D(n4350), .Z(n4306)
         );
  COND3XL U5629 ( .A(n2685), .B(n2645), .C(n4307), .D(n4306), .Z(n1037) );
  CNR2X1 U5630 ( .A(n4309), .B(n4308), .Z(n4311) );
  CENX1 U5631 ( .A(n4311), .B(n4310), .Z(n4312) );
  CND2XL U5632 ( .A(n4312), .B(n4344), .Z(n4314) );
  CANR2XL U5633 ( .A(n4363), .B(out1_2[28]), .C(acc[28]), .D(n4350), .Z(n4313)
         );
  COND3XL U5634 ( .A(n2685), .B(n2646), .C(n4314), .D(n4313), .Z(n1021) );
  CNIVX1 U5635 ( .A(out0_2[26]), .Z(n4371) );
  CEOXL U5636 ( .A(n7995), .B(n4319), .Z(n4320) );
  CND2XL U5637 ( .A(n4320), .B(n4344), .Z(n4322) );
  CANR2XL U5638 ( .A(n4363), .B(out1_2[29]), .C(acc[29]), .D(n4350), .Z(n4321)
         );
  COND3XL U5639 ( .A(n2655), .B(n2685), .C(n4322), .D(n4321), .Z(n1022) );
  CEOXL U5640 ( .A(n7953), .B(n4324), .Z(n4325) );
  CND2XL U5641 ( .A(n4325), .B(n4344), .Z(n4327) );
  CANR2XL U5642 ( .A(n4363), .B(out1_2[55]), .C(acc[55]), .D(n4350), .Z(n4326)
         );
  COND3XL U5643 ( .A(n2685), .B(n2648), .C(n4327), .D(n4326), .Z(n1048) );
  CNIVX1 U5644 ( .A(out0_2[41]), .Z(n4387) );
  CIVXL U5645 ( .A(n1368), .Z(n4332) );
  CEOXL U5646 ( .A(n7977), .B(n4328), .Z(n4329) );
  CND2XL U5647 ( .A(n4329), .B(n4344), .Z(n4331) );
  CANR2XL U5648 ( .A(n4363), .B(out1_2[41]), .C(acc[41]), .D(n4350), .Z(n4330)
         );
  COND3XL U5649 ( .A(n2685), .B(n4332), .C(n4331), .D(n4330), .Z(n1034) );
  CNIVX1 U5650 ( .A(out0_2[35]), .Z(n4388) );
  CIVXL U5651 ( .A(n1375), .Z(n4337) );
  CEOXL U5652 ( .A(n7987), .B(n4333), .Z(n4334) );
  CND2XL U5653 ( .A(n4334), .B(n4344), .Z(n4336) );
  CANR2XL U5654 ( .A(n4363), .B(out1_2[35]), .C(acc[35]), .D(n4350), .Z(n4335)
         );
  COND3XL U5655 ( .A(n2685), .B(n4337), .C(n4336), .D(n4335), .Z(n1028) );
  CNIVX1 U5656 ( .A(out0_2[47]), .Z(n4385) );
  CIVXL U5657 ( .A(n1366), .Z(n4342) );
  CEOXL U5658 ( .A(n7968), .B(n4338), .Z(n4339) );
  CND2XL U5659 ( .A(n4339), .B(n4344), .Z(n4341) );
  CANR2XL U5660 ( .A(n4363), .B(out1_2[47]), .C(acc[47]), .D(n4350), .Z(n4340)
         );
  COND3XL U5661 ( .A(n2685), .B(n4342), .C(n4341), .D(n4340), .Z(n1040) );
  CEOXL U5662 ( .A(n7983), .B(n4343), .Z(n4345) );
  CND2XL U5663 ( .A(n4345), .B(n4344), .Z(n4347) );
  CANR2XL U5664 ( .A(n4363), .B(out1_2[37]), .C(acc[37]), .D(n4350), .Z(n4346)
         );
  CEOXL U5665 ( .A(n7961), .B(n4348), .Z(n4349) );
  CND2XL U5666 ( .A(n4349), .B(n4344), .Z(n4352) );
  CANR2XL U5667 ( .A(n4363), .B(out1_2[51]), .C(acc[51]), .D(n4350), .Z(n4351)
         );
  CNIVX1 U5668 ( .A(out0_2[31]), .Z(n4369) );
  CIVXL U5669 ( .A(n1371), .Z(n4357) );
  CENX1 U5670 ( .A(n4353), .B(n7994), .Z(n4354) );
  CND2XL U5671 ( .A(n4354), .B(n4344), .Z(n4356) );
  CANR2XL U5672 ( .A(n4363), .B(out1_2[31]), .C(acc[31]), .D(n4350), .Z(n4355)
         );
  COND3XL U5673 ( .A(n4357), .B(n2685), .C(n4356), .D(n4355), .Z(n1024) );
  CIVX2 U5674 ( .A(q0[23]), .Z(n4534) );
  CIVX3 U5675 ( .A(n7867), .Z(n6460) );
  CNIVX4 U5676 ( .A(q0[26]), .Z(n4686) );
  CIVXL U5677 ( .A(n7871), .Z(n4367) );
  CMX2XL U5678 ( .A0(out0_2[20]), .A1(out1_1[20]), .S(cmd0_en_2), .Z(n1164) );
  CMX2XL U5679 ( .A0(n1387), .A1(out1_1[22]), .S(cmd0_en_2), .Z(n1162) );
  CMX2XL U5680 ( .A0(out0_2[21]), .A1(out1_1[21]), .S(cmd0_en_2), .Z(n1163) );
  CMX2XL U5681 ( .A0(n1371), .A1(out1_1[31]), .S(cmd0_en_2), .Z(n1153) );
  CMX2XL U5682 ( .A0(out0_2[30]), .A1(out1_1[30]), .S(cmd0_en_2), .Z(n1154) );
  CMX2XL U5683 ( .A0(out0_2[29]), .A1(out1_1[29]), .S(cmd0_en_2), .Z(n1155) );
  CMX2XL U5684 ( .A0(out0_2[28]), .A1(out1_1[28]), .S(cmd0_en_2), .Z(n1156) );
  CMX2XL U5685 ( .A0(n1372), .A1(out1_1[27]), .S(cmd0_en_2), .Z(n1157) );
  CMX2XL U5686 ( .A0(n1373), .A1(out1_1[26]), .S(cmd0_en_2), .Z(n1158) );
  CMX2XL U5687 ( .A0(n1377), .A1(out1_1[25]), .S(cmd0_en_2), .Z(n1159) );
  CMX2XL U5688 ( .A0(n1388), .A1(out1_1[23]), .S(cmd0_en_2), .Z(n1161) );
  CMX2XL U5689 ( .A0(n1374), .A1(out1_1[19]), .S(cmd0_en_2), .Z(n1165) );
  CMX2XL U5690 ( .A0(n4375), .A1(out1_1[7]), .S(cmd0_en_2), .Z(n1177) );
  CMX2XL U5691 ( .A0(n4376), .A1(out1_1[6]), .S(cmd0_en_2), .Z(n1178) );
  CMX2XL U5692 ( .A0(n4377), .A1(out1_1[5]), .S(cmd0_en_2), .Z(n1179) );
  CMX2XL U5693 ( .A0(h0[1]), .A1(h[1]), .S(n7682), .Z(n920) );
  CMX2XL U5694 ( .A0(n4378), .A1(out1_1[4]), .S(cmd0_en_2), .Z(n1180) );
  CMX2XL U5695 ( .A0(n4379), .A1(out1_1[3]), .S(cmd0_en_2), .Z(n1181) );
  CMX2XL U5696 ( .A0(out0_2[18]), .A1(out1_1[18]), .S(cmd0_en_2), .Z(n1166) );
  CMX2XL U5697 ( .A0(out0_2[17]), .A1(out1_1[17]), .S(cmd0_en_2), .Z(n1167) );
  CMX2XL U5698 ( .A0(out0_2[16]), .A1(out1_1[16]), .S(cmd0_en_2), .Z(n1168) );
  CMX2XL U5699 ( .A0(n4380), .A1(out1_1[15]), .S(cmd0_en_2), .Z(n1169) );
  CMX2XL U5700 ( .A0(n1376), .A1(out1_1[14]), .S(cmd0_en_2), .Z(n1170) );
  CMX2XL U5701 ( .A0(n4382), .A1(out1_1[13]), .S(cmd0_en_2), .Z(n1171) );
  CMX2XL U5702 ( .A0(n4383), .A1(out1_1[12]), .S(cmd0_en_2), .Z(n1172) );
  CMX2XL U5703 ( .A0(n4384), .A1(out1_1[11]), .S(cmd0_en_2), .Z(n1173) );
  CMX2XL U5704 ( .A0(cmd1_en_1), .A1(n8022), .S(rst), .Z(n1187) );
  CMX2XL U5705 ( .A0(n1366), .A1(out1_1[47]), .S(cmd0_en_2), .Z(n1137) );
  CMX2XL U5706 ( .A0(out0_2[45]), .A1(out1_1[45]), .S(cmd0_en_2), .Z(n1139) );
  CMX2XL U5707 ( .A0(out0_2[44]), .A1(out1_1[44]), .S(cmd0_en_2), .Z(n1140) );
  CMX2XL U5708 ( .A0(n1367), .A1(out1_1[43]), .S(cmd0_en_2), .Z(n1141) );
  CMX2XL U5709 ( .A0(n1368), .A1(out1_1[41]), .S(cmd0_en_2), .Z(n1143) );
  CMX2XL U5710 ( .A0(out0_2[34]), .A1(out1_1[34]), .S(cmd0_en_2), .Z(n1150) );
  CMX2XL U5711 ( .A0(out0_2[38]), .A1(out1_1[38]), .S(cmd0_en_2), .Z(n1146) );
  CMX2XL U5712 ( .A0(out0_2[37]), .A1(out1_1[37]), .S(cmd0_en_2), .Z(n1147) );
  CMX2XL U5713 ( .A0(n1375), .A1(out1_1[35]), .S(cmd0_en_2), .Z(n1149) );
  CMX2XL U5714 ( .A0(out0_2[39]), .A1(out1_1[39]), .S(cmd0_en_2), .Z(n1145) );
  CENX1 U5715 ( .A(n6491), .B(n6185), .Z(n4389) );
  CENX1 U5716 ( .A(h0[17]), .B(n5793), .Z(n4488) );
  CENX1 U5717 ( .A(n5793), .B(h0[18]), .Z(n4480) );
  COND2X1 U5718 ( .A(n5911), .B(n4488), .C(n5912), .D(n4480), .Z(n4413) );
  CENX1 U5719 ( .A(n2660), .B(h0[7]), .Z(n4485) );
  COND2X1 U5720 ( .A(n6703), .B(n4485), .C(n2515), .D(n4479), .Z(n4412) );
  CENX1 U5721 ( .A(n6491), .B(h0[8]), .Z(n4444) );
  COND2X1 U5722 ( .A(n6527), .B(n4444), .C(n1557), .D(n4389), .Z(n4454) );
  CIVX2 U5723 ( .A(n4396), .Z(n4391) );
  CIVX4 U5724 ( .A(n4391), .Z(n5155) );
  CIVX8 U5725 ( .A(n5155), .Z(n6972) );
  CNR2IX1 U5726 ( .B(n7539), .A(n6972), .Z(n4439) );
  CENX1 U5727 ( .A(n6409), .B(n2512), .Z(n4417) );
  COND2X2 U5728 ( .A(n6766), .B(n4392), .C(n6765), .D(n4417), .Z(n4441) );
  COND2X1 U5729 ( .A(n7537), .B(n4495), .C(n4393), .D(n5160), .Z(n4438) );
  CND2X2 U5730 ( .A(n4395), .B(n4394), .Z(n4452) );
  CIVX2 U5731 ( .A(n4396), .Z(n6639) );
  CIVX2 U5732 ( .A(q0[21]), .Z(n4397) );
  CENX1 U5733 ( .A(n4397), .B(n2464), .Z(n4663) );
  CND2X4 U5734 ( .A(n6639), .B(n4663), .Z(n6974) );
  CENX1 U5735 ( .A(n5932), .B(h0[1]), .Z(n4403) );
  COND2X1 U5736 ( .A(n6974), .B(n4398), .C(n6972), .D(n4403), .Z(n4484) );
  CND2X1 U5737 ( .A(n4399), .B(n5932), .Z(n4400) );
  COND2X1 U5738 ( .A(n6974), .B(n4397), .C(n4400), .D(n6972), .Z(n4483) );
  COND1X2 U5739 ( .A(n4454), .B(n4452), .C(n4453), .Z(n4402) );
  CND2X2 U5740 ( .A(n4452), .B(n4454), .Z(n4401) );
  CENX1 U5741 ( .A(n6409), .B(n7674), .Z(n4481) );
  CENX1 U5742 ( .A(n6409), .B(h0[5]), .Z(n4418) );
  COND2X1 U5743 ( .A(n6765), .B(n4481), .C(n4418), .D(n1582), .Z(n4472) );
  CENX1 U5744 ( .A(n5932), .B(h0[2]), .Z(n4531) );
  COND2X1 U5745 ( .A(n6974), .B(n4403), .C(n4531), .D(n6972), .Z(n4470) );
  CENXL U5746 ( .A(h0[19]), .B(n5566), .Z(n4493) );
  CENXL U5747 ( .A(h0[20]), .B(n5566), .Z(n4476) );
  COND2X1 U5748 ( .A(n5695), .B(n4493), .C(n4886), .D(n4476), .Z(n4471) );
  CENX1 U5749 ( .A(n4470), .B(n4471), .Z(n4404) );
  COND1X2 U5750 ( .A(n4464), .B(n4465), .C(n4466), .Z(n4406) );
  CND2X2 U5751 ( .A(n4406), .B(n4405), .Z(n5450) );
  CENX1 U5752 ( .A(n5923), .B(h0[16]), .Z(n4533) );
  COR2X1 U5753 ( .A(n3368), .B(n4533), .Z(n4408) );
  CENX1 U5754 ( .A(n5923), .B(h0[15]), .Z(n4487) );
  CND2X2 U5755 ( .A(n4407), .B(n4408), .Z(n4424) );
  CENX1 U5756 ( .A(h0[13]), .B(n6118), .Z(n4416) );
  CENX1 U5757 ( .A(h0[14]), .B(n4922), .Z(n4540) );
  COND2X1 U5758 ( .A(n2565), .B(n4416), .C(n2491), .D(n4540), .Z(n4426) );
  CENX1 U5759 ( .A(n6417), .B(h0[11]), .Z(n4490) );
  CENX1 U5760 ( .A(h0[12]), .B(n6417), .Z(n4530) );
  COND2X1 U5761 ( .A(n6522), .B(n4490), .C(n5984), .D(n4530), .Z(n4423) );
  COND1X2 U5762 ( .A(n4424), .B(n4426), .C(n4423), .Z(n4410) );
  CND2X2 U5763 ( .A(n4426), .B(n4424), .Z(n4409) );
  CND2X2 U5764 ( .A(n4410), .B(n4409), .Z(n5414) );
  CNR2IX1 U5765 ( .B(n7539), .A(n7114), .Z(n4429) );
  CIVX2 U5766 ( .A(n2280), .Z(n4411) );
  CENX1 U5767 ( .A(n4861), .B(h0[22]), .Z(n4475) );
  COND2X1 U5768 ( .A(n5160), .B(n4496), .C(n7537), .D(n4475), .Z(n4428) );
  CENXL U5769 ( .A(n6828), .B(h0[3]), .Z(n4422) );
  CENXL U5770 ( .A(n6828), .B(n2511), .Z(n4532) );
  COND2X1 U5771 ( .A(n6870), .B(n4422), .C(n6770), .D(n4532), .Z(n4427) );
  CFA1X1 U5772 ( .A(n4414), .B(n4413), .CI(n4412), .CO(n5415), .S(n4464) );
  CENX2 U5773 ( .A(n5414), .B(n4415), .Z(n5449) );
  CENX1 U5774 ( .A(h0[12]), .B(n6191), .Z(n4519) );
  COND2X1 U5775 ( .A(n2564), .B(n4519), .C(n2489), .D(n4416), .Z(n4504) );
  COND2X1 U5776 ( .A(n6765), .B(n4418), .C(n4417), .D(n6766), .Z(n4503) );
  CND2X1 U5777 ( .A(n4421), .B(n4420), .Z(n6831) );
  CENX1 U5778 ( .A(n6769), .B(h0[2]), .Z(n4436) );
  COND2X1 U5779 ( .A(n6831), .B(n4436), .C(n6770), .D(n4422), .Z(n4502) );
  CENX2 U5780 ( .A(n4424), .B(n4423), .Z(n4425) );
  CENX2 U5781 ( .A(n4426), .B(n4425), .Z(n4432) );
  CFA1X1 U5782 ( .A(n4429), .B(n4428), .CI(n4427), .CO(n5416), .S(n4431) );
  CENX2 U5783 ( .A(n5450), .B(n4430), .Z(n5484) );
  CENXL U5784 ( .A(h0[18]), .B(n5104), .Z(n4494) );
  COND2X1 U5785 ( .A(n5695), .B(n4434), .C(n5696), .D(n4494), .Z(n4513) );
  COND2X1 U5786 ( .A(n6703), .B(n4435), .C(n2514), .D(n4486), .Z(n4512) );
  COND2X1 U5787 ( .A(n2420), .B(n4437), .C(n6770), .D(n4436), .Z(n4511) );
  CENX1 U5788 ( .A(n4439), .B(n4438), .Z(n4440) );
  CENX2 U5789 ( .A(n4441), .B(n4440), .Z(n4601) );
  CND2X1 U5790 ( .A(n4598), .B(n4601), .Z(n4451) );
  CENX1 U5791 ( .A(h0[16]), .B(n5793), .Z(n4489) );
  COND2X1 U5792 ( .A(n4443), .B(n4442), .C(n5912), .D(n4489), .Z(n4522) );
  CIVX2 U5793 ( .A(n4522), .Z(n4449) );
  COND2X1 U5794 ( .A(n2449), .B(n4445), .C(n1556), .D(n4444), .Z(n4520) );
  CENX1 U5795 ( .A(n6417), .B(h0[10]), .Z(n4491) );
  COND2X1 U5796 ( .A(n6523), .B(n4491), .C(n6211), .D(n4446), .Z(n4521) );
  CENXL U5797 ( .A(n4520), .B(n4521), .Z(n4447) );
  CIVX1 U5798 ( .A(n4447), .Z(n4448) );
  CENX2 U5799 ( .A(n4449), .B(n4448), .Z(n4599) );
  COND1X2 U5800 ( .A(n4598), .B(n4601), .C(n4599), .Z(n4450) );
  CND2X2 U5801 ( .A(n4451), .B(n4450), .Z(n4585) );
  CEO3X2 U5802 ( .A(n4454), .B(n4453), .C(n4452), .Z(n4583) );
  CFA1X1 U5803 ( .A(n4457), .B(n4456), .CI(n4455), .CO(n4592), .S(n4594) );
  CFA1X1 U5804 ( .A(n4461), .B(n4460), .CI(n4459), .CO(n4590), .S(n4558) );
  COND1X2 U5805 ( .A(n4585), .B(n4583), .C(n4582), .Z(n4463) );
  CND2X2 U5806 ( .A(n4463), .B(n4462), .Z(n4552) );
  CENX2 U5807 ( .A(n4465), .B(n4464), .Z(n4467) );
  CENX2 U5808 ( .A(n4467), .B(n4466), .Z(n4549) );
  CND2X2 U5809 ( .A(n4469), .B(n4468), .Z(n5483) );
  CENX2 U5810 ( .A(n5484), .B(n5483), .Z(n4544) );
  COND1X1 U5811 ( .A(n4471), .B(n4472), .C(n4470), .Z(n4474) );
  CND2X1 U5812 ( .A(n4472), .B(n4471), .Z(n4473) );
  CND2X1 U5813 ( .A(n4474), .B(n4473), .Z(n5429) );
  CENX1 U5814 ( .A(n5106), .B(h0[23]), .Z(n5159) );
  COND2X1 U5815 ( .A(n4475), .B(n5160), .C(n7537), .D(n5159), .Z(n5314) );
  COND2X1 U5816 ( .A(n5695), .B(n4476), .C(n4886), .D(n5171), .Z(n5312) );
  CENX1 U5817 ( .A(n6491), .B(h0[11]), .Z(n5195) );
  COND2X1 U5818 ( .A(n2449), .B(n4477), .C(n1557), .D(n5195), .Z(n5313) );
  CENX1 U5819 ( .A(n5314), .B(n4478), .Z(n5428) );
  COND2X1 U5820 ( .A(n6703), .B(n4479), .C(n6702), .D(n5191), .Z(n5308) );
  CENX1 U5821 ( .A(n5793), .B(h0[19]), .Z(n5182) );
  COND2X1 U5822 ( .A(n5911), .B(n4480), .C(n5912), .D(n5182), .Z(n5307) );
  CENX1 U5823 ( .A(n5308), .B(n5307), .Z(n4482) );
  CENX1 U5824 ( .A(n6699), .B(h0[7]), .Z(n5183) );
  COND2X1 U5825 ( .A(n1582), .B(n4481), .C(n6765), .D(n5183), .Z(n5309) );
  CENX1 U5826 ( .A(n4482), .B(n5309), .Z(n5427) );
  CHA1X1 U5827 ( .A(n4484), .B(n4483), .CO(n4543), .S(n4453) );
  COND2X1 U5828 ( .A(n4486), .B(n6703), .C(n2515), .D(n4485), .Z(n4501) );
  CENX1 U5829 ( .A(n5923), .B(h0[14]), .Z(n4514) );
  COND2X1 U5830 ( .A(n6114), .B(n4514), .C(n3368), .D(n4487), .Z(n4500) );
  COND2X1 U5831 ( .A(n5911), .B(n4489), .C(n5912), .D(n4488), .Z(n4499) );
  COND2X1 U5832 ( .A(n6211), .B(n4491), .C(n6523), .D(n4490), .Z(n4508) );
  COND2X1 U5833 ( .A(n5695), .B(n4494), .C(n4886), .D(n4493), .Z(n4505) );
  COND2X2 U5834 ( .A(n7537), .B(n4496), .C(n5160), .D(n4495), .Z(n4506) );
  CFA1X1 U5835 ( .A(n4500), .B(n4499), .CI(n4501), .CO(n4542), .S(n4567) );
  CFA1X1 U5836 ( .A(n4504), .B(n4503), .CI(n4502), .CO(n4433), .S(n4566) );
  CENX1 U5837 ( .A(n4508), .B(n4507), .Z(n4569) );
  COND1X1 U5838 ( .A(n4567), .B(n4566), .C(n4569), .Z(n4510) );
  CND2X1 U5839 ( .A(n4566), .B(n4567), .Z(n4509) );
  CND2X2 U5840 ( .A(n4510), .B(n4509), .Z(n4545) );
  CFA1X1 U5841 ( .A(n4513), .B(n4512), .CI(n4511), .CO(n4554), .S(n4598) );
  COND2X1 U5842 ( .A(n4959), .B(n4515), .C(n3368), .D(n4514), .Z(n4557) );
  COND1XL U5843 ( .A(n4521), .B(n4522), .C(n4520), .Z(n4525) );
  CIVXL U5844 ( .A(n4521), .Z(n4523) );
  CND2IX1 U5845 ( .B(n4523), .A(n4522), .Z(n4524) );
  CND2X1 U5846 ( .A(n4525), .B(n4524), .Z(n4553) );
  COND1X2 U5847 ( .A(n4554), .B(n4556), .C(n4553), .Z(n4527) );
  CND2X1 U5848 ( .A(n4556), .B(n4554), .Z(n4526) );
  CND2X2 U5849 ( .A(n4527), .B(n4526), .Z(n4546) );
  COND1X1 U5850 ( .A(n4548), .B(n4545), .C(n4546), .Z(n4529) );
  CND2X1 U5851 ( .A(n4545), .B(n4548), .Z(n4528) );
  CND2X2 U5852 ( .A(n4529), .B(n4528), .Z(n5474) );
  CENX1 U5853 ( .A(h0[13]), .B(n6417), .Z(n5295) );
  COND2X1 U5854 ( .A(n6418), .B(n4530), .C(n6293), .D(n5295), .Z(n5298) );
  COND2X1 U5855 ( .A(n6974), .B(n4531), .C(n6972), .D(n5157), .Z(n5297) );
  CENX1 U5856 ( .A(n6828), .B(h0[5]), .Z(n5167) );
  COND2X1 U5857 ( .A(n6870), .B(n4532), .C(n6829), .D(n5167), .Z(n5296) );
  CENX1 U5858 ( .A(n5923), .B(h0[17]), .Z(n5185) );
  COND2X1 U5859 ( .A(n4959), .B(n4533), .C(n4957), .D(n5185), .Z(n5409) );
  CNIVX4 U5860 ( .A(n4534), .Z(n4711) );
  CENX1 U5861 ( .A(n7869), .B(q0[22]), .Z(n4535) );
  CND2X1 U5862 ( .A(n4399), .B(n2659), .Z(n4536) );
  COND2X1 U5863 ( .A(n4711), .B(n2293), .C(n4536), .D(n7114), .Z(n5300) );
  CIVX1 U5864 ( .A(n5300), .Z(n4539) );
  CNIVX4 U5865 ( .A(n7869), .Z(n4537) );
  CIVX8 U5866 ( .A(n4537), .Z(n7092) );
  CENX1 U5867 ( .A(n7092), .B(n7539), .Z(n4538) );
  CENX1 U5868 ( .A(n4539), .B(n5299), .Z(n5408) );
  CENX1 U5869 ( .A(h0[15]), .B(n6191), .Z(n5193) );
  COND2X1 U5870 ( .A(n2570), .B(n4540), .C(n2488), .D(n5193), .Z(n5407) );
  CFA1X1 U5871 ( .A(n4543), .B(n4542), .CI(n4541), .CO(n5445), .S(n4548) );
  CEO3X2 U5872 ( .A(n5476), .B(n5474), .C(n5475), .Z(n5485) );
  CENX2 U5873 ( .A(n4544), .B(n5485), .Z(n4577) );
  CIVX2 U5874 ( .A(n4577), .Z(n4575) );
  CENX2 U5875 ( .A(n4546), .B(n4545), .Z(n4547) );
  CENX2 U5876 ( .A(n4548), .B(n4547), .Z(n4578) );
  CENX2 U5877 ( .A(n4550), .B(n4549), .Z(n4551) );
  CENX2 U5878 ( .A(n4552), .B(n4551), .Z(n4581) );
  CENX2 U5879 ( .A(n4554), .B(n4553), .Z(n4555) );
  CENX2 U5880 ( .A(n4556), .B(n4555), .Z(n4587) );
  CND2X1 U5881 ( .A(n4560), .B(n4559), .Z(n4561) );
  CND2X2 U5882 ( .A(n4562), .B(n4561), .Z(n4611) );
  COND1X2 U5883 ( .A(n4612), .B(n4611), .C(n4610), .Z(n4565) );
  CND2X1 U5884 ( .A(n4611), .B(n4612), .Z(n4564) );
  CND2X2 U5885 ( .A(n4565), .B(n4564), .Z(n4589) );
  CENX2 U5886 ( .A(n4569), .B(n4568), .Z(n4586) );
  CND2X2 U5887 ( .A(n4571), .B(n4570), .Z(n4579) );
  CND2X2 U5888 ( .A(n4573), .B(n4572), .Z(n4576) );
  CIVX2 U5889 ( .A(n4576), .Z(n4574) );
  CND2X2 U5890 ( .A(n4575), .B(n4574), .Z(n5396) );
  CND2X2 U5891 ( .A(n4577), .B(n4576), .Z(n5393) );
  CENX2 U5892 ( .A(n4579), .B(n4578), .Z(n4580) );
  CENX2 U5893 ( .A(n4581), .B(n4580), .Z(n4645) );
  CENX2 U5894 ( .A(n4583), .B(n4582), .Z(n4584) );
  CENX2 U5895 ( .A(n4585), .B(n4584), .Z(n4607) );
  CENX2 U5896 ( .A(n4587), .B(n4586), .Z(n4588) );
  CENX2 U5897 ( .A(n4589), .B(n4588), .Z(n4609) );
  CFA1X1 U5898 ( .A(n4592), .B(n4591), .CI(n4590), .CO(n4582), .S(n4613) );
  CND2X2 U5899 ( .A(n4597), .B(n4596), .Z(n4616) );
  CENX2 U5900 ( .A(n4599), .B(n4598), .Z(n4600) );
  CENX2 U5901 ( .A(n4601), .B(n4600), .Z(n4614) );
  COND1X2 U5902 ( .A(n4613), .B(n4616), .C(n4614), .Z(n4603) );
  CND2X2 U5903 ( .A(n4616), .B(n4613), .Z(n4602) );
  CND2X2 U5904 ( .A(n4603), .B(n4602), .Z(n4606) );
  COND1X2 U5905 ( .A(n4607), .B(n4609), .C(n4606), .Z(n4605) );
  CND2X1 U5906 ( .A(n4609), .B(n4607), .Z(n4604) );
  CND2X2 U5907 ( .A(n4605), .B(n4604), .Z(n4644) );
  CNR2X2 U5908 ( .A(n4645), .B(n4644), .Z(n4648) );
  CENX2 U5909 ( .A(n4607), .B(n4606), .Z(n4608) );
  CENX2 U5910 ( .A(n4609), .B(n4608), .Z(n4643) );
  CEO3X2 U5911 ( .A(n4612), .B(n4611), .C(n4610), .Z(n4626) );
  CENX2 U5912 ( .A(n4614), .B(n4613), .Z(n4615) );
  CENX2 U5913 ( .A(n4616), .B(n4615), .Z(n4628) );
  CND2X2 U5914 ( .A(n4621), .B(n4620), .Z(n4625) );
  CND2X2 U5915 ( .A(n4623), .B(n4622), .Z(n4642) );
  CNR2X1 U5916 ( .A(n4643), .B(n4642), .Z(n4651) );
  CNR2X2 U5917 ( .A(n4648), .B(n4651), .Z(n5392) );
  CIVX2 U5918 ( .A(n4624), .Z(n6383) );
  CND2X2 U5919 ( .A(n6383), .B(n4635), .Z(n7526) );
  CENX2 U5920 ( .A(n4626), .B(n4625), .Z(n4627) );
  CENX2 U5921 ( .A(n4628), .B(n4627), .Z(n4638) );
  CND2X2 U5922 ( .A(n4633), .B(n4632), .Z(n4637) );
  CNR2X2 U5923 ( .A(n4638), .B(n4637), .Z(n7527) );
  CNR2X1 U5924 ( .A(n7526), .B(n7527), .Z(n4641) );
  CND2X2 U5925 ( .A(n6384), .B(n4634), .Z(n4636) );
  CND2X2 U5926 ( .A(n4636), .B(n4635), .Z(n7525) );
  COND1X2 U5927 ( .A(n7527), .B(n7525), .C(n7528), .Z(n4639) );
  CANR1X2 U5928 ( .A(n4641), .B(n4640), .C(n4639), .Z(n5532) );
  CIVXL U5929 ( .A(n2284), .Z(n4657) );
  CND2X2 U5930 ( .A(n4643), .B(n4642), .Z(n4655) );
  CND2X2 U5931 ( .A(n4645), .B(n4644), .Z(n4649) );
  COND1X2 U5932 ( .A(n4655), .B(n4648), .C(n4649), .Z(n5395) );
  CANR1XL U5933 ( .A(n5392), .B(n4657), .C(n5395), .Z(n4646) );
  CENXL U5934 ( .A(n4647), .B(n4646), .Z(N38) );
  CIVXL U5935 ( .A(n4648), .Z(n4650) );
  CAN2XL U5936 ( .A(n4650), .B(n4649), .Z(n4654) );
  CIVXL U5937 ( .A(n4651), .Z(n4656) );
  CIVXL U5938 ( .A(n4655), .Z(n4652) );
  CANR1XL U5939 ( .A(n4656), .B(n4657), .C(n4652), .Z(n4653) );
  CENXL U5940 ( .A(n4654), .B(n4653), .Z(N37) );
  CENX1 U5941 ( .A(n5927), .B(n2659), .Z(n4992) );
  COND2X2 U5942 ( .A(n7114), .B(n4992), .C(n4774), .D(n2293), .Z(n5035) );
  CENX1 U5943 ( .A(n6417), .B(n2280), .Z(n5050) );
  CENX2 U5944 ( .A(q0[24]), .B(q0[23]), .Z(n4683) );
  CNIVX4 U5945 ( .A(q0[25]), .Z(n6411) );
  CENX1 U5946 ( .A(n7134), .B(h0[7]), .Z(n4990) );
  COND2X1 U5947 ( .A(n6969), .B(n4771), .C(n4990), .D(n7171), .Z(n5033) );
  CENX1 U5948 ( .A(n4660), .B(n5033), .Z(n5074) );
  CENX1 U5949 ( .A(n2597), .B(h0[19]), .Z(n4761) );
  COND2X1 U5950 ( .A(n6522), .B(n4761), .C(n6293), .D(n4661), .Z(n4695) );
  CND2XL U5951 ( .A(n4663), .B(n6639), .Z(n4665) );
  CIVX2 U5952 ( .A(n4688), .Z(n4664) );
  CND2IX2 U5953 ( .B(n4665), .A(n4664), .Z(n4666) );
  CIVX2 U5954 ( .A(n6701), .Z(n4669) );
  CIVX2 U5955 ( .A(n4699), .Z(n4668) );
  CND2X2 U5956 ( .A(n4669), .B(n4668), .Z(n4672) );
  CENX1 U5957 ( .A(h0[13]), .B(n6409), .Z(n4766) );
  CND2X2 U5958 ( .A(n4672), .B(n4671), .Z(n4705) );
  CENX1 U5959 ( .A(n6118), .B(n2279), .Z(n4738) );
  CENX1 U5960 ( .A(n6118), .B(h0[20]), .Z(n4698) );
  COND2X2 U5961 ( .A(n2491), .B(n4738), .C(n2573), .D(n4698), .Z(n4702) );
  CND2X1 U5962 ( .A(n4703), .B(n4705), .Z(n4673) );
  CND2X2 U5963 ( .A(n4674), .B(n4673), .Z(n4697) );
  CENX1 U5964 ( .A(n4679), .B(q0[28]), .Z(n4676) );
  CENX1 U5965 ( .A(h0[0]), .B(n6103), .Z(n4677) );
  COND2X2 U5966 ( .A(n4722), .B(n7124), .C(n7126), .D(n4677), .Z(n4758) );
  CND2IX1 U5967 ( .B(n7539), .A(n7090), .Z(n4678) );
  COND2X1 U5968 ( .A(n7853), .B(n7126), .C(n7124), .D(n4678), .Z(n4759) );
  CND2XL U5969 ( .A(n1259), .B(n2554), .Z(n4680) );
  CIVX2 U5970 ( .A(n4680), .Z(n4694) );
  COND1X2 U5971 ( .A(n4695), .B(n4697), .C(n4694), .Z(n4682) );
  CND2X1 U5972 ( .A(n4697), .B(n4695), .Z(n4681) );
  CENX1 U5973 ( .A(n5888), .B(h0[18]), .Z(n4739) );
  CENX1 U5974 ( .A(n6490), .B(h0[19]), .Z(n5040) );
  COND2X1 U5975 ( .A(n2449), .B(n4739), .C(n1556), .D(n5040), .Z(n5069) );
  CENX1 U5976 ( .A(h0[14]), .B(n6409), .Z(n4767) );
  CENX1 U5977 ( .A(h0[15]), .B(n6409), .Z(n5048) );
  CENX1 U5978 ( .A(n5932), .B(h0[10]), .Z(n4764) );
  CENX1 U5979 ( .A(n5932), .B(h0[11]), .Z(n4989) );
  COND2X1 U5980 ( .A(n6974), .B(n4764), .C(n6972), .D(n4989), .Z(n5067) );
  CNR2IX1 U5981 ( .B(n7538), .A(n2433), .Z(n4865) );
  CENX1 U5982 ( .A(n5106), .B(h0[27]), .Z(n4862) );
  COND2X1 U5983 ( .A(n5160), .B(n4862), .C(n7537), .D(n4710), .Z(n4864) );
  CENX1 U5984 ( .A(n6460), .B(h0[3]), .Z(n4869) );
  CENX1 U5985 ( .A(n6460), .B(n2513), .Z(n4713) );
  COND2X1 U5986 ( .A(n6969), .B(n4869), .C(n7171), .D(n4713), .Z(n4863) );
  CENX1 U5987 ( .A(h0[26]), .B(n5566), .Z(n4709) );
  COND2X1 U5988 ( .A(n4846), .B(n5695), .C(n5696), .D(n4709), .Z(n4839) );
  CENX1 U5989 ( .A(n5701), .B(h0[23]), .Z(n4854) );
  CENX1 U5990 ( .A(n5701), .B(h0[24]), .Z(n4720) );
  COND2X1 U5991 ( .A(n5911), .B(n4854), .C(n5912), .D(n4720), .Z(n4838) );
  CENX1 U5992 ( .A(q0[26]), .B(q0[25]), .Z(n4687) );
  CIVX2 U5993 ( .A(n4687), .Z(n4685) );
  CENX4 U5994 ( .A(n4686), .B(n7851), .Z(n4714) );
  CND2X4 U5995 ( .A(n7218), .B(n4714), .Z(n7217) );
  CIVX8 U5996 ( .A(n4851), .Z(n7202) );
  CENX1 U5997 ( .A(n7202), .B(h0[1]), .Z(n4852) );
  CENX1 U5998 ( .A(n7202), .B(h0[2]), .Z(n4715) );
  COND2X1 U5999 ( .A(n7205), .B(n4852), .C(n7203), .D(n4715), .Z(n4837) );
  CENX1 U6000 ( .A(n2583), .B(h0[22]), .Z(n4719) );
  CENX1 U6001 ( .A(n2279), .B(n2583), .Z(n4956) );
  COND2X2 U6002 ( .A(n3368), .B(n4719), .C(n6114), .D(n4956), .Z(n4689) );
  COND2X1 U6003 ( .A(n6974), .B(n4860), .C(n6972), .D(n4688), .Z(n4833) );
  CENX1 U6004 ( .A(n7092), .B(n7674), .Z(n4712) );
  CENX1 U6005 ( .A(n7092), .B(h0[5]), .Z(n4868) );
  COND2X1 U6006 ( .A(n7114), .B(n4712), .C(n4868), .D(n2295), .Z(n4832) );
  COND1X1 U6007 ( .A(n4689), .B(n4833), .C(n4832), .Z(n4691) );
  CIVX2 U6008 ( .A(n4689), .Z(n4834) );
  CND2X2 U6009 ( .A(n4691), .B(n4690), .Z(n4826) );
  CND2X2 U6010 ( .A(n4693), .B(n4692), .Z(n4911) );
  CENX2 U6011 ( .A(n4695), .B(n4694), .Z(n4696) );
  CENX1 U6012 ( .A(n4697), .B(n4696), .Z(n4910) );
  CENX1 U6013 ( .A(n6191), .B(h0[19]), .Z(n4855) );
  COND2X2 U6014 ( .A(n2570), .B(n4855), .C(n2490), .D(n4698), .Z(n4940) );
  CENX1 U6015 ( .A(n6409), .B(h0[11]), .Z(n4844) );
  COND2X2 U6016 ( .A(n6701), .B(n4844), .C(n6765), .D(n4699), .Z(n4942) );
  CENX1 U6017 ( .A(n5927), .B(n6769), .Z(n4845) );
  COND2X1 U6018 ( .A(n2420), .B(n4845), .C(n6770), .D(n4718), .Z(n4939) );
  CND2X2 U6019 ( .A(n4701), .B(n4700), .Z(n4818) );
  CENX2 U6020 ( .A(n4705), .B(n4704), .Z(n4824) );
  CENX1 U6021 ( .A(n6417), .B(h0[18]), .Z(n4762) );
  COND2X1 U6022 ( .A(n6211), .B(n4859), .C(n5984), .D(n4762), .Z(n4831) );
  CENX1 U6023 ( .A(n5888), .B(h0[15]), .Z(n4866) );
  CENX1 U6024 ( .A(n5888), .B(h0[16]), .Z(n4708) );
  COND2X1 U6025 ( .A(n2449), .B(n4866), .C(n1556), .D(n4708), .Z(n4830) );
  CENX1 U6026 ( .A(n6647), .B(h0[13]), .Z(n4856) );
  CENX1 U6027 ( .A(n6647), .B(h0[14]), .Z(n4757) );
  COND2X1 U6028 ( .A(n6703), .B(n4856), .C(n6702), .D(n4757), .Z(n4829) );
  COND1X1 U6029 ( .A(n4818), .B(n4824), .C(n4819), .Z(n4707) );
  CENX1 U6030 ( .A(n5888), .B(h0[17]), .Z(n4740) );
  CENXL U6031 ( .A(h0[27]), .B(n2531), .Z(n4729) );
  COND2X1 U6032 ( .A(n5695), .B(n4709), .C(n5696), .D(n4729), .Z(n4745) );
  CENX1 U6033 ( .A(n5106), .B(h0[29]), .Z(n4735) );
  CIVX8 U6034 ( .A(n4711), .Z(n6970) );
  COND2X1 U6035 ( .A(n2295), .B(n4712), .C(n7114), .D(n4773), .Z(n4749) );
  COND2X1 U6036 ( .A(n6969), .B(n4713), .C(n7171), .D(n4772), .Z(n4750) );
  CENX1 U6037 ( .A(n7202), .B(h0[3]), .Z(n4736) );
  CND2X4 U6038 ( .A(n7218), .B(n4714), .Z(n7205) );
  COND1X1 U6039 ( .A(n4750), .B(n4749), .C(n2468), .Z(n4717) );
  CND2X1 U6040 ( .A(n4750), .B(n4749), .Z(n4716) );
  COND2X1 U6041 ( .A(n6831), .B(n4718), .C(n6770), .D(n4765), .Z(n4748) );
  CENX1 U6042 ( .A(n5909), .B(h0[23]), .Z(n4775) );
  COND2X1 U6043 ( .A(n6114), .B(n4719), .C(n3368), .D(n4775), .Z(n4747) );
  CENX2 U6044 ( .A(n5701), .B(h0[25]), .Z(n4726) );
  CENX2 U6045 ( .A(n4897), .B(n4895), .Z(n4721) );
  CENX2 U6046 ( .A(n4721), .B(n4896), .Z(n4977) );
  CNIVX4 U6047 ( .A(n7126), .Z(n7252) );
  CNR2X2 U6048 ( .A(n7252), .B(n4722), .Z(n4723) );
  CIVX2 U6049 ( .A(n4723), .Z(n4725) );
  CENXL U6050 ( .A(n6103), .B(h0[2]), .Z(n4803) );
  CIVX2 U6051 ( .A(n2433), .Z(n5928) );
  CND2IX1 U6052 ( .B(n4803), .A(n5928), .Z(n4724) );
  CND2X2 U6053 ( .A(n4725), .B(n4724), .Z(n4781) );
  CIVX2 U6054 ( .A(n4781), .Z(n4734) );
  COND2X4 U6055 ( .A(n5911), .B(n4726), .C(n5912), .D(n4797), .Z(n4783) );
  CIVX2 U6056 ( .A(n5696), .Z(n4727) );
  CND2IX1 U6057 ( .B(n4887), .A(n4727), .Z(n4731) );
  CIVX2 U6058 ( .A(n5695), .Z(n4728) );
  CND2IX1 U6059 ( .B(n4729), .A(n4728), .Z(n4730) );
  CND2X2 U6060 ( .A(n4731), .B(n4730), .Z(n4782) );
  CNR2IX1 U6061 ( .B(n7539), .A(n7301), .Z(n4888) );
  CENX2 U6062 ( .A(n4861), .B(h0[30]), .Z(n4798) );
  COND2X2 U6063 ( .A(n7537), .B(n4798), .C(n5160), .D(n4735), .Z(n4889) );
  CENX1 U6064 ( .A(n7202), .B(n2513), .Z(n4802) );
  COND2X1 U6065 ( .A(n7217), .B(n4736), .C(n7203), .D(n4802), .Z(n4891) );
  CEO3X2 U6066 ( .A(n4888), .B(n4889), .C(n4891), .Z(n4902) );
  CENX1 U6067 ( .A(n4922), .B(h0[22]), .Z(n4808) );
  COND2X1 U6068 ( .A(n2567), .B(n4738), .C(n2487), .D(n4808), .Z(n4881) );
  COR2X1 U6069 ( .A(n1557), .B(n4739), .Z(n4742) );
  COR2X1 U6070 ( .A(n6576), .B(n4740), .Z(n4741) );
  CND2X2 U6071 ( .A(n4742), .B(n4741), .Z(n4879) );
  CENX1 U6072 ( .A(n6647), .B(h0[15]), .Z(n4756) );
  CENX1 U6073 ( .A(n6647), .B(h0[16]), .Z(n4796) );
  CENX2 U6074 ( .A(n4881), .B(n4743), .Z(n4901) );
  CENX2 U6075 ( .A(n4902), .B(n4901), .Z(n4744) );
  CENX2 U6076 ( .A(n4903), .B(n4744), .Z(n4975) );
  CND2X1 U6077 ( .A(n4977), .B(n4975), .Z(n4753) );
  CFA1X1 U6078 ( .A(n4747), .B(n4748), .CI(n4746), .CO(n4895), .S(n4913) );
  COND1X2 U6079 ( .A(n4977), .B(n4975), .C(n4976), .Z(n4752) );
  CND2X2 U6080 ( .A(n4753), .B(n4752), .Z(n5045) );
  CENX2 U6081 ( .A(n4755), .B(n4754), .Z(n5361) );
  COND2X1 U6082 ( .A(n6473), .B(n4757), .C(n2515), .D(n4756), .Z(n4874) );
  CIVX2 U6083 ( .A(n4758), .Z(n4760) );
  CENX1 U6084 ( .A(n4760), .B(n4759), .Z(n4873) );
  COND2X1 U6085 ( .A(n4762), .B(n6418), .C(n6523), .D(n4761), .Z(n4872) );
  COND2X2 U6086 ( .A(n4764), .B(n6972), .C(n6974), .D(n4763), .Z(n4791) );
  CENX1 U6087 ( .A(n6828), .B(h0[12]), .Z(n4807) );
  COND2X1 U6088 ( .A(n2420), .B(n4765), .C(n6829), .D(n4807), .Z(n4786) );
  CENX2 U6089 ( .A(n4791), .B(n4792), .Z(n4769) );
  COND2X1 U6090 ( .A(n6765), .B(n4767), .C(n4766), .D(n1582), .Z(n4789) );
  CNIVX1 U6091 ( .A(n4789), .Z(n4768) );
  CENX2 U6092 ( .A(n4769), .B(n4768), .Z(n4817) );
  CIVX2 U6093 ( .A(n6969), .Z(n4770) );
  CIVX2 U6094 ( .A(n4770), .Z(n4991) );
  COND2X1 U6095 ( .A(n6969), .B(n4772), .C(n7171), .D(n4771), .Z(n4780) );
  COND2X1 U6096 ( .A(n4774), .B(n7114), .C(n4773), .D(n2295), .Z(n4779) );
  CENX1 U6097 ( .A(n5909), .B(h0[24]), .Z(n4806) );
  COND2X1 U6098 ( .A(n6114), .B(n4775), .C(n3368), .D(n4806), .Z(n4778) );
  CND2X2 U6099 ( .A(n4777), .B(n4776), .Z(n5005) );
  CFA1X1 U6100 ( .A(n4780), .B(n4779), .CI(n4778), .CO(n5025), .S(n4814) );
  COND1X2 U6101 ( .A(n4783), .B(n4782), .C(n4781), .Z(n4785) );
  CIVX1 U6102 ( .A(n4786), .Z(n4788) );
  CIVX2 U6103 ( .A(n4791), .Z(n4787) );
  CND2X2 U6104 ( .A(n4788), .B(n4787), .Z(n4790) );
  CND2X2 U6105 ( .A(n4790), .B(n4789), .Z(n4794) );
  CENX2 U6106 ( .A(n5023), .B(n5024), .Z(n4795) );
  CENX2 U6107 ( .A(n5025), .B(n4795), .Z(n5007) );
  CENX2 U6108 ( .A(n5007), .B(n5005), .Z(n4813) );
  CENX1 U6109 ( .A(n6647), .B(h0[17]), .Z(n5051) );
  COND2X1 U6110 ( .A(n4796), .B(n6703), .C(n6702), .D(n5051), .Z(n5066) );
  CENX1 U6111 ( .A(n5701), .B(h0[27]), .Z(n5052) );
  COND2X1 U6112 ( .A(n5911), .B(n4797), .C(n5912), .D(n5052), .Z(n5065) );
  CENX1 U6113 ( .A(n5106), .B(h0[31]), .Z(n5046) );
  CIVDX3 U6114 ( .A(q0[31]), .Z0(n4885), .Z1(n7279) );
  CIVX12 U6115 ( .A(n4885), .Z(n7173) );
  CENX1 U6116 ( .A(n7279), .B(n7539), .Z(n4801) );
  CENX1 U6117 ( .A(q0[30]), .B(n7870), .Z(n4799) );
  CND2X4 U6118 ( .A(n2516), .B(n4799), .Z(n7228) );
  COND2X2 U6119 ( .A(n5039), .B(n2382), .C(n4801), .D(n7228), .Z(n5029) );
  CENX1 U6120 ( .A(n7202), .B(h0[5]), .Z(n5047) );
  COND2X2 U6121 ( .A(n7203), .B(n5047), .C(n7205), .D(n4802), .Z(n5030) );
  CENX2 U6122 ( .A(n5029), .B(n5030), .Z(n4805) );
  CENXL U6123 ( .A(n7090), .B(h0[3]), .Z(n5055) );
  COND2X1 U6124 ( .A(n4803), .B(n2282), .C(n2433), .D(n5055), .Z(n5028) );
  CNIVX2 U6125 ( .A(n5028), .Z(n4804) );
  CENX2 U6126 ( .A(n4805), .B(n4804), .Z(n5019) );
  CENX1 U6127 ( .A(n5909), .B(h0[25]), .Z(n4997) );
  COND2X1 U6128 ( .A(n6114), .B(n4806), .C(n3368), .D(n4997), .Z(n5060) );
  CNIVX2 U6129 ( .A(n5060), .Z(n4810) );
  CENX1 U6130 ( .A(n6828), .B(h0[13]), .Z(n5056) );
  COND2X2 U6131 ( .A(n6770), .B(n5056), .C(n4807), .D(n6870), .Z(n5061) );
  CENX1 U6132 ( .A(n6118), .B(h0[23]), .Z(n4996) );
  COND2X2 U6133 ( .A(n4996), .B(n2489), .C(n2568), .D(n4808), .Z(n5059) );
  CENX2 U6134 ( .A(n5061), .B(n5059), .Z(n4809) );
  CENX2 U6135 ( .A(n4809), .B(n4810), .Z(n5020) );
  CENX2 U6136 ( .A(n5019), .B(n5020), .Z(n4811) );
  CENX2 U6137 ( .A(n5018), .B(n4811), .Z(n5006) );
  CNIVX1 U6138 ( .A(n5006), .Z(n4812) );
  CENX2 U6139 ( .A(n4813), .B(n4812), .Z(n5012) );
  CENX2 U6140 ( .A(n4817), .B(n4816), .Z(n5371) );
  CND2X1 U6141 ( .A(n4819), .B(n4818), .Z(n4822) );
  CIVX2 U6142 ( .A(n4819), .Z(n4820) );
  CND2X2 U6143 ( .A(n4821), .B(n4822), .Z(n4823) );
  CENX2 U6144 ( .A(n4824), .B(n4823), .Z(n5081) );
  CENX2 U6145 ( .A(n4826), .B(n4825), .Z(n4827) );
  CENX2 U6146 ( .A(n4828), .B(n4827), .Z(n5083) );
  CFA1X1 U6147 ( .A(n4831), .B(n4830), .CI(n4829), .CO(n4819), .S(n5087) );
  CIVX2 U6148 ( .A(n4832), .Z(n4836) );
  CENX1 U6149 ( .A(n4834), .B(n4833), .Z(n4835) );
  CENX2 U6150 ( .A(n4836), .B(n4835), .Z(n5090) );
  CFA1X1 U6151 ( .A(n4839), .B(n4838), .CI(n4837), .CO(n4828), .S(n5088) );
  CND2X2 U6152 ( .A(n4841), .B(n4840), .Z(n5080) );
  CND2X2 U6153 ( .A(n4842), .B(n4843), .Z(n5369) );
  CENX1 U6154 ( .A(n6409), .B(h0[10]), .Z(n4950) );
  COND2X2 U6155 ( .A(n6765), .B(n4844), .C(n4950), .D(n6766), .Z(n5125) );
  CENX1 U6156 ( .A(h0[8]), .B(n6769), .Z(n4951) );
  COND2X1 U6157 ( .A(n2420), .B(n4951), .C(n6829), .D(n4845), .Z(n5127) );
  CENXL U6158 ( .A(h0[24]), .B(n5104), .Z(n4952) );
  COND2X1 U6159 ( .A(n4952), .B(n5695), .C(n4846), .D(n5696), .Z(n5124) );
  CIVX2 U6160 ( .A(n5125), .Z(n4847) );
  CND2IX1 U6161 ( .B(n4847), .A(n5127), .Z(n4848) );
  CND2X2 U6162 ( .A(n4849), .B(n4848), .Z(n4919) );
  CND2X1 U6163 ( .A(n4399), .B(n7062), .Z(n4850) );
  COND2X1 U6164 ( .A(n7217), .B(n4851), .C(n4850), .D(n7203), .Z(n4968) );
  CENX1 U6165 ( .A(n7062), .B(n7539), .Z(n4853) );
  COND2X1 U6166 ( .A(n7217), .B(n4853), .C(n7203), .D(n4852), .Z(n4969) );
  CND2X1 U6167 ( .A(n4919), .B(n4921), .Z(n4858) );
  CENX1 U6168 ( .A(n5701), .B(h0[22]), .Z(n4949) );
  CENX1 U6169 ( .A(n6118), .B(h0[18]), .Z(n4923) );
  COND2X1 U6170 ( .A(n2580), .B(n4923), .C(n2489), .D(n4855), .Z(n5129) );
  COND2X1 U6171 ( .A(n6703), .B(n4946), .C(n2515), .D(n4856), .Z(n5128) );
  COND1X2 U6172 ( .A(n4921), .B(n4919), .C(n4920), .Z(n4857) );
  CND2X2 U6173 ( .A(n4858), .B(n4857), .Z(n5086) );
  CENX1 U6174 ( .A(h0[16]), .B(n6417), .Z(n4926) );
  COND2X1 U6175 ( .A(n6522), .B(n4926), .C(n6293), .D(n4859), .Z(n4934) );
  CENX1 U6176 ( .A(n5932), .B(n7674), .Z(n4953) );
  COND2X1 U6177 ( .A(n6974), .B(n4953), .C(n2477), .D(n4860), .Z(n4933) );
  CENX1 U6178 ( .A(n4861), .B(h0[26]), .Z(n4960) );
  COND2X1 U6179 ( .A(n5160), .B(n4960), .C(n7537), .D(n4862), .Z(n4932) );
  CENX1 U6180 ( .A(n5888), .B(h0[14]), .Z(n4943) );
  COND2X1 U6181 ( .A(n2449), .B(n4943), .C(n1556), .D(n4866), .Z(n4931) );
  CIVX2 U6182 ( .A(n2293), .Z(n4867) );
  COND2X2 U6183 ( .A(n7114), .B(n4868), .C(n7095), .D(n1263), .Z(n4930) );
  COND2X1 U6184 ( .A(n6969), .B(n4954), .C(n7171), .D(n4869), .Z(n4929) );
  CND2X2 U6185 ( .A(n4917), .B(n4916), .Z(n4870) );
  CND2X2 U6186 ( .A(n4871), .B(n4870), .Z(n5084) );
  CND2X2 U6187 ( .A(n4876), .B(n4875), .Z(n5370) );
  COND1X2 U6188 ( .A(n5369), .B(n5371), .C(n5370), .Z(n4878) );
  CND2X2 U6189 ( .A(n4878), .B(n4877), .Z(n5014) );
  COND1X1 U6190 ( .A(n4881), .B(n4880), .C(n4879), .Z(n4883) );
  CND2X2 U6191 ( .A(n4883), .B(n4882), .Z(n4985) );
  CND2X1 U6192 ( .A(n4399), .B(n7279), .Z(n4884) );
  COND2X1 U6193 ( .A(n7228), .B(n4885), .C(n4884), .D(n2381), .Z(n4995) );
  CENX1 U6194 ( .A(h0[29]), .B(n5104), .Z(n5054) );
  COND2X1 U6195 ( .A(n5695), .B(n4887), .C(n4886), .D(n5054), .Z(n4994) );
  CNIVX1 U6196 ( .A(n4888), .Z(n4890) );
  COND1X1 U6197 ( .A(n4890), .B(n4891), .C(n4889), .Z(n4893) );
  CND2X2 U6198 ( .A(n4893), .B(n4892), .Z(n4984) );
  CENX2 U6199 ( .A(n4986), .B(n4984), .Z(n4894) );
  CENX1 U6200 ( .A(n4985), .B(n4894), .Z(n5000) );
  CNIVX4 U6201 ( .A(n4895), .Z(n4898) );
  COND1X4 U6202 ( .A(n4897), .B(n4898), .C(n4896), .Z(n4900) );
  CND2X2 U6203 ( .A(n4900), .B(n4899), .Z(n5002) );
  CENX2 U6204 ( .A(n5000), .B(n5002), .Z(n4907) );
  CIVX2 U6205 ( .A(n4901), .Z(n4906) );
  CNR2X2 U6206 ( .A(n4903), .B(n4902), .Z(n4905) );
  CND2X1 U6207 ( .A(n4903), .B(n4902), .Z(n4904) );
  COND1X2 U6208 ( .A(n4906), .B(n4905), .C(n4904), .Z(n5001) );
  CENX2 U6209 ( .A(n4907), .B(n2483), .Z(n5013) );
  CFA1X1 U6210 ( .A(n4911), .B(n4910), .CI(n4909), .CO(n5043), .S(n5364) );
  CENX2 U6211 ( .A(n4916), .B(n4915), .Z(n4918) );
  CENX2 U6212 ( .A(n4918), .B(n4917), .Z(n5237) );
  CENX1 U6213 ( .A(h0[17]), .B(n6118), .Z(n5111) );
  COND2X1 U6214 ( .A(n2578), .B(n5111), .C(n2490), .D(n4923), .Z(n5147) );
  CNIVX4 U6215 ( .A(n6411), .Z(n6305) );
  CND2IXL U6216 ( .B(h0[0]), .A(n6305), .Z(n4924) );
  COND2X1 U6217 ( .A(n6969), .B(n7867), .C(n4924), .D(n7171), .Z(n5173) );
  CENX1 U6218 ( .A(n7539), .B(n6305), .Z(n4925) );
  COND2X1 U6219 ( .A(n6969), .B(n4925), .C(n4955), .D(n7171), .Z(n5172) );
  CENX1 U6220 ( .A(h0[15]), .B(n6417), .Z(n5098) );
  COND2X1 U6221 ( .A(n6522), .B(n5098), .C(n6293), .D(n4926), .Z(n5146) );
  COND1X1 U6222 ( .A(n5147), .B(n5149), .C(n5146), .Z(n4928) );
  CND2X1 U6223 ( .A(n5149), .B(n5147), .Z(n4927) );
  CND2X2 U6224 ( .A(n4928), .B(n4927), .Z(n5203) );
  CFA1X1 U6225 ( .A(n4931), .B(n4930), .CI(n4929), .CO(n4915), .S(n5201) );
  CFA1X1 U6226 ( .A(n4934), .B(n4933), .CI(n4932), .CO(n4916), .S(n5202) );
  CND2X2 U6227 ( .A(n4936), .B(n4935), .Z(n5236) );
  COND1X2 U6228 ( .A(n5235), .B(n5237), .C(n5236), .Z(n4937) );
  CND2X2 U6229 ( .A(n4937), .B(n4938), .Z(n5140) );
  CENX1 U6230 ( .A(n4940), .B(n4939), .Z(n4941) );
  CENX1 U6231 ( .A(n4942), .B(n4941), .Z(n5092) );
  COR2X1 U6232 ( .A(n1556), .B(n4943), .Z(n4945) );
  CENX1 U6233 ( .A(n5888), .B(h0[13]), .Z(n5114) );
  COR2X1 U6234 ( .A(n6576), .B(n5114), .Z(n4944) );
  CND2X2 U6235 ( .A(n4945), .B(n4944), .Z(n5209) );
  CENX1 U6236 ( .A(n2583), .B(h0[19]), .Z(n5119) );
  COND2X1 U6237 ( .A(n6114), .B(n5119), .C(n3368), .D(n4958), .Z(n5211) );
  CENX1 U6238 ( .A(n6647), .B(h0[11]), .Z(n5096) );
  COND1X1 U6239 ( .A(n5209), .B(n5211), .C(n2466), .Z(n4948) );
  CENX1 U6240 ( .A(n5701), .B(n2280), .Z(n5095) );
  COND2X1 U6241 ( .A(n5911), .B(n5095), .C(n5912), .D(n4949), .Z(n5152) );
  CENX1 U6242 ( .A(n6409), .B(n5927), .Z(n5216) );
  COND2X1 U6243 ( .A(n6766), .B(n5216), .C(n6765), .D(n4950), .Z(n5151) );
  CENXL U6244 ( .A(h0[23]), .B(n2531), .Z(n5105) );
  COND2X1 U6245 ( .A(n5105), .B(n5695), .C(n4886), .D(n4952), .Z(n5145) );
  CENX1 U6246 ( .A(n5932), .B(h0[5]), .Z(n5218) );
  COND2X1 U6247 ( .A(n6974), .B(n5218), .C(n2477), .D(n4953), .Z(n5144) );
  COND2X1 U6248 ( .A(n4955), .B(n6969), .C(n7171), .D(n4954), .Z(n5143) );
  COND2X1 U6249 ( .A(n4959), .B(n4958), .C(n4957), .D(n4956), .Z(n5234) );
  CNR2IX1 U6250 ( .B(n7538), .A(n7203), .Z(n5224) );
  CENX1 U6251 ( .A(n5106), .B(h0[25]), .Z(n5107) );
  COND2X1 U6252 ( .A(n5160), .B(n5107), .C(n7537), .D(n4960), .Z(n5225) );
  CIVX2 U6253 ( .A(n7114), .Z(n4963) );
  CIVX2 U6254 ( .A(n4961), .Z(n4962) );
  CND2X2 U6255 ( .A(n4963), .B(n4962), .Z(n4964) );
  COND1X2 U6256 ( .A(n5224), .B(n5225), .C(n5223), .Z(n4967) );
  CND2X2 U6257 ( .A(n4967), .B(n4966), .Z(n5233) );
  CIVX1 U6258 ( .A(n4968), .Z(n4970) );
  CENX1 U6259 ( .A(n4970), .B(n4969), .Z(n5232) );
  CND2X2 U6260 ( .A(n4972), .B(n4971), .Z(n5139) );
  COND1X2 U6261 ( .A(n5138), .B(n5140), .C(n5139), .Z(n4974) );
  CND2X2 U6262 ( .A(n4974), .B(n4973), .Z(n5366) );
  CANR1X2 U6263 ( .A(n5364), .B(n5366), .C(n5365), .Z(n4979) );
  CNR2X2 U6264 ( .A(n5366), .B(n5364), .Z(n4978) );
  CNR2X2 U6265 ( .A(n4979), .B(n4978), .Z(n5360) );
  CNIVXL U6266 ( .A(n5360), .Z(n4980) );
  COND1X1 U6267 ( .A(n4981), .B(n5363), .C(n4980), .Z(n4983) );
  CND2X2 U6268 ( .A(n4983), .B(n4982), .Z(n5077) );
  CND2X1 U6269 ( .A(n4985), .B(n4986), .Z(n4988) );
  COND1X2 U6270 ( .A(n4986), .B(n4985), .C(n4984), .Z(n4987) );
  CND2X2 U6271 ( .A(n4988), .B(n4987), .Z(n5597) );
  CENX1 U6272 ( .A(n5932), .B(h0[12]), .Z(n5634) );
  COND2X2 U6273 ( .A(n6972), .B(n5634), .C(n6974), .D(n4989), .Z(n5623) );
  CENX1 U6274 ( .A(n7134), .B(h0[8]), .Z(n5564) );
  COND2X1 U6275 ( .A(n6969), .B(n4990), .C(n5564), .D(n7171), .Z(n5622) );
  CENX1 U6276 ( .A(h0[10]), .B(n7092), .Z(n5632) );
  COND2X1 U6277 ( .A(n2294), .B(n4992), .C(n7114), .D(n5632), .Z(n5621) );
  CEO3X2 U6278 ( .A(n5623), .B(n4993), .C(n5621), .Z(n5598) );
  CENX2 U6279 ( .A(n5597), .B(n5598), .Z(n4999) );
  CHA1X1 U6280 ( .A(n4995), .B(n4994), .CO(n5589), .S(n4986) );
  CENX1 U6281 ( .A(n6118), .B(h0[24]), .Z(n5578) );
  CENX1 U6282 ( .A(h0[26]), .B(n2583), .Z(n5580) );
  COND2X1 U6283 ( .A(n6114), .B(n4997), .C(n3368), .D(n5580), .Z(n5592) );
  COND1X2 U6284 ( .A(n5002), .B(n5001), .C(n5000), .Z(n5004) );
  CENX2 U6285 ( .A(n1571), .B(n5602), .Z(n5011) );
  COND1X2 U6286 ( .A(n5007), .B(n5006), .C(n5005), .Z(n5009) );
  CND2X2 U6287 ( .A(n5007), .B(n5006), .Z(n5008) );
  CND2X2 U6288 ( .A(n5009), .B(n5008), .Z(n5604) );
  CENX2 U6289 ( .A(n5010), .B(n5011), .Z(n5664) );
  CIVX2 U6290 ( .A(n5664), .Z(n5017) );
  COND1X2 U6291 ( .A(n5013), .B(n5014), .C(n5012), .Z(n5016) );
  CND2X2 U6292 ( .A(n5016), .B(n5015), .Z(n5666) );
  CENX2 U6293 ( .A(n5017), .B(n5666), .Z(n5076) );
  COND1X1 U6294 ( .A(n5019), .B(n5020), .C(n5018), .Z(n5022) );
  CND2X2 U6295 ( .A(n5022), .B(n5021), .Z(n5648) );
  CND2X2 U6296 ( .A(n5027), .B(n5026), .Z(n5647) );
  CND2X2 U6297 ( .A(n5032), .B(n5031), .Z(n5636) );
  CIVX1 U6298 ( .A(n5033), .Z(n5037) );
  CND2X1 U6299 ( .A(n5034), .B(n5035), .Z(n5036) );
  COND2X1 U6300 ( .A(n7228), .B(n5039), .C(n5700), .D(n2382), .Z(n5617) );
  CENX1 U6301 ( .A(n6490), .B(h0[20]), .Z(n5644) );
  COND2X2 U6302 ( .A(n6576), .B(n5040), .C(n5644), .D(n1557), .Z(n5618) );
  CENX2 U6303 ( .A(n5636), .B(n5041), .Z(n5645) );
  COND1X2 U6304 ( .A(n5045), .B(n5044), .C(n5043), .Z(n5654) );
  CND2X2 U6305 ( .A(n5045), .B(n5044), .Z(n5652) );
  CND2X2 U6306 ( .A(n5654), .B(n5652), .Z(n5658) );
  CAOR1X1 U6307 ( .A(n7537), .B(n5160), .C(n5046), .Z(n5586) );
  CENX1 U6308 ( .A(n7202), .B(n7674), .Z(n5570) );
  COND2X1 U6309 ( .A(n7205), .B(n5047), .C(n7203), .D(n5570), .Z(n5584) );
  CENX1 U6310 ( .A(n5586), .B(n5584), .Z(n5049) );
  CENX1 U6311 ( .A(h0[16]), .B(n6409), .Z(n5572) );
  COND2X2 U6312 ( .A(n6765), .B(n5572), .C(n6701), .D(n5048), .Z(n5585) );
  CENX2 U6313 ( .A(n5049), .B(n5585), .Z(n5607) );
  CENX1 U6314 ( .A(n6417), .B(h0[22]), .Z(n5642) );
  COND2X1 U6315 ( .A(n6211), .B(n5050), .C(n5984), .D(n5642), .Z(n5627) );
  COND2X1 U6316 ( .A(n6703), .B(n5051), .C(n2515), .D(n5565), .Z(n5626) );
  CENX1 U6317 ( .A(n5701), .B(h0[28]), .Z(n5643) );
  COND2X1 U6318 ( .A(n5911), .B(n5052), .C(n5912), .D(n5643), .Z(n5628) );
  COND2X1 U6319 ( .A(n5695), .B(n5054), .C(n5696), .D(n5567), .Z(n5583) );
  CENX1 U6320 ( .A(n6103), .B(n2512), .Z(n5571) );
  COND2X1 U6321 ( .A(n5055), .B(n2282), .C(n2433), .D(n5571), .Z(n5582) );
  CENX1 U6322 ( .A(n6828), .B(h0[14]), .Z(n5633) );
  COND2X1 U6323 ( .A(n6870), .B(n5056), .C(n6829), .D(n5633), .Z(n5581) );
  CENX2 U6324 ( .A(n5608), .B(n5609), .Z(n5057) );
  CENX2 U6325 ( .A(n5607), .B(n5057), .Z(n5561) );
  CND2IX1 U6326 ( .B(n5058), .A(n5060), .Z(n5063) );
  CND2X2 U6327 ( .A(n5063), .B(n5062), .Z(n5613) );
  CFA1X1 U6328 ( .A(n5064), .B(n5065), .CI(n5066), .CO(n5612), .S(n5018) );
  CFA1X1 U6329 ( .A(n5069), .B(n5067), .CI(n5068), .CO(n5614), .S(n5072) );
  CNIVX2 U6330 ( .A(n5614), .Z(n5070) );
  CENX2 U6331 ( .A(n5071), .B(n5070), .Z(n5560) );
  CEO3X1 U6332 ( .A(n2292), .B(n5655), .C(n5658), .Z(n5667) );
  CIVX2 U6333 ( .A(n5667), .Z(n5075) );
  CND2X2 U6334 ( .A(n5077), .B(n5078), .Z(n7309) );
  CIVXL U6335 ( .A(n7310), .Z(n5079) );
  CENX2 U6336 ( .A(n5081), .B(n5080), .Z(n5082) );
  CEO3X2 U6337 ( .A(n5086), .B(n5085), .C(n5084), .Z(n5374) );
  CENX2 U6338 ( .A(n5094), .B(n5093), .Z(n5246) );
  CENX1 U6339 ( .A(n5701), .B(h0[20]), .Z(n5181) );
  COND2X1 U6340 ( .A(n6703), .B(n5190), .C(n2514), .D(n5096), .Z(n5254) );
  CENXL U6341 ( .A(n6828), .B(n2443), .Z(n5166) );
  COND2X1 U6342 ( .A(n5166), .B(n6870), .C(n6829), .D(n5097), .Z(n5253) );
  CIVX2 U6343 ( .A(n5098), .Z(n5100) );
  CND2X2 U6344 ( .A(n5100), .B(n5099), .Z(n5103) );
  CIVX2 U6345 ( .A(n5294), .Z(n5101) );
  CND2X2 U6346 ( .A(n5103), .B(n5102), .Z(n5108) );
  CIVX2 U6347 ( .A(n5108), .Z(n5260) );
  CENX1 U6348 ( .A(h0[22]), .B(n2531), .Z(n5170) );
  COND2X1 U6349 ( .A(n5695), .B(n5170), .C(n4886), .D(n5105), .Z(n5261) );
  CIVX1 U6350 ( .A(n5261), .Z(n5110) );
  CENX1 U6351 ( .A(n5106), .B(h0[24]), .Z(n5158) );
  COND2X1 U6352 ( .A(n5160), .B(n5158), .C(n7537), .D(n5107), .Z(n5262) );
  COND1X2 U6353 ( .A(n5108), .B(n5261), .C(n5262), .Z(n5109) );
  COND1X4 U6354 ( .A(n5260), .B(n5110), .C(n5109), .Z(n5178) );
  CENX1 U6355 ( .A(h0[16]), .B(n6191), .Z(n5192) );
  CENX1 U6356 ( .A(n5888), .B(h0[12]), .Z(n5194) );
  CIVX2 U6357 ( .A(n5194), .Z(n5113) );
  CND2X2 U6358 ( .A(n5113), .B(n5112), .Z(n5118) );
  CIVX2 U6359 ( .A(n5114), .Z(n5116) );
  CIVX2 U6360 ( .A(n1556), .Z(n5115) );
  CND2X2 U6361 ( .A(n5116), .B(n5115), .Z(n5117) );
  CND2X2 U6362 ( .A(n5118), .B(n5117), .Z(n5187) );
  CENX1 U6363 ( .A(h0[18]), .B(n5923), .Z(n5184) );
  COND2X1 U6364 ( .A(n6114), .B(n5184), .C(n3368), .D(n5119), .Z(n5186) );
  COND1X1 U6365 ( .A(n2365), .B(n5187), .C(n5186), .Z(n5121) );
  CND2X2 U6366 ( .A(n5121), .B(n5120), .Z(n5177) );
  CND2X2 U6367 ( .A(n5123), .B(n5122), .Z(n5280) );
  CENX2 U6368 ( .A(n5125), .B(n5124), .Z(n5126) );
  CENX2 U6369 ( .A(n5127), .B(n5126), .Z(n5277) );
  CFA1X1 U6370 ( .A(n5130), .B(n5129), .CI(n5128), .CO(n4920), .S(n5278) );
  CND2X2 U6371 ( .A(n5133), .B(n5132), .Z(n5247) );
  COND1X2 U6372 ( .A(n5248), .B(n5246), .C(n5247), .Z(n5135) );
  CND2X1 U6373 ( .A(n5246), .B(n5248), .Z(n5134) );
  CND2X2 U6374 ( .A(n5135), .B(n5134), .Z(n5375) );
  CNIVX4 U6375 ( .A(n5375), .Z(n5136) );
  CENX2 U6376 ( .A(n5137), .B(n5136), .Z(n5389) );
  CENX2 U6377 ( .A(n5139), .B(n5138), .Z(n5142) );
  CENX2 U6378 ( .A(n5142), .B(n5141), .Z(n5388) );
  CFA1X1 U6379 ( .A(n5143), .B(n5144), .CI(n5145), .CO(n5229), .S(n5250) );
  CENX1 U6380 ( .A(n5147), .B(n5146), .Z(n5148) );
  CENX2 U6381 ( .A(n5149), .B(n5148), .Z(n5252) );
  CFA1X1 U6382 ( .A(n5150), .B(n5151), .CI(n5152), .CO(n5230), .S(n5249) );
  CND2X2 U6383 ( .A(n5154), .B(n5153), .Z(n5293) );
  CND2IX1 U6384 ( .B(n5219), .A(n5155), .Z(n5156) );
  COND1X1 U6385 ( .A(n5157), .B(n6974), .C(n5156), .Z(n5161) );
  CND2IX2 U6386 ( .B(n5306), .A(n5303), .Z(n5165) );
  CND2IX1 U6387 ( .B(n5162), .A(n5161), .Z(n5163) );
  CND2IX2 U6388 ( .B(n5305), .A(n5163), .Z(n5164) );
  CIVX2 U6389 ( .A(n5321), .Z(n5174) );
  COND2X1 U6390 ( .A(n6870), .B(n5167), .C(n6829), .D(n5166), .Z(n5341) );
  COND2X1 U6391 ( .A(n2294), .B(n5169), .C(n2374), .D(n5212), .Z(n5340) );
  CHA1X1 U6392 ( .A(n5173), .B(n5172), .CO(n5149), .S(n5322) );
  COND1X2 U6393 ( .A(n5174), .B(n5320), .C(n5322), .Z(n5176) );
  CND2X2 U6394 ( .A(n5176), .B(n5175), .Z(n5327) );
  COND2X1 U6395 ( .A(n5182), .B(n5911), .C(n5912), .D(n5181), .Z(n5338) );
  CENX1 U6396 ( .A(n6409), .B(h0[8]), .Z(n5217) );
  COND2X1 U6397 ( .A(n6701), .B(n5183), .C(n6765), .D(n5217), .Z(n5337) );
  COND2X1 U6398 ( .A(n6114), .B(n5185), .C(n3368), .D(n5184), .Z(n5336) );
  CENX2 U6399 ( .A(n5186), .B(n5189), .Z(n5331) );
  COND2X1 U6400 ( .A(n5191), .B(n6703), .C(n6702), .D(n5190), .Z(n5344) );
  COND2X1 U6401 ( .A(n2569), .B(n5193), .C(n2487), .D(n5192), .Z(n5343) );
  COND2X1 U6402 ( .A(n2449), .B(n5195), .C(n1557), .D(n5194), .Z(n5342) );
  CND2X1 U6403 ( .A(n5331), .B(n5328), .Z(n5196) );
  CND2X2 U6404 ( .A(n5197), .B(n5196), .Z(n5326) );
  COND1X2 U6405 ( .A(n5198), .B(n5325), .C(n5326), .Z(n5200) );
  CND2X2 U6406 ( .A(n5200), .B(n5199), .Z(n5291) );
  COND1X2 U6407 ( .A(n5293), .B(n5291), .C(n5292), .Z(n5208) );
  CND2X2 U6408 ( .A(n5291), .B(n5206), .Z(n5207) );
  CND2X2 U6409 ( .A(n5208), .B(n5207), .Z(n5244) );
  CIVX1 U6410 ( .A(n5212), .Z(n5213) );
  CND2IXL U6411 ( .B(n2295), .A(n5213), .Z(n5215) );
  CND2X1 U6412 ( .A(n5215), .B(n5214), .Z(n5259) );
  COND2X1 U6413 ( .A(n6701), .B(n5217), .C(n6765), .D(n5216), .Z(n5256) );
  COND2X1 U6414 ( .A(n6974), .B(n5219), .C(n6972), .D(n5218), .Z(n5257) );
  CNIVX1 U6415 ( .A(n5225), .Z(n5226) );
  COND1X1 U6416 ( .A(n5267), .B(n5268), .C(n5270), .Z(n5228) );
  CND2X2 U6417 ( .A(n5228), .B(n5227), .Z(n5276) );
  CFA1X1 U6418 ( .A(n5231), .B(n5230), .CI(n5229), .CO(n5094), .S(n5275) );
  CFA1X1 U6419 ( .A(n5234), .B(n5233), .CI(n5232), .CO(n5091), .S(n5274) );
  CENX2 U6420 ( .A(n5235), .B(n5236), .Z(n5239) );
  CENX2 U6421 ( .A(n5238), .B(n5239), .Z(n5245) );
  CND2X2 U6422 ( .A(n5241), .B(n5240), .Z(n5387) );
  CENX2 U6423 ( .A(n5388), .B(n5387), .Z(n5242) );
  CEO3X2 U6424 ( .A(n5247), .B(n5248), .C(n2415), .Z(n5287) );
  CENX2 U6425 ( .A(n5252), .B(n5251), .Z(n5401) );
  CFA1X1 U6426 ( .A(n5254), .B(n5255), .CI(n5253), .CO(n5180), .S(n5332) );
  CENX2 U6427 ( .A(n5259), .B(n5258), .Z(n5335) );
  CIVX2 U6428 ( .A(n5260), .Z(n5264) );
  CENX1 U6429 ( .A(n5262), .B(n5261), .Z(n5263) );
  CENX2 U6430 ( .A(n5264), .B(n5263), .Z(n5333) );
  CND2X2 U6431 ( .A(n5335), .B(n5332), .Z(n5265) );
  CND2X2 U6432 ( .A(n5266), .B(n5265), .Z(n5402) );
  CND2X1 U6433 ( .A(n5401), .B(n5402), .Z(n5273) );
  CND2X1 U6434 ( .A(n5403), .B(n5401), .Z(n5272) );
  CND2X1 U6435 ( .A(n2375), .B(n5402), .Z(n5271) );
  CND3X2 U6436 ( .A(n5273), .B(n5272), .C(n5271), .Z(n5354) );
  CFA1X1 U6437 ( .A(n5276), .B(n5275), .CI(n5274), .CO(n5243), .S(n5353) );
  CND2X1 U6438 ( .A(n5354), .B(n5353), .Z(n5283) );
  CENX2 U6439 ( .A(n5278), .B(n5277), .Z(n5279) );
  CENX2 U6440 ( .A(n5280), .B(n5279), .Z(n5355) );
  CND2X1 U6441 ( .A(n5353), .B(n5355), .Z(n5282) );
  CND2X1 U6442 ( .A(n5354), .B(n5355), .Z(n5281) );
  CND3X2 U6443 ( .A(n5283), .B(n5282), .C(n5281), .Z(n5288) );
  CIVX2 U6444 ( .A(n5287), .Z(n5284) );
  CND2IX1 U6445 ( .B(n5284), .A(n5290), .Z(n5285) );
  CEO3X2 U6446 ( .A(n5293), .B(n5292), .C(n5291), .Z(n5461) );
  COND2X1 U6447 ( .A(n1262), .B(n5295), .C(n6523), .D(n5294), .Z(n5410) );
  CFA1X1 U6448 ( .A(n5298), .B(n5297), .CI(n5296), .CO(n5413), .S(n5447) );
  CAN2X2 U6449 ( .A(n5300), .B(n5299), .Z(n5411) );
  COND1X1 U6450 ( .A(n5410), .B(n5413), .C(n5411), .Z(n5302) );
  CND2X1 U6451 ( .A(n5410), .B(n5413), .Z(n5301) );
  CIVX2 U6452 ( .A(n5303), .Z(n5304) );
  CEO3X2 U6453 ( .A(n5306), .B(n5305), .C(n5304), .Z(n5421) );
  COND1X1 U6454 ( .A(n5308), .B(n5309), .C(n5307), .Z(n5311) );
  CND2X1 U6455 ( .A(n5309), .B(n5308), .Z(n5310) );
  CND2X2 U6456 ( .A(n5310), .B(n5311), .Z(n5419) );
  CND2X1 U6457 ( .A(n5421), .B(n5419), .Z(n5319) );
  COND1X1 U6458 ( .A(n5314), .B(n5313), .C(n5312), .Z(n5316) );
  CND2X1 U6459 ( .A(n5316), .B(n5315), .Z(n5420) );
  CND2X1 U6460 ( .A(n5421), .B(n5420), .Z(n5318) );
  CND2XL U6461 ( .A(n5419), .B(n5420), .Z(n5317) );
  CND3X2 U6462 ( .A(n5319), .B(n5318), .C(n5317), .Z(n5433) );
  CIVX2 U6463 ( .A(n5320), .Z(n5324) );
  CENX2 U6464 ( .A(n5322), .B(n2493), .Z(n5323) );
  CENX2 U6465 ( .A(n5324), .B(n5323), .Z(n5432) );
  CEO3X2 U6466 ( .A(n5327), .B(n5326), .C(n5325), .Z(n5397) );
  CENX2 U6467 ( .A(n2363), .B(n5330), .Z(n5438) );
  CENX2 U6468 ( .A(n5333), .B(n5332), .Z(n5334) );
  CENX2 U6469 ( .A(n5335), .B(n5334), .Z(n5440) );
  CFA1X1 U6470 ( .A(n5336), .B(n5337), .CI(n5338), .CO(n5328), .S(n5426) );
  COND1X2 U6471 ( .A(n5426), .B(n5345), .C(n5423), .Z(n5347) );
  CND2X2 U6472 ( .A(n5347), .B(n5346), .Z(n5439) );
  COND1X2 U6473 ( .A(n1258), .B(n5440), .C(n5439), .Z(n5349) );
  CND2X2 U6474 ( .A(n5440), .B(n1258), .Z(n5348) );
  CND2X2 U6475 ( .A(n5349), .B(n5348), .Z(n5400) );
  CND2X2 U6476 ( .A(n5350), .B(n5400), .Z(n5352) );
  CND2X1 U6477 ( .A(n5397), .B(n5398), .Z(n5351) );
  CND2X2 U6478 ( .A(n5352), .B(n5351), .Z(n5460) );
  CNIVXL U6479 ( .A(n5460), .Z(n5356) );
  CND2X1 U6480 ( .A(n5461), .B(n5356), .Z(n5359) );
  CEO3X2 U6481 ( .A(n5355), .B(n5354), .C(n5353), .Z(n5462) );
  CND2X1 U6482 ( .A(n2455), .B(n5461), .Z(n5358) );
  CND3X2 U6483 ( .A(n5359), .B(n5358), .C(n5357), .Z(n5517) );
  CNR2X2 U6484 ( .A(n5555), .B(n2335), .Z(n5547) );
  CENX2 U6485 ( .A(n5361), .B(n5360), .Z(n5362) );
  CENX2 U6486 ( .A(n5362), .B(n5363), .Z(n5541) );
  CIVX2 U6487 ( .A(n5366), .Z(n5367) );
  CIVX2 U6488 ( .A(n5369), .Z(n5372) );
  CND2X2 U6489 ( .A(n5377), .B(n5376), .Z(n5384) );
  CNIVX4 U6490 ( .A(n5384), .Z(n5378) );
  CND2X2 U6491 ( .A(n5379), .B(n5378), .Z(n5380) );
  COND1X2 U6492 ( .A(n5386), .B(n5381), .C(n5380), .Z(n5540) );
  CNR2X2 U6493 ( .A(n5541), .B(n5540), .Z(n5523) );
  CIVDX2 U6494 ( .A(n5382), .Z0(n5383), .Z1(n5379) );
  CENX2 U6495 ( .A(n5384), .B(n5383), .Z(n5385) );
  CENX2 U6496 ( .A(n5385), .B(n5386), .Z(n5522) );
  CND2X2 U6497 ( .A(n5391), .B(n5390), .Z(n5521) );
  CNR2X2 U6498 ( .A(n5522), .B(n5521), .Z(n5548) );
  CNR2X2 U6499 ( .A(n5523), .B(n5548), .Z(n5525) );
  CND2X2 U6500 ( .A(n5525), .B(n5547), .Z(n5528) );
  CND2X2 U6501 ( .A(n5396), .B(n5392), .Z(n5533) );
  CIVX2 U6502 ( .A(n5393), .Z(n5394) );
  CANR1X2 U6503 ( .A(n5396), .B(n5395), .C(n5394), .Z(n5531) );
  COND1X2 U6504 ( .A(n5533), .B(n5532), .C(n5531), .Z(n5516) );
  CENX2 U6505 ( .A(n5398), .B(n5397), .Z(n5399) );
  CENX2 U6506 ( .A(n5400), .B(n5399), .Z(n5506) );
  CIVX2 U6507 ( .A(n5401), .Z(n5406) );
  CIVX2 U6508 ( .A(n5402), .Z(n5404) );
  CENX2 U6509 ( .A(n5404), .B(n2375), .Z(n5405) );
  CENX2 U6510 ( .A(n5406), .B(n5405), .Z(n5464) );
  CFA1X1 U6511 ( .A(n5409), .B(n5408), .CI(n5407), .CO(n5455), .S(n5446) );
  CENX2 U6512 ( .A(n5410), .B(n5411), .Z(n5412) );
  COND1X2 U6513 ( .A(n5416), .B(n5415), .C(n5414), .Z(n5418) );
  CND2X2 U6514 ( .A(n5418), .B(n5417), .Z(n5453) );
  CEOX2 U6515 ( .A(n5420), .B(n5419), .Z(n5422) );
  CEOX2 U6516 ( .A(n5422), .B(n5421), .Z(n5470) );
  CENX2 U6517 ( .A(n5424), .B(n5423), .Z(n5425) );
  CENX2 U6518 ( .A(n5425), .B(n5426), .Z(n5469) );
  CFA1X1 U6519 ( .A(n5429), .B(n5428), .CI(n5427), .CO(n5471), .S(n5476) );
  COND1X2 U6520 ( .A(n5470), .B(n5469), .C(n5471), .Z(n5431) );
  CND2X2 U6521 ( .A(n5431), .B(n5430), .Z(n5443) );
  CENX2 U6522 ( .A(n5464), .B(n5465), .Z(n5437) );
  CENX2 U6523 ( .A(n5506), .B(n5437), .Z(n7010) );
  CEO3X2 U6524 ( .A(n5444), .B(n5443), .C(n5442), .Z(n5490) );
  CFA1X1 U6525 ( .A(n5447), .B(n5446), .CI(n5445), .CO(n5480), .S(n5475) );
  COND1X2 U6526 ( .A(n5450), .B(n5449), .C(n5448), .Z(n5452) );
  CND2X2 U6527 ( .A(n5452), .B(n5451), .Z(n5479) );
  CFA1X1 U6528 ( .A(n5455), .B(n5454), .CI(n5453), .CO(n5444), .S(n5482) );
  CND2X2 U6529 ( .A(n5459), .B(n5458), .Z(n7009) );
  CNR2X2 U6530 ( .A(n7010), .B(n7009), .Z(n5468) );
  CENX2 U6531 ( .A(n5461), .B(n5460), .Z(n5463) );
  CENX2 U6532 ( .A(n5463), .B(n5462), .Z(n5511) );
  CNIVX4 U6533 ( .A(n5465), .Z(n5505) );
  CND2X2 U6534 ( .A(n5466), .B(n5509), .Z(n5467) );
  CIVX2 U6535 ( .A(n5503), .Z(n5530) );
  CENX1 U6536 ( .A(n5471), .B(n5470), .Z(n5472) );
  CND2X2 U6537 ( .A(n5478), .B(n5477), .Z(n5493) );
  CENX2 U6538 ( .A(n2437), .B(n5481), .Z(n5495) );
  CNR2X1 U6539 ( .A(n5498), .B(n5499), .Z(n7013) );
  CIVX2 U6540 ( .A(n7013), .Z(n6381) );
  CENX2 U6541 ( .A(n5489), .B(n5488), .Z(n5491) );
  CENX2 U6542 ( .A(n5491), .B(n5490), .Z(n5501) );
  COND1X2 U6543 ( .A(n5494), .B(n5495), .C(n5493), .Z(n5497) );
  CND2X1 U6544 ( .A(n5495), .B(n5494), .Z(n5496) );
  CND2X2 U6545 ( .A(n5497), .B(n5496), .Z(n5500) );
  CNR2X2 U6546 ( .A(n5501), .B(n5500), .Z(n5502) );
  CIVX2 U6547 ( .A(n5502), .Z(n7015) );
  CND2X2 U6548 ( .A(n6381), .B(n7015), .Z(n7487) );
  CNR2X2 U6549 ( .A(n5530), .B(n7487), .Z(n5515) );
  CND2X2 U6550 ( .A(n5499), .B(n5498), .Z(n7012) );
  CND2X2 U6551 ( .A(n5501), .B(n5500), .Z(n7014) );
  COND1X2 U6552 ( .A(n7012), .B(n5502), .C(n7014), .Z(n7489) );
  CND2X2 U6553 ( .A(n7489), .B(n5503), .Z(n5514) );
  CIVX2 U6554 ( .A(n5504), .Z(n7497) );
  CND2X2 U6555 ( .A(n5511), .B(n5510), .Z(n7496) );
  CIVX2 U6556 ( .A(n7496), .Z(n5512) );
  CND2X2 U6557 ( .A(n5513), .B(n5514), .Z(n5534) );
  CND2X2 U6558 ( .A(n5518), .B(n5517), .Z(n7510) );
  CND2X1 U6559 ( .A(n5520), .B(n5519), .Z(n5554) );
  COND1X2 U6560 ( .A(n7510), .B(n5553), .C(n5554), .Z(n5546) );
  CND2X1 U6561 ( .A(n5541), .B(n5540), .Z(n5542) );
  CANR1X2 U6562 ( .A(n5546), .B(n5525), .C(n5524), .Z(n5526) );
  CIVX2 U6563 ( .A(n1257), .Z(n7475) );
  CIVXL U6564 ( .A(n2431), .Z(n5529) );
  CNR2XL U6565 ( .A(n5529), .B(n5548), .Z(n5539) );
  CNR2XL U6566 ( .A(n5530), .B(n7487), .Z(n5535) );
  COND1XL U6567 ( .A(n5533), .B(n2284), .C(n5531), .Z(n6382) );
  CANR1XL U6568 ( .A(n5535), .B(n6382), .C(n5534), .Z(n5536) );
  CIVXL U6569 ( .A(n5536), .Z(n7513) );
  CIVXL U6570 ( .A(n5546), .Z(n5537) );
  COND1XL U6571 ( .A(n5548), .B(n5537), .C(n5549), .Z(n5538) );
  CANR1XL U6572 ( .A(n5539), .B(n7513), .C(n5538), .Z(n5545) );
  COR2XL U6573 ( .A(n5540), .B(n5541), .Z(n5543) );
  CAN2XL U6574 ( .A(n5542), .B(n5543), .Z(n5544) );
  CENXL U6575 ( .A(n5544), .B(n5545), .Z(N46) );
  CANR1XL U6576 ( .A(n2431), .B(n7513), .C(n5546), .Z(n5552) );
  CIVXL U6577 ( .A(n5548), .Z(n5550) );
  CAN2XL U6578 ( .A(n5550), .B(n5549), .Z(n5551) );
  CENXL U6579 ( .A(n5551), .B(n5552), .Z(N45) );
  CNR2IXL U6580 ( .B(n5554), .A(n2335), .Z(n5558) );
  CIVXL U6581 ( .A(n5555), .Z(n7511) );
  CIVXL U6582 ( .A(n7510), .Z(n5556) );
  CANR1XL U6583 ( .A(n7511), .B(n7513), .C(n5556), .Z(n5557) );
  CENXL U6584 ( .A(n5558), .B(n5557), .Z(N44) );
  CND2X2 U6585 ( .A(n5563), .B(n5562), .Z(n5771) );
  CENX1 U6586 ( .A(n7134), .B(n5927), .Z(n5763) );
  COND2X1 U6587 ( .A(n6969), .B(n5564), .C(n7171), .D(n5763), .Z(n5742) );
  CNIVXL U6588 ( .A(n5742), .Z(n5569) );
  COND2X1 U6589 ( .A(n5565), .B(n6703), .C(n6702), .D(n5709), .Z(n5743) );
  CENXL U6590 ( .A(h0[31]), .B(n5104), .Z(n5697) );
  COND2X1 U6591 ( .A(n5695), .B(n5567), .C(n5696), .D(n5697), .Z(n5741) );
  CENX1 U6592 ( .A(h0[7]), .B(n7202), .Z(n5764) );
  COND2X2 U6593 ( .A(n7217), .B(n5570), .C(n7203), .D(n5764), .Z(n5729) );
  CENX1 U6594 ( .A(n6103), .B(h0[5]), .Z(n5756) );
  COND2X2 U6595 ( .A(n2433), .B(n5756), .C(n2282), .D(n5571), .Z(n5728) );
  CNR2X4 U6596 ( .A(n6701), .B(n5572), .Z(n5573) );
  CENX1 U6597 ( .A(h0[17]), .B(n6409), .Z(n5704) );
  CNR2X2 U6598 ( .A(n6765), .B(n5704), .Z(n5574) );
  CENX2 U6599 ( .A(n5728), .B(n2348), .Z(n5577) );
  CENX2 U6600 ( .A(n5577), .B(n5729), .Z(n5684) );
  CENX1 U6601 ( .A(n6118), .B(h0[25]), .Z(n5765) );
  COND2X1 U6602 ( .A(n7228), .B(n5700), .C(n5755), .D(n7301), .Z(n5579) );
  CIVX1 U6603 ( .A(n5579), .Z(n5721) );
  CND2X2 U6604 ( .A(n5588), .B(n5587), .Z(n5735) );
  CND2X1 U6605 ( .A(n5592), .B(n5591), .Z(n5593) );
  CNIVX2 U6606 ( .A(n5736), .Z(n5595) );
  CIVX2 U6607 ( .A(n5596), .Z(n5600) );
  COND1X2 U6608 ( .A(n5603), .B(n5604), .C(n5602), .Z(n5606) );
  CND2X1 U6609 ( .A(n5604), .B(n1571), .Z(n5605) );
  CND2X2 U6610 ( .A(n5606), .B(n5605), .Z(n5770) );
  CEO3X2 U6611 ( .A(n5771), .B(n5769), .C(n5770), .Z(n5776) );
  CIVX2 U6612 ( .A(n5776), .Z(n5663) );
  COND1X1 U6613 ( .A(n5608), .B(n5609), .C(n5607), .Z(n5611) );
  CND2X1 U6614 ( .A(n5609), .B(n5608), .Z(n5610) );
  CND2X2 U6615 ( .A(n5611), .B(n5610), .Z(n5752) );
  CND2X1 U6616 ( .A(n5614), .B(n5613), .Z(n5615) );
  CND2X2 U6617 ( .A(n5616), .B(n5615), .Z(n5748) );
  CIVX1 U6618 ( .A(n5617), .Z(n5620) );
  CIVX2 U6619 ( .A(n5618), .Z(n5619) );
  CND2X2 U6620 ( .A(n5620), .B(n5619), .Z(n5760) );
  CND2X1 U6621 ( .A(n5622), .B(n5623), .Z(n5625) );
  COND1X1 U6622 ( .A(n5623), .B(n5622), .C(n5621), .Z(n5624) );
  CND2X2 U6623 ( .A(n5625), .B(n5624), .Z(n5759) );
  COND1X1 U6624 ( .A(n5628), .B(n5627), .C(n5626), .Z(n5630) );
  CND2X1 U6625 ( .A(n5628), .B(n5627), .Z(n5629) );
  CND2X1 U6626 ( .A(n5630), .B(n5629), .Z(n5758) );
  CEO3X2 U6627 ( .A(n5760), .B(n5758), .C(n5759), .Z(n5749) );
  CENX2 U6628 ( .A(n5748), .B(n5749), .Z(n5631) );
  COND2X1 U6629 ( .A(n2294), .B(n5632), .C(n7114), .D(n5690), .Z(n5725) );
  CENX1 U6630 ( .A(n6828), .B(h0[15]), .Z(n5691) );
  COND2X1 U6631 ( .A(n6870), .B(n5633), .C(n6829), .D(n5691), .Z(n5724) );
  CENX1 U6632 ( .A(h0[13]), .B(n5932), .Z(n5692) );
  COND2X1 U6633 ( .A(n6974), .B(n5634), .C(n5692), .D(n6972), .Z(n5723) );
  CENX1 U6634 ( .A(n5725), .B(n5635), .Z(n5689) );
  CIVX2 U6635 ( .A(n5636), .Z(n5641) );
  CNR2X1 U6636 ( .A(n5637), .B(n5638), .Z(n5640) );
  CND2XL U6637 ( .A(n5638), .B(n5637), .Z(n5639) );
  COND1X1 U6638 ( .A(n5641), .B(n5640), .C(n5639), .Z(n5688) );
  COND2X1 U6639 ( .A(n6211), .B(n5642), .C(n5984), .D(n2283), .Z(n5746) );
  CENX1 U6640 ( .A(n5701), .B(h0[29]), .Z(n5702) );
  COND2X1 U6641 ( .A(n5911), .B(n5643), .C(n5912), .D(n5702), .Z(n5745) );
  CENX1 U6642 ( .A(n6490), .B(n2280), .Z(n5740) );
  COND2X1 U6643 ( .A(n6576), .B(n5644), .C(n6525), .D(n5740), .Z(n5744) );
  CNIVX1 U6644 ( .A(n5645), .Z(n5646) );
  CND2X2 U6645 ( .A(n5648), .B(n5647), .Z(n5649) );
  CND2X2 U6646 ( .A(n5650), .B(n5649), .Z(n5673) );
  CIVXL U6647 ( .A(n2291), .Z(n5653) );
  CND3X1 U6648 ( .A(n5654), .B(n5653), .C(n5652), .Z(n5656) );
  CND2X2 U6649 ( .A(n5656), .B(n5655), .Z(n5660) );
  CND2X2 U6650 ( .A(n5658), .B(n5657), .Z(n5659) );
  CENX2 U6651 ( .A(n5661), .B(n5777), .Z(n5662) );
  CENX2 U6652 ( .A(n5663), .B(n5662), .Z(n6265) );
  CNIVX4 U6653 ( .A(n5664), .Z(n5665) );
  CND2X1 U6654 ( .A(n1577), .B(n5665), .Z(n5670) );
  CNR2X2 U6655 ( .A(n5665), .B(n5666), .Z(n5668) );
  CND2IX1 U6656 ( .B(n5668), .A(n2596), .Z(n5669) );
  CND2X2 U6657 ( .A(n5670), .B(n5669), .Z(n6266) );
  CNR2X2 U6658 ( .A(n6265), .B(n6266), .Z(n7306) );
  CNR2X1 U6659 ( .A(n7306), .B(n7310), .Z(n7469) );
  CND2X2 U6660 ( .A(n5673), .B(n2358), .Z(n5674) );
  CND2X2 U6661 ( .A(n5675), .B(n5674), .Z(n5828) );
  COND1X1 U6662 ( .A(n5677), .B(n5679), .C(n5676), .Z(n5681) );
  CNIVX1 U6663 ( .A(n5677), .Z(n5678) );
  CND2X2 U6664 ( .A(n5679), .B(n5678), .Z(n5680) );
  CND2X2 U6665 ( .A(n5681), .B(n5680), .Z(n5830) );
  COND1X1 U6666 ( .A(n5683), .B(n5684), .C(n5682), .Z(n5686) );
  CND2X1 U6667 ( .A(n5683), .B(n5684), .Z(n5685) );
  CFA1X1 U6668 ( .A(n5689), .B(n5688), .CI(n5687), .CO(n5834), .S(n5672) );
  CENX1 U6669 ( .A(h0[12]), .B(n2659), .Z(n5797) );
  COND2X2 U6670 ( .A(n7114), .B(n5797), .C(n5690), .D(n2293), .Z(n5875) );
  COND2X1 U6671 ( .A(n6831), .B(n5691), .C(n6829), .D(n5866), .Z(n5874) );
  CENX1 U6672 ( .A(h0[14]), .B(n5932), .Z(n5864) );
  COR2XL U6673 ( .A(n6972), .B(n5864), .Z(n5693) );
  CND2X1 U6674 ( .A(n5694), .B(n5693), .Z(n5873) );
  CEO3X2 U6675 ( .A(n5875), .B(n5874), .C(n5873), .Z(n5804) );
  CIVX2 U6676 ( .A(n5804), .Z(n5718) );
  CND2X1 U6677 ( .A(n5696), .B(n5695), .Z(n5699) );
  CIVXL U6678 ( .A(n5697), .Z(n5698) );
  CND2X2 U6679 ( .A(n5699), .B(n5698), .Z(n5810) );
  COND2X1 U6680 ( .A(n7228), .B(n5700), .C(n5755), .D(n7301), .Z(n5812) );
  CENX1 U6681 ( .A(n5701), .B(h0[30]), .Z(n5794) );
  CENX2 U6682 ( .A(n5810), .B(n5703), .Z(n5802) );
  CENX1 U6683 ( .A(h0[18]), .B(n6409), .Z(n5791) );
  COR2X1 U6684 ( .A(n6765), .B(n5791), .Z(n5707) );
  CIVX2 U6685 ( .A(n5705), .Z(n5706) );
  CND2X2 U6686 ( .A(n5707), .B(n5706), .Z(n5850) );
  CIVX2 U6687 ( .A(n5850), .Z(n5801) );
  COND2X2 U6688 ( .A(n6523), .B(n5867), .C(n5708), .D(n6522), .Z(n5848) );
  CIVX2 U6689 ( .A(n5709), .Z(n5710) );
  CENX1 U6690 ( .A(n2660), .B(h0[20]), .Z(n5870) );
  CIVX2 U6691 ( .A(n5870), .Z(n5713) );
  CND2X2 U6692 ( .A(n5713), .B(n5712), .Z(n5714) );
  CND2X2 U6693 ( .A(n5715), .B(n5714), .Z(n5849) );
  CENX2 U6694 ( .A(n5848), .B(n5849), .Z(n5800) );
  CENX2 U6695 ( .A(n5802), .B(n5716), .Z(n5717) );
  CENX2 U6696 ( .A(n5718), .B(n5717), .Z(n5833) );
  CEO3X2 U6697 ( .A(n5835), .B(n5834), .C(n5833), .Z(n5831) );
  CENX2 U6698 ( .A(n5830), .B(n5831), .Z(n5719) );
  CENX2 U6699 ( .A(n5828), .B(n5719), .Z(n5885) );
  COND1X1 U6700 ( .A(n5724), .B(n5725), .C(n1267), .Z(n5727) );
  CND2X1 U6701 ( .A(n5725), .B(n5724), .Z(n5726) );
  CND2X2 U6702 ( .A(n5727), .B(n5726), .Z(n5805) );
  COND1X2 U6703 ( .A(n5729), .B(n2349), .C(n5728), .Z(n5732) );
  CND2X1 U6704 ( .A(n5730), .B(n5729), .Z(n5731) );
  CND2X2 U6705 ( .A(n5732), .B(n5731), .Z(n5807) );
  CENX2 U6706 ( .A(n5805), .B(n5807), .Z(n5733) );
  CENX2 U6707 ( .A(n5734), .B(n5733), .Z(n5823) );
  COND1X1 U6708 ( .A(n5736), .B(n5737), .C(n5735), .Z(n5739) );
  CND2X2 U6709 ( .A(n5739), .B(n5738), .Z(n5822) );
  COND2X1 U6710 ( .A(n2449), .B(n5740), .C(n1556), .D(n5815), .Z(n5787) );
  COND1X1 U6711 ( .A(n5743), .B(n5742), .C(n5741), .Z(n5784) );
  CND2X1 U6712 ( .A(n5743), .B(n5742), .Z(n5783) );
  CFA1X1 U6713 ( .A(n5744), .B(n5745), .CI(n5746), .CO(n5786), .S(n5687) );
  CEO3X2 U6714 ( .A(n5787), .B(n5788), .C(n5786), .Z(n5821) );
  CENX2 U6715 ( .A(n5822), .B(n5821), .Z(n5747) );
  CENX2 U6716 ( .A(n2281), .B(n5747), .Z(n5839) );
  CNIVX2 U6717 ( .A(n5839), .Z(n5768) );
  CNIVX4 U6718 ( .A(n5748), .Z(n5751) );
  CND2X2 U6719 ( .A(n5752), .B(n5751), .Z(n5753) );
  CENX1 U6720 ( .A(h0[28]), .B(n2583), .Z(n5792) );
  COND2X1 U6721 ( .A(n6114), .B(n5754), .C(n3368), .D(n5792), .Z(n5856) );
  CENX1 U6722 ( .A(n7173), .B(n2512), .Z(n5818) );
  CENX1 U6723 ( .A(n7090), .B(n2443), .Z(n5798) );
  COND2X1 U6724 ( .A(n7126), .B(n5756), .C(n2433), .D(n5798), .Z(n5854) );
  CENX1 U6725 ( .A(n1264), .B(n5857), .Z(n5757) );
  COND1X1 U6726 ( .A(n5760), .B(n5759), .C(n5758), .Z(n5762) );
  CND2X1 U6727 ( .A(n5760), .B(n5759), .Z(n5761) );
  CENX1 U6728 ( .A(n6460), .B(h0[10]), .Z(n5863) );
  CENX1 U6729 ( .A(h0[8]), .B(n7202), .Z(n5862) );
  COND2X2 U6730 ( .A(n7203), .B(n5862), .C(n7205), .D(n5764), .Z(n5843) );
  CENX1 U6731 ( .A(n4922), .B(h0[26]), .Z(n5796) );
  CENX2 U6732 ( .A(n5768), .B(n5767), .Z(n5884) );
  COND1X2 U6733 ( .A(n5771), .B(n5770), .C(n5769), .Z(n5773) );
  CND2X1 U6734 ( .A(n5770), .B(n5771), .Z(n5772) );
  CND2X2 U6735 ( .A(n5772), .B(n5773), .Z(n5883) );
  CENX2 U6736 ( .A(n5884), .B(n5883), .Z(n5774) );
  CNIVXL U6737 ( .A(n5775), .Z(n5778) );
  CND2X1 U6738 ( .A(n5776), .B(n5778), .Z(n5781) );
  CND2X1 U6739 ( .A(n5776), .B(n2609), .Z(n5780) );
  CND2X1 U6740 ( .A(n5778), .B(n2609), .Z(n5779) );
  CND3X2 U6741 ( .A(n5781), .B(n5780), .C(n5779), .Z(n6267) );
  CIVX1 U6742 ( .A(n5787), .Z(n5782) );
  CND2X1 U6743 ( .A(n5786), .B(n5785), .Z(n5790) );
  CND2X2 U6744 ( .A(n5790), .B(n5789), .Z(n6046) );
  CENX1 U6745 ( .A(n6699), .B(h0[19]), .Z(n5996) );
  COND2X1 U6746 ( .A(n6765), .B(n5996), .C(n5791), .D(n6701), .Z(n5894) );
  COND2X1 U6747 ( .A(n6114), .B(n5792), .C(n3368), .D(n5910), .Z(n5893) );
  CENX1 U6748 ( .A(n5793), .B(h0[31]), .Z(n5913) );
  COND2X1 U6749 ( .A(n5911), .B(n5794), .C(n5912), .D(n5913), .Z(n5892) );
  CENX1 U6750 ( .A(n5893), .B(n5892), .Z(n5795) );
  CENX1 U6751 ( .A(n5894), .B(n5795), .Z(n6045) );
  CENX1 U6752 ( .A(n6118), .B(h0[27]), .Z(n5908) );
  COND2X1 U6753 ( .A(n2572), .B(n5796), .C(n2487), .D(n5908), .Z(n5891) );
  CENX1 U6754 ( .A(h0[13]), .B(n2659), .Z(n6002) );
  COND2X1 U6755 ( .A(n2295), .B(n5797), .C(n7114), .D(n6002), .Z(n5890) );
  CENX1 U6756 ( .A(n6103), .B(h0[7]), .Z(n5907) );
  CENX2 U6757 ( .A(n6045), .B(n6044), .Z(n5799) );
  CENX2 U6758 ( .A(n6046), .B(n5799), .Z(n5960) );
  CND2X1 U6759 ( .A(n5802), .B(n5804), .Z(n6054) );
  CND2IX1 U6760 ( .B(n5803), .A(n5802), .Z(n6056) );
  CND2X1 U6761 ( .A(n5807), .B(n5806), .Z(n5808) );
  CND2X2 U6762 ( .A(n5809), .B(n5808), .Z(n6059) );
  CND2XL U6763 ( .A(n2333), .B(n5812), .Z(n5814) );
  COND1X1 U6764 ( .A(n5812), .B(n2334), .C(n5810), .Z(n5813) );
  CND2X2 U6765 ( .A(n5814), .B(n5813), .Z(n5940) );
  CND2X2 U6766 ( .A(n5817), .B(n5816), .Z(n5941) );
  CENX1 U6767 ( .A(n7173), .B(h0[5]), .Z(n5906) );
  CENX2 U6768 ( .A(n5941), .B(n5918), .Z(n5819) );
  CENX2 U6769 ( .A(n5940), .B(n5819), .Z(n6057) );
  CENX1 U6770 ( .A(n6059), .B(n6057), .Z(n5820) );
  COND1X2 U6771 ( .A(n5822), .B(n5823), .C(n5821), .Z(n5825) );
  CND2X1 U6772 ( .A(n5823), .B(n5822), .Z(n5824) );
  CND2X2 U6773 ( .A(n5825), .B(n5824), .Z(n5958) );
  CIVX2 U6774 ( .A(n5831), .Z(n5827) );
  CIVX2 U6775 ( .A(n5830), .Z(n5826) );
  CND2X2 U6776 ( .A(n5827), .B(n5826), .Z(n5829) );
  CND2X1 U6777 ( .A(n5831), .B(n5830), .Z(n6086) );
  CND2X2 U6778 ( .A(n2508), .B(n6086), .Z(n5832) );
  CENX2 U6779 ( .A(n6090), .B(n5832), .Z(n5882) );
  CAN2XL U6780 ( .A(n5834), .B(n2492), .Z(n5837) );
  COND1XL U6781 ( .A(n2492), .B(n5834), .C(n5833), .Z(n5836) );
  CND2IX1 U6782 ( .B(n5837), .A(n5836), .Z(n6085) );
  COND1X2 U6783 ( .A(n5840), .B(n5839), .C(n5838), .Z(n5842) );
  CND2X1 U6784 ( .A(n5840), .B(n5839), .Z(n5841) );
  CND2X2 U6785 ( .A(n5842), .B(n5841), .Z(n6083) );
  CND2X2 U6786 ( .A(n5847), .B(n5846), .Z(n5936) );
  CND2X2 U6787 ( .A(n5848), .B(n5850), .Z(n5853) );
  CND2X2 U6788 ( .A(n2440), .B(n5850), .Z(n5852) );
  CND3X4 U6789 ( .A(n5853), .B(n5852), .C(n5851), .Z(n5937) );
  CIVX2 U6790 ( .A(n5854), .Z(n5855) );
  CIVX2 U6791 ( .A(n5855), .Z(n5858) );
  COND1X2 U6792 ( .A(n5857), .B(n5858), .C(n5856), .Z(n5860) );
  CND2X2 U6793 ( .A(n5860), .B(n5859), .Z(n5938) );
  CENX1 U6794 ( .A(n5937), .B(n5938), .Z(n5861) );
  CENX1 U6795 ( .A(n5936), .B(n5861), .Z(n5957) );
  CENX1 U6796 ( .A(n5927), .B(n7202), .Z(n5991) );
  COND2X1 U6797 ( .A(n7205), .B(n5862), .C(n7203), .D(n5991), .Z(n5978) );
  CENX1 U6798 ( .A(h0[15]), .B(n5932), .Z(n6004) );
  COND2X2 U6799 ( .A(n6972), .B(n6004), .C(n5864), .D(n6974), .Z(n5976) );
  CENX1 U6800 ( .A(n6828), .B(h0[17]), .Z(n5992) );
  CNR2X2 U6801 ( .A(n5869), .B(n5868), .Z(n5900) );
  CENX1 U6802 ( .A(n2660), .B(n2279), .Z(n5995) );
  COND2X1 U6803 ( .A(n6703), .B(n5870), .C(n6702), .D(n5995), .Z(n5897) );
  CIVX2 U6804 ( .A(n5897), .Z(n5871) );
  CENX2 U6805 ( .A(n5871), .B(n5900), .Z(n5872) );
  CENX2 U6806 ( .A(n5899), .B(n5872), .Z(n5944) );
  CND2X1 U6807 ( .A(n5874), .B(n5873), .Z(n5876) );
  CENX2 U6808 ( .A(n5944), .B(n5946), .Z(n5877) );
  CENX1 U6809 ( .A(n5945), .B(n5877), .Z(n5956) );
  CFA1X1 U6810 ( .A(n5880), .B(n5879), .CI(n5878), .CO(n5955), .S(n5840) );
  CEO3X2 U6811 ( .A(n6085), .B(n6083), .C(n6084), .Z(n5881) );
  CENX2 U6812 ( .A(n5881), .B(n5882), .Z(n7466) );
  COND1X2 U6813 ( .A(n5884), .B(n5885), .C(n2608), .Z(n5887) );
  CND2X1 U6814 ( .A(n5885), .B(n5884), .Z(n5886) );
  CND2X2 U6815 ( .A(n5887), .B(n5886), .Z(n7465) );
  CNR2X2 U6816 ( .A(n2446), .B(n7460), .Z(n6270) );
  CENX1 U6817 ( .A(n5888), .B(h0[24]), .Z(n5999) );
  COND2X1 U6818 ( .A(n2449), .B(n5999), .C(n1556), .D(n6100), .Z(n6163) );
  CENX1 U6819 ( .A(n6411), .B(h0[12]), .Z(n5986) );
  CENX1 U6820 ( .A(n6305), .B(h0[13]), .Z(n6096) );
  COND2X1 U6821 ( .A(n6969), .B(n5986), .C(n7171), .D(n6096), .Z(n6162) );
  CENX1 U6822 ( .A(h0[10]), .B(n7202), .Z(n5990) );
  CENX1 U6823 ( .A(h0[11]), .B(n7202), .Z(n6105) );
  COND2X1 U6824 ( .A(n7205), .B(n5990), .C(n7203), .D(n6105), .Z(n6161) );
  CFA1X1 U6825 ( .A(n5891), .B(n5890), .CI(n5889), .CO(n5961), .S(n6044) );
  CND2XL U6826 ( .A(n5893), .B(n5894), .Z(n5896) );
  COND1X1 U6827 ( .A(n5894), .B(n5893), .C(n5892), .Z(n5895) );
  CND2X2 U6828 ( .A(n5896), .B(n5895), .Z(n5963) );
  CIVX1 U6829 ( .A(n5900), .Z(n5898) );
  COND1X1 U6830 ( .A(n5898), .B(n5899), .C(n5897), .Z(n5902) );
  CND2IX1 U6831 ( .B(n5900), .A(n5899), .Z(n5901) );
  CND2X2 U6832 ( .A(n5902), .B(n5901), .Z(n5962) );
  COND1X2 U6833 ( .A(n5961), .B(n5963), .C(n5962), .Z(n5904) );
  CND2X2 U6834 ( .A(n5904), .B(n5903), .Z(n6109) );
  CENX1 U6835 ( .A(n7173), .B(n7674), .Z(n5905) );
  CENX1 U6836 ( .A(n7173), .B(h0[7]), .Z(n6102) );
  COND2X1 U6837 ( .A(n7228), .B(n5905), .C(n6102), .D(n2381), .Z(n6239) );
  CIVX2 U6838 ( .A(n6239), .Z(n6121) );
  COND2X1 U6839 ( .A(n7228), .B(n5906), .C(n5905), .D(n2382), .Z(n5971) );
  CENXL U6840 ( .A(n7090), .B(h0[8]), .Z(n5926) );
  COND2X1 U6841 ( .A(n2282), .B(n5907), .C(n2433), .D(n5926), .Z(n5970) );
  CENX1 U6842 ( .A(n6191), .B(h0[28]), .Z(n5933) );
  COND2X2 U6843 ( .A(n3368), .B(n5924), .C(n5910), .D(n6114), .Z(n5973) );
  CNIVX1 U6844 ( .A(n5973), .Z(n5920) );
  CIVX2 U6845 ( .A(n5920), .Z(n5917) );
  CND2X2 U6846 ( .A(n5912), .B(n5911), .Z(n5915) );
  CIVX2 U6847 ( .A(n5913), .Z(n5914) );
  CND2X2 U6848 ( .A(n5915), .B(n5914), .Z(n5972) );
  CIVX2 U6849 ( .A(n5972), .Z(n5916) );
  CND2X2 U6850 ( .A(n5917), .B(n5916), .Z(n5919) );
  CIVX2 U6851 ( .A(n5918), .Z(n5974) );
  CND2X2 U6852 ( .A(n5919), .B(n5974), .Z(n5922) );
  CND2XL U6853 ( .A(n5972), .B(n5920), .Z(n5921) );
  CND2X2 U6854 ( .A(n5922), .B(n5921), .Z(n6120) );
  CEO3X2 U6855 ( .A(n6121), .B(n6122), .C(n6120), .Z(n6111) );
  CEO3X2 U6856 ( .A(n6110), .B(n6109), .C(n6111), .Z(n6170) );
  CENX1 U6857 ( .A(n6699), .B(n2280), .Z(n6146) );
  CENX1 U6858 ( .A(n6409), .B(h0[20]), .Z(n5997) );
  COND2X2 U6859 ( .A(n6765), .B(n6146), .C(n6701), .D(n5997), .Z(n6140) );
  CIVX1 U6860 ( .A(n2282), .Z(n5925) );
  CND2IX1 U6861 ( .B(n5926), .A(n5925), .Z(n5930) );
  CENX1 U6862 ( .A(n6103), .B(n5927), .Z(n6104) );
  CND2IX2 U6863 ( .B(n6104), .A(n5928), .Z(n5929) );
  CND2X2 U6864 ( .A(n5930), .B(n5929), .Z(n6141) );
  CENX2 U6865 ( .A(n6140), .B(n6141), .Z(n5931) );
  CENXL U6866 ( .A(h0[18]), .B(n6828), .Z(n5993) );
  COND2X1 U6867 ( .A(n6831), .B(n5993), .C(n6829), .D(n6145), .Z(n6155) );
  CENX1 U6868 ( .A(n2659), .B(h0[14]), .Z(n6001) );
  CENX1 U6869 ( .A(h0[15]), .B(n2659), .Z(n6108) );
  COND2X1 U6870 ( .A(n2294), .B(n6001), .C(n7114), .D(n6108), .Z(n6154) );
  CENX1 U6871 ( .A(n2660), .B(h0[22]), .Z(n5994) );
  CENX1 U6872 ( .A(n2660), .B(h0[23]), .Z(n6106) );
  COND2X1 U6873 ( .A(n5994), .B(n6703), .C(n2515), .D(n6106), .Z(n6153) );
  CENX2 U6874 ( .A(n6148), .B(n6150), .Z(n5935) );
  CENX1 U6875 ( .A(n5932), .B(h0[17]), .Z(n6107) );
  CENX1 U6876 ( .A(h0[16]), .B(n5932), .Z(n6003) );
  COND2X1 U6877 ( .A(n6972), .B(n6107), .C(n6003), .D(n6974), .Z(n6156) );
  CENX1 U6878 ( .A(n6417), .B(h0[26]), .Z(n5983) );
  CENX1 U6879 ( .A(n6417), .B(h0[27]), .Z(n6097) );
  COND2X1 U6880 ( .A(n6418), .B(n5983), .C(n6293), .D(n6097), .Z(n6157) );
  CENX1 U6881 ( .A(n6118), .B(h0[29]), .Z(n6119) );
  COND2X1 U6882 ( .A(n2569), .B(n5933), .C(n2491), .D(n6119), .Z(n6158) );
  CENX1 U6883 ( .A(n6157), .B(n6158), .Z(n5934) );
  CENX1 U6884 ( .A(n6156), .B(n5934), .Z(n6149) );
  CIVX2 U6885 ( .A(n6049), .Z(n5952) );
  CND2X2 U6886 ( .A(n5943), .B(n5942), .Z(n6050) );
  CIVX2 U6887 ( .A(n6050), .Z(n5947) );
  CND2X2 U6888 ( .A(n5949), .B(n5948), .Z(n6052) );
  CND2X2 U6889 ( .A(n6052), .B(n6050), .Z(n5950) );
  CENX2 U6890 ( .A(n5954), .B(n5953), .Z(n6173) );
  CENX1 U6891 ( .A(n5962), .B(n5961), .Z(n5964) );
  CND2X1 U6892 ( .A(n5964), .B(n5963), .Z(n5968) );
  CIVX2 U6893 ( .A(n5963), .Z(n5966) );
  CIVX2 U6894 ( .A(n5964), .Z(n5965) );
  CND2X2 U6895 ( .A(n5966), .B(n5965), .Z(n5967) );
  CND2X4 U6896 ( .A(n5968), .B(n5967), .Z(n6041) );
  CFA1X1 U6897 ( .A(n5969), .B(n5970), .CI(n5971), .CO(n6122), .S(n6038) );
  CENX2 U6898 ( .A(n5973), .B(n5972), .Z(n5975) );
  CENX2 U6899 ( .A(n5975), .B(n5974), .Z(n6032) );
  CNIVX4 U6900 ( .A(n5976), .Z(n5979) );
  COND1X1 U6901 ( .A(n5979), .B(n5978), .C(n5977), .Z(n5981) );
  CND2X2 U6902 ( .A(n5979), .B(n5978), .Z(n5980) );
  CND2X2 U6903 ( .A(n5981), .B(n5980), .Z(n6033) );
  CENX2 U6904 ( .A(n6038), .B(n6037), .Z(n5982) );
  COND2X1 U6905 ( .A(n5985), .B(n6418), .C(n6293), .D(n5983), .Z(n6028) );
  CIVX2 U6906 ( .A(n5986), .Z(n5987) );
  CND2X2 U6907 ( .A(n1548), .B(n5987), .Z(n5988) );
  COND1X1 U6908 ( .A(n5989), .B(n6969), .C(n5988), .Z(n6027) );
  COND2X1 U6909 ( .A(n7205), .B(n5991), .C(n7203), .D(n5990), .Z(n6026) );
  COND2XL U6910 ( .A(n5993), .B(n6770), .C(n5992), .D(n6831), .Z(n6016) );
  COND2X2 U6911 ( .A(n5997), .B(n6765), .C(n5996), .D(n6701), .Z(n6018) );
  CENX1 U6912 ( .A(n6017), .B(n6018), .Z(n5998) );
  CENX1 U6913 ( .A(n6016), .B(n5998), .Z(n6011) );
  COND2X1 U6914 ( .A(n2449), .B(n6000), .C(n1557), .D(n5999), .Z(n6021) );
  COND2X1 U6915 ( .A(n6974), .B(n6004), .C(n6972), .D(n6003), .Z(n6022) );
  CNIVX1 U6916 ( .A(n6022), .Z(n6005) );
  CENX2 U6917 ( .A(n6012), .B(n6006), .Z(n6040) );
  CENX2 U6918 ( .A(n6007), .B(n6040), .Z(n6071) );
  CND2X2 U6919 ( .A(n6010), .B(n6009), .Z(n6174) );
  CND2X1 U6920 ( .A(n6013), .B(n6012), .Z(n6014) );
  CND2X2 U6921 ( .A(n6015), .B(n6014), .Z(n6167) );
  COND1XL U6922 ( .A(n6017), .B(n6018), .C(n6016), .Z(n6020) );
  CND2XL U6923 ( .A(n6018), .B(n6017), .Z(n6019) );
  CND2X1 U6924 ( .A(n6020), .B(n6019), .Z(n6127) );
  CND2X2 U6925 ( .A(n6025), .B(n6024), .Z(n6125) );
  COND1X1 U6926 ( .A(n6027), .B(n6028), .C(n6026), .Z(n6030) );
  CND2XL U6927 ( .A(n6028), .B(n6027), .Z(n6029) );
  CND2X1 U6928 ( .A(n6030), .B(n6029), .Z(n6126) );
  CENX1 U6929 ( .A(n6125), .B(n6126), .Z(n6031) );
  CENX1 U6930 ( .A(n6127), .B(n6031), .Z(n6166) );
  COND1X2 U6931 ( .A(n6033), .B(n6034), .C(n6038), .Z(n6036) );
  CND2X2 U6932 ( .A(n6036), .B(n6035), .Z(n6165) );
  COND1X2 U6933 ( .A(n6041), .B(n6040), .C(n6039), .Z(n6043) );
  CND2X2 U6934 ( .A(n6041), .B(n6040), .Z(n6042) );
  CND2X4 U6935 ( .A(n6043), .B(n6042), .Z(n6136) );
  COND1X1 U6936 ( .A(n6046), .B(n6045), .C(n6044), .Z(n6048) );
  CND2X2 U6937 ( .A(n6048), .B(n6047), .Z(n6075) );
  CENX2 U6938 ( .A(n6050), .B(n6049), .Z(n6051) );
  CENX2 U6939 ( .A(n6052), .B(n6051), .Z(n6074) );
  CIVX1 U6940 ( .A(n6059), .Z(n6053) );
  CND4X1 U6941 ( .A(n6056), .B(n6055), .C(n6054), .D(n6053), .Z(n6058) );
  CND2X2 U6942 ( .A(n6058), .B(n6057), .Z(n6063) );
  CNIVXL U6943 ( .A(n6059), .Z(n6060) );
  CND2X2 U6944 ( .A(n6061), .B(n6060), .Z(n6062) );
  CND2X2 U6945 ( .A(n6063), .B(n6062), .Z(n6073) );
  COND1X2 U6946 ( .A(n6075), .B(n6074), .C(n6073), .Z(n6065) );
  CND2X2 U6947 ( .A(n6074), .B(n6075), .Z(n6064) );
  CENX2 U6948 ( .A(n6136), .B(n6135), .Z(n6066) );
  CEO3X1 U6949 ( .A(n6173), .B(n6174), .C(n6172), .Z(n6274) );
  COND1X2 U6950 ( .A(n6067), .B(n6083), .C(n6084), .Z(n6069) );
  CND2X2 U6951 ( .A(n6069), .B(n6068), .Z(n6081) );
  CIVX2 U6952 ( .A(n6081), .Z(n6079) );
  CEO3X2 U6953 ( .A(n6072), .B(n6071), .C(n6070), .Z(n6080) );
  CEO3X2 U6954 ( .A(n6075), .B(n6073), .C(n6074), .Z(n6082) );
  CNR2X2 U6955 ( .A(n6080), .B(n6082), .Z(n6078) );
  CIVXL U6956 ( .A(n6082), .Z(n6076) );
  CND2IX2 U6957 ( .B(n6076), .A(n6080), .Z(n6077) );
  COND1X2 U6958 ( .A(n6079), .B(n6078), .C(n6077), .Z(n6273) );
  CNR2X2 U6959 ( .A(n6274), .B(n6273), .Z(n7018) );
  CEO3X2 U6960 ( .A(n6082), .B(n6081), .C(n6080), .Z(n6272) );
  CND2XL U6961 ( .A(n6087), .B(n6086), .Z(n6088) );
  CND3X2 U6962 ( .A(n6093), .B(n6092), .C(n6091), .Z(n6271) );
  CIVX2 U6963 ( .A(n6209), .Z(n6094) );
  CENX1 U6964 ( .A(n6417), .B(h0[28]), .Z(n6210) );
  COR2X1 U6965 ( .A(n6418), .B(n6097), .Z(n6098) );
  CND2X2 U6966 ( .A(n6099), .B(n6098), .Z(n6233) );
  CENX1 U6967 ( .A(n6490), .B(h0[26]), .Z(n6213) );
  COND2X1 U6968 ( .A(n2449), .B(n6100), .C(n1557), .D(n6213), .Z(n6231) );
  CENX2 U6969 ( .A(n6233), .B(n6231), .Z(n6101) );
  CENX1 U6970 ( .A(n7173), .B(h0[8]), .Z(n6186) );
  COND2X1 U6971 ( .A(n7228), .B(n6102), .C(n6186), .D(n2381), .Z(n6204) );
  CENX1 U6972 ( .A(n6103), .B(h0[10]), .Z(n6194) );
  COND2X1 U6973 ( .A(n2282), .B(n6104), .C(n2433), .D(n6194), .Z(n6203) );
  CENX1 U6974 ( .A(h0[12]), .B(n7062), .Z(n6206) );
  COND2X1 U6975 ( .A(n7217), .B(n6105), .C(n7203), .D(n6206), .Z(n6202) );
  CENX1 U6976 ( .A(n2660), .B(h0[24]), .Z(n6205) );
  COND2X1 U6977 ( .A(n6703), .B(n6106), .C(n2514), .D(n6205), .Z(n6230) );
  COND2X1 U6978 ( .A(n6974), .B(n6107), .C(n6184), .D(n6972), .Z(n6229) );
  CENX1 U6979 ( .A(h0[16]), .B(n2659), .Z(n6212) );
  COND2X1 U6980 ( .A(n2295), .B(n6108), .C(n7114), .D(n6212), .Z(n6228) );
  COND1X1 U6981 ( .A(n1222), .B(n6111), .C(n6109), .Z(n6113) );
  CND2X1 U6982 ( .A(n1222), .B(n6111), .Z(n6112) );
  CND2X2 U6983 ( .A(n6113), .B(n6112), .Z(n6258) );
  CIVX2 U6984 ( .A(n6115), .Z(n6116) );
  CND2X2 U6985 ( .A(n6117), .B(n6116), .Z(n6236) );
  CENX1 U6986 ( .A(n6118), .B(h0[30]), .Z(n6192) );
  COND2X1 U6987 ( .A(n2574), .B(n6119), .C(n2490), .D(n6192), .Z(n6237) );
  CEO3X1 U6988 ( .A(n6236), .B(n6237), .C(n6239), .Z(n6197) );
  CND2X2 U6989 ( .A(n6124), .B(n6123), .Z(n6198) );
  CND2X2 U6990 ( .A(n6129), .B(n6128), .Z(n6199) );
  CEO3X2 U6991 ( .A(n6197), .B(n6198), .C(n6199), .Z(n6260) );
  CIVX2 U6992 ( .A(n6135), .Z(n6132) );
  CIVX2 U6993 ( .A(n6136), .Z(n6131) );
  CND2X2 U6994 ( .A(n6132), .B(n6131), .Z(n6133) );
  CND2X2 U6995 ( .A(n6134), .B(n6133), .Z(n6139) );
  CND2X2 U6996 ( .A(n2441), .B(n6137), .Z(n6138) );
  CND2X4 U6997 ( .A(n6139), .B(n6138), .Z(n6276) );
  CND2X1 U6998 ( .A(n6141), .B(n6142), .Z(n6144) );
  CND2X2 U6999 ( .A(n6144), .B(n6143), .Z(n6181) );
  CENX1 U7000 ( .A(n6769), .B(h0[20]), .Z(n6193) );
  COND2X1 U7001 ( .A(n2420), .B(n6145), .C(n6770), .D(n6193), .Z(n6179) );
  CENX1 U7002 ( .A(n6699), .B(h0[22]), .Z(n6188) );
  COND1X1 U7003 ( .A(n6149), .B(n6150), .C(n6148), .Z(n6152) );
  CND2X1 U7004 ( .A(n6150), .B(n6149), .Z(n6151) );
  CND2X2 U7005 ( .A(n6152), .B(n6151), .Z(n6225) );
  CFA1X1 U7006 ( .A(n6155), .B(n6154), .CI(n6153), .CO(n6245), .S(n6150) );
  CND2X2 U7007 ( .A(n6160), .B(n6159), .Z(n6246) );
  CFA1X1 U7008 ( .A(n6163), .B(n6162), .CI(n6161), .CO(n6244), .S(n6110) );
  CENX2 U7009 ( .A(n6246), .B(n6244), .Z(n6164) );
  CENX2 U7010 ( .A(n6164), .B(n6245), .Z(n6223) );
  CEO3X2 U7011 ( .A(n6224), .B(n6225), .C(n6223), .Z(n6217) );
  CND2X2 U7012 ( .A(n6170), .B(n6169), .Z(n6215) );
  CND2X2 U7013 ( .A(n6216), .B(n6215), .Z(n6220) );
  CEO3X1 U7014 ( .A(n6277), .B(n6276), .C(n2407), .Z(n6178) );
  CND2X1 U7015 ( .A(n6174), .B(n6172), .Z(n6177) );
  CND2X1 U7016 ( .A(n6174), .B(n2502), .Z(n6175) );
  CND3X2 U7017 ( .A(n6177), .B(n6176), .C(n6175), .Z(n6278) );
  CNR2X2 U7018 ( .A(n6178), .B(n6278), .Z(n7028) );
  CND2X1 U7019 ( .A(n6181), .B(n6180), .Z(n6182) );
  CND2X2 U7020 ( .A(n6183), .B(n6182), .Z(n6327) );
  CIVX2 U7021 ( .A(n6327), .Z(n6196) );
  COND2X1 U7022 ( .A(n7065), .B(n6184), .C(n2477), .D(n6302), .Z(n6319) );
  CENX1 U7023 ( .A(n7173), .B(n6185), .Z(n6310) );
  COND2X1 U7024 ( .A(n7228), .B(n6186), .C(n7301), .D(n6310), .Z(n6187) );
  COND2X2 U7025 ( .A(n6765), .B(n6300), .C(n6701), .D(n6188), .Z(n6320) );
  CENX1 U7026 ( .A(n6444), .B(n6320), .Z(n6189) );
  CIVX2 U7027 ( .A(n6189), .Z(n6190) );
  CENX1 U7028 ( .A(n6319), .B(n6190), .Z(n6324) );
  CENX1 U7029 ( .A(n6118), .B(h0[31]), .Z(n6292) );
  COND2X2 U7030 ( .A(n2489), .B(n6292), .C(n2576), .D(n6192), .Z(n6352) );
  CENX1 U7031 ( .A(n6769), .B(n2279), .Z(n6351) );
  COND2X1 U7032 ( .A(n2420), .B(n6193), .C(n6829), .D(n6351), .Z(n6353) );
  CENXL U7033 ( .A(n7090), .B(h0[11]), .Z(n6308) );
  COND2X1 U7034 ( .A(n2282), .B(n6194), .C(n2433), .D(n6308), .Z(n6354) );
  CEO3X1 U7035 ( .A(n6352), .B(n6353), .C(n6354), .Z(n6326) );
  CENX2 U7036 ( .A(n6196), .B(n6195), .Z(n6363) );
  COND1X1 U7037 ( .A(n2439), .B(n6199), .C(n6198), .Z(n6201) );
  CND2X1 U7038 ( .A(n6199), .B(n2439), .Z(n6200) );
  CND2X2 U7039 ( .A(n6201), .B(n6200), .Z(n6362) );
  CFA1X1 U7040 ( .A(n6204), .B(n6203), .CI(n6202), .CO(n6348), .S(n6251) );
  CENX1 U7041 ( .A(n2660), .B(h0[25]), .Z(n6304) );
  COND2X1 U7042 ( .A(n6703), .B(n6205), .C(n2514), .D(n6304), .Z(n6314) );
  COND2X1 U7043 ( .A(n7217), .B(n6206), .C(n7203), .D(n6309), .Z(n6312) );
  CENX1 U7044 ( .A(n6305), .B(h0[15]), .Z(n6306) );
  CIVX2 U7045 ( .A(n6306), .Z(n6207) );
  CND2X1 U7046 ( .A(n1549), .B(n6207), .Z(n6208) );
  CENX1 U7047 ( .A(n6417), .B(h0[29]), .Z(n6295) );
  COND2X1 U7048 ( .A(n6211), .B(n6210), .C(n5984), .D(n6295), .Z(n6359) );
  CENX1 U7049 ( .A(h0[17]), .B(n2659), .Z(n6301) );
  CENX1 U7050 ( .A(n6490), .B(h0[27]), .Z(n6303) );
  COND2X1 U7051 ( .A(n2449), .B(n6213), .C(n1556), .D(n6303), .Z(n6357) );
  CEO3X2 U7052 ( .A(n6348), .B(n6346), .C(n6347), .Z(n6360) );
  CND2X1 U7053 ( .A(n2614), .B(n6215), .Z(n6218) );
  CND2X1 U7054 ( .A(n6220), .B(n6219), .Z(n6221) );
  CND2X2 U7055 ( .A(n6222), .B(n6221), .Z(n6286) );
  CND2X1 U7056 ( .A(n6225), .B(n6224), .Z(n6226) );
  CND2X2 U7057 ( .A(n6227), .B(n6226), .Z(n6332) );
  CFA1X1 U7058 ( .A(n6230), .B(n6229), .CI(n6228), .CO(n6341), .S(n6250) );
  COND1X1 U7059 ( .A(n6232), .B(n6233), .C(n6231), .Z(n6235) );
  CND2X2 U7060 ( .A(n6235), .B(n6234), .Z(n6342) );
  CNIVX4 U7061 ( .A(n6236), .Z(n6238) );
  CIVX2 U7062 ( .A(n6238), .Z(n6240) );
  CND2IX1 U7063 ( .B(n6240), .A(n6239), .Z(n6241) );
  CND2X2 U7064 ( .A(n6242), .B(n6241), .Z(n6343) );
  CENX2 U7065 ( .A(n6342), .B(n6343), .Z(n6243) );
  CENX2 U7066 ( .A(n6341), .B(n6243), .Z(n6338) );
  CIVX2 U7067 ( .A(n6338), .Z(n6257) );
  CND2X2 U7068 ( .A(n6248), .B(n6247), .Z(n6337) );
  CND2X1 U7069 ( .A(n6251), .B(n6253), .Z(n6249) );
  CND2IX1 U7070 ( .B(n6250), .A(n6249), .Z(n6255) );
  CIVX2 U7071 ( .A(n6251), .Z(n6252) );
  CND2IX1 U7072 ( .B(n6253), .A(n6252), .Z(n6254) );
  CND2X2 U7073 ( .A(n6255), .B(n6254), .Z(n6335) );
  CENX2 U7074 ( .A(n6337), .B(n6335), .Z(n6256) );
  CENX2 U7075 ( .A(n6257), .B(n6256), .Z(n6330) );
  COND1X1 U7076 ( .A(n6259), .B(n6260), .C(n6258), .Z(n6262) );
  CND2X2 U7077 ( .A(n6261), .B(n6262), .Z(n6331) );
  CEO3X2 U7078 ( .A(n6332), .B(n6330), .C(n6331), .Z(n6289) );
  CEO3X1 U7079 ( .A(n6288), .B(n6286), .C(n6289), .Z(n6281) );
  COND1X1 U7080 ( .A(n6277), .B(n6275), .C(n6276), .Z(n6264) );
  CNR2X2 U7081 ( .A(n2286), .B(n6280), .Z(n7046) );
  CND2X2 U7082 ( .A(n7035), .B(n6283), .Z(n6285) );
  COND1X2 U7083 ( .A(n7306), .B(n7309), .C(n7307), .Z(n7472) );
  CND2X2 U7084 ( .A(n2308), .B(n6267), .Z(n7470) );
  COND1X2 U7085 ( .A(n7470), .B(n6268), .C(n7468), .Z(n6269) );
  CND2X2 U7086 ( .A(n6272), .B(n6271), .Z(n7021) );
  CND2X1 U7087 ( .A(n6274), .B(n6273), .Z(n7019) );
  CEO3X2 U7088 ( .A(n6277), .B(n6276), .C(n2407), .Z(n6279) );
  CND2X2 U7089 ( .A(n6279), .B(n6278), .Z(n7039) );
  COND1X2 U7090 ( .A(n7046), .B(n7039), .C(n7047), .Z(n6282) );
  CND2X1 U7091 ( .A(n6289), .B(n6288), .Z(n6290) );
  CIVX2 U7092 ( .A(n6447), .Z(n6299) );
  CENX1 U7093 ( .A(n2597), .B(h0[30]), .Z(n6419) );
  CNR2X1 U7094 ( .A(n6419), .B(n6293), .Z(n6294) );
  CIVX2 U7095 ( .A(n6294), .Z(n6297) );
  COR2X1 U7096 ( .A(n6418), .B(n6295), .Z(n6296) );
  CND2X2 U7097 ( .A(n6297), .B(n6296), .Z(n6445) );
  CENX2 U7098 ( .A(n6445), .B(n6444), .Z(n6298) );
  CENX2 U7099 ( .A(n6299), .B(n6298), .Z(n6394) );
  CENX1 U7100 ( .A(n6699), .B(h0[24]), .Z(n6410) );
  CENX1 U7101 ( .A(h0[18]), .B(n7092), .Z(n6405) );
  COND2X1 U7102 ( .A(n6301), .B(n2294), .C(n6405), .D(n7114), .Z(n6401) );
  CENX1 U7103 ( .A(n6490), .B(h0[28]), .Z(n6407) );
  COND2X1 U7104 ( .A(n2449), .B(n6303), .C(n1556), .D(n6407), .Z(n6404) );
  CENX1 U7105 ( .A(n2660), .B(h0[26]), .Z(n6406) );
  COND2X1 U7106 ( .A(n6703), .B(n6304), .C(n2514), .D(n6406), .Z(n6403) );
  CENX1 U7107 ( .A(n6305), .B(h0[16]), .Z(n6414) );
  COND2X1 U7108 ( .A(n4991), .B(n6306), .C(n7171), .D(n6414), .Z(n6402) );
  CENX1 U7109 ( .A(n6103), .B(h0[12]), .Z(n6420) );
  COND2X1 U7110 ( .A(n2282), .B(n6308), .C(n6420), .D(n7124), .Z(n6397) );
  CENX1 U7111 ( .A(h0[14]), .B(n7062), .Z(n6408) );
  COND2X2 U7112 ( .A(n7203), .B(n6408), .C(n6309), .D(n7205), .Z(n6398) );
  CENX1 U7113 ( .A(n7173), .B(h0[10]), .Z(n6442) );
  COND2X1 U7114 ( .A(n7228), .B(n6310), .C(n6442), .D(n2381), .Z(n6399) );
  CENX1 U7115 ( .A(n6398), .B(n6399), .Z(n6311) );
  CENX1 U7116 ( .A(n6397), .B(n6311), .Z(n6436) );
  CND2X2 U7117 ( .A(n6316), .B(n6315), .Z(n6435) );
  CNR2X2 U7118 ( .A(n6444), .B(n6320), .Z(n6317) );
  CIVX2 U7119 ( .A(n6317), .Z(n6318) );
  CND2X2 U7120 ( .A(n6319), .B(n6318), .Z(n6322) );
  CND2XL U7121 ( .A(n6320), .B(n6444), .Z(n6321) );
  CND2X2 U7122 ( .A(n6322), .B(n6321), .Z(n6434) );
  CENX2 U7123 ( .A(n6435), .B(n6434), .Z(n6323) );
  CENX2 U7124 ( .A(n6436), .B(n6323), .Z(n6427) );
  COND1X1 U7125 ( .A(n6326), .B(n6327), .C(n6325), .Z(n6329) );
  CND2X1 U7126 ( .A(n6327), .B(n6326), .Z(n6328) );
  CND2X2 U7127 ( .A(n6329), .B(n6328), .Z(n6426) );
  CND2X2 U7128 ( .A(n6334), .B(n6333), .Z(n6453) );
  CIVX2 U7129 ( .A(n6335), .Z(n6336) );
  COND1X2 U7130 ( .A(n6337), .B(n6338), .C(n6336), .Z(n6340) );
  CND2X2 U7131 ( .A(n6338), .B(n6337), .Z(n6339) );
  CND2X2 U7132 ( .A(n6340), .B(n6339), .Z(n6422) );
  CND2X2 U7133 ( .A(n6345), .B(n6344), .Z(n6433) );
  CENX1 U7134 ( .A(n2454), .B(h0[22]), .Z(n6443) );
  COND2X1 U7135 ( .A(n2420), .B(n6351), .C(n6829), .D(n6443), .Z(n6438) );
  COND1X1 U7136 ( .A(n6353), .B(n6354), .C(n6352), .Z(n6356) );
  CND2X2 U7137 ( .A(n6356), .B(n6355), .Z(n6437) );
  CEO3X2 U7138 ( .A(n6438), .B(n6437), .C(n6439), .Z(n6431) );
  CNIVX4 U7139 ( .A(n6360), .Z(n6361) );
  COND1X2 U7140 ( .A(n6362), .B(n6363), .C(n6361), .Z(n6365) );
  CND2X2 U7141 ( .A(n6363), .B(n6362), .Z(n6364) );
  CND2X4 U7142 ( .A(n6365), .B(n6364), .Z(n6423) );
  CEO3X2 U7143 ( .A(n6422), .B(n6421), .C(n6423), .Z(n6455) );
  CIVX2 U7144 ( .A(n6368), .Z(n6366) );
  CND2X2 U7145 ( .A(n2296), .B(n6366), .Z(n7453) );
  CAN2XL U7146 ( .A(n7453), .B(n7454), .Z(n6369) );
  CENXL U7147 ( .A(n2359), .B(n6369), .Z(N55) );
  CND2X1 U7148 ( .A(n6386), .B(n6385), .Z(n6391) );
  CANR1XL U7149 ( .A(n6389), .B(n6388), .C(n6387), .Z(n6390) );
  CEOXL U7150 ( .A(n6391), .B(n6390), .Z(N27) );
  CND2X2 U7151 ( .A(n6396), .B(n6395), .Z(n6607) );
  CND2X1 U7152 ( .A(n6399), .B(n6398), .Z(n6400) );
  CFA1X1 U7153 ( .A(n6404), .B(n6402), .CI(n6403), .CO(n6500), .S(n6392) );
  CENX1 U7154 ( .A(h0[19]), .B(n6970), .Z(n6470) );
  CENX1 U7155 ( .A(n2660), .B(h0[27]), .Z(n6472) );
  COND2X1 U7156 ( .A(n6406), .B(n6703), .C(n2515), .D(n6472), .Z(n6515) );
  CENX1 U7157 ( .A(n6490), .B(h0[29]), .Z(n6526) );
  COND2X1 U7158 ( .A(n2449), .B(n6407), .C(n1557), .D(n6526), .Z(n6514) );
  CENX1 U7159 ( .A(h0[15]), .B(n7062), .Z(n6498) );
  COND2X1 U7160 ( .A(n7205), .B(n6408), .C(n7203), .D(n6498), .Z(n6508) );
  CENX1 U7161 ( .A(n6409), .B(h0[25]), .Z(n6480) );
  COND2X1 U7162 ( .A(n1582), .B(n6410), .C(n6765), .D(n6480), .Z(n6510) );
  CENX1 U7163 ( .A(n6508), .B(n6510), .Z(n6415) );
  CENX1 U7164 ( .A(n6411), .B(h0[17]), .Z(n6467) );
  CIVX2 U7165 ( .A(n6467), .Z(n6412) );
  CND2IX1 U7166 ( .B(n7171), .A(n6412), .Z(n6413) );
  COND2X1 U7167 ( .A(n6974), .B(n6416), .C(n6972), .D(n6481), .Z(n6513) );
  CENX1 U7168 ( .A(n6417), .B(h0[31]), .Z(n6521) );
  CENX1 U7169 ( .A(n6103), .B(h0[13]), .Z(n6496) );
  COND1X2 U7170 ( .A(n6422), .B(n6423), .C(n6421), .Z(n6425) );
  CND2X2 U7171 ( .A(n6423), .B(n6422), .Z(n6424) );
  CND2X2 U7172 ( .A(n6425), .B(n6424), .Z(n6920) );
  CND2X2 U7173 ( .A(n6430), .B(n6429), .Z(n6911) );
  CFA1X1 U7174 ( .A(n6433), .B(n6432), .CI(n6431), .CO(n6910), .S(n6421) );
  CND2X2 U7175 ( .A(n6441), .B(n6440), .Z(n6597) );
  CENX1 U7176 ( .A(n7173), .B(h0[11]), .Z(n6494) );
  COND2X1 U7177 ( .A(n7228), .B(n6442), .C(n6494), .D(n2382), .Z(n6558) );
  CIVX2 U7178 ( .A(n6558), .Z(n6528) );
  CENX1 U7179 ( .A(n6769), .B(h0[23]), .Z(n6478) );
  COND2X1 U7180 ( .A(n2420), .B(n6443), .C(n6770), .D(n6478), .Z(n6504) );
  CENX1 U7181 ( .A(n6528), .B(n6504), .Z(n6450) );
  CIVX2 U7182 ( .A(n6444), .Z(n6446) );
  COND1X2 U7183 ( .A(n6447), .B(n6446), .C(n6445), .Z(n6449) );
  CND2X2 U7184 ( .A(n6449), .B(n6448), .Z(n6505) );
  CENX2 U7185 ( .A(n6450), .B(n6505), .Z(n6598) );
  CENX2 U7186 ( .A(n6597), .B(n6598), .Z(n6451) );
  CENX2 U7187 ( .A(n6596), .B(n6451), .Z(n6909) );
  CENX2 U7188 ( .A(n6910), .B(n6909), .Z(n6452) );
  CENX2 U7189 ( .A(n6911), .B(n6452), .Z(n6921) );
  CEO3X2 U7190 ( .A(n6919), .B(n6920), .C(n6921), .Z(n6931) );
  CIVX2 U7191 ( .A(n6931), .Z(n6459) );
  COND1X2 U7192 ( .A(n6454), .B(n6455), .C(n6453), .Z(n6457) );
  CND2X2 U7193 ( .A(n6457), .B(n6456), .Z(n6930) );
  CIVX2 U7194 ( .A(n6930), .Z(n6458) );
  CND2X2 U7195 ( .A(n6459), .B(n6458), .Z(n7457) );
  CND2X2 U7196 ( .A(n7453), .B(n7457), .Z(n7383) );
  CIVX2 U7197 ( .A(n7383), .Z(n7373) );
  CENX1 U7198 ( .A(n7173), .B(h0[13]), .Z(n6553) );
  CENX1 U7199 ( .A(n7173), .B(h0[14]), .Z(n6645) );
  CENX1 U7200 ( .A(n6103), .B(h0[15]), .Z(n6462) );
  CENX1 U7201 ( .A(n6103), .B(h0[16]), .Z(n6650) );
  CENX1 U7202 ( .A(h0[17]), .B(n7062), .Z(n6461) );
  CENX1 U7203 ( .A(h0[18]), .B(n7202), .Z(n6642) );
  COND2X1 U7204 ( .A(n7205), .B(n6461), .C(n7203), .D(n6642), .Z(n6620) );
  CENX1 U7205 ( .A(n6769), .B(h0[24]), .Z(n6477) );
  COND2X1 U7206 ( .A(n2420), .B(n6477), .C(n6829), .D(n6492), .Z(n6466) );
  COND2X1 U7207 ( .A(n2397), .B(n6469), .C(n7171), .D(n6583), .Z(n6465) );
  CENX1 U7208 ( .A(n2279), .B(n6970), .Z(n6585) );
  CENX1 U7209 ( .A(h0[20]), .B(n6970), .Z(n6471) );
  COND2X1 U7210 ( .A(n7114), .B(n6585), .C(n6471), .D(n2295), .Z(n6464) );
  CENX1 U7211 ( .A(h0[16]), .B(n7062), .Z(n6497) );
  CENX1 U7212 ( .A(n6699), .B(h0[27]), .Z(n6487) );
  CENX1 U7213 ( .A(n6699), .B(h0[26]), .Z(n6479) );
  CENX1 U7214 ( .A(n7090), .B(h0[14]), .Z(n6495) );
  COND2X1 U7215 ( .A(n6495), .B(n7126), .C(n2433), .D(n6462), .Z(n6539) );
  CENX1 U7216 ( .A(n6622), .B(n6624), .Z(n6463) );
  CENX1 U7217 ( .A(n6623), .B(n6463), .Z(n6653) );
  CFA1X1 U7218 ( .A(n6466), .B(n6465), .CI(n6464), .CO(n6622), .S(n6567) );
  COND2X2 U7219 ( .A(n7171), .B(n6469), .C(n4991), .D(n6467), .Z(n6530) );
  CENX1 U7220 ( .A(n2660), .B(h0[28]), .Z(n6488) );
  COND2X2 U7221 ( .A(n2514), .B(n6488), .C(n6473), .D(n6472), .Z(n6531) );
  CND2X2 U7222 ( .A(n6476), .B(n6475), .Z(n6565) );
  CIVX2 U7223 ( .A(n6565), .Z(n6483) );
  COND2X1 U7224 ( .A(n6831), .B(n6478), .C(n6770), .D(n6477), .Z(n6520) );
  COND2X1 U7225 ( .A(n6480), .B(n1582), .C(n6765), .D(n6479), .Z(n6519) );
  CIVX2 U7226 ( .A(n6564), .Z(n6482) );
  CND2X2 U7227 ( .A(n6483), .B(n6482), .Z(n6484) );
  CND2X2 U7228 ( .A(n6567), .B(n6484), .Z(n6486) );
  CND2X2 U7229 ( .A(n6486), .B(n6485), .Z(n6652) );
  CENX1 U7230 ( .A(n6699), .B(h0[28]), .Z(n6644) );
  COND2X1 U7231 ( .A(n6701), .B(n6487), .C(n6765), .D(n6644), .Z(n6629) );
  CENX1 U7232 ( .A(n2660), .B(h0[29]), .Z(n6579) );
  COND2X1 U7233 ( .A(n6703), .B(n6488), .C(n2515), .D(n6579), .Z(n6547) );
  COND2X1 U7234 ( .A(n6974), .B(n6489), .C(n6972), .D(n6584), .Z(n6546) );
  CENX1 U7235 ( .A(n6490), .B(h0[30]), .Z(n6524) );
  CENX1 U7236 ( .A(n6491), .B(h0[31]), .Z(n6575) );
  COND2X1 U7237 ( .A(n2449), .B(n6524), .C(n1556), .D(n6575), .Z(n6545) );
  CENX1 U7238 ( .A(n2454), .B(h0[26]), .Z(n6646) );
  COND2X1 U7239 ( .A(n2420), .B(n6492), .C(n6829), .D(n6646), .Z(n6627) );
  CENX1 U7240 ( .A(n7173), .B(h0[12]), .Z(n6554) );
  COND2X1 U7241 ( .A(n7228), .B(n6494), .C(n6554), .D(n2382), .Z(n6557) );
  COND2X1 U7242 ( .A(n2282), .B(n6496), .C(n7124), .D(n6495), .Z(n6556) );
  COND2X1 U7243 ( .A(n7205), .B(n6498), .C(n7203), .D(n6497), .Z(n6555) );
  CND2X2 U7244 ( .A(n6507), .B(n6506), .Z(n6601) );
  COND1X1 U7245 ( .A(n6509), .B(n6510), .C(n6508), .Z(n6512) );
  CND2X1 U7246 ( .A(n6510), .B(n6509), .Z(n6511) );
  CND2X2 U7247 ( .A(n6512), .B(n6511), .Z(n6542) );
  CFA1X1 U7248 ( .A(n6515), .B(n6516), .CI(n6514), .CO(n6541), .S(n6536) );
  CENX2 U7249 ( .A(n6540), .B(n6541), .Z(n6517) );
  CENX2 U7250 ( .A(n6542), .B(n6517), .Z(n6906) );
  CFA1X1 U7251 ( .A(n6520), .B(n6519), .CI(n6518), .CO(n6564), .S(n6570) );
  CANR1X2 U7252 ( .A(n6523), .B(n6522), .C(n6521), .Z(n6559) );
  COND2X1 U7253 ( .A(n6527), .B(n6526), .C(n1557), .D(n6524), .Z(n6560) );
  CENX1 U7254 ( .A(n6528), .B(n6560), .Z(n6529) );
  CENX1 U7255 ( .A(n6559), .B(n6529), .Z(n6568) );
  CENX2 U7256 ( .A(n2403), .B(n6532), .Z(n6569) );
  CENX2 U7257 ( .A(n6568), .B(n6569), .Z(n6533) );
  CFA1X1 U7258 ( .A(n6536), .B(n6535), .CI(n6534), .CO(n6905), .S(n6604) );
  COND1X1 U7259 ( .A(n6906), .B(n6908), .C(n6905), .Z(n6538) );
  CND2X1 U7260 ( .A(n6908), .B(n6906), .Z(n6537) );
  CND2X2 U7261 ( .A(n6538), .B(n6537), .Z(n6586) );
  COND1X2 U7262 ( .A(n6541), .B(n6542), .C(n6540), .Z(n6544) );
  CND2X2 U7263 ( .A(n6542), .B(n6541), .Z(n6543) );
  CND2X2 U7264 ( .A(n6544), .B(n6543), .Z(n6551) );
  CFA1X1 U7265 ( .A(n6547), .B(n6546), .CI(n6545), .CO(n6628), .S(n6550) );
  COND2X1 U7266 ( .A(n7228), .B(n6554), .C(n6553), .D(n2382), .Z(n6619) );
  CIVX2 U7267 ( .A(n6619), .Z(n6582) );
  CFA1X1 U7268 ( .A(n6557), .B(n6556), .CI(n6555), .CO(n6581), .S(n6603) );
  CND2IXL U7269 ( .B(n6559), .A(n6558), .Z(n6563) );
  CND2X2 U7270 ( .A(n6528), .B(n6559), .Z(n6561) );
  CND2X1 U7271 ( .A(n6561), .B(n6560), .Z(n6562) );
  CND2X2 U7272 ( .A(n6563), .B(n6562), .Z(n6580) );
  CENX2 U7273 ( .A(n6567), .B(n6566), .Z(n6591) );
  COND1X1 U7274 ( .A(n6569), .B(n6570), .C(n6568), .Z(n6572) );
  CND2X2 U7275 ( .A(n6572), .B(n6571), .Z(n6590) );
  CND2X1 U7276 ( .A(n6591), .B(n6589), .Z(n6573) );
  CND2X2 U7277 ( .A(n6574), .B(n6573), .Z(n6633) );
  CIVXL U7278 ( .A(n6575), .Z(n6578) );
  CND2X1 U7279 ( .A(n6578), .B(n6577), .Z(n6618) );
  CENX1 U7280 ( .A(n2660), .B(h0[30]), .Z(n6648) );
  COND2X1 U7281 ( .A(n6703), .B(n6579), .C(n2515), .D(n6648), .Z(n6617) );
  CFA1X1 U7282 ( .A(n6582), .B(n6581), .CI(n6580), .CO(n6637), .S(n6589) );
  CENX1 U7283 ( .A(n7134), .B(h0[20]), .Z(n6641) );
  COND2X1 U7284 ( .A(n7119), .B(n6583), .C(n7171), .D(n6641), .Z(n6616) );
  COND2X1 U7285 ( .A(n7065), .B(n6584), .C(n2477), .D(n6640), .Z(n6615) );
  CENX1 U7286 ( .A(h0[22]), .B(n6970), .Z(n6649) );
  COND2X1 U7287 ( .A(n7114), .B(n6649), .C(n6585), .D(n2294), .Z(n6614) );
  CEO3X2 U7288 ( .A(n6661), .B(n6658), .C(n6662), .Z(n6944) );
  CEO3X2 U7289 ( .A(n6588), .B(n6587), .C(n6586), .Z(n6899) );
  CENX2 U7290 ( .A(n6590), .B(n6589), .Z(n6592) );
  CENX2 U7291 ( .A(n6592), .B(n2357), .Z(n6901) );
  CIVX1 U7292 ( .A(n6597), .Z(n6594) );
  CIVX2 U7293 ( .A(n6598), .Z(n6593) );
  CND2X1 U7294 ( .A(n6594), .B(n6593), .Z(n6595) );
  CND2X1 U7295 ( .A(n6596), .B(n6595), .Z(n6600) );
  CND2X2 U7296 ( .A(n6600), .B(n6599), .Z(n6903) );
  CFA1X1 U7297 ( .A(n6603), .B(n6602), .CI(n6601), .CO(n6588), .S(n6902) );
  COR2X1 U7298 ( .A(n6903), .B(n6902), .Z(n6608) );
  CNR2X2 U7299 ( .A(n6607), .B(n6606), .Z(n6605) );
  CND2X2 U7300 ( .A(n6608), .B(n6904), .Z(n6610) );
  CND2X2 U7301 ( .A(n6610), .B(n6609), .Z(n6900) );
  COND1X2 U7302 ( .A(n6899), .B(n6901), .C(n6900), .Z(n6612) );
  CND2X2 U7303 ( .A(n6612), .B(n6611), .Z(n6943) );
  CNR2X2 U7304 ( .A(n6944), .B(n6943), .Z(n6613) );
  CIVX2 U7305 ( .A(n6613), .Z(n7439) );
  CFA1X1 U7306 ( .A(n6616), .B(n6615), .CI(n6614), .CO(n6673), .S(n6636) );
  CFA1X1 U7307 ( .A(n6619), .B(n6618), .CI(n6617), .CO(n6672), .S(n6638) );
  CENX2 U7308 ( .A(n6673), .B(n6621), .Z(n6690) );
  CND2X2 U7309 ( .A(n6626), .B(n6625), .Z(n6688) );
  CFA1X1 U7310 ( .A(n6629), .B(n6628), .CI(n6627), .CO(n6689), .S(n6651) );
  CENX2 U7311 ( .A(n6688), .B(n6689), .Z(n6630) );
  CIVX2 U7312 ( .A(n6712), .Z(n6714) );
  CND2X1 U7313 ( .A(n6635), .B(n6634), .Z(n6711) );
  CFA1X1 U7314 ( .A(n6638), .B(n6637), .CI(n6636), .CO(n6683), .S(n6631) );
  CENX1 U7315 ( .A(n7134), .B(n2280), .Z(n6669) );
  CENX1 U7316 ( .A(h0[19]), .B(n7202), .Z(n6708) );
  CENX1 U7317 ( .A(n6680), .B(n6643), .Z(n6695) );
  CENX1 U7318 ( .A(n6699), .B(h0[29]), .Z(n6700) );
  CENX1 U7319 ( .A(n7173), .B(h0[15]), .Z(n6707) );
  COND2X1 U7320 ( .A(n7228), .B(n6645), .C(n6707), .D(n7301), .Z(n6722) );
  CIVX2 U7321 ( .A(n6722), .Z(n6697) );
  CENX1 U7322 ( .A(n6769), .B(h0[27]), .Z(n6668) );
  COND2X1 U7323 ( .A(n2420), .B(n6646), .C(n6770), .D(n6668), .Z(n6696) );
  CENX1 U7324 ( .A(h0[23]), .B(n6970), .Z(n6670) );
  CENX1 U7325 ( .A(n6103), .B(h0[17]), .Z(n6709) );
  COND2X1 U7326 ( .A(n2282), .B(n6650), .C(n2433), .D(n6709), .Z(n6677) );
  CENX2 U7327 ( .A(n6683), .B(n6684), .Z(n6656) );
  COND1X1 U7328 ( .A(n6652), .B(n6653), .C(n6651), .Z(n6655) );
  CND2X2 U7329 ( .A(n6655), .B(n6654), .Z(n6685) );
  CENX2 U7330 ( .A(n6685), .B(n6656), .Z(n6713) );
  CEN3X2 U7331 ( .A(n6714), .B(n6711), .C(n6713), .Z(n6946) );
  CIVX2 U7332 ( .A(n6946), .Z(n6667) );
  CIVX2 U7333 ( .A(n6662), .Z(n6657) );
  CND2IX2 U7334 ( .B(n2445), .A(n6657), .Z(n6660) );
  CND2X2 U7335 ( .A(n6660), .B(n6659), .Z(n6665) );
  CIVX1 U7336 ( .A(n2445), .Z(n6663) );
  CND2X2 U7337 ( .A(n6665), .B(n6664), .Z(n6945) );
  CIVX2 U7338 ( .A(n6945), .Z(n6666) );
  CND2X4 U7339 ( .A(n6667), .B(n6666), .Z(n7443) );
  CENX1 U7340 ( .A(n6769), .B(h0[28]), .Z(n6729) );
  COND2X1 U7341 ( .A(n2420), .B(n6668), .C(n6770), .D(n6729), .Z(n6751) );
  COND2X1 U7342 ( .A(n7119), .B(n6669), .C(n7171), .D(n6718), .Z(n6749) );
  CENX1 U7343 ( .A(h0[24]), .B(n6970), .Z(n6731) );
  COND2X1 U7344 ( .A(n7114), .B(n6731), .C(n6670), .D(n7095), .Z(n6750) );
  CEO3X1 U7345 ( .A(n6751), .B(n6749), .C(n6750), .Z(n6738) );
  COND1X1 U7346 ( .A(n6672), .B(n6673), .C(n6671), .Z(n6675) );
  CND2X1 U7347 ( .A(n6673), .B(n6672), .Z(n6674) );
  CND2X2 U7348 ( .A(n6675), .B(n6674), .Z(n6737) );
  COND2X1 U7349 ( .A(n7065), .B(n6676), .C(n2477), .D(n6746), .Z(n6725) );
  CND2X2 U7350 ( .A(n6682), .B(n6681), .Z(n6726) );
  CEO3X2 U7351 ( .A(n6725), .B(n6724), .C(n6726), .Z(n6739) );
  CEO3X1 U7352 ( .A(n6738), .B(n6737), .C(n6739), .Z(n6761) );
  CND2X2 U7353 ( .A(n6687), .B(n6686), .Z(n6759) );
  COND1X2 U7354 ( .A(n6689), .B(n6690), .C(n6688), .Z(n6692) );
  CND2X2 U7355 ( .A(n6692), .B(n6691), .Z(n6734) );
  CFA1X1 U7356 ( .A(n6695), .B(n6694), .CI(n6693), .CO(n6733), .S(n6684) );
  CFA1X1 U7357 ( .A(n6698), .B(n6697), .CI(n6696), .CO(n6744), .S(n6694) );
  CENX1 U7358 ( .A(n6699), .B(h0[30]), .Z(n6730) );
  COND2X1 U7359 ( .A(n6701), .B(n6700), .C(n6765), .D(n6730), .Z(n6721) );
  CIVXL U7360 ( .A(n6703), .Z(n6706) );
  CIVX2 U7361 ( .A(n6704), .Z(n6705) );
  COND1X1 U7362 ( .A(n5712), .B(n6706), .C(n6705), .Z(n6720) );
  CENX1 U7363 ( .A(n7173), .B(h0[16]), .Z(n6717) );
  COND2X1 U7364 ( .A(n7228), .B(n6707), .C(n6717), .D(n2382), .Z(n6756) );
  CENX1 U7365 ( .A(h0[20]), .B(n7202), .Z(n6745) );
  COND2X1 U7366 ( .A(n7205), .B(n6708), .C(n7203), .D(n6745), .Z(n6755) );
  CENXL U7367 ( .A(n7090), .B(h0[18]), .Z(n6747) );
  COND2X1 U7368 ( .A(n7126), .B(n6709), .C(n2433), .D(n6747), .Z(n6754) );
  CENX2 U7369 ( .A(n6733), .B(n6732), .Z(n6710) );
  CENX2 U7370 ( .A(n6734), .B(n6710), .Z(n6760) );
  CEO3X2 U7371 ( .A(n6761), .B(n6759), .C(n6760), .Z(n6948) );
  CND2IX1 U7372 ( .B(n6714), .A(n6713), .Z(n6715) );
  CND2X2 U7373 ( .A(n6716), .B(n6715), .Z(n6947) );
  CNR2X2 U7374 ( .A(n6948), .B(n6947), .Z(n7325) );
  CENX1 U7375 ( .A(n7173), .B(h0[17]), .Z(n6800) );
  COND2X1 U7376 ( .A(n7228), .B(n6717), .C(n6800), .D(n2382), .Z(n6846) );
  CIVX2 U7377 ( .A(n6846), .Z(n6776) );
  CNIVXL U7378 ( .A(n6969), .Z(n6719) );
  COND2X1 U7379 ( .A(n6307), .B(n6718), .C(n7171), .D(n6773), .Z(n6778) );
  CENX1 U7380 ( .A(n6776), .B(n6778), .Z(n6723) );
  CND2X2 U7381 ( .A(n6728), .B(n6727), .Z(n6810) );
  CENX1 U7382 ( .A(n6769), .B(h0[29]), .Z(n6771) );
  COND2X1 U7383 ( .A(n2420), .B(n6729), .C(n6770), .D(n6771), .Z(n6804) );
  CENX1 U7384 ( .A(n6699), .B(h0[31]), .Z(n6764) );
  COND2X1 U7385 ( .A(n6765), .B(n6764), .C(n6730), .D(n1582), .Z(n6802) );
  CENX1 U7386 ( .A(h0[25]), .B(n2659), .Z(n6772) );
  CEO3X1 U7387 ( .A(n6804), .B(n6802), .C(n6803), .Z(n6812) );
  CND2X2 U7388 ( .A(n6736), .B(n6735), .Z(n6816) );
  COND1X2 U7389 ( .A(n6738), .B(n6739), .C(n6737), .Z(n6741) );
  CND2X2 U7390 ( .A(n6739), .B(n6738), .Z(n6740) );
  CND2X2 U7391 ( .A(n6741), .B(n6740), .Z(n6782) );
  CFA1X1 U7392 ( .A(n6744), .B(n6743), .CI(n6742), .CO(n6783), .S(n6732) );
  CENX1 U7393 ( .A(n2280), .B(n7202), .Z(n6775) );
  COND2X1 U7394 ( .A(n7205), .B(n6745), .C(n7203), .D(n6775), .Z(n6809) );
  COND2X1 U7395 ( .A(n6974), .B(n6746), .C(n6972), .D(n6793), .Z(n6808) );
  COND2X1 U7396 ( .A(n6747), .B(n7126), .C(n7124), .D(n6795), .Z(n6807) );
  CIVXL U7397 ( .A(n6751), .Z(n6748) );
  CND2IX1 U7398 ( .B(n6748), .A(n6750), .Z(n6753) );
  COND1X1 U7399 ( .A(n6751), .B(n6750), .C(n6749), .Z(n6752) );
  CND2X2 U7400 ( .A(n6753), .B(n6752), .Z(n6788) );
  CFA1X1 U7401 ( .A(n6756), .B(n6755), .CI(n6754), .CO(n6789), .S(n6742) );
  CENX2 U7402 ( .A(n6788), .B(n6789), .Z(n6757) );
  CENX2 U7403 ( .A(n2300), .B(n6757), .Z(n6784) );
  CENX2 U7404 ( .A(n6782), .B(n6758), .Z(n6817) );
  CEO3X1 U7405 ( .A(n6815), .B(n6816), .C(n6817), .Z(n6950) );
  CND2X2 U7406 ( .A(n6763), .B(n6762), .Z(n6949) );
  CNR2X2 U7407 ( .A(n6950), .B(n6949), .Z(n7332) );
  CNR2X2 U7408 ( .A(n7325), .B(n7332), .Z(n7417) );
  CIVX2 U7409 ( .A(n6764), .Z(n6768) );
  CND2IX1 U7410 ( .B(n2435), .A(n1582), .Z(n6767) );
  CENX1 U7411 ( .A(n6769), .B(h0[30]), .Z(n6830) );
  COND2X1 U7412 ( .A(n2420), .B(n6771), .C(n6770), .D(n6830), .Z(n6844) );
  CENX1 U7413 ( .A(h0[26]), .B(n6970), .Z(n6821) );
  COND2X1 U7414 ( .A(n7114), .B(n6821), .C(n6772), .D(n2295), .Z(n6820) );
  COND2X1 U7415 ( .A(n6468), .B(n6773), .C(n7171), .D(n6827), .Z(n6819) );
  CENX1 U7416 ( .A(h0[22]), .B(n7202), .Z(n6823) );
  COND2X1 U7417 ( .A(n7205), .B(n6775), .C(n7203), .D(n6823), .Z(n6818) );
  CND2X2 U7418 ( .A(n6780), .B(n6779), .Z(n6840) );
  CNIVX1 U7419 ( .A(n6840), .Z(n6781) );
  CIVX2 U7420 ( .A(n6782), .Z(n6786) );
  COND1X2 U7421 ( .A(n6787), .B(n6786), .C(n6785), .Z(n6855) );
  CENX1 U7422 ( .A(n5932), .B(h0[28]), .Z(n6824) );
  COND2X1 U7423 ( .A(n6974), .B(n6793), .C(n6972), .D(n6824), .Z(n6849) );
  CIVX2 U7424 ( .A(n7126), .Z(n6794) );
  CND2IX1 U7425 ( .B(n6795), .A(n6794), .Z(n6799) );
  CENX1 U7426 ( .A(n6103), .B(h0[20]), .Z(n6822) );
  CIVX2 U7427 ( .A(n6822), .Z(n6796) );
  CND2X2 U7428 ( .A(n6797), .B(n6796), .Z(n6798) );
  CND2X2 U7429 ( .A(n6799), .B(n6798), .Z(n6847) );
  CENX1 U7430 ( .A(n7173), .B(h0[18]), .Z(n6843) );
  COND2X1 U7431 ( .A(n7228), .B(n6800), .C(n6843), .D(n7301), .Z(n6848) );
  CENX1 U7432 ( .A(n6847), .B(n6848), .Z(n6801) );
  COND1X1 U7433 ( .A(n6804), .B(n6803), .C(n6802), .Z(n6805) );
  CND2X2 U7434 ( .A(n6806), .B(n6805), .Z(n6853) );
  CFA1X1 U7435 ( .A(n6809), .B(n6808), .CI(n6807), .CO(n6852), .S(n6790) );
  COND1X2 U7436 ( .A(n6812), .B(n6811), .C(n6810), .Z(n6814) );
  CND2X2 U7437 ( .A(n6814), .B(n6813), .Z(n6834) );
  CEO3X2 U7438 ( .A(n6832), .B(n6833), .C(n6834), .Z(n6857) );
  CNR2X2 U7439 ( .A(n6952), .B(n6951), .Z(n7420) );
  CFA1X1 U7440 ( .A(n6820), .B(n6819), .CI(n6818), .CO(n6883), .S(n6838) );
  COND2X2 U7441 ( .A(n7114), .B(n6866), .C(n6821), .D(n2295), .Z(n6864) );
  CENXL U7442 ( .A(n7090), .B(n2278), .Z(n6867) );
  COND2X1 U7443 ( .A(n2282), .B(n6822), .C(n6867), .D(n2433), .Z(n6863) );
  CENX1 U7444 ( .A(h0[23]), .B(n7202), .Z(n6891) );
  CENX1 U7445 ( .A(n5932), .B(h0[29]), .Z(n6868) );
  CENX1 U7446 ( .A(n7134), .B(h0[25]), .Z(n6887) );
  CIVX2 U7447 ( .A(n6887), .Z(n6825) );
  CENXL U7448 ( .A(h0[31]), .B(n6828), .Z(n6869) );
  COND2X1 U7449 ( .A(n6831), .B(n6830), .C(n6829), .D(n6869), .Z(n6888) );
  CNIVX4 U7450 ( .A(n6832), .Z(n6835) );
  COND1X2 U7451 ( .A(n6834), .B(n6835), .C(n6833), .Z(n6837) );
  CND2X2 U7452 ( .A(n6835), .B(n6834), .Z(n6836) );
  CND2X2 U7453 ( .A(n6837), .B(n6836), .Z(n6892) );
  COND1X2 U7454 ( .A(n6839), .B(n6840), .C(n6838), .Z(n6842) );
  CND2X1 U7455 ( .A(n6840), .B(n6839), .Z(n6841) );
  CND2X2 U7456 ( .A(n6842), .B(n6841), .Z(n6873) );
  CENX1 U7457 ( .A(n7173), .B(h0[19]), .Z(n6865) );
  COND2X1 U7458 ( .A(n7228), .B(n6843), .C(n6865), .D(n7301), .Z(n6967) );
  CIVX2 U7459 ( .A(n6967), .Z(n6878) );
  CFA1X1 U7460 ( .A(n6846), .B(n6845), .CI(n6844), .CO(n6877), .S(n6839) );
  COND1XL U7461 ( .A(n6848), .B(n6849), .C(n6847), .Z(n6851) );
  CND2X1 U7462 ( .A(n6849), .B(n6848), .Z(n6850) );
  CND2X1 U7463 ( .A(n6851), .B(n6850), .Z(n6879) );
  CEO3X2 U7464 ( .A(n6878), .B(n6877), .C(n6879), .Z(n6872) );
  CENX2 U7465 ( .A(n6872), .B(n6874), .Z(n6854) );
  CENX2 U7466 ( .A(n6873), .B(n6854), .Z(n6894) );
  CIVX2 U7467 ( .A(n6954), .Z(n6861) );
  COND1X2 U7468 ( .A(n6856), .B(n6857), .C(n6855), .Z(n6859) );
  CND2X2 U7469 ( .A(n6859), .B(n6858), .Z(n6953) );
  CIVX2 U7470 ( .A(n6953), .Z(n6860) );
  CND2X2 U7471 ( .A(n6861), .B(n6860), .Z(n7391) );
  CFA1X1 U7472 ( .A(n6864), .B(n6863), .CI(n6862), .CO(n6983), .S(n6884) );
  CENX1 U7473 ( .A(n7173), .B(h0[20]), .Z(n6977) );
  CENX1 U7474 ( .A(h0[28]), .B(n6970), .Z(n6971) );
  COND2X1 U7475 ( .A(n7114), .B(n6971), .C(n6866), .D(n2294), .Z(n6975) );
  CENXL U7476 ( .A(n7090), .B(h0[22]), .Z(n6980) );
  COND2X1 U7477 ( .A(n6974), .B(n6868), .C(n6972), .D(n6973), .Z(n6966) );
  COND1X2 U7478 ( .A(n6874), .B(n6873), .C(n6872), .Z(n6876) );
  CND2X1 U7479 ( .A(n6874), .B(n6873), .Z(n6875) );
  CND2X2 U7480 ( .A(n6876), .B(n6875), .Z(n6992) );
  CND2X1 U7481 ( .A(n6879), .B(n6878), .Z(n6880) );
  COND2X1 U7482 ( .A(n6774), .B(n6887), .C(n7171), .D(n6968), .Z(n6989) );
  CENX1 U7483 ( .A(h0[24]), .B(n7202), .Z(n6979) );
  COND2X1 U7484 ( .A(n7123), .B(n6891), .C(n7203), .D(n6979), .Z(n6987) );
  CEO3X2 U7485 ( .A(n6994), .B(n6992), .C(n6991), .Z(n6956) );
  CIVX2 U7486 ( .A(n6956), .Z(n6898) );
  CND2X2 U7487 ( .A(n6896), .B(n6895), .Z(n6955) );
  CIVX2 U7488 ( .A(n6955), .Z(n6897) );
  CND2X2 U7489 ( .A(n6898), .B(n6897), .Z(n7395) );
  CNR2X2 U7490 ( .A(n7420), .B(n6959), .Z(n6961) );
  CND2X2 U7491 ( .A(n7417), .B(n6961), .Z(n7051) );
  CNR2X4 U7492 ( .A(n7337), .B(n7051), .Z(n7151) );
  CEO3X2 U7493 ( .A(n6901), .B(n6900), .C(n6899), .Z(n6937) );
  CIVX2 U7494 ( .A(n6937), .Z(n6938) );
  CENX2 U7495 ( .A(n6906), .B(n6905), .Z(n6907) );
  CENX2 U7496 ( .A(n1265), .B(n6907), .Z(n6918) );
  COND1X2 U7497 ( .A(n6910), .B(n6911), .C(n6909), .Z(n6913) );
  CND2X2 U7498 ( .A(n6911), .B(n6910), .Z(n6912) );
  CND2X2 U7499 ( .A(n6913), .B(n6912), .Z(n6917) );
  COND1X1 U7500 ( .A(n6916), .B(n6918), .C(n6917), .Z(n6915) );
  CND2X1 U7501 ( .A(n6916), .B(n6918), .Z(n6914) );
  CND2X2 U7502 ( .A(n6915), .B(n6914), .Z(n6936) );
  CIVX2 U7503 ( .A(n6936), .Z(n6939) );
  CND2X2 U7504 ( .A(n6938), .B(n6939), .Z(n7323) );
  CEO3X1 U7505 ( .A(n6918), .B(n6917), .C(n6916), .Z(n6935) );
  CIVX2 U7506 ( .A(n6935), .Z(n6925) );
  COND1X1 U7507 ( .A(n6919), .B(n6921), .C(n6920), .Z(n6923) );
  CND2X2 U7508 ( .A(n6923), .B(n6922), .Z(n6934) );
  CIVX2 U7509 ( .A(n6934), .Z(n6924) );
  CND2X2 U7510 ( .A(n6925), .B(n6924), .Z(n7322) );
  CND2X1 U7511 ( .A(n7323), .B(n7322), .Z(n7327) );
  CIVX2 U7512 ( .A(n7327), .Z(n6926) );
  CND3X4 U7513 ( .A(n7373), .B(n7151), .C(n6926), .Z(n7281) );
  CANR1X2 U7514 ( .A(n2525), .B(n2386), .C(n2481), .Z(n7485) );
  CND2X1 U7515 ( .A(n7323), .B(n7322), .Z(n6942) );
  CIVX2 U7516 ( .A(n7454), .Z(n6933) );
  CND2X2 U7517 ( .A(n6931), .B(n6930), .Z(n7456) );
  CIVX2 U7518 ( .A(n7456), .Z(n6932) );
  CND2X1 U7519 ( .A(n6935), .B(n6934), .Z(n7374) );
  CND2X2 U7520 ( .A(n6937), .B(n6936), .Z(n7378) );
  CND2X1 U7521 ( .A(n6939), .B(n6938), .Z(n6940) );
  CND2X2 U7522 ( .A(n6944), .B(n6943), .Z(n7370) );
  CIVX2 U7523 ( .A(n7370), .Z(n7437) );
  CND2X2 U7524 ( .A(n6946), .B(n6945), .Z(n7442) );
  CIVX2 U7525 ( .A(n7442), .Z(n7328) );
  CANR1X2 U7526 ( .A(n7437), .B(n7443), .C(n7328), .Z(n6963) );
  CND2X2 U7527 ( .A(n6948), .B(n6947), .Z(n7364) );
  CND2X1 U7528 ( .A(n6950), .B(n6949), .Z(n7333) );
  COND1X2 U7529 ( .A(n7364), .B(n7332), .C(n7333), .Z(n7415) );
  CND2X2 U7530 ( .A(n6954), .B(n6953), .Z(n7349) );
  CIVX2 U7531 ( .A(n7349), .Z(n7389) );
  CND2X2 U7532 ( .A(n6956), .B(n6955), .Z(n7394) );
  CIVX2 U7533 ( .A(n7394), .Z(n6957) );
  CANR1X2 U7534 ( .A(n7395), .B(n7389), .C(n6957), .Z(n6958) );
  COND1X1 U7535 ( .A(n7340), .B(n6959), .C(n6958), .Z(n6960) );
  CIVXL U7536 ( .A(n7314), .Z(n6964) );
  COND1XL U7537 ( .A(n7281), .B(n2359), .C(n6964), .Z(n7002) );
  CFA1X1 U7538 ( .A(n6967), .B(n6966), .CI(n6965), .CO(n7069), .S(n6984) );
  CENX1 U7539 ( .A(h0[29]), .B(n6970), .Z(n7066) );
  COND2X1 U7540 ( .A(n6974), .B(n6973), .C(n6972), .D(n7064), .Z(n7059) );
  CENX1 U7541 ( .A(n7173), .B(n2279), .Z(n7060) );
  CIVX1 U7542 ( .A(n7060), .Z(n6976) );
  CIVX1 U7543 ( .A(n6977), .Z(n6978) );
  CENX1 U7544 ( .A(h0[25]), .B(n7202), .Z(n7063) );
  COND2X1 U7545 ( .A(n7123), .B(n6979), .C(n7203), .D(n7063), .Z(n7055) );
  CIVX2 U7546 ( .A(n7055), .Z(n6981) );
  CENX1 U7547 ( .A(n6103), .B(h0[23]), .Z(n7061) );
  COND2X1 U7548 ( .A(n7252), .B(n6980), .C(n7253), .D(n7061), .Z(n7054) );
  CEO3X2 U7549 ( .A(n7081), .B(n6981), .C(n7054), .Z(n7073) );
  CFA1X1 U7550 ( .A(n6989), .B(n6988), .CI(n6987), .CO(n7071), .S(n6990) );
  CNIVX4 U7551 ( .A(n6991), .Z(n6995) );
  COND1X2 U7552 ( .A(n6994), .B(n6995), .C(n6993), .Z(n6997) );
  CND2X2 U7553 ( .A(n6995), .B(n6994), .Z(n6996) );
  CND2X2 U7554 ( .A(n6997), .B(n6996), .Z(n6999) );
  CNR2X1 U7555 ( .A(n7000), .B(n6999), .Z(n6998) );
  CIVX2 U7556 ( .A(n6998), .Z(n7354) );
  CND2X1 U7557 ( .A(n7000), .B(n6999), .Z(n7152) );
  CND2X1 U7558 ( .A(n7354), .B(n7152), .Z(n7001) );
  CENXL U7559 ( .A(n7002), .B(n7001), .Z(N66) );
  CIVXL U7560 ( .A(n7003), .Z(n7023) );
  CND2XL U7561 ( .A(n7023), .B(n7021), .Z(n7007) );
  CIVXL U7562 ( .A(n2368), .Z(n7042) );
  CIVXL U7563 ( .A(n7042), .Z(n7005) );
  COND1XL U7564 ( .A(n7020), .B(n7475), .C(n7005), .Z(n7006) );
  CENXL U7565 ( .A(n7007), .B(n7006), .Z(N51) );
  COND1XL U7566 ( .A(n7013), .B(n7494), .C(n2297), .Z(n7017) );
  CND2X1 U7567 ( .A(n7015), .B(n7014), .Z(n7016) );
  CENXL U7568 ( .A(n7016), .B(n7017), .Z(N40) );
  CND2XL U7569 ( .A(n2558), .B(n7019), .Z(n7027) );
  CIVXL U7570 ( .A(n7020), .Z(n7037) );
  CND2XL U7571 ( .A(n7037), .B(n7023), .Z(n7025) );
  CIVXL U7572 ( .A(n7021), .Z(n7022) );
  CANR1XL U7573 ( .A(n7023), .B(n7042), .C(n7022), .Z(n7024) );
  COND1XL U7574 ( .A(n7475), .B(n7025), .C(n7024), .Z(n7026) );
  CENXL U7575 ( .A(n7027), .B(n7026), .Z(N52) );
  CNIVXL U7576 ( .A(n7028), .Z(n7040) );
  CIVXL U7577 ( .A(n7040), .Z(n7029) );
  CND2IX1 U7578 ( .B(n7030), .A(n7029), .Z(n7034) );
  CND2XL U7579 ( .A(n7037), .B(n2615), .Z(n7032) );
  CANR1XL U7580 ( .A(n2615), .B(n7042), .C(n2557), .Z(n7031) );
  COND1XL U7581 ( .A(n7475), .B(n7032), .C(n7031), .Z(n7033) );
  CENXL U7582 ( .A(n7034), .B(n7033), .Z(N53) );
  CIVXL U7583 ( .A(n7035), .Z(n7036) );
  CNR2XL U7584 ( .A(n7036), .B(n7040), .Z(n7043) );
  CND2XL U7585 ( .A(n7043), .B(n7037), .Z(n7045) );
  COND1XL U7586 ( .A(n7040), .B(n2607), .C(n7039), .Z(n7041) );
  CANR1XL U7587 ( .A(n7043), .B(n7042), .C(n7041), .Z(n7044) );
  CIVXL U7588 ( .A(n1261), .Z(n7048) );
  CND2XL U7589 ( .A(n7048), .B(n7047), .Z(n7049) );
  CENXL U7590 ( .A(n7050), .B(n7049), .Z(N54) );
  CNR2X2 U7591 ( .A(n7052), .B(n7337), .Z(n7132) );
  CIVX1 U7592 ( .A(n7054), .Z(n7058) );
  CNR2IX2 U7593 ( .B(n7081), .A(n7055), .Z(n7057) );
  CND2IX1 U7594 ( .B(n7081), .A(n7055), .Z(n7056) );
  COND1X1 U7595 ( .A(n7058), .B(n7057), .C(n7056), .Z(n7087) );
  CNIVX1 U7596 ( .A(n7228), .Z(n7300) );
  CENX1 U7597 ( .A(n7173), .B(h0[22]), .Z(n7082) );
  COND2X1 U7598 ( .A(n7300), .B(n7060), .C(n7082), .D(n2382), .Z(n7085) );
  CENXL U7599 ( .A(n6103), .B(h0[24]), .Z(n7091) );
  COND2X1 U7600 ( .A(n7252), .B(n7061), .C(n7253), .D(n7091), .Z(n7084) );
  CENX1 U7601 ( .A(h0[26]), .B(n7062), .Z(n7089) );
  COND2X1 U7602 ( .A(n7123), .B(n7063), .C(n7203), .D(n7089), .Z(n7083) );
  CENX1 U7603 ( .A(h0[30]), .B(n2659), .Z(n7094) );
  COND2X1 U7604 ( .A(n7114), .B(n7094), .C(n7066), .D(n7095), .Z(n7079) );
  CNR2X1 U7605 ( .A(n7154), .B(n7153), .Z(n7077) );
  CIVX2 U7606 ( .A(n7077), .Z(n7358) );
  CND2X2 U7607 ( .A(n7354), .B(n7358), .Z(n7425) );
  CFA1X1 U7608 ( .A(n7079), .B(n7080), .CI(n7081), .CO(n7108), .S(n7096) );
  CENX1 U7609 ( .A(n7173), .B(h0[23]), .Z(n7121) );
  COND2X2 U7610 ( .A(n7228), .B(n7082), .C(n2382), .D(n7121), .Z(n7145) );
  CIVX2 U7611 ( .A(n7145), .Z(n7107) );
  CFA1X1 U7612 ( .A(n7085), .B(n7084), .CI(n7083), .CO(n7112), .S(n7097) );
  CFA1X1 U7613 ( .A(n7088), .B(n7087), .CI(n7086), .CO(n7111), .S(n7103) );
  CENX1 U7614 ( .A(h0[27]), .B(n7202), .Z(n7122) );
  COND2X1 U7615 ( .A(n7123), .B(n7089), .C(n7203), .D(n7122), .Z(n7129) );
  CENXL U7616 ( .A(n6103), .B(h0[25]), .Z(n7125) );
  COND2X1 U7617 ( .A(n7252), .B(n7091), .C(n7253), .D(n7125), .Z(n7128) );
  CENX1 U7618 ( .A(h0[31]), .B(n7092), .Z(n7115) );
  COR2X1 U7619 ( .A(n7114), .B(n7115), .Z(n7093) );
  COND1X2 U7620 ( .A(n7095), .B(n7094), .C(n7093), .Z(n7127) );
  CND2X2 U7621 ( .A(n7100), .B(n7099), .Z(n7104) );
  CFA1X1 U7622 ( .A(n7103), .B(n7102), .CI(n7101), .CO(n7156), .S(n7154) );
  CNR2X2 U7623 ( .A(n7157), .B(n7156), .Z(n7432) );
  CNR2X2 U7624 ( .A(n7425), .B(n7432), .Z(n7260) );
  CFA1X1 U7625 ( .A(n7106), .B(n7105), .CI(n7104), .CO(n7162), .S(n7157) );
  CFA1X1 U7626 ( .A(n7109), .B(n7108), .CI(n7107), .CO(n7160), .S(n7106) );
  CFA1X1 U7627 ( .A(n7112), .B(n7111), .CI(n7110), .CO(n7159), .S(n7105) );
  CND2X1 U7628 ( .A(n7114), .B(n2294), .Z(n7117) );
  CIVX1 U7629 ( .A(n7115), .Z(n7116) );
  CND2X2 U7630 ( .A(n7117), .B(n7116), .Z(n7146) );
  CENX2 U7631 ( .A(n7146), .B(n7145), .Z(n7120) );
  CENX2 U7632 ( .A(n7120), .B(n7144), .Z(n7139) );
  CENX1 U7633 ( .A(n7173), .B(h0[24]), .Z(n7140) );
  COND2X1 U7634 ( .A(n7228), .B(n7121), .C(n7140), .D(n2381), .Z(n7143) );
  CENX1 U7635 ( .A(h0[28]), .B(n7202), .Z(n7133) );
  COND2X1 U7636 ( .A(n7123), .B(n7122), .C(n7203), .D(n7133), .Z(n7142) );
  CENXL U7637 ( .A(n7090), .B(h0[26]), .Z(n7136) );
  COND2X1 U7638 ( .A(n2282), .B(n7125), .C(n2433), .D(n7136), .Z(n7141) );
  CFA1X1 U7639 ( .A(n7129), .B(n7128), .CI(n7127), .CO(n7137), .S(n7110) );
  CNIVX4 U7640 ( .A(n2376), .Z(n7385) );
  CFA1X1 U7641 ( .A(n7160), .B(n7159), .CI(n7158), .CO(n7166), .S(n7130) );
  CENX1 U7642 ( .A(h0[29]), .B(n7202), .Z(n7175) );
  COND2X1 U7643 ( .A(n7205), .B(n7133), .C(n7203), .D(n7175), .Z(n7178) );
  CENXL U7644 ( .A(n7134), .B(h0[31]), .Z(n7170) );
  COND2X1 U7645 ( .A(n6774), .B(n7135), .C(n7171), .D(n7170), .Z(n7177) );
  CENXL U7646 ( .A(n7090), .B(h0[27]), .Z(n7172) );
  COND2X1 U7647 ( .A(n7252), .B(n7136), .C(n7253), .D(n7172), .Z(n7176) );
  CFA1X1 U7648 ( .A(n7139), .B(n7138), .CI(n7137), .CO(n7184), .S(n7158) );
  COND2X1 U7649 ( .A(n7300), .B(n7140), .C(n7174), .D(n2381), .Z(n7196) );
  CIVX2 U7650 ( .A(n7196), .Z(n7182) );
  CFA1X1 U7651 ( .A(n7143), .B(n7142), .CI(n7141), .CO(n7181), .S(n7138) );
  CND2X2 U7652 ( .A(n7148), .B(n7147), .Z(n7180) );
  CIVX2 U7653 ( .A(n7191), .Z(n7450) );
  CIVX2 U7654 ( .A(n7152), .Z(n7353) );
  CND2X1 U7655 ( .A(n7154), .B(n7153), .Z(n7357) );
  CIVX2 U7656 ( .A(n7357), .Z(n7155) );
  CANR1X2 U7657 ( .A(n7353), .B(n7358), .C(n7155), .Z(n7427) );
  COND1XL U7658 ( .A(n7432), .B(n2352), .C(n7433), .Z(n7259) );
  CEO3XL U7659 ( .A(n7160), .B(n7159), .C(n7158), .Z(n7161) );
  CANR1XL U7660 ( .A(n7264), .B(n7259), .C(n7234), .Z(n7163) );
  COND1XL U7661 ( .A(n7164), .B(n7352), .C(n7163), .Z(n7446) );
  CIVX2 U7662 ( .A(n7449), .Z(n7167) );
  CANR1XL U7663 ( .A(n7450), .B(n7446), .C(n7167), .Z(n7168) );
  COND1XL U7664 ( .A(n7169), .B(n7485), .C(n7168), .Z(n7190) );
  CAOR1XL U7665 ( .A(n7171), .B(n6719), .C(n7170), .Z(n7195) );
  CENXL U7666 ( .A(n6103), .B(h0[28]), .Z(n7207) );
  CENX1 U7667 ( .A(n7173), .B(h0[26]), .Z(n7206) );
  COND2X1 U7668 ( .A(n7300), .B(n7174), .C(n7206), .D(n2382), .Z(n7198) );
  CENX1 U7669 ( .A(h0[30]), .B(n7202), .Z(n7204) );
  COND2X1 U7670 ( .A(n1226), .B(n7175), .C(n7203), .D(n7204), .Z(n7197) );
  CENX1 U7671 ( .A(n7198), .B(n7197), .Z(n7179) );
  CFA1X1 U7672 ( .A(n7178), .B(n7177), .CI(n7176), .CO(n7199), .S(n7185) );
  CENX1 U7673 ( .A(n7179), .B(n7199), .Z(n7209) );
  CFA1X1 U7674 ( .A(n7182), .B(n7181), .CI(n7180), .CO(n7208), .S(n7183) );
  CFA1X1 U7675 ( .A(n7185), .B(n7184), .CI(n7183), .CO(n7186), .S(n7165) );
  CIVX2 U7676 ( .A(n7233), .Z(n7188) );
  CND2X1 U7677 ( .A(n7187), .B(n7186), .Z(n7232) );
  CND2X1 U7678 ( .A(n7188), .B(n7232), .Z(n7189) );
  CENXL U7679 ( .A(n7190), .B(n7189), .Z(N71) );
  CIVX2 U7680 ( .A(n7235), .Z(n7193) );
  CND2X2 U7681 ( .A(n7193), .B(n7192), .Z(n7236) );
  CFA1X1 U7682 ( .A(n7196), .B(n7195), .CI(n7194), .CO(n7214), .S(n7210) );
  COND1XL U7683 ( .A(n7198), .B(n7199), .C(n7197), .Z(n7201) );
  CND2X1 U7684 ( .A(n7199), .B(n7198), .Z(n7200) );
  CND2X1 U7685 ( .A(n7201), .B(n7200), .Z(n7213) );
  CENX1 U7686 ( .A(h0[31]), .B(n7202), .Z(n7216) );
  COND2X1 U7687 ( .A(n1226), .B(n7204), .C(n7203), .D(n7216), .Z(n7222) );
  CENX1 U7688 ( .A(h0[27]), .B(n7279), .Z(n7215) );
  COND2X1 U7689 ( .A(n7300), .B(n7206), .C(n7215), .D(n2381), .Z(n7226) );
  CIVX1 U7690 ( .A(n7226), .Z(n7221) );
  CENXL U7691 ( .A(n6103), .B(h0[29]), .Z(n7219) );
  CFA1X1 U7692 ( .A(n7210), .B(n7209), .CI(n7208), .CO(n7237), .S(n7187) );
  CNR2X1 U7693 ( .A(n7238), .B(n7237), .Z(n7211) );
  CIVX2 U7694 ( .A(n7211), .Z(n7319) );
  CIVX2 U7695 ( .A(n7275), .Z(n7268) );
  CFA1X1 U7696 ( .A(n7214), .B(n7213), .CI(n7212), .CO(n7240), .S(n7238) );
  CENX1 U7697 ( .A(h0[28]), .B(n7279), .Z(n7227) );
  COND2X1 U7698 ( .A(n7228), .B(n7215), .C(n7227), .D(n2382), .Z(n7231) );
  CENXL U7699 ( .A(n6103), .B(h0[30]), .Z(n7223) );
  CFA1X1 U7700 ( .A(n7222), .B(n7221), .CI(n7220), .CO(n7229), .S(n7212) );
  CNR2X1 U7701 ( .A(n7240), .B(n7239), .Z(n7274) );
  CIVX1 U7702 ( .A(n7274), .Z(n7271) );
  CND2X1 U7703 ( .A(n7268), .B(n7271), .Z(n7243) );
  CNR2X2 U7704 ( .A(n7281), .B(n7243), .Z(n7398) );
  CENXL U7705 ( .A(n6103), .B(h0[31]), .Z(n7251) );
  CFA1X1 U7706 ( .A(n7226), .B(n7225), .CI(n7224), .CO(n7249), .S(n7230) );
  CENX1 U7707 ( .A(h0[29]), .B(n7279), .Z(n7254) );
  COND2X1 U7708 ( .A(n7228), .B(n7227), .C(n7254), .D(n2382), .Z(n7278) );
  CIVX1 U7709 ( .A(n7278), .Z(n7248) );
  CFA1X1 U7710 ( .A(n7231), .B(n7230), .CI(n7229), .CO(n7244), .S(n7239) );
  COR2X1 U7711 ( .A(n7245), .B(n7244), .Z(n7403) );
  CND2XL U7712 ( .A(n7398), .B(n7403), .Z(n7247) );
  CND2IX2 U7713 ( .B(n7211), .A(n7313), .Z(n7290) );
  CND2X1 U7714 ( .A(n7238), .B(n7237), .Z(n7318) );
  CND2X1 U7715 ( .A(n7240), .B(n7239), .Z(n7288) );
  CIVXL U7716 ( .A(n7288), .Z(n7241) );
  COND1XL U7717 ( .A(n7243), .B(n7352), .C(n7242), .Z(n7399) );
  CND2X1 U7718 ( .A(n7245), .B(n7244), .Z(n7402) );
  CIVX1 U7719 ( .A(n7402), .Z(n7284) );
  CANR1XL U7720 ( .A(n7403), .B(n7399), .C(n7284), .Z(n7246) );
  COND1XL U7721 ( .A(n7247), .B(n7485), .C(n7246), .Z(n7258) );
  CFA1X1 U7722 ( .A(n7250), .B(n7249), .CI(n7248), .CO(n7256), .S(n7245) );
  CENX1 U7723 ( .A(h0[30]), .B(n7279), .Z(n7280) );
  COND2X1 U7724 ( .A(n7300), .B(n7254), .C(n7280), .D(n2381), .Z(n7276) );
  COR2X1 U7725 ( .A(n7256), .B(n7255), .Z(n7285) );
  CND2X1 U7726 ( .A(n7256), .B(n7255), .Z(n7282) );
  CND2X1 U7727 ( .A(n7285), .B(n7282), .Z(n7257) );
  CENXL U7728 ( .A(n7258), .B(n7257), .Z(N75) );
  CIVX2 U7729 ( .A(n7281), .Z(n7426) );
  CND2XL U7730 ( .A(n7426), .B(n7260), .Z(n7262) );
  CANR1XL U7731 ( .A(n7260), .B(n7314), .C(n7259), .Z(n7261) );
  COND1XL U7732 ( .A(n7262), .B(n7362), .C(n7261), .Z(n7266) );
  CND2X1 U7733 ( .A(n7264), .B(n7263), .Z(n7265) );
  CENXL U7734 ( .A(n7266), .B(n7265), .Z(N69) );
  CND2XL U7735 ( .A(n7426), .B(n7268), .Z(n7270) );
  CANR1XL U7736 ( .A(n7268), .B(n7314), .C(n7267), .Z(n7269) );
  COND1XL U7737 ( .A(n7270), .B(n2467), .C(n7269), .Z(n7273) );
  CND2XL U7738 ( .A(n7271), .B(n7288), .Z(n7272) );
  CENXL U7739 ( .A(n7273), .B(n7272), .Z(N73) );
  CND2XL U7740 ( .A(n7403), .B(n7285), .Z(n7287) );
  COR2X1 U7741 ( .A(n7274), .B(n7287), .Z(n7291) );
  CFA1X1 U7742 ( .A(n7278), .B(n7277), .CI(n7276), .CO(n7293), .S(n7255) );
  CENX1 U7743 ( .A(h0[31]), .B(n7279), .Z(n7299) );
  COND2X1 U7744 ( .A(n7300), .B(n7280), .C(n7299), .D(n2381), .Z(n7302) );
  CIVX1 U7745 ( .A(n7302), .Z(n7292) );
  COR2X1 U7746 ( .A(n7293), .B(n7292), .Z(n7411) );
  CNR2X2 U7747 ( .A(n7281), .B(n7296), .Z(n7479) );
  CIVXL U7748 ( .A(n7479), .Z(n7298) );
  CIVXL U7749 ( .A(n7282), .Z(n7283) );
  CANR1XL U7750 ( .A(n7285), .B(n7284), .C(n7283), .Z(n7286) );
  COAN1XL U7751 ( .A(n7288), .B(n7287), .C(n7286), .Z(n7289) );
  CND2X1 U7752 ( .A(n7293), .B(n7292), .Z(n7410) );
  CIVXL U7753 ( .A(n7410), .Z(n7294) );
  COND1X1 U7754 ( .A(n7296), .B(n2541), .C(n7295), .Z(n7482) );
  CIVXL U7755 ( .A(n7482), .Z(n7297) );
  COND1XL U7756 ( .A(n7298), .B(n7362), .C(n7297), .Z(n7305) );
  CAOR1X1 U7757 ( .A(n2382), .B(n7300), .C(n7299), .Z(n7303) );
  COR2XL U7758 ( .A(n7303), .B(n7302), .Z(n7483) );
  CND2XL U7759 ( .A(n7303), .B(n7302), .Z(n7480) );
  CND2XL U7760 ( .A(n7483), .B(n7480), .Z(n7304) );
  CENXL U7761 ( .A(n7305), .B(n7304), .Z(N77) );
  CIVXL U7762 ( .A(n7306), .Z(n7308) );
  CND2XL U7763 ( .A(n7307), .B(n7308), .Z(n7312) );
  COND1XL U7764 ( .A(n2509), .B(n7475), .C(n7309), .Z(n7311) );
  CENXL U7765 ( .A(n7312), .B(n7311), .Z(N48) );
  CND2XL U7766 ( .A(n7426), .B(n7315), .Z(n7317) );
  CANR1XL U7767 ( .A(n7315), .B(n7314), .C(n2351), .Z(n7316) );
  COND1XL U7768 ( .A(n7317), .B(n7362), .C(n7316), .Z(n7321) );
  CND2XL U7769 ( .A(n7319), .B(n7318), .Z(n7320) );
  CENXL U7770 ( .A(n7321), .B(n7320), .Z(N72) );
  CND2X1 U7771 ( .A(n7323), .B(n2376), .Z(n7324) );
  CNR2X2 U7772 ( .A(n7324), .B(n7383), .Z(n7436) );
  CIVX2 U7773 ( .A(n7436), .Z(n7369) );
  CNR2X1 U7774 ( .A(n7369), .B(n7337), .Z(n7414) );
  CIVXL U7775 ( .A(n7325), .Z(n7365) );
  CND2XL U7776 ( .A(n7414), .B(n7365), .Z(n7331) );
  CIVX2 U7777 ( .A(n7438), .Z(n7368) );
  CANR1X2 U7778 ( .A(n7437), .B(n7443), .C(n7328), .Z(n7339) );
  COND1X1 U7779 ( .A(n7337), .B(n7368), .C(n7339), .Z(n7416) );
  CIVXL U7780 ( .A(n7364), .Z(n7329) );
  CANR1XL U7781 ( .A(n7365), .B(n7416), .C(n7329), .Z(n7330) );
  COND1XL U7782 ( .A(n7331), .B(n2467), .C(n7330), .Z(n7336) );
  CIVXL U7783 ( .A(n7332), .Z(n7334) );
  CND2XL U7784 ( .A(n7334), .B(n7333), .Z(n7335) );
  CENXL U7785 ( .A(n7336), .B(n7335), .Z(N62) );
  CIVXL U7786 ( .A(n7337), .Z(n7338) );
  CND2X1 U7787 ( .A(n7344), .B(n7338), .Z(n7346) );
  CNR2X1 U7788 ( .A(n7369), .B(n7346), .Z(n7388) );
  CIVXL U7789 ( .A(n7388), .Z(n7348) );
  CIVX1 U7790 ( .A(n7339), .Z(n7343) );
  CND2IXL U7791 ( .B(n7420), .A(n7415), .Z(n7341) );
  CND2X1 U7792 ( .A(n7341), .B(n7421), .Z(n7342) );
  COND1X1 U7793 ( .A(n7346), .B(n7368), .C(n7345), .Z(n7390) );
  CIVXL U7794 ( .A(n7390), .Z(n7347) );
  COND1XL U7795 ( .A(n7348), .B(n7362), .C(n7347), .Z(n7351) );
  CND2X1 U7796 ( .A(n7349), .B(n7391), .Z(n7350) );
  CENXL U7797 ( .A(n7351), .B(n7350), .Z(N64) );
  CND2XL U7798 ( .A(n7426), .B(n7354), .Z(n7356) );
  CANR1XL U7799 ( .A(n7354), .B(n7314), .C(n7353), .Z(n7355) );
  COND1XL U7800 ( .A(n7356), .B(n2467), .C(n7355), .Z(n7360) );
  CND2X1 U7801 ( .A(n7358), .B(n7357), .Z(n7359) );
  CENXL U7802 ( .A(n7360), .B(n7359), .Z(N67) );
  CIVXL U7803 ( .A(n7414), .Z(n7363) );
  CIVXL U7804 ( .A(n7416), .Z(n7361) );
  COND1XL U7805 ( .A(n7363), .B(n2467), .C(n7361), .Z(n7367) );
  CND2X1 U7806 ( .A(n7365), .B(n7364), .Z(n7366) );
  CENXL U7807 ( .A(n7367), .B(n7366), .Z(N61) );
  COND1XL U7808 ( .A(n7369), .B(n7485), .C(n7368), .Z(n7372) );
  CND2X1 U7809 ( .A(n7439), .B(n7370), .Z(n7371) );
  CENXL U7810 ( .A(n7372), .B(n7371), .Z(N59) );
  CND2XL U7811 ( .A(n7373), .B(n7385), .Z(n7377) );
  CIVXL U7812 ( .A(n2391), .Z(n7375) );
  COND1XL U7813 ( .A(n7377), .B(n2359), .C(n7376), .Z(n7381) );
  CND2X1 U7814 ( .A(n7379), .B(n7378), .Z(n7380) );
  CENXL U7815 ( .A(n7381), .B(n7380), .Z(N58) );
  COND1XL U7816 ( .A(n7383), .B(n7485), .C(n2581), .Z(n7387) );
  CND2X1 U7817 ( .A(n7385), .B(n7384), .Z(n7386) );
  CENXL U7818 ( .A(n7387), .B(n7386), .Z(N57) );
  CND2XL U7819 ( .A(n7388), .B(n7391), .Z(n7393) );
  CANR1XL U7820 ( .A(n7391), .B(n7390), .C(n7389), .Z(n7392) );
  COND1XL U7821 ( .A(n7393), .B(n2623), .C(n7392), .Z(n7397) );
  CND2X1 U7822 ( .A(n7395), .B(n7394), .Z(n7396) );
  CENXL U7823 ( .A(n7397), .B(n7396), .Z(N65) );
  CIVXL U7824 ( .A(n7398), .Z(n7401) );
  CIVXL U7825 ( .A(n7399), .Z(n7400) );
  COND1XL U7826 ( .A(n7401), .B(n7485), .C(n7400), .Z(n7405) );
  CND2XL U7827 ( .A(n7403), .B(n7402), .Z(n7404) );
  CENXL U7828 ( .A(n7405), .B(n7404), .Z(N74) );
  CND2XL U7829 ( .A(n7426), .B(n7407), .Z(n7409) );
  CANR1XL U7830 ( .A(n7407), .B(n7314), .C(n7406), .Z(n7408) );
  COND1XL U7831 ( .A(n7409), .B(n2623), .C(n7408), .Z(n7413) );
  CND2X1 U7832 ( .A(n7411), .B(n7410), .Z(n7412) );
  CENXL U7833 ( .A(n7413), .B(n7412), .Z(N76) );
  CND2XL U7834 ( .A(n7414), .B(n7417), .Z(n7419) );
  CANR1XL U7835 ( .A(n7417), .B(n7416), .C(n7415), .Z(n7418) );
  COND1XL U7836 ( .A(n7419), .B(n7485), .C(n7418), .Z(n7424) );
  CIVXL U7837 ( .A(n7420), .Z(n7422) );
  CND2X1 U7838 ( .A(n7422), .B(n7421), .Z(n7423) );
  CENXL U7839 ( .A(n7424), .B(n7423), .Z(N63) );
  CIVXL U7840 ( .A(n7425), .Z(n7429) );
  CND2XL U7841 ( .A(n7426), .B(n7429), .Z(n7431) );
  CIVXL U7842 ( .A(n2352), .Z(n7428) );
  CANR1XL U7843 ( .A(n7429), .B(n7314), .C(n7428), .Z(n7430) );
  COND1XL U7844 ( .A(n7431), .B(n2623), .C(n7430), .Z(n7435) );
  CND2X1 U7845 ( .A(n7192), .B(n7433), .Z(n7434) );
  CENXL U7846 ( .A(n7435), .B(n7434), .Z(N68) );
  CND2XL U7847 ( .A(n7436), .B(n7439), .Z(n7441) );
  CANR1XL U7848 ( .A(n7439), .B(n7438), .C(n7437), .Z(n7440) );
  COND1XL U7849 ( .A(n7441), .B(n7485), .C(n7440), .Z(n7445) );
  CND2XL U7850 ( .A(n7443), .B(n7442), .Z(n7444) );
  CENXL U7851 ( .A(n7445), .B(n7444), .Z(N60) );
  CIVXL U7852 ( .A(n7446), .Z(n7447) );
  COND1XL U7853 ( .A(n7448), .B(n2623), .C(n7447), .Z(n7452) );
  CND2X1 U7854 ( .A(n7450), .B(n7449), .Z(n7451) );
  CENXL U7855 ( .A(n7452), .B(n7451), .Z(N70) );
  CIVX2 U7856 ( .A(n7453), .Z(n7455) );
  COND1XL U7857 ( .A(n7455), .B(n7485), .C(n7454), .Z(n7459) );
  CND2XL U7858 ( .A(n7457), .B(n7456), .Z(n7458) );
  CENXL U7859 ( .A(n7459), .B(n7458), .Z(N56) );
  CIVXL U7860 ( .A(n7460), .Z(n7473) );
  CND2XL U7861 ( .A(n7473), .B(n1550), .Z(n7464) );
  CIVXL U7862 ( .A(n7469), .Z(n7462) );
  CIVXL U7863 ( .A(n7472), .Z(n7461) );
  CENXL U7864 ( .A(n7464), .B(n7463), .Z(N49) );
  COR2XL U7865 ( .A(n7465), .B(n7466), .Z(n7467) );
  CND2XL U7866 ( .A(n7468), .B(n7467), .Z(n7478) );
  CND2XL U7867 ( .A(n7469), .B(n7473), .Z(n7476) );
  CIVXL U7868 ( .A(n1539), .Z(n7471) );
  CANR1XL U7869 ( .A(n7473), .B(n2530), .C(n7471), .Z(n7474) );
  CENXL U7870 ( .A(n7478), .B(n7477), .Z(N50) );
  CND2XL U7871 ( .A(n7479), .B(n7483), .Z(n7486) );
  CIVXL U7872 ( .A(n7480), .Z(n7481) );
  CANR1XL U7873 ( .A(n7483), .B(n7482), .C(n7481), .Z(n7484) );
  COAN1XL U7874 ( .A(n7486), .B(n7485), .C(n7484), .Z(N78) );
  CIVXL U7875 ( .A(n7487), .Z(n7488) );
  CND2XL U7876 ( .A(n7488), .B(n7492), .Z(n7495) );
  CIVDXL U7877 ( .A(n2314), .Z0(n7008), .Z1(n7491) );
  CENXL U7878 ( .A(n7499), .B(n7498), .Z(N42) );
  CIVXL U7879 ( .A(n7500), .Z(n7505) );
  CND2X1 U7880 ( .A(n7507), .B(n7506), .Z(n7509) );
  CENX1 U7881 ( .A(n7509), .B(n7508), .Z(N22) );
  CND2XL U7882 ( .A(n7511), .B(n7510), .Z(n7512) );
  CENXL U7883 ( .A(n7512), .B(n7513), .Z(N43) );
  CIVXL U7884 ( .A(n7514), .Z(n7532) );
  CIVX1 U7885 ( .A(n7515), .Z(n7517) );
  CND2X1 U7886 ( .A(n7517), .B(n7516), .Z(n7518) );
  CEOXL U7887 ( .A(n7519), .B(n7518), .Z(N23) );
  CIVX2 U7888 ( .A(n7520), .Z(n7522) );
  CND2X1 U7889 ( .A(n7522), .B(n7521), .Z(n7523) );
  CEOXL U7890 ( .A(n7524), .B(n7523), .Z(N21) );
  CMX2XL U7891 ( .A0(n7539), .A1(h[0]), .S(n7682), .Z(n917) );
  CIVXL U7892 ( .A(n7681), .Z(n8021) );
  CMX2XL U7893 ( .A0(h0_0[4]), .A1(n2513), .S(cmd2_en_0), .Z(n928) );
  CMX2XL U7894 ( .A0(h0_0[0]), .A1(n7539), .S(cmd2_en_0), .Z(n916) );
  CMX2XL U7895 ( .A0(h0_0[2]), .A1(h0[2]), .S(cmd2_en_0), .Z(n922) );
  CMX2XL U7896 ( .A0(h0_0[3]), .A1(n1232), .S(cmd2_en_0), .Z(n925) );
  CMX2XL U7897 ( .A0(h0_0[6]), .A1(n7674), .S(cmd2_en_0), .Z(n934) );
  CIVXL U7898 ( .A(n7540), .Z(n7698) );
  COND2XL U7899 ( .A(n7727), .B(n7713), .C(n7729), .D(n7544), .Z(n7546) );
  CANR1XL U7900 ( .A(n7726), .B(n7712), .C(n7724), .Z(n7545) );
  COND2XL U7901 ( .A(n2865), .B(n7999), .C(n7546), .D(n7545), .Z(n889) );
  COND2XL U7902 ( .A(n7727), .B(n7717), .C(n7729), .D(n7547), .Z(n7549) );
  CANR1XL U7903 ( .A(n7726), .B(n7716), .C(n7724), .Z(n7548) );
  COND2XL U7904 ( .A(n2865), .B(n7998), .C(n7549), .D(n7548), .Z(n853) );
  COND2XL U7905 ( .A(n2865), .B(n7955), .C(n7741), .D(n7722), .Z(n910) );
  CND3XL U7906 ( .A(n7551), .B(h0_1[4]), .C(n7550), .Z(n7562) );
  COND2XL U7907 ( .A(n7770), .B(n7748), .C(n7763), .D(n7765), .Z(n7555) );
  COND2XL U7908 ( .A(n7766), .B(n7552), .C(n2663), .D(n7769), .Z(n7554) );
  CNR2XL U7909 ( .A(n7553), .B(h0_1[4]), .Z(n7772) );
  CANR4CXL U7910 ( .A(n7555), .B(n7554), .C(n7772), .D(n7771), .Z(n7561) );
  COND2XL U7911 ( .A(n7758), .B(n7557), .C(n7556), .D(n7744), .Z(n7558) );
  COND4CXL U7912 ( .A(n7762), .B(n7559), .C(n7558), .D(n8020), .Z(n7560) );
  CND3XL U7913 ( .A(n7562), .B(n7561), .C(n7560), .Z(n7564) );
  CANR2XL U7914 ( .A(n7720), .B(n7780), .C(out2_2[2]), .D(n7751), .Z(n7563) );
  COND3XL U7915 ( .A(n7723), .B(n7565), .C(n7564), .D(n7563), .Z(n885) );
  CIVXL U7916 ( .A(n7566), .Z(n7568) );
  CND2XL U7917 ( .A(n7568), .B(n7567), .Z(n7572) );
  CANR1XL U7918 ( .A(n7570), .B(n7806), .C(n7569), .Z(n7571) );
  CEOXL U7919 ( .A(n7572), .B(n7571), .Z(n7573) );
  CMX2XL U7920 ( .A0(out1_2[24]), .A1(n7573), .S(cmd1_en_2), .Z(n7911) );
  CANR2XL U7921 ( .A(n7747), .B(n7575), .C(n7762), .D(n7574), .Z(n7579) );
  CANR2XL U7922 ( .A(n7582), .B(n7577), .C(n7755), .D(n7576), .Z(n7578) );
  CND2XL U7923 ( .A(n7579), .B(n7578), .Z(n7753) );
  CANR2XL U7924 ( .A(n7582), .B(n7581), .C(n7755), .D(n7580), .Z(n7586) );
  CANR2XL U7925 ( .A(n2859), .B(n7584), .C(n7747), .D(n7583), .Z(n7585) );
  CND2XL U7926 ( .A(n7586), .B(n7585), .Z(n7750) );
  COND2XL U7927 ( .A(n7727), .B(n7753), .C(n7750), .D(n7729), .Z(n7588) );
  CANR1XL U7928 ( .A(n7726), .B(n7752), .C(n7724), .Z(n7587) );
  COND2XL U7929 ( .A(n2865), .B(n8000), .C(n7588), .D(n7587), .Z(n864) );
  CIVXL U7930 ( .A(n7589), .Z(n7591) );
  CND2XL U7931 ( .A(n7591), .B(n7590), .Z(n7602) );
  CIVXL U7932 ( .A(n7592), .Z(n7617) );
  CND2XL U7933 ( .A(n7617), .B(n7596), .Z(n7598) );
  CNR2XL U7934 ( .A(n7635), .B(n7598), .Z(n7600) );
  CIVXL U7935 ( .A(n7593), .Z(n7624) );
  CIVXL U7936 ( .A(n7594), .Z(n7595) );
  CANR1XL U7937 ( .A(n7596), .B(n7624), .C(n7595), .Z(n7597) );
  COND1XL U7938 ( .A(n7598), .B(n7638), .C(n7597), .Z(n7599) );
  CANR1XL U7939 ( .A(n7600), .B(n7806), .C(n7599), .Z(n7601) );
  CEOXL U7940 ( .A(n7602), .B(n7601), .Z(n7603) );
  CMX2XL U7941 ( .A0(out1_2[29]), .A1(n7603), .S(cmd1_en_2), .Z(n7906) );
  CIVXL U7942 ( .A(n7621), .Z(n7604) );
  CND2XL U7943 ( .A(n7604), .B(n7619), .Z(n7610) );
  CND2XL U7944 ( .A(n7617), .B(n7615), .Z(n7606) );
  CNR2XL U7945 ( .A(n7635), .B(n7606), .Z(n7608) );
  CANR1XL U7946 ( .A(n7615), .B(n7624), .C(n7618), .Z(n7605) );
  COND1XL U7947 ( .A(n7606), .B(n7638), .C(n7605), .Z(n7607) );
  CANR1XL U7948 ( .A(n7608), .B(n7806), .C(n7607), .Z(n7609) );
  CEOXL U7949 ( .A(n7610), .B(n7609), .Z(n7611) );
  CMX2XL U7950 ( .A0(out1_2[30]), .A1(n7611), .S(cmd1_en_2), .Z(n7905) );
  CIVXL U7951 ( .A(n7612), .Z(n7614) );
  CND2XL U7952 ( .A(n7614), .B(n7613), .Z(n7630) );
  CIVXL U7953 ( .A(n7615), .Z(n7616) );
  CNR2XL U7954 ( .A(n7616), .B(n7621), .Z(n7623) );
  CND2XL U7955 ( .A(n7623), .B(n7617), .Z(n7626) );
  CNR2XL U7956 ( .A(n7635), .B(n7626), .Z(n7628) );
  CIVXL U7957 ( .A(n7618), .Z(n7620) );
  COND1XL U7958 ( .A(n7621), .B(n7620), .C(n7619), .Z(n7622) );
  CANR1XL U7959 ( .A(n7624), .B(n7623), .C(n7622), .Z(n7625) );
  COND1XL U7960 ( .A(n7626), .B(n7638), .C(n7625), .Z(n7627) );
  CANR1XL U7961 ( .A(n7628), .B(n7806), .C(n7627), .Z(n7629) );
  CEOXL U7962 ( .A(n7630), .B(n7629), .Z(n7631) );
  CMX2XL U7963 ( .A0(out1_2[31]), .A1(n7631), .S(cmd1_en_2), .Z(n7904) );
  CND2XL U7964 ( .A(n7633), .B(n7632), .Z(n7643) );
  CIVXL U7965 ( .A(n7634), .Z(n7639) );
  CNR2XL U7966 ( .A(n7635), .B(n7639), .Z(n7641) );
  CIVXL U7967 ( .A(n7636), .Z(n7637) );
  COND1XL U7968 ( .A(n7639), .B(n7638), .C(n7637), .Z(n7640) );
  CANR1XL U7969 ( .A(n7641), .B(n7806), .C(n7640), .Z(n7642) );
  CEOXL U7970 ( .A(n7643), .B(n7642), .Z(n7644) );
  CMX2XL U7971 ( .A0(out1_2[26]), .A1(n7644), .S(cmd1_en_2), .Z(n7909) );
  CIVXL U7972 ( .A(n7645), .Z(n7647) );
  CND2XL U7973 ( .A(n7647), .B(n7646), .Z(n7651) );
  CANR1XL U7974 ( .A(n7649), .B(n3949), .C(n7648), .Z(n7650) );
  CEOXL U7975 ( .A(n7651), .B(n7650), .Z(n7652) );
  CMX2XL U7976 ( .A0(out1_2[40]), .A1(n7652), .S(cmd1_en_2), .Z(n7895) );
  CND2XL U7977 ( .A(n7654), .B(n7653), .Z(n7664) );
  CIVXL U7978 ( .A(n7655), .Z(n7660) );
  CNR2XL U7979 ( .A(n7656), .B(n7660), .Z(n7662) );
  CIVXL U7980 ( .A(n7657), .Z(n7658) );
  COND1XL U7981 ( .A(n7660), .B(n7659), .C(n7658), .Z(n7661) );
  CANR1XL U7982 ( .A(n7662), .B(n3949), .C(n7661), .Z(n7663) );
  CEOXL U7983 ( .A(n7664), .B(n7663), .Z(n7665) );
  CMX2XL U7984 ( .A0(out1_2[42]), .A1(n7665), .S(cmd1_en_2), .Z(n7893) );
  CIVXL U7985 ( .A(n7666), .Z(n7668) );
  CND2XL U7986 ( .A(n7668), .B(n7667), .Z(n7672) );
  CANR1XL U7987 ( .A(n7670), .B(n3949), .C(n7669), .Z(n7671) );
  CEOXL U7988 ( .A(n7672), .B(n7671), .Z(n7673) );
  CMX2XL U7989 ( .A0(out1_2[34]), .A1(n7673), .S(cmd1_en_2), .Z(n7901) );
  CMX2X1 U7990 ( .A0(h0[28]), .A1(h[28]), .S(n7682), .Z(n957) );
  CMX2X1 U7991 ( .A0(h0[23]), .A1(h[23]), .S(n7682), .Z(n952) );
  CMX2X1 U7992 ( .A0(n7674), .A1(h[6]), .S(n7682), .Z(n935) );
  CMX2X1 U7993 ( .A0(h0[20]), .A1(h[20]), .S(pushin), .Z(n949) );
  CAOR2XL U7994 ( .A(out2_2[63]), .B(n7751), .C(n7700), .D(n7738), .Z(n882) );
  CIVX1 U7995 ( .A(n7675), .Z(n7696) );
  CAOR2XL U7996 ( .A(out2_2[62]), .B(n7751), .C(n7692), .D(n7738), .Z(n914) );
  CAOR2XL U7997 ( .A(out2_2[51]), .B(n7751), .C(n7705), .D(n7738), .Z(n876) );
  CND2IXL U7998 ( .B(cmd0[1]), .A(n1489), .Z(n7676) );
  CNR2IXL U7999 ( .B(n1335), .A(n7676), .Z(cmd1_en_0) );
  CMX2XL U8000 ( .A0(cmd0_en_1), .A1(cmd0_en_2), .S(rst), .Z(n1188) );
  CNR2XL U8001 ( .A(n1335), .B(n7676), .Z(cmd0_en_0) );
  CMX2XL U8002 ( .A0(out0_2[59]), .A1(out1_1[59]), .S(cmd0_en_2), .Z(n1125) );
  CMX2XL U8003 ( .A0(out0_2[42]), .A1(out1_1[42]), .S(cmd0_en_2), .Z(n1142) );
  CMX2XL U8004 ( .A0(out0_2[48]), .A1(out1_1[48]), .S(cmd0_en_2), .Z(n1136) );
  CMX2XL U8005 ( .A0(out0_2[46]), .A1(out1_1[46]), .S(cmd0_en_2), .Z(n1138) );
  CMX2XL U8006 ( .A0(out0_2[57]), .A1(out1_1[57]), .S(cmd0_en_2), .Z(n1127) );
  CMX2XL U8007 ( .A0(out0_2[36]), .A1(out1_1[36]), .S(cmd0_en_2), .Z(n1148) );
  CMX2XL U8008 ( .A0(n7677), .A1(out1_1[52]), .S(cmd0_en_2), .Z(n1132) );
  CMX2XL U8009 ( .A0(n7678), .A1(out1_1[53]), .S(cmd0_en_2), .Z(n1131) );
  CMX2XL U8010 ( .A0(n4323), .A1(out1_1[55]), .S(cmd0_en_2), .Z(n1129) );
  CMX2XL U8011 ( .A0(out0_2[56]), .A1(out1_1[56]), .S(cmd0_en_2), .Z(n1128) );
  CMX2XL U8012 ( .A0(n1369), .A1(out1_1[40]), .S(cmd0_en_2), .Z(n1144) );
  CMX2XL U8013 ( .A0(out0_2[50]), .A1(out1_1[50]), .S(cmd0_en_2), .Z(n1134) );
  CMX2XL U8014 ( .A0(out0_2[49]), .A1(out1_1[49]), .S(cmd0_en_2), .Z(n1135) );
  CMX2XL U8015 ( .A0(out0_2[51]), .A1(out1_1[51]), .S(cmd0_en_2), .Z(n1133) );
  CMX2XL U8016 ( .A0(out0_2[60]), .A1(out1_1[60]), .S(cmd0_en_2), .Z(n1124) );
  CMX2XL U8017 ( .A0(out0_2[54]), .A1(out1_1[54]), .S(cmd0_en_2), .Z(n1130) );
  CMX2XL U8018 ( .A0(out0_2[61]), .A1(out1_1[61]), .S(cmd0_en_2), .Z(n1123) );
  CMX2XL U8019 ( .A0(out0_2[62]), .A1(out1_1[62]), .S(cmd0_en_2), .Z(n1122) );
  CMX2XL U8020 ( .A0(out0_2[58]), .A1(out1_1[58]), .S(cmd0_en_2), .Z(n1126) );
  CMX2XL U8021 ( .A0(out0_2[63]), .A1(out1_1[63]), .S(cmd0_en_2), .Z(n1121) );
  CMX2XL U8022 ( .A0(h0[5]), .A1(h[5]), .S(pushin), .Z(n932) );
  CMX2XL U8023 ( .A0(n2512), .A1(h[4]), .S(pushin), .Z(n929) );
  CMX2XL U8024 ( .A0(h0[2]), .A1(h[2]), .S(pushin), .Z(n923) );
  CMX2XL U8025 ( .A0(h0_1[2]), .A1(h0_0[2]), .S(cmd2_en_1), .Z(n921) );
  CMX2XL U8026 ( .A0(n7680), .A1(h0_0[3]), .S(cmd2_en_1), .Z(n924) );
  CMX2XL U8027 ( .A0(acc[28]), .A1(z[28]), .S(n7681), .Z(n1217) );
  CMX2XL U8028 ( .A0(acc[29]), .A1(z[29]), .S(n7681), .Z(n1218) );
  CMX2XL U8029 ( .A0(acc[30]), .A1(z[30]), .S(n7681), .Z(n1219) );
  CMX2XL U8030 ( .A0(acc[31]), .A1(z[31]), .S(n7681), .Z(n1220) );
  CMX2XL U8031 ( .A0(acc[26]), .A1(z[26]), .S(n7681), .Z(n1215) );
  CMX2XL U8032 ( .A0(acc[27]), .A1(z[27]), .S(n7681), .Z(n1216) );
  CMX2XL U8033 ( .A0(acc[20]), .A1(z[20]), .S(n7681), .Z(n1209) );
  CMX2XL U8034 ( .A0(acc[21]), .A1(z[21]), .S(n7681), .Z(n1210) );
  CMX2XL U8035 ( .A0(acc[23]), .A1(z[23]), .S(n7681), .Z(n1212) );
  CMX2XL U8036 ( .A0(acc[25]), .A1(z[25]), .S(n7681), .Z(n1214) );
  CMX2XL U8037 ( .A0(acc[6]), .A1(z[6]), .S(n7681), .Z(n1195) );
  CMX2XL U8038 ( .A0(acc[7]), .A1(z[7]), .S(n7681), .Z(n1196) );
  CMX2XL U8039 ( .A0(acc[22]), .A1(z[22]), .S(n7681), .Z(n1211) );
  CMX2XL U8040 ( .A0(acc[13]), .A1(z[13]), .S(n7681), .Z(n1202) );
  CMX2XL U8041 ( .A0(acc[3]), .A1(z[3]), .S(n7681), .Z(n1192) );
  CMX2XL U8042 ( .A0(acc[5]), .A1(z[5]), .S(n7681), .Z(n1194) );
  CMX2XL U8043 ( .A0(acc[18]), .A1(z[18]), .S(n7681), .Z(n1207) );
  CMX2XL U8044 ( .A0(acc[19]), .A1(z[19]), .S(n7681), .Z(n1208) );
  CMX2XL U8045 ( .A0(acc[14]), .A1(z[14]), .S(n7681), .Z(n1203) );
  CMX2XL U8046 ( .A0(acc[15]), .A1(z[15]), .S(n7681), .Z(n1204) );
  CMX2XL U8047 ( .A0(q0[0]), .A1(q[0]), .S(n7682), .Z(n961) );
  COND2XL U8048 ( .A(n2865), .B(n7942), .C(n7683), .D(n7722), .Z(n913) );
  COND2XL U8049 ( .A(n2865), .B(n7945), .C(n7684), .D(n7722), .Z(n880) );
  COND2XL U8050 ( .A(n2865), .B(n7951), .C(n7685), .D(n7722), .Z(n911) );
  CIVXL U8051 ( .A(n7728), .Z(n7687) );
  CANR2XL U8052 ( .A(n7725), .B(n7704), .C(out2_2[41]), .D(n7751), .Z(n7686)
         );
  COND1XL U8053 ( .A(n7722), .B(n7687), .C(n7686), .Z(n862) );
  CIVXL U8054 ( .A(n7688), .Z(n7691) );
  CANR2XL U8055 ( .A(n7689), .B(n7704), .C(out2_2[37]), .D(n7751), .Z(n7690)
         );
  COND1XL U8056 ( .A(n7722), .B(n7691), .C(n7690), .Z(n870) );
  CIVXL U8057 ( .A(n7692), .Z(n7695) );
  CANR2XL U8058 ( .A(n7693), .B(n7738), .C(out2_2[46]), .D(n7751), .Z(n7694)
         );
  COND1XL U8059 ( .A(n7742), .B(n7695), .C(n7694), .Z(n906) );
  CANR2XL U8060 ( .A(n7696), .B(n7704), .C(out2_2[45]), .D(n7751), .Z(n7697)
         );
  COND1XL U8061 ( .A(n7722), .B(n7698), .C(n7697), .Z(n873) );
  CIVXL U8062 ( .A(n7699), .Z(n7702) );
  CANR2XL U8063 ( .A(n7700), .B(n7704), .C(out2_2[47]), .D(n7751), .Z(n7701)
         );
  COND1XL U8064 ( .A(n7722), .B(n7702), .C(n7701), .Z(n874) );
  CIVXL U8065 ( .A(n7703), .Z(n7707) );
  CANR2XL U8066 ( .A(n7705), .B(n7704), .C(out2_2[35]), .D(n7751), .Z(n7706)
         );
  COND1XL U8067 ( .A(n7707), .B(n7722), .C(n7706), .Z(n859) );
  CIVXL U8068 ( .A(n7752), .Z(n7709) );
  CANR2XL U8069 ( .A(n7753), .B(n7738), .C(out2_2[33]), .D(n7751), .Z(n7708)
         );
  COND1XL U8070 ( .A(n7709), .B(n7742), .C(n7708), .Z(n866) );
  CIVXL U8071 ( .A(n7779), .Z(n7711) );
  CANR2XL U8072 ( .A(n7781), .B(n7738), .C(out2_2[32]), .D(n7751), .Z(n7710)
         );
  COND1XL U8073 ( .A(n7711), .B(n7742), .C(n7710), .Z(n901) );
  CIVXL U8074 ( .A(n7712), .Z(n7715) );
  CANR2XL U8075 ( .A(n7713), .B(n7738), .C(out2_2[36]), .D(n7751), .Z(n7714)
         );
  COND1XL U8076 ( .A(n7715), .B(n7742), .C(n7714), .Z(n900) );
  CIVXL U8077 ( .A(n7716), .Z(n7719) );
  CANR2XL U8078 ( .A(n7717), .B(n7738), .C(out2_2[39]), .D(n7751), .Z(n7718)
         );
  COND1XL U8079 ( .A(n7719), .B(n7742), .C(n7718), .Z(n854) );
  COND2XL U8080 ( .A(n2865), .B(n7947), .C(n7737), .D(n7722), .Z(n912) );
  CANR2XL U8081 ( .A(n7720), .B(n7738), .C(out2_2[34]), .D(n7751), .Z(n7721)
         );
  COND1XL U8082 ( .A(n7742), .B(n7723), .C(n7721), .Z(n897) );
  COND2XL U8083 ( .A(n2865), .B(n7963), .C(n7723), .D(n7722), .Z(n905) );
  CANR1XL U8084 ( .A(n7726), .B(n7725), .C(n7724), .Z(n7734) );
  CNR2XL U8085 ( .A(n7728), .B(n7727), .Z(n7733) );
  CNR2XL U8086 ( .A(n7730), .B(n7729), .Z(n7732) );
  CND2XL U8087 ( .A(n7751), .B(out2_2[25]), .Z(n7731) );
  CANR2XL U8088 ( .A(n7735), .B(n7738), .C(out2_2[42]), .D(n7751), .Z(n7736)
         );
  COND1XL U8089 ( .A(n7742), .B(n7737), .C(n7736), .Z(n904) );
  CANR2XL U8090 ( .A(n7739), .B(n7738), .C(out2_2[38]), .D(n7751), .Z(n7740)
         );
  COND1XL U8091 ( .A(n7742), .B(n7741), .C(n7740), .Z(n902) );
  CIVXL U8092 ( .A(n7749), .Z(n7764) );
  CND3XL U8093 ( .A(n7756), .B(n7755), .C(n7754), .Z(n7757) );
  COND1XL U8094 ( .A(n7759), .B(n7758), .C(n7757), .Z(n7760) );
  COND4CXL U8095 ( .A(n7762), .B(n7761), .C(n7760), .D(n8020), .Z(n7776) );
  COND2XL U8096 ( .A(n7766), .B(n7765), .C(n7764), .D(n7763), .Z(n7774) );
  CIVXL U8097 ( .A(n7767), .Z(n7768) );
  COND2XL U8098 ( .A(n7770), .B(n7769), .C(n7768), .D(n2663), .Z(n7773) );
  CANR4CXL U8099 ( .A(n7774), .B(n7773), .C(n7772), .D(n7771), .Z(n7775) );
  COND3XL U8100 ( .A(n7777), .B(n8020), .C(n7776), .D(n7775), .Z(n7784) );
  CANR2XL U8101 ( .A(n7779), .B(n7778), .C(out2_2[0]), .D(n7751), .Z(n7783) );
  CND2XL U8102 ( .A(n7781), .B(n7780), .Z(n7782) );
  CND3XL U8103 ( .A(n7784), .B(n7783), .C(n7782), .Z(n892) );
  CIVXL U8104 ( .A(n7793), .Z(n7795) );
  CND2XL U8105 ( .A(n7795), .B(n7794), .Z(n7801) );
  CIVXL U8106 ( .A(n7807), .Z(n7796) );
  CNR2XL U8107 ( .A(n7796), .B(n7803), .Z(n7799) );
  CIVXL U8108 ( .A(n7805), .Z(n7797) );
  COND1XL U8109 ( .A(n7803), .B(n7797), .C(n7804), .Z(n7798) );
  CANR1XL U8110 ( .A(n7799), .B(n7806), .C(n7798), .Z(n7800) );
  CEOXL U8111 ( .A(n7801), .B(n7800), .Z(n7802) );
  CMX2XL U8112 ( .A0(out1_2[19]), .A1(n7802), .S(n8022), .Z(n7916) );
  CIVXL U8113 ( .A(acc[63]), .Z(n7811) );
  CANR2XL U8114 ( .A(n7808), .B(out0_2[63]), .C(out1_2[63]), .D(cmd1_en_2_d), 
        .Z(n7809) );
  COND1XL U8115 ( .A(n7811), .B(n7810), .C(n7809), .Z(n7812) );
  COR2XL U8116 ( .A(n7812), .B(out1_1[63]), .Z(n7814) );
  CND2XL U8117 ( .A(n7812), .B(out1_1[63]), .Z(n7813) );
  CND2X1 U8118 ( .A(n7814), .B(n7813), .Z(n7835) );
  CND2XL U8119 ( .A(n7815), .B(n7822), .Z(n7825) );
  CNR2XL U8120 ( .A(n7816), .B(n7825), .Z(n7828) );
  CND2XL U8121 ( .A(n7817), .B(n7828), .Z(n7831) );
  CNR2XL U8122 ( .A(n7818), .B(n7831), .Z(n7833) );
  CIVXL U8123 ( .A(n7819), .Z(n7820) );
  CANR1XL U8124 ( .A(n7822), .B(n7821), .C(n7820), .Z(n7823) );
  COND1XL U8125 ( .A(n7825), .B(n7824), .C(n7823), .Z(n7826) );
  CANR1XL U8126 ( .A(n7828), .B(n7827), .C(n7826), .Z(n7829) );
  COND1XL U8127 ( .A(n7831), .B(n7830), .C(n7829), .Z(n7832) );
  CANR1XL U8128 ( .A(n7833), .B(n3949), .C(n7832), .Z(n7834) );
  CEOXL U8129 ( .A(n7835), .B(n7834), .Z(n7836) );
  CMXI2XL U8130 ( .A0(out1_2[63]), .A1(n7836), .S(n7846), .Z(n7837) );
  CIVXL U8131 ( .A(n7837), .Z(n1057) );
endmodule

