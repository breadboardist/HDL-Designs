
module sfilt_DW01_add_0 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63;

  CAN2X1 U1 ( .A(A[39]), .B(n2), .Z(n1) );
  CAN2X1 U2 ( .A(A[38]), .B(n57), .Z(n2) );
  CAN2X1 U3 ( .A(A[31]), .B(n4), .Z(n3) );
  CAN2X1 U4 ( .A(A[30]), .B(n63), .Z(n4) );
  CAN2X1 U5 ( .A(A[28]), .B(n6), .Z(n5) );
  CAN2X1 U6 ( .A(A[27]), .B(n7), .Z(n6) );
  CAN2X1 U7 ( .A(A[26]), .B(n8), .Z(n7) );
  CAN2X1 U8 ( .A(A[25]), .B(n9), .Z(n8) );
  CAN2X1 U9 ( .A(A[24]), .B(n10), .Z(n9) );
  CAN2X1 U10 ( .A(A[23]), .B(n11), .Z(n10) );
  CAN2X1 U11 ( .A(A[22]), .B(n12), .Z(n11) );
  CAN2X1 U12 ( .A(A[21]), .B(n13), .Z(n12) );
  CAN2X1 U13 ( .A(A[20]), .B(n14), .Z(n13) );
  CAN2X1 U14 ( .A(A[19]), .B(n15), .Z(n14) );
  CAN2X1 U15 ( .A(A[18]), .B(n16), .Z(n15) );
  CAN2X1 U16 ( .A(A[17]), .B(n17), .Z(n16) );
  CAN2X1 U17 ( .A(A[16]), .B(n18), .Z(n17) );
  CAN2X1 U18 ( .A(A[15]), .B(n19), .Z(n18) );
  CAN2X1 U19 ( .A(A[14]), .B(n20), .Z(n19) );
  CAN2X1 U20 ( .A(A[13]), .B(n21), .Z(n20) );
  CAN2X1 U21 ( .A(A[12]), .B(n22), .Z(n21) );
  CAN2X1 U22 ( .A(A[11]), .B(n23), .Z(n22) );
  CAN2X1 U23 ( .A(A[10]), .B(n24), .Z(n23) );
  CAN2X1 U24 ( .A(A[9]), .B(n25), .Z(n24) );
  CAN2X1 U25 ( .A(A[8]), .B(n26), .Z(n25) );
  CAN2X1 U26 ( .A(A[7]), .B(n27), .Z(n26) );
  CAN2X1 U27 ( .A(A[6]), .B(n28), .Z(n27) );
  CAN2X1 U28 ( .A(A[5]), .B(n29), .Z(n28) );
  CAN2X1 U29 ( .A(A[4]), .B(n30), .Z(n29) );
  CAN2X1 U30 ( .A(A[3]), .B(n31), .Z(n30) );
  CAN2X1 U31 ( .A(A[2]), .B(n32), .Z(n31) );
  CAN2X1 U32 ( .A(A[1]), .B(n33), .Z(n32) );
  CAN2X1 U33 ( .A(B[0]), .B(A[0]), .Z(n33) );
  CAN2X1 U34 ( .A(A[62]), .B(n36), .Z(n34) );
  CAN2X1 U35 ( .A(A[60]), .B(n37), .Z(n35) );
  CAN2X1 U36 ( .A(A[61]), .B(n35), .Z(n36) );
  CAN2X1 U37 ( .A(A[59]), .B(n38), .Z(n37) );
  CAN2X1 U38 ( .A(A[58]), .B(n39), .Z(n38) );
  CAN2X1 U39 ( .A(A[57]), .B(n40), .Z(n39) );
  CAN2X1 U40 ( .A(A[56]), .B(n41), .Z(n40) );
  CAN2X1 U41 ( .A(A[55]), .B(n42), .Z(n41) );
  CAN2X1 U42 ( .A(A[54]), .B(n43), .Z(n42) );
  CAN2X1 U43 ( .A(A[53]), .B(n44), .Z(n43) );
  CAN2X1 U44 ( .A(A[52]), .B(n45), .Z(n44) );
  CAN2X1 U45 ( .A(A[51]), .B(n46), .Z(n45) );
  CAN2X1 U46 ( .A(A[50]), .B(n47), .Z(n46) );
  CAN2X1 U47 ( .A(A[49]), .B(n48), .Z(n47) );
  CAN2X1 U48 ( .A(A[48]), .B(n49), .Z(n48) );
  CAN2X1 U49 ( .A(A[47]), .B(n50), .Z(n49) );
  CAN2X1 U50 ( .A(A[46]), .B(n51), .Z(n50) );
  CAN2X1 U51 ( .A(A[45]), .B(n52), .Z(n51) );
  CAN2X1 U52 ( .A(A[44]), .B(n53), .Z(n52) );
  CAN2X1 U53 ( .A(A[43]), .B(n54), .Z(n53) );
  CAN2X1 U54 ( .A(A[42]), .B(n55), .Z(n54) );
  CAN2X1 U55 ( .A(A[41]), .B(n56), .Z(n55) );
  CAN2X1 U56 ( .A(A[40]), .B(n1), .Z(n56) );
  CAN2X1 U57 ( .A(A[37]), .B(n58), .Z(n57) );
  CAN2X1 U58 ( .A(A[36]), .B(n59), .Z(n58) );
  CAN2X1 U59 ( .A(A[35]), .B(n60), .Z(n59) );
  CAN2X1 U60 ( .A(A[34]), .B(n61), .Z(n60) );
  CAN2X1 U61 ( .A(A[33]), .B(n62), .Z(n61) );
  CAN2X1 U62 ( .A(A[32]), .B(n3), .Z(n62) );
  CAN2X1 U63 ( .A(A[29]), .B(n5), .Z(n63) );
  CEOX1 U64 ( .A(A[61]), .B(n35), .Z(SUM[61]) );
  CEOX1 U65 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  CEOX1 U66 ( .A(A[63]), .B(n34), .Z(SUM[63]) );
  CEOX1 U67 ( .A(A[62]), .B(n36), .Z(SUM[62]) );
  CEOX1 U68 ( .A(A[60]), .B(n37), .Z(SUM[60]) );
  CEOX1 U69 ( .A(A[59]), .B(n38), .Z(SUM[59]) );
  CEOX1 U70 ( .A(A[58]), .B(n39), .Z(SUM[58]) );
  CEOX1 U71 ( .A(A[57]), .B(n40), .Z(SUM[57]) );
  CEOX1 U72 ( .A(A[56]), .B(n41), .Z(SUM[56]) );
  CEOX1 U73 ( .A(A[55]), .B(n42), .Z(SUM[55]) );
  CEOX1 U74 ( .A(A[54]), .B(n43), .Z(SUM[54]) );
  CEOX1 U75 ( .A(A[53]), .B(n44), .Z(SUM[53]) );
  CEOX1 U76 ( .A(A[52]), .B(n45), .Z(SUM[52]) );
  CEOX1 U77 ( .A(A[51]), .B(n46), .Z(SUM[51]) );
  CEOX1 U78 ( .A(A[50]), .B(n47), .Z(SUM[50]) );
  CEOX1 U79 ( .A(A[49]), .B(n48), .Z(SUM[49]) );
  CEOX1 U80 ( .A(A[46]), .B(n51), .Z(SUM[46]) );
  CEOX1 U81 ( .A(A[48]), .B(n49), .Z(SUM[48]) );
  CEOX1 U82 ( .A(A[47]), .B(n50), .Z(SUM[47]) );
  CEOX1 U83 ( .A(A[45]), .B(n52), .Z(SUM[45]) );
  CEOX1 U84 ( .A(A[42]), .B(n55), .Z(SUM[42]) );
  CEOX1 U85 ( .A(A[44]), .B(n53), .Z(SUM[44]) );
  CEOX1 U86 ( .A(A[43]), .B(n54), .Z(SUM[43]) );
  CEOX1 U87 ( .A(A[41]), .B(n56), .Z(SUM[41]) );
  CEOX1 U88 ( .A(A[40]), .B(n1), .Z(SUM[40]) );
  CEOX1 U89 ( .A(A[39]), .B(n2), .Z(SUM[39]) );
  CEOX1 U90 ( .A(A[38]), .B(n57), .Z(SUM[38]) );
  CEOX1 U91 ( .A(A[37]), .B(n58), .Z(SUM[37]) );
  CEOX1 U92 ( .A(A[36]), .B(n59), .Z(SUM[36]) );
  CEOX1 U93 ( .A(A[35]), .B(n60), .Z(SUM[35]) );
  CEOX1 U94 ( .A(A[34]), .B(n61), .Z(SUM[34]) );
  CEOX1 U95 ( .A(A[33]), .B(n62), .Z(SUM[33]) );
  CEOX1 U96 ( .A(A[32]), .B(n3), .Z(SUM[32]) );
  CEOX1 U97 ( .A(A[30]), .B(n63), .Z(SUM[30]) );
  CEOX1 U98 ( .A(A[29]), .B(n5), .Z(SUM[29]) );
  CEOX1 U99 ( .A(A[31]), .B(n4), .Z(SUM[31]) );
  CEOX1 U100 ( .A(A[28]), .B(n6), .Z(SUM[28]) );
  CEOX1 U101 ( .A(A[26]), .B(n8), .Z(SUM[26]) );
  CEOX1 U102 ( .A(A[25]), .B(n9), .Z(SUM[25]) );
  CEOX1 U103 ( .A(A[27]), .B(n7), .Z(SUM[27]) );
  CEOX1 U104 ( .A(A[22]), .B(n12), .Z(SUM[22]) );
  CEOX1 U105 ( .A(A[21]), .B(n13), .Z(SUM[21]) );
  CEOX1 U106 ( .A(A[24]), .B(n10), .Z(SUM[24]) );
  CEOX1 U107 ( .A(A[23]), .B(n11), .Z(SUM[23]) );
  CEOX1 U108 ( .A(A[18]), .B(n16), .Z(SUM[18]) );
  CEOX1 U109 ( .A(A[20]), .B(n14), .Z(SUM[20]) );
  CEOX1 U110 ( .A(A[19]), .B(n15), .Z(SUM[19]) );
  CEOX1 U111 ( .A(A[17]), .B(n17), .Z(SUM[17]) );
  CEOX1 U112 ( .A(A[14]), .B(n20), .Z(SUM[14]) );
  CEOX1 U113 ( .A(A[16]), .B(n18), .Z(SUM[16]) );
  CEOX1 U114 ( .A(A[15]), .B(n19), .Z(SUM[15]) );
  CEOX1 U115 ( .A(A[13]), .B(n21), .Z(SUM[13]) );
  CEOX1 U116 ( .A(A[12]), .B(n22), .Z(SUM[12]) );
  CEOX1 U117 ( .A(A[11]), .B(n23), .Z(SUM[11]) );
  CEOX1 U118 ( .A(A[10]), .B(n24), .Z(SUM[10]) );
  CEOX1 U119 ( .A(A[9]), .B(n25), .Z(SUM[9]) );
  CEOX1 U120 ( .A(A[8]), .B(n26), .Z(SUM[8]) );
  CEOX1 U121 ( .A(A[7]), .B(n27), .Z(SUM[7]) );
  CEOX1 U122 ( .A(A[5]), .B(n29), .Z(SUM[5]) );
  CEOX1 U123 ( .A(A[6]), .B(n28), .Z(SUM[6]) );
  CEOX1 U124 ( .A(A[4]), .B(n30), .Z(SUM[4]) );
  CEOX1 U125 ( .A(A[3]), .B(n31), .Z(SUM[3]) );
  CEOX1 U126 ( .A(A[2]), .B(n32), .Z(SUM[2]) );
  CEOX1 U127 ( .A(A[1]), .B(n33), .Z(SUM[1]) );
endmodule


module sfilt_DW01_add_1 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [63:1] carry;

  CFA1X1 U1_63 ( .A(A[63]), .B(B[63]), .CI(carry[63]), .S(SUM[63]) );
  CFA1X1 U1_62 ( .A(A[62]), .B(B[62]), .CI(carry[62]), .CO(carry[63]), .S(
        SUM[62]) );
  CFA1X1 U1_61 ( .A(A[61]), .B(B[61]), .CI(carry[61]), .CO(carry[62]), .S(
        SUM[61]) );
  CFA1X1 U1_60 ( .A(A[60]), .B(B[60]), .CI(carry[60]), .CO(carry[61]), .S(
        SUM[60]) );
  CFA1X1 U1_59 ( .A(A[59]), .B(B[59]), .CI(carry[59]), .CO(carry[60]), .S(
        SUM[59]) );
  CFA1X1 U1_58 ( .A(A[58]), .B(B[58]), .CI(carry[58]), .CO(carry[59]), .S(
        SUM[58]) );
  CFA1X1 U1_57 ( .A(A[57]), .B(B[57]), .CI(carry[57]), .CO(carry[58]), .S(
        SUM[57]) );
  CFA1X1 U1_56 ( .A(A[56]), .B(B[56]), .CI(carry[56]), .CO(carry[57]), .S(
        SUM[56]) );
  CFA1X1 U1_55 ( .A(A[55]), .B(B[55]), .CI(carry[55]), .CO(carry[56]), .S(
        SUM[55]) );
  CFA1X1 U1_54 ( .A(A[54]), .B(B[54]), .CI(carry[54]), .CO(carry[55]), .S(
        SUM[54]) );
  CFA1X1 U1_53 ( .A(A[53]), .B(B[53]), .CI(carry[53]), .CO(carry[54]), .S(
        SUM[53]) );
  CFA1X1 U1_52 ( .A(A[52]), .B(B[52]), .CI(carry[52]), .CO(carry[53]), .S(
        SUM[52]) );
  CFA1X1 U1_51 ( .A(A[51]), .B(B[51]), .CI(carry[51]), .CO(carry[52]), .S(
        SUM[51]) );
  CFA1X1 U1_50 ( .A(A[50]), .B(B[50]), .CI(carry[50]), .CO(carry[51]), .S(
        SUM[50]) );
  CFA1X1 U1_49 ( .A(A[49]), .B(B[49]), .CI(carry[49]), .CO(carry[50]), .S(
        SUM[49]) );
  CFA1X1 U1_48 ( .A(A[48]), .B(B[48]), .CI(carry[48]), .CO(carry[49]), .S(
        SUM[48]) );
  CFA1X1 U1_47 ( .A(A[47]), .B(B[47]), .CI(carry[47]), .CO(carry[48]), .S(
        SUM[47]) );
  CFA1X1 U1_46 ( .A(A[46]), .B(B[46]), .CI(carry[46]), .CO(carry[47]), .S(
        SUM[46]) );
  CFA1X1 U1_45 ( .A(A[45]), .B(B[45]), .CI(carry[45]), .CO(carry[46]), .S(
        SUM[45]) );
  CFA1X1 U1_44 ( .A(A[44]), .B(B[44]), .CI(carry[44]), .CO(carry[45]), .S(
        SUM[44]) );
  CFA1X1 U1_43 ( .A(A[43]), .B(B[43]), .CI(carry[43]), .CO(carry[44]), .S(
        SUM[43]) );
  CFA1X1 U1_42 ( .A(A[42]), .B(B[42]), .CI(carry[42]), .CO(carry[43]), .S(
        SUM[42]) );
  CFA1X1 U1_41 ( .A(A[41]), .B(B[41]), .CI(carry[41]), .CO(carry[42]), .S(
        SUM[41]) );
  CFA1X1 U1_40 ( .A(A[40]), .B(B[40]), .CI(carry[40]), .CO(carry[41]), .S(
        SUM[40]) );
  CFA1X1 U1_39 ( .A(A[39]), .B(B[39]), .CI(carry[39]), .CO(carry[40]), .S(
        SUM[39]) );
  CFA1X1 U1_38 ( .A(A[38]), .B(B[38]), .CI(carry[38]), .CO(carry[39]), .S(
        SUM[38]) );
  CFA1X1 U1_37 ( .A(A[37]), .B(B[37]), .CI(carry[37]), .CO(carry[38]), .S(
        SUM[37]) );
  CFA1X1 U1_36 ( .A(A[36]), .B(B[36]), .CI(carry[36]), .CO(carry[37]), .S(
        SUM[36]) );
  CFA1X1 U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  CFA1X1 U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  CFA1X1 U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  CFA1X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  CFA1X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  CFA1X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  CFA1X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  CFA1X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  CFA1X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  CFA1X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  CFA1X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  CFA1X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  CFA1X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  CFA1X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  CFA1X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  CFA1X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  CFA1X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  CFA1X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  CFA1X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  CFA1X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  CFA1X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  CFA1X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  CFA1X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  CFA1X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  CFA1X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  CFA1X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  CFA1X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  CFA1X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  CFA1X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  CFA1X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  CFA1X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  CFA1X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  CFA1X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  CFA1X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  CFA1X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  CAN2X1 U1 ( .A(B[0]), .B(A[0]), .Z(n1) );
  CEOX1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module sfilt_DW_mult_tc_0 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n212, n213, n214,
         n215, n216, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089;

  CFA1X1 U149 ( .A(n210), .B(n149), .CI(n1156), .CO(n148), .S(product[62]) );
  CFA1X1 U150 ( .A(n2460), .B(n150), .CI(n212), .CO(n149), .S(product[61]) );
  CFA1X1 U151 ( .A(n213), .B(n151), .CI(n214), .CO(n150), .S(product[60]) );
  CFA1X1 U152 ( .A(n218), .B(n152), .CI(n215), .CO(n151), .S(product[59]) );
  CFA1X1 U153 ( .A(n219), .B(n153), .CI(n222), .CO(n152), .S(product[58]) );
  CFA1X1 U154 ( .A(n228), .B(n154), .CI(n223), .CO(n153), .S(product[57]) );
  CFA1X1 U155 ( .A(n234), .B(n155), .CI(n229), .CO(n154), .S(product[56]) );
  CFA1X1 U156 ( .A(n235), .B(n156), .CI(n242), .CO(n155), .S(product[55]) );
  CFA1X1 U157 ( .A(n250), .B(n157), .CI(n243), .CO(n156), .S(product[54]) );
  CFA1X1 U158 ( .A(n260), .B(n158), .CI(n251), .CO(n157), .S(product[53]) );
  CFA1X1 U159 ( .A(n270), .B(n159), .CI(n261), .CO(n158), .S(product[52]) );
  CFA1X1 U160 ( .A(n282), .B(n160), .CI(n271), .CO(n159), .S(product[51]) );
  CFA1X1 U161 ( .A(n283), .B(n161), .CI(n294), .CO(n160), .S(product[50]) );
  CFA1X1 U162 ( .A(n308), .B(n162), .CI(n295), .CO(n161), .S(product[49]) );
  CFA1X1 U163 ( .A(n322), .B(n163), .CI(n309), .CO(n162), .S(product[48]) );
  CFA1X1 U164 ( .A(n338), .B(n164), .CI(n323), .CO(n163), .S(product[47]) );
  CFA1X1 U165 ( .A(n354), .B(n165), .CI(n339), .CO(n164), .S(product[46]) );
  CFA1X1 U166 ( .A(n372), .B(n166), .CI(n355), .CO(n165), .S(product[45]) );
  CFA1X1 U167 ( .A(n390), .B(n167), .CI(n373), .CO(n166), .S(product[44]) );
  CFA1X1 U168 ( .A(n410), .B(n168), .CI(n391), .CO(n167), .S(product[43]) );
  CFA1X1 U169 ( .A(n430), .B(n169), .CI(n411), .CO(n168), .S(product[42]) );
  CFA1X1 U170 ( .A(n452), .B(n170), .CI(n431), .CO(n169), .S(product[41]) );
  CFA1X1 U171 ( .A(n474), .B(n171), .CI(n453), .CO(n170), .S(product[40]) );
  CFA1X1 U172 ( .A(n498), .B(n172), .CI(n475), .CO(n171), .S(product[39]) );
  CFA1X1 U173 ( .A(n522), .B(n173), .CI(n499), .CO(n172), .S(product[38]) );
  CFA1X1 U174 ( .A(n548), .B(n174), .CI(n523), .CO(n173), .S(product[37]) );
  CFA1X1 U175 ( .A(n574), .B(n175), .CI(n549), .CO(n174), .S(product[36]) );
  CFA1X1 U176 ( .A(n602), .B(n176), .CI(n575), .CO(n175), .S(product[35]) );
  CFA1X1 U177 ( .A(n630), .B(n177), .CI(n603), .CO(n176), .S(product[34]) );
  CFA1X1 U178 ( .A(n660), .B(n178), .CI(n631), .CO(n177), .S(product[33]) );
  CFA1X1 U179 ( .A(n690), .B(n179), .CI(n661), .CO(n178), .S(product[32]) );
  CFA1X1 U180 ( .A(n720), .B(n180), .CI(n691), .CO(n179), .S(product[31]) );
  CFA1X1 U181 ( .A(n748), .B(n181), .CI(n721), .CO(n180), .S(product[30]) );
  CFA1X1 U182 ( .A(n776), .B(n182), .CI(n749), .CO(n181), .S(product[29]) );
  CFA1X1 U183 ( .A(n802), .B(n183), .CI(n777), .CO(n182), .S(product[28]) );
  CFA1X1 U184 ( .A(n828), .B(n184), .CI(n803), .CO(n183), .S(product[27]) );
  CFA1X1 U185 ( .A(n852), .B(n185), .CI(n829), .CO(n184), .S(product[26]) );
  CFA1X1 U186 ( .A(n876), .B(n186), .CI(n853), .CO(n185), .S(product[25]) );
  CFA1X1 U187 ( .A(n898), .B(n187), .CI(n877), .CO(n186), .S(product[24]) );
  CFA1X1 U188 ( .A(n920), .B(n188), .CI(n899), .CO(n187), .S(product[23]) );
  CFA1X1 U189 ( .A(n940), .B(n189), .CI(n921), .CO(n188), .S(product[22]) );
  CFA1X1 U190 ( .A(n960), .B(n190), .CI(n941), .CO(n189), .S(product[21]) );
  CFA1X1 U191 ( .A(n978), .B(n191), .CI(n961), .CO(n190), .S(product[20]) );
  CFA1X1 U192 ( .A(n996), .B(n192), .CI(n979), .CO(n191), .S(product[19]) );
  CFA1X1 U193 ( .A(n1012), .B(n193), .CI(n997), .CO(n192), .S(product[18]) );
  CFA1X1 U194 ( .A(n1028), .B(n194), .CI(n1013), .CO(n193), .S(product[17]) );
  CFA1X1 U195 ( .A(n1042), .B(n195), .CI(n1029), .CO(n194), .S(product[16]) );
  CFA1X1 U196 ( .A(n1056), .B(n196), .CI(n1043), .CO(n195), .S(product[15]) );
  CFA1X1 U197 ( .A(n1068), .B(n197), .CI(n1057), .CO(n196), .S(product[14]) );
  CFA1X1 U198 ( .A(n1080), .B(n198), .CI(n1069), .CO(n197), .S(product[13]) );
  CFA1X1 U199 ( .A(n1090), .B(n199), .CI(n1081), .CO(n198), .S(product[12]) );
  CFA1X1 U200 ( .A(n1100), .B(n200), .CI(n1091), .CO(n199), .S(product[11]) );
  CFA1X1 U201 ( .A(n1108), .B(n201), .CI(n1101), .CO(n200), .S(product[10]) );
  CFA1X1 U202 ( .A(n1116), .B(n202), .CI(n1109), .CO(n201), .S(product[9]) );
  CFA1X1 U203 ( .A(n1122), .B(n203), .CI(n1117), .CO(n202), .S(product[8]) );
  CFA1X1 U204 ( .A(n1128), .B(n204), .CI(n1123), .CO(n203), .S(product[7]) );
  CFA1X1 U205 ( .A(n1132), .B(n205), .CI(n1129), .CO(n204), .S(product[6]) );
  CFA1X1 U206 ( .A(n1136), .B(n206), .CI(n1133), .CO(n205), .S(product[5]) );
  CFA1X1 U207 ( .A(n1138), .B(n207), .CI(n1137), .CO(n206), .S(product[4]) );
  CFA1X1 U208 ( .A(n1154), .B(n208), .CI(n1139), .CO(n207), .S(product[3]) );
  CFA1X1 U209 ( .A(n1635), .B(n209), .CI(n1666), .CO(n208), .S(product[2]) );
  CHA1X1 U210 ( .A(n1155), .B(n1667), .CO(n209), .S(product[1]) );
  CFA1X1 U212 ( .A(n216), .B(n1188), .CI(n1157), .CO(n212), .S(n213) );
  CFA1X1 U213 ( .A(n1158), .B(n220), .CI(n2462), .CO(n214), .S(n215) );
  CFA1X1 U215 ( .A(n1159), .B(n221), .CI(n224), .CO(n218), .S(n219) );
  CFA1X1 U216 ( .A(n226), .B(n1220), .CI(n1189), .CO(n220), .S(n221) );
  CFA1X1 U217 ( .A(n232), .B(n230), .CI(n225), .CO(n222), .S(n223) );
  CFA1X1 U218 ( .A(n1190), .B(n2464), .CI(n1160), .CO(n224), .S(n225) );
  CFA1X1 U220 ( .A(n233), .B(n231), .CI(n236), .CO(n228), .S(n229) );
  CFA1X1 U221 ( .A(n1221), .B(n238), .CI(n240), .CO(n230), .S(n231) );
  CFA1X1 U222 ( .A(n1161), .B(n1252), .CI(n1191), .CO(n232), .S(n233) );
  CFA1X1 U223 ( .A(n239), .B(n244), .CI(n237), .CO(n234), .S(n235) );
  CFA1X1 U224 ( .A(n2466), .B(n246), .CI(n248), .CO(n236), .S(n237) );
  CFA1X1 U225 ( .A(n1192), .B(n1222), .CI(n1162), .CO(n238), .S(n239) );
  CFA1X1 U227 ( .A(n254), .B(n252), .CI(n245), .CO(n242), .S(n243) );
  CFA1X1 U228 ( .A(n256), .B(n249), .CI(n247), .CO(n244), .S(n245) );
  CFA1X1 U229 ( .A(n258), .B(n1223), .CI(n1193), .CO(n246), .S(n247) );
  CFA1X1 U230 ( .A(n1163), .B(n1284), .CI(n1253), .CO(n248), .S(n249) );
  CFA1X1 U231 ( .A(n255), .B(n253), .CI(n262), .CO(n250), .S(n251) );
  CFA1X1 U232 ( .A(n266), .B(n264), .CI(n257), .CO(n252), .S(n253) );
  CFA1X1 U233 ( .A(n1224), .B(n268), .CI(n2468), .CO(n254), .S(n255) );
  CFA1X1 U234 ( .A(n1194), .B(n1164), .CI(n1254), .CO(n256), .S(n257) );
  CFA1X1 U236 ( .A(n265), .B(n263), .CI(n272), .CO(n260), .S(n261) );
  CFA1X1 U237 ( .A(n267), .B(n274), .CI(n269), .CO(n262), .S(n263) );
  CFA1X1 U238 ( .A(n1255), .B(n276), .CI(n278), .CO(n264), .S(n265) );
  CFA1X1 U239 ( .A(n1285), .B(n1225), .CI(n1195), .CO(n266), .S(n267) );
  CFA1X1 U240 ( .A(n1165), .B(n1316), .CI(n280), .CO(n268), .S(n269) );
  CFA1X1 U241 ( .A(n275), .B(n273), .CI(n284), .CO(n270), .S(n271) );
  CFA1X1 U242 ( .A(n277), .B(n286), .CI(n288), .CO(n272), .S(n273) );
  CFA1X1 U243 ( .A(n292), .B(n279), .CI(n290), .CO(n274), .S(n275) );
  CFA1X1 U244 ( .A(n1196), .B(n2470), .CI(n1166), .CO(n276), .S(n277) );
  CFA1X1 U245 ( .A(n1226), .B(n1256), .CI(n1286), .CO(n278), .S(n279) );
  CFA1X1 U247 ( .A(n287), .B(n285), .CI(n296), .CO(n282), .S(n283) );
  CFA1X1 U248 ( .A(n300), .B(n298), .CI(n289), .CO(n284), .S(n285) );
  CFA1X1 U249 ( .A(n302), .B(n293), .CI(n291), .CO(n286), .S(n287) );
  CFA1X1 U250 ( .A(n1257), .B(n304), .CI(n1227), .CO(n288), .S(n289) );
  CFA1X1 U251 ( .A(n1317), .B(n1287), .CI(n1197), .CO(n290), .S(n291) );
  CFA1X1 U252 ( .A(n1167), .B(n1348), .CI(n306), .CO(n292), .S(n293) );
  CFA1X1 U253 ( .A(n299), .B(n297), .CI(n310), .CO(n294), .S(n295) );
  CFA1X1 U254 ( .A(n314), .B(n312), .CI(n301), .CO(n296), .S(n297) );
  CFA1X1 U255 ( .A(n316), .B(n305), .CI(n303), .CO(n298), .S(n299) );
  CFA1X1 U256 ( .A(n2472), .B(n318), .CI(n320), .CO(n300), .S(n301) );
  CFA1X1 U257 ( .A(n1318), .B(n1288), .CI(n1258), .CO(n302), .S(n303) );
  CFA1X1 U258 ( .A(n1228), .B(n1198), .CI(n1168), .CO(n304), .S(n305) );
  CFA1X1 U260 ( .A(n313), .B(n311), .CI(n324), .CO(n308), .S(n309) );
  CFA1X1 U261 ( .A(n328), .B(n326), .CI(n315), .CO(n310), .S(n311) );
  CFA1X1 U262 ( .A(n319), .B(n330), .CI(n321), .CO(n312), .S(n313) );
  CFA1X1 U263 ( .A(n334), .B(n317), .CI(n332), .CO(n314), .S(n315) );
  CFA1X1 U264 ( .A(n1289), .B(n1259), .CI(n1229), .CO(n316), .S(n317) );
  CFA1X1 U265 ( .A(n1349), .B(n1319), .CI(n1199), .CO(n318), .S(n319) );
  CFA1X1 U266 ( .A(n1169), .B(n1380), .CI(n336), .CO(n320), .S(n321) );
  CFA1X1 U267 ( .A(n327), .B(n325), .CI(n340), .CO(n322), .S(n323) );
  CFA1X1 U268 ( .A(n344), .B(n342), .CI(n329), .CO(n324), .S(n325) );
  CFA1X1 U269 ( .A(n335), .B(n331), .CI(n346), .CO(n326), .S(n327) );
  CFA1X1 U270 ( .A(n350), .B(n333), .CI(n348), .CO(n328), .S(n329) );
  CFA1X1 U271 ( .A(n1260), .B(n352), .CI(n2474), .CO(n330), .S(n331) );
  CFA1X1 U272 ( .A(n1290), .B(n1200), .CI(n1170), .CO(n332), .S(n333) );
  CFA1X1 U273 ( .A(n1230), .B(n1320), .CI(n1350), .CO(n334), .S(n335) );
  CFA1X1 U275 ( .A(n343), .B(n341), .CI(n356), .CO(n338), .S(n339) );
  CFA1X1 U276 ( .A(n360), .B(n358), .CI(n345), .CO(n340), .S(n341) );
  CFA1X1 U277 ( .A(n353), .B(n347), .CI(n362), .CO(n342), .S(n343) );
  CFA1X1 U278 ( .A(n364), .B(n351), .CI(n349), .CO(n344), .S(n345) );
  CFA1X1 U279 ( .A(n1291), .B(n366), .CI(n368), .CO(n346), .S(n347) );
  CFA1X1 U280 ( .A(n1321), .B(n1261), .CI(n1231), .CO(n348), .S(n349) );
  CFA1X1 U281 ( .A(n1351), .B(n1201), .CI(n370), .CO(n350), .S(n351) );
  CFA1X1 U282 ( .A(n1171), .B(n1412), .CI(n1381), .CO(n352), .S(n353) );
  CFA1X1 U283 ( .A(n359), .B(n357), .CI(n374), .CO(n354), .S(n355) );
  CFA1X1 U284 ( .A(n361), .B(n376), .CI(n378), .CO(n356), .S(n357) );
  CFA1X1 U285 ( .A(n382), .B(n363), .CI(n380), .CO(n358), .S(n359) );
  CFA1X1 U286 ( .A(n367), .B(n365), .CI(n369), .CO(n360), .S(n361) );
  CFA1X1 U287 ( .A(n388), .B(n386), .CI(n384), .CO(n362), .S(n363) );
  CFA1X1 U288 ( .A(n1382), .B(n2476), .CI(n1352), .CO(n364), .S(n365) );
  CFA1X1 U289 ( .A(n1232), .B(n1322), .CI(n1292), .CO(n366), .S(n367) );
  CFA1X1 U290 ( .A(n1262), .B(n1202), .CI(n1172), .CO(n368), .S(n369) );
  CFA1X1 U292 ( .A(n377), .B(n375), .CI(n392), .CO(n372), .S(n373) );
  CFA1X1 U293 ( .A(n396), .B(n394), .CI(n379), .CO(n374), .S(n375) );
  CFA1X1 U294 ( .A(n398), .B(n381), .CI(n383), .CO(n376), .S(n377) );
  CFA1X1 U295 ( .A(n387), .B(n400), .CI(n389), .CO(n378), .S(n379) );
  CFA1X1 U296 ( .A(n404), .B(n385), .CI(n402), .CO(n380), .S(n381) );
  CFA1X1 U297 ( .A(n1353), .B(n406), .CI(n1323), .CO(n382), .S(n383) );
  CFA1X1 U298 ( .A(n1233), .B(n1293), .CI(n1263), .CO(n384), .S(n385) );
  CFA1X1 U299 ( .A(n1383), .B(n1203), .CI(n408), .CO(n386), .S(n387) );
  CFA1X1 U300 ( .A(n1173), .B(n1444), .CI(n1413), .CO(n388), .S(n389) );
  CFA1X1 U301 ( .A(n395), .B(n393), .CI(n412), .CO(n390), .S(n391) );
  CFA1X1 U302 ( .A(n416), .B(n414), .CI(n397), .CO(n392), .S(n393) );
  CFA1X1 U303 ( .A(n401), .B(n399), .CI(n418), .CO(n394), .S(n395) );
  CFA1X1 U304 ( .A(n405), .B(n420), .CI(n407), .CO(n396), .S(n397) );
  CFA1X1 U305 ( .A(n424), .B(n403), .CI(n422), .CO(n398), .S(n399) );
  CFA1X1 U306 ( .A(n2478), .B(n426), .CI(n428), .CO(n400), .S(n401) );
  CFA1X1 U307 ( .A(n1354), .B(n1324), .CI(n1234), .CO(n402), .S(n403) );
  CFA1X1 U308 ( .A(n1294), .B(n1204), .CI(n1384), .CO(n404), .S(n405) );
  CFA1X1 U309 ( .A(n1264), .B(n1414), .CI(n1174), .CO(n406), .S(n407) );
  CFA1X1 U311 ( .A(n415), .B(n413), .CI(n432), .CO(n410), .S(n411) );
  CFA1X1 U312 ( .A(n436), .B(n434), .CI(n417), .CO(n412), .S(n413) );
  CFA1X1 U313 ( .A(n438), .B(n419), .CI(n421), .CO(n414), .S(n415) );
  CFA1X1 U314 ( .A(n425), .B(n440), .CI(n442), .CO(n416), .S(n417) );
  CFA1X1 U315 ( .A(n423), .B(n427), .CI(n429), .CO(n418), .S(n419) );
  CFA1X1 U316 ( .A(n448), .B(n446), .CI(n444), .CO(n420), .S(n421) );
  CFA1X1 U317 ( .A(n1355), .B(n1325), .CI(n1295), .CO(n422), .S(n423) );
  CFA1X1 U318 ( .A(n1235), .B(n1265), .CI(n1385), .CO(n424), .S(n425) );
  CFA1X1 U319 ( .A(n1415), .B(n1205), .CI(n450), .CO(n426), .S(n427) );
  CFA1X1 U320 ( .A(n1175), .B(n1476), .CI(n1445), .CO(n428), .S(n429) );
  CFA1X1 U321 ( .A(n435), .B(n433), .CI(n454), .CO(n430), .S(n431) );
  CFA1X1 U322 ( .A(n458), .B(n456), .CI(n437), .CO(n432), .S(n433) );
  CFA1X1 U323 ( .A(n460), .B(n439), .CI(n441), .CO(n434), .S(n435) );
  CFA1X1 U324 ( .A(n464), .B(n443), .CI(n462), .CO(n436), .S(n437) );
  CFA1X1 U325 ( .A(n445), .B(n447), .CI(n449), .CO(n438), .S(n439) );
  CFA1X1 U326 ( .A(n470), .B(n468), .CI(n466), .CO(n440), .S(n441) );
  CFA1X1 U327 ( .A(n1356), .B(n472), .CI(n2480), .CO(n442), .S(n443) );
  CFA1X1 U328 ( .A(n1386), .B(n1326), .CI(n1236), .CO(n444), .S(n445) );
  CFA1X1 U329 ( .A(n1266), .B(n1416), .CI(n1206), .CO(n446), .S(n447) );
  CFA1X1 U330 ( .A(n1296), .B(n1446), .CI(n1176), .CO(n448), .S(n449) );
  CFA1X1 U332 ( .A(n457), .B(n455), .CI(n476), .CO(n452), .S(n453) );
  CFA1X1 U333 ( .A(n480), .B(n478), .CI(n459), .CO(n454), .S(n455) );
  CFA1X1 U334 ( .A(n463), .B(n461), .CI(n482), .CO(n456), .S(n457) );
  CFA1X1 U335 ( .A(n486), .B(n484), .CI(n465), .CO(n458), .S(n459) );
  CFA1X1 U336 ( .A(n469), .B(n471), .CI(n473), .CO(n460), .S(n461) );
  CFA1X1 U337 ( .A(n490), .B(n467), .CI(n488), .CO(n462), .S(n463) );
  CFA1X1 U338 ( .A(n1357), .B(n492), .CI(n494), .CO(n464), .S(n465) );
  CFA1X1 U339 ( .A(n1387), .B(n1327), .CI(n1297), .CO(n466), .S(n467) );
  CFA1X1 U340 ( .A(n1447), .B(n1417), .CI(n1267), .CO(n468), .S(n469) );
  CFA1X1 U341 ( .A(n1477), .B(n1237), .CI(n1207), .CO(n470), .S(n471) );
  CFA1X1 U342 ( .A(n1177), .B(n1508), .CI(n496), .CO(n472), .S(n473) );
  CFA1X1 U343 ( .A(n479), .B(n477), .CI(n500), .CO(n474), .S(n475) );
  CFA1X1 U344 ( .A(n504), .B(n502), .CI(n481), .CO(n476), .S(n477) );
  CFA1X1 U345 ( .A(n485), .B(n483), .CI(n506), .CO(n478), .S(n479) );
  CFA1X1 U346 ( .A(n510), .B(n487), .CI(n508), .CO(n480), .S(n481) );
  CFA1X1 U347 ( .A(n495), .B(n512), .CI(n489), .CO(n482), .S(n483) );
  CFA1X1 U348 ( .A(n518), .B(n493), .CI(n491), .CO(n484), .S(n485) );
  CFA1X1 U349 ( .A(n520), .B(n516), .CI(n514), .CO(n486), .S(n487) );
  CFA1X1 U350 ( .A(n1388), .B(n2482), .CI(n1298), .CO(n488), .S(n489) );
  CFA1X1 U351 ( .A(n1418), .B(n1268), .CI(n1238), .CO(n490), .S(n491) );
  CFA1X1 U352 ( .A(n1358), .B(n1448), .CI(n1478), .CO(n492), .S(n493) );
  CFA1X1 U353 ( .A(n1328), .B(n1208), .CI(n1178), .CO(n494), .S(n495) );
  CFA1X1 U355 ( .A(n503), .B(n501), .CI(n524), .CO(n498), .S(n499) );
  CFA1X1 U356 ( .A(n528), .B(n526), .CI(n505), .CO(n500), .S(n501) );
  CFA1X1 U357 ( .A(n509), .B(n507), .CI(n530), .CO(n502), .S(n503) );
  CFA1X1 U358 ( .A(n513), .B(n511), .CI(n532), .CO(n504), .S(n505) );
  CFA1X1 U359 ( .A(n517), .B(n534), .CI(n536), .CO(n506), .S(n507) );
  CFA1X1 U360 ( .A(n515), .B(n519), .CI(n521), .CO(n508), .S(n509) );
  CFA1X1 U361 ( .A(n538), .B(n542), .CI(n540), .CO(n510), .S(n511) );
  CFA1X1 U362 ( .A(n1389), .B(n544), .CI(n1359), .CO(n512), .S(n513) );
  CFA1X1 U363 ( .A(n1419), .B(n1299), .CI(n1269), .CO(n514), .S(n515) );
  CFA1X1 U364 ( .A(n1479), .B(n1449), .CI(n1239), .CO(n516), .S(n517) );
  CFA1X1 U365 ( .A(n1329), .B(n1209), .CI(n546), .CO(n518), .S(n519) );
  CFA1X1 U366 ( .A(n1179), .B(n1540), .CI(n1509), .CO(n520), .S(n521) );
  CFA1X1 U367 ( .A(n527), .B(n525), .CI(n550), .CO(n522), .S(n523) );
  CFA1X1 U368 ( .A(n554), .B(n552), .CI(n529), .CO(n524), .S(n525) );
  CFA1X1 U369 ( .A(n533), .B(n531), .CI(n556), .CO(n526), .S(n527) );
  CFA1X1 U370 ( .A(n560), .B(n535), .CI(n558), .CO(n528), .S(n529) );
  CFA1X1 U371 ( .A(n541), .B(n537), .CI(n562), .CO(n530), .S(n531) );
  CFA1X1 U372 ( .A(n539), .B(n543), .CI(n545), .CO(n532), .S(n533) );
  CFA1X1 U373 ( .A(n564), .B(n568), .CI(n566), .CO(n534), .S(n535) );
  CFA1X1 U374 ( .A(n2484), .B(n570), .CI(n572), .CO(n536), .S(n537) );
  CFA1X1 U375 ( .A(n1360), .B(n1300), .CI(n1240), .CO(n538), .S(n539) );
  CFA1X1 U376 ( .A(n1390), .B(n1210), .CI(n1180), .CO(n540), .S(n541) );
  CFA1X1 U377 ( .A(n1270), .B(n1420), .CI(n1450), .CO(n542), .S(n543) );
  CFA1X1 U378 ( .A(n1330), .B(n1480), .CI(n1510), .CO(n544), .S(n545) );
  CFA1X1 U380 ( .A(n553), .B(n551), .CI(n576), .CO(n548), .S(n549) );
  CFA1X1 U381 ( .A(n580), .B(n578), .CI(n555), .CO(n550), .S(n551) );
  CFA1X1 U382 ( .A(n584), .B(n557), .CI(n582), .CO(n552), .S(n553) );
  CFA1X1 U383 ( .A(n563), .B(n559), .CI(n561), .CO(n554), .S(n555) );
  CFA1X1 U384 ( .A(n590), .B(n586), .CI(n588), .CO(n556), .S(n557) );
  CFA1X1 U385 ( .A(n571), .B(n573), .CI(n569), .CO(n558), .S(n559) );
  CFA1X1 U386 ( .A(n594), .B(n567), .CI(n565), .CO(n560), .S(n561) );
  CFA1X1 U387 ( .A(n598), .B(n596), .CI(n592), .CO(n562), .S(n563) );
  CFA1X1 U388 ( .A(n1421), .B(n1391), .CI(n1331), .CO(n564), .S(n565) );
  CFA1X1 U389 ( .A(n1451), .B(n1301), .CI(n1271), .CO(n566), .S(n567) );
  CFA1X1 U390 ( .A(n1481), .B(n1241), .CI(n1211), .CO(n568), .S(n569) );
  CFA1X1 U391 ( .A(n1361), .B(n600), .CI(n1511), .CO(n570), .S(n571) );
  CFA1X1 U392 ( .A(n1181), .B(n1572), .CI(n1541), .CO(n572), .S(n573) );
  CFA1X1 U393 ( .A(n579), .B(n577), .CI(n604), .CO(n574), .S(n575) );
  CFA1X1 U394 ( .A(n608), .B(n606), .CI(n581), .CO(n576), .S(n577) );
  CFA1X1 U395 ( .A(n585), .B(n583), .CI(n610), .CO(n578), .S(n579) );
  CFA1X1 U396 ( .A(n589), .B(n612), .CI(n587), .CO(n580), .S(n581) );
  CFA1X1 U397 ( .A(n616), .B(n614), .CI(n591), .CO(n582), .S(n583) );
  CFA1X1 U398 ( .A(n597), .B(n618), .CI(n599), .CO(n584), .S(n585) );
  CFA1X1 U399 ( .A(n624), .B(n595), .CI(n593), .CO(n586), .S(n587) );
  CFA1X1 U400 ( .A(n622), .B(n620), .CI(n626), .CO(n588), .S(n589) );
  CFA1X1 U401 ( .A(n1482), .B(n628), .CI(n2486), .CO(n590), .S(n591) );
  CFA1X1 U402 ( .A(n1512), .B(n1452), .CI(n1422), .CO(n592), .S(n593) );
  CFA1X1 U403 ( .A(n1272), .B(n1392), .CI(n1302), .CO(n594), .S(n595) );
  CFA1X1 U404 ( .A(n1332), .B(n1242), .CI(n1212), .CO(n596), .S(n597) );
  CFA1X1 U405 ( .A(n1362), .B(n1542), .CI(n1182), .CO(n598), .S(n599) );
  CFA1X1 U407 ( .A(n607), .B(n605), .CI(n632), .CO(n602), .S(n603) );
  CFA1X1 U408 ( .A(n636), .B(n634), .CI(n609), .CO(n604), .S(n605) );
  CFA1X1 U409 ( .A(n613), .B(n611), .CI(n638), .CO(n606), .S(n607) );
  CFA1X1 U410 ( .A(n617), .B(n640), .CI(n615), .CO(n608), .S(n609) );
  CFA1X1 U411 ( .A(n644), .B(n642), .CI(n619), .CO(n610), .S(n611) );
  CFA1X1 U412 ( .A(n623), .B(n646), .CI(n625), .CO(n612), .S(n613) );
  CFA1X1 U413 ( .A(n621), .B(n627), .CI(n629), .CO(n614), .S(n615) );
  CFA1X1 U414 ( .A(n652), .B(n648), .CI(n650), .CO(n616), .S(n617) );
  CFA1X1 U415 ( .A(n1483), .B(n654), .CI(n656), .CO(n618), .S(n619) );
  CFA1X1 U416 ( .A(n1513), .B(n1453), .CI(n1423), .CO(n620), .S(n621) );
  CFA1X1 U417 ( .A(n1303), .B(n1363), .CI(n1333), .CO(n622), .S(n623) );
  CFA1X1 U418 ( .A(n1543), .B(n1273), .CI(n1243), .CO(n624), .S(n625) );
  CFA1X1 U419 ( .A(n1393), .B(n1213), .CI(n1573), .CO(n626), .S(n627) );
  CFA1X1 U420 ( .A(n1183), .B(n1604), .CI(n658), .CO(n628), .S(n629) );
  CFA1X1 U421 ( .A(n635), .B(n633), .CI(n662), .CO(n630), .S(n631) );
  CFA1X1 U422 ( .A(n666), .B(n664), .CI(n637), .CO(n632), .S(n633) );
  CFA1X1 U423 ( .A(n641), .B(n639), .CI(n668), .CO(n634), .S(n635) );
  CFA1X1 U424 ( .A(n645), .B(n643), .CI(n670), .CO(n636), .S(n637) );
  CFA1X1 U425 ( .A(n674), .B(n672), .CI(n647), .CO(n638), .S(n639) );
  CFA1X1 U426 ( .A(n651), .B(n676), .CI(n653), .CO(n640), .S(n641) );
  CFA1X1 U427 ( .A(n655), .B(n649), .CI(n657), .CO(n642), .S(n643) );
  CFA1X1 U428 ( .A(n684), .B(n678), .CI(n686), .CO(n644), .S(n645) );
  CFA1X1 U429 ( .A(n688), .B(n682), .CI(n680), .CO(n646), .S(n647) );
  CFA1X1 U430 ( .A(n1484), .B(n2488), .CI(n1514), .CO(n648), .S(n649) );
  CFA1X1 U431 ( .A(n1544), .B(n1454), .CI(n1424), .CO(n650), .S(n651) );
  CFA1X1 U432 ( .A(n1304), .B(n1334), .CI(n1274), .CO(n652), .S(n653) );
  CFA1X1 U433 ( .A(n1394), .B(n1244), .CI(n1574), .CO(n654), .S(n655) );
  CFA1X1 U434 ( .A(n1364), .B(n1214), .CI(n1184), .CO(n656), .S(n657) );
  CFA1X1 U436 ( .A(n665), .B(n663), .CI(n692), .CO(n660), .S(n661) );
  CFA1X1 U437 ( .A(n669), .B(n694), .CI(n667), .CO(n662), .S(n663) );
  CFA1X1 U438 ( .A(n671), .B(n696), .CI(n698), .CO(n664), .S(n665) );
  CFA1X1 U439 ( .A(n675), .B(n673), .CI(n700), .CO(n666), .S(n667) );
  CFA1X1 U440 ( .A(n704), .B(n702), .CI(n677), .CO(n668), .S(n669) );
  CFA1X1 U441 ( .A(n683), .B(n706), .CI(n679), .CO(n670), .S(n671) );
  CFA1X1 U442 ( .A(n685), .B(n681), .CI(n687), .CO(n672), .S(n673) );
  CFA1X1 U443 ( .A(n708), .B(n712), .CI(n714), .CO(n674), .S(n675) );
  CFA1X1 U444 ( .A(n689), .B(n716), .CI(n710), .CO(n676), .S(n677) );
  CFA1X1 U445 ( .A(n1515), .B(n718), .CI(n1545), .CO(n678), .S(n679) );
  CFA1X1 U446 ( .A(n1575), .B(n1485), .CI(n1425), .CO(n680), .S(n681) );
  CFA1X1 U447 ( .A(n1335), .B(n1305), .CI(n1275), .CO(n682), .S(n683) );
  CFA1X1 U448 ( .A(n1365), .B(n1245), .CI(n1605), .CO(n684), .S(n685) );
  CFA1X1 U449 ( .A(n1395), .B(n1636), .CI(n1185), .CO(n686), .S(n687) );
  CFA1X1 U452 ( .A(n695), .B(n693), .CI(n722), .CO(n690), .S(n691) );
  CFA1X1 U453 ( .A(n699), .B(n724), .CI(n697), .CO(n692), .S(n693) );
  CFA1X1 U454 ( .A(n701), .B(n726), .CI(n728), .CO(n694), .S(n695) );
  CFA1X1 U455 ( .A(n705), .B(n703), .CI(n730), .CO(n696), .S(n697) );
  CFA1X1 U456 ( .A(n734), .B(n732), .CI(n707), .CO(n698), .S(n699) );
  CFA1X1 U457 ( .A(n711), .B(n736), .CI(n713), .CO(n700), .S(n701) );
  CFA1X1 U458 ( .A(n709), .B(n715), .CI(n717), .CO(n702), .S(n703) );
  CFA1X1 U459 ( .A(n738), .B(n740), .CI(n742), .CO(n704), .S(n705) );
  CFA1X1 U460 ( .A(n719), .B(n744), .CI(n746), .CO(n706), .S(n707) );
  CFA1X1 U461 ( .A(n1336), .B(n1396), .CI(n1486), .CO(n708), .S(n709) );
  CFA1X1 U462 ( .A(n1516), .B(n1306), .CI(n1276), .CO(n710), .S(n711) );
  CFA1X1 U463 ( .A(n1366), .B(n1546), .CI(n1576), .CO(n712), .S(n713) );
  CFA1X1 U464 ( .A(n1456), .B(n1606), .CI(n1637), .CO(n714), .S(n715) );
  CFA1X1 U465 ( .A(n1426), .B(n1246), .CI(n1216), .CO(n716), .S(n717) );
  CHA1X1 U466 ( .A(n1186), .B(n1140), .CO(n718), .S(n719) );
  CFA1X1 U467 ( .A(n725), .B(n723), .CI(n750), .CO(n720), .S(n721) );
  CFA1X1 U468 ( .A(n729), .B(n752), .CI(n727), .CO(n722), .S(n723) );
  CFA1X1 U469 ( .A(n731), .B(n754), .CI(n756), .CO(n724), .S(n725) );
  CFA1X1 U470 ( .A(n758), .B(n733), .CI(n735), .CO(n726), .S(n727) );
  CFA1X1 U471 ( .A(n762), .B(n737), .CI(n760), .CO(n728), .S(n729) );
  CFA1X1 U472 ( .A(n743), .B(n764), .CI(n741), .CO(n730), .S(n731) );
  CFA1X1 U473 ( .A(n747), .B(n745), .CI(n739), .CO(n732), .S(n733) );
  CFA1X1 U474 ( .A(n768), .B(n770), .CI(n772), .CO(n734), .S(n735) );
  CFA1X1 U475 ( .A(n1487), .B(n766), .CI(n774), .CO(n736), .S(n737) );
  CFA1X1 U476 ( .A(n1517), .B(n1457), .CI(n1427), .CO(n738), .S(n739) );
  CFA1X1 U477 ( .A(n1337), .B(n1397), .CI(n1367), .CO(n740), .S(n741) );
  CFA1X1 U478 ( .A(n1547), .B(n1307), .CI(n1277), .CO(n742), .S(n743) );
  CFA1X1 U479 ( .A(n1607), .B(n1577), .CI(n1217), .CO(n744), .S(n745) );
  CFA1X1 U480 ( .A(n1187), .B(n1638), .CI(n1247), .CO(n746), .S(n747) );
  CFA1X1 U481 ( .A(n753), .B(n751), .CI(n778), .CO(n748), .S(n749) );
  CFA1X1 U482 ( .A(n757), .B(n780), .CI(n755), .CO(n750), .S(n751) );
  CFA1X1 U483 ( .A(n759), .B(n782), .CI(n784), .CO(n752), .S(n753) );
  CFA1X1 U484 ( .A(n763), .B(n761), .CI(n786), .CO(n754), .S(n755) );
  CFA1X1 U485 ( .A(n790), .B(n788), .CI(n765), .CO(n756), .S(n757) );
  CFA1X1 U486 ( .A(n771), .B(n773), .CI(n769), .CO(n758), .S(n759) );
  CFA1X1 U487 ( .A(n794), .B(n767), .CI(n792), .CO(n760), .S(n761) );
  CFA1X1 U488 ( .A(n800), .B(n796), .CI(n798), .CO(n762), .S(n763) );
  CFA1X1 U489 ( .A(n1428), .B(n775), .CI(n1488), .CO(n764), .S(n765) );
  CFA1X1 U490 ( .A(n1518), .B(n1398), .CI(n1338), .CO(n766), .S(n767) );
  CFA1X1 U491 ( .A(n1308), .B(n1278), .CI(n1248), .CO(n768), .S(n769) );
  CFA1X1 U492 ( .A(n1368), .B(n1548), .CI(n1578), .CO(n770), .S(n771) );
  CFA1X1 U493 ( .A(n1458), .B(n1608), .CI(n1639), .CO(n772), .S(n773) );
  CHA1X1 U494 ( .A(n1218), .B(n1141), .CO(n774), .S(n775) );
  CFA1X1 U495 ( .A(n781), .B(n779), .CI(n804), .CO(n776), .S(n777) );
  CFA1X1 U496 ( .A(n808), .B(n806), .CI(n783), .CO(n778), .S(n779) );
  CFA1X1 U497 ( .A(n787), .B(n785), .CI(n810), .CO(n780), .S(n781) );
  CFA1X1 U498 ( .A(n791), .B(n789), .CI(n812), .CO(n782), .S(n783) );
  CFA1X1 U499 ( .A(n795), .B(n814), .CI(n816), .CO(n784), .S(n785) );
  CFA1X1 U500 ( .A(n793), .B(n797), .CI(n799), .CO(n786), .S(n787) );
  CFA1X1 U501 ( .A(n822), .B(n801), .CI(n824), .CO(n788), .S(n789) );
  CFA1X1 U502 ( .A(n826), .B(n820), .CI(n818), .CO(n790), .S(n791) );
  CFA1X1 U503 ( .A(n1489), .B(n1459), .CI(n1429), .CO(n792), .S(n793) );
  CFA1X1 U504 ( .A(n1519), .B(n1399), .CI(n1369), .CO(n794), .S(n795) );
  CFA1X1 U505 ( .A(n1549), .B(n1339), .CI(n1309), .CO(n796), .S(n797) );
  CFA1X1 U506 ( .A(n1609), .B(n1579), .CI(n1249), .CO(n798), .S(n799) );
  CFA1X1 U507 ( .A(n1219), .B(n1640), .CI(n1279), .CO(n800), .S(n801) );
  CFA1X1 U508 ( .A(n807), .B(n805), .CI(n830), .CO(n802), .S(n803) );
  CFA1X1 U509 ( .A(n811), .B(n832), .CI(n809), .CO(n804), .S(n805) );
  CFA1X1 U510 ( .A(n836), .B(n834), .CI(n813), .CO(n806), .S(n807) );
  CFA1X1 U511 ( .A(n817), .B(n815), .CI(n838), .CO(n808), .S(n809) );
  CFA1X1 U512 ( .A(n821), .B(n840), .CI(n819), .CO(n810), .S(n811) );
  CFA1X1 U513 ( .A(n842), .B(n823), .CI(n825), .CO(n812), .S(n813) );
  CFA1X1 U514 ( .A(n844), .B(n848), .CI(n846), .CO(n814), .S(n815) );
  CFA1X1 U515 ( .A(n1550), .B(n850), .CI(n827), .CO(n816), .S(n817) );
  CFA1X1 U516 ( .A(n1580), .B(n1520), .CI(n1430), .CO(n818), .S(n819) );
  CFA1X1 U517 ( .A(n1400), .B(n1370), .CI(n1610), .CO(n820), .S(n821) );
  CFA1X1 U518 ( .A(n1490), .B(n1641), .CI(n1340), .CO(n822), .S(n823) );
  CFA1X1 U519 ( .A(n1460), .B(n1310), .CI(n1280), .CO(n824), .S(n825) );
  CHA1X1 U520 ( .A(n1250), .B(n1142), .CO(n826), .S(n827) );
  CFA1X1 U521 ( .A(n833), .B(n831), .CI(n854), .CO(n828), .S(n829) );
  CFA1X1 U522 ( .A(n858), .B(n835), .CI(n856), .CO(n830), .S(n831) );
  CFA1X1 U523 ( .A(n841), .B(n837), .CI(n839), .CO(n832), .S(n833) );
  CFA1X1 U524 ( .A(n864), .B(n860), .CI(n862), .CO(n834), .S(n835) );
  CFA1X1 U525 ( .A(n847), .B(n843), .CI(n849), .CO(n836), .S(n837) );
  CFA1X1 U526 ( .A(n870), .B(n845), .CI(n851), .CO(n838), .S(n839) );
  CFA1X1 U527 ( .A(n872), .B(n868), .CI(n866), .CO(n840), .S(n841) );
  CFA1X1 U528 ( .A(n1521), .B(n874), .CI(n1491), .CO(n842), .S(n843) );
  CFA1X1 U529 ( .A(n1551), .B(n1461), .CI(n1431), .CO(n844), .S(n845) );
  CFA1X1 U530 ( .A(n1581), .B(n1401), .CI(n1371), .CO(n846), .S(n847) );
  CFA1X1 U531 ( .A(n1611), .B(n1341), .CI(n1281), .CO(n848), .S(n849) );
  CFA1X1 U532 ( .A(n1251), .B(n1642), .CI(n1311), .CO(n850), .S(n851) );
  CFA1X1 U533 ( .A(n857), .B(n855), .CI(n878), .CO(n852), .S(n853) );
  CFA1X1 U534 ( .A(n882), .B(n880), .CI(n859), .CO(n854), .S(n855) );
  CFA1X1 U535 ( .A(n884), .B(n861), .CI(n863), .CO(n856), .S(n857) );
  CFA1X1 U536 ( .A(n888), .B(n865), .CI(n886), .CO(n858), .S(n859) );
  CFA1X1 U537 ( .A(n869), .B(n871), .CI(n873), .CO(n860), .S(n861) );
  CFA1X1 U538 ( .A(n892), .B(n867), .CI(n890), .CO(n862), .S(n863) );
  CFA1X1 U539 ( .A(n875), .B(n894), .CI(n896), .CO(n864), .S(n865) );
  CFA1X1 U540 ( .A(n1552), .B(n1522), .CI(n1462), .CO(n866), .S(n867) );
  CFA1X1 U541 ( .A(n1582), .B(n1432), .CI(n1372), .CO(n868), .S(n869) );
  CFA1X1 U542 ( .A(n1402), .B(n1342), .CI(n1312), .CO(n870), .S(n871) );
  CFA1X1 U543 ( .A(n1492), .B(n1612), .CI(n1643), .CO(n872), .S(n873) );
  CHA1X1 U544 ( .A(n1282), .B(n1143), .CO(n874), .S(n875) );
  CFA1X1 U545 ( .A(n881), .B(n879), .CI(n900), .CO(n876), .S(n877) );
  CFA1X1 U546 ( .A(n904), .B(n902), .CI(n883), .CO(n878), .S(n879) );
  CFA1X1 U547 ( .A(n906), .B(n885), .CI(n887), .CO(n880), .S(n881) );
  CFA1X1 U548 ( .A(n910), .B(n889), .CI(n908), .CO(n882), .S(n883) );
  CFA1X1 U549 ( .A(n891), .B(n893), .CI(n895), .CO(n884), .S(n885) );
  CFA1X1 U550 ( .A(n914), .B(n897), .CI(n912), .CO(n886), .S(n887) );
  CFA1X1 U551 ( .A(n1493), .B(n916), .CI(n918), .CO(n888), .S(n889) );
  CFA1X1 U552 ( .A(n1523), .B(n1463), .CI(n1433), .CO(n890), .S(n891) );
  CFA1X1 U553 ( .A(n1583), .B(n1553), .CI(n1403), .CO(n892), .S(n893) );
  CFA1X1 U554 ( .A(n1613), .B(n1373), .CI(n1313), .CO(n894), .S(n895) );
  CFA1X1 U555 ( .A(n1283), .B(n1644), .CI(n1343), .CO(n896), .S(n897) );
  CFA1X1 U556 ( .A(n903), .B(n901), .CI(n922), .CO(n898), .S(n899) );
  CFA1X1 U557 ( .A(n907), .B(n905), .CI(n924), .CO(n900), .S(n901) );
  CFA1X1 U558 ( .A(n928), .B(n926), .CI(n909), .CO(n902), .S(n903) );
  CFA1X1 U559 ( .A(n917), .B(n911), .CI(n930), .CO(n904), .S(n905) );
  CFA1X1 U560 ( .A(n936), .B(n915), .CI(n913), .CO(n906), .S(n907) );
  CFA1X1 U561 ( .A(n938), .B(n934), .CI(n932), .CO(n908), .S(n909) );
  CFA1X1 U562 ( .A(n1554), .B(n919), .CI(n1524), .CO(n910), .S(n911) );
  CFA1X1 U563 ( .A(n1584), .B(n1434), .CI(n1404), .CO(n912), .S(n913) );
  CFA1X1 U564 ( .A(n1464), .B(n1614), .CI(n1645), .CO(n914), .S(n915) );
  CFA1X1 U565 ( .A(n1494), .B(n1374), .CI(n1344), .CO(n916), .S(n917) );
  CHA1X1 U566 ( .A(n1314), .B(n1144), .CO(n918), .S(n919) );
  CFA1X1 U567 ( .A(n925), .B(n923), .CI(n942), .CO(n920), .S(n921) );
  CFA1X1 U568 ( .A(n929), .B(n944), .CI(n927), .CO(n922), .S(n923) );
  CFA1X1 U569 ( .A(n948), .B(n946), .CI(n931), .CO(n924), .S(n925) );
  CFA1X1 U570 ( .A(n935), .B(n950), .CI(n937), .CO(n926), .S(n927) );
  CFA1X1 U571 ( .A(n952), .B(n933), .CI(n939), .CO(n928), .S(n929) );
  CFA1X1 U572 ( .A(n958), .B(n954), .CI(n956), .CO(n930), .S(n931) );
  CFA1X1 U573 ( .A(n1555), .B(n1525), .CI(n1495), .CO(n932), .S(n933) );
  CFA1X1 U574 ( .A(n1585), .B(n1465), .CI(n1435), .CO(n934), .S(n935) );
  CFA1X1 U575 ( .A(n1615), .B(n1405), .CI(n1345), .CO(n936), .S(n937) );
  CFA1X1 U576 ( .A(n1315), .B(n1646), .CI(n1375), .CO(n938), .S(n939) );
  CFA1X1 U577 ( .A(n945), .B(n943), .CI(n962), .CO(n940), .S(n941) );
  CFA1X1 U578 ( .A(n949), .B(n964), .CI(n947), .CO(n942), .S(n943) );
  CFA1X1 U579 ( .A(n968), .B(n966), .CI(n951), .CO(n944), .S(n945) );
  CFA1X1 U580 ( .A(n953), .B(n955), .CI(n957), .CO(n946), .S(n947) );
  CFA1X1 U581 ( .A(n974), .B(n970), .CI(n972), .CO(n948), .S(n949) );
  CFA1X1 U582 ( .A(n1466), .B(n976), .CI(n959), .CO(n950), .S(n951) );
  CFA1X1 U583 ( .A(n1526), .B(n1406), .CI(n1376), .CO(n952), .S(n953) );
  CFA1X1 U584 ( .A(n1436), .B(n1556), .CI(n1586), .CO(n954), .S(n955) );
  CFA1X1 U585 ( .A(n1496), .B(n1616), .CI(n1647), .CO(n956), .S(n957) );
  CHA1X1 U586 ( .A(n1346), .B(n1145), .CO(n958), .S(n959) );
  CFA1X1 U587 ( .A(n965), .B(n963), .CI(n980), .CO(n960), .S(n961) );
  CFA1X1 U588 ( .A(n969), .B(n982), .CI(n967), .CO(n962), .S(n963) );
  CFA1X1 U589 ( .A(n971), .B(n984), .CI(n986), .CO(n964), .S(n965) );
  CFA1X1 U590 ( .A(n977), .B(n975), .CI(n973), .CO(n966), .S(n967) );
  CFA1X1 U591 ( .A(n992), .B(n990), .CI(n988), .CO(n968), .S(n969) );
  CFA1X1 U592 ( .A(n1557), .B(n994), .CI(n1527), .CO(n970), .S(n971) );
  CFA1X1 U593 ( .A(n1587), .B(n1497), .CI(n1467), .CO(n972), .S(n973) );
  CFA1X1 U594 ( .A(n1617), .B(n1437), .CI(n1377), .CO(n974), .S(n975) );
  CFA1X1 U595 ( .A(n1347), .B(n1648), .CI(n1407), .CO(n976), .S(n977) );
  CFA1X1 U596 ( .A(n983), .B(n981), .CI(n998), .CO(n978), .S(n979) );
  CFA1X1 U597 ( .A(n987), .B(n1000), .CI(n985), .CO(n980), .S(n981) );
  CFA1X1 U598 ( .A(n993), .B(n1002), .CI(n1004), .CO(n982), .S(n983) );
  CFA1X1 U599 ( .A(n1006), .B(n991), .CI(n989), .CO(n984), .S(n985) );
  CFA1X1 U600 ( .A(n995), .B(n1008), .CI(n1010), .CO(n986), .S(n987) );
  CFA1X1 U601 ( .A(n1618), .B(n1588), .CI(n1498), .CO(n988), .S(n989) );
  CFA1X1 U602 ( .A(n1558), .B(n1468), .CI(n1649), .CO(n990), .S(n991) );
  CFA1X1 U603 ( .A(n1528), .B(n1438), .CI(n1408), .CO(n992), .S(n993) );
  CHA1X1 U604 ( .A(n1378), .B(n1146), .CO(n994), .S(n995) );
  CFA1X1 U605 ( .A(n1001), .B(n999), .CI(n1014), .CO(n996), .S(n997) );
  CFA1X1 U606 ( .A(n1005), .B(n1016), .CI(n1003), .CO(n998), .S(n999) );
  CFA1X1 U607 ( .A(n1009), .B(n1018), .CI(n1020), .CO(n1000), .S(n1001) );
  CFA1X1 U608 ( .A(n1022), .B(n1007), .CI(n1011), .CO(n1002), .S(n1003) );
  CFA1X1 U609 ( .A(n1559), .B(n1024), .CI(n1026), .CO(n1004), .S(n1005) );
  CFA1X1 U610 ( .A(n1589), .B(n1529), .CI(n1499), .CO(n1006), .S(n1007) );
  CFA1X1 U611 ( .A(n1619), .B(n1469), .CI(n1409), .CO(n1008), .S(n1009) );
  CFA1X1 U612 ( .A(n1379), .B(n1650), .CI(n1439), .CO(n1010), .S(n1011) );
  CFA1X1 U613 ( .A(n1017), .B(n1015), .CI(n1030), .CO(n1012), .S(n1013) );
  CFA1X1 U614 ( .A(n1021), .B(n1032), .CI(n1019), .CO(n1014), .S(n1015) );
  CFA1X1 U615 ( .A(n1023), .B(n1034), .CI(n1025), .CO(n1016), .S(n1017) );
  CFA1X1 U616 ( .A(n1040), .B(n1038), .CI(n1036), .CO(n1018), .S(n1019) );
  CFA1X1 U617 ( .A(n1590), .B(n1027), .CI(n1560), .CO(n1020), .S(n1021) );
  CFA1X1 U618 ( .A(n1470), .B(n1500), .CI(n1440), .CO(n1022), .S(n1023) );
  CFA1X1 U619 ( .A(n1530), .B(n1620), .CI(n1651), .CO(n1024), .S(n1025) );
  CHA1X1 U620 ( .A(n1410), .B(n1147), .CO(n1026), .S(n1027) );
  CFA1X1 U621 ( .A(n1033), .B(n1031), .CI(n1044), .CO(n1028), .S(n1029) );
  CFA1X1 U622 ( .A(n1048), .B(n1035), .CI(n1046), .CO(n1030), .S(n1031) );
  CFA1X1 U623 ( .A(n1041), .B(n1039), .CI(n1037), .CO(n1032), .S(n1033) );
  CFA1X1 U624 ( .A(n1054), .B(n1050), .CI(n1052), .CO(n1034), .S(n1035) );
  CFA1X1 U625 ( .A(n1591), .B(n1561), .CI(n1531), .CO(n1036), .S(n1037) );
  CFA1X1 U626 ( .A(n1621), .B(n1501), .CI(n1441), .CO(n1038), .S(n1039) );
  CFA1X1 U627 ( .A(n1411), .B(n1652), .CI(n1471), .CO(n1040), .S(n1041) );
  CFA1X1 U628 ( .A(n1047), .B(n1045), .CI(n1058), .CO(n1042), .S(n1043) );
  CFA1X1 U629 ( .A(n1053), .B(n1049), .CI(n1060), .CO(n1044), .S(n1045) );
  CFA1X1 U630 ( .A(n1064), .B(n1051), .CI(n1062), .CO(n1046), .S(n1047) );
  CFA1X1 U631 ( .A(n1622), .B(n1066), .CI(n1055), .CO(n1048), .S(n1049) );
  CFA1X1 U632 ( .A(n1532), .B(n1592), .CI(n1653), .CO(n1050), .S(n1051) );
  CFA1X1 U633 ( .A(n1562), .B(n1502), .CI(n1472), .CO(n1052), .S(n1053) );
  CHA1X1 U634 ( .A(n1442), .B(n1148), .CO(n1054), .S(n1055) );
  CFA1X1 U635 ( .A(n1061), .B(n1059), .CI(n1070), .CO(n1056), .S(n1057) );
  CFA1X1 U636 ( .A(n1065), .B(n1072), .CI(n1063), .CO(n1058), .S(n1059) );
  CFA1X1 U637 ( .A(n1076), .B(n1067), .CI(n1074), .CO(n1060), .S(n1061) );
  CFA1X1 U638 ( .A(n1593), .B(n1078), .CI(n1563), .CO(n1062), .S(n1063) );
  CFA1X1 U639 ( .A(n1623), .B(n1533), .CI(n1473), .CO(n1064), .S(n1065) );
  CFA1X1 U640 ( .A(n1443), .B(n1654), .CI(n1503), .CO(n1066), .S(n1067) );
  CFA1X1 U641 ( .A(n1073), .B(n1071), .CI(n1082), .CO(n1068), .S(n1069) );
  CFA1X1 U642 ( .A(n1075), .B(n1084), .CI(n1077), .CO(n1070), .S(n1071) );
  CFA1X1 U643 ( .A(n1079), .B(n1086), .CI(n1088), .CO(n1072), .S(n1073) );
  CFA1X1 U644 ( .A(n1594), .B(n1534), .CI(n1504), .CO(n1074), .S(n1075) );
  CFA1X1 U645 ( .A(n1564), .B(n1624), .CI(n1655), .CO(n1076), .S(n1077) );
  CHA1X1 U646 ( .A(n1474), .B(n1149), .CO(n1078), .S(n1079) );
  CFA1X1 U647 ( .A(n1092), .B(n1083), .CI(n1085), .CO(n1080), .S(n1081) );
  CFA1X1 U648 ( .A(n1089), .B(n1094), .CI(n1087), .CO(n1082), .S(n1083) );
  CFA1X1 U649 ( .A(n1595), .B(n1096), .CI(n1098), .CO(n1084), .S(n1085) );
  CFA1X1 U650 ( .A(n1625), .B(n1565), .CI(n1505), .CO(n1086), .S(n1087) );
  CFA1X1 U651 ( .A(n1475), .B(n1656), .CI(n1535), .CO(n1088), .S(n1089) );
  CFA1X1 U652 ( .A(n1095), .B(n1093), .CI(n1102), .CO(n1090), .S(n1091) );
  CFA1X1 U653 ( .A(n1106), .B(n1097), .CI(n1104), .CO(n1092), .S(n1093) );
  CFA1X1 U654 ( .A(n1626), .B(n1099), .CI(n1566), .CO(n1094), .S(n1095) );
  CFA1X1 U655 ( .A(n1596), .B(n1657), .CI(n1536), .CO(n1096), .S(n1097) );
  CHA1X1 U656 ( .A(n1506), .B(n1150), .CO(n1098), .S(n1099) );
  CFA1X1 U657 ( .A(n1105), .B(n1103), .CI(n1110), .CO(n1100), .S(n1101) );
  CFA1X1 U658 ( .A(n1114), .B(n1107), .CI(n1112), .CO(n1102), .S(n1103) );
  CFA1X1 U659 ( .A(n1627), .B(n1597), .CI(n1537), .CO(n1104), .S(n1105) );
  CFA1X1 U660 ( .A(n1507), .B(n1658), .CI(n1567), .CO(n1106), .S(n1107) );
  CFA1X1 U661 ( .A(n1118), .B(n1111), .CI(n1113), .CO(n1108), .S(n1109) );
  CFA1X1 U662 ( .A(n1659), .B(n1120), .CI(n1115), .CO(n1110), .S(n1111) );
  CFA1X1 U663 ( .A(n1598), .B(n1628), .CI(n1568), .CO(n1112), .S(n1113) );
  CHA1X1 U664 ( .A(n1538), .B(n1151), .CO(n1114), .S(n1115) );
  CFA1X1 U665 ( .A(n1124), .B(n1119), .CI(n1121), .CO(n1116), .S(n1117) );
  CFA1X1 U666 ( .A(n1629), .B(n1126), .CI(n1569), .CO(n1118), .S(n1119) );
  CFA1X1 U667 ( .A(n1539), .B(n1660), .CI(n1599), .CO(n1120), .S(n1121) );
  CFA1X1 U668 ( .A(n1127), .B(n1125), .CI(n1130), .CO(n1122), .S(n1123) );
  CFA1X1 U669 ( .A(n1661), .B(n1630), .CI(n1600), .CO(n1124), .S(n1125) );
  CHA1X1 U670 ( .A(n1570), .B(n1152), .CO(n1126), .S(n1127) );
  CFA1X1 U671 ( .A(n1601), .B(n1131), .CI(n1134), .CO(n1128), .S(n1129) );
  CFA1X1 U672 ( .A(n1571), .B(n1631), .CI(n1662), .CO(n1130), .S(n1131) );
  CFA1X1 U673 ( .A(n1663), .B(n1135), .CI(n1632), .CO(n1132), .S(n1133) );
  CHA1X1 U674 ( .A(n1602), .B(n1153), .CO(n1134), .S(n1135) );
  CFA1X1 U675 ( .A(n1603), .B(n1633), .CI(n1664), .CO(n1136), .S(n1137) );
  CHA1X1 U676 ( .A(n1665), .B(n1634), .CO(n1138), .S(n1139) );
  CIVX2 U1861 ( .A(b[1]), .Z(n2453) );
  CIVX2 U1862 ( .A(b[3]), .Z(n2455) );
  CIVX2 U1863 ( .A(b[6]), .Z(n2458) );
  CIVX2 U1864 ( .A(b[2]), .Z(n2454) );
  CIVX2 U1865 ( .A(b[4]), .Z(n2456) );
  CIVX2 U1866 ( .A(b[5]), .Z(n2457) );
  CIVX2 U1867 ( .A(a[5]), .Z(n2487) );
  CIVX2 U1868 ( .A(a[3]), .Z(n2489) );
  CND2X1 U1869 ( .A(n2440), .B(n3065), .Z(n2535) );
  CND2X1 U1870 ( .A(n2439), .B(n3063), .Z(n2531) );
  CND2X1 U1871 ( .A(n2438), .B(n3061), .Z(n2527) );
  CND2X1 U1872 ( .A(a[1]), .B(n2491), .Z(n2582) );
  CIVX2 U1873 ( .A(a[1]), .Z(n2490) );
  CIVX2 U1874 ( .A(b[0]), .Z(n2515) );
  CIVX2 U1875 ( .A(a[0]), .Z(n2491) );
  CNIVX1 U1876 ( .A(n2536), .Z(n2440) );
  CEOX1 U1877 ( .A(n2487), .B(a[6]), .Z(n2536) );
  CNIVX1 U1878 ( .A(n2532), .Z(n2439) );
  CEOX1 U1879 ( .A(n2489), .B(a[4]), .Z(n2532) );
  CNIVX1 U1880 ( .A(n2528), .Z(n2438) );
  CEOX1 U1881 ( .A(n2490), .B(a[2]), .Z(n2528) );
  CIVX2 U1882 ( .A(a[11]), .Z(n2481) );
  CIVX2 U1883 ( .A(a[9]), .Z(n2483) );
  CIVX2 U1884 ( .A(a[7]), .Z(n2485) );
  CND2X1 U1885 ( .A(n2442), .B(n3069), .Z(n2543) );
  CND2X1 U1886 ( .A(n2441), .B(n3067), .Z(n2539) );
  CIVX2 U1887 ( .A(b[10]), .Z(n2511) );
  CIVX2 U1888 ( .A(b[9]), .Z(n2512) );
  CIVX2 U1889 ( .A(b[7]), .Z(n2514) );
  CIVX2 U1890 ( .A(b[8]), .Z(n2513) );
  CNIVX1 U1891 ( .A(n2544), .Z(n2442) );
  CEOX1 U1892 ( .A(n2483), .B(a[10]), .Z(n2544) );
  CNIVX1 U1893 ( .A(n2540), .Z(n2441) );
  CEOX1 U1894 ( .A(n2485), .B(a[8]), .Z(n2540) );
  CIVX2 U1895 ( .A(a[15]), .Z(n2477) );
  CIVX2 U1896 ( .A(a[13]), .Z(n2479) );
  CND2X1 U1897 ( .A(n2444), .B(n3073), .Z(n2549) );
  CND2X1 U1898 ( .A(n2443), .B(n3071), .Z(n2523) );
  CIVX2 U1899 ( .A(b[13]), .Z(n2508) );
  CIVX2 U1900 ( .A(b[12]), .Z(n2509) );
  CIVX2 U1901 ( .A(b[11]), .Z(n2510) );
  CNIVX1 U1902 ( .A(n2550), .Z(n2444) );
  CEOX1 U1903 ( .A(n2479), .B(a[14]), .Z(n2550) );
  CNIVX1 U1904 ( .A(n2525), .Z(n2443) );
  CEOX1 U1905 ( .A(n2481), .B(a[12]), .Z(n2525) );
  CIVX2 U1906 ( .A(a[19]), .Z(n2473) );
  CIVX2 U1907 ( .A(a[17]), .Z(n2475) );
  CND2X1 U1908 ( .A(n2445), .B(n3075), .Z(n2553) );
  CND2X1 U1909 ( .A(n2446), .B(n3077), .Z(n2557) );
  CIVX2 U1910 ( .A(b[18]), .Z(n2503) );
  CIVX2 U1911 ( .A(b[17]), .Z(n2504) );
  CIVX2 U1912 ( .A(b[14]), .Z(n2507) );
  CIVX2 U1913 ( .A(b[16]), .Z(n2505) );
  CIVX2 U1914 ( .A(b[15]), .Z(n2506) );
  CNIVX1 U1915 ( .A(n2554), .Z(n2445) );
  CEOX1 U1916 ( .A(n2477), .B(a[16]), .Z(n2554) );
  CNIVX1 U1917 ( .A(n2558), .Z(n2446) );
  CEOX1 U1918 ( .A(n2475), .B(a[18]), .Z(n2558) );
  CIVX2 U1919 ( .A(a[21]), .Z(n2471) );
  CIVX2 U1920 ( .A(a[23]), .Z(n2469) );
  CND2X1 U1921 ( .A(n2447), .B(n3079), .Z(n2561) );
  CND2X1 U1922 ( .A(n2448), .B(n3081), .Z(n2565) );
  CIVX2 U1923 ( .A(b[22]), .Z(n2499) );
  CIVX2 U1924 ( .A(b[20]), .Z(n2501) );
  CIVX2 U1925 ( .A(b[21]), .Z(n2500) );
  CIVX2 U1926 ( .A(b[19]), .Z(n2502) );
  CNIVX1 U1927 ( .A(n2562), .Z(n2447) );
  CEOX1 U1928 ( .A(n2473), .B(a[20]), .Z(n2562) );
  CNIVX1 U1929 ( .A(n2566), .Z(n2448) );
  CEOX1 U1930 ( .A(n2471), .B(a[22]), .Z(n2566) );
  CIVX2 U1931 ( .A(a[25]), .Z(n2467) );
  CIVX2 U1932 ( .A(a[27]), .Z(n2465) );
  CND2X1 U1933 ( .A(n2450), .B(n3085), .Z(n2573) );
  CND2X1 U1934 ( .A(n2449), .B(n3083), .Z(n2569) );
  CIVX2 U1935 ( .A(b[24]), .Z(n2497) );
  CIVX2 U1936 ( .A(b[25]), .Z(n2496) );
  CIVX2 U1937 ( .A(b[23]), .Z(n2498) );
  CNIVX1 U1938 ( .A(n2574), .Z(n2450) );
  CEOX1 U1939 ( .A(n2467), .B(a[26]), .Z(n2574) );
  CNIVX1 U1940 ( .A(n2570), .Z(n2449) );
  CEOX1 U1941 ( .A(n2469), .B(a[24]), .Z(n2570) );
  CIVX2 U1942 ( .A(a[29]), .Z(n2463) );
  CND2X1 U1943 ( .A(n2452), .B(n3089), .Z(n2579) );
  CND2X1 U1944 ( .A(n2451), .B(n3087), .Z(n2519) );
  CIVX2 U1945 ( .A(a[31]), .Z(n2461) );
  CIVX2 U1946 ( .A(b[29]), .Z(n2492) );
  CIVX2 U1947 ( .A(b[28]), .Z(n2493) );
  CIVX2 U1948 ( .A(b[27]), .Z(n2494) );
  CIVX2 U1949 ( .A(b[26]), .Z(n2495) );
  CNIVX1 U1950 ( .A(n2580), .Z(n2452) );
  CEOX1 U1951 ( .A(n2463), .B(a[30]), .Z(n2580) );
  CNIVX1 U1952 ( .A(n2520), .Z(n2451) );
  CEOX1 U1953 ( .A(n2465), .B(a[28]), .Z(n2520) );
  CIVX2 U1954 ( .A(n148), .Z(product[63]) );
  CIVX2 U1955 ( .A(n210), .Z(n2460) );
  CIVX2 U1956 ( .A(n216), .Z(n2462) );
  CIVX2 U1957 ( .A(n226), .Z(n2464) );
  CIVX2 U1958 ( .A(n240), .Z(n2466) );
  CIVX2 U1959 ( .A(n258), .Z(n2468) );
  CIVX2 U1960 ( .A(n280), .Z(n2470) );
  CIVX2 U1961 ( .A(n306), .Z(n2472) );
  CIVX2 U1962 ( .A(n336), .Z(n2474) );
  CIVX2 U1963 ( .A(n370), .Z(n2476) );
  CIVX2 U1964 ( .A(n408), .Z(n2478) );
  CIVX2 U1965 ( .A(n450), .Z(n2480) );
  CIVX2 U1966 ( .A(n496), .Z(n2482) );
  CIVX2 U1967 ( .A(n546), .Z(n2484) );
  CIVX2 U1968 ( .A(n600), .Z(n2486) );
  CIVX2 U1969 ( .A(n658), .Z(n2488) );
  CNR2X1 U1970 ( .A(n2491), .B(n2515), .Z(product[0]) );
  CENX1 U1971 ( .A(n2516), .B(n2517), .Z(n689) );
  COR2X1 U1972 ( .A(n2517), .B(n2516), .Z(n688) );
  COND2X1 U1973 ( .A(n2518), .B(n2519), .C(n2451), .D(n2521), .Z(n2516) );
  COND2X1 U1974 ( .A(n2522), .B(n2523), .C(n2524), .D(n2443), .Z(n2517) );
  COND2X1 U1975 ( .A(n2526), .B(n2527), .C(n2438), .D(n2529), .Z(n658) );
  COND2X1 U1976 ( .A(n2530), .B(n2531), .C(n2439), .D(n2533), .Z(n600) );
  COND2X1 U1977 ( .A(n2534), .B(n2535), .C(n2440), .D(n2537), .Z(n546) );
  COND2X1 U1978 ( .A(n2538), .B(n2539), .C(n2441), .D(n2541), .Z(n496) );
  COND2X1 U1979 ( .A(n2542), .B(n2543), .C(n2442), .D(n2545), .Z(n450) );
  COND2X1 U1980 ( .A(n2546), .B(n2523), .C(n2443), .D(n2547), .Z(n408) );
  COND2X1 U1981 ( .A(n2548), .B(n2549), .C(n2444), .D(n2551), .Z(n370) );
  COND2X1 U1982 ( .A(n2552), .B(n2553), .C(n2445), .D(n2555), .Z(n336) );
  COND2X1 U1983 ( .A(n2556), .B(n2557), .C(n2446), .D(n2559), .Z(n306) );
  COND2X1 U1984 ( .A(n2560), .B(n2561), .C(n2447), .D(n2563), .Z(n280) );
  COND2X1 U1985 ( .A(n2564), .B(n2565), .C(n2448), .D(n2567), .Z(n258) );
  COND2X1 U1986 ( .A(n2568), .B(n2569), .C(n2449), .D(n2571), .Z(n240) );
  COND2X1 U1987 ( .A(n2572), .B(n2573), .C(n2450), .D(n2575), .Z(n226) );
  COND2X1 U1988 ( .A(n2576), .B(n2519), .C(n2451), .D(n2577), .Z(n216) );
  COND2X1 U1989 ( .A(n2578), .B(n2579), .C(n2452), .D(n2581), .Z(n210) );
  COND2X1 U1990 ( .A(b[0]), .B(n2582), .C(n2583), .D(n2491), .Z(n1667) );
  COND2X1 U1991 ( .A(n2583), .B(n2582), .C(n2584), .D(n2491), .Z(n1666) );
  CENX1 U1992 ( .A(n2490), .B(n2453), .Z(n2583) );
  COND2X1 U1993 ( .A(n2584), .B(n2582), .C(n2585), .D(n2491), .Z(n1665) );
  CENX1 U1994 ( .A(n2490), .B(n2454), .Z(n2584) );
  COND2X1 U1995 ( .A(n2585), .B(n2582), .C(n2586), .D(n2491), .Z(n1664) );
  CENX1 U1996 ( .A(n2490), .B(n2455), .Z(n2585) );
  COND2X1 U1997 ( .A(n2586), .B(n2582), .C(n2587), .D(n2491), .Z(n1663) );
  CENX1 U1998 ( .A(n2490), .B(n2456), .Z(n2586) );
  COND2X1 U1999 ( .A(n2587), .B(n2582), .C(n2588), .D(n2491), .Z(n1662) );
  CENX1 U2000 ( .A(n2490), .B(n2457), .Z(n2587) );
  COND2X1 U2001 ( .A(n2588), .B(n2582), .C(n2589), .D(n2491), .Z(n1661) );
  CENX1 U2002 ( .A(n2490), .B(n2458), .Z(n2588) );
  COND2X1 U2003 ( .A(n2589), .B(n2582), .C(n2590), .D(n2491), .Z(n1660) );
  CENX1 U2004 ( .A(n2490), .B(n2514), .Z(n2589) );
  COND2X1 U2005 ( .A(n2590), .B(n2582), .C(n2591), .D(n2491), .Z(n1659) );
  CENX1 U2006 ( .A(n2490), .B(n2513), .Z(n2590) );
  COND2X1 U2007 ( .A(n2591), .B(n2582), .C(n2592), .D(n2491), .Z(n1658) );
  CENX1 U2008 ( .A(n2490), .B(n2512), .Z(n2591) );
  COND2X1 U2009 ( .A(n2592), .B(n2582), .C(n2593), .D(n2491), .Z(n1657) );
  CENX1 U2010 ( .A(n2490), .B(n2511), .Z(n2592) );
  COND2X1 U2011 ( .A(n2593), .B(n2582), .C(n2594), .D(n2491), .Z(n1656) );
  CENX1 U2012 ( .A(n2490), .B(n2510), .Z(n2593) );
  COND2X1 U2013 ( .A(n2594), .B(n2582), .C(n2595), .D(n2491), .Z(n1655) );
  CENX1 U2014 ( .A(n2490), .B(n2509), .Z(n2594) );
  COND2X1 U2015 ( .A(n2595), .B(n2582), .C(n2596), .D(n2491), .Z(n1654) );
  CENX1 U2016 ( .A(n2490), .B(n2508), .Z(n2595) );
  COND2X1 U2017 ( .A(n2596), .B(n2582), .C(n2597), .D(n2491), .Z(n1653) );
  CENX1 U2018 ( .A(n2490), .B(n2507), .Z(n2596) );
  COND2X1 U2019 ( .A(n2597), .B(n2582), .C(n2598), .D(n2491), .Z(n1652) );
  CENX1 U2020 ( .A(n2490), .B(n2506), .Z(n2597) );
  COND2X1 U2021 ( .A(n2598), .B(n2582), .C(n2599), .D(n2491), .Z(n1651) );
  CENX1 U2022 ( .A(n2490), .B(n2505), .Z(n2598) );
  COND2X1 U2023 ( .A(n2599), .B(n2582), .C(n2600), .D(n2491), .Z(n1650) );
  CENX1 U2024 ( .A(n2490), .B(n2504), .Z(n2599) );
  COND2X1 U2025 ( .A(n2600), .B(n2582), .C(n2601), .D(n2491), .Z(n1649) );
  CENX1 U2026 ( .A(n2490), .B(n2503), .Z(n2600) );
  COND2X1 U2027 ( .A(n2601), .B(n2582), .C(n2602), .D(n2491), .Z(n1648) );
  CENX1 U2028 ( .A(n2490), .B(n2502), .Z(n2601) );
  COND2X1 U2029 ( .A(n2602), .B(n2582), .C(n2603), .D(n2491), .Z(n1647) );
  CENX1 U2030 ( .A(n2490), .B(n2501), .Z(n2602) );
  COND2X1 U2031 ( .A(n2603), .B(n2582), .C(n2604), .D(n2491), .Z(n1646) );
  CENX1 U2032 ( .A(n2490), .B(n2500), .Z(n2603) );
  COND2X1 U2033 ( .A(n2604), .B(n2582), .C(n2605), .D(n2491), .Z(n1645) );
  CENX1 U2034 ( .A(n2490), .B(n2499), .Z(n2604) );
  COND2X1 U2035 ( .A(n2605), .B(n2582), .C(n2606), .D(n2491), .Z(n1644) );
  CENX1 U2036 ( .A(n2490), .B(n2498), .Z(n2605) );
  COND2X1 U2037 ( .A(n2606), .B(n2582), .C(n2607), .D(n2491), .Z(n1643) );
  CENX1 U2038 ( .A(n2490), .B(n2497), .Z(n2606) );
  COND2X1 U2039 ( .A(n2607), .B(n2582), .C(n2608), .D(n2491), .Z(n1642) );
  CENX1 U2040 ( .A(n2490), .B(n2496), .Z(n2607) );
  COND2X1 U2041 ( .A(n2608), .B(n2582), .C(n2609), .D(n2491), .Z(n1641) );
  CENX1 U2042 ( .A(n2490), .B(n2495), .Z(n2608) );
  COND2X1 U2043 ( .A(n2609), .B(n2582), .C(n2610), .D(n2491), .Z(n1640) );
  CENX1 U2044 ( .A(n2490), .B(n2494), .Z(n2609) );
  COND2X1 U2045 ( .A(n2610), .B(n2582), .C(n2611), .D(n2491), .Z(n1639) );
  CENX1 U2046 ( .A(n2490), .B(n2493), .Z(n2610) );
  COND2X1 U2047 ( .A(n2611), .B(n2582), .C(n2612), .D(n2491), .Z(n1638) );
  CENX1 U2048 ( .A(n2490), .B(n2492), .Z(n2611) );
  COND2X1 U2049 ( .A(n2612), .B(n2582), .C(n2613), .D(n2491), .Z(n1637) );
  CENX1 U2050 ( .A(a[1]), .B(b[30]), .Z(n2612) );
  CAOR1X1 U2051 ( .A(n2491), .B(n2582), .C(n2613), .Z(n1636) );
  CENX1 U2052 ( .A(a[1]), .B(b[31]), .Z(n2613) );
  CNR2X1 U2053 ( .A(n2438), .B(n2515), .Z(n1635) );
  COND2X1 U2054 ( .A(n2614), .B(n2527), .C(n2438), .D(n2615), .Z(n1634) );
  CENX1 U2055 ( .A(n2515), .B(n2489), .Z(n2614) );
  COND2X1 U2056 ( .A(n2615), .B(n2527), .C(n2438), .D(n2616), .Z(n1633) );
  CENX1 U2057 ( .A(n2489), .B(n2453), .Z(n2615) );
  COND2X1 U2058 ( .A(n2616), .B(n2527), .C(n2438), .D(n2617), .Z(n1632) );
  CENX1 U2059 ( .A(n2489), .B(n2454), .Z(n2616) );
  COND2X1 U2060 ( .A(n2617), .B(n2527), .C(n2438), .D(n2618), .Z(n1631) );
  CENX1 U2061 ( .A(n2489), .B(n2455), .Z(n2617) );
  COND2X1 U2062 ( .A(n2618), .B(n2527), .C(n2438), .D(n2619), .Z(n1630) );
  CENX1 U2063 ( .A(n2489), .B(n2456), .Z(n2618) );
  COND2X1 U2064 ( .A(n2619), .B(n2527), .C(n2438), .D(n2620), .Z(n1629) );
  CENX1 U2065 ( .A(n2489), .B(n2457), .Z(n2619) );
  COND2X1 U2066 ( .A(n2620), .B(n2527), .C(n2438), .D(n2621), .Z(n1628) );
  CENX1 U2067 ( .A(n2489), .B(n2458), .Z(n2620) );
  COND2X1 U2068 ( .A(n2621), .B(n2527), .C(n2438), .D(n2622), .Z(n1627) );
  CENX1 U2069 ( .A(n2489), .B(n2514), .Z(n2621) );
  COND2X1 U2070 ( .A(n2622), .B(n2527), .C(n2438), .D(n2623), .Z(n1626) );
  CENX1 U2071 ( .A(n2489), .B(n2513), .Z(n2622) );
  COND2X1 U2072 ( .A(n2623), .B(n2527), .C(n2438), .D(n2624), .Z(n1625) );
  CENX1 U2073 ( .A(n2489), .B(n2512), .Z(n2623) );
  COND2X1 U2074 ( .A(n2624), .B(n2527), .C(n2438), .D(n2625), .Z(n1624) );
  CENX1 U2075 ( .A(n2489), .B(n2511), .Z(n2624) );
  COND2X1 U2076 ( .A(n2625), .B(n2527), .C(n2438), .D(n2626), .Z(n1623) );
  CENX1 U2077 ( .A(n2489), .B(n2510), .Z(n2625) );
  COND2X1 U2078 ( .A(n2626), .B(n2527), .C(n2438), .D(n2627), .Z(n1622) );
  CENX1 U2079 ( .A(n2489), .B(n2509), .Z(n2626) );
  COND2X1 U2080 ( .A(n2627), .B(n2527), .C(n2438), .D(n2628), .Z(n1621) );
  CENX1 U2081 ( .A(n2489), .B(n2508), .Z(n2627) );
  COND2X1 U2082 ( .A(n2628), .B(n2527), .C(n2438), .D(n2629), .Z(n1620) );
  CENX1 U2083 ( .A(n2489), .B(n2507), .Z(n2628) );
  COND2X1 U2084 ( .A(n2629), .B(n2527), .C(n2438), .D(n2630), .Z(n1619) );
  CENX1 U2085 ( .A(n2489), .B(n2506), .Z(n2629) );
  COND2X1 U2086 ( .A(n2630), .B(n2527), .C(n2438), .D(n2631), .Z(n1618) );
  CENX1 U2087 ( .A(n2489), .B(n2505), .Z(n2630) );
  COND2X1 U2088 ( .A(n2631), .B(n2527), .C(n2438), .D(n2632), .Z(n1617) );
  CENX1 U2089 ( .A(n2489), .B(n2504), .Z(n2631) );
  COND2X1 U2090 ( .A(n2632), .B(n2527), .C(n2438), .D(n2633), .Z(n1616) );
  CENX1 U2091 ( .A(n2489), .B(n2503), .Z(n2632) );
  COND2X1 U2092 ( .A(n2633), .B(n2527), .C(n2438), .D(n2634), .Z(n1615) );
  CENX1 U2093 ( .A(n2489), .B(n2502), .Z(n2633) );
  COND2X1 U2094 ( .A(n2634), .B(n2527), .C(n2438), .D(n2635), .Z(n1614) );
  CENX1 U2095 ( .A(n2489), .B(n2501), .Z(n2634) );
  COND2X1 U2096 ( .A(n2635), .B(n2527), .C(n2438), .D(n2636), .Z(n1613) );
  CENX1 U2097 ( .A(n2489), .B(n2500), .Z(n2635) );
  COND2X1 U2098 ( .A(n2636), .B(n2527), .C(n2438), .D(n2637), .Z(n1612) );
  CENX1 U2099 ( .A(n2489), .B(n2499), .Z(n2636) );
  COND2X1 U2100 ( .A(n2637), .B(n2527), .C(n2438), .D(n2638), .Z(n1611) );
  CENX1 U2101 ( .A(n2489), .B(n2498), .Z(n2637) );
  COND2X1 U2102 ( .A(n2638), .B(n2527), .C(n2438), .D(n2639), .Z(n1610) );
  CENX1 U2103 ( .A(n2489), .B(n2497), .Z(n2638) );
  COND2X1 U2104 ( .A(n2639), .B(n2527), .C(n2438), .D(n2640), .Z(n1609) );
  CENX1 U2105 ( .A(n2489), .B(n2496), .Z(n2639) );
  COND2X1 U2106 ( .A(n2640), .B(n2527), .C(n2438), .D(n2641), .Z(n1608) );
  CENX1 U2107 ( .A(n2489), .B(n2495), .Z(n2640) );
  COND2X1 U2108 ( .A(n2641), .B(n2527), .C(n2438), .D(n2642), .Z(n1607) );
  CENX1 U2109 ( .A(n2489), .B(n2494), .Z(n2641) );
  COND2X1 U2110 ( .A(n2642), .B(n2527), .C(n2438), .D(n2643), .Z(n1606) );
  CENX1 U2111 ( .A(n2489), .B(n2493), .Z(n2642) );
  COND2X1 U2112 ( .A(n2643), .B(n2527), .C(n2438), .D(n2526), .Z(n1605) );
  CEOX1 U2113 ( .A(n2489), .B(b[30]), .Z(n2526) );
  CENX1 U2114 ( .A(n2489), .B(n2492), .Z(n2643) );
  CAOR1X1 U2115 ( .A(n2527), .B(n2438), .C(n2529), .Z(n1604) );
  CEOX1 U2116 ( .A(n2489), .B(b[31]), .Z(n2529) );
  CNR2X1 U2117 ( .A(n2439), .B(n2515), .Z(n1603) );
  COND2X1 U2118 ( .A(n2644), .B(n2531), .C(n2439), .D(n2645), .Z(n1602) );
  CENX1 U2119 ( .A(n2515), .B(n2487), .Z(n2644) );
  COND2X1 U2120 ( .A(n2645), .B(n2531), .C(n2439), .D(n2646), .Z(n1601) );
  CENX1 U2121 ( .A(n2487), .B(n2453), .Z(n2645) );
  COND2X1 U2122 ( .A(n2646), .B(n2531), .C(n2439), .D(n2647), .Z(n1600) );
  CENX1 U2123 ( .A(n2487), .B(n2454), .Z(n2646) );
  COND2X1 U2124 ( .A(n2647), .B(n2531), .C(n2439), .D(n2648), .Z(n1599) );
  CENX1 U2125 ( .A(n2487), .B(n2455), .Z(n2647) );
  COND2X1 U2126 ( .A(n2648), .B(n2531), .C(n2439), .D(n2649), .Z(n1598) );
  CENX1 U2127 ( .A(n2487), .B(n2456), .Z(n2648) );
  COND2X1 U2128 ( .A(n2649), .B(n2531), .C(n2439), .D(n2650), .Z(n1597) );
  CENX1 U2129 ( .A(n2487), .B(n2457), .Z(n2649) );
  COND2X1 U2130 ( .A(n2650), .B(n2531), .C(n2439), .D(n2651), .Z(n1596) );
  CENX1 U2131 ( .A(n2487), .B(n2458), .Z(n2650) );
  COND2X1 U2132 ( .A(n2651), .B(n2531), .C(n2439), .D(n2652), .Z(n1595) );
  CENX1 U2133 ( .A(n2487), .B(n2514), .Z(n2651) );
  COND2X1 U2134 ( .A(n2652), .B(n2531), .C(n2439), .D(n2653), .Z(n1594) );
  CENX1 U2135 ( .A(n2487), .B(n2513), .Z(n2652) );
  COND2X1 U2136 ( .A(n2653), .B(n2531), .C(n2439), .D(n2654), .Z(n1593) );
  CENX1 U2137 ( .A(n2487), .B(n2512), .Z(n2653) );
  COND2X1 U2138 ( .A(n2654), .B(n2531), .C(n2439), .D(n2655), .Z(n1592) );
  CENX1 U2139 ( .A(n2487), .B(n2511), .Z(n2654) );
  COND2X1 U2140 ( .A(n2655), .B(n2531), .C(n2439), .D(n2656), .Z(n1591) );
  CENX1 U2141 ( .A(n2487), .B(n2510), .Z(n2655) );
  COND2X1 U2142 ( .A(n2656), .B(n2531), .C(n2439), .D(n2657), .Z(n1590) );
  CENX1 U2143 ( .A(n2487), .B(n2509), .Z(n2656) );
  COND2X1 U2144 ( .A(n2657), .B(n2531), .C(n2439), .D(n2658), .Z(n1589) );
  CENX1 U2145 ( .A(n2487), .B(n2508), .Z(n2657) );
  COND2X1 U2146 ( .A(n2658), .B(n2531), .C(n2439), .D(n2659), .Z(n1588) );
  CENX1 U2147 ( .A(n2487), .B(n2507), .Z(n2658) );
  COND2X1 U2148 ( .A(n2659), .B(n2531), .C(n2439), .D(n2660), .Z(n1587) );
  CENX1 U2149 ( .A(n2487), .B(n2506), .Z(n2659) );
  COND2X1 U2150 ( .A(n2660), .B(n2531), .C(n2439), .D(n2661), .Z(n1586) );
  CENX1 U2151 ( .A(n2487), .B(n2505), .Z(n2660) );
  COND2X1 U2152 ( .A(n2661), .B(n2531), .C(n2439), .D(n2662), .Z(n1585) );
  CENX1 U2153 ( .A(n2487), .B(n2504), .Z(n2661) );
  COND2X1 U2154 ( .A(n2662), .B(n2531), .C(n2439), .D(n2663), .Z(n1584) );
  CENX1 U2155 ( .A(n2487), .B(n2503), .Z(n2662) );
  COND2X1 U2156 ( .A(n2663), .B(n2531), .C(n2439), .D(n2664), .Z(n1583) );
  CENX1 U2157 ( .A(n2487), .B(n2502), .Z(n2663) );
  COND2X1 U2158 ( .A(n2664), .B(n2531), .C(n2439), .D(n2665), .Z(n1582) );
  CENX1 U2159 ( .A(n2487), .B(n2501), .Z(n2664) );
  COND2X1 U2160 ( .A(n2665), .B(n2531), .C(n2439), .D(n2666), .Z(n1581) );
  CENX1 U2161 ( .A(n2487), .B(n2500), .Z(n2665) );
  COND2X1 U2162 ( .A(n2666), .B(n2531), .C(n2439), .D(n2667), .Z(n1580) );
  CENX1 U2163 ( .A(n2487), .B(n2499), .Z(n2666) );
  COND2X1 U2164 ( .A(n2667), .B(n2531), .C(n2439), .D(n2668), .Z(n1579) );
  CENX1 U2165 ( .A(n2487), .B(n2498), .Z(n2667) );
  COND2X1 U2166 ( .A(n2668), .B(n2531), .C(n2439), .D(n2669), .Z(n1578) );
  CENX1 U2167 ( .A(n2487), .B(n2497), .Z(n2668) );
  COND2X1 U2168 ( .A(n2669), .B(n2531), .C(n2439), .D(n2670), .Z(n1577) );
  CENX1 U2169 ( .A(n2487), .B(n2496), .Z(n2669) );
  COND2X1 U2170 ( .A(n2670), .B(n2531), .C(n2439), .D(n2671), .Z(n1576) );
  CENX1 U2171 ( .A(n2487), .B(n2495), .Z(n2670) );
  COND2X1 U2172 ( .A(n2671), .B(n2531), .C(n2439), .D(n2672), .Z(n1575) );
  CENX1 U2173 ( .A(n2487), .B(n2494), .Z(n2671) );
  COND2X1 U2174 ( .A(n2672), .B(n2531), .C(n2439), .D(n2673), .Z(n1574) );
  CENX1 U2175 ( .A(n2487), .B(n2493), .Z(n2672) );
  COND2X1 U2176 ( .A(n2673), .B(n2531), .C(n2439), .D(n2530), .Z(n1573) );
  CEOX1 U2177 ( .A(n2487), .B(b[30]), .Z(n2530) );
  CENX1 U2178 ( .A(n2487), .B(n2492), .Z(n2673) );
  CAOR1X1 U2179 ( .A(n2531), .B(n2439), .C(n2533), .Z(n1572) );
  CEOX1 U2180 ( .A(n2487), .B(b[31]), .Z(n2533) );
  CNR2X1 U2181 ( .A(n2440), .B(n2515), .Z(n1571) );
  COND2X1 U2182 ( .A(n2674), .B(n2535), .C(n2440), .D(n2675), .Z(n1570) );
  CENX1 U2183 ( .A(n2515), .B(n2485), .Z(n2674) );
  COND2X1 U2184 ( .A(n2675), .B(n2535), .C(n2440), .D(n2676), .Z(n1569) );
  CENX1 U2185 ( .A(n2485), .B(n2453), .Z(n2675) );
  COND2X1 U2186 ( .A(n2676), .B(n2535), .C(n2440), .D(n2677), .Z(n1568) );
  CENX1 U2187 ( .A(n2485), .B(n2454), .Z(n2676) );
  COND2X1 U2188 ( .A(n2677), .B(n2535), .C(n2440), .D(n2678), .Z(n1567) );
  CENX1 U2189 ( .A(n2485), .B(n2455), .Z(n2677) );
  COND2X1 U2190 ( .A(n2678), .B(n2535), .C(n2440), .D(n2679), .Z(n1566) );
  CENX1 U2191 ( .A(n2485), .B(n2456), .Z(n2678) );
  COND2X1 U2192 ( .A(n2679), .B(n2535), .C(n2440), .D(n2680), .Z(n1565) );
  CENX1 U2193 ( .A(n2485), .B(n2457), .Z(n2679) );
  COND2X1 U2194 ( .A(n2680), .B(n2535), .C(n2440), .D(n2681), .Z(n1564) );
  CENX1 U2195 ( .A(n2485), .B(n2458), .Z(n2680) );
  COND2X1 U2196 ( .A(n2681), .B(n2535), .C(n2440), .D(n2682), .Z(n1563) );
  CENX1 U2197 ( .A(n2485), .B(n2514), .Z(n2681) );
  COND2X1 U2198 ( .A(n2682), .B(n2535), .C(n2440), .D(n2683), .Z(n1562) );
  CENX1 U2199 ( .A(n2485), .B(n2513), .Z(n2682) );
  COND2X1 U2200 ( .A(n2683), .B(n2535), .C(n2440), .D(n2684), .Z(n1561) );
  CENX1 U2201 ( .A(n2485), .B(n2512), .Z(n2683) );
  COND2X1 U2202 ( .A(n2684), .B(n2535), .C(n2440), .D(n2685), .Z(n1560) );
  CENX1 U2203 ( .A(n2485), .B(n2511), .Z(n2684) );
  COND2X1 U2204 ( .A(n2685), .B(n2535), .C(n2440), .D(n2686), .Z(n1559) );
  CENX1 U2205 ( .A(n2485), .B(n2510), .Z(n2685) );
  COND2X1 U2206 ( .A(n2686), .B(n2535), .C(n2440), .D(n2687), .Z(n1558) );
  CENX1 U2207 ( .A(n2485), .B(n2509), .Z(n2686) );
  COND2X1 U2208 ( .A(n2687), .B(n2535), .C(n2440), .D(n2688), .Z(n1557) );
  CENX1 U2209 ( .A(n2485), .B(n2508), .Z(n2687) );
  COND2X1 U2210 ( .A(n2688), .B(n2535), .C(n2440), .D(n2689), .Z(n1556) );
  CENX1 U2211 ( .A(n2485), .B(n2507), .Z(n2688) );
  COND2X1 U2212 ( .A(n2689), .B(n2535), .C(n2440), .D(n2690), .Z(n1555) );
  CENX1 U2213 ( .A(n2485), .B(n2506), .Z(n2689) );
  COND2X1 U2214 ( .A(n2690), .B(n2535), .C(n2440), .D(n2691), .Z(n1554) );
  CENX1 U2215 ( .A(n2485), .B(n2505), .Z(n2690) );
  COND2X1 U2216 ( .A(n2691), .B(n2535), .C(n2440), .D(n2692), .Z(n1553) );
  CENX1 U2217 ( .A(n2485), .B(n2504), .Z(n2691) );
  COND2X1 U2218 ( .A(n2692), .B(n2535), .C(n2440), .D(n2693), .Z(n1552) );
  CENX1 U2219 ( .A(n2485), .B(n2503), .Z(n2692) );
  COND2X1 U2220 ( .A(n2693), .B(n2535), .C(n2440), .D(n2694), .Z(n1551) );
  CENX1 U2221 ( .A(n2485), .B(n2502), .Z(n2693) );
  COND2X1 U2222 ( .A(n2694), .B(n2535), .C(n2440), .D(n2695), .Z(n1550) );
  CENX1 U2223 ( .A(n2485), .B(n2501), .Z(n2694) );
  COND2X1 U2224 ( .A(n2695), .B(n2535), .C(n2440), .D(n2696), .Z(n1549) );
  CENX1 U2225 ( .A(n2485), .B(n2500), .Z(n2695) );
  COND2X1 U2226 ( .A(n2696), .B(n2535), .C(n2440), .D(n2697), .Z(n1548) );
  CENX1 U2227 ( .A(n2485), .B(n2499), .Z(n2696) );
  COND2X1 U2228 ( .A(n2697), .B(n2535), .C(n2440), .D(n2698), .Z(n1547) );
  CENX1 U2229 ( .A(n2485), .B(n2498), .Z(n2697) );
  COND2X1 U2230 ( .A(n2698), .B(n2535), .C(n2440), .D(n2699), .Z(n1546) );
  CENX1 U2231 ( .A(n2485), .B(n2497), .Z(n2698) );
  COND2X1 U2232 ( .A(n2699), .B(n2535), .C(n2440), .D(n2700), .Z(n1545) );
  CENX1 U2233 ( .A(n2485), .B(n2496), .Z(n2699) );
  COND2X1 U2234 ( .A(n2700), .B(n2535), .C(n2440), .D(n2701), .Z(n1544) );
  CENX1 U2235 ( .A(n2485), .B(n2495), .Z(n2700) );
  COND2X1 U2236 ( .A(n2701), .B(n2535), .C(n2440), .D(n2702), .Z(n1543) );
  CENX1 U2237 ( .A(n2485), .B(n2494), .Z(n2701) );
  COND2X1 U2238 ( .A(n2702), .B(n2535), .C(n2440), .D(n2703), .Z(n1542) );
  CENX1 U2239 ( .A(n2485), .B(n2493), .Z(n2702) );
  COND2X1 U2240 ( .A(n2703), .B(n2535), .C(n2440), .D(n2534), .Z(n1541) );
  CEOX1 U2241 ( .A(n2485), .B(b[30]), .Z(n2534) );
  CENX1 U2242 ( .A(n2485), .B(n2492), .Z(n2703) );
  CAOR1X1 U2243 ( .A(n2535), .B(n2440), .C(n2537), .Z(n1540) );
  CEOX1 U2244 ( .A(n2485), .B(b[31]), .Z(n2537) );
  CNR2X1 U2245 ( .A(n2441), .B(n2515), .Z(n1539) );
  COND2X1 U2246 ( .A(n2704), .B(n2539), .C(n2441), .D(n2705), .Z(n1538) );
  CENX1 U2247 ( .A(n2515), .B(n2483), .Z(n2704) );
  COND2X1 U2248 ( .A(n2705), .B(n2539), .C(n2441), .D(n2706), .Z(n1537) );
  CENX1 U2249 ( .A(n2483), .B(n2453), .Z(n2705) );
  COND2X1 U2250 ( .A(n2706), .B(n2539), .C(n2441), .D(n2707), .Z(n1536) );
  CENX1 U2251 ( .A(n2483), .B(n2454), .Z(n2706) );
  COND2X1 U2252 ( .A(n2707), .B(n2539), .C(n2441), .D(n2708), .Z(n1535) );
  CENX1 U2253 ( .A(n2483), .B(n2455), .Z(n2707) );
  COND2X1 U2254 ( .A(n2708), .B(n2539), .C(n2441), .D(n2709), .Z(n1534) );
  CENX1 U2255 ( .A(n2483), .B(n2456), .Z(n2708) );
  COND2X1 U2256 ( .A(n2709), .B(n2539), .C(n2441), .D(n2710), .Z(n1533) );
  CENX1 U2257 ( .A(n2483), .B(n2457), .Z(n2709) );
  COND2X1 U2258 ( .A(n2710), .B(n2539), .C(n2441), .D(n2711), .Z(n1532) );
  CENX1 U2259 ( .A(n2483), .B(n2458), .Z(n2710) );
  COND2X1 U2260 ( .A(n2711), .B(n2539), .C(n2441), .D(n2712), .Z(n1531) );
  CENX1 U2261 ( .A(n2483), .B(n2514), .Z(n2711) );
  COND2X1 U2262 ( .A(n2712), .B(n2539), .C(n2441), .D(n2713), .Z(n1530) );
  CENX1 U2263 ( .A(n2483), .B(n2513), .Z(n2712) );
  COND2X1 U2264 ( .A(n2713), .B(n2539), .C(n2441), .D(n2714), .Z(n1529) );
  CENX1 U2265 ( .A(n2483), .B(n2512), .Z(n2713) );
  COND2X1 U2266 ( .A(n2714), .B(n2539), .C(n2441), .D(n2715), .Z(n1528) );
  CENX1 U2267 ( .A(n2483), .B(n2511), .Z(n2714) );
  COND2X1 U2268 ( .A(n2715), .B(n2539), .C(n2441), .D(n2716), .Z(n1527) );
  CENX1 U2269 ( .A(n2483), .B(n2510), .Z(n2715) );
  COND2X1 U2270 ( .A(n2716), .B(n2539), .C(n2441), .D(n2717), .Z(n1526) );
  CENX1 U2271 ( .A(n2483), .B(n2509), .Z(n2716) );
  COND2X1 U2272 ( .A(n2717), .B(n2539), .C(n2441), .D(n2718), .Z(n1525) );
  CENX1 U2273 ( .A(n2483), .B(n2508), .Z(n2717) );
  COND2X1 U2274 ( .A(n2718), .B(n2539), .C(n2441), .D(n2719), .Z(n1524) );
  CENX1 U2275 ( .A(n2483), .B(n2507), .Z(n2718) );
  COND2X1 U2276 ( .A(n2719), .B(n2539), .C(n2441), .D(n2720), .Z(n1523) );
  CENX1 U2277 ( .A(n2483), .B(n2506), .Z(n2719) );
  COND2X1 U2278 ( .A(n2720), .B(n2539), .C(n2441), .D(n2721), .Z(n1522) );
  CENX1 U2279 ( .A(n2483), .B(n2505), .Z(n2720) );
  COND2X1 U2280 ( .A(n2721), .B(n2539), .C(n2441), .D(n2722), .Z(n1521) );
  CENX1 U2281 ( .A(n2483), .B(n2504), .Z(n2721) );
  COND2X1 U2282 ( .A(n2722), .B(n2539), .C(n2441), .D(n2723), .Z(n1520) );
  CENX1 U2283 ( .A(n2483), .B(n2503), .Z(n2722) );
  COND2X1 U2284 ( .A(n2723), .B(n2539), .C(n2441), .D(n2724), .Z(n1519) );
  CENX1 U2285 ( .A(n2483), .B(n2502), .Z(n2723) );
  COND2X1 U2286 ( .A(n2724), .B(n2539), .C(n2441), .D(n2725), .Z(n1518) );
  CENX1 U2287 ( .A(n2483), .B(n2501), .Z(n2724) );
  COND2X1 U2288 ( .A(n2725), .B(n2539), .C(n2441), .D(n2726), .Z(n1517) );
  CENX1 U2289 ( .A(n2483), .B(n2500), .Z(n2725) );
  COND2X1 U2290 ( .A(n2726), .B(n2539), .C(n2441), .D(n2727), .Z(n1516) );
  CENX1 U2291 ( .A(n2483), .B(n2499), .Z(n2726) );
  COND2X1 U2292 ( .A(n2727), .B(n2539), .C(n2441), .D(n2728), .Z(n1515) );
  CENX1 U2293 ( .A(n2483), .B(n2498), .Z(n2727) );
  COND2X1 U2294 ( .A(n2728), .B(n2539), .C(n2441), .D(n2729), .Z(n1514) );
  CENX1 U2295 ( .A(n2483), .B(n2497), .Z(n2728) );
  COND2X1 U2296 ( .A(n2729), .B(n2539), .C(n2441), .D(n2730), .Z(n1513) );
  CENX1 U2297 ( .A(n2483), .B(n2496), .Z(n2729) );
  COND2X1 U2298 ( .A(n2730), .B(n2539), .C(n2441), .D(n2731), .Z(n1512) );
  CENX1 U2299 ( .A(n2483), .B(n2495), .Z(n2730) );
  COND2X1 U2300 ( .A(n2731), .B(n2539), .C(n2441), .D(n2732), .Z(n1511) );
  CENX1 U2301 ( .A(n2483), .B(n2494), .Z(n2731) );
  COND2X1 U2302 ( .A(n2732), .B(n2539), .C(n2441), .D(n2733), .Z(n1510) );
  CENX1 U2303 ( .A(n2483), .B(n2493), .Z(n2732) );
  COND2X1 U2304 ( .A(n2733), .B(n2539), .C(n2441), .D(n2538), .Z(n1509) );
  CEOX1 U2305 ( .A(n2483), .B(b[30]), .Z(n2538) );
  CENX1 U2306 ( .A(n2483), .B(n2492), .Z(n2733) );
  CAOR1X1 U2307 ( .A(n2539), .B(n2441), .C(n2541), .Z(n1508) );
  CEOX1 U2308 ( .A(n2483), .B(b[31]), .Z(n2541) );
  CNR2X1 U2309 ( .A(n2442), .B(n2515), .Z(n1507) );
  COND2X1 U2310 ( .A(n2734), .B(n2543), .C(n2442), .D(n2735), .Z(n1506) );
  CENX1 U2311 ( .A(n2515), .B(n2481), .Z(n2734) );
  COND2X1 U2312 ( .A(n2735), .B(n2543), .C(n2442), .D(n2736), .Z(n1505) );
  CENX1 U2313 ( .A(n2481), .B(n2453), .Z(n2735) );
  COND2X1 U2314 ( .A(n2736), .B(n2543), .C(n2442), .D(n2737), .Z(n1504) );
  CENX1 U2315 ( .A(n2481), .B(n2454), .Z(n2736) );
  COND2X1 U2316 ( .A(n2737), .B(n2543), .C(n2442), .D(n2738), .Z(n1503) );
  CENX1 U2317 ( .A(n2481), .B(n2455), .Z(n2737) );
  COND2X1 U2318 ( .A(n2738), .B(n2543), .C(n2442), .D(n2739), .Z(n1502) );
  CENX1 U2319 ( .A(n2481), .B(n2456), .Z(n2738) );
  COND2X1 U2320 ( .A(n2739), .B(n2543), .C(n2442), .D(n2740), .Z(n1501) );
  CENX1 U2321 ( .A(n2481), .B(n2457), .Z(n2739) );
  COND2X1 U2322 ( .A(n2740), .B(n2543), .C(n2442), .D(n2741), .Z(n1500) );
  CENX1 U2323 ( .A(n2481), .B(n2458), .Z(n2740) );
  COND2X1 U2324 ( .A(n2741), .B(n2543), .C(n2442), .D(n2742), .Z(n1499) );
  CENX1 U2325 ( .A(n2481), .B(n2514), .Z(n2741) );
  COND2X1 U2326 ( .A(n2742), .B(n2543), .C(n2442), .D(n2743), .Z(n1498) );
  CENX1 U2327 ( .A(n2481), .B(n2513), .Z(n2742) );
  COND2X1 U2328 ( .A(n2743), .B(n2543), .C(n2442), .D(n2744), .Z(n1497) );
  CENX1 U2329 ( .A(n2481), .B(n2512), .Z(n2743) );
  COND2X1 U2330 ( .A(n2744), .B(n2543), .C(n2442), .D(n2745), .Z(n1496) );
  CENX1 U2331 ( .A(n2481), .B(n2511), .Z(n2744) );
  COND2X1 U2332 ( .A(n2745), .B(n2543), .C(n2442), .D(n2746), .Z(n1495) );
  CENX1 U2333 ( .A(n2481), .B(n2510), .Z(n2745) );
  COND2X1 U2334 ( .A(n2746), .B(n2543), .C(n2442), .D(n2747), .Z(n1494) );
  CENX1 U2335 ( .A(n2481), .B(n2509), .Z(n2746) );
  COND2X1 U2336 ( .A(n2747), .B(n2543), .C(n2442), .D(n2748), .Z(n1493) );
  CENX1 U2337 ( .A(n2481), .B(n2508), .Z(n2747) );
  COND2X1 U2338 ( .A(n2748), .B(n2543), .C(n2442), .D(n2749), .Z(n1492) );
  CENX1 U2339 ( .A(n2481), .B(n2507), .Z(n2748) );
  COND2X1 U2340 ( .A(n2749), .B(n2543), .C(n2442), .D(n2750), .Z(n1491) );
  CENX1 U2341 ( .A(n2481), .B(n2506), .Z(n2749) );
  COND2X1 U2342 ( .A(n2750), .B(n2543), .C(n2442), .D(n2751), .Z(n1490) );
  CENX1 U2343 ( .A(n2481), .B(n2505), .Z(n2750) );
  COND2X1 U2344 ( .A(n2751), .B(n2543), .C(n2442), .D(n2752), .Z(n1489) );
  CENX1 U2345 ( .A(n2481), .B(n2504), .Z(n2751) );
  COND2X1 U2346 ( .A(n2752), .B(n2543), .C(n2442), .D(n2753), .Z(n1488) );
  CENX1 U2347 ( .A(n2481), .B(n2503), .Z(n2752) );
  COND2X1 U2348 ( .A(n2753), .B(n2543), .C(n2442), .D(n2754), .Z(n1487) );
  CENX1 U2349 ( .A(n2481), .B(n2502), .Z(n2753) );
  COND2X1 U2350 ( .A(n2754), .B(n2543), .C(n2442), .D(n2755), .Z(n1486) );
  CENX1 U2351 ( .A(n2481), .B(n2501), .Z(n2754) );
  COND2X1 U2352 ( .A(n2755), .B(n2543), .C(n2442), .D(n2756), .Z(n1485) );
  CENX1 U2353 ( .A(n2481), .B(n2500), .Z(n2755) );
  COND2X1 U2354 ( .A(n2756), .B(n2543), .C(n2442), .D(n2757), .Z(n1484) );
  CENX1 U2355 ( .A(n2481), .B(n2499), .Z(n2756) );
  COND2X1 U2356 ( .A(n2757), .B(n2543), .C(n2442), .D(n2758), .Z(n1483) );
  CENX1 U2357 ( .A(n2481), .B(n2498), .Z(n2757) );
  COND2X1 U2358 ( .A(n2758), .B(n2543), .C(n2442), .D(n2759), .Z(n1482) );
  CENX1 U2359 ( .A(n2481), .B(n2497), .Z(n2758) );
  COND2X1 U2360 ( .A(n2759), .B(n2543), .C(n2442), .D(n2760), .Z(n1481) );
  CENX1 U2361 ( .A(n2481), .B(n2496), .Z(n2759) );
  COND2X1 U2362 ( .A(n2760), .B(n2543), .C(n2442), .D(n2761), .Z(n1480) );
  CENX1 U2363 ( .A(n2481), .B(n2495), .Z(n2760) );
  COND2X1 U2364 ( .A(n2761), .B(n2543), .C(n2442), .D(n2762), .Z(n1479) );
  CENX1 U2365 ( .A(n2481), .B(n2494), .Z(n2761) );
  COND2X1 U2366 ( .A(n2762), .B(n2543), .C(n2442), .D(n2763), .Z(n1478) );
  CENX1 U2367 ( .A(n2481), .B(n2493), .Z(n2762) );
  COND2X1 U2368 ( .A(n2763), .B(n2543), .C(n2442), .D(n2542), .Z(n1477) );
  CEOX1 U2369 ( .A(n2481), .B(b[30]), .Z(n2542) );
  CENX1 U2370 ( .A(n2481), .B(n2492), .Z(n2763) );
  CAOR1X1 U2371 ( .A(n2543), .B(n2442), .C(n2545), .Z(n1476) );
  CEOX1 U2372 ( .A(n2481), .B(b[31]), .Z(n2545) );
  CNR2X1 U2373 ( .A(n2443), .B(n2515), .Z(n1475) );
  COND2X1 U2374 ( .A(n2764), .B(n2523), .C(n2443), .D(n2765), .Z(n1474) );
  CENX1 U2375 ( .A(n2515), .B(n2479), .Z(n2764) );
  COND2X1 U2376 ( .A(n2765), .B(n2523), .C(n2443), .D(n2766), .Z(n1473) );
  CENX1 U2377 ( .A(n2479), .B(n2453), .Z(n2765) );
  COND2X1 U2378 ( .A(n2766), .B(n2523), .C(n2443), .D(n2767), .Z(n1472) );
  CENX1 U2379 ( .A(n2479), .B(n2454), .Z(n2766) );
  COND2X1 U2380 ( .A(n2767), .B(n2523), .C(n2443), .D(n2768), .Z(n1471) );
  CENX1 U2381 ( .A(n2479), .B(n2455), .Z(n2767) );
  COND2X1 U2382 ( .A(n2768), .B(n2523), .C(n2443), .D(n2769), .Z(n1470) );
  CENX1 U2383 ( .A(n2479), .B(n2456), .Z(n2768) );
  COND2X1 U2384 ( .A(n2769), .B(n2523), .C(n2443), .D(n2770), .Z(n1469) );
  CENX1 U2385 ( .A(n2479), .B(n2457), .Z(n2769) );
  COND2X1 U2386 ( .A(n2770), .B(n2523), .C(n2443), .D(n2771), .Z(n1468) );
  CENX1 U2387 ( .A(n2479), .B(n2458), .Z(n2770) );
  COND2X1 U2388 ( .A(n2771), .B(n2523), .C(n2443), .D(n2772), .Z(n1467) );
  CENX1 U2389 ( .A(n2479), .B(n2514), .Z(n2771) );
  COND2X1 U2390 ( .A(n2772), .B(n2523), .C(n2443), .D(n2773), .Z(n1466) );
  CENX1 U2391 ( .A(n2479), .B(n2513), .Z(n2772) );
  COND2X1 U2392 ( .A(n2773), .B(n2523), .C(n2443), .D(n2774), .Z(n1465) );
  CENX1 U2393 ( .A(n2479), .B(n2512), .Z(n2773) );
  COND2X1 U2394 ( .A(n2774), .B(n2523), .C(n2443), .D(n2775), .Z(n1464) );
  CENX1 U2395 ( .A(n2479), .B(n2511), .Z(n2774) );
  COND2X1 U2396 ( .A(n2775), .B(n2523), .C(n2443), .D(n2776), .Z(n1463) );
  CENX1 U2397 ( .A(n2479), .B(n2510), .Z(n2775) );
  COND2X1 U2398 ( .A(n2776), .B(n2523), .C(n2443), .D(n2777), .Z(n1462) );
  CENX1 U2399 ( .A(n2479), .B(n2509), .Z(n2776) );
  COND2X1 U2400 ( .A(n2777), .B(n2523), .C(n2443), .D(n2778), .Z(n1461) );
  CENX1 U2401 ( .A(n2479), .B(n2508), .Z(n2777) );
  COND2X1 U2402 ( .A(n2778), .B(n2523), .C(n2443), .D(n2779), .Z(n1460) );
  CENX1 U2403 ( .A(n2479), .B(n2507), .Z(n2778) );
  COND2X1 U2404 ( .A(n2779), .B(n2523), .C(n2443), .D(n2780), .Z(n1459) );
  CENX1 U2405 ( .A(n2479), .B(n2506), .Z(n2779) );
  COND2X1 U2406 ( .A(n2780), .B(n2523), .C(n2443), .D(n2781), .Z(n1458) );
  CENX1 U2407 ( .A(n2479), .B(n2505), .Z(n2780) );
  COND2X1 U2408 ( .A(n2781), .B(n2523), .C(n2443), .D(n2782), .Z(n1457) );
  CENX1 U2409 ( .A(n2479), .B(n2504), .Z(n2781) );
  COND2X1 U2410 ( .A(n2782), .B(n2523), .C(n2443), .D(n2522), .Z(n1456) );
  CENX1 U2411 ( .A(n2479), .B(n2502), .Z(n2522) );
  CENX1 U2412 ( .A(n2479), .B(n2503), .Z(n2782) );
  COND2X1 U2413 ( .A(n2524), .B(n2523), .C(n2443), .D(n2783), .Z(n1454) );
  CENX1 U2414 ( .A(n2479), .B(n2501), .Z(n2524) );
  COND2X1 U2415 ( .A(n2783), .B(n2523), .C(n2443), .D(n2784), .Z(n1453) );
  CENX1 U2416 ( .A(n2479), .B(n2500), .Z(n2783) );
  COND2X1 U2417 ( .A(n2784), .B(n2523), .C(n2443), .D(n2785), .Z(n1452) );
  CENX1 U2418 ( .A(n2479), .B(n2499), .Z(n2784) );
  COND2X1 U2419 ( .A(n2785), .B(n2523), .C(n2443), .D(n2786), .Z(n1451) );
  CENX1 U2420 ( .A(n2479), .B(n2498), .Z(n2785) );
  COND2X1 U2421 ( .A(n2786), .B(n2523), .C(n2443), .D(n2787), .Z(n1450) );
  CENX1 U2422 ( .A(n2479), .B(n2497), .Z(n2786) );
  COND2X1 U2423 ( .A(n2787), .B(n2523), .C(n2443), .D(n2788), .Z(n1449) );
  CENX1 U2424 ( .A(n2479), .B(n2496), .Z(n2787) );
  COND2X1 U2425 ( .A(n2788), .B(n2523), .C(n2443), .D(n2789), .Z(n1448) );
  CENX1 U2426 ( .A(n2479), .B(n2495), .Z(n2788) );
  COND2X1 U2427 ( .A(n2789), .B(n2523), .C(n2443), .D(n2790), .Z(n1447) );
  CENX1 U2428 ( .A(n2479), .B(n2494), .Z(n2789) );
  COND2X1 U2429 ( .A(n2790), .B(n2523), .C(n2443), .D(n2791), .Z(n1446) );
  CENX1 U2430 ( .A(n2479), .B(n2493), .Z(n2790) );
  COND2X1 U2431 ( .A(n2791), .B(n2523), .C(n2443), .D(n2546), .Z(n1445) );
  CEOX1 U2432 ( .A(n2479), .B(b[30]), .Z(n2546) );
  CENX1 U2433 ( .A(n2479), .B(n2492), .Z(n2791) );
  CAOR1X1 U2434 ( .A(n2523), .B(n2443), .C(n2547), .Z(n1444) );
  CEOX1 U2435 ( .A(n2479), .B(b[31]), .Z(n2547) );
  CNR2X1 U2436 ( .A(n2444), .B(n2515), .Z(n1443) );
  COND2X1 U2437 ( .A(n2792), .B(n2549), .C(n2444), .D(n2793), .Z(n1442) );
  CENX1 U2438 ( .A(n2515), .B(n2477), .Z(n2792) );
  COND2X1 U2439 ( .A(n2793), .B(n2549), .C(n2444), .D(n2794), .Z(n1441) );
  CENX1 U2440 ( .A(n2477), .B(n2453), .Z(n2793) );
  COND2X1 U2441 ( .A(n2794), .B(n2549), .C(n2444), .D(n2795), .Z(n1440) );
  CENX1 U2442 ( .A(n2477), .B(n2454), .Z(n2794) );
  COND2X1 U2443 ( .A(n2795), .B(n2549), .C(n2444), .D(n2796), .Z(n1439) );
  CENX1 U2444 ( .A(n2477), .B(n2455), .Z(n2795) );
  COND2X1 U2445 ( .A(n2796), .B(n2549), .C(n2444), .D(n2797), .Z(n1438) );
  CENX1 U2446 ( .A(n2477), .B(n2456), .Z(n2796) );
  COND2X1 U2447 ( .A(n2797), .B(n2549), .C(n2444), .D(n2798), .Z(n1437) );
  CENX1 U2448 ( .A(n2477), .B(n2457), .Z(n2797) );
  COND2X1 U2449 ( .A(n2798), .B(n2549), .C(n2444), .D(n2799), .Z(n1436) );
  CENX1 U2450 ( .A(n2477), .B(n2458), .Z(n2798) );
  COND2X1 U2451 ( .A(n2799), .B(n2549), .C(n2444), .D(n2800), .Z(n1435) );
  CENX1 U2452 ( .A(n2477), .B(n2514), .Z(n2799) );
  COND2X1 U2453 ( .A(n2800), .B(n2549), .C(n2444), .D(n2801), .Z(n1434) );
  CENX1 U2454 ( .A(n2477), .B(n2513), .Z(n2800) );
  COND2X1 U2455 ( .A(n2801), .B(n2549), .C(n2444), .D(n2802), .Z(n1433) );
  CENX1 U2456 ( .A(n2477), .B(n2512), .Z(n2801) );
  COND2X1 U2457 ( .A(n2802), .B(n2549), .C(n2444), .D(n2803), .Z(n1432) );
  CENX1 U2458 ( .A(n2477), .B(n2511), .Z(n2802) );
  COND2X1 U2459 ( .A(n2803), .B(n2549), .C(n2444), .D(n2804), .Z(n1431) );
  CENX1 U2460 ( .A(n2477), .B(n2510), .Z(n2803) );
  COND2X1 U2461 ( .A(n2804), .B(n2549), .C(n2444), .D(n2805), .Z(n1430) );
  CENX1 U2462 ( .A(n2477), .B(n2509), .Z(n2804) );
  COND2X1 U2463 ( .A(n2805), .B(n2549), .C(n2444), .D(n2806), .Z(n1429) );
  CENX1 U2464 ( .A(n2477), .B(n2508), .Z(n2805) );
  COND2X1 U2465 ( .A(n2806), .B(n2549), .C(n2444), .D(n2807), .Z(n1428) );
  CENX1 U2466 ( .A(n2477), .B(n2507), .Z(n2806) );
  COND2X1 U2467 ( .A(n2807), .B(n2549), .C(n2444), .D(n2808), .Z(n1427) );
  CENX1 U2468 ( .A(n2477), .B(n2506), .Z(n2807) );
  COND2X1 U2469 ( .A(n2808), .B(n2549), .C(n2444), .D(n2809), .Z(n1426) );
  CENX1 U2470 ( .A(n2477), .B(n2505), .Z(n2808) );
  COND2X1 U2471 ( .A(n2809), .B(n2549), .C(n2444), .D(n2810), .Z(n1425) );
  CENX1 U2472 ( .A(n2477), .B(n2504), .Z(n2809) );
  COND2X1 U2473 ( .A(n2810), .B(n2549), .C(n2444), .D(n2811), .Z(n1424) );
  CENX1 U2474 ( .A(n2477), .B(n2503), .Z(n2810) );
  COND2X1 U2475 ( .A(n2811), .B(n2549), .C(n2444), .D(n2812), .Z(n1423) );
  CENX1 U2476 ( .A(n2477), .B(n2502), .Z(n2811) );
  COND2X1 U2477 ( .A(n2812), .B(n2549), .C(n2444), .D(n2813), .Z(n1422) );
  CENX1 U2478 ( .A(n2477), .B(n2501), .Z(n2812) );
  COND2X1 U2479 ( .A(n2813), .B(n2549), .C(n2444), .D(n2814), .Z(n1421) );
  CENX1 U2480 ( .A(n2477), .B(n2500), .Z(n2813) );
  COND2X1 U2481 ( .A(n2814), .B(n2549), .C(n2444), .D(n2815), .Z(n1420) );
  CENX1 U2482 ( .A(n2477), .B(n2499), .Z(n2814) );
  COND2X1 U2483 ( .A(n2815), .B(n2549), .C(n2444), .D(n2816), .Z(n1419) );
  CENX1 U2484 ( .A(n2477), .B(n2498), .Z(n2815) );
  COND2X1 U2485 ( .A(n2816), .B(n2549), .C(n2444), .D(n2817), .Z(n1418) );
  CENX1 U2486 ( .A(n2477), .B(n2497), .Z(n2816) );
  COND2X1 U2487 ( .A(n2817), .B(n2549), .C(n2444), .D(n2818), .Z(n1417) );
  CENX1 U2488 ( .A(n2477), .B(n2496), .Z(n2817) );
  COND2X1 U2489 ( .A(n2818), .B(n2549), .C(n2444), .D(n2819), .Z(n1416) );
  CENX1 U2490 ( .A(n2477), .B(n2495), .Z(n2818) );
  COND2X1 U2491 ( .A(n2819), .B(n2549), .C(n2444), .D(n2820), .Z(n1415) );
  CENX1 U2492 ( .A(n2477), .B(n2494), .Z(n2819) );
  COND2X1 U2493 ( .A(n2820), .B(n2549), .C(n2444), .D(n2821), .Z(n1414) );
  CENX1 U2494 ( .A(n2477), .B(n2493), .Z(n2820) );
  COND2X1 U2495 ( .A(n2821), .B(n2549), .C(n2444), .D(n2548), .Z(n1413) );
  CEOX1 U2496 ( .A(n2477), .B(b[30]), .Z(n2548) );
  CENX1 U2497 ( .A(n2477), .B(n2492), .Z(n2821) );
  CAOR1X1 U2498 ( .A(n2549), .B(n2444), .C(n2551), .Z(n1412) );
  CEOX1 U2499 ( .A(n2477), .B(b[31]), .Z(n2551) );
  CNR2X1 U2500 ( .A(n2445), .B(n2515), .Z(n1411) );
  COND2X1 U2501 ( .A(n2822), .B(n2553), .C(n2445), .D(n2823), .Z(n1410) );
  CENX1 U2502 ( .A(n2515), .B(n2475), .Z(n2822) );
  COND2X1 U2503 ( .A(n2823), .B(n2553), .C(n2445), .D(n2824), .Z(n1409) );
  CENX1 U2504 ( .A(n2475), .B(n2453), .Z(n2823) );
  COND2X1 U2505 ( .A(n2824), .B(n2553), .C(n2445), .D(n2825), .Z(n1408) );
  CENX1 U2506 ( .A(n2475), .B(n2454), .Z(n2824) );
  COND2X1 U2507 ( .A(n2825), .B(n2553), .C(n2445), .D(n2826), .Z(n1407) );
  CENX1 U2508 ( .A(n2475), .B(n2455), .Z(n2825) );
  COND2X1 U2509 ( .A(n2826), .B(n2553), .C(n2445), .D(n2827), .Z(n1406) );
  CENX1 U2510 ( .A(n2475), .B(n2456), .Z(n2826) );
  COND2X1 U2511 ( .A(n2827), .B(n2553), .C(n2445), .D(n2828), .Z(n1405) );
  CENX1 U2512 ( .A(n2475), .B(n2457), .Z(n2827) );
  COND2X1 U2513 ( .A(n2828), .B(n2553), .C(n2445), .D(n2829), .Z(n1404) );
  CENX1 U2514 ( .A(n2475), .B(n2458), .Z(n2828) );
  COND2X1 U2515 ( .A(n2829), .B(n2553), .C(n2445), .D(n2830), .Z(n1403) );
  CENX1 U2516 ( .A(n2475), .B(n2514), .Z(n2829) );
  COND2X1 U2517 ( .A(n2830), .B(n2553), .C(n2445), .D(n2831), .Z(n1402) );
  CENX1 U2518 ( .A(n2475), .B(n2513), .Z(n2830) );
  COND2X1 U2519 ( .A(n2831), .B(n2553), .C(n2445), .D(n2832), .Z(n1401) );
  CENX1 U2520 ( .A(n2475), .B(n2512), .Z(n2831) );
  COND2X1 U2521 ( .A(n2832), .B(n2553), .C(n2445), .D(n2833), .Z(n1400) );
  CENX1 U2522 ( .A(n2475), .B(n2511), .Z(n2832) );
  COND2X1 U2523 ( .A(n2833), .B(n2553), .C(n2445), .D(n2834), .Z(n1399) );
  CENX1 U2524 ( .A(n2475), .B(n2510), .Z(n2833) );
  COND2X1 U2525 ( .A(n2834), .B(n2553), .C(n2445), .D(n2835), .Z(n1398) );
  CENX1 U2526 ( .A(n2475), .B(n2509), .Z(n2834) );
  COND2X1 U2527 ( .A(n2835), .B(n2553), .C(n2445), .D(n2836), .Z(n1397) );
  CENX1 U2528 ( .A(n2475), .B(n2508), .Z(n2835) );
  COND2X1 U2529 ( .A(n2836), .B(n2553), .C(n2445), .D(n2837), .Z(n1396) );
  CENX1 U2530 ( .A(n2475), .B(n2507), .Z(n2836) );
  COND2X1 U2531 ( .A(n2837), .B(n2553), .C(n2445), .D(n2838), .Z(n1395) );
  CENX1 U2532 ( .A(n2475), .B(n2506), .Z(n2837) );
  COND2X1 U2533 ( .A(n2838), .B(n2553), .C(n2445), .D(n2839), .Z(n1394) );
  CENX1 U2534 ( .A(n2475), .B(n2505), .Z(n2838) );
  COND2X1 U2535 ( .A(n2839), .B(n2553), .C(n2445), .D(n2840), .Z(n1393) );
  CENX1 U2536 ( .A(n2475), .B(n2504), .Z(n2839) );
  COND2X1 U2537 ( .A(n2840), .B(n2553), .C(n2445), .D(n2841), .Z(n1392) );
  CENX1 U2538 ( .A(n2475), .B(n2503), .Z(n2840) );
  COND2X1 U2539 ( .A(n2841), .B(n2553), .C(n2445), .D(n2842), .Z(n1391) );
  CENX1 U2540 ( .A(n2475), .B(n2502), .Z(n2841) );
  COND2X1 U2541 ( .A(n2842), .B(n2553), .C(n2445), .D(n2843), .Z(n1390) );
  CENX1 U2542 ( .A(n2475), .B(n2501), .Z(n2842) );
  COND2X1 U2543 ( .A(n2843), .B(n2553), .C(n2445), .D(n2844), .Z(n1389) );
  CENX1 U2544 ( .A(n2475), .B(n2500), .Z(n2843) );
  COND2X1 U2545 ( .A(n2844), .B(n2553), .C(n2445), .D(n2845), .Z(n1388) );
  CENX1 U2546 ( .A(n2475), .B(n2499), .Z(n2844) );
  COND2X1 U2547 ( .A(n2845), .B(n2553), .C(n2445), .D(n2846), .Z(n1387) );
  CENX1 U2548 ( .A(n2475), .B(n2498), .Z(n2845) );
  COND2X1 U2549 ( .A(n2846), .B(n2553), .C(n2445), .D(n2847), .Z(n1386) );
  CENX1 U2550 ( .A(n2475), .B(n2497), .Z(n2846) );
  COND2X1 U2551 ( .A(n2847), .B(n2553), .C(n2445), .D(n2848), .Z(n1385) );
  CENX1 U2552 ( .A(n2475), .B(n2496), .Z(n2847) );
  COND2X1 U2553 ( .A(n2848), .B(n2553), .C(n2445), .D(n2849), .Z(n1384) );
  CENX1 U2554 ( .A(n2475), .B(n2495), .Z(n2848) );
  COND2X1 U2555 ( .A(n2849), .B(n2553), .C(n2445), .D(n2850), .Z(n1383) );
  CENX1 U2556 ( .A(n2475), .B(n2494), .Z(n2849) );
  COND2X1 U2557 ( .A(n2850), .B(n2553), .C(n2445), .D(n2851), .Z(n1382) );
  CENX1 U2558 ( .A(n2475), .B(n2493), .Z(n2850) );
  COND2X1 U2559 ( .A(n2851), .B(n2553), .C(n2445), .D(n2552), .Z(n1381) );
  CEOX1 U2560 ( .A(n2475), .B(b[30]), .Z(n2552) );
  CENX1 U2561 ( .A(n2475), .B(n2492), .Z(n2851) );
  CAOR1X1 U2562 ( .A(n2553), .B(n2445), .C(n2555), .Z(n1380) );
  CEOX1 U2563 ( .A(n2475), .B(b[31]), .Z(n2555) );
  CNR2X1 U2564 ( .A(n2446), .B(n2515), .Z(n1379) );
  COND2X1 U2565 ( .A(n2852), .B(n2557), .C(n2446), .D(n2853), .Z(n1378) );
  CENX1 U2566 ( .A(n2515), .B(n2473), .Z(n2852) );
  COND2X1 U2567 ( .A(n2853), .B(n2557), .C(n2446), .D(n2854), .Z(n1377) );
  CENX1 U2568 ( .A(n2473), .B(n2453), .Z(n2853) );
  COND2X1 U2569 ( .A(n2854), .B(n2557), .C(n2446), .D(n2855), .Z(n1376) );
  CENX1 U2570 ( .A(n2473), .B(n2454), .Z(n2854) );
  COND2X1 U2571 ( .A(n2855), .B(n2557), .C(n2446), .D(n2856), .Z(n1375) );
  CENX1 U2572 ( .A(n2473), .B(n2455), .Z(n2855) );
  COND2X1 U2573 ( .A(n2856), .B(n2557), .C(n2446), .D(n2857), .Z(n1374) );
  CENX1 U2574 ( .A(n2473), .B(n2456), .Z(n2856) );
  COND2X1 U2575 ( .A(n2857), .B(n2557), .C(n2446), .D(n2858), .Z(n1373) );
  CENX1 U2576 ( .A(n2473), .B(n2457), .Z(n2857) );
  COND2X1 U2577 ( .A(n2858), .B(n2557), .C(n2446), .D(n2859), .Z(n1372) );
  CENX1 U2578 ( .A(n2473), .B(n2458), .Z(n2858) );
  COND2X1 U2579 ( .A(n2859), .B(n2557), .C(n2446), .D(n2860), .Z(n1371) );
  CENX1 U2580 ( .A(n2473), .B(n2514), .Z(n2859) );
  COND2X1 U2581 ( .A(n2860), .B(n2557), .C(n2446), .D(n2861), .Z(n1370) );
  CENX1 U2582 ( .A(n2473), .B(n2513), .Z(n2860) );
  COND2X1 U2583 ( .A(n2861), .B(n2557), .C(n2446), .D(n2862), .Z(n1369) );
  CENX1 U2584 ( .A(n2473), .B(n2512), .Z(n2861) );
  COND2X1 U2585 ( .A(n2862), .B(n2557), .C(n2446), .D(n2863), .Z(n1368) );
  CENX1 U2586 ( .A(n2473), .B(n2511), .Z(n2862) );
  COND2X1 U2587 ( .A(n2863), .B(n2557), .C(n2446), .D(n2864), .Z(n1367) );
  CENX1 U2588 ( .A(n2473), .B(n2510), .Z(n2863) );
  COND2X1 U2589 ( .A(n2864), .B(n2557), .C(n2446), .D(n2865), .Z(n1366) );
  CENX1 U2590 ( .A(n2473), .B(n2509), .Z(n2864) );
  COND2X1 U2591 ( .A(n2865), .B(n2557), .C(n2446), .D(n2866), .Z(n1365) );
  CENX1 U2592 ( .A(n2473), .B(n2508), .Z(n2865) );
  COND2X1 U2593 ( .A(n2866), .B(n2557), .C(n2446), .D(n2867), .Z(n1364) );
  CENX1 U2594 ( .A(n2473), .B(n2507), .Z(n2866) );
  COND2X1 U2595 ( .A(n2867), .B(n2557), .C(n2446), .D(n2868), .Z(n1363) );
  CENX1 U2596 ( .A(n2473), .B(n2506), .Z(n2867) );
  COND2X1 U2597 ( .A(n2868), .B(n2557), .C(n2446), .D(n2869), .Z(n1362) );
  CENX1 U2598 ( .A(n2473), .B(n2505), .Z(n2868) );
  COND2X1 U2599 ( .A(n2869), .B(n2557), .C(n2446), .D(n2870), .Z(n1361) );
  CENX1 U2600 ( .A(n2473), .B(n2504), .Z(n2869) );
  COND2X1 U2601 ( .A(n2870), .B(n2557), .C(n2446), .D(n2871), .Z(n1360) );
  CENX1 U2602 ( .A(n2473), .B(n2503), .Z(n2870) );
  COND2X1 U2603 ( .A(n2871), .B(n2557), .C(n2446), .D(n2872), .Z(n1359) );
  CENX1 U2604 ( .A(n2473), .B(n2502), .Z(n2871) );
  COND2X1 U2605 ( .A(n2872), .B(n2557), .C(n2446), .D(n2873), .Z(n1358) );
  CENX1 U2606 ( .A(n2473), .B(n2501), .Z(n2872) );
  COND2X1 U2607 ( .A(n2873), .B(n2557), .C(n2446), .D(n2874), .Z(n1357) );
  CENX1 U2608 ( .A(n2473), .B(n2500), .Z(n2873) );
  COND2X1 U2609 ( .A(n2874), .B(n2557), .C(n2446), .D(n2875), .Z(n1356) );
  CENX1 U2610 ( .A(n2473), .B(n2499), .Z(n2874) );
  COND2X1 U2611 ( .A(n2875), .B(n2557), .C(n2446), .D(n2876), .Z(n1355) );
  CENX1 U2612 ( .A(n2473), .B(n2498), .Z(n2875) );
  COND2X1 U2613 ( .A(n2876), .B(n2557), .C(n2446), .D(n2877), .Z(n1354) );
  CENX1 U2614 ( .A(n2473), .B(n2497), .Z(n2876) );
  COND2X1 U2615 ( .A(n2877), .B(n2557), .C(n2446), .D(n2878), .Z(n1353) );
  CENX1 U2616 ( .A(n2473), .B(n2496), .Z(n2877) );
  COND2X1 U2617 ( .A(n2878), .B(n2557), .C(n2446), .D(n2879), .Z(n1352) );
  CENX1 U2618 ( .A(n2473), .B(n2495), .Z(n2878) );
  COND2X1 U2619 ( .A(n2879), .B(n2557), .C(n2446), .D(n2880), .Z(n1351) );
  CENX1 U2620 ( .A(n2473), .B(n2494), .Z(n2879) );
  COND2X1 U2621 ( .A(n2880), .B(n2557), .C(n2446), .D(n2881), .Z(n1350) );
  CENX1 U2622 ( .A(n2473), .B(n2493), .Z(n2880) );
  COND2X1 U2623 ( .A(n2881), .B(n2557), .C(n2446), .D(n2556), .Z(n1349) );
  CEOX1 U2624 ( .A(n2473), .B(b[30]), .Z(n2556) );
  CENX1 U2625 ( .A(n2473), .B(n2492), .Z(n2881) );
  CAOR1X1 U2626 ( .A(n2557), .B(n2446), .C(n2559), .Z(n1348) );
  CEOX1 U2627 ( .A(n2473), .B(b[31]), .Z(n2559) );
  CNR2X1 U2628 ( .A(n2447), .B(n2515), .Z(n1347) );
  COND2X1 U2629 ( .A(n2882), .B(n2561), .C(n2447), .D(n2883), .Z(n1346) );
  CENX1 U2630 ( .A(n2515), .B(n2471), .Z(n2882) );
  COND2X1 U2631 ( .A(n2883), .B(n2561), .C(n2447), .D(n2884), .Z(n1345) );
  CENX1 U2632 ( .A(n2471), .B(n2453), .Z(n2883) );
  COND2X1 U2633 ( .A(n2884), .B(n2561), .C(n2447), .D(n2885), .Z(n1344) );
  CENX1 U2634 ( .A(n2471), .B(n2454), .Z(n2884) );
  COND2X1 U2635 ( .A(n2885), .B(n2561), .C(n2447), .D(n2886), .Z(n1343) );
  CENX1 U2636 ( .A(n2471), .B(n2455), .Z(n2885) );
  COND2X1 U2637 ( .A(n2886), .B(n2561), .C(n2447), .D(n2887), .Z(n1342) );
  CENX1 U2638 ( .A(n2471), .B(n2456), .Z(n2886) );
  COND2X1 U2639 ( .A(n2887), .B(n2561), .C(n2447), .D(n2888), .Z(n1341) );
  CENX1 U2640 ( .A(n2471), .B(n2457), .Z(n2887) );
  COND2X1 U2641 ( .A(n2888), .B(n2561), .C(n2447), .D(n2889), .Z(n1340) );
  CENX1 U2642 ( .A(n2471), .B(n2458), .Z(n2888) );
  COND2X1 U2643 ( .A(n2889), .B(n2561), .C(n2447), .D(n2890), .Z(n1339) );
  CENX1 U2644 ( .A(n2471), .B(n2514), .Z(n2889) );
  COND2X1 U2645 ( .A(n2890), .B(n2561), .C(n2447), .D(n2891), .Z(n1338) );
  CENX1 U2646 ( .A(n2471), .B(n2513), .Z(n2890) );
  COND2X1 U2647 ( .A(n2891), .B(n2561), .C(n2447), .D(n2892), .Z(n1337) );
  CENX1 U2648 ( .A(n2471), .B(n2512), .Z(n2891) );
  COND2X1 U2649 ( .A(n2892), .B(n2561), .C(n2447), .D(n2893), .Z(n1336) );
  CENX1 U2650 ( .A(n2471), .B(n2511), .Z(n2892) );
  COND2X1 U2651 ( .A(n2893), .B(n2561), .C(n2447), .D(n2894), .Z(n1335) );
  CENX1 U2652 ( .A(n2471), .B(n2510), .Z(n2893) );
  COND2X1 U2653 ( .A(n2894), .B(n2561), .C(n2447), .D(n2895), .Z(n1334) );
  CENX1 U2654 ( .A(n2471), .B(n2509), .Z(n2894) );
  COND2X1 U2655 ( .A(n2895), .B(n2561), .C(n2447), .D(n2896), .Z(n1333) );
  CENX1 U2656 ( .A(n2471), .B(n2508), .Z(n2895) );
  COND2X1 U2657 ( .A(n2896), .B(n2561), .C(n2447), .D(n2897), .Z(n1332) );
  CENX1 U2658 ( .A(n2471), .B(n2507), .Z(n2896) );
  COND2X1 U2659 ( .A(n2897), .B(n2561), .C(n2447), .D(n2898), .Z(n1331) );
  CENX1 U2660 ( .A(n2471), .B(n2506), .Z(n2897) );
  COND2X1 U2661 ( .A(n2898), .B(n2561), .C(n2447), .D(n2899), .Z(n1330) );
  CENX1 U2662 ( .A(n2471), .B(n2505), .Z(n2898) );
  COND2X1 U2663 ( .A(n2899), .B(n2561), .C(n2447), .D(n2900), .Z(n1329) );
  CENX1 U2664 ( .A(n2471), .B(n2504), .Z(n2899) );
  COND2X1 U2665 ( .A(n2900), .B(n2561), .C(n2447), .D(n2901), .Z(n1328) );
  CENX1 U2666 ( .A(n2471), .B(n2503), .Z(n2900) );
  COND2X1 U2667 ( .A(n2901), .B(n2561), .C(n2447), .D(n2902), .Z(n1327) );
  CENX1 U2668 ( .A(n2471), .B(n2502), .Z(n2901) );
  COND2X1 U2669 ( .A(n2902), .B(n2561), .C(n2447), .D(n2903), .Z(n1326) );
  CENX1 U2670 ( .A(n2471), .B(n2501), .Z(n2902) );
  COND2X1 U2671 ( .A(n2903), .B(n2561), .C(n2447), .D(n2904), .Z(n1325) );
  CENX1 U2672 ( .A(n2471), .B(n2500), .Z(n2903) );
  COND2X1 U2673 ( .A(n2904), .B(n2561), .C(n2447), .D(n2905), .Z(n1324) );
  CENX1 U2674 ( .A(n2471), .B(n2499), .Z(n2904) );
  COND2X1 U2675 ( .A(n2905), .B(n2561), .C(n2447), .D(n2906), .Z(n1323) );
  CENX1 U2676 ( .A(n2471), .B(n2498), .Z(n2905) );
  COND2X1 U2677 ( .A(n2906), .B(n2561), .C(n2447), .D(n2907), .Z(n1322) );
  CENX1 U2678 ( .A(n2471), .B(n2497), .Z(n2906) );
  COND2X1 U2679 ( .A(n2907), .B(n2561), .C(n2447), .D(n2908), .Z(n1321) );
  CENX1 U2680 ( .A(n2471), .B(n2496), .Z(n2907) );
  COND2X1 U2681 ( .A(n2908), .B(n2561), .C(n2447), .D(n2909), .Z(n1320) );
  CENX1 U2682 ( .A(n2471), .B(n2495), .Z(n2908) );
  COND2X1 U2683 ( .A(n2909), .B(n2561), .C(n2447), .D(n2910), .Z(n1319) );
  CENX1 U2684 ( .A(n2471), .B(n2494), .Z(n2909) );
  COND2X1 U2685 ( .A(n2910), .B(n2561), .C(n2447), .D(n2911), .Z(n1318) );
  CENX1 U2686 ( .A(n2471), .B(n2493), .Z(n2910) );
  COND2X1 U2687 ( .A(n2911), .B(n2561), .C(n2447), .D(n2560), .Z(n1317) );
  CEOX1 U2688 ( .A(n2471), .B(b[30]), .Z(n2560) );
  CENX1 U2689 ( .A(n2471), .B(n2492), .Z(n2911) );
  CAOR1X1 U2690 ( .A(n2561), .B(n2447), .C(n2563), .Z(n1316) );
  CEOX1 U2691 ( .A(n2471), .B(b[31]), .Z(n2563) );
  CNR2X1 U2692 ( .A(n2448), .B(n2515), .Z(n1315) );
  COND2X1 U2693 ( .A(n2912), .B(n2565), .C(n2448), .D(n2913), .Z(n1314) );
  CENX1 U2694 ( .A(n2515), .B(n2469), .Z(n2912) );
  COND2X1 U2695 ( .A(n2913), .B(n2565), .C(n2448), .D(n2914), .Z(n1313) );
  CENX1 U2696 ( .A(n2469), .B(n2453), .Z(n2913) );
  COND2X1 U2697 ( .A(n2914), .B(n2565), .C(n2448), .D(n2915), .Z(n1312) );
  CENX1 U2698 ( .A(n2469), .B(n2454), .Z(n2914) );
  COND2X1 U2699 ( .A(n2915), .B(n2565), .C(n2448), .D(n2916), .Z(n1311) );
  CENX1 U2700 ( .A(n2469), .B(n2455), .Z(n2915) );
  COND2X1 U2701 ( .A(n2916), .B(n2565), .C(n2448), .D(n2917), .Z(n1310) );
  CENX1 U2702 ( .A(n2469), .B(n2456), .Z(n2916) );
  COND2X1 U2703 ( .A(n2917), .B(n2565), .C(n2448), .D(n2918), .Z(n1309) );
  CENX1 U2704 ( .A(n2469), .B(n2457), .Z(n2917) );
  COND2X1 U2705 ( .A(n2918), .B(n2565), .C(n2448), .D(n2919), .Z(n1308) );
  CENX1 U2706 ( .A(n2469), .B(n2458), .Z(n2918) );
  COND2X1 U2707 ( .A(n2919), .B(n2565), .C(n2448), .D(n2920), .Z(n1307) );
  CENX1 U2708 ( .A(n2469), .B(n2514), .Z(n2919) );
  COND2X1 U2709 ( .A(n2920), .B(n2565), .C(n2448), .D(n2921), .Z(n1306) );
  CENX1 U2710 ( .A(n2469), .B(n2513), .Z(n2920) );
  COND2X1 U2711 ( .A(n2921), .B(n2565), .C(n2448), .D(n2922), .Z(n1305) );
  CENX1 U2712 ( .A(n2469), .B(n2512), .Z(n2921) );
  COND2X1 U2713 ( .A(n2922), .B(n2565), .C(n2448), .D(n2923), .Z(n1304) );
  CENX1 U2714 ( .A(n2469), .B(n2511), .Z(n2922) );
  COND2X1 U2715 ( .A(n2923), .B(n2565), .C(n2448), .D(n2924), .Z(n1303) );
  CENX1 U2716 ( .A(n2469), .B(n2510), .Z(n2923) );
  COND2X1 U2717 ( .A(n2924), .B(n2565), .C(n2448), .D(n2925), .Z(n1302) );
  CENX1 U2718 ( .A(n2469), .B(n2509), .Z(n2924) );
  COND2X1 U2719 ( .A(n2925), .B(n2565), .C(n2448), .D(n2926), .Z(n1301) );
  CENX1 U2720 ( .A(n2469), .B(n2508), .Z(n2925) );
  COND2X1 U2721 ( .A(n2926), .B(n2565), .C(n2448), .D(n2927), .Z(n1300) );
  CENX1 U2722 ( .A(n2469), .B(n2507), .Z(n2926) );
  COND2X1 U2723 ( .A(n2927), .B(n2565), .C(n2448), .D(n2928), .Z(n1299) );
  CENX1 U2724 ( .A(n2469), .B(n2506), .Z(n2927) );
  COND2X1 U2725 ( .A(n2928), .B(n2565), .C(n2448), .D(n2929), .Z(n1298) );
  CENX1 U2726 ( .A(n2469), .B(n2505), .Z(n2928) );
  COND2X1 U2727 ( .A(n2929), .B(n2565), .C(n2448), .D(n2930), .Z(n1297) );
  CENX1 U2728 ( .A(n2469), .B(n2504), .Z(n2929) );
  COND2X1 U2729 ( .A(n2930), .B(n2565), .C(n2448), .D(n2931), .Z(n1296) );
  CENX1 U2730 ( .A(n2469), .B(n2503), .Z(n2930) );
  COND2X1 U2731 ( .A(n2931), .B(n2565), .C(n2448), .D(n2932), .Z(n1295) );
  CENX1 U2732 ( .A(n2469), .B(n2502), .Z(n2931) );
  COND2X1 U2733 ( .A(n2932), .B(n2565), .C(n2448), .D(n2933), .Z(n1294) );
  CENX1 U2734 ( .A(n2469), .B(n2501), .Z(n2932) );
  COND2X1 U2735 ( .A(n2933), .B(n2565), .C(n2448), .D(n2934), .Z(n1293) );
  CENX1 U2736 ( .A(n2469), .B(n2500), .Z(n2933) );
  COND2X1 U2737 ( .A(n2934), .B(n2565), .C(n2448), .D(n2935), .Z(n1292) );
  CENX1 U2738 ( .A(n2469), .B(n2499), .Z(n2934) );
  COND2X1 U2739 ( .A(n2935), .B(n2565), .C(n2448), .D(n2936), .Z(n1291) );
  CENX1 U2740 ( .A(n2469), .B(n2498), .Z(n2935) );
  COND2X1 U2741 ( .A(n2936), .B(n2565), .C(n2448), .D(n2937), .Z(n1290) );
  CENX1 U2742 ( .A(n2469), .B(n2497), .Z(n2936) );
  COND2X1 U2743 ( .A(n2937), .B(n2565), .C(n2448), .D(n2938), .Z(n1289) );
  CENX1 U2744 ( .A(n2469), .B(n2496), .Z(n2937) );
  COND2X1 U2745 ( .A(n2938), .B(n2565), .C(n2448), .D(n2939), .Z(n1288) );
  CENX1 U2746 ( .A(n2469), .B(n2495), .Z(n2938) );
  COND2X1 U2747 ( .A(n2939), .B(n2565), .C(n2448), .D(n2940), .Z(n1287) );
  CENX1 U2748 ( .A(n2469), .B(n2494), .Z(n2939) );
  COND2X1 U2749 ( .A(n2940), .B(n2565), .C(n2448), .D(n2941), .Z(n1286) );
  CENX1 U2750 ( .A(n2469), .B(n2493), .Z(n2940) );
  COND2X1 U2751 ( .A(n2941), .B(n2565), .C(n2448), .D(n2564), .Z(n1285) );
  CEOX1 U2752 ( .A(n2469), .B(b[30]), .Z(n2564) );
  CENX1 U2753 ( .A(n2469), .B(n2492), .Z(n2941) );
  CAOR1X1 U2754 ( .A(n2565), .B(n2448), .C(n2567), .Z(n1284) );
  CEOX1 U2755 ( .A(n2469), .B(b[31]), .Z(n2567) );
  CNR2X1 U2756 ( .A(n2449), .B(n2515), .Z(n1283) );
  COND2X1 U2757 ( .A(n2942), .B(n2569), .C(n2449), .D(n2943), .Z(n1282) );
  CENX1 U2758 ( .A(n2515), .B(n2467), .Z(n2942) );
  COND2X1 U2759 ( .A(n2943), .B(n2569), .C(n2449), .D(n2944), .Z(n1281) );
  CENX1 U2760 ( .A(n2467), .B(n2453), .Z(n2943) );
  COND2X1 U2761 ( .A(n2944), .B(n2569), .C(n2449), .D(n2945), .Z(n1280) );
  CENX1 U2762 ( .A(n2467), .B(n2454), .Z(n2944) );
  COND2X1 U2763 ( .A(n2945), .B(n2569), .C(n2449), .D(n2946), .Z(n1279) );
  CENX1 U2764 ( .A(n2467), .B(n2455), .Z(n2945) );
  COND2X1 U2765 ( .A(n2946), .B(n2569), .C(n2449), .D(n2947), .Z(n1278) );
  CENX1 U2766 ( .A(n2467), .B(n2456), .Z(n2946) );
  COND2X1 U2767 ( .A(n2947), .B(n2569), .C(n2449), .D(n2948), .Z(n1277) );
  CENX1 U2768 ( .A(n2467), .B(n2457), .Z(n2947) );
  COND2X1 U2769 ( .A(n2948), .B(n2569), .C(n2449), .D(n2949), .Z(n1276) );
  CENX1 U2770 ( .A(n2467), .B(n2458), .Z(n2948) );
  COND2X1 U2771 ( .A(n2949), .B(n2569), .C(n2449), .D(n2950), .Z(n1275) );
  CENX1 U2772 ( .A(n2467), .B(n2514), .Z(n2949) );
  COND2X1 U2773 ( .A(n2950), .B(n2569), .C(n2449), .D(n2951), .Z(n1274) );
  CENX1 U2774 ( .A(n2467), .B(n2513), .Z(n2950) );
  COND2X1 U2775 ( .A(n2951), .B(n2569), .C(n2449), .D(n2952), .Z(n1273) );
  CENX1 U2776 ( .A(n2467), .B(n2512), .Z(n2951) );
  COND2X1 U2777 ( .A(n2952), .B(n2569), .C(n2449), .D(n2953), .Z(n1272) );
  CENX1 U2778 ( .A(n2467), .B(n2511), .Z(n2952) );
  COND2X1 U2779 ( .A(n2953), .B(n2569), .C(n2449), .D(n2954), .Z(n1271) );
  CENX1 U2780 ( .A(n2467), .B(n2510), .Z(n2953) );
  COND2X1 U2781 ( .A(n2954), .B(n2569), .C(n2449), .D(n2955), .Z(n1270) );
  CENX1 U2782 ( .A(n2467), .B(n2509), .Z(n2954) );
  COND2X1 U2783 ( .A(n2955), .B(n2569), .C(n2449), .D(n2956), .Z(n1269) );
  CENX1 U2784 ( .A(n2467), .B(n2508), .Z(n2955) );
  COND2X1 U2785 ( .A(n2956), .B(n2569), .C(n2449), .D(n2957), .Z(n1268) );
  CENX1 U2786 ( .A(n2467), .B(n2507), .Z(n2956) );
  COND2X1 U2787 ( .A(n2957), .B(n2569), .C(n2449), .D(n2958), .Z(n1267) );
  CENX1 U2788 ( .A(n2467), .B(n2506), .Z(n2957) );
  COND2X1 U2789 ( .A(n2958), .B(n2569), .C(n2449), .D(n2959), .Z(n1266) );
  CENX1 U2790 ( .A(n2467), .B(n2505), .Z(n2958) );
  COND2X1 U2791 ( .A(n2959), .B(n2569), .C(n2449), .D(n2960), .Z(n1265) );
  CENX1 U2792 ( .A(n2467), .B(n2504), .Z(n2959) );
  COND2X1 U2793 ( .A(n2960), .B(n2569), .C(n2449), .D(n2961), .Z(n1264) );
  CENX1 U2794 ( .A(n2467), .B(n2503), .Z(n2960) );
  COND2X1 U2795 ( .A(n2961), .B(n2569), .C(n2449), .D(n2962), .Z(n1263) );
  CENX1 U2796 ( .A(n2467), .B(n2502), .Z(n2961) );
  COND2X1 U2797 ( .A(n2962), .B(n2569), .C(n2449), .D(n2963), .Z(n1262) );
  CENX1 U2798 ( .A(n2467), .B(n2501), .Z(n2962) );
  COND2X1 U2799 ( .A(n2963), .B(n2569), .C(n2449), .D(n2964), .Z(n1261) );
  CENX1 U2800 ( .A(n2467), .B(n2500), .Z(n2963) );
  COND2X1 U2801 ( .A(n2964), .B(n2569), .C(n2449), .D(n2965), .Z(n1260) );
  CENX1 U2802 ( .A(n2467), .B(n2499), .Z(n2964) );
  COND2X1 U2803 ( .A(n2965), .B(n2569), .C(n2449), .D(n2966), .Z(n1259) );
  CENX1 U2804 ( .A(n2467), .B(n2498), .Z(n2965) );
  COND2X1 U2805 ( .A(n2966), .B(n2569), .C(n2449), .D(n2967), .Z(n1258) );
  CENX1 U2806 ( .A(n2467), .B(n2497), .Z(n2966) );
  COND2X1 U2807 ( .A(n2967), .B(n2569), .C(n2449), .D(n2968), .Z(n1257) );
  CENX1 U2808 ( .A(n2467), .B(n2496), .Z(n2967) );
  COND2X1 U2809 ( .A(n2968), .B(n2569), .C(n2449), .D(n2969), .Z(n1256) );
  CENX1 U2810 ( .A(n2467), .B(n2495), .Z(n2968) );
  COND2X1 U2811 ( .A(n2969), .B(n2569), .C(n2449), .D(n2970), .Z(n1255) );
  CENX1 U2812 ( .A(n2467), .B(n2494), .Z(n2969) );
  COND2X1 U2813 ( .A(n2970), .B(n2569), .C(n2449), .D(n2971), .Z(n1254) );
  CENX1 U2814 ( .A(n2467), .B(n2493), .Z(n2970) );
  COND2X1 U2815 ( .A(n2971), .B(n2569), .C(n2449), .D(n2568), .Z(n1253) );
  CEOX1 U2816 ( .A(n2467), .B(b[30]), .Z(n2568) );
  CENX1 U2817 ( .A(n2467), .B(n2492), .Z(n2971) );
  CAOR1X1 U2818 ( .A(n2569), .B(n2449), .C(n2571), .Z(n1252) );
  CEOX1 U2819 ( .A(n2467), .B(b[31]), .Z(n2571) );
  CNR2X1 U2820 ( .A(n2450), .B(n2515), .Z(n1251) );
  COND2X1 U2821 ( .A(n2972), .B(n2573), .C(n2450), .D(n2973), .Z(n1250) );
  CENX1 U2822 ( .A(n2515), .B(n2465), .Z(n2972) );
  COND2X1 U2823 ( .A(n2973), .B(n2573), .C(n2450), .D(n2974), .Z(n1249) );
  CENX1 U2824 ( .A(n2465), .B(n2453), .Z(n2973) );
  COND2X1 U2825 ( .A(n2974), .B(n2573), .C(n2450), .D(n2975), .Z(n1248) );
  CENX1 U2826 ( .A(n2465), .B(n2454), .Z(n2974) );
  COND2X1 U2827 ( .A(n2975), .B(n2573), .C(n2450), .D(n2976), .Z(n1247) );
  CENX1 U2828 ( .A(n2465), .B(n2455), .Z(n2975) );
  COND2X1 U2829 ( .A(n2976), .B(n2573), .C(n2450), .D(n2977), .Z(n1246) );
  CENX1 U2830 ( .A(n2465), .B(n2456), .Z(n2976) );
  COND2X1 U2831 ( .A(n2977), .B(n2573), .C(n2450), .D(n2978), .Z(n1245) );
  CENX1 U2832 ( .A(n2465), .B(n2457), .Z(n2977) );
  COND2X1 U2833 ( .A(n2978), .B(n2573), .C(n2450), .D(n2979), .Z(n1244) );
  CENX1 U2834 ( .A(n2465), .B(n2458), .Z(n2978) );
  COND2X1 U2835 ( .A(n2979), .B(n2573), .C(n2450), .D(n2980), .Z(n1243) );
  CENX1 U2836 ( .A(n2465), .B(n2514), .Z(n2979) );
  COND2X1 U2837 ( .A(n2980), .B(n2573), .C(n2450), .D(n2981), .Z(n1242) );
  CENX1 U2838 ( .A(n2465), .B(n2513), .Z(n2980) );
  COND2X1 U2839 ( .A(n2981), .B(n2573), .C(n2450), .D(n2982), .Z(n1241) );
  CENX1 U2840 ( .A(n2465), .B(n2512), .Z(n2981) );
  COND2X1 U2841 ( .A(n2982), .B(n2573), .C(n2450), .D(n2983), .Z(n1240) );
  CENX1 U2842 ( .A(n2465), .B(n2511), .Z(n2982) );
  COND2X1 U2843 ( .A(n2983), .B(n2573), .C(n2450), .D(n2984), .Z(n1239) );
  CENX1 U2844 ( .A(n2465), .B(n2510), .Z(n2983) );
  COND2X1 U2845 ( .A(n2984), .B(n2573), .C(n2450), .D(n2985), .Z(n1238) );
  CENX1 U2846 ( .A(n2465), .B(n2509), .Z(n2984) );
  COND2X1 U2847 ( .A(n2985), .B(n2573), .C(n2450), .D(n2986), .Z(n1237) );
  CENX1 U2848 ( .A(n2465), .B(n2508), .Z(n2985) );
  COND2X1 U2849 ( .A(n2986), .B(n2573), .C(n2450), .D(n2987), .Z(n1236) );
  CENX1 U2850 ( .A(n2465), .B(n2507), .Z(n2986) );
  COND2X1 U2851 ( .A(n2987), .B(n2573), .C(n2450), .D(n2988), .Z(n1235) );
  CENX1 U2852 ( .A(n2465), .B(n2506), .Z(n2987) );
  COND2X1 U2853 ( .A(n2988), .B(n2573), .C(n2450), .D(n2989), .Z(n1234) );
  CENX1 U2854 ( .A(n2465), .B(n2505), .Z(n2988) );
  COND2X1 U2855 ( .A(n2989), .B(n2573), .C(n2450), .D(n2990), .Z(n1233) );
  CENX1 U2856 ( .A(n2465), .B(n2504), .Z(n2989) );
  COND2X1 U2857 ( .A(n2990), .B(n2573), .C(n2450), .D(n2991), .Z(n1232) );
  CENX1 U2858 ( .A(n2465), .B(n2503), .Z(n2990) );
  COND2X1 U2859 ( .A(n2991), .B(n2573), .C(n2450), .D(n2992), .Z(n1231) );
  CENX1 U2860 ( .A(n2465), .B(n2502), .Z(n2991) );
  COND2X1 U2861 ( .A(n2992), .B(n2573), .C(n2450), .D(n2993), .Z(n1230) );
  CENX1 U2862 ( .A(n2465), .B(n2501), .Z(n2992) );
  COND2X1 U2863 ( .A(n2993), .B(n2573), .C(n2450), .D(n2994), .Z(n1229) );
  CENX1 U2864 ( .A(n2465), .B(n2500), .Z(n2993) );
  COND2X1 U2865 ( .A(n2994), .B(n2573), .C(n2450), .D(n2995), .Z(n1228) );
  CENX1 U2866 ( .A(n2465), .B(n2499), .Z(n2994) );
  COND2X1 U2867 ( .A(n2995), .B(n2573), .C(n2450), .D(n2996), .Z(n1227) );
  CENX1 U2868 ( .A(n2465), .B(n2498), .Z(n2995) );
  COND2X1 U2869 ( .A(n2996), .B(n2573), .C(n2450), .D(n2997), .Z(n1226) );
  CENX1 U2870 ( .A(n2465), .B(n2497), .Z(n2996) );
  COND2X1 U2871 ( .A(n2997), .B(n2573), .C(n2450), .D(n2998), .Z(n1225) );
  CENX1 U2872 ( .A(n2465), .B(n2496), .Z(n2997) );
  COND2X1 U2873 ( .A(n2998), .B(n2573), .C(n2450), .D(n2999), .Z(n1224) );
  CENX1 U2874 ( .A(n2465), .B(n2495), .Z(n2998) );
  COND2X1 U2875 ( .A(n2999), .B(n2573), .C(n2450), .D(n3000), .Z(n1223) );
  CENX1 U2876 ( .A(n2465), .B(n2494), .Z(n2999) );
  COND2X1 U2877 ( .A(n3000), .B(n2573), .C(n2450), .D(n3001), .Z(n1222) );
  CENX1 U2878 ( .A(n2465), .B(n2493), .Z(n3000) );
  COND2X1 U2879 ( .A(n3001), .B(n2573), .C(n2450), .D(n2572), .Z(n1221) );
  CEOX1 U2880 ( .A(n2465), .B(b[30]), .Z(n2572) );
  CENX1 U2881 ( .A(n2465), .B(n2492), .Z(n3001) );
  CAOR1X1 U2882 ( .A(n2573), .B(n2450), .C(n2575), .Z(n1220) );
  CEOX1 U2883 ( .A(n2465), .B(b[31]), .Z(n2575) );
  CNR2X1 U2884 ( .A(n2451), .B(n2515), .Z(n1219) );
  COND2X1 U2885 ( .A(n3002), .B(n2519), .C(n2451), .D(n3003), .Z(n1218) );
  CENX1 U2886 ( .A(n2515), .B(n2463), .Z(n3002) );
  COND2X1 U2887 ( .A(n3003), .B(n2519), .C(n2451), .D(n3004), .Z(n1217) );
  CENX1 U2888 ( .A(n2463), .B(n2453), .Z(n3003) );
  COND2X1 U2889 ( .A(n3004), .B(n2519), .C(n2451), .D(n2518), .Z(n1216) );
  CENX1 U2890 ( .A(n2463), .B(n2455), .Z(n2518) );
  CENX1 U2891 ( .A(n2463), .B(n2454), .Z(n3004) );
  COND2X1 U2892 ( .A(n2521), .B(n2519), .C(n2451), .D(n3005), .Z(n1214) );
  CENX1 U2893 ( .A(n2463), .B(n2456), .Z(n2521) );
  COND2X1 U2894 ( .A(n3005), .B(n2519), .C(n2451), .D(n3006), .Z(n1213) );
  CENX1 U2895 ( .A(n2463), .B(n2457), .Z(n3005) );
  COND2X1 U2896 ( .A(n3006), .B(n2519), .C(n2451), .D(n3007), .Z(n1212) );
  CENX1 U2897 ( .A(n2463), .B(n2458), .Z(n3006) );
  COND2X1 U2898 ( .A(n3007), .B(n2519), .C(n2451), .D(n3008), .Z(n1211) );
  CENX1 U2899 ( .A(n2463), .B(n2514), .Z(n3007) );
  COND2X1 U2900 ( .A(n3008), .B(n2519), .C(n2451), .D(n3009), .Z(n1210) );
  CENX1 U2901 ( .A(n2463), .B(n2513), .Z(n3008) );
  COND2X1 U2902 ( .A(n3009), .B(n2519), .C(n2451), .D(n3010), .Z(n1209) );
  CENX1 U2903 ( .A(n2463), .B(n2512), .Z(n3009) );
  COND2X1 U2904 ( .A(n3010), .B(n2519), .C(n2451), .D(n3011), .Z(n1208) );
  CENX1 U2905 ( .A(n2463), .B(n2511), .Z(n3010) );
  COND2X1 U2906 ( .A(n3011), .B(n2519), .C(n2451), .D(n3012), .Z(n1207) );
  CENX1 U2907 ( .A(n2463), .B(n2510), .Z(n3011) );
  COND2X1 U2908 ( .A(n3012), .B(n2519), .C(n2451), .D(n3013), .Z(n1206) );
  CENX1 U2909 ( .A(n2463), .B(n2509), .Z(n3012) );
  COND2X1 U2910 ( .A(n3013), .B(n2519), .C(n2451), .D(n3014), .Z(n1205) );
  CENX1 U2911 ( .A(n2463), .B(n2508), .Z(n3013) );
  COND2X1 U2912 ( .A(n3014), .B(n2519), .C(n2451), .D(n3015), .Z(n1204) );
  CENX1 U2913 ( .A(n2463), .B(n2507), .Z(n3014) );
  COND2X1 U2914 ( .A(n3015), .B(n2519), .C(n2451), .D(n3016), .Z(n1203) );
  CENX1 U2915 ( .A(n2463), .B(n2506), .Z(n3015) );
  COND2X1 U2916 ( .A(n3016), .B(n2519), .C(n2451), .D(n3017), .Z(n1202) );
  CENX1 U2917 ( .A(n2463), .B(n2505), .Z(n3016) );
  COND2X1 U2918 ( .A(n3017), .B(n2519), .C(n2451), .D(n3018), .Z(n1201) );
  CENX1 U2919 ( .A(n2463), .B(n2504), .Z(n3017) );
  COND2X1 U2920 ( .A(n3018), .B(n2519), .C(n2451), .D(n3019), .Z(n1200) );
  CENX1 U2921 ( .A(n2463), .B(n2503), .Z(n3018) );
  COND2X1 U2922 ( .A(n3019), .B(n2519), .C(n2451), .D(n3020), .Z(n1199) );
  CENX1 U2923 ( .A(n2463), .B(n2502), .Z(n3019) );
  COND2X1 U2924 ( .A(n3020), .B(n2519), .C(n2451), .D(n3021), .Z(n1198) );
  CENX1 U2925 ( .A(n2463), .B(n2501), .Z(n3020) );
  COND2X1 U2926 ( .A(n3021), .B(n2519), .C(n2451), .D(n3022), .Z(n1197) );
  CENX1 U2927 ( .A(n2463), .B(n2500), .Z(n3021) );
  COND2X1 U2928 ( .A(n3022), .B(n2519), .C(n2451), .D(n3023), .Z(n1196) );
  CENX1 U2929 ( .A(n2463), .B(n2499), .Z(n3022) );
  COND2X1 U2930 ( .A(n3023), .B(n2519), .C(n2451), .D(n3024), .Z(n1195) );
  CENX1 U2931 ( .A(n2463), .B(n2498), .Z(n3023) );
  COND2X1 U2932 ( .A(n3024), .B(n2519), .C(n2451), .D(n3025), .Z(n1194) );
  CENX1 U2933 ( .A(n2463), .B(n2497), .Z(n3024) );
  COND2X1 U2934 ( .A(n3025), .B(n2519), .C(n2451), .D(n3026), .Z(n1193) );
  CENX1 U2935 ( .A(n2463), .B(n2496), .Z(n3025) );
  COND2X1 U2936 ( .A(n3026), .B(n2519), .C(n2451), .D(n3027), .Z(n1192) );
  CENX1 U2937 ( .A(n2463), .B(n2495), .Z(n3026) );
  COND2X1 U2938 ( .A(n3027), .B(n2519), .C(n2451), .D(n3028), .Z(n1191) );
  CENX1 U2939 ( .A(n2463), .B(n2494), .Z(n3027) );
  COND2X1 U2940 ( .A(n3028), .B(n2519), .C(n2451), .D(n3029), .Z(n1190) );
  CENX1 U2941 ( .A(n2463), .B(n2493), .Z(n3028) );
  COND2X1 U2942 ( .A(n3029), .B(n2519), .C(n2451), .D(n2576), .Z(n1189) );
  CEOX1 U2943 ( .A(n2463), .B(b[30]), .Z(n2576) );
  CENX1 U2944 ( .A(n2463), .B(n2492), .Z(n3029) );
  CAOR1X1 U2945 ( .A(n2519), .B(n2451), .C(n2577), .Z(n1188) );
  CEOX1 U2946 ( .A(n2463), .B(b[31]), .Z(n2577) );
  CNR2X1 U2947 ( .A(n2452), .B(n2515), .Z(n1187) );
  COND2X1 U2948 ( .A(n3030), .B(n2579), .C(n2452), .D(n3031), .Z(n1186) );
  CENX1 U2949 ( .A(n2515), .B(n2461), .Z(n3030) );
  COND2X1 U2950 ( .A(n3031), .B(n2579), .C(n2452), .D(n3032), .Z(n1185) );
  CENX1 U2951 ( .A(n2461), .B(n2453), .Z(n3031) );
  COND2X1 U2952 ( .A(n3032), .B(n2579), .C(n2452), .D(n3033), .Z(n1184) );
  CENX1 U2953 ( .A(n2461), .B(n2454), .Z(n3032) );
  COND2X1 U2954 ( .A(n3033), .B(n2579), .C(n2452), .D(n3034), .Z(n1183) );
  CENX1 U2955 ( .A(n2461), .B(n2455), .Z(n3033) );
  COND2X1 U2956 ( .A(n3034), .B(n2579), .C(n2452), .D(n3035), .Z(n1182) );
  CENX1 U2957 ( .A(n2461), .B(n2456), .Z(n3034) );
  COND2X1 U2958 ( .A(n3035), .B(n2579), .C(n2452), .D(n3036), .Z(n1181) );
  CENX1 U2959 ( .A(n2461), .B(n2457), .Z(n3035) );
  COND2X1 U2960 ( .A(n3036), .B(n2579), .C(n2452), .D(n3037), .Z(n1180) );
  CENX1 U2961 ( .A(n2461), .B(n2458), .Z(n3036) );
  COND2X1 U2962 ( .A(n3037), .B(n2579), .C(n2452), .D(n3038), .Z(n1179) );
  CENX1 U2963 ( .A(n2461), .B(n2514), .Z(n3037) );
  COND2X1 U2964 ( .A(n3038), .B(n2579), .C(n2452), .D(n3039), .Z(n1178) );
  CENX1 U2965 ( .A(n2461), .B(n2513), .Z(n3038) );
  COND2X1 U2966 ( .A(n3039), .B(n2579), .C(n2452), .D(n3040), .Z(n1177) );
  CENX1 U2967 ( .A(n2461), .B(n2512), .Z(n3039) );
  COND2X1 U2968 ( .A(n3040), .B(n2579), .C(n2452), .D(n3041), .Z(n1176) );
  CENX1 U2969 ( .A(n2461), .B(n2511), .Z(n3040) );
  COND2X1 U2970 ( .A(n3041), .B(n2579), .C(n2452), .D(n3042), .Z(n1175) );
  CENX1 U2971 ( .A(n2461), .B(n2510), .Z(n3041) );
  COND2X1 U2972 ( .A(n3042), .B(n2579), .C(n2452), .D(n3043), .Z(n1174) );
  CENX1 U2973 ( .A(n2461), .B(n2509), .Z(n3042) );
  COND2X1 U2974 ( .A(n3043), .B(n2579), .C(n2452), .D(n3044), .Z(n1173) );
  CENX1 U2975 ( .A(n2461), .B(n2508), .Z(n3043) );
  COND2X1 U2976 ( .A(n3044), .B(n2579), .C(n2452), .D(n3045), .Z(n1172) );
  CENX1 U2977 ( .A(n2461), .B(n2507), .Z(n3044) );
  COND2X1 U2978 ( .A(n3045), .B(n2579), .C(n2452), .D(n3046), .Z(n1171) );
  CENX1 U2979 ( .A(n2461), .B(n2506), .Z(n3045) );
  COND2X1 U2980 ( .A(n3046), .B(n2579), .C(n2452), .D(n3047), .Z(n1170) );
  CENX1 U2981 ( .A(n2461), .B(n2505), .Z(n3046) );
  COND2X1 U2982 ( .A(n3047), .B(n2579), .C(n2452), .D(n3048), .Z(n1169) );
  CENX1 U2983 ( .A(n2461), .B(n2504), .Z(n3047) );
  COND2X1 U2984 ( .A(n3048), .B(n2579), .C(n2452), .D(n3049), .Z(n1168) );
  CENX1 U2985 ( .A(n2461), .B(n2503), .Z(n3048) );
  COND2X1 U2986 ( .A(n3049), .B(n2579), .C(n2452), .D(n3050), .Z(n1167) );
  CENX1 U2987 ( .A(n2461), .B(n2502), .Z(n3049) );
  COND2X1 U2988 ( .A(n3050), .B(n2579), .C(n2452), .D(n3051), .Z(n1166) );
  CENX1 U2989 ( .A(n2461), .B(n2501), .Z(n3050) );
  COND2X1 U2990 ( .A(n3051), .B(n2579), .C(n2452), .D(n3052), .Z(n1165) );
  CENX1 U2991 ( .A(n2461), .B(n2500), .Z(n3051) );
  COND2X1 U2992 ( .A(n3052), .B(n2579), .C(n2452), .D(n3053), .Z(n1164) );
  CENX1 U2993 ( .A(n2461), .B(n2499), .Z(n3052) );
  COND2X1 U2994 ( .A(n3053), .B(n2579), .C(n2452), .D(n3054), .Z(n1163) );
  CENX1 U2995 ( .A(n2461), .B(n2498), .Z(n3053) );
  COND2X1 U2996 ( .A(n3054), .B(n2579), .C(n2452), .D(n3055), .Z(n1162) );
  CENX1 U2997 ( .A(n2461), .B(n2497), .Z(n3054) );
  COND2X1 U2998 ( .A(n3055), .B(n2579), .C(n2452), .D(n3056), .Z(n1161) );
  CENX1 U2999 ( .A(n2461), .B(n2496), .Z(n3055) );
  COND2X1 U3000 ( .A(n3056), .B(n2579), .C(n2452), .D(n3057), .Z(n1160) );
  CENX1 U3001 ( .A(n2461), .B(n2495), .Z(n3056) );
  COND2X1 U3002 ( .A(n3057), .B(n2579), .C(n2452), .D(n3058), .Z(n1159) );
  CENX1 U3003 ( .A(n2461), .B(n2494), .Z(n3057) );
  COND2X1 U3004 ( .A(n3058), .B(n2579), .C(n2452), .D(n3059), .Z(n1158) );
  CENX1 U3005 ( .A(n2461), .B(n2493), .Z(n3058) );
  COND2X1 U3006 ( .A(n3059), .B(n2579), .C(n2452), .D(n2578), .Z(n1157) );
  CEOX1 U3007 ( .A(n2461), .B(b[30]), .Z(n2578) );
  CENX1 U3008 ( .A(n2461), .B(n2492), .Z(n3059) );
  CAOR1X1 U3009 ( .A(n2579), .B(n2452), .C(n2581), .Z(n1156) );
  CEOX1 U3010 ( .A(n2461), .B(b[31]), .Z(n2581) );
  COND1XL U3011 ( .A(b[0]), .B(n2490), .C(n2582), .Z(n1155) );
  COND11X1 U3012 ( .A(n2489), .B(b[0]), .C(n2438), .D(n3060), .Z(n1154) );
  CND2IX1 U3013 ( .B(n2527), .A(a[3]), .Z(n3060) );
  CENX1 U3014 ( .A(n2489), .B(a[2]), .Z(n3061) );
  COND11X1 U3015 ( .A(n2487), .B(b[0]), .C(n2439), .D(n3062), .Z(n1153) );
  CND2IX1 U3016 ( .B(n2531), .A(a[5]), .Z(n3062) );
  CENX1 U3017 ( .A(n2487), .B(a[4]), .Z(n3063) );
  COND11X1 U3018 ( .A(n2485), .B(b[0]), .C(n2440), .D(n3064), .Z(n1152) );
  CND2IX1 U3019 ( .B(n2535), .A(a[7]), .Z(n3064) );
  CENX1 U3020 ( .A(n2485), .B(a[6]), .Z(n3065) );
  COND11X1 U3021 ( .A(n2483), .B(b[0]), .C(n2441), .D(n3066), .Z(n1151) );
  CND2IX1 U3022 ( .B(n2539), .A(a[9]), .Z(n3066) );
  CENX1 U3023 ( .A(n2483), .B(a[8]), .Z(n3067) );
  COND11X1 U3024 ( .A(n2481), .B(b[0]), .C(n2442), .D(n3068), .Z(n1150) );
  CND2IX1 U3025 ( .B(n2543), .A(a[11]), .Z(n3068) );
  CENX1 U3026 ( .A(n2481), .B(a[10]), .Z(n3069) );
  COND11X1 U3027 ( .A(n2479), .B(b[0]), .C(n2443), .D(n3070), .Z(n1149) );
  CND2IX1 U3028 ( .B(n2523), .A(a[13]), .Z(n3070) );
  CENX1 U3029 ( .A(n2479), .B(a[12]), .Z(n3071) );
  COND11X1 U3030 ( .A(n2477), .B(b[0]), .C(n2444), .D(n3072), .Z(n1148) );
  CND2IX1 U3031 ( .B(n2549), .A(a[15]), .Z(n3072) );
  CENX1 U3032 ( .A(n2477), .B(a[14]), .Z(n3073) );
  COND11X1 U3033 ( .A(n2475), .B(b[0]), .C(n2445), .D(n3074), .Z(n1147) );
  CND2IX1 U3034 ( .B(n2553), .A(a[17]), .Z(n3074) );
  CENX1 U3035 ( .A(n2475), .B(a[16]), .Z(n3075) );
  COND11X1 U3036 ( .A(n2473), .B(b[0]), .C(n2446), .D(n3076), .Z(n1146) );
  CND2IX1 U3037 ( .B(n2557), .A(a[19]), .Z(n3076) );
  CENX1 U3038 ( .A(n2473), .B(a[18]), .Z(n3077) );
  COND11X1 U3039 ( .A(n2471), .B(b[0]), .C(n2447), .D(n3078), .Z(n1145) );
  CND2IX1 U3040 ( .B(n2561), .A(a[21]), .Z(n3078) );
  CENX1 U3041 ( .A(n2471), .B(a[20]), .Z(n3079) );
  COND11X1 U3042 ( .A(n2469), .B(b[0]), .C(n2448), .D(n3080), .Z(n1144) );
  CND2IX1 U3043 ( .B(n2565), .A(a[23]), .Z(n3080) );
  CENX1 U3044 ( .A(n2469), .B(a[22]), .Z(n3081) );
  COND11X1 U3045 ( .A(n2467), .B(b[0]), .C(n2449), .D(n3082), .Z(n1143) );
  CND2IX1 U3046 ( .B(n2569), .A(a[25]), .Z(n3082) );
  CENX1 U3047 ( .A(n2467), .B(a[24]), .Z(n3083) );
  COND11X1 U3048 ( .A(n2465), .B(b[0]), .C(n2450), .D(n3084), .Z(n1142) );
  CND2IX1 U3049 ( .B(n2573), .A(a[27]), .Z(n3084) );
  CENX1 U3050 ( .A(n2465), .B(a[26]), .Z(n3085) );
  COND11X1 U3051 ( .A(n2463), .B(b[0]), .C(n2451), .D(n3086), .Z(n1141) );
  CND2IX1 U3052 ( .B(n2519), .A(a[29]), .Z(n3086) );
  CENX1 U3053 ( .A(n2463), .B(a[28]), .Z(n3087) );
  COND11X1 U3054 ( .A(n2461), .B(b[0]), .C(n2452), .D(n3088), .Z(n1140) );
  CND2IX1 U3055 ( .B(n2579), .A(a[31]), .Z(n3088) );
  CENX1 U3056 ( .A(n2461), .B(a[30]), .Z(n3089) );
endmodule


module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push0, _pushout_d, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39,
         N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53,
         N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67,
         N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, n8, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] acc;
  wire   [1:0] cmd0;

  CAOR2X1 U3 ( .A(q[2]), .B(n420), .C(q0[2]), .D(n433), .Z(n245) );
  CAOR2X1 U4 ( .A(q[3]), .B(n420), .C(q0[3]), .D(n446), .Z(n246) );
  CAOR2X1 U8 ( .A(q[4]), .B(n420), .C(q0[4]), .D(n431), .Z(n247) );
  CAOR2X1 U9 ( .A(q[5]), .B(n420), .C(q0[5]), .D(n432), .Z(n248) );
  CAOR2X1 U10 ( .A(q[6]), .B(n419), .C(q0[6]), .D(n429), .Z(n249) );
  CAOR2X1 U11 ( .A(q[7]), .B(n419), .C(q0[7]), .D(n430), .Z(n250) );
  CAOR2X1 U12 ( .A(q[8]), .B(n419), .C(q0[8]), .D(n427), .Z(n251) );
  CAOR2X1 U13 ( .A(q[9]), .B(n419), .C(q0[9]), .D(n428), .Z(n252) );
  CAOR2X1 U14 ( .A(q[10]), .B(n419), .C(q0[10]), .D(n425), .Z(n253) );
  CAOR2X1 U15 ( .A(q[11]), .B(n419), .C(q0[11]), .D(n426), .Z(n254) );
  CAOR2X1 U16 ( .A(q[12]), .B(n419), .C(q0[12]), .D(n421), .Z(n255) );
  CAOR2X1 U17 ( .A(q[13]), .B(n419), .C(q0[13]), .D(n421), .Z(n256) );
  CAOR2X1 U18 ( .A(q[14]), .B(n419), .C(q0[14]), .D(n422), .Z(n257) );
  CAOR2X1 U19 ( .A(q[15]), .B(n419), .C(q0[15]), .D(n422), .Z(n258) );
  CAOR2X1 U20 ( .A(q[16]), .B(n419), .C(q0[16]), .D(n423), .Z(n259) );
  CAOR2X1 U21 ( .A(q[17]), .B(n419), .C(q0[17]), .D(n423), .Z(n260) );
  CAOR2X1 U22 ( .A(q[18]), .B(n418), .C(q0[18]), .D(n424), .Z(n261) );
  CAOR2X1 U23 ( .A(q[19]), .B(n418), .C(q0[19]), .D(n424), .Z(n262) );
  CAOR2X1 U24 ( .A(q[20]), .B(n418), .C(q0[20]), .D(n425), .Z(n263) );
  CAOR2X1 U25 ( .A(q[21]), .B(n418), .C(q0[21]), .D(n425), .Z(n264) );
  CAOR2X1 U26 ( .A(q[22]), .B(n418), .C(q0[22]), .D(n426), .Z(n265) );
  CAOR2X1 U27 ( .A(q[23]), .B(n418), .C(q0[23]), .D(n426), .Z(n266) );
  CAOR2X1 U28 ( .A(q[24]), .B(n418), .C(q0[24]), .D(n427), .Z(n267) );
  CAOR2X1 U29 ( .A(q[25]), .B(n418), .C(q0[25]), .D(n427), .Z(n268) );
  CAOR2X1 U30 ( .A(q[26]), .B(n418), .C(q0[26]), .D(n428), .Z(n269) );
  CAOR2X1 U31 ( .A(q[27]), .B(n418), .C(q0[27]), .D(n428), .Z(n270) );
  CAOR2X1 U32 ( .A(q[28]), .B(n418), .C(q0[28]), .D(n429), .Z(n271) );
  CAOR2X1 U33 ( .A(q[29]), .B(n418), .C(q0[29]), .D(n429), .Z(n272) );
  CAOR2X1 U34 ( .A(q[30]), .B(n417), .C(q0[30]), .D(n430), .Z(n273) );
  CAOR2X1 U35 ( .A(q[31]), .B(n417), .C(q0[31]), .D(n430), .Z(n274) );
  CAOR2X1 U269 ( .A(h[0]), .B(n417), .C(h0[0]), .D(n431), .Z(n211) );
  CAOR2X1 U270 ( .A(h[1]), .B(n417), .C(n399), .D(n431), .Z(n212) );
  CAOR2X1 U271 ( .A(h[2]), .B(n417), .C(n351), .D(n432), .Z(n213) );
  CAOR2X1 U272 ( .A(h[3]), .B(n417), .C(n405), .D(n432), .Z(n214) );
  CAOR2X1 U273 ( .A(h[4]), .B(n417), .C(n356), .D(n433), .Z(n215) );
  CAOR2X1 U274 ( .A(h[5]), .B(n417), .C(n410), .D(n433), .Z(n216) );
  CAOR2X1 U275 ( .A(h[6]), .B(n417), .C(n414), .D(n434), .Z(n217) );
  CAOR2X1 U299 ( .A(h[30]), .B(n415), .C(h0[30]), .D(n446), .Z(n241) );
  CAOR2X1 U300 ( .A(h[31]), .B(n415), .C(h0[31]), .D(n446), .Z(n242) );
  CAOR2X1 U302 ( .A(q[1]), .B(n415), .C(q0[1]), .D(n447), .Z(n244) );
  sfilt_DW01_add_0 add_43 ( .A({N272, N271, N270, N269, N268, N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, 
        N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, 
        N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, 
        N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, 
        N216, N215, N214, N213, N212, N211, N210, N209}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        N208}), .CI(1'b0), .SUM({N336, N335, N334, N333, N332, N331, N330, 
        N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, 
        N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, 
        N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, 
        N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280, N279, N278, N277, N276, N275, N274, N273}) );
  sfilt_DW01_add_1 add_39 ( .A({N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16}), .B(
        acc), .CI(1'b0), .SUM({N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, 
        N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, 
        N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, 
        N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, 
        N151, N150, N149, N148, N147, N146, N145, N144}) );
  sfilt_DW_mult_tc_0 r300 ( .a(q0), .b({h0[31:7], n414, n410, n356, n405, n353, 
        n399, h0[0]}), .product({N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16}) );
  CFD2QXL \dout_reg[31]  ( .D(n307), .CP(clk), .CD(n372), .Q(z[31]) );
  CFD2QXL \dout_reg[30]  ( .D(n306), .CP(clk), .CD(n372), .Q(z[30]) );
  CFD2QXL \dout_reg[29]  ( .D(n305), .CP(clk), .CD(n372), .Q(z[29]) );
  CFD2QXL \dout_reg[28]  ( .D(n304), .CP(clk), .CD(n372), .Q(z[28]) );
  CFD2QXL \dout_reg[27]  ( .D(n303), .CP(clk), .CD(n372), .Q(z[27]) );
  CFD2QXL \dout_reg[26]  ( .D(n302), .CP(clk), .CD(n372), .Q(z[26]) );
  CFD2QXL \dout_reg[25]  ( .D(n301), .CP(clk), .CD(n372), .Q(z[25]) );
  CFD2QXL \dout_reg[24]  ( .D(n300), .CP(clk), .CD(n372), .Q(z[24]) );
  CFD2QXL \dout_reg[23]  ( .D(n299), .CP(clk), .CD(n372), .Q(z[23]) );
  CFD2QXL \dout_reg[22]  ( .D(n298), .CP(clk), .CD(n372), .Q(z[22]) );
  CFD2QXL \dout_reg[21]  ( .D(n297), .CP(clk), .CD(n372), .Q(z[21]) );
  CFD2QXL \dout_reg[20]  ( .D(n296), .CP(clk), .CD(n373), .Q(z[20]) );
  CFD2QXL \dout_reg[19]  ( .D(n295), .CP(clk), .CD(n373), .Q(z[19]) );
  CFD2QXL \dout_reg[18]  ( .D(n294), .CP(clk), .CD(n373), .Q(z[18]) );
  CFD2QXL \dout_reg[17]  ( .D(n293), .CP(clk), .CD(n373), .Q(z[17]) );
  CFD2QXL \dout_reg[16]  ( .D(n292), .CP(clk), .CD(n373), .Q(z[16]) );
  CFD2QXL \dout_reg[15]  ( .D(n291), .CP(clk), .CD(n373), .Q(z[15]) );
  CFD2QXL \dout_reg[14]  ( .D(n290), .CP(clk), .CD(n373), .Q(z[14]) );
  CFD2QXL \dout_reg[13]  ( .D(n289), .CP(clk), .CD(n373), .Q(z[13]) );
  CFD2QXL \dout_reg[12]  ( .D(n288), .CP(clk), .CD(n373), .Q(z[12]) );
  CFD2QXL \dout_reg[11]  ( .D(n287), .CP(clk), .CD(n373), .Q(z[11]) );
  CFD2QXL \dout_reg[10]  ( .D(n286), .CP(clk), .CD(n373), .Q(z[10]) );
  CFD2QXL \dout_reg[9]  ( .D(n285), .CP(clk), .CD(n373), .Q(z[9]) );
  CFD2QXL \dout_reg[8]  ( .D(n284), .CP(clk), .CD(n373), .Q(z[8]) );
  CFD2QXL \dout_reg[7]  ( .D(n283), .CP(clk), .CD(n374), .Q(z[7]) );
  CFD2QXL \dout_reg[6]  ( .D(n282), .CP(clk), .CD(n374), .Q(z[6]) );
  CFD2QXL \dout_reg[5]  ( .D(n281), .CP(clk), .CD(n374), .Q(z[5]) );
  CFD2QXL \dout_reg[4]  ( .D(n280), .CP(clk), .CD(n374), .Q(z[4]) );
  CFD2QXL \dout_reg[3]  ( .D(n279), .CP(clk), .CD(n374), .Q(z[3]) );
  CFD2QXL \dout_reg[2]  ( .D(n278), .CP(clk), .CD(n374), .Q(z[2]) );
  CFD2QXL \dout_reg[1]  ( .D(n277), .CP(clk), .CD(n374), .Q(z[1]) );
  CFD2QXL \dout_reg[0]  ( .D(n276), .CP(clk), .CD(n374), .Q(z[0]) );
  CFD2QXL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n362), .Q(cmd0[0]) );
  CFD2QXL push0_reg ( .D(n420), .CP(clk), .CD(n362), .Q(push0) );
  CFD2QXL \acc_reg[32]  ( .D(n177), .CP(clk), .CD(n369), .Q(acc[32]) );
  CFD2QXL \acc_reg[33]  ( .D(n176), .CP(clk), .CD(n369), .Q(acc[33]) );
  CFD2QXL \acc_reg[34]  ( .D(n175), .CP(clk), .CD(n369), .Q(acc[34]) );
  CFD2QXL \acc_reg[35]  ( .D(n174), .CP(clk), .CD(n370), .Q(acc[35]) );
  CFD2QXL \acc_reg[36]  ( .D(n173), .CP(clk), .CD(n370), .Q(acc[36]) );
  CFD2QXL \acc_reg[37]  ( .D(n172), .CP(clk), .CD(n370), .Q(acc[37]) );
  CFD2QXL \acc_reg[38]  ( .D(n171), .CP(clk), .CD(n370), .Q(acc[38]) );
  CFD2QXL \acc_reg[39]  ( .D(n170), .CP(clk), .CD(n370), .Q(acc[39]) );
  CFD2QXL \acc_reg[40]  ( .D(n169), .CP(clk), .CD(n370), .Q(acc[40]) );
  CFD2QXL \acc_reg[41]  ( .D(n168), .CP(clk), .CD(n370), .Q(acc[41]) );
  CFD2QXL \acc_reg[42]  ( .D(n167), .CP(clk), .CD(n370), .Q(acc[42]) );
  CFD2QXL \acc_reg[43]  ( .D(n166), .CP(clk), .CD(n370), .Q(acc[43]) );
  CFD2QXL \acc_reg[44]  ( .D(n165), .CP(clk), .CD(n370), .Q(acc[44]) );
  CFD2QXL \acc_reg[45]  ( .D(n164), .CP(clk), .CD(n370), .Q(acc[45]) );
  CFD2QXL \acc_reg[46]  ( .D(n163), .CP(clk), .CD(n370), .Q(acc[46]) );
  CFD2QXL \acc_reg[47]  ( .D(n162), .CP(clk), .CD(n370), .Q(acc[47]) );
  CFD2QXL \acc_reg[48]  ( .D(n161), .CP(clk), .CD(n371), .Q(acc[48]) );
  CFD2QXL \acc_reg[49]  ( .D(n160), .CP(clk), .CD(n371), .Q(acc[49]) );
  CFD2QXL \acc_reg[50]  ( .D(n159), .CP(clk), .CD(n371), .Q(acc[50]) );
  CFD2QXL \acc_reg[51]  ( .D(n158), .CP(clk), .CD(n371), .Q(acc[51]) );
  CFD2QXL \acc_reg[52]  ( .D(n157), .CP(clk), .CD(n371), .Q(acc[52]) );
  CFD2QXL \acc_reg[53]  ( .D(n156), .CP(clk), .CD(n371), .Q(acc[53]) );
  CFD2QXL \acc_reg[54]  ( .D(n155), .CP(clk), .CD(n371), .Q(acc[54]) );
  CFD2QXL \acc_reg[55]  ( .D(n154), .CP(clk), .CD(n371), .Q(acc[55]) );
  CFD2QXL \acc_reg[56]  ( .D(n153), .CP(clk), .CD(n371), .Q(acc[56]) );
  CFD2QXL \acc_reg[57]  ( .D(n152), .CP(clk), .CD(n371), .Q(acc[57]) );
  CFD2QXL \acc_reg[58]  ( .D(n151), .CP(clk), .CD(n371), .Q(acc[58]) );
  CFD2QXL \acc_reg[59]  ( .D(n150), .CP(clk), .CD(n371), .Q(acc[59]) );
  CFD2QXL \acc_reg[60]  ( .D(n149), .CP(clk), .CD(n371), .Q(acc[60]) );
  CFD2QXL \acc_reg[61]  ( .D(n148), .CP(clk), .CD(n372), .Q(acc[61]) );
  CFD2QXL \acc_reg[62]  ( .D(n147), .CP(clk), .CD(n372), .Q(acc[62]) );
  CFD2QXL \acc_reg[63]  ( .D(n210), .CP(clk), .CD(n367), .Q(acc[63]) );
  CFD2QXL \acc_reg[28]  ( .D(n181), .CP(clk), .CD(n369), .Q(acc[28]) );
  CFD2QXL \acc_reg[29]  ( .D(n180), .CP(clk), .CD(n369), .Q(acc[29]) );
  CFD2QXL \acc_reg[30]  ( .D(n179), .CP(clk), .CD(n369), .Q(acc[30]) );
  CFD2QXL \acc_reg[31]  ( .D(n178), .CP(clk), .CD(n369), .Q(acc[31]) );
  CFD2QXL \acc_reg[25]  ( .D(n184), .CP(clk), .CD(n369), .Q(acc[25]) );
  CFD2QXL \acc_reg[26]  ( .D(n183), .CP(clk), .CD(n369), .Q(acc[26]) );
  CFD2QXL \acc_reg[27]  ( .D(n182), .CP(clk), .CD(n369), .Q(acc[27]) );
  CFD2QXL \acc_reg[21]  ( .D(n188), .CP(clk), .CD(n368), .Q(acc[21]) );
  CFD2QXL \acc_reg[22]  ( .D(n187), .CP(clk), .CD(n369), .Q(acc[22]) );
  CFD2QXL \acc_reg[23]  ( .D(n186), .CP(clk), .CD(n369), .Q(acc[23]) );
  CFD2QXL \acc_reg[24]  ( .D(n185), .CP(clk), .CD(n369), .Q(acc[24]) );
  CFD2QXL \h0_reg[31]  ( .D(n242), .CP(clk), .CD(n364), .Q(h0[31]) );
  CFD2QXL \q0_reg[30]  ( .D(n273), .CP(clk), .CD(n362), .Q(q0[30]) );
  CFD2QXL \q0_reg[28]  ( .D(n271), .CP(clk), .CD(n362), .Q(q0[28]) );
  CFD2QXL \acc_reg[18]  ( .D(n191), .CP(clk), .CD(n368), .Q(acc[18]) );
  CFD2QXL \acc_reg[19]  ( .D(n190), .CP(clk), .CD(n368), .Q(acc[19]) );
  CFD2QXL \acc_reg[20]  ( .D(n189), .CP(clk), .CD(n368), .Q(acc[20]) );
  CFD2QXL \h0_reg[29]  ( .D(n240), .CP(clk), .CD(n364), .Q(h0[29]) );
  CFD2QXL \h0_reg[28]  ( .D(n239), .CP(clk), .CD(n365), .Q(h0[28]) );
  CFD2QXL \h0_reg[27]  ( .D(n238), .CP(clk), .CD(n365), .Q(h0[27]) );
  CFD2QXL \h0_reg[26]  ( .D(n237), .CP(clk), .CD(n365), .Q(h0[26]) );
  CFD2QXL \q0_reg[31]  ( .D(n274), .CP(clk), .CD(n362), .Q(q0[31]) );
  CFD2QXL \q0_reg[29]  ( .D(n272), .CP(clk), .CD(n362), .Q(q0[29]) );
  CFD2QXL \h0_reg[30]  ( .D(n241), .CP(clk), .CD(n364), .Q(h0[30]) );
  CFD2QXL \q0_reg[26]  ( .D(n269), .CP(clk), .CD(n362), .Q(q0[26]) );
  CFD2QXL \q0_reg[24]  ( .D(n267), .CP(clk), .CD(n362), .Q(q0[24]) );
  CFD2QXL \acc_reg[14]  ( .D(n195), .CP(clk), .CD(n368), .Q(acc[14]) );
  CFD2QXL \acc_reg[15]  ( .D(n194), .CP(clk), .CD(n368), .Q(acc[15]) );
  CFD2QXL \acc_reg[16]  ( .D(n193), .CP(clk), .CD(n368), .Q(acc[16]) );
  CFD2QXL \acc_reg[17]  ( .D(n192), .CP(clk), .CD(n368), .Q(acc[17]) );
  CFD2QXL \h0_reg[25]  ( .D(n236), .CP(clk), .CD(n365), .Q(h0[25]) );
  CFD2QXL \h0_reg[24]  ( .D(n235), .CP(clk), .CD(n365), .Q(h0[24]) );
  CFD2QXL \h0_reg[23]  ( .D(n234), .CP(clk), .CD(n365), .Q(h0[23]) );
  CFD2QXL \q0_reg[27]  ( .D(n270), .CP(clk), .CD(n362), .Q(q0[27]) );
  CFD2QXL \q0_reg[25]  ( .D(n268), .CP(clk), .CD(n362), .Q(q0[25]) );
  CFD2QXL \q0_reg[22]  ( .D(n265), .CP(clk), .CD(n363), .Q(q0[22]) );
  CFD2QXL \q0_reg[20]  ( .D(n263), .CP(clk), .CD(n363), .Q(q0[20]) );
  CFD2QXL \acc_reg[11]  ( .D(n198), .CP(clk), .CD(n368), .Q(acc[11]) );
  CFD2QXL \acc_reg[12]  ( .D(n197), .CP(clk), .CD(n368), .Q(acc[12]) );
  CFD2QXL \acc_reg[13]  ( .D(n196), .CP(clk), .CD(n368), .Q(acc[13]) );
  CFD2QXL \h0_reg[22]  ( .D(n233), .CP(clk), .CD(n365), .Q(h0[22]) );
  CFD2QXL \h0_reg[21]  ( .D(n232), .CP(clk), .CD(n365), .Q(h0[21]) );
  CFD2QXL \h0_reg[20]  ( .D(n231), .CP(clk), .CD(n365), .Q(h0[20]) );
  CFD2QXL \h0_reg[19]  ( .D(n230), .CP(clk), .CD(n365), .Q(h0[19]) );
  CFD2QXL \q0_reg[23]  ( .D(n266), .CP(clk), .CD(n362), .Q(q0[23]) );
  CFD2QXL \q0_reg[21]  ( .D(n264), .CP(clk), .CD(n363), .Q(q0[21]) );
  CFD2QXL \q0_reg[18]  ( .D(n261), .CP(clk), .CD(n363), .Q(q0[18]) );
  CFD2QXL \q0_reg[16]  ( .D(n259), .CP(clk), .CD(n363), .Q(q0[16]) );
  CFD2QXL \acc_reg[8]  ( .D(n201), .CP(clk), .CD(n367), .Q(acc[8]) );
  CFD2QXL \acc_reg[9]  ( .D(n200), .CP(clk), .CD(n368), .Q(acc[9]) );
  CFD2QXL \acc_reg[10]  ( .D(n199), .CP(clk), .CD(n368), .Q(acc[10]) );
  CFD2QXL \h0_reg[18]  ( .D(n229), .CP(clk), .CD(n365), .Q(h0[18]) );
  CFD2QXL \h0_reg[17]  ( .D(n228), .CP(clk), .CD(n365), .Q(h0[17]) );
  CFD2QXL \h0_reg[16]  ( .D(n227), .CP(clk), .CD(n365), .Q(h0[16]) );
  CFD2QXL \h0_reg[15]  ( .D(n226), .CP(clk), .CD(n366), .Q(h0[15]) );
  CFD2QXL \h0_reg[14]  ( .D(n225), .CP(clk), .CD(n366), .Q(h0[14]) );
  CFD2QXL \q0_reg[19]  ( .D(n262), .CP(clk), .CD(n363), .Q(q0[19]) );
  CFD2QXL \q0_reg[17]  ( .D(n260), .CP(clk), .CD(n363), .Q(q0[17]) );
  CFD2QXL \q0_reg[14]  ( .D(n257), .CP(clk), .CD(n363), .Q(q0[14]) );
  CFD2QXL \q0_reg[12]  ( .D(n255), .CP(clk), .CD(n363), .Q(q0[12]) );
  CFD2QXL \acc_reg[4]  ( .D(n205), .CP(clk), .CD(n367), .Q(acc[4]) );
  CFD2QXL \acc_reg[5]  ( .D(n204), .CP(clk), .CD(n367), .Q(acc[5]) );
  CFD2QXL \acc_reg[6]  ( .D(n203), .CP(clk), .CD(n367), .Q(acc[6]) );
  CFD2QXL \acc_reg[7]  ( .D(n202), .CP(clk), .CD(n367), .Q(acc[7]) );
  CFD2QXL \h0_reg[13]  ( .D(n224), .CP(clk), .CD(n366), .Q(h0[13]) );
  CFD2QXL \h0_reg[12]  ( .D(n223), .CP(clk), .CD(n366), .Q(h0[12]) );
  CFD2QXL \h0_reg[11]  ( .D(n222), .CP(clk), .CD(n366), .Q(h0[11]) );
  CFD2QXL \q0_reg[15]  ( .D(n258), .CP(clk), .CD(n363), .Q(q0[15]) );
  CFD2QXL \q0_reg[13]  ( .D(n256), .CP(clk), .CD(n363), .Q(q0[13]) );
  CFD2QXL \q0_reg[10]  ( .D(n253), .CP(clk), .CD(n363), .Q(q0[10]) );
  CFD2QXL \q0_reg[8]  ( .D(n251), .CP(clk), .CD(n364), .Q(q0[8]) );
  CFD2QXL \q0_reg[6]  ( .D(n249), .CP(clk), .CD(n364), .Q(q0[6]) );
  CFD2QXL \acc_reg[1]  ( .D(n208), .CP(clk), .CD(n367), .Q(acc[1]) );
  CFD2QXL \acc_reg[2]  ( .D(n207), .CP(clk), .CD(n367), .Q(acc[2]) );
  CFD2QXL \acc_reg[3]  ( .D(n206), .CP(clk), .CD(n367), .Q(acc[3]) );
  CFD2QXL \h0_reg[10]  ( .D(n221), .CP(clk), .CD(n366), .Q(h0[10]) );
  CFD2QXL \h0_reg[9]  ( .D(n220), .CP(clk), .CD(n366), .Q(h0[9]) );
  CFD2QXL \h0_reg[8]  ( .D(n219), .CP(clk), .CD(n366), .Q(h0[8]) );
  CFD2QXL \h0_reg[7]  ( .D(n218), .CP(clk), .CD(n366), .Q(h0[7]) );
  CFD2QXL \q0_reg[11]  ( .D(n254), .CP(clk), .CD(n363), .Q(q0[11]) );
  CFD2QXL \q0_reg[9]  ( .D(n252), .CP(clk), .CD(n364), .Q(q0[9]) );
  CFD2QXL \q0_reg[7]  ( .D(n250), .CP(clk), .CD(n364), .Q(q0[7]) );
  CFD2QXL \acc_reg[0]  ( .D(n209), .CP(clk), .CD(n367), .Q(acc[0]) );
  CFD2QXL \h0_reg[3]  ( .D(n214), .CP(clk), .CD(n366), .Q(h0[3]) );
  CFD2QXL \q0_reg[4]  ( .D(n247), .CP(clk), .CD(n364), .Q(q0[4]) );
  CFD2QXL \q0_reg[2]  ( .D(n245), .CP(clk), .CD(n364), .Q(q0[2]) );
  CFD2QXL \h0_reg[2]  ( .D(n213), .CP(clk), .CD(n367), .Q(h0[2]) );
  CFD2QXL \q0_reg[0]  ( .D(n243), .CP(clk), .CD(n364), .Q(q0[0]) );
  CFD2QXL \h0_reg[4]  ( .D(n215), .CP(clk), .CD(n366), .Q(h0[4]) );
  CFD2QXL \q0_reg[5]  ( .D(n248), .CP(clk), .CD(n364), .Q(q0[5]) );
  CFD2QXL \q0_reg[3]  ( .D(n246), .CP(clk), .CD(n364), .Q(q0[3]) );
  CFD2QXL \h0_reg[6]  ( .D(n217), .CP(clk), .CD(n366), .Q(h0[6]) );
  CFD2QXL \h0_reg[5]  ( .D(n216), .CP(clk), .CD(n366), .Q(h0[5]) );
  CFD2QXL \q0_reg[1]  ( .D(n244), .CP(clk), .CD(n364), .Q(q0[1]) );
  CFD2QXL \h0_reg[1]  ( .D(n212), .CP(clk), .CD(n367), .Q(h0[1]) );
  CFD2QXL \h0_reg[0]  ( .D(n211), .CP(clk), .CD(n367), .Q(h0[0]) );
  CFD2QXL _pushout_reg ( .D(n308), .CP(clk), .CD(n362), .Q(pushout) );
  CFD2XL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n450), .Q(cmd0[1]), .QN(
        n451) );
  CAOR2X2 U308 ( .A(q[0]), .B(n415), .C(q0[0]), .D(n447), .Z(n243) );
  CAOR2X2 U309 ( .A(h[7]), .B(n417), .C(h0[7]), .D(n434), .Z(n218) );
  CAOR2X2 U310 ( .A(h[8]), .B(n417), .C(h0[8]), .D(n435), .Z(n219) );
  CAOR2X2 U311 ( .A(h[9]), .B(n417), .C(h0[9]), .D(n435), .Z(n220) );
  CAOR2X2 U312 ( .A(h[10]), .B(n416), .C(h0[10]), .D(n436), .Z(n221) );
  CAOR2X2 U313 ( .A(h[11]), .B(n416), .C(h0[11]), .D(n436), .Z(n222) );
  CAOR2X2 U314 ( .A(h[12]), .B(n416), .C(h0[12]), .D(n437), .Z(n223) );
  CAOR2X2 U315 ( .A(h[13]), .B(n416), .C(h0[13]), .D(n437), .Z(n224) );
  CAOR2X2 U316 ( .A(h[14]), .B(n416), .C(h0[14]), .D(n438), .Z(n225) );
  CAOR2X2 U317 ( .A(h[15]), .B(n416), .C(h0[15]), .D(n438), .Z(n226) );
  CAOR2X2 U318 ( .A(h[16]), .B(n416), .C(h0[16]), .D(n439), .Z(n227) );
  CAOR2X2 U319 ( .A(h[17]), .B(n416), .C(h0[17]), .D(n439), .Z(n228) );
  CAOR2X2 U320 ( .A(h[18]), .B(n416), .C(h0[18]), .D(n440), .Z(n229) );
  CAOR2X2 U321 ( .A(h[19]), .B(n416), .C(h0[19]), .D(n440), .Z(n230) );
  CAOR2X2 U322 ( .A(h[20]), .B(n416), .C(h0[20]), .D(n441), .Z(n231) );
  CAOR2X2 U323 ( .A(h[21]), .B(n416), .C(h0[21]), .D(n441), .Z(n232) );
  CAOR2X2 U324 ( .A(h[22]), .B(n415), .C(h0[22]), .D(n442), .Z(n233) );
  CAOR2X2 U325 ( .A(h[23]), .B(n415), .C(h0[23]), .D(n442), .Z(n234) );
  CAOR2X2 U326 ( .A(h[24]), .B(n415), .C(h0[24]), .D(n443), .Z(n235) );
  CAOR2X2 U327 ( .A(h[25]), .B(n415), .C(h0[25]), .D(n443), .Z(n236) );
  CAOR2X2 U328 ( .A(h[26]), .B(n415), .C(h0[26]), .D(n444), .Z(n237) );
  CAOR2X2 U329 ( .A(h[27]), .B(n415), .C(h0[27]), .D(n444), .Z(n238) );
  CAOR2X2 U330 ( .A(h[28]), .B(n415), .C(h0[28]), .D(n445), .Z(n239) );
  CAOR2X2 U331 ( .A(h[29]), .B(n415), .C(h0[29]), .D(n445), .Z(n240) );
  CAOR2X4 U332 ( .A(acc[0]), .B(n381), .C(z[0]), .D(n382), .Z(n276) );
  CAOR2X4 U333 ( .A(acc[1]), .B(n381), .C(z[1]), .D(n382), .Z(n277) );
  CAOR2X4 U334 ( .A(acc[2]), .B(n381), .C(z[2]), .D(n383), .Z(n278) );
  CAOR2X4 U335 ( .A(acc[3]), .B(n381), .C(z[3]), .D(n383), .Z(n279) );
  CAOR2X4 U336 ( .A(acc[4]), .B(n381), .C(z[4]), .D(n384), .Z(n280) );
  CAOR2X4 U337 ( .A(acc[5]), .B(n381), .C(z[5]), .D(n384), .Z(n281) );
  CAOR2X4 U338 ( .A(acc[6]), .B(n381), .C(z[6]), .D(n384), .Z(n282) );
  CAOR2X4 U339 ( .A(acc[7]), .B(n381), .C(z[7]), .D(n383), .Z(n283) );
  CAOR2X4 U340 ( .A(acc[8]), .B(n380), .C(z[8]), .D(n385), .Z(n284) );
  CAOR2X4 U341 ( .A(acc[9]), .B(n380), .C(z[9]), .D(n385), .Z(n285) );
  CAOR2X4 U342 ( .A(acc[10]), .B(n380), .C(z[10]), .D(n386), .Z(n286) );
  CAOR2X4 U343 ( .A(acc[11]), .B(n380), .C(z[11]), .D(n386), .Z(n287) );
  CAOR2X4 U344 ( .A(acc[12]), .B(n380), .C(z[12]), .D(n386), .Z(n288) );
  CAOR2X4 U345 ( .A(acc[13]), .B(n380), .C(z[13]), .D(n385), .Z(n289) );
  CAOR2X4 U346 ( .A(acc[14]), .B(n380), .C(z[14]), .D(n387), .Z(n290) );
  CAOR2X4 U347 ( .A(acc[15]), .B(n380), .C(z[15]), .D(n387), .Z(n291) );
  CAOR2X4 U348 ( .A(acc[16]), .B(n380), .C(z[16]), .D(n388), .Z(n292) );
  CAOR2X4 U349 ( .A(acc[17]), .B(n380), .C(z[17]), .D(n388), .Z(n293) );
  CAOR2X4 U350 ( .A(acc[18]), .B(n380), .C(z[18]), .D(n388), .Z(n294) );
  CAOR2X4 U351 ( .A(acc[19]), .B(n380), .C(z[19]), .D(n387), .Z(n295) );
  CAOR2X4 U352 ( .A(acc[20]), .B(n379), .C(z[20]), .D(n389), .Z(n296) );
  CAOR2X4 U353 ( .A(acc[21]), .B(n379), .C(z[21]), .D(n389), .Z(n297) );
  CAOR2X4 U354 ( .A(acc[22]), .B(n379), .C(z[22]), .D(n390), .Z(n298) );
  CAOR2X4 U355 ( .A(acc[23]), .B(n379), .C(z[23]), .D(n390), .Z(n299) );
  CAOR2X4 U356 ( .A(acc[24]), .B(n379), .C(z[24]), .D(n390), .Z(n300) );
  CAOR2X4 U357 ( .A(acc[25]), .B(n379), .C(z[25]), .D(n389), .Z(n301) );
  CAOR2X4 U358 ( .A(acc[26]), .B(n379), .C(z[26]), .D(n391), .Z(n302) );
  CAOR2X4 U359 ( .A(acc[27]), .B(n379), .C(z[27]), .D(n391), .Z(n303) );
  CAOR2X4 U360 ( .A(acc[28]), .B(n379), .C(z[28]), .D(n392), .Z(n304) );
  CAOR2X4 U361 ( .A(acc[29]), .B(n379), .C(z[29]), .D(n392), .Z(n305) );
  CAOR2X4 U362 ( .A(acc[30]), .B(n379), .C(z[30]), .D(n392), .Z(n306) );
  CAOR2X4 U363 ( .A(acc[31]), .B(n379), .C(z[31]), .D(n391), .Z(n307) );
  CNIVX1 U364 ( .A(_pushout_d), .Z(n308) );
  CIVX2 U365 ( .A(n406), .Z(n405) );
  CIVX2 U366 ( .A(n400), .Z(n398) );
  CIVX2 U367 ( .A(n400), .Z(n397) );
  CIVX2 U368 ( .A(n400), .Z(n395) );
  CIVX2 U369 ( .A(n400), .Z(n396) );
  CIVX2 U370 ( .A(n406), .Z(n403) );
  CIVX2 U371 ( .A(n406), .Z(n402) );
  CNR2X1 U372 ( .A(n581), .B(n351), .Z(n658) );
  CNR2X1 U373 ( .A(n537), .B(n354), .Z(n672) );
  CNR2X1 U374 ( .A(n596), .B(n355), .Z(n665) );
  CNR2X1 U375 ( .A(n613), .B(n352), .Z(n651) );
  CNR2X1 U376 ( .A(n600), .B(n358), .Z(n717) );
  CIVX2 U377 ( .A(n400), .Z(n394) );
  CIVX2 U378 ( .A(n406), .Z(n401) );
  CND2X1 U379 ( .A(n519), .B(n400), .Z(n537) );
  CND2X1 U380 ( .A(n565), .B(n400), .Z(n596) );
  CND2X1 U381 ( .A(n672), .B(n406), .Z(n600) );
  CIVX2 U382 ( .A(n406), .Z(n404) );
  CND2X1 U383 ( .A(n658), .B(n406), .Z(n711) );
  CND2X1 U384 ( .A(n651), .B(n406), .Z(n695) );
  CND2X1 U385 ( .A(n644), .B(n406), .Z(n691) );
  CND2X1 U386 ( .A(n627), .B(n406), .Z(n687) );
  CND2X1 U387 ( .A(n620), .B(n406), .Z(n683) );
  CND2X1 U388 ( .A(n679), .B(n406), .Z(n744) );
  CNR2X1 U389 ( .A(n725), .B(n361), .Z(n765) );
  CNR2X1 U390 ( .A(n723), .B(n357), .Z(n764) );
  CNR2X1 U391 ( .A(n721), .B(n361), .Z(n763) );
  CNR2X1 U392 ( .A(n706), .B(n356), .Z(n762) );
  CNR2X1 U393 ( .A(n637), .B(n357), .Z(n753) );
  CND2X1 U394 ( .A(n665), .B(n406), .Z(n715) );
  CNR2X1 U395 ( .A(n691), .B(n356), .Z(n780) );
  CNR2X1 U396 ( .A(n687), .B(n360), .Z(n771) );
  CNR2X1 U397 ( .A(n683), .B(n356), .Z(n770) );
  CNR2X1 U398 ( .A(n744), .B(n357), .Z(n769) );
  CNR2X1 U399 ( .A(n742), .B(n358), .Z(n768) );
  CNR2X1 U400 ( .A(n729), .B(n359), .Z(n767) );
  CNR2X1 U401 ( .A(n727), .B(n360), .Z(n766) );
  CNR3XL U402 ( .A(n464), .B(n411), .C(n409), .Z(N241) );
  CNR2X1 U403 ( .A(n711), .B(n360), .Z(n782) );
  CNR2X1 U404 ( .A(n715), .B(n359), .Z(n783) );
  CNR2X1 U405 ( .A(n695), .B(n361), .Z(n781) );
  CNR3XL U406 ( .A(n478), .B(n413), .C(n409), .Z(N243) );
  CNR3XL U407 ( .A(n475), .B(n413), .C(n409), .Z(N242) );
  CNR3XL U408 ( .A(n484), .B(n413), .C(n408), .Z(N249) );
  CNR3XL U409 ( .A(n483), .B(n412), .C(n408), .Z(N248) );
  CNR3XL U410 ( .A(n482), .B(n413), .C(n409), .Z(N247) );
  CNR3XL U411 ( .A(n481), .B(n413), .C(n409), .Z(N246) );
  CNR3XL U412 ( .A(n480), .B(n413), .C(n409), .Z(N245) );
  CNR3XL U413 ( .A(n454), .B(n412), .C(n408), .Z(N250) );
  CNR3XL U414 ( .A(n479), .B(n413), .C(n409), .Z(N244) );
  CNR3XL U415 ( .A(n461), .B(n412), .C(n408), .Z(N257) );
  CNR3XL U416 ( .A(n460), .B(n412), .C(n408), .Z(N256) );
  CNR3XL U417 ( .A(n459), .B(n412), .C(n408), .Z(N255) );
  CNR3XL U418 ( .A(n458), .B(n412), .C(n408), .Z(N254) );
  CNR3XL U419 ( .A(n457), .B(n412), .C(n408), .Z(N253) );
  CNR3XL U420 ( .A(n456), .B(n412), .C(n408), .Z(N252) );
  CNR3XL U421 ( .A(n455), .B(n412), .C(n408), .Z(N251) );
  CNR3XL U422 ( .A(n469), .B(n411), .C(n407), .Z(N264) );
  CNR3XL U423 ( .A(n468), .B(n411), .C(n407), .Z(N263) );
  CNR3XL U424 ( .A(n467), .B(n411), .C(n407), .Z(N262) );
  CNR3XL U425 ( .A(n466), .B(n412), .C(n407), .Z(N261) );
  CNR3XL U426 ( .A(n465), .B(n411), .C(n407), .Z(N260) );
  CNR3XL U427 ( .A(n463), .B(n412), .C(n408), .Z(N259) );
  CNR3XL U428 ( .A(n462), .B(n412), .C(n408), .Z(N258) );
  CNR3XL U429 ( .A(n476), .B(n411), .C(n407), .Z(N270) );
  CNR3XL U430 ( .A(n473), .B(n411), .C(n407), .Z(N268) );
  CNR3XL U431 ( .A(n472), .B(n411), .C(n407), .Z(N267) );
  CNR3XL U432 ( .A(n471), .B(n411), .C(n407), .Z(N266) );
  CNR3XL U433 ( .A(n470), .B(n411), .C(n407), .Z(N265) );
  CNR3XL U434 ( .A(n474), .B(n411), .C(n407), .Z(N269) );
  CNR4X1 U435 ( .A(n375), .B(n11), .C(n12), .D(n13), .Z(n8) );
  CNR2X1 U436 ( .A(n413), .B(n784), .Z(N272) );
  CNIVX1 U437 ( .A(n453), .Z(n375) );
  CNIVX1 U438 ( .A(n337), .Z(n339) );
  CNIVX1 U439 ( .A(n337), .Z(n340) );
  CNIVX1 U440 ( .A(n337), .Z(n341) );
  CNIVX1 U441 ( .A(n337), .Z(n342) );
  CNR3XL U442 ( .A(n477), .B(n411), .C(n407), .Z(N271) );
  CNR3XL U443 ( .A(n375), .B(n451), .C(n452), .Z(_pushout_d) );
  CNIVX1 U444 ( .A(n453), .Z(n377) );
  CNIVX1 U445 ( .A(n453), .Z(n376) );
  CNIVX1 U446 ( .A(n323), .Z(n325) );
  CNIVX1 U447 ( .A(n309), .Z(n311) );
  CNIVX1 U448 ( .A(n323), .Z(n326) );
  CNIVX1 U449 ( .A(n309), .Z(n312) );
  CNIVX1 U450 ( .A(n323), .Z(n327) );
  CNIVX1 U451 ( .A(n309), .Z(n313) );
  CNIVX1 U452 ( .A(n323), .Z(n328) );
  CNIVX1 U453 ( .A(n309), .Z(n314) );
  CNIVX1 U454 ( .A(n338), .Z(n343) );
  CNIVX1 U455 ( .A(n338), .Z(n344) );
  CNIVX1 U456 ( .A(n338), .Z(n345) );
  CNIVX1 U457 ( .A(n338), .Z(n346) );
  CNIVX1 U458 ( .A(n17), .Z(n347) );
  CNIVX1 U459 ( .A(n17), .Z(n348) );
  CNIVX1 U460 ( .A(n17), .Z(n349) );
  CNIVX1 U461 ( .A(n17), .Z(n350) );
  CNIVX1 U462 ( .A(n324), .Z(n329) );
  CNIVX1 U463 ( .A(n310), .Z(n315) );
  CNIVX1 U464 ( .A(n324), .Z(n330) );
  CNIVX1 U465 ( .A(n310), .Z(n316) );
  CNIVX1 U466 ( .A(n324), .Z(n331) );
  CNIVX1 U467 ( .A(n310), .Z(n317) );
  CNIVX1 U468 ( .A(n324), .Z(n332) );
  CNIVX1 U469 ( .A(n310), .Z(n318) );
  CNIVX1 U470 ( .A(n16), .Z(n333) );
  CNIVX1 U471 ( .A(n18), .Z(n319) );
  CNIVX1 U472 ( .A(n18), .Z(n320) );
  CNIVX1 U473 ( .A(n16), .Z(n334) );
  CNIVX1 U474 ( .A(n18), .Z(n321) );
  CNIVX1 U475 ( .A(n16), .Z(n335) );
  CNIVX1 U476 ( .A(n16), .Z(n336) );
  CNIVX1 U477 ( .A(n18), .Z(n322) );
  CNIVX1 U478 ( .A(n450), .Z(n373) );
  CNIVX1 U479 ( .A(n450), .Z(n372) );
  CNIVX1 U480 ( .A(n450), .Z(n371) );
  CNIVX1 U481 ( .A(n450), .Z(n370) );
  CNIVX1 U482 ( .A(n450), .Z(n369) );
  CNIVX1 U483 ( .A(n450), .Z(n368) );
  CNIVX1 U484 ( .A(n450), .Z(n367) );
  CNIVX1 U485 ( .A(n450), .Z(n366) );
  CNIVX1 U486 ( .A(n450), .Z(n365) );
  CNIVX1 U487 ( .A(n450), .Z(n364) );
  CNIVX1 U488 ( .A(n450), .Z(n363) );
  CNIVX1 U489 ( .A(n450), .Z(n362) );
  CNIVX1 U490 ( .A(n450), .Z(n374) );
  CND2X1 U491 ( .A(n143), .B(n144), .Z(n210) );
  CANR2X1 U492 ( .A(N336), .B(n322), .C(acc[63]), .D(n375), .Z(n143) );
  CANR2X1 U493 ( .A(N79), .B(n336), .C(N207), .D(n350), .Z(n144) );
  CNIVX1 U494 ( .A(h0[5]), .Z(n410) );
  CNIVX1 U495 ( .A(h0[2]), .Z(n353) );
  CNIVX1 U496 ( .A(h0[4]), .Z(n356) );
  CND2X1 U497 ( .A(n14), .B(n15), .Z(n147) );
  CANR2X1 U498 ( .A(N335), .B(n311), .C(acc[62]), .D(n375), .Z(n14) );
  CANR2X1 U499 ( .A(N78), .B(n325), .C(N206), .D(n339), .Z(n15) );
  CND2X1 U500 ( .A(n19), .B(n20), .Z(n148) );
  CANR2X1 U501 ( .A(N334), .B(n312), .C(acc[61]), .D(n378), .Z(n19) );
  CANR2X1 U502 ( .A(N77), .B(n326), .C(N205), .D(n340), .Z(n20) );
  CNIVX1 U503 ( .A(n453), .Z(n378) );
  CND2X1 U504 ( .A(n21), .B(n22), .Z(n149) );
  CANR2X1 U505 ( .A(N333), .B(n313), .C(acc[60]), .D(n377), .Z(n21) );
  CANR2X1 U506 ( .A(N76), .B(n327), .C(N204), .D(n341), .Z(n22) );
  CND2X1 U507 ( .A(n23), .B(n24), .Z(n150) );
  CANR2X1 U508 ( .A(N332), .B(n314), .C(acc[59]), .D(n377), .Z(n23) );
  CANR2X1 U509 ( .A(N75), .B(n328), .C(N203), .D(n342), .Z(n24) );
  CNIVX1 U510 ( .A(h0[6]), .Z(n414) );
  CND2X1 U511 ( .A(n25), .B(n26), .Z(n151) );
  CANR2X1 U512 ( .A(N331), .B(n311), .C(acc[58]), .D(n377), .Z(n25) );
  CANR2X1 U513 ( .A(N74), .B(n325), .C(N202), .D(n339), .Z(n26) );
  CND2X1 U514 ( .A(n27), .B(n28), .Z(n152) );
  CANR2X1 U515 ( .A(N330), .B(n312), .C(acc[57]), .D(n377), .Z(n27) );
  CANR2X1 U516 ( .A(N73), .B(n326), .C(N201), .D(n340), .Z(n28) );
  CND2X1 U517 ( .A(n29), .B(n30), .Z(n153) );
  CANR2X1 U518 ( .A(N329), .B(n313), .C(acc[56]), .D(n377), .Z(n29) );
  CANR2X1 U519 ( .A(N72), .B(n327), .C(N200), .D(n341), .Z(n30) );
  CND2X1 U520 ( .A(n31), .B(n32), .Z(n154) );
  CANR2X1 U521 ( .A(N328), .B(n314), .C(acc[55]), .D(n377), .Z(n31) );
  CANR2X1 U522 ( .A(N71), .B(n328), .C(N199), .D(n342), .Z(n32) );
  CND2X1 U523 ( .A(n33), .B(n34), .Z(n155) );
  CANR2X1 U524 ( .A(N327), .B(n315), .C(acc[54]), .D(n377), .Z(n33) );
  CANR2X1 U525 ( .A(N70), .B(n329), .C(N198), .D(n343), .Z(n34) );
  CND2X1 U526 ( .A(n35), .B(n36), .Z(n156) );
  CANR2X1 U527 ( .A(N326), .B(n316), .C(acc[53]), .D(n377), .Z(n35) );
  CANR2X1 U528 ( .A(N69), .B(n330), .C(N197), .D(n344), .Z(n36) );
  CND2X1 U529 ( .A(n37), .B(n38), .Z(n157) );
  CANR2X1 U530 ( .A(N325), .B(n317), .C(acc[52]), .D(n377), .Z(n37) );
  CANR2X1 U531 ( .A(N68), .B(n331), .C(N196), .D(n345), .Z(n38) );
  CND2X1 U532 ( .A(n39), .B(n40), .Z(n158) );
  CANR2X1 U533 ( .A(N324), .B(n318), .C(acc[51]), .D(n377), .Z(n39) );
  CANR2X1 U534 ( .A(N67), .B(n332), .C(N195), .D(n346), .Z(n40) );
  CND2X1 U535 ( .A(n41), .B(n42), .Z(n159) );
  CANR2X1 U536 ( .A(N323), .B(n315), .C(acc[50]), .D(n377), .Z(n41) );
  CANR2X1 U537 ( .A(N66), .B(n329), .C(N194), .D(n343), .Z(n42) );
  CND2X1 U538 ( .A(n43), .B(n44), .Z(n160) );
  CANR2X1 U539 ( .A(N322), .B(n316), .C(acc[49]), .D(n377), .Z(n43) );
  CANR2X1 U540 ( .A(N65), .B(n330), .C(N193), .D(n344), .Z(n44) );
  CND2X1 U541 ( .A(n49), .B(n50), .Z(n163) );
  CANR2X1 U542 ( .A(N319), .B(n319), .C(acc[46]), .D(n377), .Z(n49) );
  CANR2X1 U543 ( .A(N62), .B(n333), .C(N190), .D(n347), .Z(n50) );
  CND2X1 U544 ( .A(n45), .B(n46), .Z(n161) );
  CANR2X1 U545 ( .A(N321), .B(n317), .C(acc[48]), .D(n377), .Z(n45) );
  CANR2X1 U546 ( .A(N64), .B(n331), .C(N192), .D(n345), .Z(n46) );
  CND2X1 U547 ( .A(n47), .B(n48), .Z(n162) );
  CANR2X1 U548 ( .A(N320), .B(n318), .C(acc[47]), .D(n377), .Z(n47) );
  CANR2X1 U549 ( .A(N63), .B(n332), .C(N191), .D(n346), .Z(n48) );
  CND2X1 U550 ( .A(n51), .B(n52), .Z(n164) );
  CANR2X1 U551 ( .A(N318), .B(n320), .C(acc[45]), .D(n377), .Z(n51) );
  CANR2X1 U552 ( .A(N61), .B(n334), .C(N189), .D(n348), .Z(n52) );
  CND2X1 U553 ( .A(n57), .B(n58), .Z(n167) );
  CANR2X1 U554 ( .A(N315), .B(n311), .C(acc[42]), .D(n377), .Z(n57) );
  CANR2X1 U555 ( .A(N58), .B(n325), .C(N186), .D(n339), .Z(n58) );
  CND2X1 U556 ( .A(n53), .B(n54), .Z(n165) );
  CANR2X1 U557 ( .A(N317), .B(n321), .C(acc[44]), .D(n377), .Z(n53) );
  CANR2X1 U558 ( .A(N60), .B(n335), .C(N188), .D(n349), .Z(n54) );
  CND2X1 U559 ( .A(n55), .B(n56), .Z(n166) );
  CANR2X1 U560 ( .A(N316), .B(n322), .C(acc[43]), .D(n377), .Z(n55) );
  CANR2X1 U561 ( .A(N59), .B(n336), .C(N187), .D(n350), .Z(n56) );
  CND2X1 U562 ( .A(n59), .B(n60), .Z(n168) );
  CANR2X1 U563 ( .A(N314), .B(n312), .C(acc[41]), .D(n377), .Z(n59) );
  CANR2X1 U564 ( .A(N57), .B(n326), .C(N185), .D(n340), .Z(n60) );
  CND2X1 U565 ( .A(n61), .B(n62), .Z(n169) );
  CANR2X1 U566 ( .A(N313), .B(n313), .C(acc[40]), .D(n377), .Z(n61) );
  CANR2X1 U567 ( .A(N56), .B(n327), .C(N184), .D(n341), .Z(n62) );
  CND2X1 U568 ( .A(n63), .B(n64), .Z(n170) );
  CANR2X1 U569 ( .A(N312), .B(n314), .C(acc[39]), .D(n377), .Z(n63) );
  CANR2X1 U570 ( .A(N55), .B(n328), .C(N183), .D(n342), .Z(n64) );
  CND2X1 U571 ( .A(n65), .B(n66), .Z(n171) );
  CANR2X1 U572 ( .A(N311), .B(n319), .C(acc[38]), .D(n376), .Z(n65) );
  CANR2X1 U573 ( .A(N54), .B(n333), .C(N182), .D(n347), .Z(n66) );
  CND2X1 U574 ( .A(n67), .B(n68), .Z(n172) );
  CANR2X1 U575 ( .A(N310), .B(n320), .C(acc[37]), .D(n376), .Z(n67) );
  CANR2X1 U576 ( .A(N53), .B(n334), .C(N181), .D(n348), .Z(n68) );
  CND2X1 U577 ( .A(n69), .B(n70), .Z(n173) );
  CANR2X1 U578 ( .A(N309), .B(n321), .C(acc[36]), .D(n376), .Z(n69) );
  CANR2X1 U579 ( .A(N52), .B(n335), .C(N180), .D(n349), .Z(n70) );
  CND2X1 U580 ( .A(n71), .B(n72), .Z(n174) );
  CANR2X1 U581 ( .A(N308), .B(n322), .C(acc[35]), .D(n376), .Z(n71) );
  CANR2X1 U582 ( .A(N51), .B(n336), .C(N179), .D(n350), .Z(n72) );
  CIVX2 U583 ( .A(h0[0]), .Z(n485) );
  CND2X1 U584 ( .A(n73), .B(n74), .Z(n175) );
  CANR2X1 U585 ( .A(N307), .B(n315), .C(acc[34]), .D(n376), .Z(n73) );
  CANR2X1 U586 ( .A(N50), .B(n329), .C(N178), .D(n343), .Z(n74) );
  CND2X1 U587 ( .A(n75), .B(n76), .Z(n176) );
  CANR2X1 U588 ( .A(N306), .B(n316), .C(acc[33]), .D(n376), .Z(n75) );
  CANR2X1 U589 ( .A(N49), .B(n330), .C(N177), .D(n344), .Z(n76) );
  CAN2X1 U590 ( .A(acc[0]), .B(h0[0]), .Z(n486) );
  CND2X1 U591 ( .A(n77), .B(n78), .Z(n177) );
  CANR2X1 U592 ( .A(N305), .B(n317), .C(acc[32]), .D(n376), .Z(n77) );
  CANR2X1 U593 ( .A(N48), .B(n331), .C(N176), .D(n345), .Z(n78) );
  CND2X1 U594 ( .A(n81), .B(n82), .Z(n179) );
  CANR2X1 U595 ( .A(N303), .B(n319), .C(acc[30]), .D(n376), .Z(n81) );
  CANR2X1 U596 ( .A(N46), .B(n333), .C(N174), .D(n347), .Z(n82) );
  CND2X1 U597 ( .A(n83), .B(n84), .Z(n180) );
  CANR2X1 U598 ( .A(N302), .B(n320), .C(acc[29]), .D(n376), .Z(n83) );
  CANR2X1 U599 ( .A(N45), .B(n334), .C(N173), .D(n348), .Z(n84) );
  CNIVX1 U600 ( .A(h0[2]), .Z(n352) );
  CNIVX1 U601 ( .A(h0[2]), .Z(n351) );
  CNIVX1 U602 ( .A(h0[2]), .Z(n355) );
  CNIVX1 U603 ( .A(h0[2]), .Z(n354) );
  CNIVX1 U604 ( .A(h0[4]), .Z(n360) );
  CNIVX1 U605 ( .A(h0[4]), .Z(n357) );
  CNIVX1 U606 ( .A(h0[4]), .Z(n358) );
  CNIVX1 U607 ( .A(h0[4]), .Z(n359) );
  CNIVX1 U608 ( .A(h0[5]), .Z(n409) );
  CNR2IX1 U609 ( .B(acc[63]), .A(h0[0]), .Z(n519) );
  CNIVX1 U610 ( .A(h0[6]), .Z(n413) );
  CND2X1 U611 ( .A(n79), .B(n80), .Z(n178) );
  CANR2X1 U612 ( .A(N304), .B(n318), .C(acc[31]), .D(n376), .Z(n79) );
  CANR2X1 U613 ( .A(N47), .B(n332), .C(N175), .D(n346), .Z(n80) );
  CND2X1 U614 ( .A(n85), .B(n86), .Z(n181) );
  CANR2X1 U615 ( .A(N301), .B(n321), .C(acc[28]), .D(n376), .Z(n85) );
  CANR2X1 U616 ( .A(N44), .B(n335), .C(N172), .D(n349), .Z(n86) );
  CND2X1 U617 ( .A(n89), .B(n90), .Z(n183) );
  CANR2X1 U618 ( .A(N299), .B(n311), .C(acc[26]), .D(n376), .Z(n89) );
  CANR2X1 U619 ( .A(N42), .B(n325), .C(N170), .D(n339), .Z(n90) );
  CND2X1 U620 ( .A(n91), .B(n92), .Z(n184) );
  CANR2X1 U621 ( .A(N298), .B(n312), .C(acc[25]), .D(n376), .Z(n91) );
  CANR2X1 U622 ( .A(N41), .B(n326), .C(N169), .D(n340), .Z(n92) );
  CNIVX1 U623 ( .A(h0[4]), .Z(n361) );
  CND2X1 U624 ( .A(n87), .B(n88), .Z(n182) );
  CANR2X1 U625 ( .A(N300), .B(n322), .C(acc[27]), .D(n376), .Z(n87) );
  CANR2X1 U626 ( .A(N43), .B(n336), .C(N171), .D(n350), .Z(n88) );
  CND2X1 U627 ( .A(n97), .B(n98), .Z(n187) );
  CANR2X1 U628 ( .A(N295), .B(n311), .C(acc[22]), .D(n376), .Z(n97) );
  CANR2X1 U629 ( .A(N38), .B(n325), .C(N166), .D(n339), .Z(n98) );
  CND2X1 U630 ( .A(n99), .B(n100), .Z(n188) );
  CANR2X1 U631 ( .A(N294), .B(n312), .C(acc[21]), .D(n376), .Z(n99) );
  CANR2X1 U632 ( .A(N37), .B(n326), .C(N165), .D(n340), .Z(n100) );
  CND2X1 U633 ( .A(n93), .B(n94), .Z(n185) );
  CANR2X1 U634 ( .A(N297), .B(n313), .C(acc[24]), .D(n376), .Z(n93) );
  CANR2X1 U635 ( .A(N40), .B(n327), .C(N168), .D(n341), .Z(n94) );
  CND2X1 U636 ( .A(n95), .B(n96), .Z(n186) );
  CANR2X1 U637 ( .A(N296), .B(n314), .C(acc[23]), .D(n376), .Z(n95) );
  CANR2X1 U638 ( .A(N39), .B(n328), .C(N167), .D(n342), .Z(n96) );
  CND2X1 U639 ( .A(n105), .B(n106), .Z(n191) );
  CANR2X1 U640 ( .A(N291), .B(n315), .C(acc[18]), .D(n376), .Z(n105) );
  CANR2X1 U641 ( .A(N34), .B(n329), .C(N162), .D(n343), .Z(n106) );
  CND2X1 U642 ( .A(n101), .B(n102), .Z(n189) );
  CANR2X1 U643 ( .A(N293), .B(n313), .C(acc[20]), .D(n376), .Z(n101) );
  CANR2X1 U644 ( .A(N36), .B(n327), .C(N164), .D(n341), .Z(n102) );
  CND2X1 U645 ( .A(n103), .B(n104), .Z(n190) );
  CANR2X1 U646 ( .A(N292), .B(n314), .C(acc[19]), .D(n376), .Z(n103) );
  CANR2X1 U647 ( .A(N35), .B(n328), .C(N163), .D(n342), .Z(n104) );
  CND2X1 U648 ( .A(n107), .B(n108), .Z(n192) );
  CANR2X1 U649 ( .A(N290), .B(n316), .C(acc[17]), .D(n375), .Z(n107) );
  CANR2X1 U650 ( .A(N33), .B(n330), .C(N161), .D(n344), .Z(n108) );
  CND2X1 U651 ( .A(n113), .B(n114), .Z(n195) );
  CANR2X1 U652 ( .A(N287), .B(n315), .C(acc[14]), .D(n376), .Z(n113) );
  CANR2X1 U653 ( .A(N30), .B(n329), .C(N158), .D(n343), .Z(n114) );
  CND2X1 U654 ( .A(n109), .B(n110), .Z(n193) );
  CANR2X1 U655 ( .A(N289), .B(n317), .C(acc[16]), .D(n375), .Z(n109) );
  CANR2X1 U656 ( .A(N32), .B(n331), .C(N160), .D(n345), .Z(n110) );
  CND2X1 U657 ( .A(n111), .B(n112), .Z(n194) );
  CANR2X1 U658 ( .A(N288), .B(n318), .C(acc[15]), .D(n375), .Z(n111) );
  CANR2X1 U659 ( .A(N31), .B(n332), .C(N159), .D(n346), .Z(n112) );
  CND2X1 U660 ( .A(n115), .B(n116), .Z(n196) );
  CANR2X1 U661 ( .A(N286), .B(n316), .C(acc[13]), .D(n375), .Z(n115) );
  CANR2X1 U662 ( .A(N29), .B(n330), .C(N157), .D(n344), .Z(n116) );
  CNIVX1 U663 ( .A(h0[6]), .Z(n411) );
  CND2X1 U664 ( .A(n117), .B(n118), .Z(n197) );
  CANR2X1 U665 ( .A(N285), .B(n317), .C(acc[12]), .D(n375), .Z(n117) );
  CANR2X1 U666 ( .A(N28), .B(n331), .C(N156), .D(n345), .Z(n118) );
  CND2X1 U667 ( .A(n119), .B(n120), .Z(n198) );
  CANR2X1 U668 ( .A(N284), .B(n318), .C(acc[11]), .D(n375), .Z(n119) );
  CANR2X1 U669 ( .A(N27), .B(n332), .C(N155), .D(n346), .Z(n120) );
  CNIVX1 U670 ( .A(h0[5]), .Z(n408) );
  CNIVX1 U671 ( .A(h0[6]), .Z(n412) );
  CND2X1 U672 ( .A(n121), .B(n122), .Z(n199) );
  CANR2X1 U673 ( .A(N283), .B(n319), .C(acc[10]), .D(n375), .Z(n121) );
  CANR2X1 U674 ( .A(N26), .B(n333), .C(N154), .D(n347), .Z(n122) );
  CND2X1 U675 ( .A(n123), .B(n124), .Z(n200) );
  CANR2X1 U676 ( .A(N282), .B(n320), .C(acc[9]), .D(n375), .Z(n123) );
  CANR2X1 U677 ( .A(N25), .B(n334), .C(N153), .D(n348), .Z(n124) );
  CND2X1 U678 ( .A(n125), .B(n126), .Z(n201) );
  CANR2X1 U679 ( .A(N281), .B(n321), .C(acc[8]), .D(n375), .Z(n125) );
  CANR2X1 U680 ( .A(N24), .B(n335), .C(N152), .D(n349), .Z(n126) );
  CND2X1 U681 ( .A(n127), .B(n128), .Z(n202) );
  CANR2X1 U682 ( .A(N280), .B(n322), .C(acc[7]), .D(n375), .Z(n127) );
  CANR2X1 U683 ( .A(N23), .B(n336), .C(N151), .D(n350), .Z(n128) );
  CND2X1 U684 ( .A(n131), .B(n132), .Z(n204) );
  CANR2X1 U685 ( .A(N278), .B(n312), .C(acc[5]), .D(n375), .Z(n131) );
  CANR2X1 U686 ( .A(N21), .B(n326), .C(N149), .D(n340), .Z(n132) );
  CND2X1 U687 ( .A(n129), .B(n130), .Z(n203) );
  CANR2X1 U688 ( .A(N279), .B(n311), .C(acc[6]), .D(n375), .Z(n129) );
  CANR2X1 U689 ( .A(N22), .B(n325), .C(N150), .D(n339), .Z(n130) );
  CND2X1 U690 ( .A(n133), .B(n134), .Z(n205) );
  CANR2X1 U691 ( .A(N277), .B(n313), .C(acc[4]), .D(n375), .Z(n133) );
  CANR2X1 U692 ( .A(N20), .B(n327), .C(N148), .D(n341), .Z(n134) );
  CND2X1 U693 ( .A(n141), .B(n142), .Z(n209) );
  CANR2X1 U694 ( .A(N16), .B(n335), .C(N144), .D(n349), .Z(n142) );
  CANR2X1 U695 ( .A(N273), .B(n321), .C(acc[0]), .D(n375), .Z(n141) );
  CNIVX1 U696 ( .A(h0[5]), .Z(n407) );
  CND2X1 U697 ( .A(n135), .B(n136), .Z(n206) );
  CANR2X1 U698 ( .A(N276), .B(n314), .C(acc[3]), .D(n375), .Z(n135) );
  CANR2X1 U699 ( .A(N19), .B(n328), .C(N147), .D(n342), .Z(n136) );
  CND2X1 U700 ( .A(n137), .B(n138), .Z(n207) );
  CANR2X1 U701 ( .A(N275), .B(n319), .C(acc[2]), .D(n375), .Z(n137) );
  CANR2X1 U702 ( .A(N18), .B(n333), .C(N146), .D(n347), .Z(n138) );
  CND2X1 U703 ( .A(n139), .B(n140), .Z(n208) );
  CANR2X1 U704 ( .A(N17), .B(n334), .C(N145), .D(n348), .Z(n140) );
  CANR2X1 U705 ( .A(N274), .B(n320), .C(acc[1]), .D(n375), .Z(n139) );
  CNR2X1 U706 ( .A(n451), .B(cmd0[0]), .Z(n13) );
  CNR2X1 U707 ( .A(n452), .B(cmd0[1]), .Z(n12) );
  CNR2X1 U708 ( .A(cmd0[0]), .B(cmd0[1]), .Z(n11) );
  CAN2X1 U709 ( .A(n12), .B(push0), .Z(n337) );
  CAN2X1 U710 ( .A(n12), .B(push0), .Z(n338) );
  CAN2X1 U711 ( .A(n11), .B(push0), .Z(n324) );
  CAN2X1 U712 ( .A(n13), .B(push0), .Z(n310) );
  CAN2X1 U713 ( .A(n11), .B(push0), .Z(n323) );
  CAN2X1 U714 ( .A(n13), .B(push0), .Z(n309) );
  CAN2X1 U715 ( .A(n12), .B(push0), .Z(n17) );
  CAN2X1 U716 ( .A(n11), .B(push0), .Z(n16) );
  CAN2X1 U717 ( .A(n13), .B(push0), .Z(n18) );
  CIVX2 U718 ( .A(rst), .Z(n450) );
  CIVX2 U719 ( .A(n393), .Z(n379) );
  CIVX2 U720 ( .A(n393), .Z(n380) );
  CIVX2 U721 ( .A(n448), .Z(n415) );
  CIVX2 U722 ( .A(n448), .Z(n416) );
  CIVX2 U723 ( .A(n448), .Z(n417) );
  CIVX2 U724 ( .A(n449), .Z(n418) );
  CIVX2 U725 ( .A(n449), .Z(n419) );
  CIVXL U726 ( .A(n393), .Z(n381) );
  CIVXL U727 ( .A(n8), .Z(n382) );
  CIVXL U728 ( .A(n8), .Z(n383) );
  CIVXL U729 ( .A(n8), .Z(n384) );
  CIVXL U730 ( .A(n8), .Z(n385) );
  CIVXL U731 ( .A(n8), .Z(n386) );
  CIVXL U732 ( .A(n8), .Z(n387) );
  CIVXL U733 ( .A(n8), .Z(n388) );
  CIVXL U734 ( .A(n8), .Z(n389) );
  CIVXL U735 ( .A(n8), .Z(n390) );
  CIVXL U736 ( .A(n8), .Z(n391) );
  CIVXL U737 ( .A(n8), .Z(n392) );
  CIVXL U738 ( .A(n8), .Z(n393) );
  CIVXL U739 ( .A(n400), .Z(n399) );
  CIVX2 U740 ( .A(h0[1]), .Z(n400) );
  CIVX2 U741 ( .A(h0[3]), .Z(n406) );
  CIVXL U742 ( .A(n449), .Z(n420) );
  CIVXL U743 ( .A(pushin), .Z(n421) );
  CIVXL U744 ( .A(pushin), .Z(n422) );
  CIVXL U745 ( .A(pushin), .Z(n423) );
  CIVXL U746 ( .A(pushin), .Z(n424) );
  CIVXL U747 ( .A(pushin), .Z(n425) );
  CIVXL U748 ( .A(pushin), .Z(n426) );
  CIVXL U749 ( .A(pushin), .Z(n427) );
  CIVXL U750 ( .A(pushin), .Z(n428) );
  CIVXL U751 ( .A(pushin), .Z(n429) );
  CIVXL U752 ( .A(pushin), .Z(n430) );
  CIVXL U753 ( .A(pushin), .Z(n431) );
  CIVXL U754 ( .A(pushin), .Z(n432) );
  CIVXL U755 ( .A(pushin), .Z(n433) );
  CIVXL U756 ( .A(pushin), .Z(n434) );
  CIVXL U757 ( .A(pushin), .Z(n435) );
  CIVXL U758 ( .A(pushin), .Z(n436) );
  CIVXL U759 ( .A(pushin), .Z(n437) );
  CIVXL U760 ( .A(pushin), .Z(n438) );
  CIVXL U761 ( .A(pushin), .Z(n439) );
  CIVXL U762 ( .A(pushin), .Z(n440) );
  CIVXL U763 ( .A(pushin), .Z(n441) );
  CIVXL U764 ( .A(pushin), .Z(n442) );
  CIVXL U765 ( .A(pushin), .Z(n443) );
  CIVXL U766 ( .A(pushin), .Z(n444) );
  CIVXL U767 ( .A(pushin), .Z(n445) );
  CIVXL U768 ( .A(pushin), .Z(n446) );
  CIVXL U769 ( .A(pushin), .Z(n447) );
  CIVXL U770 ( .A(pushin), .Z(n448) );
  CIVXL U771 ( .A(pushin), .Z(n449) );
  CIVX2 U772 ( .A(cmd0[0]), .Z(n452) );
  CIVX2 U773 ( .A(push0), .Z(n453) );
  CIVX2 U774 ( .A(n746), .Z(n454) );
  CIVX2 U775 ( .A(n747), .Z(n455) );
  CIVX2 U776 ( .A(n748), .Z(n456) );
  CIVX2 U777 ( .A(n749), .Z(n457) );
  CIVX2 U778 ( .A(n750), .Z(n458) );
  CIVX2 U779 ( .A(n751), .Z(n459) );
  CIVX2 U780 ( .A(n752), .Z(n460) );
  CIVX2 U781 ( .A(n753), .Z(n461) );
  CIVX2 U782 ( .A(n762), .Z(n462) );
  CIVX2 U783 ( .A(n763), .Z(n463) );
  CIVX2 U784 ( .A(n719), .Z(n464) );
  CIVX2 U785 ( .A(n764), .Z(n465) );
  CIVX2 U786 ( .A(n765), .Z(n466) );
  CIVX2 U787 ( .A(n766), .Z(n467) );
  CIVX2 U788 ( .A(n767), .Z(n468) );
  CIVX2 U789 ( .A(n768), .Z(n469) );
  CIVX2 U790 ( .A(n769), .Z(n470) );
  CIVX2 U791 ( .A(n770), .Z(n471) );
  CIVX2 U792 ( .A(n771), .Z(n472) );
  CIVX2 U793 ( .A(n780), .Z(n473) );
  CIVX2 U794 ( .A(n781), .Z(n474) );
  CIVX2 U795 ( .A(n720), .Z(n475) );
  CIVX2 U796 ( .A(n782), .Z(n476) );
  CIVX2 U797 ( .A(n783), .Z(n477) );
  CIVX2 U798 ( .A(n740), .Z(n478) );
  CIVX2 U799 ( .A(n760), .Z(n479) );
  CIVX2 U800 ( .A(n778), .Z(n480) );
  CIVX2 U801 ( .A(n791), .Z(n481) );
  CIVX2 U802 ( .A(n799), .Z(n482) );
  CIVX2 U803 ( .A(n805), .Z(n483) );
  CIVX2 U804 ( .A(n811), .Z(n484) );
  CMX2X1 U805 ( .A0(acc[2]), .A1(acc[1]), .S(n485), .Z(n698) );
  CMXI2X1 U806 ( .A0(n486), .A1(n698), .S(n399), .Z(n487) );
  CMX2X1 U807 ( .A0(acc[4]), .A1(acc[3]), .S(n485), .Z(n697) );
  CMX2X1 U808 ( .A0(acc[6]), .A1(acc[5]), .S(n485), .Z(n700) );
  CMXI2X1 U809 ( .A0(n697), .A1(n700), .S(n399), .Z(n755) );
  CMXI2X1 U810 ( .A0(n487), .A1(n755), .S(n355), .Z(n488) );
  CMX2X1 U811 ( .A0(acc[8]), .A1(acc[7]), .S(n485), .Z(n699) );
  CMX2X1 U812 ( .A0(acc[10]), .A1(acc[9]), .S(n485), .Z(n493) );
  CMXI2X1 U813 ( .A0(n699), .A1(n493), .S(n399), .Z(n754) );
  CMX2X1 U814 ( .A0(acc[12]), .A1(acc[11]), .S(n485), .Z(n492) );
  CMX2X1 U815 ( .A0(acc[14]), .A1(acc[13]), .S(n485), .Z(n495) );
  CMXI2X1 U816 ( .A0(n492), .A1(n495), .S(n398), .Z(n525) );
  CMXI2X1 U817 ( .A0(n754), .A1(n525), .S(n354), .Z(n802) );
  CMXI2X1 U818 ( .A0(n488), .A1(n802), .S(n405), .Z(n489) );
  CMX2X1 U819 ( .A0(acc[16]), .A1(acc[15]), .S(n485), .Z(n494) );
  CMX2X1 U820 ( .A0(acc[18]), .A1(acc[17]), .S(n485), .Z(n497) );
  CMXI2X1 U821 ( .A0(n494), .A1(n497), .S(n398), .Z(n524) );
  CMX2X1 U822 ( .A0(acc[20]), .A1(acc[19]), .S(n485), .Z(n496) );
  CMX2X1 U823 ( .A0(acc[22]), .A1(acc[21]), .S(n485), .Z(n499) );
  CMXI2X1 U824 ( .A0(n496), .A1(n499), .S(n398), .Z(n527) );
  CMXI2X1 U825 ( .A0(n524), .A1(n527), .S(n355), .Z(n801) );
  CMX2X1 U826 ( .A0(acc[24]), .A1(acc[23]), .S(n485), .Z(n498) );
  CMX2X1 U827 ( .A0(acc[26]), .A1(acc[25]), .S(n485), .Z(n501) );
  CMXI2X1 U828 ( .A0(n498), .A1(n501), .S(n398), .Z(n526) );
  CMX2X1 U829 ( .A0(acc[28]), .A1(acc[27]), .S(n485), .Z(n500) );
  CMX2X1 U830 ( .A0(acc[30]), .A1(acc[29]), .S(n485), .Z(n503) );
  CMXI2X1 U831 ( .A0(n500), .A1(n503), .S(n398), .Z(n529) );
  CMXI2X1 U832 ( .A0(n526), .A1(n529), .S(n351), .Z(n669) );
  CMXI2X1 U833 ( .A0(n801), .A1(n669), .S(n405), .Z(n599) );
  CMXI2X1 U834 ( .A0(n489), .A1(n599), .S(n359), .Z(n490) );
  CMX2X1 U835 ( .A0(acc[32]), .A1(acc[31]), .S(n485), .Z(n502) );
  CMX2X1 U836 ( .A0(acc[34]), .A1(acc[33]), .S(n485), .Z(n505) );
  CMXI2X1 U837 ( .A0(n502), .A1(n505), .S(n398), .Z(n528) );
  CMX2X1 U838 ( .A0(acc[36]), .A1(acc[35]), .S(n485), .Z(n504) );
  CMX2X1 U839 ( .A0(acc[38]), .A1(acc[37]), .S(n485), .Z(n507) );
  CMXI2X1 U840 ( .A0(n504), .A1(n507), .S(n398), .Z(n531) );
  CMXI2X1 U841 ( .A0(n528), .A1(n531), .S(n352), .Z(n668) );
  CMX2X1 U842 ( .A0(acc[40]), .A1(acc[39]), .S(n485), .Z(n506) );
  CMX2X1 U843 ( .A0(acc[42]), .A1(acc[41]), .S(n485), .Z(n510) );
  CMXI2X1 U844 ( .A0(n506), .A1(n510), .S(n398), .Z(n530) );
  CMX2X1 U845 ( .A0(acc[44]), .A1(acc[43]), .S(n485), .Z(n509) );
  CMX2X1 U846 ( .A0(acc[46]), .A1(acc[45]), .S(n485), .Z(n512) );
  CMXI2X1 U847 ( .A0(n509), .A1(n512), .S(n398), .Z(n534) );
  CMXI2X1 U848 ( .A0(n530), .A1(n534), .S(n351), .Z(n671) );
  CMXI2X1 U849 ( .A0(n668), .A1(n671), .S(n405), .Z(n598) );
  CMX2X1 U850 ( .A0(acc[48]), .A1(acc[47]), .S(n485), .Z(n511) );
  CMX2X1 U851 ( .A0(acc[50]), .A1(acc[49]), .S(n485), .Z(n514) );
  CMXI2X1 U852 ( .A0(n511), .A1(n514), .S(n398), .Z(n533) );
  CMX2X1 U853 ( .A0(acc[52]), .A1(acc[51]), .S(n485), .Z(n513) );
  CMX2X1 U854 ( .A0(acc[54]), .A1(acc[53]), .S(n485), .Z(n516) );
  CMXI2X1 U855 ( .A0(n513), .A1(n516), .S(n398), .Z(n536) );
  CMXI2X1 U856 ( .A0(n533), .A1(n536), .S(n352), .Z(n670) );
  CMX2X1 U857 ( .A0(acc[56]), .A1(acc[55]), .S(n485), .Z(n515) );
  CMX2X1 U858 ( .A0(acc[58]), .A1(acc[57]), .S(n485), .Z(n518) );
  CMXI2X1 U859 ( .A0(n515), .A1(n518), .S(n398), .Z(n535) );
  CMX2X1 U860 ( .A0(acc[60]), .A1(acc[59]), .S(n485), .Z(n517) );
  CMX2X1 U861 ( .A0(acc[62]), .A1(acc[61]), .S(n485), .Z(n520) );
  CMXI2X1 U862 ( .A0(n517), .A1(n520), .S(n397), .Z(n538) );
  CMXI2X1 U863 ( .A0(n535), .A1(n538), .S(n353), .Z(n673) );
  CMXI2X1 U864 ( .A0(n670), .A1(n673), .S(n405), .Z(n601) );
  CMXI2X1 U865 ( .A0(n598), .A1(n601), .S(n357), .Z(n718) );
  CMXI2X1 U866 ( .A0(n490), .A1(n718), .S(n410), .Z(n491) );
  CND2IX1 U867 ( .B(n410), .A(n717), .Z(n784) );
  CMXI2X1 U868 ( .A0(n491), .A1(n784), .S(n413), .Z(N208) );
  CMXI2X1 U869 ( .A0(n493), .A1(n492), .S(n397), .Z(n785) );
  CMXI2X1 U870 ( .A0(n495), .A1(n494), .S(n397), .Z(n569) );
  CMXI2X1 U871 ( .A0(n785), .A1(n569), .S(n354), .Z(n702) );
  CMXI2X1 U872 ( .A0(n497), .A1(n496), .S(n397), .Z(n568) );
  CMXI2X1 U873 ( .A0(n499), .A1(n498), .S(n397), .Z(n571) );
  CMXI2X1 U874 ( .A0(n568), .A1(n571), .S(n353), .Z(n617) );
  CMXI2X1 U875 ( .A0(n702), .A1(n617), .S(n405), .Z(n508) );
  CMXI2X1 U876 ( .A0(n501), .A1(n500), .S(n397), .Z(n570) );
  CMXI2X1 U877 ( .A0(n503), .A1(n502), .S(n397), .Z(n573) );
  CMXI2X1 U878 ( .A0(n570), .A1(n573), .S(n352), .Z(n616) );
  CMXI2X1 U879 ( .A0(n505), .A1(n504), .S(n397), .Z(n572) );
  CMXI2X1 U880 ( .A0(n507), .A1(n506), .S(n397), .Z(n575) );
  CMXI2X1 U881 ( .A0(n572), .A1(n575), .S(n355), .Z(n619) );
  CMXI2X1 U882 ( .A0(n616), .A1(n619), .S(n405), .Z(n682) );
  CMXI2X1 U883 ( .A0(n508), .A1(n682), .S(n358), .Z(n521) );
  CMXI2X1 U884 ( .A0(n510), .A1(n509), .S(n397), .Z(n574) );
  CMXI2X1 U885 ( .A0(n512), .A1(n511), .S(n397), .Z(n578) );
  CMXI2X1 U886 ( .A0(n574), .A1(n578), .S(n351), .Z(n618) );
  CMXI2X1 U887 ( .A0(n514), .A1(n513), .S(n397), .Z(n577) );
  CMXI2X1 U888 ( .A0(n516), .A1(n515), .S(n396), .Z(n580) );
  CMXI2X1 U889 ( .A0(n577), .A1(n580), .S(n352), .Z(n621) );
  CMXI2X1 U890 ( .A0(n618), .A1(n621), .S(n405), .Z(n681) );
  CMXI2X1 U891 ( .A0(n518), .A1(n517), .S(n396), .Z(n579) );
  CMXI2X1 U892 ( .A0(n520), .A1(n519), .S(n396), .Z(n581) );
  CMXI2X1 U893 ( .A0(n579), .A1(n581), .S(n354), .Z(n620) );
  CMXI2X1 U894 ( .A0(n681), .A1(n683), .S(n359), .Z(n746) );
  CMX2GX1 U895 ( .GN(n413), .A0(n521), .A1(n746), .S(n410), .Z(N218) );
  CMX2X1 U896 ( .A0(acc[11]), .A1(acc[10]), .S(n485), .Z(n632) );
  CMX2X1 U897 ( .A0(acc[13]), .A1(acc[12]), .S(n485), .Z(n541) );
  CMXI2X1 U898 ( .A0(n632), .A1(n541), .S(n396), .Z(n793) );
  CMX2X1 U899 ( .A0(acc[15]), .A1(acc[14]), .S(n485), .Z(n540) );
  CMX2X1 U900 ( .A0(acc[17]), .A1(acc[16]), .S(n485), .Z(n543) );
  CMXI2X1 U901 ( .A0(n540), .A1(n543), .S(n396), .Z(n584) );
  CMXI2X1 U902 ( .A0(n793), .A1(n584), .S(n353), .Z(n736) );
  CMX2X1 U903 ( .A0(acc[19]), .A1(acc[18]), .S(n485), .Z(n542) );
  CMX2X1 U904 ( .A0(acc[21]), .A1(acc[20]), .S(n485), .Z(n545) );
  CMXI2X1 U905 ( .A0(n542), .A1(n545), .S(n396), .Z(n583) );
  CMX2X1 U906 ( .A0(acc[23]), .A1(acc[22]), .S(n485), .Z(n544) );
  CMX2X1 U907 ( .A0(acc[25]), .A1(acc[24]), .S(n485), .Z(n547) );
  CMXI2X1 U908 ( .A0(n544), .A1(n547), .S(n396), .Z(n586) );
  CMXI2X1 U909 ( .A0(n583), .A1(n586), .S(n353), .Z(n624) );
  CMXI2X1 U910 ( .A0(n736), .A1(n624), .S(n405), .Z(n522) );
  CMX2X1 U911 ( .A0(acc[27]), .A1(acc[26]), .S(n485), .Z(n546) );
  CMX2X1 U912 ( .A0(acc[29]), .A1(acc[28]), .S(n485), .Z(n549) );
  CMXI2X1 U913 ( .A0(n546), .A1(n549), .S(n396), .Z(n585) );
  CMX2X1 U914 ( .A0(acc[31]), .A1(acc[30]), .S(n485), .Z(n548) );
  CMX2X1 U915 ( .A0(acc[33]), .A1(acc[32]), .S(n485), .Z(n551) );
  CMXI2X1 U916 ( .A0(n548), .A1(n551), .S(n396), .Z(n588) );
  CMXI2X1 U917 ( .A0(n585), .A1(n588), .S(n354), .Z(n623) );
  CMX2X1 U918 ( .A0(acc[35]), .A1(acc[34]), .S(n485), .Z(n550) );
  CMX2X1 U919 ( .A0(acc[37]), .A1(acc[36]), .S(n485), .Z(n553) );
  CMXI2X1 U920 ( .A0(n550), .A1(n553), .S(n396), .Z(n587) );
  CMX2X1 U921 ( .A0(acc[39]), .A1(acc[38]), .S(n485), .Z(n552) );
  CMX2X1 U922 ( .A0(acc[41]), .A1(acc[40]), .S(n485), .Z(n555) );
  CMXI2X1 U923 ( .A0(n552), .A1(n555), .S(n396), .Z(n590) );
  CMXI2X1 U924 ( .A0(n587), .A1(n590), .S(n355), .Z(n626) );
  CMXI2X1 U925 ( .A0(n623), .A1(n626), .S(n405), .Z(n686) );
  CMXI2X1 U926 ( .A0(n522), .A1(n686), .S(n360), .Z(n523) );
  CMX2X1 U927 ( .A0(acc[43]), .A1(acc[42]), .S(n485), .Z(n554) );
  CMX2X1 U928 ( .A0(acc[45]), .A1(acc[44]), .S(n485), .Z(n558) );
  CMXI2X1 U929 ( .A0(n554), .A1(n558), .S(n395), .Z(n589) );
  CMX2X1 U930 ( .A0(acc[47]), .A1(acc[46]), .S(n485), .Z(n557) );
  CMX2X1 U931 ( .A0(acc[49]), .A1(acc[48]), .S(n485), .Z(n560) );
  CMXI2X1 U932 ( .A0(n557), .A1(n560), .S(n395), .Z(n593) );
  CMXI2X1 U933 ( .A0(n589), .A1(n593), .S(n355), .Z(n625) );
  CMX2X1 U934 ( .A0(acc[51]), .A1(acc[50]), .S(n485), .Z(n559) );
  CMX2X1 U935 ( .A0(acc[53]), .A1(acc[52]), .S(n485), .Z(n562) );
  CMXI2X1 U936 ( .A0(n559), .A1(n562), .S(n395), .Z(n592) );
  CMX2X1 U937 ( .A0(acc[55]), .A1(acc[54]), .S(n485), .Z(n561) );
  CMX2X1 U938 ( .A0(acc[57]), .A1(acc[56]), .S(n485), .Z(n564) );
  CMXI2X1 U939 ( .A0(n561), .A1(n564), .S(n395), .Z(n595) );
  CMXI2X1 U940 ( .A0(n592), .A1(n595), .S(n354), .Z(n628) );
  CMXI2X1 U941 ( .A0(n625), .A1(n628), .S(n404), .Z(n685) );
  CMX2X1 U942 ( .A0(acc[59]), .A1(acc[58]), .S(n485), .Z(n563) );
  CMX2X1 U943 ( .A0(acc[61]), .A1(acc[60]), .S(n485), .Z(n566) );
  CMXI2X1 U944 ( .A0(n563), .A1(n566), .S(n395), .Z(n594) );
  CMX2X1 U945 ( .A0(acc[63]), .A1(acc[62]), .S(n485), .Z(n565) );
  CMXI2X1 U946 ( .A0(n594), .A1(n596), .S(n351), .Z(n627) );
  CMXI2X1 U947 ( .A0(n685), .A1(n687), .S(n358), .Z(n747) );
  CMX2GX1 U948 ( .GN(n413), .A0(n523), .A1(n747), .S(n410), .Z(N219) );
  CMXI2X1 U949 ( .A0(n525), .A1(n524), .S(n352), .Z(n756) );
  CMXI2X1 U950 ( .A0(n527), .A1(n526), .S(n353), .Z(n641) );
  CMXI2X1 U951 ( .A0(n756), .A1(n641), .S(n404), .Z(n532) );
  CMXI2X1 U952 ( .A0(n529), .A1(n528), .S(n351), .Z(n640) );
  CMXI2X1 U953 ( .A0(n531), .A1(n530), .S(n355), .Z(n643) );
  CMXI2X1 U954 ( .A0(n640), .A1(n643), .S(n404), .Z(n690) );
  CMXI2X1 U955 ( .A0(n532), .A1(n690), .S(n360), .Z(n539) );
  CMXI2X1 U956 ( .A0(n534), .A1(n533), .S(n354), .Z(n642) );
  CMXI2X1 U957 ( .A0(n536), .A1(n535), .S(n355), .Z(n645) );
  CMXI2X1 U958 ( .A0(n642), .A1(n645), .S(n404), .Z(n689) );
  CMXI2X1 U959 ( .A0(n538), .A1(n537), .S(n351), .Z(n644) );
  CMXI2X1 U960 ( .A0(n689), .A1(n691), .S(n361), .Z(n748) );
  CMX2GX1 U961 ( .GN(n413), .A0(n539), .A1(n748), .S(n410), .Z(N220) );
  CMXI2X1 U962 ( .A0(n541), .A1(n540), .S(n395), .Z(n633) );
  CMXI2X1 U963 ( .A0(n543), .A1(n542), .S(n395), .Z(n604) );
  CMXI2X1 U964 ( .A0(n633), .A1(n604), .S(n352), .Z(n774) );
  CMXI2X1 U965 ( .A0(n545), .A1(n544), .S(n395), .Z(n603) );
  CMXI2X1 U966 ( .A0(n547), .A1(n546), .S(n395), .Z(n606) );
  CMXI2X1 U967 ( .A0(n603), .A1(n606), .S(n351), .Z(n648) );
  CMXI2X1 U968 ( .A0(n774), .A1(n648), .S(n404), .Z(n556) );
  CMXI2X1 U969 ( .A0(n549), .A1(n548), .S(n396), .Z(n605) );
  CMXI2X1 U970 ( .A0(n551), .A1(n550), .S(n395), .Z(n608) );
  CMXI2X1 U971 ( .A0(n605), .A1(n608), .S(n352), .Z(n647) );
  CMXI2X1 U972 ( .A0(n553), .A1(n552), .S(n395), .Z(n607) );
  CMXI2X1 U973 ( .A0(n555), .A1(n554), .S(n395), .Z(n610) );
  CMXI2X1 U974 ( .A0(n607), .A1(n610), .S(n353), .Z(n650) );
  CMXI2X1 U975 ( .A0(n647), .A1(n650), .S(n404), .Z(n694) );
  CMXI2X1 U976 ( .A0(n556), .A1(n694), .S(n356), .Z(n567) );
  CMXI2X1 U977 ( .A0(n558), .A1(n557), .S(n394), .Z(n609) );
  CMXI2X1 U978 ( .A0(n560), .A1(n559), .S(n394), .Z(n612) );
  CMXI2X1 U979 ( .A0(n609), .A1(n612), .S(n354), .Z(n649) );
  CMXI2X1 U980 ( .A0(n562), .A1(n561), .S(n394), .Z(n611) );
  CMXI2X1 U981 ( .A0(n564), .A1(n563), .S(n394), .Z(n614) );
  CMXI2X1 U982 ( .A0(n611), .A1(n614), .S(n353), .Z(n652) );
  CMXI2X1 U983 ( .A0(n649), .A1(n652), .S(n404), .Z(n693) );
  CMXI2X1 U984 ( .A0(n566), .A1(n565), .S(n394), .Z(n613) );
  CMXI2X1 U985 ( .A0(n693), .A1(n695), .S(n357), .Z(n749) );
  CMX2GX1 U986 ( .GN(n413), .A0(n567), .A1(n749), .S(n410), .Z(N221) );
  CMXI2X1 U987 ( .A0(n569), .A1(n568), .S(n352), .Z(n787) );
  CMXI2X1 U988 ( .A0(n571), .A1(n570), .S(n355), .Z(n655) );
  CMXI2X1 U989 ( .A0(n787), .A1(n655), .S(n404), .Z(n576) );
  CMXI2X1 U990 ( .A0(n573), .A1(n572), .S(n351), .Z(n654) );
  CMXI2X1 U991 ( .A0(n575), .A1(n574), .S(n352), .Z(n657) );
  CMXI2X1 U992 ( .A0(n654), .A1(n657), .S(n404), .Z(n710) );
  CMXI2X1 U993 ( .A0(n576), .A1(n710), .S(n358), .Z(n582) );
  CMXI2X1 U994 ( .A0(n578), .A1(n577), .S(n354), .Z(n656) );
  CMXI2X1 U995 ( .A0(n580), .A1(n579), .S(n353), .Z(n659) );
  CMXI2X1 U996 ( .A0(n656), .A1(n659), .S(n404), .Z(n709) );
  CMXI2X1 U997 ( .A0(n709), .A1(n711), .S(n359), .Z(n750) );
  CMX2GX1 U998 ( .GN(n413), .A0(n582), .A1(n750), .S(n410), .Z(N222) );
  CMXI2X1 U999 ( .A0(n584), .A1(n583), .S(n353), .Z(n795) );
  CMXI2X1 U1000 ( .A0(n586), .A1(n585), .S(n354), .Z(n662) );
  CMXI2X1 U1001 ( .A0(n795), .A1(n662), .S(n404), .Z(n591) );
  CMXI2X1 U1002 ( .A0(n588), .A1(n587), .S(n355), .Z(n661) );
  CMXI2X1 U1003 ( .A0(n590), .A1(n589), .S(n355), .Z(n664) );
  CMXI2X1 U1004 ( .A0(n661), .A1(n664), .S(n404), .Z(n714) );
  CMXI2X1 U1005 ( .A0(n591), .A1(n714), .S(n361), .Z(n597) );
  CMXI2X1 U1006 ( .A0(n593), .A1(n592), .S(n354), .Z(n663) );
  CMXI2X1 U1007 ( .A0(n595), .A1(n594), .S(n351), .Z(n666) );
  CMXI2X1 U1008 ( .A0(n663), .A1(n666), .S(n403), .Z(n713) );
  CMXI2X1 U1009 ( .A0(n713), .A1(n715), .S(n359), .Z(n751) );
  CMX2GX1 U1010 ( .GN(n413), .A0(n597), .A1(n751), .S(n410), .Z(N223) );
  CMXI2X1 U1011 ( .A0(n599), .A1(n598), .S(n360), .Z(n602) );
  CMXI2X1 U1012 ( .A0(n601), .A1(n600), .S(n361), .Z(n752) );
  CMX2GX1 U1013 ( .GN(n413), .A0(n602), .A1(n752), .S(n410), .Z(N224) );
  CMXI2X1 U1014 ( .A0(n604), .A1(n603), .S(n352), .Z(n807) );
  CMXI2X1 U1015 ( .A0(n606), .A1(n605), .S(n353), .Z(n676) );
  CMXI2X1 U1016 ( .A0(n807), .A1(n676), .S(n403), .Z(n635) );
  CMXI2X1 U1017 ( .A0(n608), .A1(n607), .S(n351), .Z(n675) );
  CMXI2X1 U1018 ( .A0(n610), .A1(n609), .S(n355), .Z(n678) );
  CMXI2X1 U1019 ( .A0(n675), .A1(n678), .S(n403), .Z(n638) );
  CMXI2X1 U1020 ( .A0(n635), .A1(n638), .S(n356), .Z(n615) );
  CMXI2X1 U1021 ( .A0(n612), .A1(n611), .S(n354), .Z(n677) );
  CMXI2X1 U1022 ( .A0(n614), .A1(n613), .S(n355), .Z(n679) );
  CMXI2X1 U1023 ( .A0(n677), .A1(n679), .S(n403), .Z(n637) );
  CMX2GX1 U1024 ( .GN(n413), .A0(n615), .A1(n753), .S(n410), .Z(N225) );
  CMXI2X1 U1025 ( .A0(n617), .A1(n616), .S(n403), .Z(n704) );
  CMXI2X1 U1026 ( .A0(n619), .A1(n618), .S(n403), .Z(n707) );
  CMXI2X1 U1027 ( .A0(n704), .A1(n707), .S(n360), .Z(n622) );
  CMXI2X1 U1028 ( .A0(n621), .A1(n620), .S(n403), .Z(n706) );
  CMX2GX1 U1029 ( .GN(n413), .A0(n622), .A1(n762), .S(n410), .Z(N226) );
  CMXI2X1 U1030 ( .A0(n624), .A1(n623), .S(n403), .Z(n738) );
  CMXI2X1 U1031 ( .A0(n626), .A1(n625), .S(n403), .Z(n722) );
  CMXI2X1 U1032 ( .A0(n738), .A1(n722), .S(n356), .Z(n629) );
  CMXI2X1 U1033 ( .A0(n628), .A1(n627), .S(n403), .Z(n721) );
  CMX2GX1 U1034 ( .GN(n413), .A0(n629), .A1(n763), .S(n410), .Z(N227) );
  CMX2X1 U1035 ( .A0(acc[1]), .A1(acc[0]), .S(n485), .Z(n630) );
  CMX2X1 U1036 ( .A0(acc[3]), .A1(acc[2]), .S(n485), .Z(n732) );
  CMXI2X1 U1037 ( .A0(n630), .A1(n732), .S(n394), .Z(n631) );
  CMX2X1 U1038 ( .A0(acc[5]), .A1(acc[4]), .S(n485), .Z(n731) );
  CMX2X1 U1039 ( .A0(acc[7]), .A1(acc[6]), .S(n485), .Z(n734) );
  CMXI2X1 U1040 ( .A0(n731), .A1(n734), .S(n394), .Z(n773) );
  CMXI2X1 U1041 ( .A0(n631), .A1(n773), .S(n351), .Z(n634) );
  CMX2X1 U1042 ( .A0(acc[9]), .A1(acc[8]), .S(n485), .Z(n733) );
  CMXI2X1 U1043 ( .A0(n733), .A1(n632), .S(n394), .Z(n772) );
  CMXI2X1 U1044 ( .A0(n772), .A1(n633), .S(n352), .Z(n808) );
  CMXI2X1 U1045 ( .A0(n634), .A1(n808), .S(n403), .Z(n636) );
  CMXI2X1 U1046 ( .A0(n636), .A1(n635), .S(n357), .Z(n639) );
  CMXI2X1 U1047 ( .A0(n638), .A1(n637), .S(n358), .Z(n719) );
  CMX2GX1 U1048 ( .GN(n413), .A0(n639), .A1(n719), .S(n410), .Z(N209) );
  CMXI2X1 U1049 ( .A0(n641), .A1(n640), .S(n402), .Z(n758) );
  CMXI2X1 U1050 ( .A0(n643), .A1(n642), .S(n402), .Z(n724) );
  CMXI2X1 U1051 ( .A0(n758), .A1(n724), .S(n359), .Z(n646) );
  CMXI2X1 U1052 ( .A0(n645), .A1(n644), .S(n402), .Z(n723) );
  CMX2GX1 U1053 ( .GN(n413), .A0(n646), .A1(n764), .S(n410), .Z(N228) );
  CMXI2X1 U1054 ( .A0(n648), .A1(n647), .S(n402), .Z(n776) );
  CMXI2X1 U1055 ( .A0(n650), .A1(n649), .S(n402), .Z(n726) );
  CMXI2X1 U1056 ( .A0(n776), .A1(n726), .S(n360), .Z(n653) );
  CMXI2X1 U1057 ( .A0(n652), .A1(n651), .S(n402), .Z(n725) );
  CMX2GX1 U1058 ( .GN(n413), .A0(n653), .A1(n765), .S(n410), .Z(N229) );
  CMXI2X1 U1059 ( .A0(n655), .A1(n654), .S(n402), .Z(n789) );
  CMXI2X1 U1060 ( .A0(n657), .A1(n656), .S(n402), .Z(n728) );
  CMXI2X1 U1061 ( .A0(n789), .A1(n728), .S(n361), .Z(n660) );
  CMXI2X1 U1062 ( .A0(n659), .A1(n658), .S(n402), .Z(n727) );
  CMX2GX1 U1063 ( .GN(n413), .A0(n660), .A1(n766), .S(n410), .Z(N230) );
  CMXI2X1 U1064 ( .A0(n662), .A1(n661), .S(n402), .Z(n797) );
  CMXI2X1 U1065 ( .A0(n664), .A1(n663), .S(n402), .Z(n730) );
  CMXI2X1 U1066 ( .A0(n797), .A1(n730), .S(n357), .Z(n667) );
  CMXI2X1 U1067 ( .A0(n666), .A1(n665), .S(n403), .Z(n729) );
  CMX2GX1 U1068 ( .GN(n413), .A0(n667), .A1(n767), .S(n410), .Z(N231) );
  CMXI2X1 U1069 ( .A0(n669), .A1(n668), .S(n402), .Z(n803) );
  CMXI2X1 U1070 ( .A0(n671), .A1(n670), .S(n401), .Z(n743) );
  CMXI2X1 U1071 ( .A0(n803), .A1(n743), .S(n361), .Z(n674) );
  CMXI2X1 U1072 ( .A0(n673), .A1(n672), .S(n401), .Z(n742) );
  CMX2GX1 U1073 ( .GN(n413), .A0(n674), .A1(n768), .S(n410), .Z(N232) );
  CMXI2X1 U1074 ( .A0(n676), .A1(n675), .S(n401), .Z(n809) );
  CMXI2X1 U1075 ( .A0(n678), .A1(n677), .S(n401), .Z(n745) );
  CMXI2X1 U1076 ( .A0(n809), .A1(n745), .S(n356), .Z(n680) );
  CMX2GX1 U1077 ( .GN(n413), .A0(n680), .A1(n769), .S(n410), .Z(N233) );
  CMXI2X1 U1078 ( .A0(n682), .A1(n681), .S(n357), .Z(n684) );
  CMX2GX1 U1079 ( .GN(n413), .A0(n684), .A1(n770), .S(n409), .Z(N234) );
  CMXI2X1 U1080 ( .A0(n686), .A1(n685), .S(n358), .Z(n688) );
  CMX2GX1 U1081 ( .GN(n414), .A0(n688), .A1(n771), .S(n409), .Z(N235) );
  CMXI2X1 U1082 ( .A0(n690), .A1(n689), .S(n356), .Z(n692) );
  CMX2GX1 U1083 ( .GN(n414), .A0(n692), .A1(n780), .S(n409), .Z(N236) );
  CMXI2X1 U1084 ( .A0(n694), .A1(n693), .S(n358), .Z(n696) );
  CMX2GX1 U1085 ( .GN(n414), .A0(n696), .A1(n781), .S(n409), .Z(N237) );
  CMXI2X1 U1086 ( .A0(n698), .A1(n697), .S(n394), .Z(n701) );
  CMXI2X1 U1087 ( .A0(n700), .A1(n699), .S(n394), .Z(n786) );
  CMXI2X1 U1088 ( .A0(n701), .A1(n786), .S(n351), .Z(n703) );
  CMXI2X1 U1089 ( .A0(n703), .A1(n702), .S(n401), .Z(n705) );
  CMXI2X1 U1090 ( .A0(n705), .A1(n704), .S(n359), .Z(n708) );
  CMXI2X1 U1091 ( .A0(n707), .A1(n706), .S(n360), .Z(n720) );
  CMX2GX1 U1092 ( .GN(n414), .A0(n708), .A1(n720), .S(n409), .Z(N210) );
  CMXI2X1 U1093 ( .A0(n710), .A1(n709), .S(n361), .Z(n712) );
  CMX2GX1 U1094 ( .GN(n414), .A0(n712), .A1(n782), .S(n409), .Z(N238) );
  CMXI2X1 U1095 ( .A0(n714), .A1(n713), .S(n356), .Z(n716) );
  CMX2GX1 U1096 ( .GN(n414), .A0(n716), .A1(n783), .S(n409), .Z(N239) );
  CMX2GX1 U1097 ( .GN(n414), .A0(n718), .A1(n717), .S(n409), .Z(N240) );
  CMXI2X1 U1098 ( .A0(n722), .A1(n721), .S(n357), .Z(n740) );
  CMXI2X1 U1099 ( .A0(n724), .A1(n723), .S(n359), .Z(n760) );
  CMXI2X1 U1100 ( .A0(n726), .A1(n725), .S(n357), .Z(n778) );
  CMXI2X1 U1101 ( .A0(n728), .A1(n727), .S(n358), .Z(n791) );
  CMXI2X1 U1102 ( .A0(n730), .A1(n729), .S(n359), .Z(n799) );
  CMXI2X1 U1103 ( .A0(n732), .A1(n731), .S(n394), .Z(n735) );
  CMXI2X1 U1104 ( .A0(n734), .A1(n733), .S(n394), .Z(n794) );
  CMXI2X1 U1105 ( .A0(n735), .A1(n794), .S(n352), .Z(n737) );
  CMXI2X1 U1106 ( .A0(n737), .A1(n736), .S(n401), .Z(n739) );
  CMXI2X1 U1107 ( .A0(n739), .A1(n738), .S(n360), .Z(n741) );
  CMX2GX1 U1108 ( .GN(n414), .A0(n741), .A1(n740), .S(n409), .Z(N211) );
  CMXI2X1 U1109 ( .A0(n743), .A1(n742), .S(n358), .Z(n805) );
  CMXI2X1 U1110 ( .A0(n745), .A1(n744), .S(n360), .Z(n811) );
  CMXI2X1 U1111 ( .A0(n755), .A1(n754), .S(n353), .Z(n757) );
  CMXI2X1 U1112 ( .A0(n757), .A1(n756), .S(n401), .Z(n759) );
  CMXI2X1 U1113 ( .A0(n759), .A1(n758), .S(n361), .Z(n761) );
  CMX2GX1 U1114 ( .GN(n414), .A0(n761), .A1(n760), .S(n409), .Z(N212) );
  CMXI2X1 U1115 ( .A0(n773), .A1(n772), .S(n354), .Z(n775) );
  CMXI2X1 U1116 ( .A0(n775), .A1(n774), .S(n401), .Z(n777) );
  CMXI2X1 U1117 ( .A0(n777), .A1(n776), .S(n356), .Z(n779) );
  CMX2GX1 U1118 ( .GN(n414), .A0(n779), .A1(n778), .S(n409), .Z(N213) );
  CMXI2X1 U1119 ( .A0(n786), .A1(n785), .S(n353), .Z(n788) );
  CMXI2X1 U1120 ( .A0(n788), .A1(n787), .S(n401), .Z(n790) );
  CMXI2X1 U1121 ( .A0(n790), .A1(n789), .S(n357), .Z(n792) );
  CMX2GX1 U1122 ( .GN(n414), .A0(n792), .A1(n791), .S(n409), .Z(N214) );
  CMXI2X1 U1123 ( .A0(n794), .A1(n793), .S(n352), .Z(n796) );
  CMXI2X1 U1124 ( .A0(n796), .A1(n795), .S(n401), .Z(n798) );
  CMXI2X1 U1125 ( .A0(n798), .A1(n797), .S(n358), .Z(n800) );
  CMX2GX1 U1126 ( .GN(n414), .A0(n800), .A1(n799), .S(n409), .Z(N215) );
  CMXI2X1 U1127 ( .A0(n802), .A1(n801), .S(n401), .Z(n804) );
  CMXI2X1 U1128 ( .A0(n804), .A1(n803), .S(n359), .Z(n806) );
  CMX2GX1 U1129 ( .GN(n414), .A0(n806), .A1(n805), .S(n409), .Z(N216) );
  CMXI2X1 U1130 ( .A0(n808), .A1(n807), .S(n401), .Z(n810) );
  CMXI2X1 U1131 ( .A0(n810), .A1(n809), .S(n361), .Z(n812) );
  CMX2GX1 U1132 ( .GN(n414), .A0(n812), .A1(n811), .S(n409), .Z(N217) );
endmodule

