
module poly5_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   \carry[16] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75;

  AND2X2 U1 ( .A(n17), .B(n35), .Y(n1) );
  AND2X2 U2 ( .A(n18), .B(n37), .Y(n2) );
  AND2X2 U3 ( .A(n19), .B(n39), .Y(n3) );
  AND2X2 U4 ( .A(n20), .B(n41), .Y(n4) );
  AND2X2 U5 ( .A(n21), .B(n43), .Y(n5) );
  AND2X2 U6 ( .A(n22), .B(n45), .Y(n6) );
  AND2X2 U7 ( .A(n23), .B(n47), .Y(n7) );
  AND2X2 U8 ( .A(n24), .B(n49), .Y(n8) );
  AND2X2 U9 ( .A(n25), .B(n51), .Y(n9) );
  AND2X2 U10 ( .A(n26), .B(n53), .Y(n10) );
  AND2X2 U11 ( .A(n27), .B(n55), .Y(n11) );
  AND2X2 U12 ( .A(n28), .B(n57), .Y(n12) );
  AND2X2 U13 ( .A(n29), .B(n59), .Y(n13) );
  AND2X2 U14 ( .A(n30), .B(n61), .Y(n14) );
  AND2X2 U15 ( .A(\carry[16] ), .B(n63), .Y(n15) );
  AND2X2 U16 ( .A(n1), .B(n34), .Y(n16) );
  AND2X2 U17 ( .A(n2), .B(n36), .Y(n17) );
  AND2X2 U18 ( .A(n3), .B(n38), .Y(n18) );
  AND2X2 U19 ( .A(n4), .B(n40), .Y(n19) );
  AND2X2 U20 ( .A(n5), .B(n42), .Y(n20) );
  AND2X2 U21 ( .A(n6), .B(n44), .Y(n21) );
  AND2X2 U22 ( .A(n7), .B(n46), .Y(n22) );
  AND2X2 U23 ( .A(n8), .B(n48), .Y(n23) );
  AND2X2 U24 ( .A(n9), .B(n50), .Y(n24) );
  AND2X2 U25 ( .A(n10), .B(n52), .Y(n25) );
  AND2X2 U26 ( .A(n11), .B(n54), .Y(n26) );
  AND2X2 U27 ( .A(n12), .B(n56), .Y(n27) );
  AND2X2 U28 ( .A(n13), .B(n58), .Y(n28) );
  AND2X2 U29 ( .A(n14), .B(n60), .Y(n29) );
  AND2X2 U30 ( .A(n15), .B(n62), .Y(n30) );
  AND2X2 U31 ( .A(n16), .B(n33), .Y(n31) );
  XOR2X1 U32 ( .A(n32), .B(n31), .Y(DIFF[47]) );
  XOR2X1 U33 ( .A(n16), .B(n33), .Y(DIFF[46]) );
  XOR2X1 U34 ( .A(n1), .B(n34), .Y(DIFF[45]) );
  XOR2X1 U35 ( .A(n17), .B(n35), .Y(DIFF[44]) );
  XOR2X1 U36 ( .A(n2), .B(n36), .Y(DIFF[43]) );
  XOR2X1 U37 ( .A(n18), .B(n37), .Y(DIFF[42]) );
  XOR2X1 U38 ( .A(n3), .B(n38), .Y(DIFF[41]) );
  XOR2X1 U39 ( .A(n19), .B(n39), .Y(DIFF[40]) );
  XOR2X1 U40 ( .A(n4), .B(n40), .Y(DIFF[39]) );
  XOR2X1 U41 ( .A(n20), .B(n41), .Y(DIFF[38]) );
  XOR2X1 U42 ( .A(n5), .B(n42), .Y(DIFF[37]) );
  XOR2X1 U43 ( .A(n21), .B(n43), .Y(DIFF[36]) );
  XOR2X1 U44 ( .A(n6), .B(n44), .Y(DIFF[35]) );
  XOR2X1 U45 ( .A(n22), .B(n45), .Y(DIFF[34]) );
  XOR2X1 U46 ( .A(n7), .B(n46), .Y(DIFF[33]) );
  XOR2X1 U47 ( .A(n23), .B(n47), .Y(DIFF[32]) );
  XOR2X1 U48 ( .A(n8), .B(n48), .Y(DIFF[31]) );
  XOR2X1 U49 ( .A(n24), .B(n49), .Y(DIFF[30]) );
  XOR2X1 U50 ( .A(n9), .B(n50), .Y(DIFF[29]) );
  XOR2X1 U51 ( .A(n25), .B(n51), .Y(DIFF[28]) );
  XOR2X1 U52 ( .A(n10), .B(n52), .Y(DIFF[27]) );
  XOR2X1 U53 ( .A(n26), .B(n53), .Y(DIFF[26]) );
  XOR2X1 U54 ( .A(n11), .B(n54), .Y(DIFF[25]) );
  XOR2X1 U55 ( .A(n27), .B(n55), .Y(DIFF[24]) );
  XOR2X1 U56 ( .A(n12), .B(n56), .Y(DIFF[23]) );
  XOR2X1 U57 ( .A(n28), .B(n57), .Y(DIFF[22]) );
  XOR2X1 U58 ( .A(n13), .B(n58), .Y(DIFF[21]) );
  XOR2X1 U59 ( .A(n29), .B(n59), .Y(DIFF[20]) );
  XOR2X1 U60 ( .A(n14), .B(n60), .Y(DIFF[19]) );
  XOR2X1 U61 ( .A(n30), .B(n61), .Y(DIFF[18]) );
  XOR2X1 U62 ( .A(n15), .B(n62), .Y(DIFF[17]) );
  XOR2X1 U63 ( .A(\carry[16] ), .B(n63), .Y(DIFF[16]) );
  INVX2 U64 ( .A(B[47]), .Y(n32) );
  INVX2 U65 ( .A(B[46]), .Y(n33) );
  INVX2 U66 ( .A(B[45]), .Y(n34) );
  INVX2 U67 ( .A(B[44]), .Y(n35) );
  INVX2 U68 ( .A(B[43]), .Y(n36) );
  INVX2 U69 ( .A(B[42]), .Y(n37) );
  INVX2 U70 ( .A(B[41]), .Y(n38) );
  INVX2 U71 ( .A(B[40]), .Y(n39) );
  INVX2 U72 ( .A(B[39]), .Y(n40) );
  INVX2 U73 ( .A(B[38]), .Y(n41) );
  INVX2 U74 ( .A(B[37]), .Y(n42) );
  INVX2 U75 ( .A(B[36]), .Y(n43) );
  INVX2 U76 ( .A(B[35]), .Y(n44) );
  INVX2 U77 ( .A(B[34]), .Y(n45) );
  INVX2 U78 ( .A(B[33]), .Y(n46) );
  INVX2 U79 ( .A(B[32]), .Y(n47) );
  INVX2 U80 ( .A(B[31]), .Y(n48) );
  INVX2 U81 ( .A(B[30]), .Y(n49) );
  INVX2 U82 ( .A(B[29]), .Y(n50) );
  INVX2 U83 ( .A(B[28]), .Y(n51) );
  INVX2 U84 ( .A(B[27]), .Y(n52) );
  INVX2 U85 ( .A(B[26]), .Y(n53) );
  INVX2 U86 ( .A(B[25]), .Y(n54) );
  INVX2 U87 ( .A(B[24]), .Y(n55) );
  INVX2 U88 ( .A(B[23]), .Y(n56) );
  INVX2 U89 ( .A(B[22]), .Y(n57) );
  INVX2 U90 ( .A(B[21]), .Y(n58) );
  INVX2 U91 ( .A(B[20]), .Y(n59) );
  INVX2 U92 ( .A(B[19]), .Y(n60) );
  INVX2 U93 ( .A(B[18]), .Y(n61) );
  INVX2 U94 ( .A(B[17]), .Y(n62) );
  INVX2 U95 ( .A(B[16]), .Y(n63) );
  NOR2X1 U96 ( .A(n64), .B(n65), .Y(\carry[16] ) );
  NAND3X1 U97 ( .A(n66), .B(n67), .C(n68), .Y(n65) );
  AND2X1 U98 ( .A(n69), .B(n70), .Y(n68) );
  NOR2X1 U99 ( .A(B[1]), .B(B[15]), .Y(n70) );
  NOR2X1 U100 ( .A(B[14]), .B(B[13]), .Y(n69) );
  NOR2X1 U101 ( .A(B[12]), .B(B[11]), .Y(n67) );
  NOR2X1 U102 ( .A(B[10]), .B(B[0]), .Y(n66) );
  NAND3X1 U103 ( .A(n71), .B(n72), .C(n73), .Y(n64) );
  AND2X1 U104 ( .A(n74), .B(n75), .Y(n73) );
  NOR2X1 U105 ( .A(B[9]), .B(B[8]), .Y(n75) );
  NOR2X1 U106 ( .A(B[7]), .B(B[6]), .Y(n74) );
  NOR2X1 U107 ( .A(B[5]), .B(B[4]), .Y(n72) );
  NOR2X1 U108 ( .A(B[3]), .B(B[2]), .Y(n71) );
endmodule


module poly5_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND2X2 U1 ( .A(n15), .B(n33), .Y(n1) );
  AND2X2 U2 ( .A(n16), .B(n35), .Y(n2) );
  AND2X2 U3 ( .A(n17), .B(n37), .Y(n3) );
  AND2X2 U4 ( .A(n18), .B(n39), .Y(n4) );
  AND2X2 U5 ( .A(n19), .B(n41), .Y(n5) );
  AND2X2 U6 ( .A(n20), .B(n43), .Y(n6) );
  AND2X2 U7 ( .A(n21), .B(n45), .Y(n7) );
  AND2X2 U8 ( .A(n22), .B(n47), .Y(n8) );
  AND2X2 U9 ( .A(n23), .B(n49), .Y(n9) );
  AND2X2 U10 ( .A(n24), .B(n51), .Y(n10) );
  AND2X2 U11 ( .A(n25), .B(n53), .Y(n11) );
  AND2X2 U12 ( .A(n26), .B(n55), .Y(n12) );
  AND2X2 U13 ( .A(n27), .B(n57), .Y(n13) );
  AND2X2 U14 ( .A(n28), .B(n59), .Y(n14) );
  AND2X2 U15 ( .A(n2), .B(n34), .Y(n15) );
  AND2X2 U16 ( .A(n3), .B(n36), .Y(n16) );
  AND2X2 U17 ( .A(n4), .B(n38), .Y(n17) );
  AND2X2 U18 ( .A(n5), .B(n40), .Y(n18) );
  AND2X2 U19 ( .A(n6), .B(n42), .Y(n19) );
  AND2X2 U20 ( .A(n7), .B(n44), .Y(n20) );
  AND2X2 U21 ( .A(n8), .B(n46), .Y(n21) );
  AND2X2 U22 ( .A(n9), .B(n48), .Y(n22) );
  AND2X2 U23 ( .A(n10), .B(n50), .Y(n23) );
  AND2X2 U24 ( .A(n11), .B(n52), .Y(n24) );
  AND2X2 U25 ( .A(n12), .B(n54), .Y(n25) );
  AND2X2 U26 ( .A(n13), .B(n56), .Y(n26) );
  AND2X2 U27 ( .A(n14), .B(n58), .Y(n27) );
  AND2X2 U28 ( .A(n61), .B(n60), .Y(n28) );
  AND2X2 U29 ( .A(n1), .B(n32), .Y(n29) );
  XOR2X1 U30 ( .A(B[31]), .B(n30), .Y(DIFF[31]) );
  XOR2X1 U31 ( .A(n29), .B(n31), .Y(DIFF[30]) );
  NAND2X1 U32 ( .A(n29), .B(n31), .Y(n30) );
  XOR2X1 U33 ( .A(n1), .B(n32), .Y(DIFF[29]) );
  XOR2X1 U34 ( .A(n15), .B(n33), .Y(DIFF[28]) );
  XOR2X1 U35 ( .A(n2), .B(n34), .Y(DIFF[27]) );
  XOR2X1 U36 ( .A(n16), .B(n35), .Y(DIFF[26]) );
  XOR2X1 U37 ( .A(n3), .B(n36), .Y(DIFF[25]) );
  XOR2X1 U38 ( .A(n17), .B(n37), .Y(DIFF[24]) );
  XOR2X1 U39 ( .A(n4), .B(n38), .Y(DIFF[23]) );
  XOR2X1 U40 ( .A(n18), .B(n39), .Y(DIFF[22]) );
  XOR2X1 U41 ( .A(n5), .B(n40), .Y(DIFF[21]) );
  XOR2X1 U42 ( .A(n19), .B(n41), .Y(DIFF[20]) );
  XOR2X1 U43 ( .A(n6), .B(n42), .Y(DIFF[19]) );
  XOR2X1 U44 ( .A(n20), .B(n43), .Y(DIFF[18]) );
  XOR2X1 U45 ( .A(n7), .B(n44), .Y(DIFF[17]) );
  XOR2X1 U46 ( .A(n21), .B(n45), .Y(DIFF[16]) );
  XOR2X1 U47 ( .A(n8), .B(n46), .Y(DIFF[15]) );
  XOR2X1 U48 ( .A(n22), .B(n47), .Y(DIFF[14]) );
  XOR2X1 U49 ( .A(n9), .B(n48), .Y(DIFF[13]) );
  XOR2X1 U50 ( .A(n23), .B(n49), .Y(DIFF[12]) );
  XOR2X1 U51 ( .A(n10), .B(n50), .Y(DIFF[11]) );
  XOR2X1 U52 ( .A(n24), .B(n51), .Y(DIFF[10]) );
  XOR2X1 U53 ( .A(n11), .B(n52), .Y(DIFF[9]) );
  XOR2X1 U54 ( .A(n25), .B(n53), .Y(DIFF[8]) );
  XOR2X1 U55 ( .A(n12), .B(n54), .Y(DIFF[7]) );
  XOR2X1 U56 ( .A(n26), .B(n55), .Y(DIFF[6]) );
  XOR2X1 U57 ( .A(n13), .B(n56), .Y(DIFF[5]) );
  XOR2X1 U58 ( .A(n27), .B(n57), .Y(DIFF[4]) );
  XOR2X1 U59 ( .A(n14), .B(n58), .Y(DIFF[3]) );
  XOR2X1 U60 ( .A(n28), .B(n59), .Y(DIFF[2]) );
  XOR2X1 U61 ( .A(n61), .B(n60), .Y(DIFF[1]) );
  INVX2 U62 ( .A(B[30]), .Y(n31) );
  INVX2 U63 ( .A(B[29]), .Y(n32) );
  INVX2 U64 ( .A(B[28]), .Y(n33) );
  INVX2 U65 ( .A(B[27]), .Y(n34) );
  INVX2 U66 ( .A(B[26]), .Y(n35) );
  INVX2 U67 ( .A(B[25]), .Y(n36) );
  INVX2 U68 ( .A(B[24]), .Y(n37) );
  INVX2 U69 ( .A(B[23]), .Y(n38) );
  INVX2 U70 ( .A(B[22]), .Y(n39) );
  INVX2 U71 ( .A(B[21]), .Y(n40) );
  INVX2 U72 ( .A(B[20]), .Y(n41) );
  INVX2 U73 ( .A(B[19]), .Y(n42) );
  INVX2 U74 ( .A(B[18]), .Y(n43) );
  INVX2 U75 ( .A(B[17]), .Y(n44) );
  INVX2 U76 ( .A(B[16]), .Y(n45) );
  INVX2 U77 ( .A(B[15]), .Y(n46) );
  INVX2 U78 ( .A(B[14]), .Y(n47) );
  INVX2 U79 ( .A(B[13]), .Y(n48) );
  INVX2 U80 ( .A(B[12]), .Y(n49) );
  INVX2 U81 ( .A(B[11]), .Y(n50) );
  INVX2 U82 ( .A(B[10]), .Y(n51) );
  INVX2 U83 ( .A(B[9]), .Y(n52) );
  INVX2 U84 ( .A(B[8]), .Y(n53) );
  INVX2 U85 ( .A(B[7]), .Y(n54) );
  INVX2 U86 ( .A(B[6]), .Y(n55) );
  INVX2 U87 ( .A(B[5]), .Y(n56) );
  INVX2 U88 ( .A(B[4]), .Y(n57) );
  INVX2 U89 ( .A(B[3]), .Y(n58) );
  INVX2 U90 ( .A(B[2]), .Y(n59) );
  INVX2 U91 ( .A(B[1]), .Y(n60) );
  INVX2 U92 ( .A(\B[0] ), .Y(n61) );
endmodule


module poly5_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   \carry[16] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75;

  AND2X2 U1 ( .A(n17), .B(n35), .Y(n1) );
  AND2X2 U2 ( .A(n18), .B(n37), .Y(n2) );
  AND2X2 U3 ( .A(n19), .B(n39), .Y(n3) );
  AND2X2 U4 ( .A(n20), .B(n41), .Y(n4) );
  AND2X2 U5 ( .A(n21), .B(n43), .Y(n5) );
  AND2X2 U6 ( .A(n22), .B(n45), .Y(n6) );
  AND2X2 U7 ( .A(n23), .B(n47), .Y(n7) );
  AND2X2 U8 ( .A(n24), .B(n49), .Y(n8) );
  AND2X2 U9 ( .A(n25), .B(n51), .Y(n9) );
  AND2X2 U10 ( .A(n26), .B(n53), .Y(n10) );
  AND2X2 U11 ( .A(n27), .B(n55), .Y(n11) );
  AND2X2 U12 ( .A(n28), .B(n57), .Y(n12) );
  AND2X2 U13 ( .A(n29), .B(n59), .Y(n13) );
  AND2X2 U14 ( .A(n30), .B(n61), .Y(n14) );
  AND2X2 U15 ( .A(\carry[16] ), .B(n63), .Y(n15) );
  AND2X2 U16 ( .A(n1), .B(n34), .Y(n16) );
  AND2X2 U17 ( .A(n2), .B(n36), .Y(n17) );
  AND2X2 U18 ( .A(n3), .B(n38), .Y(n18) );
  AND2X2 U19 ( .A(n4), .B(n40), .Y(n19) );
  AND2X2 U20 ( .A(n5), .B(n42), .Y(n20) );
  AND2X2 U21 ( .A(n6), .B(n44), .Y(n21) );
  AND2X2 U22 ( .A(n7), .B(n46), .Y(n22) );
  AND2X2 U23 ( .A(n8), .B(n48), .Y(n23) );
  AND2X2 U24 ( .A(n9), .B(n50), .Y(n24) );
  AND2X2 U25 ( .A(n10), .B(n52), .Y(n25) );
  AND2X2 U26 ( .A(n11), .B(n54), .Y(n26) );
  AND2X2 U27 ( .A(n12), .B(n56), .Y(n27) );
  AND2X2 U28 ( .A(n13), .B(n58), .Y(n28) );
  AND2X2 U29 ( .A(n14), .B(n60), .Y(n29) );
  AND2X2 U30 ( .A(n15), .B(n62), .Y(n30) );
  AND2X2 U31 ( .A(n16), .B(n33), .Y(n31) );
  XOR2X1 U32 ( .A(n32), .B(n31), .Y(DIFF[47]) );
  XOR2X1 U33 ( .A(n16), .B(n33), .Y(DIFF[46]) );
  XOR2X1 U34 ( .A(n1), .B(n34), .Y(DIFF[45]) );
  XOR2X1 U35 ( .A(n17), .B(n35), .Y(DIFF[44]) );
  XOR2X1 U36 ( .A(n2), .B(n36), .Y(DIFF[43]) );
  XOR2X1 U37 ( .A(n18), .B(n37), .Y(DIFF[42]) );
  XOR2X1 U38 ( .A(n3), .B(n38), .Y(DIFF[41]) );
  XOR2X1 U39 ( .A(n19), .B(n39), .Y(DIFF[40]) );
  XOR2X1 U40 ( .A(n4), .B(n40), .Y(DIFF[39]) );
  XOR2X1 U41 ( .A(n20), .B(n41), .Y(DIFF[38]) );
  XOR2X1 U42 ( .A(n5), .B(n42), .Y(DIFF[37]) );
  XOR2X1 U43 ( .A(n21), .B(n43), .Y(DIFF[36]) );
  XOR2X1 U44 ( .A(n6), .B(n44), .Y(DIFF[35]) );
  XOR2X1 U45 ( .A(n22), .B(n45), .Y(DIFF[34]) );
  XOR2X1 U46 ( .A(n7), .B(n46), .Y(DIFF[33]) );
  XOR2X1 U47 ( .A(n23), .B(n47), .Y(DIFF[32]) );
  XOR2X1 U48 ( .A(n8), .B(n48), .Y(DIFF[31]) );
  XOR2X1 U49 ( .A(n24), .B(n49), .Y(DIFF[30]) );
  XOR2X1 U50 ( .A(n9), .B(n50), .Y(DIFF[29]) );
  XOR2X1 U51 ( .A(n25), .B(n51), .Y(DIFF[28]) );
  XOR2X1 U52 ( .A(n10), .B(n52), .Y(DIFF[27]) );
  XOR2X1 U53 ( .A(n26), .B(n53), .Y(DIFF[26]) );
  XOR2X1 U54 ( .A(n11), .B(n54), .Y(DIFF[25]) );
  XOR2X1 U55 ( .A(n27), .B(n55), .Y(DIFF[24]) );
  XOR2X1 U56 ( .A(n12), .B(n56), .Y(DIFF[23]) );
  XOR2X1 U57 ( .A(n28), .B(n57), .Y(DIFF[22]) );
  XOR2X1 U58 ( .A(n13), .B(n58), .Y(DIFF[21]) );
  XOR2X1 U59 ( .A(n29), .B(n59), .Y(DIFF[20]) );
  XOR2X1 U60 ( .A(n14), .B(n60), .Y(DIFF[19]) );
  XOR2X1 U61 ( .A(n30), .B(n61), .Y(DIFF[18]) );
  XOR2X1 U62 ( .A(n15), .B(n62), .Y(DIFF[17]) );
  XOR2X1 U63 ( .A(\carry[16] ), .B(n63), .Y(DIFF[16]) );
  INVX2 U64 ( .A(B[47]), .Y(n32) );
  INVX2 U65 ( .A(B[46]), .Y(n33) );
  INVX2 U66 ( .A(B[45]), .Y(n34) );
  INVX2 U67 ( .A(B[44]), .Y(n35) );
  INVX2 U68 ( .A(B[43]), .Y(n36) );
  INVX2 U69 ( .A(B[42]), .Y(n37) );
  INVX2 U70 ( .A(B[41]), .Y(n38) );
  INVX2 U71 ( .A(B[40]), .Y(n39) );
  INVX2 U72 ( .A(B[39]), .Y(n40) );
  INVX2 U73 ( .A(B[38]), .Y(n41) );
  INVX2 U74 ( .A(B[37]), .Y(n42) );
  INVX2 U75 ( .A(B[36]), .Y(n43) );
  INVX2 U76 ( .A(B[35]), .Y(n44) );
  INVX2 U77 ( .A(B[34]), .Y(n45) );
  INVX2 U78 ( .A(B[33]), .Y(n46) );
  INVX2 U79 ( .A(B[32]), .Y(n47) );
  INVX2 U80 ( .A(B[31]), .Y(n48) );
  INVX2 U81 ( .A(B[30]), .Y(n49) );
  INVX2 U82 ( .A(B[29]), .Y(n50) );
  INVX2 U83 ( .A(B[28]), .Y(n51) );
  INVX2 U84 ( .A(B[27]), .Y(n52) );
  INVX2 U85 ( .A(B[26]), .Y(n53) );
  INVX2 U86 ( .A(B[25]), .Y(n54) );
  INVX2 U87 ( .A(B[24]), .Y(n55) );
  INVX2 U88 ( .A(B[23]), .Y(n56) );
  INVX2 U89 ( .A(B[22]), .Y(n57) );
  INVX2 U90 ( .A(B[21]), .Y(n58) );
  INVX2 U91 ( .A(B[20]), .Y(n59) );
  INVX2 U92 ( .A(B[19]), .Y(n60) );
  INVX2 U93 ( .A(B[18]), .Y(n61) );
  INVX2 U94 ( .A(B[17]), .Y(n62) );
  INVX2 U95 ( .A(B[16]), .Y(n63) );
  NOR2X1 U96 ( .A(n64), .B(n65), .Y(\carry[16] ) );
  NAND3X1 U97 ( .A(n66), .B(n67), .C(n68), .Y(n65) );
  AND2X1 U98 ( .A(n69), .B(n70), .Y(n68) );
  NOR2X1 U99 ( .A(B[1]), .B(B[15]), .Y(n70) );
  NOR2X1 U100 ( .A(B[14]), .B(B[13]), .Y(n69) );
  NOR2X1 U101 ( .A(B[12]), .B(B[11]), .Y(n67) );
  NOR2X1 U102 ( .A(B[10]), .B(B[0]), .Y(n66) );
  NAND3X1 U103 ( .A(n71), .B(n72), .C(n73), .Y(n64) );
  AND2X1 U104 ( .A(n74), .B(n75), .Y(n73) );
  NOR2X1 U105 ( .A(B[9]), .B(B[8]), .Y(n75) );
  NOR2X1 U106 ( .A(B[7]), .B(B[6]), .Y(n74) );
  NOR2X1 U107 ( .A(B[5]), .B(B[4]), .Y(n72) );
  NOR2X1 U108 ( .A(B[3]), .B(B[2]), .Y(n71) );
endmodule


module poly5_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND2X2 U1 ( .A(n15), .B(n33), .Y(n1) );
  AND2X2 U2 ( .A(n16), .B(n35), .Y(n2) );
  AND2X2 U3 ( .A(n17), .B(n37), .Y(n3) );
  AND2X2 U4 ( .A(n18), .B(n39), .Y(n4) );
  AND2X2 U5 ( .A(n19), .B(n41), .Y(n5) );
  AND2X2 U6 ( .A(n20), .B(n43), .Y(n6) );
  AND2X2 U7 ( .A(n21), .B(n45), .Y(n7) );
  AND2X2 U8 ( .A(n22), .B(n47), .Y(n8) );
  AND2X2 U9 ( .A(n23), .B(n49), .Y(n9) );
  AND2X2 U10 ( .A(n24), .B(n51), .Y(n10) );
  AND2X2 U11 ( .A(n25), .B(n53), .Y(n11) );
  AND2X2 U12 ( .A(n26), .B(n55), .Y(n12) );
  AND2X2 U13 ( .A(n27), .B(n57), .Y(n13) );
  AND2X2 U14 ( .A(n28), .B(n59), .Y(n14) );
  AND2X2 U15 ( .A(n2), .B(n34), .Y(n15) );
  AND2X2 U16 ( .A(n3), .B(n36), .Y(n16) );
  AND2X2 U17 ( .A(n4), .B(n38), .Y(n17) );
  AND2X2 U18 ( .A(n5), .B(n40), .Y(n18) );
  AND2X2 U19 ( .A(n6), .B(n42), .Y(n19) );
  AND2X2 U20 ( .A(n7), .B(n44), .Y(n20) );
  AND2X2 U21 ( .A(n8), .B(n46), .Y(n21) );
  AND2X2 U22 ( .A(n9), .B(n48), .Y(n22) );
  AND2X2 U23 ( .A(n10), .B(n50), .Y(n23) );
  AND2X2 U24 ( .A(n11), .B(n52), .Y(n24) );
  AND2X2 U25 ( .A(n12), .B(n54), .Y(n25) );
  AND2X2 U26 ( .A(n13), .B(n56), .Y(n26) );
  AND2X2 U27 ( .A(n14), .B(n58), .Y(n27) );
  AND2X2 U28 ( .A(n61), .B(n60), .Y(n28) );
  AND2X2 U29 ( .A(n1), .B(n32), .Y(n29) );
  XOR2X1 U30 ( .A(B[31]), .B(n30), .Y(DIFF[31]) );
  XOR2X1 U31 ( .A(n29), .B(n31), .Y(DIFF[30]) );
  NAND2X1 U32 ( .A(n29), .B(n31), .Y(n30) );
  XOR2X1 U33 ( .A(n1), .B(n32), .Y(DIFF[29]) );
  XOR2X1 U34 ( .A(n15), .B(n33), .Y(DIFF[28]) );
  XOR2X1 U35 ( .A(n2), .B(n34), .Y(DIFF[27]) );
  XOR2X1 U36 ( .A(n16), .B(n35), .Y(DIFF[26]) );
  XOR2X1 U37 ( .A(n3), .B(n36), .Y(DIFF[25]) );
  XOR2X1 U38 ( .A(n17), .B(n37), .Y(DIFF[24]) );
  XOR2X1 U39 ( .A(n4), .B(n38), .Y(DIFF[23]) );
  XOR2X1 U40 ( .A(n18), .B(n39), .Y(DIFF[22]) );
  XOR2X1 U41 ( .A(n5), .B(n40), .Y(DIFF[21]) );
  XOR2X1 U42 ( .A(n19), .B(n41), .Y(DIFF[20]) );
  XOR2X1 U43 ( .A(n6), .B(n42), .Y(DIFF[19]) );
  XOR2X1 U44 ( .A(n20), .B(n43), .Y(DIFF[18]) );
  XOR2X1 U45 ( .A(n7), .B(n44), .Y(DIFF[17]) );
  XOR2X1 U46 ( .A(n21), .B(n45), .Y(DIFF[16]) );
  XOR2X1 U47 ( .A(n8), .B(n46), .Y(DIFF[15]) );
  XOR2X1 U48 ( .A(n22), .B(n47), .Y(DIFF[14]) );
  XOR2X1 U49 ( .A(n9), .B(n48), .Y(DIFF[13]) );
  XOR2X1 U50 ( .A(n23), .B(n49), .Y(DIFF[12]) );
  XOR2X1 U51 ( .A(n10), .B(n50), .Y(DIFF[11]) );
  XOR2X1 U52 ( .A(n24), .B(n51), .Y(DIFF[10]) );
  XOR2X1 U53 ( .A(n11), .B(n52), .Y(DIFF[9]) );
  XOR2X1 U54 ( .A(n25), .B(n53), .Y(DIFF[8]) );
  XOR2X1 U55 ( .A(n12), .B(n54), .Y(DIFF[7]) );
  XOR2X1 U56 ( .A(n26), .B(n55), .Y(DIFF[6]) );
  XOR2X1 U57 ( .A(n13), .B(n56), .Y(DIFF[5]) );
  XOR2X1 U58 ( .A(n27), .B(n57), .Y(DIFF[4]) );
  XOR2X1 U59 ( .A(n14), .B(n58), .Y(DIFF[3]) );
  XOR2X1 U60 ( .A(n28), .B(n59), .Y(DIFF[2]) );
  XOR2X1 U61 ( .A(n61), .B(n60), .Y(DIFF[1]) );
  INVX2 U62 ( .A(B[30]), .Y(n31) );
  INVX2 U63 ( .A(B[29]), .Y(n32) );
  INVX2 U64 ( .A(B[28]), .Y(n33) );
  INVX2 U65 ( .A(B[27]), .Y(n34) );
  INVX2 U66 ( .A(B[26]), .Y(n35) );
  INVX2 U67 ( .A(B[25]), .Y(n36) );
  INVX2 U68 ( .A(B[24]), .Y(n37) );
  INVX2 U69 ( .A(B[23]), .Y(n38) );
  INVX2 U70 ( .A(B[22]), .Y(n39) );
  INVX2 U71 ( .A(B[21]), .Y(n40) );
  INVX2 U72 ( .A(B[20]), .Y(n41) );
  INVX2 U73 ( .A(B[19]), .Y(n42) );
  INVX2 U74 ( .A(B[18]), .Y(n43) );
  INVX2 U75 ( .A(B[17]), .Y(n44) );
  INVX2 U76 ( .A(B[16]), .Y(n45) );
  INVX2 U77 ( .A(B[15]), .Y(n46) );
  INVX2 U78 ( .A(B[14]), .Y(n47) );
  INVX2 U79 ( .A(B[13]), .Y(n48) );
  INVX2 U80 ( .A(B[12]), .Y(n49) );
  INVX2 U81 ( .A(B[11]), .Y(n50) );
  INVX2 U82 ( .A(B[10]), .Y(n51) );
  INVX2 U83 ( .A(B[9]), .Y(n52) );
  INVX2 U84 ( .A(B[8]), .Y(n53) );
  INVX2 U85 ( .A(B[7]), .Y(n54) );
  INVX2 U86 ( .A(B[6]), .Y(n55) );
  INVX2 U87 ( .A(B[5]), .Y(n56) );
  INVX2 U88 ( .A(B[4]), .Y(n57) );
  INVX2 U89 ( .A(B[3]), .Y(n58) );
  INVX2 U90 ( .A(B[2]), .Y(n59) );
  INVX2 U91 ( .A(B[1]), .Y(n60) );
  INVX2 U92 ( .A(\B[0] ), .Y(n61) );
endmodule


module poly5_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   \carry[16] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75;

  AND2X2 U1 ( .A(n17), .B(n35), .Y(n1) );
  AND2X2 U2 ( .A(n18), .B(n37), .Y(n2) );
  AND2X2 U3 ( .A(n19), .B(n39), .Y(n3) );
  AND2X2 U4 ( .A(n20), .B(n41), .Y(n4) );
  AND2X2 U5 ( .A(n21), .B(n43), .Y(n5) );
  AND2X2 U6 ( .A(n22), .B(n45), .Y(n6) );
  AND2X2 U7 ( .A(n23), .B(n47), .Y(n7) );
  AND2X2 U8 ( .A(n24), .B(n49), .Y(n8) );
  AND2X2 U9 ( .A(n25), .B(n51), .Y(n9) );
  AND2X2 U10 ( .A(n26), .B(n53), .Y(n10) );
  AND2X2 U11 ( .A(n27), .B(n55), .Y(n11) );
  AND2X2 U12 ( .A(n28), .B(n57), .Y(n12) );
  AND2X2 U13 ( .A(n29), .B(n59), .Y(n13) );
  AND2X2 U14 ( .A(n30), .B(n61), .Y(n14) );
  AND2X2 U15 ( .A(\carry[16] ), .B(n63), .Y(n15) );
  AND2X2 U16 ( .A(n1), .B(n34), .Y(n16) );
  AND2X2 U17 ( .A(n2), .B(n36), .Y(n17) );
  AND2X2 U18 ( .A(n3), .B(n38), .Y(n18) );
  AND2X2 U19 ( .A(n4), .B(n40), .Y(n19) );
  AND2X2 U20 ( .A(n5), .B(n42), .Y(n20) );
  AND2X2 U21 ( .A(n6), .B(n44), .Y(n21) );
  AND2X2 U22 ( .A(n7), .B(n46), .Y(n22) );
  AND2X2 U23 ( .A(n8), .B(n48), .Y(n23) );
  AND2X2 U24 ( .A(n9), .B(n50), .Y(n24) );
  AND2X2 U25 ( .A(n10), .B(n52), .Y(n25) );
  AND2X2 U26 ( .A(n11), .B(n54), .Y(n26) );
  AND2X2 U27 ( .A(n12), .B(n56), .Y(n27) );
  AND2X2 U28 ( .A(n13), .B(n58), .Y(n28) );
  AND2X2 U29 ( .A(n14), .B(n60), .Y(n29) );
  AND2X2 U30 ( .A(n15), .B(n62), .Y(n30) );
  AND2X2 U31 ( .A(n16), .B(n33), .Y(n31) );
  XOR2X1 U32 ( .A(n32), .B(n31), .Y(DIFF[47]) );
  XOR2X1 U33 ( .A(n16), .B(n33), .Y(DIFF[46]) );
  XOR2X1 U34 ( .A(n1), .B(n34), .Y(DIFF[45]) );
  XOR2X1 U35 ( .A(n17), .B(n35), .Y(DIFF[44]) );
  XOR2X1 U36 ( .A(n2), .B(n36), .Y(DIFF[43]) );
  XOR2X1 U37 ( .A(n18), .B(n37), .Y(DIFF[42]) );
  XOR2X1 U38 ( .A(n3), .B(n38), .Y(DIFF[41]) );
  XOR2X1 U39 ( .A(n19), .B(n39), .Y(DIFF[40]) );
  XOR2X1 U40 ( .A(n4), .B(n40), .Y(DIFF[39]) );
  XOR2X1 U41 ( .A(n20), .B(n41), .Y(DIFF[38]) );
  XOR2X1 U42 ( .A(n5), .B(n42), .Y(DIFF[37]) );
  XOR2X1 U43 ( .A(n21), .B(n43), .Y(DIFF[36]) );
  XOR2X1 U44 ( .A(n6), .B(n44), .Y(DIFF[35]) );
  XOR2X1 U45 ( .A(n22), .B(n45), .Y(DIFF[34]) );
  XOR2X1 U46 ( .A(n7), .B(n46), .Y(DIFF[33]) );
  XOR2X1 U47 ( .A(n23), .B(n47), .Y(DIFF[32]) );
  XOR2X1 U48 ( .A(n8), .B(n48), .Y(DIFF[31]) );
  XOR2X1 U49 ( .A(n24), .B(n49), .Y(DIFF[30]) );
  XOR2X1 U50 ( .A(n9), .B(n50), .Y(DIFF[29]) );
  XOR2X1 U51 ( .A(n25), .B(n51), .Y(DIFF[28]) );
  XOR2X1 U52 ( .A(n10), .B(n52), .Y(DIFF[27]) );
  XOR2X1 U53 ( .A(n26), .B(n53), .Y(DIFF[26]) );
  XOR2X1 U54 ( .A(n11), .B(n54), .Y(DIFF[25]) );
  XOR2X1 U55 ( .A(n27), .B(n55), .Y(DIFF[24]) );
  XOR2X1 U56 ( .A(n12), .B(n56), .Y(DIFF[23]) );
  XOR2X1 U57 ( .A(n28), .B(n57), .Y(DIFF[22]) );
  XOR2X1 U58 ( .A(n13), .B(n58), .Y(DIFF[21]) );
  XOR2X1 U59 ( .A(n29), .B(n59), .Y(DIFF[20]) );
  XOR2X1 U60 ( .A(n14), .B(n60), .Y(DIFF[19]) );
  XOR2X1 U61 ( .A(n30), .B(n61), .Y(DIFF[18]) );
  XOR2X1 U62 ( .A(n15), .B(n62), .Y(DIFF[17]) );
  XOR2X1 U63 ( .A(\carry[16] ), .B(n63), .Y(DIFF[16]) );
  INVX2 U64 ( .A(B[47]), .Y(n32) );
  INVX2 U65 ( .A(B[46]), .Y(n33) );
  INVX2 U66 ( .A(B[45]), .Y(n34) );
  INVX2 U67 ( .A(B[44]), .Y(n35) );
  INVX2 U68 ( .A(B[43]), .Y(n36) );
  INVX2 U69 ( .A(B[42]), .Y(n37) );
  INVX2 U70 ( .A(B[41]), .Y(n38) );
  INVX2 U71 ( .A(B[40]), .Y(n39) );
  INVX2 U72 ( .A(B[39]), .Y(n40) );
  INVX2 U73 ( .A(B[38]), .Y(n41) );
  INVX2 U74 ( .A(B[37]), .Y(n42) );
  INVX2 U75 ( .A(B[36]), .Y(n43) );
  INVX2 U76 ( .A(B[35]), .Y(n44) );
  INVX2 U77 ( .A(B[34]), .Y(n45) );
  INVX2 U78 ( .A(B[33]), .Y(n46) );
  INVX2 U79 ( .A(B[32]), .Y(n47) );
  INVX2 U80 ( .A(B[31]), .Y(n48) );
  INVX2 U81 ( .A(B[30]), .Y(n49) );
  INVX2 U82 ( .A(B[29]), .Y(n50) );
  INVX2 U83 ( .A(B[28]), .Y(n51) );
  INVX2 U84 ( .A(B[27]), .Y(n52) );
  INVX2 U85 ( .A(B[26]), .Y(n53) );
  INVX2 U86 ( .A(B[25]), .Y(n54) );
  INVX2 U87 ( .A(B[24]), .Y(n55) );
  INVX2 U88 ( .A(B[23]), .Y(n56) );
  INVX2 U89 ( .A(B[22]), .Y(n57) );
  INVX2 U90 ( .A(B[21]), .Y(n58) );
  INVX2 U91 ( .A(B[20]), .Y(n59) );
  INVX2 U92 ( .A(B[19]), .Y(n60) );
  INVX2 U93 ( .A(B[18]), .Y(n61) );
  INVX2 U94 ( .A(B[17]), .Y(n62) );
  INVX2 U95 ( .A(B[16]), .Y(n63) );
  NOR2X1 U96 ( .A(n64), .B(n65), .Y(\carry[16] ) );
  NAND3X1 U97 ( .A(n66), .B(n67), .C(n68), .Y(n65) );
  AND2X1 U98 ( .A(n69), .B(n70), .Y(n68) );
  NOR2X1 U99 ( .A(B[1]), .B(B[15]), .Y(n70) );
  NOR2X1 U100 ( .A(B[14]), .B(B[13]), .Y(n69) );
  NOR2X1 U101 ( .A(B[12]), .B(B[11]), .Y(n67) );
  NOR2X1 U102 ( .A(B[10]), .B(B[0]), .Y(n66) );
  NAND3X1 U103 ( .A(n71), .B(n72), .C(n73), .Y(n64) );
  AND2X1 U104 ( .A(n74), .B(n75), .Y(n73) );
  NOR2X1 U105 ( .A(B[9]), .B(B[8]), .Y(n75) );
  NOR2X1 U106 ( .A(B[7]), .B(B[6]), .Y(n74) );
  NOR2X1 U107 ( .A(B[5]), .B(B[4]), .Y(n72) );
  NOR2X1 U108 ( .A(B[3]), .B(B[2]), .Y(n71) );
endmodule


module poly5_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND2X2 U1 ( .A(n15), .B(n33), .Y(n1) );
  AND2X2 U2 ( .A(n16), .B(n35), .Y(n2) );
  AND2X2 U3 ( .A(n17), .B(n37), .Y(n3) );
  AND2X2 U4 ( .A(n18), .B(n39), .Y(n4) );
  AND2X2 U5 ( .A(n19), .B(n41), .Y(n5) );
  AND2X2 U6 ( .A(n20), .B(n43), .Y(n6) );
  AND2X2 U7 ( .A(n21), .B(n45), .Y(n7) );
  AND2X2 U8 ( .A(n22), .B(n47), .Y(n8) );
  AND2X2 U9 ( .A(n23), .B(n49), .Y(n9) );
  AND2X2 U10 ( .A(n24), .B(n51), .Y(n10) );
  AND2X2 U11 ( .A(n25), .B(n53), .Y(n11) );
  AND2X2 U12 ( .A(n26), .B(n55), .Y(n12) );
  AND2X2 U13 ( .A(n27), .B(n57), .Y(n13) );
  AND2X2 U14 ( .A(n28), .B(n59), .Y(n14) );
  AND2X2 U15 ( .A(n2), .B(n34), .Y(n15) );
  AND2X2 U16 ( .A(n3), .B(n36), .Y(n16) );
  AND2X2 U17 ( .A(n4), .B(n38), .Y(n17) );
  AND2X2 U18 ( .A(n5), .B(n40), .Y(n18) );
  AND2X2 U19 ( .A(n6), .B(n42), .Y(n19) );
  AND2X2 U20 ( .A(n7), .B(n44), .Y(n20) );
  AND2X2 U21 ( .A(n8), .B(n46), .Y(n21) );
  AND2X2 U22 ( .A(n9), .B(n48), .Y(n22) );
  AND2X2 U23 ( .A(n10), .B(n50), .Y(n23) );
  AND2X2 U24 ( .A(n11), .B(n52), .Y(n24) );
  AND2X2 U25 ( .A(n12), .B(n54), .Y(n25) );
  AND2X2 U26 ( .A(n13), .B(n56), .Y(n26) );
  AND2X2 U27 ( .A(n14), .B(n58), .Y(n27) );
  AND2X2 U28 ( .A(n61), .B(n60), .Y(n28) );
  AND2X2 U29 ( .A(n1), .B(n32), .Y(n29) );
  XOR2X1 U30 ( .A(B[31]), .B(n30), .Y(DIFF[31]) );
  XOR2X1 U31 ( .A(n29), .B(n31), .Y(DIFF[30]) );
  NAND2X1 U32 ( .A(n29), .B(n31), .Y(n30) );
  XOR2X1 U33 ( .A(n1), .B(n32), .Y(DIFF[29]) );
  XOR2X1 U34 ( .A(n15), .B(n33), .Y(DIFF[28]) );
  XOR2X1 U35 ( .A(n2), .B(n34), .Y(DIFF[27]) );
  XOR2X1 U36 ( .A(n16), .B(n35), .Y(DIFF[26]) );
  XOR2X1 U37 ( .A(n3), .B(n36), .Y(DIFF[25]) );
  XOR2X1 U38 ( .A(n17), .B(n37), .Y(DIFF[24]) );
  XOR2X1 U39 ( .A(n4), .B(n38), .Y(DIFF[23]) );
  XOR2X1 U40 ( .A(n18), .B(n39), .Y(DIFF[22]) );
  XOR2X1 U41 ( .A(n5), .B(n40), .Y(DIFF[21]) );
  XOR2X1 U42 ( .A(n19), .B(n41), .Y(DIFF[20]) );
  XOR2X1 U43 ( .A(n6), .B(n42), .Y(DIFF[19]) );
  XOR2X1 U44 ( .A(n20), .B(n43), .Y(DIFF[18]) );
  XOR2X1 U45 ( .A(n7), .B(n44), .Y(DIFF[17]) );
  XOR2X1 U46 ( .A(n21), .B(n45), .Y(DIFF[16]) );
  XOR2X1 U47 ( .A(n8), .B(n46), .Y(DIFF[15]) );
  XOR2X1 U48 ( .A(n22), .B(n47), .Y(DIFF[14]) );
  XOR2X1 U49 ( .A(n9), .B(n48), .Y(DIFF[13]) );
  XOR2X1 U50 ( .A(n23), .B(n49), .Y(DIFF[12]) );
  XOR2X1 U51 ( .A(n10), .B(n50), .Y(DIFF[11]) );
  XOR2X1 U52 ( .A(n24), .B(n51), .Y(DIFF[10]) );
  XOR2X1 U53 ( .A(n11), .B(n52), .Y(DIFF[9]) );
  XOR2X1 U54 ( .A(n25), .B(n53), .Y(DIFF[8]) );
  XOR2X1 U55 ( .A(n12), .B(n54), .Y(DIFF[7]) );
  XOR2X1 U56 ( .A(n26), .B(n55), .Y(DIFF[6]) );
  XOR2X1 U57 ( .A(n13), .B(n56), .Y(DIFF[5]) );
  XOR2X1 U58 ( .A(n27), .B(n57), .Y(DIFF[4]) );
  XOR2X1 U59 ( .A(n14), .B(n58), .Y(DIFF[3]) );
  XOR2X1 U60 ( .A(n28), .B(n59), .Y(DIFF[2]) );
  XOR2X1 U61 ( .A(n61), .B(n60), .Y(DIFF[1]) );
  INVX2 U62 ( .A(B[30]), .Y(n31) );
  INVX2 U63 ( .A(B[29]), .Y(n32) );
  INVX2 U64 ( .A(B[28]), .Y(n33) );
  INVX2 U65 ( .A(B[27]), .Y(n34) );
  INVX2 U66 ( .A(B[26]), .Y(n35) );
  INVX2 U67 ( .A(B[25]), .Y(n36) );
  INVX2 U68 ( .A(B[24]), .Y(n37) );
  INVX2 U69 ( .A(B[23]), .Y(n38) );
  INVX2 U70 ( .A(B[22]), .Y(n39) );
  INVX2 U71 ( .A(B[21]), .Y(n40) );
  INVX2 U72 ( .A(B[20]), .Y(n41) );
  INVX2 U73 ( .A(B[19]), .Y(n42) );
  INVX2 U74 ( .A(B[18]), .Y(n43) );
  INVX2 U75 ( .A(B[17]), .Y(n44) );
  INVX2 U76 ( .A(B[16]), .Y(n45) );
  INVX2 U77 ( .A(B[15]), .Y(n46) );
  INVX2 U78 ( .A(B[14]), .Y(n47) );
  INVX2 U79 ( .A(B[13]), .Y(n48) );
  INVX2 U80 ( .A(B[12]), .Y(n49) );
  INVX2 U81 ( .A(B[11]), .Y(n50) );
  INVX2 U82 ( .A(B[10]), .Y(n51) );
  INVX2 U83 ( .A(B[9]), .Y(n52) );
  INVX2 U84 ( .A(B[8]), .Y(n53) );
  INVX2 U85 ( .A(B[7]), .Y(n54) );
  INVX2 U86 ( .A(B[6]), .Y(n55) );
  INVX2 U87 ( .A(B[5]), .Y(n56) );
  INVX2 U88 ( .A(B[4]), .Y(n57) );
  INVX2 U89 ( .A(B[3]), .Y(n58) );
  INVX2 U90 ( .A(B[2]), .Y(n59) );
  INVX2 U91 ( .A(B[1]), .Y(n60) );
  INVX2 U92 ( .A(\B[0] ), .Y(n61) );
endmodule


module poly5_DW01_sub_6 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   \carry[16] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75;

  AND2X2 U1 ( .A(n11), .B(n39), .Y(n1) );
  AND2X2 U2 ( .A(n9), .B(n43), .Y(n2) );
  AND2X2 U3 ( .A(n10), .B(n45), .Y(n3) );
  AND2X2 U4 ( .A(n12), .B(n41), .Y(n4) );
  AND2X2 U5 ( .A(n14), .B(n35), .Y(n5) );
  AND2X2 U6 ( .A(n8), .B(n37), .Y(n6) );
  AND2X2 U7 ( .A(n18), .B(n47), .Y(n7) );
  AND2X2 U8 ( .A(n1), .B(n38), .Y(n8) );
  AND2X2 U9 ( .A(n3), .B(n44), .Y(n9) );
  AND2X2 U10 ( .A(n7), .B(n46), .Y(n10) );
  AND2X2 U11 ( .A(n4), .B(n40), .Y(n11) );
  AND2X2 U12 ( .A(n2), .B(n42), .Y(n12) );
  AND2X2 U13 ( .A(n5), .B(n34), .Y(n13) );
  AND2X2 U14 ( .A(n6), .B(n36), .Y(n14) );
  AND2X2 U15 ( .A(n13), .B(n33), .Y(n15) );
  AND2X1 U16 ( .A(n19), .B(n50), .Y(n16) );
  AND2X2 U17 ( .A(n16), .B(n49), .Y(n17) );
  AND2X2 U18 ( .A(n17), .B(n48), .Y(n18) );
  AND2X1 U19 ( .A(n21), .B(n51), .Y(n19) );
  AND2X2 U20 ( .A(n25), .B(n58), .Y(n24) );
  AND2X2 U21 ( .A(n24), .B(n57), .Y(n26) );
  AND2X2 U22 ( .A(n26), .B(n56), .Y(n27) );
  AND2X2 U23 ( .A(n28), .B(n59), .Y(n25) );
  AND2X2 U24 ( .A(n27), .B(n55), .Y(n23) );
  AND2X2 U25 ( .A(n23), .B(n54), .Y(n20) );
  AND2X1 U26 ( .A(n22), .B(n52), .Y(n21) );
  AND2X2 U27 ( .A(n20), .B(n53), .Y(n22) );
  AND2X2 U28 ( .A(n29), .B(n60), .Y(n28) );
  AND2X2 U29 ( .A(n30), .B(n61), .Y(n29) );
  AND2X2 U30 ( .A(n31), .B(n62), .Y(n30) );
  AND2X2 U31 ( .A(\carry[16] ), .B(n63), .Y(n31) );
  XOR2X1 U32 ( .A(n32), .B(n15), .Y(DIFF[47]) );
  XOR2X1 U33 ( .A(n13), .B(n33), .Y(DIFF[46]) );
  XOR2X1 U34 ( .A(n5), .B(n34), .Y(DIFF[45]) );
  XOR2X1 U35 ( .A(n14), .B(n35), .Y(DIFF[44]) );
  XOR2X1 U36 ( .A(n6), .B(n36), .Y(DIFF[43]) );
  XOR2X1 U37 ( .A(n8), .B(n37), .Y(DIFF[42]) );
  XOR2X1 U38 ( .A(n1), .B(n38), .Y(DIFF[41]) );
  XOR2X1 U39 ( .A(n11), .B(n39), .Y(DIFF[40]) );
  XOR2X1 U40 ( .A(n4), .B(n40), .Y(DIFF[39]) );
  XOR2X1 U41 ( .A(n12), .B(n41), .Y(DIFF[38]) );
  XOR2X1 U42 ( .A(n2), .B(n42), .Y(DIFF[37]) );
  XOR2X1 U43 ( .A(n9), .B(n43), .Y(DIFF[36]) );
  XOR2X1 U44 ( .A(n3), .B(n44), .Y(DIFF[35]) );
  XOR2X1 U45 ( .A(n10), .B(n45), .Y(DIFF[34]) );
  XOR2X1 U46 ( .A(n7), .B(n46), .Y(DIFF[33]) );
  XOR2X1 U47 ( .A(n18), .B(n47), .Y(DIFF[32]) );
  XOR2X1 U48 ( .A(n17), .B(n48), .Y(DIFF[31]) );
  XOR2X1 U49 ( .A(n16), .B(n49), .Y(DIFF[30]) );
  XOR2X1 U50 ( .A(n19), .B(n50), .Y(DIFF[29]) );
  XOR2X1 U51 ( .A(n21), .B(n51), .Y(DIFF[28]) );
  XOR2X1 U52 ( .A(n22), .B(n52), .Y(DIFF[27]) );
  XOR2X1 U53 ( .A(n20), .B(n53), .Y(DIFF[26]) );
  XOR2X1 U54 ( .A(n23), .B(n54), .Y(DIFF[25]) );
  XOR2X1 U55 ( .A(n27), .B(n55), .Y(DIFF[24]) );
  XOR2X1 U56 ( .A(n26), .B(n56), .Y(DIFF[23]) );
  XOR2X1 U57 ( .A(n24), .B(n57), .Y(DIFF[22]) );
  XOR2X1 U58 ( .A(n25), .B(n58), .Y(DIFF[21]) );
  XOR2X1 U59 ( .A(n28), .B(n59), .Y(DIFF[20]) );
  XOR2X1 U60 ( .A(n29), .B(n60), .Y(DIFF[19]) );
  XOR2X1 U61 ( .A(n30), .B(n61), .Y(DIFF[18]) );
  XOR2X1 U62 ( .A(n31), .B(n62), .Y(DIFF[17]) );
  XOR2X1 U63 ( .A(\carry[16] ), .B(n63), .Y(DIFF[16]) );
  INVX2 U64 ( .A(B[47]), .Y(n32) );
  INVX2 U65 ( .A(B[46]), .Y(n33) );
  INVX2 U66 ( .A(B[45]), .Y(n34) );
  INVX2 U67 ( .A(B[44]), .Y(n35) );
  INVX2 U68 ( .A(B[43]), .Y(n36) );
  INVX2 U69 ( .A(B[42]), .Y(n37) );
  INVX2 U70 ( .A(B[41]), .Y(n38) );
  INVX2 U71 ( .A(B[40]), .Y(n39) );
  INVX2 U72 ( .A(B[39]), .Y(n40) );
  INVX2 U73 ( .A(B[38]), .Y(n41) );
  INVX2 U74 ( .A(B[37]), .Y(n42) );
  INVX2 U75 ( .A(B[36]), .Y(n43) );
  INVX2 U76 ( .A(B[35]), .Y(n44) );
  INVX2 U77 ( .A(B[34]), .Y(n45) );
  INVX2 U78 ( .A(B[33]), .Y(n46) );
  INVX2 U79 ( .A(B[32]), .Y(n47) );
  INVX2 U80 ( .A(B[31]), .Y(n48) );
  INVX2 U81 ( .A(B[30]), .Y(n49) );
  INVX2 U82 ( .A(B[29]), .Y(n50) );
  INVX2 U83 ( .A(B[28]), .Y(n51) );
  INVX2 U84 ( .A(B[27]), .Y(n52) );
  INVX2 U85 ( .A(B[26]), .Y(n53) );
  INVX2 U86 ( .A(B[25]), .Y(n54) );
  INVX2 U87 ( .A(B[24]), .Y(n55) );
  INVX2 U88 ( .A(B[23]), .Y(n56) );
  INVX2 U89 ( .A(B[22]), .Y(n57) );
  INVX2 U90 ( .A(B[21]), .Y(n58) );
  INVX2 U91 ( .A(B[20]), .Y(n59) );
  INVX2 U92 ( .A(B[19]), .Y(n60) );
  INVX2 U93 ( .A(B[18]), .Y(n61) );
  INVX2 U94 ( .A(B[17]), .Y(n62) );
  INVX2 U95 ( .A(B[16]), .Y(n63) );
  NOR2X1 U96 ( .A(n64), .B(n65), .Y(\carry[16] ) );
  NAND3X1 U97 ( .A(n66), .B(n67), .C(n68), .Y(n65) );
  AND2X1 U98 ( .A(n70), .B(n69), .Y(n68) );
  NOR2X1 U99 ( .A(B[1]), .B(B[15]), .Y(n70) );
  NOR2X1 U100 ( .A(B[14]), .B(B[13]), .Y(n69) );
  NOR2X1 U101 ( .A(B[12]), .B(B[11]), .Y(n67) );
  NOR2X1 U102 ( .A(B[10]), .B(B[0]), .Y(n66) );
  NAND3X1 U103 ( .A(n71), .B(n72), .C(n73), .Y(n64) );
  AND2X1 U104 ( .A(n74), .B(n75), .Y(n73) );
  NOR2X1 U105 ( .A(B[9]), .B(B[8]), .Y(n75) );
  NOR2X1 U106 ( .A(B[7]), .B(B[6]), .Y(n74) );
  NOR2X1 U107 ( .A(B[5]), .B(B[4]), .Y(n72) );
  NOR2X1 U108 ( .A(B[3]), .B(B[2]), .Y(n71) );
endmodule


module poly5_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND2X2 U1 ( .A(n17), .B(n45), .Y(n1) );
  AND2X2 U2 ( .A(n18), .B(n47), .Y(n2) );
  AND2X2 U3 ( .A(n19), .B(n49), .Y(n3) );
  AND2X2 U4 ( .A(n20), .B(n51), .Y(n4) );
  AND2X2 U5 ( .A(n21), .B(n53), .Y(n5) );
  AND2X2 U6 ( .A(n22), .B(n55), .Y(n6) );
  AND2X2 U7 ( .A(n23), .B(n57), .Y(n7) );
  AND2X2 U8 ( .A(n24), .B(n59), .Y(n8) );
  AND2X2 U9 ( .A(n26), .B(n33), .Y(n9) );
  AND2X2 U10 ( .A(n27), .B(n35), .Y(n10) );
  AND2X2 U11 ( .A(n28), .B(n37), .Y(n11) );
  AND2X2 U12 ( .A(n29), .B(n39), .Y(n12) );
  AND2X2 U13 ( .A(n15), .B(n41), .Y(n13) );
  AND2X2 U14 ( .A(n16), .B(n43), .Y(n14) );
  AND2X2 U15 ( .A(n14), .B(n42), .Y(n15) );
  AND2X2 U16 ( .A(n1), .B(n44), .Y(n16) );
  AND2X2 U17 ( .A(n2), .B(n46), .Y(n17) );
  AND2X2 U18 ( .A(n3), .B(n48), .Y(n18) );
  AND2X2 U19 ( .A(n4), .B(n50), .Y(n19) );
  AND2X2 U20 ( .A(n5), .B(n52), .Y(n20) );
  AND2X2 U21 ( .A(n6), .B(n54), .Y(n21) );
  AND2X2 U22 ( .A(n7), .B(n56), .Y(n22) );
  AND2X2 U23 ( .A(n8), .B(n58), .Y(n23) );
  AND2X2 U24 ( .A(n61), .B(n60), .Y(n24) );
  AND2X2 U25 ( .A(n9), .B(n32), .Y(n25) );
  AND2X2 U26 ( .A(n10), .B(n34), .Y(n26) );
  AND2X2 U27 ( .A(n11), .B(n36), .Y(n27) );
  AND2X2 U28 ( .A(n12), .B(n38), .Y(n28) );
  AND2X2 U29 ( .A(n13), .B(n40), .Y(n29) );
  XOR2X1 U30 ( .A(B[31]), .B(n30), .Y(DIFF[31]) );
  XOR2X1 U31 ( .A(n25), .B(n31), .Y(DIFF[30]) );
  NAND2X1 U32 ( .A(n25), .B(n31), .Y(n30) );
  XOR2X1 U33 ( .A(n9), .B(n32), .Y(DIFF[29]) );
  XOR2X1 U34 ( .A(n26), .B(n33), .Y(DIFF[28]) );
  XOR2X1 U35 ( .A(n10), .B(n34), .Y(DIFF[27]) );
  XOR2X1 U36 ( .A(n27), .B(n35), .Y(DIFF[26]) );
  XOR2X1 U37 ( .A(n11), .B(n36), .Y(DIFF[25]) );
  XOR2X1 U38 ( .A(n28), .B(n37), .Y(DIFF[24]) );
  XOR2X1 U39 ( .A(n12), .B(n38), .Y(DIFF[23]) );
  XOR2X1 U40 ( .A(n29), .B(n39), .Y(DIFF[22]) );
  XOR2X1 U41 ( .A(n13), .B(n40), .Y(DIFF[21]) );
  XOR2X1 U42 ( .A(n15), .B(n41), .Y(DIFF[20]) );
  XOR2X1 U43 ( .A(n14), .B(n42), .Y(DIFF[19]) );
  XOR2X1 U44 ( .A(n16), .B(n43), .Y(DIFF[18]) );
  XOR2X1 U45 ( .A(n1), .B(n44), .Y(DIFF[17]) );
  XOR2X1 U46 ( .A(n17), .B(n45), .Y(DIFF[16]) );
  XOR2X1 U47 ( .A(n2), .B(n46), .Y(DIFF[15]) );
  XOR2X1 U48 ( .A(n18), .B(n47), .Y(DIFF[14]) );
  XOR2X1 U49 ( .A(n3), .B(n48), .Y(DIFF[13]) );
  XOR2X1 U50 ( .A(n19), .B(n49), .Y(DIFF[12]) );
  XOR2X1 U51 ( .A(n4), .B(n50), .Y(DIFF[11]) );
  XOR2X1 U52 ( .A(n20), .B(n51), .Y(DIFF[10]) );
  XOR2X1 U53 ( .A(n5), .B(n52), .Y(DIFF[9]) );
  XOR2X1 U54 ( .A(n21), .B(n53), .Y(DIFF[8]) );
  XOR2X1 U55 ( .A(n6), .B(n54), .Y(DIFF[7]) );
  XOR2X1 U56 ( .A(n22), .B(n55), .Y(DIFF[6]) );
  XOR2X1 U57 ( .A(n7), .B(n56), .Y(DIFF[5]) );
  XOR2X1 U58 ( .A(n23), .B(n57), .Y(DIFF[4]) );
  XOR2X1 U59 ( .A(n8), .B(n58), .Y(DIFF[3]) );
  XOR2X1 U60 ( .A(n24), .B(n59), .Y(DIFF[2]) );
  XOR2X1 U61 ( .A(n61), .B(n60), .Y(DIFF[1]) );
  INVX2 U62 ( .A(B[30]), .Y(n31) );
  INVX2 U63 ( .A(B[29]), .Y(n32) );
  INVX2 U64 ( .A(B[28]), .Y(n33) );
  INVX2 U65 ( .A(B[27]), .Y(n34) );
  INVX2 U66 ( .A(B[26]), .Y(n35) );
  INVX2 U67 ( .A(B[25]), .Y(n36) );
  INVX2 U68 ( .A(B[24]), .Y(n37) );
  INVX2 U69 ( .A(B[23]), .Y(n38) );
  INVX2 U70 ( .A(B[22]), .Y(n39) );
  INVX2 U71 ( .A(B[21]), .Y(n40) );
  INVX2 U72 ( .A(B[20]), .Y(n41) );
  INVX2 U73 ( .A(B[19]), .Y(n42) );
  INVX2 U74 ( .A(B[18]), .Y(n43) );
  INVX2 U75 ( .A(B[17]), .Y(n44) );
  INVX2 U76 ( .A(B[16]), .Y(n45) );
  INVX2 U77 ( .A(B[15]), .Y(n46) );
  INVX2 U78 ( .A(B[14]), .Y(n47) );
  INVX2 U79 ( .A(B[13]), .Y(n48) );
  INVX2 U80 ( .A(B[12]), .Y(n49) );
  INVX2 U81 ( .A(B[11]), .Y(n50) );
  INVX2 U82 ( .A(B[10]), .Y(n51) );
  INVX2 U83 ( .A(B[9]), .Y(n52) );
  INVX2 U84 ( .A(B[8]), .Y(n53) );
  INVX2 U85 ( .A(B[7]), .Y(n54) );
  INVX2 U86 ( .A(B[6]), .Y(n55) );
  INVX2 U87 ( .A(B[5]), .Y(n56) );
  INVX2 U88 ( .A(B[4]), .Y(n57) );
  INVX2 U89 ( .A(B[3]), .Y(n58) );
  INVX2 U90 ( .A(B[2]), .Y(n59) );
  INVX2 U91 ( .A(B[1]), .Y(n60) );
  INVX2 U92 ( .A(\B[0] ), .Y(n61) );
endmodule


module poly5_DW01_sub_10 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  AND2X2 U1 ( .A(n16), .B(n33), .Y(n1) );
  AND2X2 U2 ( .A(n17), .B(n35), .Y(n2) );
  AND2X2 U3 ( .A(n18), .B(n37), .Y(n3) );
  AND2X2 U4 ( .A(n19), .B(n39), .Y(n4) );
  AND2X2 U5 ( .A(n20), .B(n41), .Y(n5) );
  AND2X2 U6 ( .A(n21), .B(n43), .Y(n6) );
  AND2X2 U7 ( .A(n22), .B(n45), .Y(n7) );
  AND2X2 U8 ( .A(n23), .B(n47), .Y(n8) );
  AND2X2 U9 ( .A(n24), .B(n49), .Y(n9) );
  AND2X2 U10 ( .A(n25), .B(n51), .Y(n10) );
  AND2X2 U11 ( .A(n26), .B(n53), .Y(n11) );
  AND2X2 U12 ( .A(n27), .B(n55), .Y(n12) );
  AND2X2 U13 ( .A(n28), .B(n57), .Y(n13) );
  AND2X2 U14 ( .A(n29), .B(n59), .Y(n14) );
  AND2X2 U15 ( .A(n1), .B(n32), .Y(n15) );
  AND2X2 U16 ( .A(n2), .B(n34), .Y(n16) );
  AND2X2 U17 ( .A(n3), .B(n36), .Y(n17) );
  AND2X2 U18 ( .A(n4), .B(n38), .Y(n18) );
  AND2X2 U19 ( .A(n5), .B(n40), .Y(n19) );
  AND2X2 U20 ( .A(n6), .B(n42), .Y(n20) );
  AND2X2 U21 ( .A(n7), .B(n44), .Y(n21) );
  AND2X2 U22 ( .A(n8), .B(n46), .Y(n22) );
  AND2X2 U23 ( .A(n9), .B(n48), .Y(n23) );
  AND2X2 U24 ( .A(n10), .B(n50), .Y(n24) );
  AND2X2 U25 ( .A(n11), .B(n52), .Y(n25) );
  AND2X2 U26 ( .A(n12), .B(n54), .Y(n26) );
  AND2X2 U27 ( .A(n13), .B(n56), .Y(n27) );
  AND2X2 U28 ( .A(n14), .B(n58), .Y(n28) );
  AND2X2 U29 ( .A(n61), .B(n60), .Y(n29) );
  XOR2X1 U30 ( .A(B[31]), .B(n30), .Y(DIFF[31]) );
  XOR2X1 U31 ( .A(n15), .B(n31), .Y(DIFF[30]) );
  NAND2X1 U32 ( .A(n15), .B(n31), .Y(n30) );
  XOR2X1 U33 ( .A(n1), .B(n32), .Y(DIFF[29]) );
  XOR2X1 U34 ( .A(n16), .B(n33), .Y(DIFF[28]) );
  XOR2X1 U35 ( .A(n2), .B(n34), .Y(DIFF[27]) );
  XOR2X1 U36 ( .A(n17), .B(n35), .Y(DIFF[26]) );
  XOR2X1 U37 ( .A(n3), .B(n36), .Y(DIFF[25]) );
  XOR2X1 U38 ( .A(n18), .B(n37), .Y(DIFF[24]) );
  XOR2X1 U39 ( .A(n4), .B(n38), .Y(DIFF[23]) );
  XOR2X1 U40 ( .A(n19), .B(n39), .Y(DIFF[22]) );
  XOR2X1 U41 ( .A(n5), .B(n40), .Y(DIFF[21]) );
  XOR2X1 U42 ( .A(n20), .B(n41), .Y(DIFF[20]) );
  XOR2X1 U43 ( .A(n6), .B(n42), .Y(DIFF[19]) );
  XOR2X1 U44 ( .A(n21), .B(n43), .Y(DIFF[18]) );
  XOR2X1 U45 ( .A(n7), .B(n44), .Y(DIFF[17]) );
  XOR2X1 U46 ( .A(n22), .B(n45), .Y(DIFF[16]) );
  XOR2X1 U47 ( .A(n8), .B(n46), .Y(DIFF[15]) );
  XOR2X1 U48 ( .A(n23), .B(n47), .Y(DIFF[14]) );
  XOR2X1 U49 ( .A(n9), .B(n48), .Y(DIFF[13]) );
  XOR2X1 U50 ( .A(n24), .B(n49), .Y(DIFF[12]) );
  XOR2X1 U51 ( .A(n10), .B(n50), .Y(DIFF[11]) );
  XOR2X1 U52 ( .A(n25), .B(n51), .Y(DIFF[10]) );
  XOR2X1 U53 ( .A(n11), .B(n52), .Y(DIFF[9]) );
  XOR2X1 U54 ( .A(n26), .B(n53), .Y(DIFF[8]) );
  XOR2X1 U55 ( .A(n12), .B(n54), .Y(DIFF[7]) );
  XOR2X1 U56 ( .A(n27), .B(n55), .Y(DIFF[6]) );
  XOR2X1 U57 ( .A(n13), .B(n56), .Y(DIFF[5]) );
  XOR2X1 U58 ( .A(n28), .B(n57), .Y(DIFF[4]) );
  XOR2X1 U59 ( .A(n14), .B(n58), .Y(DIFF[3]) );
  XOR2X1 U60 ( .A(n29), .B(n59), .Y(DIFF[2]) );
  XOR2X1 U61 ( .A(n61), .B(n60), .Y(DIFF[1]) );
  INVX2 U62 ( .A(B[30]), .Y(n31) );
  INVX2 U63 ( .A(B[29]), .Y(n32) );
  INVX2 U64 ( .A(B[28]), .Y(n33) );
  INVX2 U65 ( .A(B[27]), .Y(n34) );
  INVX2 U66 ( .A(B[26]), .Y(n35) );
  INVX2 U67 ( .A(B[25]), .Y(n36) );
  INVX2 U68 ( .A(B[24]), .Y(n37) );
  INVX2 U69 ( .A(B[23]), .Y(n38) );
  INVX2 U70 ( .A(B[22]), .Y(n39) );
  INVX2 U71 ( .A(B[21]), .Y(n40) );
  INVX2 U72 ( .A(B[20]), .Y(n41) );
  INVX2 U73 ( .A(B[19]), .Y(n42) );
  INVX2 U74 ( .A(B[18]), .Y(n43) );
  INVX2 U75 ( .A(B[17]), .Y(n44) );
  INVX2 U76 ( .A(B[16]), .Y(n45) );
  INVX2 U77 ( .A(B[15]), .Y(n46) );
  INVX2 U78 ( .A(B[14]), .Y(n47) );
  INVX2 U79 ( .A(B[13]), .Y(n48) );
  INVX2 U80 ( .A(B[12]), .Y(n49) );
  INVX2 U81 ( .A(B[11]), .Y(n50) );
  INVX2 U82 ( .A(B[10]), .Y(n51) );
  INVX2 U83 ( .A(B[9]), .Y(n52) );
  INVX2 U84 ( .A(B[8]), .Y(n53) );
  INVX2 U85 ( .A(B[7]), .Y(n54) );
  INVX2 U86 ( .A(B[6]), .Y(n55) );
  INVX2 U87 ( .A(B[5]), .Y(n56) );
  INVX2 U88 ( .A(B[4]), .Y(n57) );
  INVX2 U89 ( .A(B[3]), .Y(n58) );
  INVX2 U90 ( .A(B[2]), .Y(n59) );
  INVX2 U91 ( .A(B[1]), .Y(n60) );
  INVX2 U92 ( .A(\B[0] ), .Y(n61) );
endmodule


module poly5_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module poly5_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module poly5_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(B[1]), .C(n1), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module poly5_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FAX1 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .YS(SUM[31]) );
  FAX1 U1_30 ( .A(A[30]), .B(B[30]), .C(carry[30]), .YC(carry[31]), .YS(
        SUM[30]) );
  FAX1 U1_29 ( .A(A[29]), .B(B[29]), .C(carry[29]), .YC(carry[30]), .YS(
        SUM[29]) );
  FAX1 U1_28 ( .A(A[28]), .B(B[28]), .C(carry[28]), .YC(carry[29]), .YS(
        SUM[28]) );
  FAX1 U1_27 ( .A(A[27]), .B(B[27]), .C(carry[27]), .YC(carry[28]), .YS(
        SUM[27]) );
  FAX1 U1_26 ( .A(A[26]), .B(B[26]), .C(carry[26]), .YC(carry[27]), .YS(
        SUM[26]) );
  FAX1 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .YC(carry[26]), .YS(
        SUM[25]) );
  FAX1 U1_24 ( .A(A[24]), .B(B[24]), .C(carry[24]), .YC(carry[25]), .YS(
        SUM[24]) );
  FAX1 U1_23 ( .A(A[23]), .B(B[23]), .C(carry[23]), .YC(carry[24]), .YS(
        SUM[23]) );
  FAX1 U1_22 ( .A(A[22]), .B(B[22]), .C(carry[22]), .YC(carry[23]), .YS(
        SUM[22]) );
  FAX1 U1_21 ( .A(A[21]), .B(B[21]), .C(carry[21]), .YC(carry[22]), .YS(
        SUM[21]) );
  FAX1 U1_20 ( .A(A[20]), .B(B[20]), .C(carry[20]), .YC(carry[21]), .YS(
        SUM[20]) );
  FAX1 U1_19 ( .A(A[19]), .B(B[19]), .C(carry[19]), .YC(carry[20]), .YS(
        SUM[19]) );
  FAX1 U1_18 ( .A(A[18]), .B(B[18]), .C(carry[18]), .YC(carry[19]), .YS(
        SUM[18]) );
  FAX1 U1_17 ( .A(A[17]), .B(B[17]), .C(carry[17]), .YC(carry[18]), .YS(
        SUM[17]) );
  FAX1 U1_16 ( .A(A[16]), .B(B[16]), .C(carry[16]), .YC(carry[17]), .YS(
        SUM[16]) );
  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YC(carry[16]), .YS(
        SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  FAX1 U1_4 ( .A(A[4]), .B(B[4]), .C(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  FAX1 U1_3 ( .A(A[3]), .B(B[3]), .C(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  FAX1 U1_2 ( .A(A[2]), .B(B[2]), .C(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  FAX1 U1_1 ( .A(A[1]), .B(n1), .C(B[1]), .YC(carry[2]), .YS(SUM[1]) );
  AND2X2 U1 ( .A(B[0]), .B(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(B[0]), .B(A[0]), .Y(SUM[0]) );
endmodule


module poly5_DW_mult_uns_4 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n2132, n2135, n2138, n2141, n2144, n2147, n2150, n2153, n2156, n2159,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732;
  assign n2132 = a[2];
  assign n2135 = a[5];
  assign n2138 = a[8];
  assign n2141 = a[11];
  assign n2144 = a[14];
  assign n2147 = a[17];
  assign n2150 = a[20];
  assign n2153 = a[23];
  assign n2156 = a[26];
  assign n2159 = a[29];

  FAX1 U336 ( .A(n2406), .B(n2417), .C(n2353), .YC(n2352), .YS(product[46]) );
  FAX1 U337 ( .A(n2431), .B(n2418), .C(n2354), .YC(n2353), .YS(product[45]) );
  FAX1 U338 ( .A(n2444), .B(n2432), .C(n2355), .YC(n2354), .YS(product[44]) );
  FAX1 U339 ( .A(n2445), .B(n2458), .C(n2356), .YC(n2355), .YS(product[43]) );
  FAX1 U340 ( .A(n2474), .B(n2459), .C(n2357), .YC(n2356), .YS(product[42]) );
  FAX1 U341 ( .A(n2489), .B(n2475), .C(n2358), .YC(n2357), .YS(product[41]) );
  FAX1 U342 ( .A(n2490), .B(n2504), .C(n2359), .YC(n2358), .YS(product[40]) );
  FAX1 U343 ( .A(n2522), .B(n2505), .C(n2360), .YC(n2359), .YS(product[39]) );
  FAX1 U344 ( .A(n2539), .B(n2523), .C(n2361), .YC(n2360), .YS(product[38]) );
  FAX1 U345 ( .A(n2540), .B(n2556), .C(n2362), .YC(n2361), .YS(product[37]) );
  FAX1 U346 ( .A(n2574), .B(n2557), .C(n2363), .YC(n2362), .YS(product[36]) );
  FAX1 U347 ( .A(n2592), .B(n2575), .C(n2364), .YC(n2363), .YS(product[35]) );
  FAX1 U348 ( .A(n2593), .B(n2610), .C(n2365), .YC(n2364), .YS(product[34]) );
  FAX1 U349 ( .A(n2628), .B(n2611), .C(n2366), .YC(n2365), .YS(product[33]) );
  FAX1 U350 ( .A(n3629), .B(n2629), .C(n2367), .YC(n2366), .YS(product[32]) );
  FAX1 U351 ( .A(n2647), .B(n3630), .C(n2368), .YC(n2367), .YS(product[31]) );
  FAX1 U352 ( .A(n2665), .B(n3631), .C(n2369), .YC(n2368), .YS(product[30]) );
  FAX1 U353 ( .A(n2683), .B(n3632), .C(n2370), .YC(n2369), .YS(product[29]) );
  FAX1 U354 ( .A(n2701), .B(n3633), .C(n2371), .YC(n2370), .YS(product[28]) );
  FAX1 U355 ( .A(n2719), .B(n3634), .C(n2372), .YC(n2371), .YS(product[27]) );
  FAX1 U356 ( .A(n2737), .B(n3635), .C(n2373), .YC(n2372), .YS(product[26]) );
  FAX1 U357 ( .A(n2753), .B(n3636), .C(n2374), .YC(n2373), .YS(product[25]) );
  FAX1 U358 ( .A(n2769), .B(n3637), .C(n2375), .YC(n2374), .YS(product[24]) );
  FAX1 U359 ( .A(n2785), .B(n3638), .C(n2376), .YC(n2375), .YS(product[23]) );
  FAX1 U360 ( .A(n2799), .B(n3639), .C(n2377), .YC(n2376), .YS(product[22]) );
  FAX1 U361 ( .A(n2813), .B(n3640), .C(n2378), .YC(n2377), .YS(product[21]) );
  FAX1 U362 ( .A(n2827), .B(n3641), .C(n2379), .YC(n2378), .YS(product[20]) );
  FAX1 U363 ( .A(n2839), .B(n3642), .C(n2380), .YC(n2379), .YS(product[19]) );
  FAX1 U364 ( .A(n2851), .B(n3643), .C(n2381), .YC(n2380), .YS(product[18]) );
  FAX1 U365 ( .A(n2863), .B(n3644), .C(n2382), .YC(n2381), .YS(product[17]) );
  FAX1 U366 ( .A(n2873), .B(n3645), .C(n2383), .YC(n2382), .YS(product[16]) );
  FAX1 U367 ( .A(n2883), .B(n3646), .C(n2384), .YC(n2383), .YS(product[15]) );
  FAX1 U368 ( .A(n2893), .B(n3647), .C(n2385), .YC(n2384), .YS(product[14]) );
  FAX1 U369 ( .A(n2901), .B(n3648), .C(n2386), .YC(n2385), .YS(product[13]) );
  FAX1 U370 ( .A(n2909), .B(n3649), .C(n2387), .YC(n2386), .YS(product[12]) );
  FAX1 U371 ( .A(n2917), .B(n3650), .C(n2388), .YC(n2387), .YS(product[11]) );
  FAX1 U372 ( .A(n2923), .B(n3651), .C(n2389), .YC(n2388), .YS(product[10]) );
  FAX1 U373 ( .A(n2929), .B(n3652), .C(n2390), .YC(n2389), .YS(product[9]) );
  FAX1 U374 ( .A(n2935), .B(n3653), .C(n2391), .YC(n2390), .YS(product[8]) );
  FAX1 U375 ( .A(n2939), .B(n3654), .C(n2392), .YC(n2391), .YS(product[7]) );
  FAX1 U376 ( .A(n2943), .B(n3655), .C(n2393), .YC(n2392), .YS(product[6]) );
  FAX1 U377 ( .A(n2947), .B(n3656), .C(n2394), .YC(n2393), .YS(product[5]) );
  FAX1 U378 ( .A(n3657), .B(n2949), .C(n2395), .YC(n2394), .YS(product[4]) );
  FAX1 U379 ( .A(n2951), .B(n3658), .C(n2396), .YC(n2395), .YS(product[3]) );
  HAX1 U380 ( .A(n3659), .B(n2397), .YC(n2396), .YS(product[2]) );
  HAX1 U381 ( .A(n2398), .B(n3660), .YC(n2397), .YS(product[1]) );
  HAX1 U382 ( .A(n2132), .B(n3661), .YC(n2398), .YS(product[0]) );
  FAX1 U384 ( .A(n2408), .B(n3455), .C(n2419), .YC(n2405), .YS(n2406) );
  FAX1 U385 ( .A(n2410), .B(n2421), .C(n3425), .YC(n2407), .YS(n2408) );
  FAX1 U386 ( .A(n2412), .B(n3398), .C(n2423), .YC(n2409), .YS(n2410) );
  FAX1 U387 ( .A(n2414), .B(n2425), .C(n3374), .YC(n2411), .YS(n2412) );
  FAX1 U388 ( .A(n2416), .B(n3353), .C(n2427), .YC(n2413), .YS(n2414) );
  FAX1 U389 ( .A(n4644), .B(n2429), .C(n3336), .YC(n2415), .YS(n2416) );
  FAX1 U390 ( .A(n3456), .B(n2420), .C(n3488), .YC(n2417), .YS(n2418) );
  FAX1 U391 ( .A(n2435), .B(n2422), .C(n2433), .YC(n2419), .YS(n2420) );
  FAX1 U392 ( .A(n3399), .B(n2424), .C(n3426), .YC(n2421), .YS(n2422) );
  FAX1 U393 ( .A(n2439), .B(n2426), .C(n2437), .YC(n2423), .YS(n2424) );
  FAX1 U394 ( .A(n2441), .B(n2428), .C(n3375), .YC(n2425), .YS(n2426) );
  FAX1 U395 ( .A(n4709), .B(n3337), .C(n3354), .YC(n2427), .YS(n2428) );
  FAX1 U397 ( .A(n2446), .B(n2434), .C(n3489), .YC(n2431), .YS(n2432) );
  FAX1 U398 ( .A(n2448), .B(n2436), .C(n3457), .YC(n2433), .YS(n2434) );
  FAX1 U399 ( .A(n2450), .B(n2438), .C(n3427), .YC(n2435), .YS(n2436) );
  FAX1 U400 ( .A(n2452), .B(n2440), .C(n3400), .YC(n2437), .YS(n2438) );
  FAX1 U401 ( .A(n2454), .B(n2442), .C(n3376), .YC(n2439), .YS(n2440) );
  FAX1 U402 ( .A(n2456), .B(n4709), .C(n3355), .YC(n2441), .YS(n2442) );
  FAX1 U404 ( .A(n2447), .B(n3490), .C(n2460), .YC(n2444), .YS(n2445) );
  FAX1 U405 ( .A(n2449), .B(n2462), .C(n3458), .YC(n2446), .YS(n2447) );
  FAX1 U406 ( .A(n2451), .B(n3428), .C(n2464), .YC(n2448), .YS(n2449) );
  FAX1 U407 ( .A(n2453), .B(n2466), .C(n3401), .YC(n2450), .YS(n2451) );
  FAX1 U408 ( .A(n2455), .B(n3377), .C(n2468), .YC(n2452), .YS(n2453) );
  FAX1 U409 ( .A(n2457), .B(n3356), .C(n2470), .YC(n2454), .YS(n2455) );
  FAX1 U410 ( .A(n4649), .B(n2472), .C(n3338), .YC(n2456), .YS(n2457) );
  FAX1 U411 ( .A(n3491), .B(n2461), .C(n3523), .YC(n2458), .YS(n2459) );
  FAX1 U412 ( .A(n2478), .B(n2463), .C(n2476), .YC(n2460), .YS(n2461) );
  FAX1 U413 ( .A(n3429), .B(n2465), .C(n3459), .YC(n2462), .YS(n2463) );
  FAX1 U414 ( .A(n2482), .B(n2467), .C(n2480), .YC(n2464), .YS(n2465) );
  FAX1 U415 ( .A(n2484), .B(n2469), .C(n3402), .YC(n2466), .YS(n2467) );
  FAX1 U416 ( .A(n2486), .B(n2471), .C(n3378), .YC(n2468), .YS(n2469) );
  FAX1 U417 ( .A(n4714), .B(n3339), .C(n3357), .YC(n2470), .YS(n2471) );
  FAX1 U419 ( .A(n2491), .B(n2477), .C(n3524), .YC(n2474), .YS(n2475) );
  FAX1 U420 ( .A(n2493), .B(n2479), .C(n3492), .YC(n2476), .YS(n2477) );
  FAX1 U421 ( .A(n2495), .B(n2481), .C(n3460), .YC(n2478), .YS(n2479) );
  FAX1 U422 ( .A(n2497), .B(n2483), .C(n3430), .YC(n2480), .YS(n2481) );
  FAX1 U423 ( .A(n2499), .B(n2485), .C(n3403), .YC(n2482), .YS(n2483) );
  FAX1 U424 ( .A(n2501), .B(n2487), .C(n3379), .YC(n2484), .YS(n2485) );
  FAX1 U425 ( .A(n3340), .B(n4714), .C(n3358), .YC(n2486), .YS(n2487) );
  FAX1 U427 ( .A(n2492), .B(n3525), .C(n2506), .YC(n2489), .YS(n2490) );
  FAX1 U428 ( .A(n2494), .B(n2508), .C(n3493), .YC(n2491), .YS(n2492) );
  FAX1 U429 ( .A(n2496), .B(n3461), .C(n2510), .YC(n2493), .YS(n2494) );
  FAX1 U430 ( .A(n2498), .B(n2512), .C(n3431), .YC(n2495), .YS(n2496) );
  FAX1 U431 ( .A(n2500), .B(n3404), .C(n2514), .YC(n2497), .YS(n2498) );
  FAX1 U432 ( .A(n2502), .B(n3380), .C(n2516), .YC(n2499), .YS(n2500) );
  FAX1 U433 ( .A(n2503), .B(n2518), .C(n3359), .YC(n2501), .YS(n2502) );
  FAX1 U434 ( .A(n4654), .B(n2520), .C(n3341), .YC(n2472), .YS(n2503) );
  FAX1 U435 ( .A(n3526), .B(n2507), .C(n3558), .YC(n2504), .YS(n2505) );
  FAX1 U436 ( .A(n2526), .B(n2509), .C(n2524), .YC(n2506), .YS(n2507) );
  FAX1 U437 ( .A(n3462), .B(n2511), .C(n3494), .YC(n2508), .YS(n2509) );
  FAX1 U438 ( .A(n2530), .B(n2513), .C(n2528), .YC(n2510), .YS(n2511) );
  FAX1 U439 ( .A(n2532), .B(n2515), .C(n3432), .YC(n2512), .YS(n2513) );
  FAX1 U440 ( .A(n2534), .B(n2517), .C(n3405), .YC(n2514), .YS(n2515) );
  FAX1 U441 ( .A(n3360), .B(n2519), .C(n3381), .YC(n2516), .YS(n2517) );
  FAX1 U442 ( .A(n4718), .B(n3342), .C(n2536), .YC(n2518), .YS(n2519) );
  FAX1 U444 ( .A(n2541), .B(n2525), .C(n3559), .YC(n2522), .YS(n2523) );
  FAX1 U445 ( .A(n2543), .B(n2527), .C(n3527), .YC(n2524), .YS(n2525) );
  FAX1 U446 ( .A(n2545), .B(n2529), .C(n3495), .YC(n2526), .YS(n2527) );
  FAX1 U447 ( .A(n2547), .B(n2531), .C(n3463), .YC(n2528), .YS(n2529) );
  FAX1 U448 ( .A(n2549), .B(n2533), .C(n3433), .YC(n2530), .YS(n2531) );
  FAX1 U449 ( .A(n2551), .B(n2535), .C(n3406), .YC(n2532), .YS(n2533) );
  FAX1 U450 ( .A(n2553), .B(n2537), .C(n3382), .YC(n2534), .YS(n2535) );
  FAX1 U451 ( .A(n3343), .B(n4718), .C(n3361), .YC(n2536), .YS(n2537) );
  FAX1 U453 ( .A(n2542), .B(n3560), .C(n2558), .YC(n2539), .YS(n2540) );
  FAX1 U454 ( .A(n2544), .B(n2560), .C(n3528), .YC(n2541), .YS(n2542) );
  FAX1 U455 ( .A(n2546), .B(n3496), .C(n2562), .YC(n2543), .YS(n2544) );
  FAX1 U456 ( .A(n2548), .B(n2564), .C(n3464), .YC(n2545), .YS(n2546) );
  FAX1 U457 ( .A(n2550), .B(n3434), .C(n2566), .YC(n2547), .YS(n2548) );
  FAX1 U458 ( .A(n2552), .B(n3407), .C(n2568), .YC(n2549), .YS(n2550) );
  FAX1 U459 ( .A(n2554), .B(n2570), .C(n3383), .YC(n2551), .YS(n2552) );
  FAX1 U460 ( .A(n2555), .B(n2572), .C(n3362), .YC(n2553), .YS(n2554) );
  FAX1 U461 ( .A(n4746), .B(n4659), .C(n3344), .YC(n2520), .YS(n2555) );
  FAX1 U462 ( .A(n3561), .B(n2559), .C(n3593), .YC(n2556), .YS(n2557) );
  FAX1 U463 ( .A(n2578), .B(n2561), .C(n2576), .YC(n2558), .YS(n2559) );
  FAX1 U464 ( .A(n3497), .B(n2563), .C(n3529), .YC(n2560), .YS(n2561) );
  FAX1 U465 ( .A(n2582), .B(n2565), .C(n2580), .YC(n2562), .YS(n2563) );
  FAX1 U466 ( .A(n2584), .B(n2567), .C(n3465), .YC(n2564), .YS(n2565) );
  FAX1 U467 ( .A(n2586), .B(n2569), .C(n3435), .YC(n2566), .YS(n2567) );
  FAX1 U468 ( .A(n3384), .B(n2571), .C(n3408), .YC(n2568), .YS(n2569) );
  FAX1 U469 ( .A(n3363), .B(n2573), .C(n2588), .YC(n2570), .YS(n2571) );
  FAX1 U470 ( .A(n2132), .B(n3345), .C(n2590), .YC(n2572), .YS(n2573) );
  FAX1 U471 ( .A(n2594), .B(n2577), .C(n3594), .YC(n2574), .YS(n2575) );
  FAX1 U472 ( .A(n3530), .B(n2579), .C(n3562), .YC(n2576), .YS(n2577) );
  FAX1 U473 ( .A(n2598), .B(n2581), .C(n2596), .YC(n2578), .YS(n2579) );
  FAX1 U474 ( .A(n3466), .B(n2583), .C(n3498), .YC(n2580), .YS(n2581) );
  FAX1 U475 ( .A(n3436), .B(n2585), .C(n2600), .YC(n2582), .YS(n2583) );
  FAX1 U476 ( .A(n2604), .B(n2587), .C(n2602), .YC(n2584), .YS(n2585) );
  FAX1 U477 ( .A(n3385), .B(n2589), .C(n3409), .YC(n2586), .YS(n2587) );
  FAX1 U478 ( .A(n3364), .B(n2591), .C(n2606), .YC(n2588), .YS(n2589) );
  FAX1 U479 ( .A(n2132), .B(n3346), .C(n2608), .YC(n2590), .YS(n2591) );
  FAX1 U480 ( .A(n2595), .B(n2612), .C(n3595), .YC(n2592), .YS(n2593) );
  FAX1 U481 ( .A(n2597), .B(n2614), .C(n3563), .YC(n2594), .YS(n2595) );
  FAX1 U482 ( .A(n2599), .B(n2616), .C(n3531), .YC(n2596), .YS(n2597) );
  FAX1 U483 ( .A(n2601), .B(n2618), .C(n3499), .YC(n2598), .YS(n2599) );
  FAX1 U484 ( .A(n2603), .B(n2620), .C(n3467), .YC(n2600), .YS(n2601) );
  FAX1 U485 ( .A(n2605), .B(n2622), .C(n3437), .YC(n2602), .YS(n2603) );
  FAX1 U486 ( .A(n2607), .B(n2624), .C(n3410), .YC(n2604), .YS(n2605) );
  FAX1 U487 ( .A(n2609), .B(n2626), .C(n3386), .YC(n2606), .YS(n2607) );
  FAX1 U488 ( .A(n2132), .B(n3347), .C(n3365), .YC(n2608), .YS(n2609) );
  FAX1 U489 ( .A(n2613), .B(n3596), .C(n3628), .YC(n2610), .YS(n2611) );
  FAX1 U490 ( .A(n2615), .B(n3564), .C(n2630), .YC(n2612), .YS(n2613) );
  FAX1 U491 ( .A(n2617), .B(n3532), .C(n2632), .YC(n2614), .YS(n2615) );
  FAX1 U492 ( .A(n2619), .B(n3500), .C(n2634), .YC(n2616), .YS(n2617) );
  FAX1 U493 ( .A(n2621), .B(n3468), .C(n2636), .YC(n2618), .YS(n2619) );
  FAX1 U494 ( .A(n2623), .B(n3438), .C(n2638), .YC(n2620), .YS(n2621) );
  FAX1 U495 ( .A(n2625), .B(n3411), .C(n2640), .YC(n2622), .YS(n2623) );
  FAX1 U496 ( .A(n2627), .B(n3387), .C(n2642), .YC(n2624), .YS(n2625) );
  FAX1 U497 ( .A(n3348), .B(n3366), .C(n2644), .YC(n2626), .YS(n2627) );
  FAX1 U498 ( .A(n2631), .B(n3597), .C(n2646), .YC(n2628), .YS(n2629) );
  FAX1 U499 ( .A(n2633), .B(n3565), .C(n2648), .YC(n2630), .YS(n2631) );
  FAX1 U500 ( .A(n2635), .B(n3533), .C(n2650), .YC(n2632), .YS(n2633) );
  FAX1 U501 ( .A(n2637), .B(n3501), .C(n2652), .YC(n2634), .YS(n2635) );
  FAX1 U502 ( .A(n2639), .B(n3469), .C(n2654), .YC(n2636), .YS(n2637) );
  FAX1 U503 ( .A(n2641), .B(n3439), .C(n2656), .YC(n2638), .YS(n2639) );
  FAX1 U504 ( .A(n2643), .B(n3412), .C(n2658), .YC(n2640), .YS(n2641) );
  FAX1 U505 ( .A(n2645), .B(n3388), .C(n2660), .YC(n2642), .YS(n2643) );
  FAX1 U506 ( .A(n3349), .B(n3367), .C(n2662), .YC(n2644), .YS(n2645) );
  FAX1 U507 ( .A(n2649), .B(n3598), .C(n2664), .YC(n2646), .YS(n2647) );
  FAX1 U508 ( .A(n2651), .B(n3566), .C(n2666), .YC(n2648), .YS(n2649) );
  FAX1 U509 ( .A(n2653), .B(n3534), .C(n2668), .YC(n2650), .YS(n2651) );
  FAX1 U510 ( .A(n2655), .B(n3502), .C(n2670), .YC(n2652), .YS(n2653) );
  FAX1 U511 ( .A(n2657), .B(n3470), .C(n2672), .YC(n2654), .YS(n2655) );
  FAX1 U512 ( .A(n2659), .B(n3440), .C(n2674), .YC(n2656), .YS(n2657) );
  FAX1 U513 ( .A(n2661), .B(n3413), .C(n2676), .YC(n2658), .YS(n2659) );
  FAX1 U514 ( .A(n2663), .B(n3389), .C(n2678), .YC(n2660), .YS(n2661) );
  FAX1 U515 ( .A(n3350), .B(n3368), .C(n2680), .YC(n2662), .YS(n2663) );
  FAX1 U516 ( .A(n2667), .B(n3599), .C(n2682), .YC(n2664), .YS(n2665) );
  FAX1 U517 ( .A(n2669), .B(n3567), .C(n2684), .YC(n2666), .YS(n2667) );
  FAX1 U518 ( .A(n2671), .B(n3535), .C(n2686), .YC(n2668), .YS(n2669) );
  FAX1 U519 ( .A(n2673), .B(n3503), .C(n2688), .YC(n2670), .YS(n2671) );
  FAX1 U520 ( .A(n2675), .B(n3471), .C(n2690), .YC(n2672), .YS(n2673) );
  FAX1 U521 ( .A(n2677), .B(n3441), .C(n2692), .YC(n2674), .YS(n2675) );
  FAX1 U522 ( .A(n2679), .B(n3414), .C(n2694), .YC(n2676), .YS(n2677) );
  FAX1 U523 ( .A(n2681), .B(n3390), .C(n2696), .YC(n2678), .YS(n2679) );
  FAX1 U524 ( .A(n3351), .B(n3369), .C(n2698), .YC(n2680), .YS(n2681) );
  FAX1 U525 ( .A(n2685), .B(n3600), .C(n2700), .YC(n2682), .YS(n2683) );
  FAX1 U526 ( .A(n2687), .B(n3568), .C(n2702), .YC(n2684), .YS(n2685) );
  FAX1 U527 ( .A(n2689), .B(n3536), .C(n2704), .YC(n2686), .YS(n2687) );
  FAX1 U528 ( .A(n2691), .B(n3504), .C(n2706), .YC(n2688), .YS(n2689) );
  FAX1 U529 ( .A(n2693), .B(n3472), .C(n2708), .YC(n2690), .YS(n2691) );
  FAX1 U530 ( .A(n2695), .B(n3442), .C(n2710), .YC(n2692), .YS(n2693) );
  FAX1 U531 ( .A(n2697), .B(n3415), .C(n2712), .YC(n2694), .YS(n2695) );
  FAX1 U532 ( .A(n2699), .B(n3391), .C(n2714), .YC(n2696), .YS(n2697) );
  HAX1 U533 ( .A(n3370), .B(n2716), .YC(n2698), .YS(n2699) );
  FAX1 U534 ( .A(n2703), .B(n3601), .C(n2718), .YC(n2700), .YS(n2701) );
  FAX1 U535 ( .A(n2705), .B(n3569), .C(n2720), .YC(n2702), .YS(n2703) );
  FAX1 U536 ( .A(n2707), .B(n3537), .C(n2722), .YC(n2704), .YS(n2705) );
  FAX1 U537 ( .A(n2709), .B(n3505), .C(n2724), .YC(n2706), .YS(n2707) );
  FAX1 U538 ( .A(n2711), .B(n3473), .C(n2726), .YC(n2708), .YS(n2709) );
  FAX1 U539 ( .A(n2713), .B(n3443), .C(n2728), .YC(n2710), .YS(n2711) );
  FAX1 U540 ( .A(n2715), .B(n3416), .C(n2730), .YC(n2712), .YS(n2713) );
  FAX1 U541 ( .A(n3392), .B(n2717), .C(n2732), .YC(n2714), .YS(n2715) );
  HAX1 U542 ( .A(n2734), .B(n3371), .YC(n2716), .YS(n2717) );
  FAX1 U543 ( .A(n2721), .B(n3602), .C(n2736), .YC(n2718), .YS(n2719) );
  FAX1 U544 ( .A(n2723), .B(n3570), .C(n2738), .YC(n2720), .YS(n2721) );
  FAX1 U545 ( .A(n2725), .B(n3538), .C(n2740), .YC(n2722), .YS(n2723) );
  FAX1 U546 ( .A(n2727), .B(n3506), .C(n2742), .YC(n2724), .YS(n2725) );
  FAX1 U547 ( .A(n2729), .B(n3474), .C(n2744), .YC(n2726), .YS(n2727) );
  FAX1 U548 ( .A(n2731), .B(n3444), .C(n2746), .YC(n2728), .YS(n2729) );
  FAX1 U549 ( .A(n2733), .B(n3417), .C(n2748), .YC(n2730), .YS(n2731) );
  FAX1 U550 ( .A(n2735), .B(n3393), .C(n2750), .YC(n2732), .YS(n2733) );
  HAX1 U551 ( .A(n2159), .B(n3372), .YC(n2734), .YS(n2735) );
  FAX1 U552 ( .A(n2739), .B(n3603), .C(n2752), .YC(n2736), .YS(n2737) );
  FAX1 U553 ( .A(n2741), .B(n3571), .C(n2754), .YC(n2738), .YS(n2739) );
  FAX1 U554 ( .A(n2743), .B(n3539), .C(n2756), .YC(n2740), .YS(n2741) );
  FAX1 U555 ( .A(n2745), .B(n3507), .C(n2758), .YC(n2742), .YS(n2743) );
  FAX1 U556 ( .A(n2747), .B(n3475), .C(n2760), .YC(n2744), .YS(n2745) );
  FAX1 U557 ( .A(n2749), .B(n3445), .C(n2762), .YC(n2746), .YS(n2747) );
  FAX1 U558 ( .A(n2751), .B(n3418), .C(n2764), .YC(n2748), .YS(n2749) );
  HAX1 U559 ( .A(n3394), .B(n2766), .YC(n2750), .YS(n2751) );
  FAX1 U560 ( .A(n2755), .B(n3604), .C(n2768), .YC(n2752), .YS(n2753) );
  FAX1 U561 ( .A(n2757), .B(n3572), .C(n2770), .YC(n2754), .YS(n2755) );
  FAX1 U562 ( .A(n2759), .B(n3540), .C(n2772), .YC(n2756), .YS(n2757) );
  FAX1 U563 ( .A(n2761), .B(n3508), .C(n2774), .YC(n2758), .YS(n2759) );
  FAX1 U564 ( .A(n2763), .B(n3476), .C(n2776), .YC(n2760), .YS(n2761) );
  FAX1 U565 ( .A(n2765), .B(n3446), .C(n2778), .YC(n2762), .YS(n2763) );
  FAX1 U566 ( .A(n3419), .B(n2767), .C(n2780), .YC(n2764), .YS(n2765) );
  HAX1 U567 ( .A(n2782), .B(n3395), .YC(n2766), .YS(n2767) );
  FAX1 U568 ( .A(n2771), .B(n3605), .C(n2784), .YC(n2768), .YS(n2769) );
  FAX1 U569 ( .A(n2773), .B(n3573), .C(n2786), .YC(n2770), .YS(n2771) );
  FAX1 U570 ( .A(n2775), .B(n3541), .C(n2788), .YC(n2772), .YS(n2773) );
  FAX1 U571 ( .A(n2777), .B(n3509), .C(n2790), .YC(n2774), .YS(n2775) );
  FAX1 U572 ( .A(n2779), .B(n3477), .C(n2792), .YC(n2776), .YS(n2777) );
  FAX1 U573 ( .A(n2781), .B(n3447), .C(n2794), .YC(n2778), .YS(n2779) );
  FAX1 U574 ( .A(n2783), .B(n3420), .C(n2796), .YC(n2780), .YS(n2781) );
  HAX1 U575 ( .A(n2156), .B(n3396), .YC(n2782), .YS(n2783) );
  FAX1 U576 ( .A(n2787), .B(n3606), .C(n2798), .YC(n2784), .YS(n2785) );
  FAX1 U577 ( .A(n2789), .B(n3574), .C(n2800), .YC(n2786), .YS(n2787) );
  FAX1 U578 ( .A(n2791), .B(n3542), .C(n2802), .YC(n2788), .YS(n2789) );
  FAX1 U579 ( .A(n2793), .B(n3510), .C(n2804), .YC(n2790), .YS(n2791) );
  FAX1 U580 ( .A(n2795), .B(n3478), .C(n2806), .YC(n2792), .YS(n2793) );
  FAX1 U581 ( .A(n2797), .B(n3448), .C(n2808), .YC(n2794), .YS(n2795) );
  HAX1 U582 ( .A(n3421), .B(n2810), .YC(n2796), .YS(n2797) );
  FAX1 U583 ( .A(n2801), .B(n3607), .C(n2812), .YC(n2798), .YS(n2799) );
  FAX1 U584 ( .A(n2803), .B(n3575), .C(n2814), .YC(n2800), .YS(n2801) );
  FAX1 U585 ( .A(n2805), .B(n3543), .C(n2816), .YC(n2802), .YS(n2803) );
  FAX1 U586 ( .A(n2807), .B(n3511), .C(n2818), .YC(n2804), .YS(n2805) );
  FAX1 U587 ( .A(n2809), .B(n3479), .C(n2820), .YC(n2806), .YS(n2807) );
  FAX1 U588 ( .A(n3449), .B(n2811), .C(n2822), .YC(n2808), .YS(n2809) );
  HAX1 U589 ( .A(n2824), .B(n3422), .YC(n2810), .YS(n2811) );
  FAX1 U590 ( .A(n2815), .B(n3608), .C(n2826), .YC(n2812), .YS(n2813) );
  FAX1 U591 ( .A(n2817), .B(n3576), .C(n2828), .YC(n2814), .YS(n2815) );
  FAX1 U592 ( .A(n2819), .B(n3544), .C(n2830), .YC(n2816), .YS(n2817) );
  FAX1 U593 ( .A(n2821), .B(n3512), .C(n2832), .YC(n2818), .YS(n2819) );
  FAX1 U594 ( .A(n2823), .B(n3480), .C(n2834), .YC(n2820), .YS(n2821) );
  FAX1 U595 ( .A(n2825), .B(n3450), .C(n2836), .YC(n2822), .YS(n2823) );
  HAX1 U596 ( .A(n4676), .B(n3423), .YC(n2824), .YS(n2825) );
  FAX1 U597 ( .A(n2829), .B(n3609), .C(n2838), .YC(n2826), .YS(n2827) );
  FAX1 U598 ( .A(n2831), .B(n3577), .C(n2840), .YC(n2828), .YS(n2829) );
  FAX1 U599 ( .A(n2833), .B(n3545), .C(n2842), .YC(n2830), .YS(n2831) );
  FAX1 U600 ( .A(n2835), .B(n3513), .C(n2844), .YC(n2832), .YS(n2833) );
  FAX1 U601 ( .A(n2837), .B(n3481), .C(n2846), .YC(n2834), .YS(n2835) );
  HAX1 U602 ( .A(n3451), .B(n2848), .YC(n2836), .YS(n2837) );
  FAX1 U603 ( .A(n2841), .B(n3610), .C(n2850), .YC(n2838), .YS(n2839) );
  FAX1 U604 ( .A(n2843), .B(n3578), .C(n2852), .YC(n2840), .YS(n2841) );
  FAX1 U605 ( .A(n2845), .B(n3546), .C(n2854), .YC(n2842), .YS(n2843) );
  FAX1 U606 ( .A(n2847), .B(n3514), .C(n2856), .YC(n2844), .YS(n2845) );
  FAX1 U607 ( .A(n3482), .B(n2849), .C(n2858), .YC(n2846), .YS(n2847) );
  HAX1 U608 ( .A(n2860), .B(n3452), .YC(n2848), .YS(n2849) );
  FAX1 U609 ( .A(n2853), .B(n3611), .C(n2862), .YC(n2850), .YS(n2851) );
  FAX1 U610 ( .A(n2855), .B(n3579), .C(n2864), .YC(n2852), .YS(n2853) );
  FAX1 U611 ( .A(n2857), .B(n3547), .C(n2866), .YC(n2854), .YS(n2855) );
  FAX1 U612 ( .A(n2859), .B(n3515), .C(n2868), .YC(n2856), .YS(n2857) );
  FAX1 U613 ( .A(n2861), .B(n3483), .C(n2870), .YC(n2858), .YS(n2859) );
  HAX1 U614 ( .A(n4678), .B(n3453), .YC(n2860), .YS(n2861) );
  FAX1 U615 ( .A(n2865), .B(n3612), .C(n2872), .YC(n2862), .YS(n2863) );
  FAX1 U616 ( .A(n2867), .B(n3580), .C(n2874), .YC(n2864), .YS(n2865) );
  FAX1 U617 ( .A(n2869), .B(n3548), .C(n2876), .YC(n2866), .YS(n2867) );
  FAX1 U618 ( .A(n2871), .B(n3516), .C(n2878), .YC(n2868), .YS(n2869) );
  HAX1 U619 ( .A(n3484), .B(n2880), .YC(n2870), .YS(n2871) );
  FAX1 U620 ( .A(n2875), .B(n3613), .C(n2882), .YC(n2872), .YS(n2873) );
  FAX1 U621 ( .A(n2877), .B(n3581), .C(n2884), .YC(n2874), .YS(n2875) );
  FAX1 U622 ( .A(n2879), .B(n3549), .C(n2886), .YC(n2876), .YS(n2877) );
  FAX1 U623 ( .A(n3517), .B(n2881), .C(n2888), .YC(n2878), .YS(n2879) );
  HAX1 U624 ( .A(n2890), .B(n3485), .YC(n2880), .YS(n2881) );
  FAX1 U625 ( .A(n2885), .B(n3614), .C(n2892), .YC(n2882), .YS(n2883) );
  FAX1 U626 ( .A(n2887), .B(n3582), .C(n2894), .YC(n2884), .YS(n2885) );
  FAX1 U627 ( .A(n2889), .B(n3550), .C(n2896), .YC(n2886), .YS(n2887) );
  FAX1 U628 ( .A(n2891), .B(n3518), .C(n2898), .YC(n2888), .YS(n2889) );
  HAX1 U629 ( .A(n2147), .B(n3486), .YC(n2890), .YS(n2891) );
  FAX1 U630 ( .A(n2895), .B(n3615), .C(n2900), .YC(n2892), .YS(n2893) );
  FAX1 U631 ( .A(n2897), .B(n3583), .C(n2902), .YC(n2894), .YS(n2895) );
  FAX1 U632 ( .A(n2899), .B(n3551), .C(n2904), .YC(n2896), .YS(n2897) );
  HAX1 U633 ( .A(n3519), .B(n2906), .YC(n2898), .YS(n2899) );
  FAX1 U634 ( .A(n2903), .B(n3616), .C(n2908), .YC(n2900), .YS(n2901) );
  FAX1 U635 ( .A(n2905), .B(n3584), .C(n2910), .YC(n2902), .YS(n2903) );
  FAX1 U636 ( .A(n3552), .B(n2907), .C(n2912), .YC(n2904), .YS(n2905) );
  HAX1 U637 ( .A(n2914), .B(n3520), .YC(n2906), .YS(n2907) );
  FAX1 U638 ( .A(n2911), .B(n3617), .C(n2916), .YC(n2908), .YS(n2909) );
  FAX1 U639 ( .A(n2913), .B(n3585), .C(n2918), .YC(n2910), .YS(n2911) );
  FAX1 U640 ( .A(n2915), .B(n3553), .C(n2920), .YC(n2912), .YS(n2913) );
  HAX1 U641 ( .A(n2144), .B(n3521), .YC(n2914), .YS(n2915) );
  FAX1 U642 ( .A(n2919), .B(n3618), .C(n2922), .YC(n2916), .YS(n2917) );
  FAX1 U643 ( .A(n2921), .B(n3586), .C(n2924), .YC(n2918), .YS(n2919) );
  HAX1 U644 ( .A(n3554), .B(n2926), .YC(n2920), .YS(n2921) );
  FAX1 U645 ( .A(n2925), .B(n3619), .C(n2928), .YC(n2922), .YS(n2923) );
  FAX1 U646 ( .A(n3587), .B(n2927), .C(n2930), .YC(n2924), .YS(n2925) );
  HAX1 U647 ( .A(n2932), .B(n3555), .YC(n2926), .YS(n2927) );
  FAX1 U648 ( .A(n2931), .B(n3620), .C(n2934), .YC(n2928), .YS(n2929) );
  FAX1 U649 ( .A(n2933), .B(n3588), .C(n2936), .YC(n2930), .YS(n2931) );
  HAX1 U650 ( .A(n2141), .B(n3556), .YC(n2932), .YS(n2933) );
  FAX1 U651 ( .A(n2937), .B(n3621), .C(n2938), .YC(n2934), .YS(n2935) );
  HAX1 U652 ( .A(n3589), .B(n2940), .YC(n2936), .YS(n2937) );
  FAX1 U653 ( .A(n3622), .B(n2941), .C(n2942), .YC(n2938), .YS(n2939) );
  HAX1 U654 ( .A(n2944), .B(n3590), .YC(n2940), .YS(n2941) );
  FAX1 U655 ( .A(n2945), .B(n3623), .C(n2946), .YC(n2942), .YS(n2943) );
  HAX1 U656 ( .A(n2138), .B(n3591), .YC(n2944), .YS(n2945) );
  HAX1 U657 ( .A(n3624), .B(n2948), .YC(n2946), .YS(n2947) );
  HAX1 U658 ( .A(n2950), .B(n3625), .YC(n2948), .YS(n2949) );
  HAX1 U659 ( .A(n2135), .B(n3626), .YC(n2950), .YS(n2951) );
  HAX1 U1990 ( .A(b[31]), .B(n3270), .YC(n3301), .YS(n3302) );
  FAX1 U1991 ( .A(b[31]), .B(n4633), .C(n3271), .YC(n3270), .YS(n3303) );
  FAX1 U1992 ( .A(n4633), .B(n4631), .C(n3272), .YC(n3271), .YS(n3304) );
  FAX1 U1993 ( .A(n4631), .B(n4629), .C(n3273), .YC(n3272), .YS(n3305) );
  FAX1 U1994 ( .A(n4629), .B(n4627), .C(n3274), .YC(n3273), .YS(n3306) );
  FAX1 U1995 ( .A(n4627), .B(n4625), .C(n3275), .YC(n3274), .YS(n3307) );
  FAX1 U1996 ( .A(n4625), .B(n4623), .C(n3276), .YC(n3275), .YS(n3308) );
  FAX1 U1997 ( .A(n4623), .B(n4621), .C(n3277), .YC(n3276), .YS(n3309) );
  FAX1 U1998 ( .A(b[24]), .B(n4619), .C(n3278), .YC(n3277), .YS(n3310) );
  FAX1 U1999 ( .A(n4619), .B(n4617), .C(n3279), .YC(n3278), .YS(n3311) );
  FAX1 U2000 ( .A(b[22]), .B(n4615), .C(n3280), .YC(n3279), .YS(n3312) );
  FAX1 U2001 ( .A(n4614), .B(n4612), .C(n3281), .YC(n3280), .YS(n3313) );
  FAX1 U2002 ( .A(n4612), .B(n4610), .C(n3282), .YC(n3281), .YS(n3314) );
  FAX1 U2003 ( .A(n4609), .B(n4607), .C(n3283), .YC(n3282), .YS(n3315) );
  FAX1 U2004 ( .A(b[18]), .B(n4604), .C(n3284), .YC(n3283), .YS(n3316) );
  FAX1 U2005 ( .A(n4604), .B(n4602), .C(n3285), .YC(n3284), .YS(n3317) );
  FAX1 U2006 ( .A(b[16]), .B(b[15]), .C(n3286), .YC(n3285), .YS(n3318) );
  FAX1 U2007 ( .A(n4600), .B(b[14]), .C(n3287), .YC(n3286), .YS(n3319) );
  FAX1 U2008 ( .A(n4598), .B(n4596), .C(n3288), .YC(n3287), .YS(n3320) );
  FAX1 U2009 ( .A(n4595), .B(b[12]), .C(n3289), .YC(n3288), .YS(n3321) );
  FAX1 U2010 ( .A(n4593), .B(n4591), .C(n3290), .YC(n3289), .YS(n3322) );
  FAX1 U2011 ( .A(n4590), .B(b[10]), .C(n3291), .YC(n3290), .YS(n3323) );
  FAX1 U2012 ( .A(n4588), .B(n4586), .C(n3292), .YC(n3291), .YS(n3324) );
  FAX1 U2013 ( .A(n4585), .B(b[8]), .C(n3293), .YC(n3292), .YS(n3325) );
  FAX1 U2014 ( .A(n4583), .B(b[7]), .C(n3294), .YC(n3293), .YS(n3326) );
  FAX1 U2015 ( .A(n4581), .B(b[6]), .C(n3295), .YC(n3294), .YS(n3327) );
  FAX1 U2016 ( .A(n4579), .B(n4577), .C(n3296), .YC(n3295), .YS(n3328) );
  FAX1 U2017 ( .A(n4576), .B(b[4]), .C(n3297), .YC(n3296), .YS(n3329) );
  FAX1 U2018 ( .A(n4574), .B(n4572), .C(n3298), .YC(n3297), .YS(n3330) );
  FAX1 U2019 ( .A(n4571), .B(b[2]), .C(n3299), .YC(n3298), .YS(n3331) );
  FAX1 U2020 ( .A(n4569), .B(n4680), .C(n3300), .YC(n3299), .YS(n3332) );
  HAX1 U2021 ( .A(n4680), .B(n4682), .YC(n3300), .YS(n3333) );
  OR2X2 U2024 ( .A(n4741), .B(n5388), .Y(n4552) );
  OR2X2 U2025 ( .A(n4876), .B(n4748), .Y(n4553) );
  OR2X2 U2026 ( .A(n5389), .B(n5390), .Y(n4554) );
  NAND2X1 U2027 ( .A(n5561), .B(n5559), .Y(n4555) );
  NAND2X1 U2028 ( .A(n4737), .B(n5632), .Y(n4556) );
  NAND2X1 U2029 ( .A(n4734), .B(n5695), .Y(n4557) );
  NAND2X1 U2030 ( .A(a[31]), .B(n4730), .Y(n4558) );
  INVX2 U2031 ( .A(n3332), .Y(n4724) );
  INVX2 U2032 ( .A(n3330), .Y(n4722) );
  INVX2 U2033 ( .A(n3320), .Y(n4710) );
  INVX2 U2034 ( .A(n3326), .Y(n4717) );
  INVX2 U2035 ( .A(n3318), .Y(n4707) );
  INVX2 U2036 ( .A(n3329), .Y(n4721) );
  INVX2 U2037 ( .A(n3328), .Y(n4720) );
  INVX2 U2038 ( .A(n3327), .Y(n4719) );
  INVX2 U2039 ( .A(n3331), .Y(n4723) );
  INVX2 U2040 ( .A(n3325), .Y(n4716) );
  INVX2 U2041 ( .A(n3324), .Y(n4715) );
  INVX2 U2042 ( .A(n3321), .Y(n4711) );
  INVX2 U2043 ( .A(n3323), .Y(n4713) );
  INVX2 U2044 ( .A(n3322), .Y(n4712) );
  INVX2 U2045 ( .A(n3319), .Y(n4708) );
  INVX2 U2046 ( .A(n3317), .Y(n4706) );
  INVX2 U2047 ( .A(n3316), .Y(n4705) );
  INVX2 U2048 ( .A(n3315), .Y(n4704) );
  INVX2 U2049 ( .A(n3314), .Y(n4703) );
  INVX2 U2050 ( .A(n3312), .Y(n4701) );
  INVX2 U2051 ( .A(n3313), .Y(n4702) );
  INVX2 U2052 ( .A(n3333), .Y(n4725) );
  INVX2 U2053 ( .A(n3311), .Y(n4700) );
  INVX2 U2054 ( .A(n4598), .Y(n4726) );
  INVX2 U2055 ( .A(n4681), .Y(n4680) );
  INVX2 U2056 ( .A(n4570), .Y(n4571) );
  INVX2 U2057 ( .A(n4580), .Y(n4581) );
  INVX2 U2058 ( .A(n4570), .Y(n4572) );
  INVX2 U2059 ( .A(n4575), .Y(n4576) );
  INVX2 U2060 ( .A(n4568), .Y(n4569) );
  INVX2 U2061 ( .A(n4578), .Y(n4579) );
  INVX2 U2062 ( .A(n4573), .Y(n4574) );
  INVX2 U2063 ( .A(n4683), .Y(n4686) );
  INVX2 U2064 ( .A(n4575), .Y(n4577) );
  INVX2 U2065 ( .A(n4582), .Y(n4583) );
  INVX2 U2066 ( .A(n4587), .Y(n4588) );
  INVX2 U2067 ( .A(n4584), .Y(n4585) );
  INVX2 U2068 ( .A(n4584), .Y(n4586) );
  INVX2 U2069 ( .A(n4594), .Y(n4595) );
  INVX2 U2070 ( .A(n4599), .Y(n4600) );
  INVX2 U2071 ( .A(n4594), .Y(n4596) );
  INVX2 U2072 ( .A(n4592), .Y(n4593) );
  INVX2 U2073 ( .A(n4597), .Y(n4598) );
  INVX2 U2074 ( .A(n4589), .Y(n4590) );
  INVX2 U2075 ( .A(n4589), .Y(n4591) );
  INVX2 U2076 ( .A(n4603), .Y(n4604) );
  INVX2 U2077 ( .A(n4608), .Y(n4609) );
  INVX2 U2078 ( .A(n4613), .Y(n4614) );
  INVX2 U2079 ( .A(n4601), .Y(n4602) );
  INVX2 U2080 ( .A(n4613), .Y(n4615) );
  INVX2 U2081 ( .A(n4608), .Y(n4610) );
  INVX2 U2082 ( .A(n4611), .Y(n4612) );
  INVX2 U2083 ( .A(n4603), .Y(n4605) );
  INVX2 U2084 ( .A(n4606), .Y(n4607) );
  INVX2 U2085 ( .A(n4616), .Y(n4617) );
  INVX2 U2086 ( .A(n4620), .Y(n4621) );
  BUFX2 U2087 ( .A(b[0]), .Y(n4682) );
  BUFX2 U2088 ( .A(b[0]), .Y(n4684) );
  BUFX2 U2089 ( .A(b[0]), .Y(n4683) );
  INVX1 U2090 ( .A(b[5]), .Y(n4575) );
  INVX1 U2091 ( .A(b[6]), .Y(n4578) );
  INVX1 U2092 ( .A(b[2]), .Y(n4568) );
  INVX1 U2093 ( .A(b[4]), .Y(n4573) );
  BUFX2 U2094 ( .A(b[0]), .Y(n4685) );
  INVX1 U2095 ( .A(b[8]), .Y(n4582) );
  INVX1 U2096 ( .A(b[10]), .Y(n4587) );
  INVX1 U2097 ( .A(b[9]), .Y(n4584) );
  INVX1 U2098 ( .A(b[12]), .Y(n4592) );
  INVX1 U2099 ( .A(b[14]), .Y(n4597) );
  INVX1 U2100 ( .A(b[11]), .Y(n4589) );
  INVX1 U2101 ( .A(b[20]), .Y(n4611) );
  INVX1 U2102 ( .A(b[18]), .Y(n4606) );
  INVX2 U2103 ( .A(n4618), .Y(n4619) );
  INVX2 U2104 ( .A(n4622), .Y(n4623) );
  INVX2 U2105 ( .A(n4624), .Y(n4625) );
  INVX1 U2106 ( .A(b[26]), .Y(n4624) );
  INVX1 U2107 ( .A(b[22]), .Y(n4616) );
  INVX2 U2108 ( .A(n4626), .Y(n4627) );
  INVX2 U2109 ( .A(n4630), .Y(n4631) );
  INVX2 U2110 ( .A(n4628), .Y(n4629) );
  INVX1 U2111 ( .A(b[28]), .Y(n4628) );
  INVX2 U2112 ( .A(n4632), .Y(n4633) );
  INVX1 U2113 ( .A(b[30]), .Y(n4632) );
  INVX2 U2114 ( .A(n5395), .Y(n4638) );
  INVX2 U2115 ( .A(n5484), .Y(n4634) );
  INVX2 U2116 ( .A(n4885), .Y(n4661) );
  INVX2 U2117 ( .A(n5194), .Y(n4646) );
  INVX2 U2118 ( .A(n5485), .Y(n4636) );
  INVX2 U2119 ( .A(n5085), .Y(n4652) );
  INVX2 U2120 ( .A(n5188), .Y(n4647) );
  INVX2 U2121 ( .A(n5291), .Y(n4642) );
  INVX2 U2122 ( .A(n4989), .Y(n4653) );
  INVX2 U2123 ( .A(n5092), .Y(n4648) );
  INVX2 U2124 ( .A(n4886), .Y(n4658) );
  INVX2 U2125 ( .A(n5195), .Y(n4643) );
  INVX2 U2126 ( .A(n4988), .Y(n4656) );
  INVX2 U2127 ( .A(n5091), .Y(n4651) );
  INVX2 U2128 ( .A(n4982), .Y(n4657) );
  INVX2 U2129 ( .A(n5637), .Y(n4731) );
  INVX2 U2130 ( .A(n5566), .Y(n4736) );
  INVX2 U2131 ( .A(n5638), .Y(n4733) );
  INVX2 U2132 ( .A(n5698), .Y(n4728) );
  INVX2 U2133 ( .A(n5699), .Y(n4729) );
  INVX2 U2134 ( .A(n5565), .Y(n4735) );
  INVX2 U2135 ( .A(n4559), .Y(n4668) );
  INVX2 U2136 ( .A(n4560), .Y(n4669) );
  INVX2 U2137 ( .A(n4562), .Y(n4670) );
  INVX2 U2138 ( .A(n4564), .Y(n4671) );
  INVX2 U2139 ( .A(n4561), .Y(n4664) );
  INVX2 U2140 ( .A(n4563), .Y(n4665) );
  INVX2 U2141 ( .A(n5558), .Y(n4635) );
  INVX2 U2142 ( .A(n5630), .Y(n4567) );
  INVX2 U2143 ( .A(n4880), .Y(n4662) );
  INVX2 U2144 ( .A(n5387), .Y(n4639) );
  INVX2 U2145 ( .A(n5477), .Y(n4637) );
  INVX2 U2146 ( .A(n5693), .Y(n4732) );
  AND2X1 U2147 ( .A(n4745), .B(n4977), .Y(n4559) );
  AND2X1 U2148 ( .A(n4744), .B(n5080), .Y(n4560) );
  INVX2 U2149 ( .A(n2135), .Y(n4660) );
  INVX2 U2150 ( .A(n2132), .Y(n4663) );
  INVX2 U2151 ( .A(n2138), .Y(n4655) );
  INVX2 U2152 ( .A(n2141), .Y(n4650) );
  INVX2 U2153 ( .A(n2144), .Y(n4645) );
  INVX2 U2154 ( .A(n2147), .Y(n4640) );
  INVX2 U2155 ( .A(n2147), .Y(n4641) );
  AND2X1 U2156 ( .A(n4741), .B(n5389), .Y(n4561) );
  AND2X1 U2157 ( .A(n4743), .B(n5183), .Y(n4562) );
  AND2X1 U2158 ( .A(n4740), .B(n5479), .Y(n4563) );
  AND2X1 U2159 ( .A(n4742), .B(n5286), .Y(n4564) );
  INVX2 U2160 ( .A(n2138), .Y(n4654) );
  INVX2 U2161 ( .A(n2141), .Y(n4649) );
  INVX2 U2162 ( .A(n2144), .Y(n4644) );
  INVX2 U2163 ( .A(n2135), .Y(n4659) );
  INVX2 U2164 ( .A(n5730), .Y(n4727) );
  INVX2 U2165 ( .A(n4565), .Y(n4667) );
  INVX2 U2166 ( .A(n4673), .Y(n4672) );
  INVX2 U2167 ( .A(n4675), .Y(n4674) );
  INVX2 U2168 ( .A(n4679), .Y(n4678) );
  INVX2 U2169 ( .A(n4677), .Y(n4676) );
  AND2X1 U2170 ( .A(a[1]), .B(n4748), .Y(n4565) );
  INVX2 U2171 ( .A(n4566), .Y(n4666) );
  INVX2 U2172 ( .A(n2159), .Y(n4673) );
  INVX2 U2173 ( .A(n2150), .Y(n4679) );
  AND2X1 U2174 ( .A(a[0]), .B(n4876), .Y(n4566) );
  INVX2 U2175 ( .A(n2153), .Y(n4677) );
  INVX2 U2176 ( .A(n2156), .Y(n4675) );
  INVX1 U2177 ( .A(b[3]), .Y(n4570) );
  INVX1 U2178 ( .A(b[19]), .Y(n4608) );
  INVX1 U2179 ( .A(b[24]), .Y(n4620) );
  INVX1 U2180 ( .A(b[25]), .Y(n4622) );
  INVX1 U2181 ( .A(b[1]), .Y(n4681) );
  INVX1 U2182 ( .A(b[16]), .Y(n4601) );
  INVX1 U2183 ( .A(b[23]), .Y(n4618) );
  INVX1 U2184 ( .A(b[7]), .Y(n4580) );
  INVX1 U2185 ( .A(b[13]), .Y(n4594) );
  INVX1 U2186 ( .A(b[31]), .Y(n4687) );
  INVX1 U2187 ( .A(b[17]), .Y(n4603) );
  INVX1 U2188 ( .A(b[15]), .Y(n4599) );
  INVX1 U2189 ( .A(b[27]), .Y(n4626) );
  INVX1 U2190 ( .A(b[21]), .Y(n4613) );
  INVX1 U2191 ( .A(b[29]), .Y(n4630) );
  INVX2 U2192 ( .A(n3301), .Y(n4688) );
  INVX2 U2193 ( .A(n3302), .Y(n4689) );
  INVX2 U2194 ( .A(n3303), .Y(n4690) );
  INVX2 U2195 ( .A(n5296), .Y(n4691) );
  INVX2 U2196 ( .A(n4785), .Y(n4692) );
  INVX2 U2197 ( .A(n3304), .Y(n4693) );
  INVX2 U2198 ( .A(n3305), .Y(n4694) );
  INVX2 U2199 ( .A(n3306), .Y(n4695) );
  INVX2 U2200 ( .A(n3307), .Y(n4696) );
  INVX2 U2201 ( .A(n3308), .Y(n4697) );
  INVX2 U2202 ( .A(n3309), .Y(n4698) );
  INVX2 U2203 ( .A(n3310), .Y(n4699) );
  INVX2 U2204 ( .A(n2429), .Y(n4709) );
  INVX2 U2205 ( .A(n2472), .Y(n4714) );
  INVX2 U2206 ( .A(n2520), .Y(n4718) );
  INVX2 U2207 ( .A(n5731), .Y(n4730) );
  INVX2 U2208 ( .A(n5694), .Y(n4734) );
  INVX2 U2209 ( .A(n5631), .Y(n4737) );
  INVX2 U2210 ( .A(n5561), .Y(n4738) );
  INVX2 U2211 ( .A(n5394), .Y(n4739) );
  INVX2 U2212 ( .A(n5478), .Y(n4740) );
  INVX2 U2213 ( .A(n5390), .Y(n4741) );
  INVX2 U2214 ( .A(n5287), .Y(n4742) );
  INVX2 U2215 ( .A(n5184), .Y(n4743) );
  INVX2 U2216 ( .A(n5081), .Y(n4744) );
  INVX2 U2217 ( .A(n4978), .Y(n4745) );
  INVX2 U2218 ( .A(n2132), .Y(n4746) );
  INVX2 U2219 ( .A(a[1]), .Y(n4747) );
  INVX2 U2220 ( .A(a[0]), .Y(n4748) );
  XOR2X1 U2221 ( .A(n4749), .B(n4750), .Y(product[47]) );
  XOR2X1 U2222 ( .A(n4751), .B(n4752), .Y(n4750) );
  XOR2X1 U2223 ( .A(n2405), .B(n2352), .Y(n4752) );
  XOR2X1 U2224 ( .A(n2409), .B(n2407), .Y(n4751) );
  XOR2X1 U2225 ( .A(n4753), .B(n4754), .Y(n4749) );
  XOR2X1 U2226 ( .A(n4676), .B(n4678), .Y(n4754) );
  XOR2X1 U2227 ( .A(n4755), .B(n4756), .Y(n4753) );
  XOR2X1 U2228 ( .A(n4757), .B(n4758), .Y(n4756) );
  XOR2X1 U2229 ( .A(n4759), .B(n4760), .Y(n4758) );
  XOR2X1 U2230 ( .A(n4761), .B(n4762), .Y(n4760) );
  XOR2X1 U2231 ( .A(n2411), .B(n2159), .Y(n4762) );
  XOR2X1 U2232 ( .A(n2415), .B(n2413), .Y(n4761) );
  XOR2X1 U2233 ( .A(n4763), .B(n4764), .Y(n4759) );
  XOR2X1 U2234 ( .A(n4765), .B(n4766), .Y(n4764) );
  OAI21X1 U2235 ( .A(n4558), .B(n4706), .C(n4767), .Y(n4766) );
  OAI22X1 U2236 ( .A(b[15]), .B(n4768), .C(n4727), .D(n4768), .Y(n4767) );
  OAI22X1 U2237 ( .A(n4728), .B(n4603), .C(n4729), .D(n4601), .Y(n4768) );
  OAI21X1 U2238 ( .A(n4557), .B(n4703), .C(n4769), .Y(n4765) );
  OAI22X1 U2239 ( .A(n4607), .B(n4770), .C(n4732), .D(n4770), .Y(n4769) );
  OAI22X1 U2240 ( .A(n4731), .B(n4611), .C(n4733), .D(n4608), .Y(n4770) );
  XOR2X1 U2241 ( .A(n4771), .B(n2156), .Y(n4763) );
  OAI21X1 U2242 ( .A(n4556), .B(n4700), .C(n4772), .Y(n4771) );
  OAI22X1 U2243 ( .A(n4615), .B(n4773), .C(n4567), .D(n4773), .Y(n4772) );
  OAI22X1 U2244 ( .A(n4735), .B(n4618), .C(n4736), .D(n4616), .Y(n4773) );
  OAI21X1 U2245 ( .A(n4555), .B(n4697), .C(n4774), .Y(n4757) );
  OAI22X1 U2246 ( .A(n4621), .B(n4775), .C(n4635), .D(n4775), .Y(n4774) );
  OAI22X1 U2247 ( .A(n4634), .B(n4624), .C(n4636), .D(n4622), .Y(n4775) );
  XOR2X1 U2248 ( .A(n4776), .B(n4777), .Y(n4755) );
  XNOR2X1 U2249 ( .A(n2147), .B(n4778), .Y(n4777) );
  OAI21X1 U2250 ( .A(n4664), .B(n4689), .C(n4779), .Y(n4778) );
  OAI22X1 U2251 ( .A(n4633), .B(n4780), .C(n4639), .D(n4780), .Y(n4779) );
  NOR2X1 U2252 ( .A(n4687), .B(n4552), .Y(n4780) );
  OAI21X1 U2253 ( .A(n4665), .B(n4694), .C(n4781), .Y(n4776) );
  OAI22X1 U2254 ( .A(n4627), .B(n4782), .C(n4637), .D(n4782), .Y(n4781) );
  OAI22X1 U2255 ( .A(n4739), .B(n4630), .C(n4638), .D(n4628), .Y(n4782) );
  XNOR2X1 U2256 ( .A(n4783), .B(n4663), .Y(n3661) );
  OAI22X1 U2257 ( .A(n4686), .B(n4553), .C(n4666), .D(n4686), .Y(n4783) );
  XNOR2X1 U2258 ( .A(n4784), .B(n4663), .Y(n3660) );
  OAI21X1 U2259 ( .A(n4666), .B(n4725), .C(n4692), .Y(n4784) );
  OAI22X1 U2260 ( .A(n4667), .B(n4686), .C(n4681), .D(n4553), .Y(n4785) );
  XNOR2X1 U2261 ( .A(n4786), .B(n4746), .Y(n3659) );
  OAI21X1 U2262 ( .A(n4666), .B(n4724), .C(n4787), .Y(n4786) );
  OAI22X1 U2263 ( .A(n4684), .B(n4788), .C(n4662), .D(n4788), .Y(n4787) );
  OAI22X1 U2264 ( .A(n4667), .B(n4681), .C(n4553), .D(n4568), .Y(n4788) );
  XNOR2X1 U2265 ( .A(n4789), .B(n4746), .Y(n3658) );
  OAI21X1 U2266 ( .A(n4666), .B(n4723), .C(n4790), .Y(n4789) );
  OAI22X1 U2267 ( .A(n4680), .B(n4791), .C(n4662), .D(n4791), .Y(n4790) );
  OAI22X1 U2268 ( .A(n4667), .B(n4568), .C(n4553), .D(n4570), .Y(n4791) );
  XNOR2X1 U2269 ( .A(n4792), .B(n4746), .Y(n3657) );
  OAI21X1 U2270 ( .A(n4666), .B(n4722), .C(n4793), .Y(n4792) );
  OAI22X1 U2271 ( .A(b[2]), .B(n4794), .C(n4662), .D(n4794), .Y(n4793) );
  OAI22X1 U2272 ( .A(n4667), .B(n4570), .C(n4553), .D(n4573), .Y(n4794) );
  XNOR2X1 U2273 ( .A(n4795), .B(n4746), .Y(n3656) );
  OAI21X1 U2274 ( .A(n4666), .B(n4721), .C(n4796), .Y(n4795) );
  OAI22X1 U2275 ( .A(n4572), .B(n4797), .C(n4662), .D(n4797), .Y(n4796) );
  OAI22X1 U2276 ( .A(n4667), .B(n4573), .C(n4553), .D(n4575), .Y(n4797) );
  XNOR2X1 U2277 ( .A(n4798), .B(n4746), .Y(n3655) );
  OAI21X1 U2278 ( .A(n4666), .B(n4720), .C(n4799), .Y(n4798) );
  OAI22X1 U2279 ( .A(b[4]), .B(n4800), .C(n4662), .D(n4800), .Y(n4799) );
  OAI22X1 U2280 ( .A(n4667), .B(n4575), .C(n4553), .D(n4578), .Y(n4800) );
  XNOR2X1 U2281 ( .A(n4801), .B(n4746), .Y(n3654) );
  OAI21X1 U2282 ( .A(n4666), .B(n4719), .C(n4802), .Y(n4801) );
  OAI22X1 U2283 ( .A(n4577), .B(n4803), .C(n4662), .D(n4803), .Y(n4802) );
  OAI22X1 U2284 ( .A(n4667), .B(n4578), .C(n4553), .D(n4580), .Y(n4803) );
  XNOR2X1 U2285 ( .A(n4804), .B(n4746), .Y(n3653) );
  OAI21X1 U2286 ( .A(n4666), .B(n4717), .C(n4805), .Y(n4804) );
  OAI22X1 U2287 ( .A(b[6]), .B(n4806), .C(n4662), .D(n4806), .Y(n4805) );
  OAI22X1 U2288 ( .A(n4667), .B(n4580), .C(n4553), .D(n4582), .Y(n4806) );
  XNOR2X1 U2289 ( .A(n4807), .B(n4746), .Y(n3652) );
  OAI21X1 U2290 ( .A(n4666), .B(n4716), .C(n4808), .Y(n4807) );
  OAI22X1 U2291 ( .A(b[7]), .B(n4809), .C(n4662), .D(n4809), .Y(n4808) );
  OAI22X1 U2292 ( .A(n4667), .B(n4582), .C(n4553), .D(n4584), .Y(n4809) );
  XNOR2X1 U2293 ( .A(n4810), .B(n4746), .Y(n3651) );
  OAI21X1 U2294 ( .A(n4666), .B(n4715), .C(n4811), .Y(n4810) );
  OAI22X1 U2295 ( .A(b[8]), .B(n4812), .C(n4662), .D(n4812), .Y(n4811) );
  OAI22X1 U2296 ( .A(n4667), .B(n4584), .C(n4553), .D(n4587), .Y(n4812) );
  XNOR2X1 U2297 ( .A(n4813), .B(n4746), .Y(n3650) );
  OAI21X1 U2298 ( .A(n4666), .B(n4713), .C(n4814), .Y(n4813) );
  OAI22X1 U2299 ( .A(n4586), .B(n4815), .C(n4662), .D(n4815), .Y(n4814) );
  OAI22X1 U2300 ( .A(n4667), .B(n4587), .C(n4553), .D(n4589), .Y(n4815) );
  XNOR2X1 U2301 ( .A(n4816), .B(n4746), .Y(n3649) );
  OAI21X1 U2302 ( .A(n4666), .B(n4712), .C(n4817), .Y(n4816) );
  OAI22X1 U2303 ( .A(b[10]), .B(n4818), .C(n4662), .D(n4818), .Y(n4817) );
  OAI22X1 U2304 ( .A(n4667), .B(n4589), .C(n4553), .D(n4592), .Y(n4818) );
  XNOR2X1 U2305 ( .A(n4819), .B(n4746), .Y(n3648) );
  OAI21X1 U2306 ( .A(n4666), .B(n4711), .C(n4820), .Y(n4819) );
  OAI22X1 U2307 ( .A(n4591), .B(n4821), .C(n4662), .D(n4821), .Y(n4820) );
  OAI22X1 U2308 ( .A(n4667), .B(n4592), .C(n4553), .D(n4594), .Y(n4821) );
  XNOR2X1 U2309 ( .A(n4822), .B(n4746), .Y(n3647) );
  OAI21X1 U2310 ( .A(n4666), .B(n4710), .C(n4823), .Y(n4822) );
  OAI22X1 U2311 ( .A(b[12]), .B(n4824), .C(n4662), .D(n4824), .Y(n4823) );
  OAI22X1 U2312 ( .A(n4667), .B(n4594), .C(n4553), .D(n4726), .Y(n4824) );
  XNOR2X1 U2313 ( .A(n4825), .B(n4746), .Y(n3646) );
  OAI21X1 U2314 ( .A(n4666), .B(n4708), .C(n4826), .Y(n4825) );
  OAI22X1 U2315 ( .A(n4596), .B(n4827), .C(n4662), .D(n4827), .Y(n4826) );
  OAI22X1 U2316 ( .A(n4667), .B(n4726), .C(n4553), .D(n4599), .Y(n4827) );
  XNOR2X1 U2317 ( .A(n4828), .B(n4746), .Y(n3645) );
  OAI21X1 U2318 ( .A(n4666), .B(n4707), .C(n4829), .Y(n4828) );
  OAI22X1 U2319 ( .A(b[14]), .B(n4830), .C(n4662), .D(n4830), .Y(n4829) );
  OAI22X1 U2320 ( .A(n4667), .B(n4599), .C(n4601), .D(n4553), .Y(n4830) );
  XNOR2X1 U2321 ( .A(n4831), .B(n4746), .Y(n3644) );
  OAI21X1 U2322 ( .A(n4706), .B(n4666), .C(n4832), .Y(n4831) );
  OAI22X1 U2323 ( .A(n4600), .B(n4833), .C(n4662), .D(n4833), .Y(n4832) );
  OAI22X1 U2324 ( .A(n4601), .B(n4667), .C(n4603), .D(n4553), .Y(n4833) );
  XNOR2X1 U2325 ( .A(n4834), .B(n4746), .Y(n3643) );
  OAI21X1 U2326 ( .A(n4666), .B(n4705), .C(n4835), .Y(n4834) );
  OAI22X1 U2327 ( .A(n4602), .B(n4836), .C(n4662), .D(n4836), .Y(n4835) );
  OAI22X1 U2328 ( .A(n4603), .B(n4667), .C(n4553), .D(n4606), .Y(n4836) );
  XNOR2X1 U2329 ( .A(n4837), .B(n4746), .Y(n3642) );
  OAI21X1 U2330 ( .A(n4666), .B(n4704), .C(n4838), .Y(n4837) );
  OAI22X1 U2331 ( .A(n4604), .B(n4839), .C(n4662), .D(n4839), .Y(n4838) );
  OAI22X1 U2332 ( .A(n4667), .B(n4606), .C(n4608), .D(n4553), .Y(n4839) );
  XNOR2X1 U2333 ( .A(n4840), .B(n4663), .Y(n3641) );
  OAI21X1 U2334 ( .A(n4703), .B(n4666), .C(n4841), .Y(n4840) );
  OAI22X1 U2335 ( .A(n4607), .B(n4842), .C(n4662), .D(n4842), .Y(n4841) );
  OAI22X1 U2336 ( .A(n4608), .B(n4667), .C(n4611), .D(n4553), .Y(n4842) );
  XNOR2X1 U2337 ( .A(n4843), .B(n4663), .Y(n3640) );
  OAI21X1 U2338 ( .A(n4666), .B(n4702), .C(n4844), .Y(n4843) );
  OAI22X1 U2339 ( .A(n4610), .B(n4845), .C(n4662), .D(n4845), .Y(n4844) );
  OAI22X1 U2340 ( .A(n4611), .B(n4667), .C(n4553), .D(n4613), .Y(n4845) );
  XNOR2X1 U2341 ( .A(n4846), .B(n4663), .Y(n3639) );
  OAI21X1 U2342 ( .A(n4666), .B(n4701), .C(n4847), .Y(n4846) );
  OAI22X1 U2343 ( .A(b[20]), .B(n4848), .C(n4662), .D(n4848), .Y(n4847) );
  OAI22X1 U2344 ( .A(n4667), .B(n4613), .C(n4616), .D(n4553), .Y(n4848) );
  XNOR2X1 U2345 ( .A(n4849), .B(n4663), .Y(n3638) );
  OAI21X1 U2346 ( .A(n4700), .B(n4666), .C(n4850), .Y(n4849) );
  OAI22X1 U2347 ( .A(n4614), .B(n4851), .C(n4662), .D(n4851), .Y(n4850) );
  OAI22X1 U2348 ( .A(n4616), .B(n4667), .C(n4618), .D(n4553), .Y(n4851) );
  XNOR2X1 U2349 ( .A(n4852), .B(n4663), .Y(n3637) );
  OAI21X1 U2350 ( .A(n4666), .B(n4699), .C(n4853), .Y(n4852) );
  OAI22X1 U2351 ( .A(n4617), .B(n4854), .C(n4662), .D(n4854), .Y(n4853) );
  OAI22X1 U2352 ( .A(n4618), .B(n4667), .C(n4553), .D(n4620), .Y(n4854) );
  XNOR2X1 U2353 ( .A(n4855), .B(n4663), .Y(n3636) );
  OAI21X1 U2354 ( .A(n4666), .B(n4698), .C(n4856), .Y(n4855) );
  OAI22X1 U2355 ( .A(n4619), .B(n4857), .C(n4662), .D(n4857), .Y(n4856) );
  OAI22X1 U2356 ( .A(n4667), .B(n4620), .C(n4622), .D(n4553), .Y(n4857) );
  XNOR2X1 U2357 ( .A(n4858), .B(n4663), .Y(n3635) );
  OAI21X1 U2358 ( .A(n4697), .B(n4666), .C(n4859), .Y(n4858) );
  OAI22X1 U2359 ( .A(n4621), .B(n4860), .C(n4662), .D(n4860), .Y(n4859) );
  OAI22X1 U2360 ( .A(n4622), .B(n4667), .C(n4624), .D(n4553), .Y(n4860) );
  XNOR2X1 U2361 ( .A(n4861), .B(n4663), .Y(n3634) );
  OAI21X1 U2362 ( .A(n4666), .B(n4696), .C(n4862), .Y(n4861) );
  OAI22X1 U2363 ( .A(n4623), .B(n4863), .C(n4662), .D(n4863), .Y(n4862) );
  OAI22X1 U2364 ( .A(n4624), .B(n4667), .C(n4553), .D(n4626), .Y(n4863) );
  XNOR2X1 U2365 ( .A(n4864), .B(n4663), .Y(n3633) );
  OAI21X1 U2366 ( .A(n4666), .B(n4695), .C(n4865), .Y(n4864) );
  OAI22X1 U2367 ( .A(n4625), .B(n4866), .C(n4662), .D(n4866), .Y(n4865) );
  OAI22X1 U2368 ( .A(n4667), .B(n4626), .C(n4628), .D(n4553), .Y(n4866) );
  XNOR2X1 U2369 ( .A(n4867), .B(n4663), .Y(n3632) );
  OAI21X1 U2370 ( .A(n4694), .B(n4666), .C(n4868), .Y(n4867) );
  OAI22X1 U2371 ( .A(n4627), .B(n4869), .C(n4662), .D(n4869), .Y(n4868) );
  OAI22X1 U2372 ( .A(n4628), .B(n4667), .C(n4630), .D(n4553), .Y(n4869) );
  XNOR2X1 U2373 ( .A(n4870), .B(n4663), .Y(n3631) );
  OAI21X1 U2374 ( .A(n4666), .B(n4693), .C(n4871), .Y(n4870) );
  OAI22X1 U2375 ( .A(n4629), .B(n4872), .C(n4662), .D(n4872), .Y(n4871) );
  OAI22X1 U2376 ( .A(n4630), .B(n4667), .C(n4553), .D(n4632), .Y(n4872) );
  XNOR2X1 U2377 ( .A(n4873), .B(n4663), .Y(n3630) );
  OAI21X1 U2378 ( .A(n4666), .B(n4690), .C(n4874), .Y(n4873) );
  OAI22X1 U2379 ( .A(n4631), .B(n4875), .C(n4662), .D(n4875), .Y(n4874) );
  OAI22X1 U2380 ( .A(n4667), .B(n4632), .C(n4687), .D(n4553), .Y(n4875) );
  XNOR2X1 U2381 ( .A(n4877), .B(n4663), .Y(n3629) );
  OAI21X1 U2382 ( .A(n4689), .B(n4666), .C(n4878), .Y(n4877) );
  OAI22X1 U2383 ( .A(n4633), .B(n4879), .C(n4662), .D(n4879), .Y(n4878) );
  NOR2X1 U2384 ( .A(n4667), .B(n4687), .Y(n4879) );
  XNOR2X1 U2385 ( .A(n4881), .B(n4663), .Y(n3628) );
  OAI22X1 U2386 ( .A(n4687), .B(n4880), .C(n4666), .D(n4688), .Y(n4881) );
  NAND3X1 U2387 ( .A(n4876), .B(n4748), .C(n4747), .Y(n4880) );
  XNOR2X1 U2388 ( .A(a[1]), .B(n4663), .Y(n4876) );
  XNOR2X1 U2389 ( .A(n4882), .B(n4659), .Y(n3626) );
  OAI22X1 U2390 ( .A(n4686), .B(n4658), .C(n4686), .D(n4668), .Y(n4882) );
  XNOR2X1 U2391 ( .A(n4883), .B(n4659), .Y(n3625) );
  OAI21X1 U2392 ( .A(n4725), .B(n4668), .C(n4884), .Y(n4883) );
  AOI22X1 U2393 ( .A(n4885), .B(n4684), .C(n4886), .D(n4680), .Y(n4884) );
  XNOR2X1 U2394 ( .A(n4887), .B(n4659), .Y(n3624) );
  OAI21X1 U2395 ( .A(n4724), .B(n4668), .C(n4888), .Y(n4887) );
  OAI22X1 U2396 ( .A(n4684), .B(n4889), .C(n4657), .D(n4889), .Y(n4888) );
  OAI22X1 U2397 ( .A(n4681), .B(n4661), .C(n4568), .D(n4658), .Y(n4889) );
  XNOR2X1 U2398 ( .A(n4890), .B(n4659), .Y(n3623) );
  OAI21X1 U2399 ( .A(n4723), .B(n4668), .C(n4891), .Y(n4890) );
  OAI22X1 U2400 ( .A(n4680), .B(n4892), .C(n4657), .D(n4892), .Y(n4891) );
  OAI22X1 U2401 ( .A(n4568), .B(n4661), .C(n4570), .D(n4658), .Y(n4892) );
  XNOR2X1 U2402 ( .A(n4893), .B(n4659), .Y(n3622) );
  OAI21X1 U2403 ( .A(n4722), .B(n4668), .C(n4894), .Y(n4893) );
  OAI22X1 U2404 ( .A(n4569), .B(n4895), .C(n4657), .D(n4895), .Y(n4894) );
  OAI22X1 U2405 ( .A(n4570), .B(n4661), .C(n4573), .D(n4658), .Y(n4895) );
  XNOR2X1 U2406 ( .A(n4896), .B(n4659), .Y(n3621) );
  OAI21X1 U2407 ( .A(n4721), .B(n4668), .C(n4897), .Y(n4896) );
  OAI22X1 U2408 ( .A(n4571), .B(n4898), .C(n4657), .D(n4898), .Y(n4897) );
  OAI22X1 U2409 ( .A(n4573), .B(n4661), .C(n4575), .D(n4658), .Y(n4898) );
  XNOR2X1 U2410 ( .A(n4899), .B(n4659), .Y(n3620) );
  OAI21X1 U2411 ( .A(n4720), .B(n4668), .C(n4900), .Y(n4899) );
  OAI22X1 U2412 ( .A(n4574), .B(n4901), .C(n4657), .D(n4901), .Y(n4900) );
  OAI22X1 U2413 ( .A(n4575), .B(n4661), .C(n4578), .D(n4658), .Y(n4901) );
  XNOR2X1 U2414 ( .A(n4902), .B(n4659), .Y(n3619) );
  OAI21X1 U2415 ( .A(n4719), .B(n4668), .C(n4903), .Y(n4902) );
  OAI22X1 U2416 ( .A(n4576), .B(n4904), .C(n4657), .D(n4904), .Y(n4903) );
  OAI22X1 U2417 ( .A(n4578), .B(n4661), .C(n4580), .D(n4658), .Y(n4904) );
  XNOR2X1 U2418 ( .A(n4905), .B(n4659), .Y(n3618) );
  OAI21X1 U2419 ( .A(n4717), .B(n4668), .C(n4906), .Y(n4905) );
  OAI22X1 U2420 ( .A(n4579), .B(n4907), .C(n4657), .D(n4907), .Y(n4906) );
  OAI22X1 U2421 ( .A(n4580), .B(n4661), .C(n4582), .D(n4658), .Y(n4907) );
  XNOR2X1 U2422 ( .A(n4908), .B(n4659), .Y(n3617) );
  OAI21X1 U2423 ( .A(n4716), .B(n4668), .C(n4909), .Y(n4908) );
  OAI22X1 U2424 ( .A(n4581), .B(n4910), .C(n4657), .D(n4910), .Y(n4909) );
  OAI22X1 U2425 ( .A(n4582), .B(n4661), .C(n4584), .D(n4658), .Y(n4910) );
  XNOR2X1 U2426 ( .A(n4911), .B(n4659), .Y(n3616) );
  OAI21X1 U2427 ( .A(n4715), .B(n4668), .C(n4912), .Y(n4911) );
  OAI22X1 U2428 ( .A(n4583), .B(n4913), .C(n4657), .D(n4913), .Y(n4912) );
  OAI22X1 U2429 ( .A(n4584), .B(n4661), .C(n4587), .D(n4658), .Y(n4913) );
  XNOR2X1 U2430 ( .A(n4914), .B(n4659), .Y(n3615) );
  OAI21X1 U2431 ( .A(n4713), .B(n4668), .C(n4915), .Y(n4914) );
  OAI22X1 U2432 ( .A(n4585), .B(n4916), .C(n4657), .D(n4916), .Y(n4915) );
  OAI22X1 U2433 ( .A(n4587), .B(n4661), .C(n4589), .D(n4658), .Y(n4916) );
  XNOR2X1 U2434 ( .A(n4917), .B(n4659), .Y(n3614) );
  OAI21X1 U2435 ( .A(n4712), .B(n4668), .C(n4918), .Y(n4917) );
  OAI22X1 U2436 ( .A(n4588), .B(n4919), .C(n4657), .D(n4919), .Y(n4918) );
  OAI22X1 U2437 ( .A(n4589), .B(n4661), .C(n4592), .D(n4658), .Y(n4919) );
  XNOR2X1 U2438 ( .A(n4920), .B(n4659), .Y(n3613) );
  OAI21X1 U2439 ( .A(n4711), .B(n4668), .C(n4921), .Y(n4920) );
  OAI22X1 U2440 ( .A(n4590), .B(n4922), .C(n4657), .D(n4922), .Y(n4921) );
  OAI22X1 U2441 ( .A(n4592), .B(n4661), .C(n4594), .D(n4658), .Y(n4922) );
  XNOR2X1 U2442 ( .A(n4923), .B(n4659), .Y(n3612) );
  OAI21X1 U2443 ( .A(n4710), .B(n4668), .C(n4924), .Y(n4923) );
  OAI22X1 U2444 ( .A(n4593), .B(n4925), .C(n4657), .D(n4925), .Y(n4924) );
  OAI22X1 U2445 ( .A(n4594), .B(n4661), .C(n4726), .D(n4658), .Y(n4925) );
  XNOR2X1 U2446 ( .A(n4926), .B(n4659), .Y(n3611) );
  OAI21X1 U2447 ( .A(n4708), .B(n4668), .C(n4927), .Y(n4926) );
  OAI22X1 U2448 ( .A(n4595), .B(n4928), .C(n4657), .D(n4928), .Y(n4927) );
  OAI22X1 U2449 ( .A(n4726), .B(n4661), .C(n4599), .D(n4658), .Y(n4928) );
  XNOR2X1 U2450 ( .A(n4929), .B(n4659), .Y(n3610) );
  OAI21X1 U2451 ( .A(n4707), .B(n4668), .C(n4930), .Y(n4929) );
  OAI22X1 U2452 ( .A(n4598), .B(n4931), .C(n4657), .D(n4931), .Y(n4930) );
  OAI22X1 U2453 ( .A(n4599), .B(n4661), .C(n4601), .D(n4658), .Y(n4931) );
  XNOR2X1 U2454 ( .A(n4932), .B(n4659), .Y(n3609) );
  OAI21X1 U2455 ( .A(n4706), .B(n4668), .C(n4933), .Y(n4932) );
  OAI22X1 U2456 ( .A(b[15]), .B(n4934), .C(n4657), .D(n4934), .Y(n4933) );
  OAI22X1 U2457 ( .A(n4601), .B(n4661), .C(n4603), .D(n4658), .Y(n4934) );
  XNOR2X1 U2458 ( .A(n4935), .B(n4659), .Y(n3608) );
  OAI21X1 U2459 ( .A(n4705), .B(n4668), .C(n4936), .Y(n4935) );
  OAI22X1 U2460 ( .A(n4602), .B(n4937), .C(n4657), .D(n4937), .Y(n4936) );
  OAI22X1 U2461 ( .A(n4603), .B(n4661), .C(n4606), .D(n4658), .Y(n4937) );
  XNOR2X1 U2462 ( .A(n4938), .B(n4660), .Y(n3607) );
  OAI21X1 U2463 ( .A(n4704), .B(n4668), .C(n4939), .Y(n4938) );
  OAI22X1 U2464 ( .A(n4605), .B(n4940), .C(n4657), .D(n4940), .Y(n4939) );
  OAI22X1 U2465 ( .A(n4606), .B(n4661), .C(n4608), .D(n4658), .Y(n4940) );
  XNOR2X1 U2466 ( .A(n4941), .B(n4660), .Y(n3606) );
  OAI21X1 U2467 ( .A(n4703), .B(n4668), .C(n4942), .Y(n4941) );
  OAI22X1 U2468 ( .A(n4607), .B(n4943), .C(n4657), .D(n4943), .Y(n4942) );
  OAI22X1 U2469 ( .A(n4608), .B(n4661), .C(n4611), .D(n4658), .Y(n4943) );
  XNOR2X1 U2470 ( .A(n4944), .B(n4660), .Y(n3605) );
  OAI21X1 U2471 ( .A(n4702), .B(n4668), .C(n4945), .Y(n4944) );
  OAI22X1 U2472 ( .A(n4609), .B(n4946), .C(n4657), .D(n4946), .Y(n4945) );
  OAI22X1 U2473 ( .A(n4611), .B(n4661), .C(n4613), .D(n4658), .Y(n4946) );
  XNOR2X1 U2474 ( .A(n4947), .B(n4660), .Y(n3604) );
  OAI21X1 U2475 ( .A(n4701), .B(n4668), .C(n4948), .Y(n4947) );
  OAI22X1 U2476 ( .A(n4612), .B(n4949), .C(n4657), .D(n4949), .Y(n4948) );
  OAI22X1 U2477 ( .A(n4613), .B(n4661), .C(n4616), .D(n4658), .Y(n4949) );
  XNOR2X1 U2478 ( .A(n4950), .B(n4660), .Y(n3603) );
  OAI21X1 U2479 ( .A(n4700), .B(n4668), .C(n4951), .Y(n4950) );
  OAI22X1 U2480 ( .A(n4615), .B(n4952), .C(n4657), .D(n4952), .Y(n4951) );
  OAI22X1 U2481 ( .A(n4616), .B(n4661), .C(n4618), .D(n4658), .Y(n4952) );
  XNOR2X1 U2482 ( .A(n4953), .B(n4660), .Y(n3602) );
  OAI21X1 U2483 ( .A(n4699), .B(n4668), .C(n4954), .Y(n4953) );
  OAI22X1 U2484 ( .A(n4617), .B(n4955), .C(n4657), .D(n4955), .Y(n4954) );
  OAI22X1 U2485 ( .A(n4618), .B(n4661), .C(n4620), .D(n4658), .Y(n4955) );
  XNOR2X1 U2486 ( .A(n4956), .B(n4660), .Y(n3601) );
  OAI21X1 U2487 ( .A(n4698), .B(n4668), .C(n4957), .Y(n4956) );
  OAI22X1 U2488 ( .A(n4619), .B(n4958), .C(n4657), .D(n4958), .Y(n4957) );
  OAI22X1 U2489 ( .A(n4620), .B(n4661), .C(n4622), .D(n4658), .Y(n4958) );
  XNOR2X1 U2490 ( .A(n4959), .B(n4660), .Y(n3600) );
  OAI21X1 U2491 ( .A(n4697), .B(n4668), .C(n4960), .Y(n4959) );
  OAI22X1 U2492 ( .A(n4621), .B(n4961), .C(n4657), .D(n4961), .Y(n4960) );
  OAI22X1 U2493 ( .A(n4622), .B(n4661), .C(n4624), .D(n4658), .Y(n4961) );
  XNOR2X1 U2494 ( .A(n4962), .B(n4660), .Y(n3599) );
  OAI21X1 U2495 ( .A(n4696), .B(n4668), .C(n4963), .Y(n4962) );
  OAI22X1 U2496 ( .A(n4623), .B(n4964), .C(n4657), .D(n4964), .Y(n4963) );
  OAI22X1 U2497 ( .A(n4624), .B(n4661), .C(n4626), .D(n4658), .Y(n4964) );
  XNOR2X1 U2498 ( .A(n4965), .B(n4660), .Y(n3598) );
  OAI21X1 U2499 ( .A(n4695), .B(n4668), .C(n4966), .Y(n4965) );
  OAI22X1 U2500 ( .A(n4625), .B(n4967), .C(n4657), .D(n4967), .Y(n4966) );
  OAI22X1 U2501 ( .A(n4626), .B(n4661), .C(n4628), .D(n4658), .Y(n4967) );
  XNOR2X1 U2502 ( .A(n4968), .B(n4660), .Y(n3597) );
  OAI21X1 U2503 ( .A(n4694), .B(n4668), .C(n4969), .Y(n4968) );
  OAI22X1 U2504 ( .A(n4627), .B(n4970), .C(n4657), .D(n4970), .Y(n4969) );
  OAI22X1 U2505 ( .A(n4628), .B(n4661), .C(n4630), .D(n4658), .Y(n4970) );
  XNOR2X1 U2506 ( .A(n4971), .B(n4660), .Y(n3596) );
  OAI21X1 U2507 ( .A(n4693), .B(n4668), .C(n4972), .Y(n4971) );
  OAI22X1 U2508 ( .A(n4629), .B(n4973), .C(n4657), .D(n4973), .Y(n4972) );
  OAI22X1 U2509 ( .A(n4630), .B(n4661), .C(n4632), .D(n4658), .Y(n4973) );
  XNOR2X1 U2510 ( .A(n4974), .B(n4660), .Y(n3595) );
  OAI21X1 U2511 ( .A(n4690), .B(n4668), .C(n4975), .Y(n4974) );
  OAI22X1 U2512 ( .A(n4631), .B(n4976), .C(n4657), .D(n4976), .Y(n4975) );
  OAI22X1 U2513 ( .A(n4632), .B(n4661), .C(n4687), .D(n4658), .Y(n4976) );
  NOR2X1 U2514 ( .A(n4977), .B(n4978), .Y(n4886) );
  XNOR2X1 U2515 ( .A(n4979), .B(n4660), .Y(n3594) );
  OAI21X1 U2516 ( .A(n4689), .B(n4668), .C(n4980), .Y(n4979) );
  OAI22X1 U2517 ( .A(n4633), .B(n4981), .C(n4657), .D(n4981), .Y(n4980) );
  NOR2X1 U2518 ( .A(n4661), .B(n4687), .Y(n4981) );
  NOR2X1 U2519 ( .A(n4745), .B(n4983), .Y(n4885) );
  XNOR2X1 U2520 ( .A(n4984), .B(n4660), .Y(n3593) );
  OAI22X1 U2521 ( .A(n4687), .B(n4982), .C(n4688), .D(n4668), .Y(n4984) );
  NAND3X1 U2522 ( .A(n4978), .B(n4977), .C(n4983), .Y(n4982) );
  XNOR2X1 U2523 ( .A(a[3]), .B(a[4]), .Y(n4983) );
  XNOR2X1 U2524 ( .A(a[4]), .B(n4660), .Y(n4977) );
  XOR2X1 U2525 ( .A(a[3]), .B(n4663), .Y(n4978) );
  XNOR2X1 U2526 ( .A(n4985), .B(n4654), .Y(n3591) );
  OAI22X1 U2527 ( .A(n4686), .B(n4653), .C(n4686), .D(n4669), .Y(n4985) );
  XNOR2X1 U2528 ( .A(n4986), .B(n4654), .Y(n3590) );
  OAI21X1 U2529 ( .A(n4725), .B(n4669), .C(n4987), .Y(n4986) );
  AOI22X1 U2530 ( .A(n4988), .B(n4684), .C(n4989), .D(n4680), .Y(n4987) );
  XNOR2X1 U2531 ( .A(n4990), .B(n4654), .Y(n3589) );
  OAI21X1 U2532 ( .A(n4724), .B(n4669), .C(n4991), .Y(n4990) );
  OAI22X1 U2533 ( .A(n4684), .B(n4992), .C(n4652), .D(n4992), .Y(n4991) );
  OAI22X1 U2534 ( .A(n4681), .B(n4656), .C(n4568), .D(n4653), .Y(n4992) );
  XNOR2X1 U2535 ( .A(n4993), .B(n4654), .Y(n3588) );
  OAI21X1 U2536 ( .A(n4723), .B(n4669), .C(n4994), .Y(n4993) );
  OAI22X1 U2537 ( .A(n4680), .B(n4995), .C(n4652), .D(n4995), .Y(n4994) );
  OAI22X1 U2538 ( .A(n4568), .B(n4656), .C(n4570), .D(n4653), .Y(n4995) );
  XNOR2X1 U2539 ( .A(n4996), .B(n4654), .Y(n3587) );
  OAI21X1 U2540 ( .A(n4722), .B(n4669), .C(n4997), .Y(n4996) );
  OAI22X1 U2541 ( .A(b[2]), .B(n4998), .C(n4652), .D(n4998), .Y(n4997) );
  OAI22X1 U2542 ( .A(n4570), .B(n4656), .C(n4573), .D(n4653), .Y(n4998) );
  XNOR2X1 U2543 ( .A(n4999), .B(n4654), .Y(n3586) );
  OAI21X1 U2544 ( .A(n4721), .B(n4669), .C(n5000), .Y(n4999) );
  OAI22X1 U2545 ( .A(n4572), .B(n5001), .C(n4652), .D(n5001), .Y(n5000) );
  OAI22X1 U2546 ( .A(n4573), .B(n4656), .C(n4575), .D(n4653), .Y(n5001) );
  XNOR2X1 U2547 ( .A(n5002), .B(n4654), .Y(n3585) );
  OAI21X1 U2548 ( .A(n4720), .B(n4669), .C(n5003), .Y(n5002) );
  OAI22X1 U2549 ( .A(b[4]), .B(n5004), .C(n4652), .D(n5004), .Y(n5003) );
  OAI22X1 U2550 ( .A(n4575), .B(n4656), .C(n4578), .D(n4653), .Y(n5004) );
  XNOR2X1 U2551 ( .A(n5005), .B(n4654), .Y(n3584) );
  OAI21X1 U2552 ( .A(n4719), .B(n4669), .C(n5006), .Y(n5005) );
  OAI22X1 U2553 ( .A(n4577), .B(n5007), .C(n4652), .D(n5007), .Y(n5006) );
  OAI22X1 U2554 ( .A(n4578), .B(n4656), .C(n4580), .D(n4653), .Y(n5007) );
  XNOR2X1 U2555 ( .A(n5008), .B(n4654), .Y(n3583) );
  OAI21X1 U2556 ( .A(n4717), .B(n4669), .C(n5009), .Y(n5008) );
  OAI22X1 U2557 ( .A(b[6]), .B(n5010), .C(n4652), .D(n5010), .Y(n5009) );
  OAI22X1 U2558 ( .A(n4580), .B(n4656), .C(n4582), .D(n4653), .Y(n5010) );
  XNOR2X1 U2559 ( .A(n5011), .B(n4654), .Y(n3582) );
  OAI21X1 U2560 ( .A(n4716), .B(n4669), .C(n5012), .Y(n5011) );
  OAI22X1 U2561 ( .A(b[7]), .B(n5013), .C(n4652), .D(n5013), .Y(n5012) );
  OAI22X1 U2562 ( .A(n4582), .B(n4656), .C(n4584), .D(n4653), .Y(n5013) );
  XNOR2X1 U2563 ( .A(n5014), .B(n4654), .Y(n3581) );
  OAI21X1 U2564 ( .A(n4715), .B(n4669), .C(n5015), .Y(n5014) );
  OAI22X1 U2565 ( .A(b[8]), .B(n5016), .C(n4652), .D(n5016), .Y(n5015) );
  OAI22X1 U2566 ( .A(n4584), .B(n4656), .C(n4587), .D(n4653), .Y(n5016) );
  XNOR2X1 U2567 ( .A(n5017), .B(n4654), .Y(n3580) );
  OAI21X1 U2568 ( .A(n4713), .B(n4669), .C(n5018), .Y(n5017) );
  OAI22X1 U2569 ( .A(n4586), .B(n5019), .C(n4652), .D(n5019), .Y(n5018) );
  OAI22X1 U2570 ( .A(n4587), .B(n4656), .C(n4589), .D(n4653), .Y(n5019) );
  XNOR2X1 U2571 ( .A(n5020), .B(n4654), .Y(n3579) );
  OAI21X1 U2572 ( .A(n4712), .B(n4669), .C(n5021), .Y(n5020) );
  OAI22X1 U2573 ( .A(b[10]), .B(n5022), .C(n4652), .D(n5022), .Y(n5021) );
  OAI22X1 U2574 ( .A(n4589), .B(n4656), .C(n4592), .D(n4653), .Y(n5022) );
  XNOR2X1 U2575 ( .A(n5023), .B(n4654), .Y(n3578) );
  OAI21X1 U2576 ( .A(n4711), .B(n4669), .C(n5024), .Y(n5023) );
  OAI22X1 U2577 ( .A(n4591), .B(n5025), .C(n4652), .D(n5025), .Y(n5024) );
  OAI22X1 U2578 ( .A(n4592), .B(n4656), .C(n4594), .D(n4653), .Y(n5025) );
  XNOR2X1 U2579 ( .A(n5026), .B(n4654), .Y(n3577) );
  OAI21X1 U2580 ( .A(n4710), .B(n4669), .C(n5027), .Y(n5026) );
  OAI22X1 U2581 ( .A(b[12]), .B(n5028), .C(n4652), .D(n5028), .Y(n5027) );
  OAI22X1 U2582 ( .A(n4594), .B(n4656), .C(n4726), .D(n4653), .Y(n5028) );
  XNOR2X1 U2583 ( .A(n5029), .B(n4654), .Y(n3576) );
  OAI21X1 U2584 ( .A(n4708), .B(n4669), .C(n5030), .Y(n5029) );
  OAI22X1 U2585 ( .A(n4596), .B(n5031), .C(n4652), .D(n5031), .Y(n5030) );
  OAI22X1 U2586 ( .A(n4726), .B(n4656), .C(n4599), .D(n4653), .Y(n5031) );
  XNOR2X1 U2587 ( .A(n5032), .B(n4654), .Y(n3575) );
  OAI21X1 U2588 ( .A(n4707), .B(n4669), .C(n5033), .Y(n5032) );
  OAI22X1 U2589 ( .A(b[14]), .B(n5034), .C(n4652), .D(n5034), .Y(n5033) );
  OAI22X1 U2590 ( .A(n4599), .B(n4656), .C(n4601), .D(n4653), .Y(n5034) );
  XNOR2X1 U2591 ( .A(n5035), .B(n4654), .Y(n3574) );
  OAI21X1 U2592 ( .A(n4706), .B(n4669), .C(n5036), .Y(n5035) );
  OAI22X1 U2593 ( .A(n4600), .B(n5037), .C(n4652), .D(n5037), .Y(n5036) );
  OAI22X1 U2594 ( .A(n4601), .B(n4656), .C(n4603), .D(n4653), .Y(n5037) );
  XNOR2X1 U2595 ( .A(n5038), .B(n4654), .Y(n3573) );
  OAI21X1 U2596 ( .A(n4705), .B(n4669), .C(n5039), .Y(n5038) );
  OAI22X1 U2597 ( .A(n4602), .B(n5040), .C(n4652), .D(n5040), .Y(n5039) );
  OAI22X1 U2598 ( .A(n4603), .B(n4656), .C(n4606), .D(n4653), .Y(n5040) );
  XNOR2X1 U2599 ( .A(n5041), .B(n4654), .Y(n3572) );
  OAI21X1 U2600 ( .A(n4704), .B(n4669), .C(n5042), .Y(n5041) );
  OAI22X1 U2601 ( .A(n4605), .B(n5043), .C(n4652), .D(n5043), .Y(n5042) );
  OAI22X1 U2602 ( .A(n4606), .B(n4656), .C(n4608), .D(n4653), .Y(n5043) );
  XNOR2X1 U2603 ( .A(n5044), .B(n4655), .Y(n3571) );
  OAI21X1 U2604 ( .A(n4703), .B(n4669), .C(n5045), .Y(n5044) );
  OAI22X1 U2605 ( .A(n4607), .B(n5046), .C(n4652), .D(n5046), .Y(n5045) );
  OAI22X1 U2606 ( .A(n4608), .B(n4656), .C(n4611), .D(n4653), .Y(n5046) );
  XNOR2X1 U2607 ( .A(n5047), .B(n4655), .Y(n3570) );
  OAI21X1 U2608 ( .A(n4702), .B(n4669), .C(n5048), .Y(n5047) );
  OAI22X1 U2609 ( .A(n4610), .B(n5049), .C(n4652), .D(n5049), .Y(n5048) );
  OAI22X1 U2610 ( .A(n4611), .B(n4656), .C(n4613), .D(n4653), .Y(n5049) );
  XNOR2X1 U2611 ( .A(n5050), .B(n4655), .Y(n3569) );
  OAI21X1 U2612 ( .A(n4701), .B(n4669), .C(n5051), .Y(n5050) );
  OAI22X1 U2613 ( .A(b[20]), .B(n5052), .C(n4652), .D(n5052), .Y(n5051) );
  OAI22X1 U2614 ( .A(n4613), .B(n4656), .C(n4616), .D(n4653), .Y(n5052) );
  XNOR2X1 U2615 ( .A(n5053), .B(n4655), .Y(n3568) );
  OAI21X1 U2616 ( .A(n4700), .B(n4669), .C(n5054), .Y(n5053) );
  OAI22X1 U2617 ( .A(n4614), .B(n5055), .C(n4652), .D(n5055), .Y(n5054) );
  OAI22X1 U2618 ( .A(n4616), .B(n4656), .C(n4618), .D(n4653), .Y(n5055) );
  XNOR2X1 U2619 ( .A(n5056), .B(n4655), .Y(n3567) );
  OAI21X1 U2620 ( .A(n4699), .B(n4669), .C(n5057), .Y(n5056) );
  OAI22X1 U2621 ( .A(n4617), .B(n5058), .C(n4652), .D(n5058), .Y(n5057) );
  OAI22X1 U2622 ( .A(n4618), .B(n4656), .C(n4620), .D(n4653), .Y(n5058) );
  XNOR2X1 U2623 ( .A(n5059), .B(n4655), .Y(n3566) );
  OAI21X1 U2624 ( .A(n4698), .B(n4669), .C(n5060), .Y(n5059) );
  OAI22X1 U2625 ( .A(n4619), .B(n5061), .C(n4652), .D(n5061), .Y(n5060) );
  OAI22X1 U2626 ( .A(n4620), .B(n4656), .C(n4622), .D(n4653), .Y(n5061) );
  XNOR2X1 U2627 ( .A(n5062), .B(n4655), .Y(n3565) );
  OAI21X1 U2628 ( .A(n4697), .B(n4669), .C(n5063), .Y(n5062) );
  OAI22X1 U2629 ( .A(n4621), .B(n5064), .C(n4652), .D(n5064), .Y(n5063) );
  OAI22X1 U2630 ( .A(n4622), .B(n4656), .C(n4624), .D(n4653), .Y(n5064) );
  XNOR2X1 U2631 ( .A(n5065), .B(n4655), .Y(n3564) );
  OAI21X1 U2632 ( .A(n4696), .B(n4669), .C(n5066), .Y(n5065) );
  OAI22X1 U2633 ( .A(n4623), .B(n5067), .C(n4652), .D(n5067), .Y(n5066) );
  OAI22X1 U2634 ( .A(n4624), .B(n4656), .C(n4626), .D(n4653), .Y(n5067) );
  XNOR2X1 U2635 ( .A(n5068), .B(n4655), .Y(n3563) );
  OAI21X1 U2636 ( .A(n4695), .B(n4669), .C(n5069), .Y(n5068) );
  OAI22X1 U2637 ( .A(n4625), .B(n5070), .C(n4652), .D(n5070), .Y(n5069) );
  OAI22X1 U2638 ( .A(n4626), .B(n4656), .C(n4628), .D(n4653), .Y(n5070) );
  XNOR2X1 U2639 ( .A(n5071), .B(n4655), .Y(n3562) );
  OAI21X1 U2640 ( .A(n4694), .B(n4669), .C(n5072), .Y(n5071) );
  OAI22X1 U2641 ( .A(n4627), .B(n5073), .C(n4652), .D(n5073), .Y(n5072) );
  OAI22X1 U2642 ( .A(n4628), .B(n4656), .C(n4630), .D(n4653), .Y(n5073) );
  XNOR2X1 U2643 ( .A(n5074), .B(n4655), .Y(n3561) );
  OAI21X1 U2644 ( .A(n4693), .B(n4669), .C(n5075), .Y(n5074) );
  OAI22X1 U2645 ( .A(n4629), .B(n5076), .C(n4652), .D(n5076), .Y(n5075) );
  OAI22X1 U2646 ( .A(n4630), .B(n4656), .C(n4632), .D(n4653), .Y(n5076) );
  XNOR2X1 U2647 ( .A(n5077), .B(n4655), .Y(n3560) );
  OAI21X1 U2648 ( .A(n4690), .B(n4669), .C(n5078), .Y(n5077) );
  OAI22X1 U2649 ( .A(n4631), .B(n5079), .C(n4652), .D(n5079), .Y(n5078) );
  OAI22X1 U2650 ( .A(n4632), .B(n4656), .C(n4687), .D(n4653), .Y(n5079) );
  NOR2X1 U2651 ( .A(n5080), .B(n5081), .Y(n4989) );
  XNOR2X1 U2652 ( .A(n5082), .B(n4655), .Y(n3559) );
  OAI21X1 U2653 ( .A(n4689), .B(n4669), .C(n5083), .Y(n5082) );
  OAI22X1 U2654 ( .A(n4633), .B(n5084), .C(n4652), .D(n5084), .Y(n5083) );
  NOR2X1 U2655 ( .A(n4656), .B(n4687), .Y(n5084) );
  NOR2X1 U2656 ( .A(n4744), .B(n5086), .Y(n4988) );
  XNOR2X1 U2657 ( .A(n5087), .B(n4655), .Y(n3558) );
  OAI22X1 U2658 ( .A(n4687), .B(n5085), .C(n4688), .D(n4669), .Y(n5087) );
  NAND3X1 U2659 ( .A(n5081), .B(n5080), .C(n5086), .Y(n5085) );
  XNOR2X1 U2660 ( .A(a[6]), .B(a[7]), .Y(n5086) );
  XNOR2X1 U2661 ( .A(a[7]), .B(n4655), .Y(n5080) );
  XOR2X1 U2662 ( .A(a[6]), .B(n4660), .Y(n5081) );
  XNOR2X1 U2663 ( .A(n5088), .B(n4649), .Y(n3556) );
  OAI22X1 U2664 ( .A(n4686), .B(n4648), .C(n4686), .D(n4670), .Y(n5088) );
  XNOR2X1 U2665 ( .A(n5089), .B(n4649), .Y(n3555) );
  OAI21X1 U2666 ( .A(n4725), .B(n4670), .C(n5090), .Y(n5089) );
  AOI22X1 U2667 ( .A(n5091), .B(n4684), .C(n5092), .D(n4680), .Y(n5090) );
  XNOR2X1 U2668 ( .A(n5093), .B(n4649), .Y(n3554) );
  OAI21X1 U2669 ( .A(n4724), .B(n4670), .C(n5094), .Y(n5093) );
  OAI22X1 U2670 ( .A(n4685), .B(n5095), .C(n4647), .D(n5095), .Y(n5094) );
  OAI22X1 U2671 ( .A(n4681), .B(n4651), .C(n4568), .D(n4648), .Y(n5095) );
  XNOR2X1 U2672 ( .A(n5096), .B(n4649), .Y(n3553) );
  OAI21X1 U2673 ( .A(n4723), .B(n4670), .C(n5097), .Y(n5096) );
  OAI22X1 U2674 ( .A(n4680), .B(n5098), .C(n4647), .D(n5098), .Y(n5097) );
  OAI22X1 U2675 ( .A(n4568), .B(n4651), .C(n4570), .D(n4648), .Y(n5098) );
  XNOR2X1 U2676 ( .A(n5099), .B(n4649), .Y(n3552) );
  OAI21X1 U2677 ( .A(n4722), .B(n4670), .C(n5100), .Y(n5099) );
  OAI22X1 U2678 ( .A(n4569), .B(n5101), .C(n4647), .D(n5101), .Y(n5100) );
  OAI22X1 U2679 ( .A(n4570), .B(n4651), .C(n4573), .D(n4648), .Y(n5101) );
  XNOR2X1 U2680 ( .A(n5102), .B(n4649), .Y(n3551) );
  OAI21X1 U2681 ( .A(n4721), .B(n4670), .C(n5103), .Y(n5102) );
  OAI22X1 U2682 ( .A(n4571), .B(n5104), .C(n4647), .D(n5104), .Y(n5103) );
  OAI22X1 U2683 ( .A(n4573), .B(n4651), .C(n4575), .D(n4648), .Y(n5104) );
  XNOR2X1 U2684 ( .A(n5105), .B(n4649), .Y(n3550) );
  OAI21X1 U2685 ( .A(n4720), .B(n4670), .C(n5106), .Y(n5105) );
  OAI22X1 U2686 ( .A(n4574), .B(n5107), .C(n4647), .D(n5107), .Y(n5106) );
  OAI22X1 U2687 ( .A(n4575), .B(n4651), .C(n4578), .D(n4648), .Y(n5107) );
  XNOR2X1 U2688 ( .A(n5108), .B(n4649), .Y(n3549) );
  OAI21X1 U2689 ( .A(n4719), .B(n4670), .C(n5109), .Y(n5108) );
  OAI22X1 U2690 ( .A(n4576), .B(n5110), .C(n4647), .D(n5110), .Y(n5109) );
  OAI22X1 U2691 ( .A(n4578), .B(n4651), .C(n4580), .D(n4648), .Y(n5110) );
  XNOR2X1 U2692 ( .A(n5111), .B(n4649), .Y(n3548) );
  OAI21X1 U2693 ( .A(n4717), .B(n4670), .C(n5112), .Y(n5111) );
  OAI22X1 U2694 ( .A(n4579), .B(n5113), .C(n4647), .D(n5113), .Y(n5112) );
  OAI22X1 U2695 ( .A(n4580), .B(n4651), .C(n4582), .D(n4648), .Y(n5113) );
  XNOR2X1 U2696 ( .A(n5114), .B(n4649), .Y(n3547) );
  OAI21X1 U2697 ( .A(n4716), .B(n4670), .C(n5115), .Y(n5114) );
  OAI22X1 U2698 ( .A(n4581), .B(n5116), .C(n4647), .D(n5116), .Y(n5115) );
  OAI22X1 U2699 ( .A(n4582), .B(n4651), .C(n4584), .D(n4648), .Y(n5116) );
  XNOR2X1 U2700 ( .A(n5117), .B(n4649), .Y(n3546) );
  OAI21X1 U2701 ( .A(n4715), .B(n4670), .C(n5118), .Y(n5117) );
  OAI22X1 U2702 ( .A(n4583), .B(n5119), .C(n4647), .D(n5119), .Y(n5118) );
  OAI22X1 U2703 ( .A(n4584), .B(n4651), .C(n4587), .D(n4648), .Y(n5119) );
  XNOR2X1 U2704 ( .A(n5120), .B(n4649), .Y(n3545) );
  OAI21X1 U2705 ( .A(n4713), .B(n4670), .C(n5121), .Y(n5120) );
  OAI22X1 U2706 ( .A(n4585), .B(n5122), .C(n4647), .D(n5122), .Y(n5121) );
  OAI22X1 U2707 ( .A(n4587), .B(n4651), .C(n4589), .D(n4648), .Y(n5122) );
  XNOR2X1 U2708 ( .A(n5123), .B(n4649), .Y(n3544) );
  OAI21X1 U2709 ( .A(n4712), .B(n4670), .C(n5124), .Y(n5123) );
  OAI22X1 U2710 ( .A(n4588), .B(n5125), .C(n4647), .D(n5125), .Y(n5124) );
  OAI22X1 U2711 ( .A(n4589), .B(n4651), .C(n4592), .D(n4648), .Y(n5125) );
  XNOR2X1 U2712 ( .A(n5126), .B(n4649), .Y(n3543) );
  OAI21X1 U2713 ( .A(n4711), .B(n4670), .C(n5127), .Y(n5126) );
  OAI22X1 U2714 ( .A(n4590), .B(n5128), .C(n4647), .D(n5128), .Y(n5127) );
  OAI22X1 U2715 ( .A(n4592), .B(n4651), .C(n4594), .D(n4648), .Y(n5128) );
  XNOR2X1 U2716 ( .A(n5129), .B(n4649), .Y(n3542) );
  OAI21X1 U2717 ( .A(n4710), .B(n4670), .C(n5130), .Y(n5129) );
  OAI22X1 U2718 ( .A(n4593), .B(n5131), .C(n4647), .D(n5131), .Y(n5130) );
  OAI22X1 U2719 ( .A(n4594), .B(n4651), .C(n4726), .D(n4648), .Y(n5131) );
  XNOR2X1 U2720 ( .A(n5132), .B(n4649), .Y(n3541) );
  OAI21X1 U2721 ( .A(n4708), .B(n4670), .C(n5133), .Y(n5132) );
  OAI22X1 U2722 ( .A(n4595), .B(n5134), .C(n4647), .D(n5134), .Y(n5133) );
  OAI22X1 U2723 ( .A(n4726), .B(n4651), .C(n4599), .D(n4648), .Y(n5134) );
  XNOR2X1 U2724 ( .A(n5135), .B(n4649), .Y(n3540) );
  OAI21X1 U2725 ( .A(n4707), .B(n4670), .C(n5136), .Y(n5135) );
  OAI22X1 U2726 ( .A(n4598), .B(n5137), .C(n4647), .D(n5137), .Y(n5136) );
  OAI22X1 U2727 ( .A(n4599), .B(n4651), .C(n4601), .D(n4648), .Y(n5137) );
  XNOR2X1 U2728 ( .A(n5138), .B(n4649), .Y(n3539) );
  OAI21X1 U2729 ( .A(n4706), .B(n4670), .C(n5139), .Y(n5138) );
  OAI22X1 U2730 ( .A(b[15]), .B(n5140), .C(n4647), .D(n5140), .Y(n5139) );
  OAI22X1 U2731 ( .A(n4601), .B(n4651), .C(n4603), .D(n4648), .Y(n5140) );
  XNOR2X1 U2732 ( .A(n5141), .B(n4649), .Y(n3538) );
  OAI21X1 U2733 ( .A(n4705), .B(n4670), .C(n5142), .Y(n5141) );
  OAI22X1 U2734 ( .A(n4602), .B(n5143), .C(n4647), .D(n5143), .Y(n5142) );
  OAI22X1 U2735 ( .A(n4603), .B(n4651), .C(n4606), .D(n4648), .Y(n5143) );
  XNOR2X1 U2736 ( .A(n5144), .B(n4649), .Y(n3537) );
  OAI21X1 U2737 ( .A(n4704), .B(n4670), .C(n5145), .Y(n5144) );
  OAI22X1 U2738 ( .A(n4605), .B(n5146), .C(n4647), .D(n5146), .Y(n5145) );
  OAI22X1 U2739 ( .A(n4606), .B(n4651), .C(n4608), .D(n4648), .Y(n5146) );
  XNOR2X1 U2740 ( .A(n5147), .B(n4650), .Y(n3536) );
  OAI21X1 U2741 ( .A(n4703), .B(n4670), .C(n5148), .Y(n5147) );
  OAI22X1 U2742 ( .A(n4607), .B(n5149), .C(n4647), .D(n5149), .Y(n5148) );
  OAI22X1 U2743 ( .A(n4608), .B(n4651), .C(n4611), .D(n4648), .Y(n5149) );
  XNOR2X1 U2744 ( .A(n5150), .B(n4650), .Y(n3535) );
  OAI21X1 U2745 ( .A(n4702), .B(n4670), .C(n5151), .Y(n5150) );
  OAI22X1 U2746 ( .A(n4609), .B(n5152), .C(n4647), .D(n5152), .Y(n5151) );
  OAI22X1 U2747 ( .A(n4611), .B(n4651), .C(n4613), .D(n4648), .Y(n5152) );
  XNOR2X1 U2748 ( .A(n5153), .B(n4650), .Y(n3534) );
  OAI21X1 U2749 ( .A(n4701), .B(n4670), .C(n5154), .Y(n5153) );
  OAI22X1 U2750 ( .A(n4612), .B(n5155), .C(n4647), .D(n5155), .Y(n5154) );
  OAI22X1 U2751 ( .A(n4613), .B(n4651), .C(n4616), .D(n4648), .Y(n5155) );
  XNOR2X1 U2752 ( .A(n5156), .B(n4650), .Y(n3533) );
  OAI21X1 U2753 ( .A(n4700), .B(n4670), .C(n5157), .Y(n5156) );
  OAI22X1 U2754 ( .A(n4615), .B(n5158), .C(n4647), .D(n5158), .Y(n5157) );
  OAI22X1 U2755 ( .A(n4616), .B(n4651), .C(n4618), .D(n4648), .Y(n5158) );
  XNOR2X1 U2756 ( .A(n5159), .B(n4650), .Y(n3532) );
  OAI21X1 U2757 ( .A(n4699), .B(n4670), .C(n5160), .Y(n5159) );
  OAI22X1 U2758 ( .A(n4617), .B(n5161), .C(n4647), .D(n5161), .Y(n5160) );
  OAI22X1 U2759 ( .A(n4618), .B(n4651), .C(n4620), .D(n4648), .Y(n5161) );
  XNOR2X1 U2760 ( .A(n5162), .B(n4650), .Y(n3531) );
  OAI21X1 U2761 ( .A(n4698), .B(n4670), .C(n5163), .Y(n5162) );
  OAI22X1 U2762 ( .A(n4619), .B(n5164), .C(n4647), .D(n5164), .Y(n5163) );
  OAI22X1 U2763 ( .A(n4620), .B(n4651), .C(n4622), .D(n4648), .Y(n5164) );
  XNOR2X1 U2764 ( .A(n5165), .B(n4650), .Y(n3530) );
  OAI21X1 U2765 ( .A(n4697), .B(n4670), .C(n5166), .Y(n5165) );
  OAI22X1 U2766 ( .A(n4621), .B(n5167), .C(n4647), .D(n5167), .Y(n5166) );
  OAI22X1 U2767 ( .A(n4622), .B(n4651), .C(n4624), .D(n4648), .Y(n5167) );
  XNOR2X1 U2768 ( .A(n5168), .B(n4650), .Y(n3529) );
  OAI21X1 U2769 ( .A(n4696), .B(n4670), .C(n5169), .Y(n5168) );
  OAI22X1 U2770 ( .A(n4623), .B(n5170), .C(n4647), .D(n5170), .Y(n5169) );
  OAI22X1 U2771 ( .A(n4624), .B(n4651), .C(n4626), .D(n4648), .Y(n5170) );
  XNOR2X1 U2772 ( .A(n5171), .B(n4650), .Y(n3528) );
  OAI21X1 U2773 ( .A(n4695), .B(n4670), .C(n5172), .Y(n5171) );
  OAI22X1 U2774 ( .A(n4625), .B(n5173), .C(n4647), .D(n5173), .Y(n5172) );
  OAI22X1 U2775 ( .A(n4626), .B(n4651), .C(n4628), .D(n4648), .Y(n5173) );
  XNOR2X1 U2776 ( .A(n5174), .B(n4650), .Y(n3527) );
  OAI21X1 U2777 ( .A(n4694), .B(n4670), .C(n5175), .Y(n5174) );
  OAI22X1 U2778 ( .A(n4627), .B(n5176), .C(n4647), .D(n5176), .Y(n5175) );
  OAI22X1 U2779 ( .A(n4628), .B(n4651), .C(n4630), .D(n4648), .Y(n5176) );
  XNOR2X1 U2780 ( .A(n5177), .B(n4650), .Y(n3526) );
  OAI21X1 U2781 ( .A(n4693), .B(n4670), .C(n5178), .Y(n5177) );
  OAI22X1 U2782 ( .A(n4629), .B(n5179), .C(n4647), .D(n5179), .Y(n5178) );
  OAI22X1 U2783 ( .A(n4630), .B(n4651), .C(n4632), .D(n4648), .Y(n5179) );
  XNOR2X1 U2784 ( .A(n5180), .B(n4650), .Y(n3525) );
  OAI21X1 U2785 ( .A(n4690), .B(n4670), .C(n5181), .Y(n5180) );
  OAI22X1 U2786 ( .A(n4631), .B(n5182), .C(n4647), .D(n5182), .Y(n5181) );
  OAI22X1 U2787 ( .A(n4632), .B(n4651), .C(n4687), .D(n4648), .Y(n5182) );
  NOR2X1 U2788 ( .A(n5183), .B(n5184), .Y(n5092) );
  XNOR2X1 U2789 ( .A(n5185), .B(n4650), .Y(n3524) );
  OAI21X1 U2790 ( .A(n4689), .B(n4670), .C(n5186), .Y(n5185) );
  OAI22X1 U2791 ( .A(n4633), .B(n5187), .C(n4647), .D(n5187), .Y(n5186) );
  NOR2X1 U2792 ( .A(n4651), .B(n4687), .Y(n5187) );
  NOR2X1 U2793 ( .A(n4743), .B(n5189), .Y(n5091) );
  XNOR2X1 U2794 ( .A(n5190), .B(n4650), .Y(n3523) );
  OAI22X1 U2795 ( .A(n4687), .B(n5188), .C(n4688), .D(n4670), .Y(n5190) );
  NAND3X1 U2796 ( .A(n5184), .B(n5183), .C(n5189), .Y(n5188) );
  XNOR2X1 U2797 ( .A(a[10]), .B(a[9]), .Y(n5189) );
  XNOR2X1 U2798 ( .A(a[10]), .B(n4650), .Y(n5183) );
  XOR2X1 U2799 ( .A(a[9]), .B(n4655), .Y(n5184) );
  XNOR2X1 U2800 ( .A(n5191), .B(n4644), .Y(n3521) );
  OAI22X1 U2801 ( .A(n4686), .B(n4643), .C(n4686), .D(n4671), .Y(n5191) );
  XNOR2X1 U2802 ( .A(n5192), .B(n4644), .Y(n3520) );
  OAI21X1 U2803 ( .A(n4725), .B(n4671), .C(n5193), .Y(n5192) );
  AOI22X1 U2804 ( .A(n5194), .B(n4684), .C(n5195), .D(n4680), .Y(n5193) );
  XNOR2X1 U2805 ( .A(n5196), .B(n4644), .Y(n3519) );
  OAI21X1 U2806 ( .A(n4724), .B(n4671), .C(n5197), .Y(n5196) );
  OAI22X1 U2807 ( .A(n4685), .B(n5198), .C(n4642), .D(n5198), .Y(n5197) );
  OAI22X1 U2808 ( .A(n4681), .B(n4646), .C(n4568), .D(n4643), .Y(n5198) );
  XNOR2X1 U2809 ( .A(n5199), .B(n4644), .Y(n3518) );
  OAI21X1 U2810 ( .A(n4723), .B(n4671), .C(n5200), .Y(n5199) );
  OAI22X1 U2811 ( .A(n4680), .B(n5201), .C(n4642), .D(n5201), .Y(n5200) );
  OAI22X1 U2812 ( .A(n4568), .B(n4646), .C(n4570), .D(n4643), .Y(n5201) );
  XNOR2X1 U2813 ( .A(n5202), .B(n4644), .Y(n3517) );
  OAI21X1 U2814 ( .A(n4722), .B(n4671), .C(n5203), .Y(n5202) );
  OAI22X1 U2815 ( .A(b[2]), .B(n5204), .C(n4642), .D(n5204), .Y(n5203) );
  OAI22X1 U2816 ( .A(n4570), .B(n4646), .C(n4573), .D(n4643), .Y(n5204) );
  XNOR2X1 U2817 ( .A(n5205), .B(n4644), .Y(n3516) );
  OAI21X1 U2818 ( .A(n4721), .B(n4671), .C(n5206), .Y(n5205) );
  OAI22X1 U2819 ( .A(n4572), .B(n5207), .C(n4642), .D(n5207), .Y(n5206) );
  OAI22X1 U2820 ( .A(n4573), .B(n4646), .C(n4575), .D(n4643), .Y(n5207) );
  XNOR2X1 U2821 ( .A(n5208), .B(n4644), .Y(n3515) );
  OAI21X1 U2822 ( .A(n4720), .B(n4671), .C(n5209), .Y(n5208) );
  OAI22X1 U2823 ( .A(b[4]), .B(n5210), .C(n4642), .D(n5210), .Y(n5209) );
  OAI22X1 U2824 ( .A(n4575), .B(n4646), .C(n4578), .D(n4643), .Y(n5210) );
  XNOR2X1 U2825 ( .A(n5211), .B(n4644), .Y(n3514) );
  OAI21X1 U2826 ( .A(n4719), .B(n4671), .C(n5212), .Y(n5211) );
  OAI22X1 U2827 ( .A(n4577), .B(n5213), .C(n4642), .D(n5213), .Y(n5212) );
  OAI22X1 U2828 ( .A(n4578), .B(n4646), .C(n4580), .D(n4643), .Y(n5213) );
  XNOR2X1 U2829 ( .A(n5214), .B(n4644), .Y(n3513) );
  OAI21X1 U2830 ( .A(n4717), .B(n4671), .C(n5215), .Y(n5214) );
  OAI22X1 U2831 ( .A(b[6]), .B(n5216), .C(n4642), .D(n5216), .Y(n5215) );
  OAI22X1 U2832 ( .A(n4580), .B(n4646), .C(n4582), .D(n4643), .Y(n5216) );
  XNOR2X1 U2833 ( .A(n5217), .B(n4644), .Y(n3512) );
  OAI21X1 U2834 ( .A(n4716), .B(n4671), .C(n5218), .Y(n5217) );
  OAI22X1 U2835 ( .A(b[7]), .B(n5219), .C(n4642), .D(n5219), .Y(n5218) );
  OAI22X1 U2836 ( .A(n4582), .B(n4646), .C(n4584), .D(n4643), .Y(n5219) );
  XNOR2X1 U2837 ( .A(n5220), .B(n4644), .Y(n3511) );
  OAI21X1 U2838 ( .A(n4715), .B(n4671), .C(n5221), .Y(n5220) );
  OAI22X1 U2839 ( .A(b[8]), .B(n5222), .C(n4642), .D(n5222), .Y(n5221) );
  OAI22X1 U2840 ( .A(n4584), .B(n4646), .C(n4587), .D(n4643), .Y(n5222) );
  XNOR2X1 U2841 ( .A(n5223), .B(n4644), .Y(n3510) );
  OAI21X1 U2842 ( .A(n4713), .B(n4671), .C(n5224), .Y(n5223) );
  OAI22X1 U2843 ( .A(n4586), .B(n5225), .C(n4642), .D(n5225), .Y(n5224) );
  OAI22X1 U2844 ( .A(n4587), .B(n4646), .C(n4589), .D(n4643), .Y(n5225) );
  XNOR2X1 U2845 ( .A(n5226), .B(n4644), .Y(n3509) );
  OAI21X1 U2846 ( .A(n4712), .B(n4671), .C(n5227), .Y(n5226) );
  OAI22X1 U2847 ( .A(b[10]), .B(n5228), .C(n4642), .D(n5228), .Y(n5227) );
  OAI22X1 U2848 ( .A(n4589), .B(n4646), .C(n4592), .D(n4643), .Y(n5228) );
  XNOR2X1 U2849 ( .A(n5229), .B(n4644), .Y(n3508) );
  OAI21X1 U2850 ( .A(n4711), .B(n4671), .C(n5230), .Y(n5229) );
  OAI22X1 U2851 ( .A(n4591), .B(n5231), .C(n4642), .D(n5231), .Y(n5230) );
  OAI22X1 U2852 ( .A(n4592), .B(n4646), .C(n4594), .D(n4643), .Y(n5231) );
  XNOR2X1 U2853 ( .A(n5232), .B(n4644), .Y(n3507) );
  OAI21X1 U2854 ( .A(n4710), .B(n4671), .C(n5233), .Y(n5232) );
  OAI22X1 U2855 ( .A(b[12]), .B(n5234), .C(n4642), .D(n5234), .Y(n5233) );
  OAI22X1 U2856 ( .A(n4594), .B(n4646), .C(n4726), .D(n4643), .Y(n5234) );
  XNOR2X1 U2857 ( .A(n5235), .B(n4644), .Y(n3506) );
  OAI21X1 U2858 ( .A(n4708), .B(n4671), .C(n5236), .Y(n5235) );
  OAI22X1 U2859 ( .A(n4596), .B(n5237), .C(n4642), .D(n5237), .Y(n5236) );
  OAI22X1 U2860 ( .A(n4726), .B(n4646), .C(n4599), .D(n4643), .Y(n5237) );
  XNOR2X1 U2861 ( .A(n5238), .B(n4644), .Y(n3505) );
  OAI21X1 U2862 ( .A(n4707), .B(n4671), .C(n5239), .Y(n5238) );
  OAI22X1 U2863 ( .A(b[14]), .B(n5240), .C(n4642), .D(n5240), .Y(n5239) );
  OAI22X1 U2864 ( .A(n4599), .B(n4646), .C(n4601), .D(n4643), .Y(n5240) );
  XNOR2X1 U2865 ( .A(n5241), .B(n4644), .Y(n3504) );
  OAI21X1 U2866 ( .A(n4706), .B(n4671), .C(n5242), .Y(n5241) );
  OAI22X1 U2867 ( .A(n4600), .B(n5243), .C(n4642), .D(n5243), .Y(n5242) );
  OAI22X1 U2868 ( .A(n4601), .B(n4646), .C(n4603), .D(n4643), .Y(n5243) );
  XNOR2X1 U2869 ( .A(n5244), .B(n4644), .Y(n3503) );
  OAI21X1 U2870 ( .A(n4705), .B(n4671), .C(n5245), .Y(n5244) );
  OAI22X1 U2871 ( .A(n4602), .B(n5246), .C(n4642), .D(n5246), .Y(n5245) );
  OAI22X1 U2872 ( .A(n4603), .B(n4646), .C(n4606), .D(n4643), .Y(n5246) );
  XNOR2X1 U2873 ( .A(n5247), .B(n4644), .Y(n3502) );
  OAI21X1 U2874 ( .A(n4704), .B(n4671), .C(n5248), .Y(n5247) );
  OAI22X1 U2875 ( .A(n4605), .B(n5249), .C(n4642), .D(n5249), .Y(n5248) );
  OAI22X1 U2876 ( .A(n4606), .B(n4646), .C(n4608), .D(n4643), .Y(n5249) );
  XNOR2X1 U2877 ( .A(n5250), .B(n4645), .Y(n3501) );
  OAI21X1 U2878 ( .A(n4703), .B(n4671), .C(n5251), .Y(n5250) );
  OAI22X1 U2879 ( .A(n4607), .B(n5252), .C(n4642), .D(n5252), .Y(n5251) );
  OAI22X1 U2880 ( .A(n4608), .B(n4646), .C(n4611), .D(n4643), .Y(n5252) );
  XNOR2X1 U2881 ( .A(n5253), .B(n4645), .Y(n3500) );
  OAI21X1 U2882 ( .A(n4702), .B(n4671), .C(n5254), .Y(n5253) );
  OAI22X1 U2883 ( .A(n4610), .B(n5255), .C(n4642), .D(n5255), .Y(n5254) );
  OAI22X1 U2884 ( .A(n4611), .B(n4646), .C(n4613), .D(n4643), .Y(n5255) );
  XNOR2X1 U2885 ( .A(n5256), .B(n4645), .Y(n3499) );
  OAI21X1 U2886 ( .A(n4701), .B(n4671), .C(n5257), .Y(n5256) );
  OAI22X1 U2887 ( .A(b[20]), .B(n5258), .C(n4642), .D(n5258), .Y(n5257) );
  OAI22X1 U2888 ( .A(n4613), .B(n4646), .C(n4616), .D(n4643), .Y(n5258) );
  XNOR2X1 U2889 ( .A(n5259), .B(n4645), .Y(n3498) );
  OAI21X1 U2890 ( .A(n4700), .B(n4671), .C(n5260), .Y(n5259) );
  OAI22X1 U2891 ( .A(n4614), .B(n5261), .C(n4642), .D(n5261), .Y(n5260) );
  OAI22X1 U2892 ( .A(n4616), .B(n4646), .C(n4618), .D(n4643), .Y(n5261) );
  XNOR2X1 U2893 ( .A(n5262), .B(n4645), .Y(n3497) );
  OAI21X1 U2894 ( .A(n4699), .B(n4671), .C(n5263), .Y(n5262) );
  OAI22X1 U2895 ( .A(n4617), .B(n5264), .C(n4642), .D(n5264), .Y(n5263) );
  OAI22X1 U2896 ( .A(n4618), .B(n4646), .C(n4620), .D(n4643), .Y(n5264) );
  XNOR2X1 U2897 ( .A(n5265), .B(n4645), .Y(n3496) );
  OAI21X1 U2898 ( .A(n4698), .B(n4671), .C(n5266), .Y(n5265) );
  OAI22X1 U2899 ( .A(n4619), .B(n5267), .C(n4642), .D(n5267), .Y(n5266) );
  OAI22X1 U2900 ( .A(n4620), .B(n4646), .C(n4622), .D(n4643), .Y(n5267) );
  XNOR2X1 U2901 ( .A(n5268), .B(n4645), .Y(n3495) );
  OAI21X1 U2902 ( .A(n4697), .B(n4671), .C(n5269), .Y(n5268) );
  OAI22X1 U2903 ( .A(n4621), .B(n5270), .C(n4642), .D(n5270), .Y(n5269) );
  OAI22X1 U2904 ( .A(n4622), .B(n4646), .C(n4624), .D(n4643), .Y(n5270) );
  XNOR2X1 U2905 ( .A(n5271), .B(n4645), .Y(n3494) );
  OAI21X1 U2906 ( .A(n4696), .B(n4671), .C(n5272), .Y(n5271) );
  OAI22X1 U2907 ( .A(n4623), .B(n5273), .C(n4642), .D(n5273), .Y(n5272) );
  OAI22X1 U2908 ( .A(n4624), .B(n4646), .C(n4626), .D(n4643), .Y(n5273) );
  XNOR2X1 U2909 ( .A(n5274), .B(n4645), .Y(n3493) );
  OAI21X1 U2910 ( .A(n4695), .B(n4671), .C(n5275), .Y(n5274) );
  OAI22X1 U2911 ( .A(n4625), .B(n5276), .C(n4642), .D(n5276), .Y(n5275) );
  OAI22X1 U2912 ( .A(n4626), .B(n4646), .C(n4628), .D(n4643), .Y(n5276) );
  XNOR2X1 U2913 ( .A(n5277), .B(n4645), .Y(n3492) );
  OAI21X1 U2914 ( .A(n4694), .B(n4671), .C(n5278), .Y(n5277) );
  OAI22X1 U2915 ( .A(n4627), .B(n5279), .C(n4642), .D(n5279), .Y(n5278) );
  OAI22X1 U2916 ( .A(n4628), .B(n4646), .C(n4630), .D(n4643), .Y(n5279) );
  XNOR2X1 U2917 ( .A(n5280), .B(n4645), .Y(n3491) );
  OAI21X1 U2918 ( .A(n4693), .B(n4671), .C(n5281), .Y(n5280) );
  OAI22X1 U2919 ( .A(n4629), .B(n5282), .C(n4642), .D(n5282), .Y(n5281) );
  OAI22X1 U2920 ( .A(n4630), .B(n4646), .C(n4632), .D(n4643), .Y(n5282) );
  XNOR2X1 U2921 ( .A(n5283), .B(n4645), .Y(n3490) );
  OAI21X1 U2922 ( .A(n4690), .B(n4671), .C(n5284), .Y(n5283) );
  OAI22X1 U2923 ( .A(n4631), .B(n5285), .C(n4642), .D(n5285), .Y(n5284) );
  OAI22X1 U2924 ( .A(n4632), .B(n4646), .C(n4687), .D(n4643), .Y(n5285) );
  NOR2X1 U2925 ( .A(n5286), .B(n5287), .Y(n5195) );
  XNOR2X1 U2926 ( .A(n5288), .B(n4645), .Y(n3489) );
  OAI21X1 U2927 ( .A(n4689), .B(n4671), .C(n5289), .Y(n5288) );
  OAI22X1 U2928 ( .A(n4633), .B(n5290), .C(n4642), .D(n5290), .Y(n5289) );
  NOR2X1 U2929 ( .A(n4646), .B(n4687), .Y(n5290) );
  NOR2X1 U2930 ( .A(n4742), .B(n5292), .Y(n5194) );
  XNOR2X1 U2931 ( .A(n5293), .B(n4645), .Y(n3488) );
  OAI22X1 U2932 ( .A(n4687), .B(n5291), .C(n4688), .D(n4671), .Y(n5293) );
  NAND3X1 U2933 ( .A(n5287), .B(n5286), .C(n5292), .Y(n5291) );
  XNOR2X1 U2934 ( .A(a[12]), .B(a[13]), .Y(n5292) );
  XNOR2X1 U2935 ( .A(a[13]), .B(n4645), .Y(n5286) );
  XOR2X1 U2936 ( .A(a[12]), .B(n4650), .Y(n5287) );
  XNOR2X1 U2937 ( .A(n5294), .B(n4640), .Y(n3486) );
  OAI22X1 U2938 ( .A(n4686), .B(n4554), .C(n4664), .D(n4686), .Y(n5294) );
  XNOR2X1 U2939 ( .A(n5295), .B(n4640), .Y(n3485) );
  OAI21X1 U2940 ( .A(n4664), .B(n4725), .C(n4691), .Y(n5295) );
  OAI22X1 U2941 ( .A(n4686), .B(n4552), .C(n4554), .D(n4681), .Y(n5296) );
  XNOR2X1 U2942 ( .A(n5297), .B(n4640), .Y(n3484) );
  OAI21X1 U2943 ( .A(n4664), .B(n4724), .C(n5298), .Y(n5297) );
  OAI22X1 U2944 ( .A(n4685), .B(n5299), .C(n4639), .D(n5299), .Y(n5298) );
  OAI22X1 U2945 ( .A(n4568), .B(n4554), .C(n4552), .D(n4681), .Y(n5299) );
  XNOR2X1 U2946 ( .A(n5300), .B(n4640), .Y(n3483) );
  OAI21X1 U2947 ( .A(n4664), .B(n4723), .C(n5301), .Y(n5300) );
  OAI22X1 U2948 ( .A(n4680), .B(n5302), .C(n4639), .D(n5302), .Y(n5301) );
  OAI22X1 U2949 ( .A(n4570), .B(n4554), .C(n4552), .D(n4568), .Y(n5302) );
  XNOR2X1 U2950 ( .A(n5303), .B(n4640), .Y(n3482) );
  OAI21X1 U2951 ( .A(n4664), .B(n4722), .C(n5304), .Y(n5303) );
  OAI22X1 U2952 ( .A(n4569), .B(n5305), .C(n4639), .D(n5305), .Y(n5304) );
  OAI22X1 U2953 ( .A(n4573), .B(n4554), .C(n4552), .D(n4570), .Y(n5305) );
  XNOR2X1 U2954 ( .A(n5306), .B(n4640), .Y(n3481) );
  OAI21X1 U2955 ( .A(n4664), .B(n4721), .C(n5307), .Y(n5306) );
  OAI22X1 U2956 ( .A(n4571), .B(n5308), .C(n4639), .D(n5308), .Y(n5307) );
  OAI22X1 U2957 ( .A(n4575), .B(n4554), .C(n4552), .D(n4573), .Y(n5308) );
  XNOR2X1 U2958 ( .A(n5309), .B(n4640), .Y(n3480) );
  OAI21X1 U2959 ( .A(n4664), .B(n4720), .C(n5310), .Y(n5309) );
  OAI22X1 U2960 ( .A(n4574), .B(n5311), .C(n4639), .D(n5311), .Y(n5310) );
  OAI22X1 U2961 ( .A(n4578), .B(n4554), .C(n4552), .D(n4575), .Y(n5311) );
  XNOR2X1 U2962 ( .A(n5312), .B(n4640), .Y(n3479) );
  OAI21X1 U2963 ( .A(n4664), .B(n4719), .C(n5313), .Y(n5312) );
  OAI22X1 U2964 ( .A(n4576), .B(n5314), .C(n4639), .D(n5314), .Y(n5313) );
  OAI22X1 U2965 ( .A(n4580), .B(n4554), .C(n4552), .D(n4578), .Y(n5314) );
  XNOR2X1 U2966 ( .A(n5315), .B(n4640), .Y(n3478) );
  OAI21X1 U2967 ( .A(n4664), .B(n4717), .C(n5316), .Y(n5315) );
  OAI22X1 U2968 ( .A(n4579), .B(n5317), .C(n4639), .D(n5317), .Y(n5316) );
  OAI22X1 U2969 ( .A(n4582), .B(n4554), .C(n4552), .D(n4580), .Y(n5317) );
  XNOR2X1 U2970 ( .A(n5318), .B(n4640), .Y(n3477) );
  OAI21X1 U2971 ( .A(n4664), .B(n4716), .C(n5319), .Y(n5318) );
  OAI22X1 U2972 ( .A(n4581), .B(n5320), .C(n4639), .D(n5320), .Y(n5319) );
  OAI22X1 U2973 ( .A(n4584), .B(n4554), .C(n4552), .D(n4582), .Y(n5320) );
  XNOR2X1 U2974 ( .A(n5321), .B(n4640), .Y(n3476) );
  OAI21X1 U2975 ( .A(n4664), .B(n4715), .C(n5322), .Y(n5321) );
  OAI22X1 U2976 ( .A(n4583), .B(n5323), .C(n4639), .D(n5323), .Y(n5322) );
  OAI22X1 U2977 ( .A(n4587), .B(n4554), .C(n4552), .D(n4584), .Y(n5323) );
  XNOR2X1 U2978 ( .A(n5324), .B(n4640), .Y(n3475) );
  OAI21X1 U2979 ( .A(n4664), .B(n4713), .C(n5325), .Y(n5324) );
  OAI22X1 U2980 ( .A(n4585), .B(n5326), .C(n4639), .D(n5326), .Y(n5325) );
  OAI22X1 U2981 ( .A(n4589), .B(n4554), .C(n4552), .D(n4587), .Y(n5326) );
  XNOR2X1 U2982 ( .A(n5327), .B(n4640), .Y(n3474) );
  OAI21X1 U2983 ( .A(n4664), .B(n4712), .C(n5328), .Y(n5327) );
  OAI22X1 U2984 ( .A(n4588), .B(n5329), .C(n4639), .D(n5329), .Y(n5328) );
  OAI22X1 U2985 ( .A(n4592), .B(n4554), .C(n4552), .D(n4589), .Y(n5329) );
  XNOR2X1 U2986 ( .A(n5330), .B(n4640), .Y(n3473) );
  OAI21X1 U2987 ( .A(n4664), .B(n4711), .C(n5331), .Y(n5330) );
  OAI22X1 U2988 ( .A(n4590), .B(n5332), .C(n4639), .D(n5332), .Y(n5331) );
  OAI22X1 U2989 ( .A(n4594), .B(n4554), .C(n4552), .D(n4592), .Y(n5332) );
  XNOR2X1 U2990 ( .A(n5333), .B(n4640), .Y(n3472) );
  OAI21X1 U2991 ( .A(n4664), .B(n4710), .C(n5334), .Y(n5333) );
  OAI22X1 U2992 ( .A(n4593), .B(n5335), .C(n4639), .D(n5335), .Y(n5334) );
  OAI22X1 U2993 ( .A(n4726), .B(n4554), .C(n4552), .D(n4594), .Y(n5335) );
  XNOR2X1 U2994 ( .A(n5336), .B(n4640), .Y(n3471) );
  OAI21X1 U2995 ( .A(n4664), .B(n4708), .C(n5337), .Y(n5336) );
  OAI22X1 U2996 ( .A(n4595), .B(n5338), .C(n4639), .D(n5338), .Y(n5337) );
  OAI22X1 U2997 ( .A(n4599), .B(n4554), .C(n4552), .D(n4726), .Y(n5338) );
  XNOR2X1 U2998 ( .A(n5339), .B(n4640), .Y(n3470) );
  OAI21X1 U2999 ( .A(n4664), .B(n4707), .C(n5340), .Y(n5339) );
  OAI22X1 U3000 ( .A(n4598), .B(n5341), .C(n4639), .D(n5341), .Y(n5340) );
  OAI22X1 U3001 ( .A(n4601), .B(n4554), .C(n4552), .D(n4599), .Y(n5341) );
  XNOR2X1 U3002 ( .A(n5342), .B(n4640), .Y(n3469) );
  OAI21X1 U3003 ( .A(n4706), .B(n4664), .C(n5343), .Y(n5342) );
  OAI22X1 U3004 ( .A(b[15]), .B(n5344), .C(n4639), .D(n5344), .Y(n5343) );
  OAI22X1 U3005 ( .A(n4603), .B(n4554), .C(n4601), .D(n4552), .Y(n5344) );
  XNOR2X1 U3006 ( .A(n5345), .B(n4640), .Y(n3468) );
  OAI21X1 U3007 ( .A(n4664), .B(n4705), .C(n5346), .Y(n5345) );
  OAI22X1 U3008 ( .A(n4602), .B(n5347), .C(n4639), .D(n5347), .Y(n5346) );
  OAI22X1 U3009 ( .A(n4606), .B(n4554), .C(n4603), .D(n4552), .Y(n5347) );
  XNOR2X1 U3010 ( .A(n5348), .B(n4640), .Y(n3467) );
  OAI21X1 U3011 ( .A(n4664), .B(n4704), .C(n5349), .Y(n5348) );
  OAI22X1 U3012 ( .A(n4605), .B(n5350), .C(n4639), .D(n5350), .Y(n5349) );
  OAI22X1 U3013 ( .A(n4608), .B(n4554), .C(n4552), .D(n4606), .Y(n5350) );
  XNOR2X1 U3014 ( .A(n5351), .B(n4640), .Y(n3466) );
  OAI21X1 U3015 ( .A(n4703), .B(n4664), .C(n5352), .Y(n5351) );
  OAI22X1 U3016 ( .A(n4607), .B(n5353), .C(n4639), .D(n5353), .Y(n5352) );
  OAI22X1 U3017 ( .A(n4611), .B(n4554), .C(n4608), .D(n4552), .Y(n5353) );
  XNOR2X1 U3018 ( .A(n5354), .B(n4640), .Y(n3465) );
  OAI21X1 U3019 ( .A(n4664), .B(n4702), .C(n5355), .Y(n5354) );
  OAI22X1 U3020 ( .A(n4609), .B(n5356), .C(n4639), .D(n5356), .Y(n5355) );
  OAI22X1 U3021 ( .A(n4613), .B(n4554), .C(n4611), .D(n4552), .Y(n5356) );
  XNOR2X1 U3022 ( .A(n5357), .B(n4640), .Y(n3464) );
  OAI21X1 U3023 ( .A(n4664), .B(n4701), .C(n5358), .Y(n5357) );
  OAI22X1 U3024 ( .A(n4612), .B(n5359), .C(n4639), .D(n5359), .Y(n5358) );
  OAI22X1 U3025 ( .A(n4616), .B(n4554), .C(n4552), .D(n4613), .Y(n5359) );
  XNOR2X1 U3026 ( .A(n5360), .B(n4640), .Y(n3463) );
  OAI21X1 U3027 ( .A(n4700), .B(n4664), .C(n5361), .Y(n5360) );
  OAI22X1 U3028 ( .A(n4615), .B(n5362), .C(n4639), .D(n5362), .Y(n5361) );
  OAI22X1 U3029 ( .A(n4618), .B(n4554), .C(n4616), .D(n4552), .Y(n5362) );
  XNOR2X1 U3030 ( .A(n5363), .B(n4641), .Y(n3462) );
  OAI21X1 U3031 ( .A(n4664), .B(n4699), .C(n5364), .Y(n5363) );
  OAI22X1 U3032 ( .A(n4617), .B(n5365), .C(n4639), .D(n5365), .Y(n5364) );
  OAI22X1 U3033 ( .A(n4620), .B(n4554), .C(n4618), .D(n4552), .Y(n5365) );
  XNOR2X1 U3034 ( .A(n5366), .B(n4641), .Y(n3461) );
  OAI21X1 U3035 ( .A(n4664), .B(n4698), .C(n5367), .Y(n5366) );
  OAI22X1 U3036 ( .A(n4619), .B(n5368), .C(n4639), .D(n5368), .Y(n5367) );
  OAI22X1 U3037 ( .A(n4622), .B(n4554), .C(n4552), .D(n4620), .Y(n5368) );
  XNOR2X1 U3038 ( .A(n5369), .B(n4641), .Y(n3460) );
  OAI21X1 U3039 ( .A(n4697), .B(n4664), .C(n5370), .Y(n5369) );
  OAI22X1 U3040 ( .A(n4621), .B(n5371), .C(n4639), .D(n5371), .Y(n5370) );
  OAI22X1 U3041 ( .A(n4624), .B(n4554), .C(n4622), .D(n4552), .Y(n5371) );
  XNOR2X1 U3042 ( .A(n5372), .B(n4641), .Y(n3459) );
  OAI21X1 U3043 ( .A(n4664), .B(n4696), .C(n5373), .Y(n5372) );
  OAI22X1 U3044 ( .A(n4623), .B(n5374), .C(n4639), .D(n5374), .Y(n5373) );
  OAI22X1 U3045 ( .A(n4626), .B(n4554), .C(n4624), .D(n4552), .Y(n5374) );
  XNOR2X1 U3046 ( .A(n5375), .B(n4641), .Y(n3458) );
  OAI21X1 U3047 ( .A(n4664), .B(n4695), .C(n5376), .Y(n5375) );
  OAI22X1 U3048 ( .A(n4625), .B(n5377), .C(n4639), .D(n5377), .Y(n5376) );
  OAI22X1 U3049 ( .A(n4628), .B(n4554), .C(n4552), .D(n4626), .Y(n5377) );
  XNOR2X1 U3050 ( .A(n5378), .B(n4641), .Y(n3457) );
  OAI21X1 U3051 ( .A(n4694), .B(n4664), .C(n5379), .Y(n5378) );
  OAI22X1 U3052 ( .A(n4627), .B(n5380), .C(n4639), .D(n5380), .Y(n5379) );
  OAI22X1 U3053 ( .A(n4630), .B(n4554), .C(n4628), .D(n4552), .Y(n5380) );
  XNOR2X1 U3054 ( .A(n5381), .B(n4641), .Y(n3456) );
  OAI21X1 U3055 ( .A(n4664), .B(n4693), .C(n5382), .Y(n5381) );
  OAI22X1 U3056 ( .A(n4629), .B(n5383), .C(n4639), .D(n5383), .Y(n5382) );
  OAI22X1 U3057 ( .A(n4630), .B(n4552), .C(n4632), .D(n4554), .Y(n5383) );
  XNOR2X1 U3058 ( .A(n5384), .B(n4641), .Y(n3455) );
  OAI21X1 U3059 ( .A(n4664), .B(n4690), .C(n5385), .Y(n5384) );
  OAI22X1 U3060 ( .A(n4631), .B(n5386), .C(n4639), .D(n5386), .Y(n5385) );
  NAND3X1 U3061 ( .A(n5388), .B(n5389), .C(n5390), .Y(n5387) );
  OAI22X1 U3062 ( .A(n4552), .B(n4632), .C(n4687), .D(n4554), .Y(n5386) );
  XNOR2X1 U3063 ( .A(a[15]), .B(a[16]), .Y(n5388) );
  XNOR2X1 U3064 ( .A(a[16]), .B(n4641), .Y(n5389) );
  XOR2X1 U3065 ( .A(a[15]), .B(n4645), .Y(n5390) );
  XOR2X1 U3066 ( .A(n5391), .B(n4678), .Y(n3453) );
  OAI22X1 U3067 ( .A(n4739), .B(n4686), .C(n4665), .D(n4686), .Y(n5391) );
  XOR2X1 U3068 ( .A(n5392), .B(n4678), .Y(n3452) );
  OAI21X1 U3069 ( .A(n4665), .B(n4725), .C(n5393), .Y(n5392) );
  AOI22X1 U3070 ( .A(n4680), .B(n5394), .C(n4683), .D(n5395), .Y(n5393) );
  XOR2X1 U3071 ( .A(n5396), .B(n4678), .Y(n3451) );
  OAI21X1 U3072 ( .A(n4665), .B(n4724), .C(n5397), .Y(n5396) );
  OAI22X1 U3073 ( .A(n4685), .B(n5398), .C(n4637), .D(n5398), .Y(n5397) );
  OAI22X1 U3074 ( .A(n4638), .B(n4681), .C(n4739), .D(n4568), .Y(n5398) );
  XOR2X1 U3075 ( .A(n5399), .B(n4678), .Y(n3450) );
  OAI21X1 U3076 ( .A(n4665), .B(n4723), .C(n5400), .Y(n5399) );
  OAI22X1 U3077 ( .A(n4680), .B(n5401), .C(n4637), .D(n5401), .Y(n5400) );
  OAI22X1 U3078 ( .A(n4638), .B(n4568), .C(n4739), .D(n4570), .Y(n5401) );
  XOR2X1 U3079 ( .A(n5402), .B(n4678), .Y(n3449) );
  OAI21X1 U3080 ( .A(n4665), .B(n4722), .C(n5403), .Y(n5402) );
  OAI22X1 U3081 ( .A(b[2]), .B(n5404), .C(n4637), .D(n5404), .Y(n5403) );
  OAI22X1 U3082 ( .A(n4638), .B(n4570), .C(n4739), .D(n4573), .Y(n5404) );
  XOR2X1 U3083 ( .A(n5405), .B(n4678), .Y(n3448) );
  OAI21X1 U3084 ( .A(n4665), .B(n4721), .C(n5406), .Y(n5405) );
  OAI22X1 U3085 ( .A(n4572), .B(n5407), .C(n4637), .D(n5407), .Y(n5406) );
  OAI22X1 U3086 ( .A(n4638), .B(n4573), .C(n4739), .D(n4575), .Y(n5407) );
  XOR2X1 U3087 ( .A(n5408), .B(n4678), .Y(n3447) );
  OAI21X1 U3088 ( .A(n4665), .B(n4720), .C(n5409), .Y(n5408) );
  OAI22X1 U3089 ( .A(b[4]), .B(n5410), .C(n4637), .D(n5410), .Y(n5409) );
  OAI22X1 U3090 ( .A(n4638), .B(n4575), .C(n4739), .D(n4578), .Y(n5410) );
  XOR2X1 U3091 ( .A(n5411), .B(n4678), .Y(n3446) );
  OAI21X1 U3092 ( .A(n4665), .B(n4719), .C(n5412), .Y(n5411) );
  OAI22X1 U3093 ( .A(n4577), .B(n5413), .C(n4637), .D(n5413), .Y(n5412) );
  OAI22X1 U3094 ( .A(n4638), .B(n4578), .C(n4739), .D(n4580), .Y(n5413) );
  XOR2X1 U3095 ( .A(n5414), .B(n4678), .Y(n3445) );
  OAI21X1 U3096 ( .A(n4665), .B(n4717), .C(n5415), .Y(n5414) );
  OAI22X1 U3097 ( .A(b[6]), .B(n5416), .C(n4637), .D(n5416), .Y(n5415) );
  OAI22X1 U3098 ( .A(n4638), .B(n4580), .C(n4739), .D(n4582), .Y(n5416) );
  XOR2X1 U3099 ( .A(n5417), .B(n4678), .Y(n3444) );
  OAI21X1 U3100 ( .A(n4665), .B(n4716), .C(n5418), .Y(n5417) );
  OAI22X1 U3101 ( .A(b[7]), .B(n5419), .C(n4637), .D(n5419), .Y(n5418) );
  OAI22X1 U3102 ( .A(n4638), .B(n4582), .C(n4739), .D(n4584), .Y(n5419) );
  XOR2X1 U3103 ( .A(n5420), .B(n4678), .Y(n3443) );
  OAI21X1 U3104 ( .A(n4665), .B(n4715), .C(n5421), .Y(n5420) );
  OAI22X1 U3105 ( .A(b[8]), .B(n5422), .C(n4637), .D(n5422), .Y(n5421) );
  OAI22X1 U3106 ( .A(n4638), .B(n4584), .C(n4739), .D(n4587), .Y(n5422) );
  XOR2X1 U3107 ( .A(n5423), .B(n4678), .Y(n3442) );
  OAI21X1 U3108 ( .A(n4665), .B(n4713), .C(n5424), .Y(n5423) );
  OAI22X1 U3109 ( .A(n4586), .B(n5425), .C(n4637), .D(n5425), .Y(n5424) );
  OAI22X1 U3110 ( .A(n4638), .B(n4587), .C(n4739), .D(n4589), .Y(n5425) );
  XOR2X1 U3111 ( .A(n5426), .B(n4678), .Y(n3441) );
  OAI21X1 U3112 ( .A(n4665), .B(n4712), .C(n5427), .Y(n5426) );
  OAI22X1 U3113 ( .A(b[10]), .B(n5428), .C(n4637), .D(n5428), .Y(n5427) );
  OAI22X1 U3114 ( .A(n4638), .B(n4589), .C(n4739), .D(n4592), .Y(n5428) );
  XOR2X1 U3115 ( .A(n5429), .B(n4678), .Y(n3440) );
  OAI21X1 U3116 ( .A(n4665), .B(n4711), .C(n5430), .Y(n5429) );
  OAI22X1 U3117 ( .A(n4591), .B(n5431), .C(n4637), .D(n5431), .Y(n5430) );
  OAI22X1 U3118 ( .A(n4638), .B(n4592), .C(n4739), .D(n4594), .Y(n5431) );
  XOR2X1 U3119 ( .A(n5432), .B(n4678), .Y(n3439) );
  OAI21X1 U3120 ( .A(n4665), .B(n4710), .C(n5433), .Y(n5432) );
  OAI22X1 U3121 ( .A(b[12]), .B(n5434), .C(n4637), .D(n5434), .Y(n5433) );
  OAI22X1 U3122 ( .A(n4638), .B(n4594), .C(n4739), .D(n4726), .Y(n5434) );
  XOR2X1 U3123 ( .A(n5435), .B(n4678), .Y(n3438) );
  OAI21X1 U3124 ( .A(n4665), .B(n4708), .C(n5436), .Y(n5435) );
  OAI22X1 U3125 ( .A(n4596), .B(n5437), .C(n4637), .D(n5437), .Y(n5436) );
  OAI22X1 U3126 ( .A(n4739), .B(n4599), .C(n4638), .D(n4726), .Y(n5437) );
  XOR2X1 U3127 ( .A(n5438), .B(n4678), .Y(n3437) );
  OAI21X1 U3128 ( .A(n4665), .B(n4707), .C(n5439), .Y(n5438) );
  OAI22X1 U3129 ( .A(b[14]), .B(n5440), .C(n4637), .D(n5440), .Y(n5439) );
  OAI22X1 U3130 ( .A(n4638), .B(n4599), .C(n4739), .D(n4601), .Y(n5440) );
  XOR2X1 U3131 ( .A(n5441), .B(n4678), .Y(n3436) );
  OAI21X1 U3132 ( .A(n4665), .B(n4706), .C(n5442), .Y(n5441) );
  OAI22X1 U3133 ( .A(n4600), .B(n5443), .C(n4637), .D(n5443), .Y(n5442) );
  OAI22X1 U3134 ( .A(n4739), .B(n4603), .C(n4638), .D(n4601), .Y(n5443) );
  XOR2X1 U3135 ( .A(n5444), .B(n4678), .Y(n3435) );
  OAI21X1 U3136 ( .A(n4665), .B(n4705), .C(n5445), .Y(n5444) );
  OAI22X1 U3137 ( .A(n4602), .B(n5446), .C(n4637), .D(n5446), .Y(n5445) );
  OAI22X1 U3138 ( .A(n4638), .B(n4603), .C(n4739), .D(n4606), .Y(n5446) );
  XOR2X1 U3139 ( .A(n5447), .B(n4678), .Y(n3434) );
  OAI21X1 U3140 ( .A(n4665), .B(n4704), .C(n5448), .Y(n5447) );
  OAI22X1 U3141 ( .A(n4605), .B(n5449), .C(n4637), .D(n5449), .Y(n5448) );
  OAI22X1 U3142 ( .A(n4638), .B(n4606), .C(n4739), .D(n4608), .Y(n5449) );
  XOR2X1 U3143 ( .A(n5450), .B(n2150), .Y(n3433) );
  OAI21X1 U3144 ( .A(n4665), .B(n4703), .C(n5451), .Y(n5450) );
  OAI22X1 U3145 ( .A(n4607), .B(n5452), .C(n4637), .D(n5452), .Y(n5451) );
  OAI22X1 U3146 ( .A(n4739), .B(n4611), .C(n4638), .D(n4608), .Y(n5452) );
  XOR2X1 U3147 ( .A(n5453), .B(n2150), .Y(n3432) );
  OAI21X1 U3148 ( .A(n4665), .B(n4702), .C(n5454), .Y(n5453) );
  OAI22X1 U3149 ( .A(n4610), .B(n5455), .C(n4637), .D(n5455), .Y(n5454) );
  OAI22X1 U3150 ( .A(n4638), .B(n4611), .C(n4739), .D(n4613), .Y(n5455) );
  XOR2X1 U3151 ( .A(n5456), .B(n2150), .Y(n3431) );
  OAI21X1 U3152 ( .A(n4665), .B(n4701), .C(n5457), .Y(n5456) );
  OAI22X1 U3153 ( .A(b[20]), .B(n5458), .C(n4637), .D(n5458), .Y(n5457) );
  OAI22X1 U3154 ( .A(n4638), .B(n4613), .C(n4739), .D(n4616), .Y(n5458) );
  XOR2X1 U3155 ( .A(n5459), .B(n2150), .Y(n3430) );
  OAI21X1 U3156 ( .A(n4665), .B(n4700), .C(n5460), .Y(n5459) );
  OAI22X1 U3157 ( .A(n4614), .B(n5461), .C(n4637), .D(n5461), .Y(n5460) );
  OAI22X1 U3158 ( .A(n4739), .B(n4618), .C(n4638), .D(n4616), .Y(n5461) );
  XOR2X1 U3159 ( .A(n5462), .B(n2150), .Y(n3429) );
  OAI21X1 U3160 ( .A(n4665), .B(n4699), .C(n5463), .Y(n5462) );
  OAI22X1 U3161 ( .A(n4617), .B(n5464), .C(n4637), .D(n5464), .Y(n5463) );
  OAI22X1 U3162 ( .A(n4638), .B(n4618), .C(n4739), .D(n4620), .Y(n5464) );
  XOR2X1 U3163 ( .A(n5465), .B(n2150), .Y(n3428) );
  OAI21X1 U3164 ( .A(n4665), .B(n4698), .C(n5466), .Y(n5465) );
  OAI22X1 U3165 ( .A(n4619), .B(n5467), .C(n4637), .D(n5467), .Y(n5466) );
  OAI22X1 U3166 ( .A(n4638), .B(n4620), .C(n4739), .D(n4622), .Y(n5467) );
  XOR2X1 U3167 ( .A(n5468), .B(n2150), .Y(n3427) );
  OAI21X1 U3168 ( .A(n4665), .B(n4697), .C(n5469), .Y(n5468) );
  OAI22X1 U3169 ( .A(n4621), .B(n5470), .C(n4637), .D(n5470), .Y(n5469) );
  OAI22X1 U3170 ( .A(n4739), .B(n4624), .C(n4638), .D(n4622), .Y(n5470) );
  XOR2X1 U3171 ( .A(n5471), .B(n2150), .Y(n3426) );
  OAI21X1 U3172 ( .A(n4665), .B(n4696), .C(n5472), .Y(n5471) );
  OAI22X1 U3173 ( .A(n4623), .B(n5473), .C(n4637), .D(n5473), .Y(n5472) );
  OAI22X1 U3174 ( .A(n4638), .B(n4624), .C(n4739), .D(n4626), .Y(n5473) );
  XOR2X1 U3175 ( .A(n5474), .B(n2150), .Y(n3425) );
  OAI21X1 U3176 ( .A(n4665), .B(n4695), .C(n5475), .Y(n5474) );
  OAI22X1 U3177 ( .A(n4625), .B(n5476), .C(n4637), .D(n5476), .Y(n5475) );
  NAND3X1 U3178 ( .A(n5478), .B(n5479), .C(n5480), .Y(n5477) );
  OAI22X1 U3179 ( .A(n4638), .B(n4626), .C(n4628), .D(n4739), .Y(n5476) );
  NOR2X1 U3180 ( .A(n5479), .B(n5478), .Y(n5394) );
  NOR2X1 U3181 ( .A(n4740), .B(n5480), .Y(n5395) );
  XNOR2X1 U3182 ( .A(a[18]), .B(a[19]), .Y(n5480) );
  XOR2X1 U3183 ( .A(a[19]), .B(n2150), .Y(n5479) );
  XOR2X1 U3184 ( .A(a[18]), .B(n4641), .Y(n5478) );
  XOR2X1 U3185 ( .A(n4676), .B(n5481), .Y(n3423) );
  OAI22X1 U3186 ( .A(n4686), .B(n4555), .C(n4686), .D(n4634), .Y(n5481) );
  XOR2X1 U3187 ( .A(n5482), .B(n4676), .Y(n3422) );
  OAI21X1 U3188 ( .A(n4555), .B(n4725), .C(n5483), .Y(n5482) );
  AOI22X1 U3189 ( .A(n4680), .B(n5484), .C(n4683), .D(n5485), .Y(n5483) );
  XOR2X1 U3190 ( .A(n5486), .B(n4676), .Y(n3421) );
  OAI21X1 U3191 ( .A(n4555), .B(n4724), .C(n5487), .Y(n5486) );
  OAI22X1 U3192 ( .A(n4685), .B(n5488), .C(n4635), .D(n5488), .Y(n5487) );
  OAI22X1 U3193 ( .A(n4636), .B(n4681), .C(n4634), .D(n4568), .Y(n5488) );
  XOR2X1 U3194 ( .A(n5489), .B(n4676), .Y(n3420) );
  OAI21X1 U3195 ( .A(n4555), .B(n4723), .C(n5490), .Y(n5489) );
  OAI22X1 U3196 ( .A(n4680), .B(n5491), .C(n4635), .D(n5491), .Y(n5490) );
  OAI22X1 U3197 ( .A(n4636), .B(n4568), .C(n4634), .D(n4570), .Y(n5491) );
  XOR2X1 U3198 ( .A(n5492), .B(n4676), .Y(n3419) );
  OAI21X1 U3199 ( .A(n4555), .B(n4722), .C(n5493), .Y(n5492) );
  OAI22X1 U3200 ( .A(n4569), .B(n5494), .C(n4635), .D(n5494), .Y(n5493) );
  OAI22X1 U3201 ( .A(n4636), .B(n4570), .C(n4634), .D(n4573), .Y(n5494) );
  XOR2X1 U3202 ( .A(n5495), .B(n4676), .Y(n3418) );
  OAI21X1 U3203 ( .A(n4555), .B(n4721), .C(n5496), .Y(n5495) );
  OAI22X1 U3204 ( .A(n4571), .B(n5497), .C(n4635), .D(n5497), .Y(n5496) );
  OAI22X1 U3205 ( .A(n4636), .B(n4573), .C(n4634), .D(n4575), .Y(n5497) );
  XOR2X1 U3206 ( .A(n5498), .B(n4676), .Y(n3417) );
  OAI21X1 U3207 ( .A(n4555), .B(n4720), .C(n5499), .Y(n5498) );
  OAI22X1 U3208 ( .A(n4574), .B(n5500), .C(n4635), .D(n5500), .Y(n5499) );
  OAI22X1 U3209 ( .A(n4636), .B(n4575), .C(n4634), .D(n4578), .Y(n5500) );
  XOR2X1 U3210 ( .A(n5501), .B(n4676), .Y(n3416) );
  OAI21X1 U3211 ( .A(n4555), .B(n4719), .C(n5502), .Y(n5501) );
  OAI22X1 U3212 ( .A(n4576), .B(n5503), .C(n4635), .D(n5503), .Y(n5502) );
  OAI22X1 U3213 ( .A(n4636), .B(n4578), .C(n4634), .D(n4580), .Y(n5503) );
  XOR2X1 U3214 ( .A(n5504), .B(n4676), .Y(n3415) );
  OAI21X1 U3215 ( .A(n4555), .B(n4717), .C(n5505), .Y(n5504) );
  OAI22X1 U3216 ( .A(n4579), .B(n5506), .C(n4635), .D(n5506), .Y(n5505) );
  OAI22X1 U3217 ( .A(n4636), .B(n4580), .C(n4634), .D(n4582), .Y(n5506) );
  XOR2X1 U3218 ( .A(n5507), .B(n4676), .Y(n3414) );
  OAI21X1 U3219 ( .A(n4555), .B(n4716), .C(n5508), .Y(n5507) );
  OAI22X1 U3220 ( .A(n4581), .B(n5509), .C(n4635), .D(n5509), .Y(n5508) );
  OAI22X1 U3221 ( .A(n4636), .B(n4582), .C(n4634), .D(n4584), .Y(n5509) );
  XOR2X1 U3222 ( .A(n5510), .B(n4676), .Y(n3413) );
  OAI21X1 U3223 ( .A(n4555), .B(n4715), .C(n5511), .Y(n5510) );
  OAI22X1 U3224 ( .A(n4583), .B(n5512), .C(n4635), .D(n5512), .Y(n5511) );
  OAI22X1 U3225 ( .A(n4636), .B(n4584), .C(n4634), .D(n4587), .Y(n5512) );
  XOR2X1 U3226 ( .A(n5513), .B(n4676), .Y(n3412) );
  OAI21X1 U3227 ( .A(n4555), .B(n4713), .C(n5514), .Y(n5513) );
  OAI22X1 U3228 ( .A(n4585), .B(n5515), .C(n4635), .D(n5515), .Y(n5514) );
  OAI22X1 U3229 ( .A(n4636), .B(n4587), .C(n4634), .D(n4589), .Y(n5515) );
  XOR2X1 U3230 ( .A(n5516), .B(n4676), .Y(n3411) );
  OAI21X1 U3231 ( .A(n4555), .B(n4712), .C(n5517), .Y(n5516) );
  OAI22X1 U3232 ( .A(n4588), .B(n5518), .C(n4635), .D(n5518), .Y(n5517) );
  OAI22X1 U3233 ( .A(n4636), .B(n4589), .C(n4634), .D(n4592), .Y(n5518) );
  XOR2X1 U3234 ( .A(n5519), .B(n4676), .Y(n3410) );
  OAI21X1 U3235 ( .A(n4555), .B(n4711), .C(n5520), .Y(n5519) );
  OAI22X1 U3236 ( .A(n4590), .B(n5521), .C(n4635), .D(n5521), .Y(n5520) );
  OAI22X1 U3237 ( .A(n4636), .B(n4592), .C(n4634), .D(n4594), .Y(n5521) );
  XOR2X1 U3238 ( .A(n5522), .B(n4676), .Y(n3409) );
  OAI21X1 U3239 ( .A(n4555), .B(n4710), .C(n5523), .Y(n5522) );
  OAI22X1 U3240 ( .A(n4593), .B(n5524), .C(n4635), .D(n5524), .Y(n5523) );
  OAI22X1 U3241 ( .A(n4636), .B(n4594), .C(n4634), .D(n4726), .Y(n5524) );
  XOR2X1 U3242 ( .A(n5525), .B(n4676), .Y(n3408) );
  OAI21X1 U3243 ( .A(n4555), .B(n4708), .C(n5526), .Y(n5525) );
  OAI22X1 U3244 ( .A(n4595), .B(n5527), .C(n4635), .D(n5527), .Y(n5526) );
  OAI22X1 U3245 ( .A(n4634), .B(n4599), .C(n4636), .D(n4726), .Y(n5527) );
  XOR2X1 U3246 ( .A(n5528), .B(n4676), .Y(n3407) );
  OAI21X1 U3247 ( .A(n4555), .B(n4707), .C(n5529), .Y(n5528) );
  OAI22X1 U3248 ( .A(n4598), .B(n5530), .C(n4635), .D(n5530), .Y(n5529) );
  OAI22X1 U3249 ( .A(n4636), .B(n4599), .C(n4634), .D(n4601), .Y(n5530) );
  XOR2X1 U3250 ( .A(n5531), .B(n4676), .Y(n3406) );
  OAI21X1 U3251 ( .A(n4555), .B(n4706), .C(n5532), .Y(n5531) );
  OAI22X1 U3252 ( .A(b[15]), .B(n5533), .C(n4635), .D(n5533), .Y(n5532) );
  OAI22X1 U3253 ( .A(n4634), .B(n4603), .C(n4636), .D(n4601), .Y(n5533) );
  XOR2X1 U3254 ( .A(n5534), .B(n4676), .Y(n3405) );
  OAI21X1 U3255 ( .A(n4555), .B(n4705), .C(n5535), .Y(n5534) );
  OAI22X1 U3256 ( .A(n4602), .B(n5536), .C(n4635), .D(n5536), .Y(n5535) );
  OAI22X1 U3257 ( .A(n4636), .B(n4603), .C(n4634), .D(n4606), .Y(n5536) );
  XOR2X1 U3258 ( .A(n5537), .B(n4676), .Y(n3404) );
  OAI21X1 U3259 ( .A(n4555), .B(n4704), .C(n5538), .Y(n5537) );
  OAI22X1 U3260 ( .A(n4605), .B(n5539), .C(n4635), .D(n5539), .Y(n5538) );
  OAI22X1 U3261 ( .A(n4636), .B(n4606), .C(n4634), .D(n4608), .Y(n5539) );
  XOR2X1 U3262 ( .A(n5540), .B(n2153), .Y(n3403) );
  OAI21X1 U3263 ( .A(n4555), .B(n4703), .C(n5541), .Y(n5540) );
  OAI22X1 U3264 ( .A(n4607), .B(n5542), .C(n4635), .D(n5542), .Y(n5541) );
  OAI22X1 U3265 ( .A(n4634), .B(n4611), .C(n4636), .D(n4608), .Y(n5542) );
  XOR2X1 U3266 ( .A(n5543), .B(n2153), .Y(n3402) );
  OAI21X1 U3267 ( .A(n4555), .B(n4702), .C(n5544), .Y(n5543) );
  OAI22X1 U3268 ( .A(n4609), .B(n5545), .C(n4635), .D(n5545), .Y(n5544) );
  OAI22X1 U3269 ( .A(n4636), .B(n4611), .C(n4634), .D(n4613), .Y(n5545) );
  XOR2X1 U3270 ( .A(n5546), .B(n2153), .Y(n3401) );
  OAI21X1 U3271 ( .A(n4555), .B(n4701), .C(n5547), .Y(n5546) );
  OAI22X1 U3272 ( .A(n4612), .B(n5548), .C(n4635), .D(n5548), .Y(n5547) );
  OAI22X1 U3273 ( .A(n4636), .B(n4613), .C(n4634), .D(n4616), .Y(n5548) );
  XOR2X1 U3274 ( .A(n5549), .B(n2153), .Y(n3400) );
  OAI21X1 U3275 ( .A(n4555), .B(n4700), .C(n5550), .Y(n5549) );
  OAI22X1 U3276 ( .A(n4615), .B(n5551), .C(n4635), .D(n5551), .Y(n5550) );
  OAI22X1 U3277 ( .A(n4634), .B(n4618), .C(n4636), .D(n4616), .Y(n5551) );
  XOR2X1 U3278 ( .A(n5552), .B(n2153), .Y(n3399) );
  OAI21X1 U3279 ( .A(n4555), .B(n4699), .C(n5553), .Y(n5552) );
  OAI22X1 U3280 ( .A(n4617), .B(n5554), .C(n4635), .D(n5554), .Y(n5553) );
  OAI22X1 U3281 ( .A(n4636), .B(n4618), .C(n4634), .D(n4620), .Y(n5554) );
  XOR2X1 U3282 ( .A(n5555), .B(n2153), .Y(n3398) );
  OAI21X1 U3283 ( .A(n4555), .B(n4698), .C(n5556), .Y(n5555) );
  OAI22X1 U3284 ( .A(n4619), .B(n5557), .C(n4635), .D(n5557), .Y(n5556) );
  NAND3X1 U3285 ( .A(n4738), .B(n5559), .C(n5560), .Y(n5558) );
  OAI22X1 U3286 ( .A(n4636), .B(n4620), .C(n4622), .D(n4634), .Y(n5557) );
  NOR2X1 U3287 ( .A(n5559), .B(n4738), .Y(n5484) );
  NOR2X1 U3288 ( .A(n5561), .B(n5560), .Y(n5485) );
  XNOR2X1 U3289 ( .A(a[21]), .B(a[22]), .Y(n5560) );
  XOR2X1 U3290 ( .A(a[22]), .B(n2153), .Y(n5559) );
  XOR2X1 U3291 ( .A(a[21]), .B(n2150), .Y(n5561) );
  XOR2X1 U3292 ( .A(n4674), .B(n5562), .Y(n3396) );
  OAI22X1 U3293 ( .A(n4686), .B(n4556), .C(n4686), .D(n4735), .Y(n5562) );
  XOR2X1 U3294 ( .A(n5563), .B(n2156), .Y(n3395) );
  OAI21X1 U3295 ( .A(n4556), .B(n4725), .C(n5564), .Y(n5563) );
  AOI22X1 U3296 ( .A(n4680), .B(n5565), .C(n4683), .D(n5566), .Y(n5564) );
  XOR2X1 U3297 ( .A(n5567), .B(n2156), .Y(n3394) );
  OAI21X1 U3298 ( .A(n4556), .B(n4724), .C(n5568), .Y(n5567) );
  OAI22X1 U3299 ( .A(n4685), .B(n5569), .C(n4567), .D(n5569), .Y(n5568) );
  OAI22X1 U3300 ( .A(n4736), .B(n4681), .C(n4735), .D(n4568), .Y(n5569) );
  XOR2X1 U3301 ( .A(n5570), .B(n2156), .Y(n3393) );
  OAI21X1 U3302 ( .A(n4556), .B(n4723), .C(n5571), .Y(n5570) );
  OAI22X1 U3303 ( .A(n4680), .B(n5572), .C(n4567), .D(n5572), .Y(n5571) );
  OAI22X1 U3304 ( .A(n4736), .B(n4568), .C(n4735), .D(n4570), .Y(n5572) );
  XOR2X1 U3305 ( .A(n5573), .B(n2156), .Y(n3392) );
  OAI21X1 U3306 ( .A(n4556), .B(n4722), .C(n5574), .Y(n5573) );
  OAI22X1 U3307 ( .A(b[2]), .B(n5575), .C(n4567), .D(n5575), .Y(n5574) );
  OAI22X1 U3308 ( .A(n4736), .B(n4570), .C(n4735), .D(n4573), .Y(n5575) );
  XOR2X1 U3309 ( .A(n5576), .B(n2156), .Y(n3391) );
  OAI21X1 U3310 ( .A(n4556), .B(n4721), .C(n5577), .Y(n5576) );
  OAI22X1 U3311 ( .A(n4572), .B(n5578), .C(n4567), .D(n5578), .Y(n5577) );
  OAI22X1 U3312 ( .A(n4736), .B(n4573), .C(n4735), .D(n4575), .Y(n5578) );
  XOR2X1 U3313 ( .A(n5579), .B(n2156), .Y(n3390) );
  OAI21X1 U3314 ( .A(n4556), .B(n4720), .C(n5580), .Y(n5579) );
  OAI22X1 U3315 ( .A(b[4]), .B(n5581), .C(n4567), .D(n5581), .Y(n5580) );
  OAI22X1 U3316 ( .A(n4736), .B(n4575), .C(n4735), .D(n4578), .Y(n5581) );
  XOR2X1 U3317 ( .A(n5582), .B(n2156), .Y(n3389) );
  OAI21X1 U3318 ( .A(n4556), .B(n4719), .C(n5583), .Y(n5582) );
  OAI22X1 U3319 ( .A(n4577), .B(n5584), .C(n4567), .D(n5584), .Y(n5583) );
  OAI22X1 U3320 ( .A(n4736), .B(n4578), .C(n4735), .D(n4580), .Y(n5584) );
  XOR2X1 U3321 ( .A(n5585), .B(n2156), .Y(n3388) );
  OAI21X1 U3322 ( .A(n4556), .B(n4717), .C(n5586), .Y(n5585) );
  OAI22X1 U3323 ( .A(b[6]), .B(n5587), .C(n4567), .D(n5587), .Y(n5586) );
  OAI22X1 U3324 ( .A(n4736), .B(n4580), .C(n4735), .D(n4582), .Y(n5587) );
  XOR2X1 U3325 ( .A(n5588), .B(n2156), .Y(n3387) );
  OAI21X1 U3326 ( .A(n4556), .B(n4716), .C(n5589), .Y(n5588) );
  OAI22X1 U3327 ( .A(b[7]), .B(n5590), .C(n4567), .D(n5590), .Y(n5589) );
  OAI22X1 U3328 ( .A(n4736), .B(n4582), .C(n4735), .D(n4584), .Y(n5590) );
  XOR2X1 U3329 ( .A(n5591), .B(n2156), .Y(n3386) );
  OAI21X1 U3330 ( .A(n4556), .B(n4715), .C(n5592), .Y(n5591) );
  OAI22X1 U3331 ( .A(b[8]), .B(n5593), .C(n4567), .D(n5593), .Y(n5592) );
  OAI22X1 U3332 ( .A(n4736), .B(n4584), .C(n4735), .D(n4587), .Y(n5593) );
  XOR2X1 U3333 ( .A(n5594), .B(n4674), .Y(n3385) );
  OAI21X1 U3334 ( .A(n4556), .B(n4713), .C(n5595), .Y(n5594) );
  OAI22X1 U3335 ( .A(n4586), .B(n5596), .C(n4567), .D(n5596), .Y(n5595) );
  OAI22X1 U3336 ( .A(n4736), .B(n4587), .C(n4735), .D(n4589), .Y(n5596) );
  XOR2X1 U3337 ( .A(n5597), .B(n4674), .Y(n3384) );
  OAI21X1 U3338 ( .A(n4556), .B(n4712), .C(n5598), .Y(n5597) );
  OAI22X1 U3339 ( .A(b[10]), .B(n5599), .C(n4567), .D(n5599), .Y(n5598) );
  OAI22X1 U3340 ( .A(n4736), .B(n4589), .C(n4735), .D(n4592), .Y(n5599) );
  XOR2X1 U3341 ( .A(n5600), .B(n4674), .Y(n3383) );
  OAI21X1 U3342 ( .A(n4556), .B(n4711), .C(n5601), .Y(n5600) );
  OAI22X1 U3343 ( .A(n4591), .B(n5602), .C(n4567), .D(n5602), .Y(n5601) );
  OAI22X1 U3344 ( .A(n4736), .B(n4592), .C(n4735), .D(n4594), .Y(n5602) );
  XOR2X1 U3345 ( .A(n5603), .B(n4674), .Y(n3382) );
  OAI21X1 U3346 ( .A(n4556), .B(n4710), .C(n5604), .Y(n5603) );
  OAI22X1 U3347 ( .A(b[12]), .B(n5605), .C(n4567), .D(n5605), .Y(n5604) );
  OAI22X1 U3348 ( .A(n4736), .B(n4594), .C(n4735), .D(n4726), .Y(n5605) );
  XOR2X1 U3349 ( .A(n5606), .B(n4674), .Y(n3381) );
  OAI21X1 U3350 ( .A(n4556), .B(n4708), .C(n5607), .Y(n5606) );
  OAI22X1 U3351 ( .A(n4596), .B(n5608), .C(n4567), .D(n5608), .Y(n5607) );
  OAI22X1 U3352 ( .A(n4735), .B(n4599), .C(n4736), .D(n4726), .Y(n5608) );
  XOR2X1 U3353 ( .A(n5609), .B(n4674), .Y(n3380) );
  OAI21X1 U3354 ( .A(n4556), .B(n4707), .C(n5610), .Y(n5609) );
  OAI22X1 U3355 ( .A(b[14]), .B(n5611), .C(n4567), .D(n5611), .Y(n5610) );
  OAI22X1 U3356 ( .A(n4736), .B(n4599), .C(n4735), .D(n4601), .Y(n5611) );
  XOR2X1 U3357 ( .A(n5612), .B(n4674), .Y(n3379) );
  OAI21X1 U3358 ( .A(n4556), .B(n4706), .C(n5613), .Y(n5612) );
  OAI22X1 U3359 ( .A(n4600), .B(n5614), .C(n4567), .D(n5614), .Y(n5613) );
  OAI22X1 U3360 ( .A(n4735), .B(n4603), .C(n4736), .D(n4601), .Y(n5614) );
  XOR2X1 U3361 ( .A(n5615), .B(n2156), .Y(n3378) );
  OAI21X1 U3362 ( .A(n4556), .B(n4705), .C(n5616), .Y(n5615) );
  OAI22X1 U3363 ( .A(n4602), .B(n5617), .C(n4567), .D(n5617), .Y(n5616) );
  OAI22X1 U3364 ( .A(n4736), .B(n4603), .C(n4735), .D(n4606), .Y(n5617) );
  XOR2X1 U3365 ( .A(n5618), .B(n4674), .Y(n3377) );
  OAI21X1 U3366 ( .A(n4556), .B(n4704), .C(n5619), .Y(n5618) );
  OAI22X1 U3367 ( .A(n4605), .B(n5620), .C(n4567), .D(n5620), .Y(n5619) );
  OAI22X1 U3368 ( .A(n4736), .B(n4606), .C(n4735), .D(n4608), .Y(n5620) );
  XOR2X1 U3369 ( .A(n5621), .B(n4674), .Y(n3376) );
  OAI21X1 U3370 ( .A(n4556), .B(n4703), .C(n5622), .Y(n5621) );
  OAI22X1 U3371 ( .A(n4607), .B(n5623), .C(n4567), .D(n5623), .Y(n5622) );
  OAI22X1 U3372 ( .A(n4735), .B(n4611), .C(n4736), .D(n4608), .Y(n5623) );
  XOR2X1 U3373 ( .A(n5624), .B(n4674), .Y(n3375) );
  OAI21X1 U3374 ( .A(n4556), .B(n4702), .C(n5625), .Y(n5624) );
  OAI22X1 U3375 ( .A(n4610), .B(n5626), .C(n4567), .D(n5626), .Y(n5625) );
  OAI22X1 U3376 ( .A(n4736), .B(n4611), .C(n4735), .D(n4613), .Y(n5626) );
  XOR2X1 U3377 ( .A(n5627), .B(n4674), .Y(n3374) );
  OAI21X1 U3378 ( .A(n4556), .B(n4701), .C(n5628), .Y(n5627) );
  OAI22X1 U3379 ( .A(b[20]), .B(n5629), .C(n4567), .D(n5629), .Y(n5628) );
  NAND3X1 U3380 ( .A(n5631), .B(n5632), .C(n5633), .Y(n5630) );
  OAI22X1 U3381 ( .A(n4736), .B(n4613), .C(n4616), .D(n4735), .Y(n5629) );
  NOR2X1 U3382 ( .A(n5632), .B(n5631), .Y(n5565) );
  NOR2X1 U3383 ( .A(n4737), .B(n5633), .Y(n5566) );
  XNOR2X1 U3384 ( .A(a[24]), .B(a[25]), .Y(n5633) );
  XOR2X1 U3385 ( .A(a[25]), .B(n4674), .Y(n5632) );
  XNOR2X1 U3386 ( .A(a[24]), .B(n2153), .Y(n5631) );
  XOR2X1 U3387 ( .A(n4672), .B(n5634), .Y(n3372) );
  OAI22X1 U3388 ( .A(n4686), .B(n4557), .C(n4686), .D(n4731), .Y(n5634) );
  XOR2X1 U3389 ( .A(n5635), .B(n2159), .Y(n3371) );
  OAI21X1 U3390 ( .A(n4557), .B(n4725), .C(n5636), .Y(n5635) );
  AOI22X1 U3391 ( .A(n4680), .B(n5637), .C(n4682), .D(n5638), .Y(n5636) );
  XOR2X1 U3392 ( .A(n5639), .B(n2159), .Y(n3370) );
  OAI21X1 U3393 ( .A(n4557), .B(n4724), .C(n5640), .Y(n5639) );
  OAI22X1 U3394 ( .A(n4685), .B(n5641), .C(n4732), .D(n5641), .Y(n5640) );
  OAI22X1 U3395 ( .A(n4733), .B(n4681), .C(n4731), .D(n4568), .Y(n5641) );
  XOR2X1 U3396 ( .A(n5642), .B(n2159), .Y(n3369) );
  OAI21X1 U3397 ( .A(n4557), .B(n4723), .C(n5643), .Y(n5642) );
  OAI22X1 U3398 ( .A(n4680), .B(n5644), .C(n4732), .D(n5644), .Y(n5643) );
  OAI22X1 U3399 ( .A(n4733), .B(n4568), .C(n4731), .D(n4570), .Y(n5644) );
  XOR2X1 U3400 ( .A(n5645), .B(n2159), .Y(n3368) );
  OAI21X1 U3401 ( .A(n4557), .B(n4722), .C(n5646), .Y(n5645) );
  OAI22X1 U3402 ( .A(n4569), .B(n5647), .C(n4732), .D(n5647), .Y(n5646) );
  OAI22X1 U3403 ( .A(n4733), .B(n4570), .C(n4731), .D(n4573), .Y(n5647) );
  XOR2X1 U3404 ( .A(n5648), .B(n2159), .Y(n3367) );
  OAI21X1 U3405 ( .A(n4557), .B(n4721), .C(n5649), .Y(n5648) );
  OAI22X1 U3406 ( .A(n4571), .B(n5650), .C(n4732), .D(n5650), .Y(n5649) );
  OAI22X1 U3407 ( .A(n4733), .B(n4573), .C(n4731), .D(n4575), .Y(n5650) );
  XOR2X1 U3408 ( .A(n5651), .B(n2159), .Y(n3366) );
  OAI21X1 U3409 ( .A(n4557), .B(n4720), .C(n5652), .Y(n5651) );
  OAI22X1 U3410 ( .A(n4574), .B(n5653), .C(n4732), .D(n5653), .Y(n5652) );
  OAI22X1 U3411 ( .A(n4733), .B(n4575), .C(n4731), .D(n4578), .Y(n5653) );
  XOR2X1 U3412 ( .A(n5654), .B(n2159), .Y(n3365) );
  OAI21X1 U3413 ( .A(n4557), .B(n4719), .C(n5655), .Y(n5654) );
  OAI22X1 U3414 ( .A(n4576), .B(n5656), .C(n4732), .D(n5656), .Y(n5655) );
  OAI22X1 U3415 ( .A(n4733), .B(n4578), .C(n4731), .D(n4580), .Y(n5656) );
  XOR2X1 U3416 ( .A(n5657), .B(n2159), .Y(n3364) );
  OAI21X1 U3417 ( .A(n4557), .B(n4717), .C(n5658), .Y(n5657) );
  OAI22X1 U3418 ( .A(n4579), .B(n5659), .C(n4732), .D(n5659), .Y(n5658) );
  OAI22X1 U3419 ( .A(n4733), .B(n4580), .C(n4731), .D(n4582), .Y(n5659) );
  XOR2X1 U3420 ( .A(n5660), .B(n4672), .Y(n3363) );
  OAI21X1 U3421 ( .A(n4557), .B(n4716), .C(n5661), .Y(n5660) );
  OAI22X1 U3422 ( .A(n4581), .B(n5662), .C(n4732), .D(n5662), .Y(n5661) );
  OAI22X1 U3423 ( .A(n4733), .B(n4582), .C(n4731), .D(n4584), .Y(n5662) );
  XOR2X1 U3424 ( .A(n5663), .B(n4672), .Y(n3362) );
  OAI21X1 U3425 ( .A(n4557), .B(n4715), .C(n5664), .Y(n5663) );
  OAI22X1 U3426 ( .A(n4583), .B(n5665), .C(n4732), .D(n5665), .Y(n5664) );
  OAI22X1 U3427 ( .A(n4733), .B(n4584), .C(n4731), .D(n4587), .Y(n5665) );
  XOR2X1 U3428 ( .A(n5666), .B(n4672), .Y(n3361) );
  OAI21X1 U3429 ( .A(n4557), .B(n4713), .C(n5667), .Y(n5666) );
  OAI22X1 U3430 ( .A(n4585), .B(n5668), .C(n4732), .D(n5668), .Y(n5667) );
  OAI22X1 U3431 ( .A(n4733), .B(n4587), .C(n4731), .D(n4589), .Y(n5668) );
  XOR2X1 U3432 ( .A(n5669), .B(n4672), .Y(n3360) );
  OAI21X1 U3433 ( .A(n4557), .B(n4712), .C(n5670), .Y(n5669) );
  OAI22X1 U3434 ( .A(n4588), .B(n5671), .C(n4732), .D(n5671), .Y(n5670) );
  OAI22X1 U3435 ( .A(n4733), .B(n4589), .C(n4731), .D(n4592), .Y(n5671) );
  XOR2X1 U3436 ( .A(n5672), .B(n4672), .Y(n3359) );
  OAI21X1 U3437 ( .A(n4557), .B(n4711), .C(n5673), .Y(n5672) );
  OAI22X1 U3438 ( .A(n4590), .B(n5674), .C(n4732), .D(n5674), .Y(n5673) );
  OAI22X1 U3439 ( .A(n4733), .B(n4592), .C(n4731), .D(n4594), .Y(n5674) );
  XOR2X1 U3440 ( .A(n5675), .B(n4672), .Y(n3358) );
  OAI21X1 U3441 ( .A(n4557), .B(n4710), .C(n5676), .Y(n5675) );
  OAI22X1 U3442 ( .A(n4593), .B(n5677), .C(n4732), .D(n5677), .Y(n5676) );
  OAI22X1 U3443 ( .A(n4733), .B(n4594), .C(n4731), .D(n4726), .Y(n5677) );
  XOR2X1 U3444 ( .A(n5678), .B(n4672), .Y(n3357) );
  OAI21X1 U3445 ( .A(n4557), .B(n4708), .C(n5679), .Y(n5678) );
  OAI22X1 U3446 ( .A(n4595), .B(n5680), .C(n4732), .D(n5680), .Y(n5679) );
  OAI22X1 U3447 ( .A(n4731), .B(n4599), .C(n4733), .D(n4726), .Y(n5680) );
  XOR2X1 U3448 ( .A(n5681), .B(n4672), .Y(n3356) );
  OAI21X1 U3449 ( .A(n4557), .B(n4707), .C(n5682), .Y(n5681) );
  OAI22X1 U3450 ( .A(n4598), .B(n5683), .C(n4732), .D(n5683), .Y(n5682) );
  OAI22X1 U3451 ( .A(n4733), .B(n4599), .C(n4731), .D(n4601), .Y(n5683) );
  XOR2X1 U3452 ( .A(n5684), .B(n4672), .Y(n3355) );
  OAI21X1 U3453 ( .A(n4557), .B(n4706), .C(n5685), .Y(n5684) );
  OAI22X1 U3454 ( .A(b[15]), .B(n5686), .C(n4732), .D(n5686), .Y(n5685) );
  OAI22X1 U3455 ( .A(n4731), .B(n4603), .C(n4733), .D(n4601), .Y(n5686) );
  XOR2X1 U3456 ( .A(n5687), .B(n4672), .Y(n3354) );
  OAI21X1 U3457 ( .A(n4557), .B(n4705), .C(n5688), .Y(n5687) );
  OAI22X1 U3458 ( .A(n4602), .B(n5689), .C(n4732), .D(n5689), .Y(n5688) );
  OAI22X1 U3459 ( .A(n4733), .B(n4603), .C(n4731), .D(n4606), .Y(n5689) );
  XOR2X1 U3460 ( .A(n5690), .B(n4672), .Y(n3353) );
  OAI21X1 U3461 ( .A(n4557), .B(n4704), .C(n5691), .Y(n5690) );
  OAI22X1 U3462 ( .A(n4605), .B(n5692), .C(n4732), .D(n5692), .Y(n5691) );
  NAND3X1 U3463 ( .A(n5694), .B(n5695), .C(n5696), .Y(n5693) );
  OAI22X1 U3464 ( .A(n4733), .B(n4606), .C(n4608), .D(n4731), .Y(n5692) );
  NOR2X1 U3465 ( .A(n5695), .B(n5694), .Y(n5637) );
  NOR2X1 U3466 ( .A(n4734), .B(n5696), .Y(n5638) );
  XNOR2X1 U3467 ( .A(a[27]), .B(a[28]), .Y(n5696) );
  XOR2X1 U3468 ( .A(a[28]), .B(n4672), .Y(n5695) );
  XNOR2X1 U3469 ( .A(a[27]), .B(n4674), .Y(n5694) );
  OAI22X1 U3470 ( .A(n4728), .B(n4686), .C(n4558), .D(n4686), .Y(n3351) );
  OAI21X1 U3471 ( .A(n4558), .B(n4725), .C(n5697), .Y(n3350) );
  AOI22X1 U3472 ( .A(n4680), .B(n5698), .C(n4682), .D(n5699), .Y(n5697) );
  OAI21X1 U3473 ( .A(n4558), .B(n4724), .C(n5700), .Y(n3349) );
  OAI22X1 U3474 ( .A(n4684), .B(n5701), .C(n4727), .D(n5701), .Y(n5700) );
  OAI22X1 U3475 ( .A(n4729), .B(n4681), .C(n4728), .D(n4568), .Y(n5701) );
  OAI21X1 U3476 ( .A(n4558), .B(n4723), .C(n5702), .Y(n3348) );
  OAI22X1 U3477 ( .A(n4680), .B(n5703), .C(n4727), .D(n5703), .Y(n5702) );
  OAI22X1 U3478 ( .A(n4729), .B(n4568), .C(n4728), .D(n4570), .Y(n5703) );
  OAI21X1 U3479 ( .A(n4558), .B(n4722), .C(n5704), .Y(n3347) );
  OAI22X1 U3480 ( .A(b[2]), .B(n5705), .C(n4727), .D(n5705), .Y(n5704) );
  OAI22X1 U3481 ( .A(n4729), .B(n4570), .C(n4728), .D(n4573), .Y(n5705) );
  OAI21X1 U3482 ( .A(n4558), .B(n4721), .C(n5706), .Y(n3346) );
  OAI22X1 U3483 ( .A(n4572), .B(n5707), .C(n4727), .D(n5707), .Y(n5706) );
  OAI22X1 U3484 ( .A(n4729), .B(n4573), .C(n4728), .D(n4575), .Y(n5707) );
  OAI21X1 U3485 ( .A(n4558), .B(n4720), .C(n5708), .Y(n3345) );
  OAI22X1 U3486 ( .A(b[4]), .B(n5709), .C(n4727), .D(n5709), .Y(n5708) );
  OAI22X1 U3487 ( .A(n4729), .B(n4575), .C(n4728), .D(n4578), .Y(n5709) );
  OAI21X1 U3488 ( .A(n4558), .B(n4719), .C(n5710), .Y(n3344) );
  OAI22X1 U3489 ( .A(n4577), .B(n5711), .C(n4727), .D(n5711), .Y(n5710) );
  OAI22X1 U3490 ( .A(n4729), .B(n4578), .C(n4728), .D(n4580), .Y(n5711) );
  OAI21X1 U3491 ( .A(n4558), .B(n4717), .C(n5712), .Y(n3343) );
  OAI22X1 U3492 ( .A(b[6]), .B(n5713), .C(n4727), .D(n5713), .Y(n5712) );
  OAI22X1 U3493 ( .A(n4729), .B(n4580), .C(n4728), .D(n4582), .Y(n5713) );
  OAI21X1 U3494 ( .A(n4558), .B(n4716), .C(n5714), .Y(n3342) );
  OAI22X1 U3495 ( .A(b[7]), .B(n5715), .C(n4727), .D(n5715), .Y(n5714) );
  OAI22X1 U3496 ( .A(n4729), .B(n4582), .C(n4728), .D(n4584), .Y(n5715) );
  OAI21X1 U3497 ( .A(n4558), .B(n4715), .C(n5716), .Y(n3341) );
  OAI22X1 U3498 ( .A(b[8]), .B(n5717), .C(n4727), .D(n5717), .Y(n5716) );
  OAI22X1 U3499 ( .A(n4729), .B(n4584), .C(n4728), .D(n4587), .Y(n5717) );
  OAI21X1 U3500 ( .A(n4558), .B(n4713), .C(n5718), .Y(n3340) );
  OAI22X1 U3501 ( .A(n4586), .B(n5719), .C(n4727), .D(n5719), .Y(n5718) );
  OAI22X1 U3502 ( .A(n4729), .B(n4587), .C(n4728), .D(n4589), .Y(n5719) );
  OAI21X1 U3503 ( .A(n4558), .B(n4712), .C(n5720), .Y(n3339) );
  OAI22X1 U3504 ( .A(b[10]), .B(n5721), .C(n4727), .D(n5721), .Y(n5720) );
  OAI22X1 U3505 ( .A(n4729), .B(n4589), .C(n4728), .D(n4592), .Y(n5721) );
  OAI21X1 U3506 ( .A(n4558), .B(n4711), .C(n5722), .Y(n3338) );
  OAI22X1 U3507 ( .A(n4591), .B(n5723), .C(n4727), .D(n5723), .Y(n5722) );
  OAI22X1 U3508 ( .A(n4729), .B(n4592), .C(n4728), .D(n4594), .Y(n5723) );
  OAI21X1 U3509 ( .A(n4558), .B(n4708), .C(n5724), .Y(n3337) );
  OAI22X1 U3510 ( .A(n4596), .B(n5725), .C(n4727), .D(n5725), .Y(n5724) );
  OAI22X1 U3511 ( .A(n4728), .B(n4599), .C(n4729), .D(n4726), .Y(n5725) );
  OAI21X1 U3512 ( .A(n4558), .B(n4707), .C(n5726), .Y(n3336) );
  OAI22X1 U3513 ( .A(b[14]), .B(n5727), .C(n4727), .D(n5727), .Y(n5726) );
  OAI22X1 U3514 ( .A(n4729), .B(n4599), .C(n4601), .D(n4728), .Y(n5727) );
  OAI21X1 U3515 ( .A(n4558), .B(n4710), .C(n5728), .Y(n2429) );
  OAI22X1 U3516 ( .A(b[12]), .B(n5729), .C(n4727), .D(n5729), .Y(n5728) );
  NAND3X1 U3517 ( .A(n5731), .B(a[31]), .C(n5732), .Y(n5730) );
  OAI22X1 U3518 ( .A(n4729), .B(n4594), .C(n4728), .D(n4726), .Y(n5729) );
  NOR2X1 U3519 ( .A(n5731), .B(a[31]), .Y(n5698) );
  NOR2X1 U3520 ( .A(n4730), .B(n5732), .Y(n5699) );
  XNOR2X1 U3521 ( .A(a[30]), .B(a[31]), .Y(n5732) );
  XNOR2X1 U3522 ( .A(a[30]), .B(n4672), .Y(n5731) );
endmodule


module poly5_DW_mult_uns_3 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n2132, n2135, n2138, n2141, n2144, n2147, n2150, n2153, n2156, n2159,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774;
  assign n2132 = a[2];
  assign n2135 = a[5];
  assign n2138 = a[8];
  assign n2141 = a[11];
  assign n2144 = a[14];
  assign n2147 = a[17];
  assign n2150 = a[20];
  assign n2153 = a[23];
  assign n2156 = a[26];
  assign n2159 = a[29];

  FAX1 U336 ( .A(n2406), .B(n2417), .C(n2353), .YC(n2352), .YS(product[46]) );
  FAX1 U337 ( .A(n2431), .B(n2418), .C(n2354), .YC(n2353), .YS(product[45]) );
  FAX1 U338 ( .A(n2444), .B(n2432), .C(n2355), .YC(n2354), .YS(product[44]) );
  FAX1 U339 ( .A(n2445), .B(n2458), .C(n2356), .YC(n2355), .YS(product[43]) );
  FAX1 U340 ( .A(n2474), .B(n2459), .C(n2357), .YC(n2356), .YS(product[42]) );
  FAX1 U341 ( .A(n2489), .B(n2475), .C(n2358), .YC(n2357), .YS(product[41]) );
  FAX1 U342 ( .A(n2490), .B(n2504), .C(n2359), .YC(n2358), .YS(product[40]) );
  FAX1 U343 ( .A(n2522), .B(n2505), .C(n2360), .YC(n2359), .YS(product[39]) );
  FAX1 U344 ( .A(n2539), .B(n2523), .C(n2361), .YC(n2360), .YS(product[38]) );
  FAX1 U345 ( .A(n2540), .B(n2556), .C(n2362), .YC(n2361), .YS(product[37]) );
  FAX1 U346 ( .A(n2574), .B(n2557), .C(n2363), .YC(n2362), .YS(product[36]) );
  FAX1 U347 ( .A(n2592), .B(n2575), .C(n2364), .YC(n2363), .YS(product[35]) );
  FAX1 U348 ( .A(n2593), .B(n2610), .C(n2365), .YC(n2364), .YS(product[34]) );
  FAX1 U349 ( .A(n2628), .B(n2611), .C(n2366), .YC(n2365), .YS(product[33]) );
  FAX1 U350 ( .A(n3629), .B(n2629), .C(n2367), .YC(n2366), .YS(product[32]) );
  FAX1 U351 ( .A(n2647), .B(n3630), .C(n2368), .YC(n2367), .YS(product[31]) );
  FAX1 U352 ( .A(n2665), .B(n3631), .C(n2369), .YC(n2368), .YS(product[30]) );
  FAX1 U353 ( .A(n2683), .B(n3632), .C(n2370), .YC(n2369), .YS(product[29]) );
  FAX1 U354 ( .A(n2701), .B(n3633), .C(n2371), .YC(n2370), .YS(product[28]) );
  FAX1 U355 ( .A(n2719), .B(n3634), .C(n2372), .YC(n2371), .YS(product[27]) );
  FAX1 U356 ( .A(n2737), .B(n3635), .C(n2373), .YC(n2372), .YS(product[26]) );
  FAX1 U357 ( .A(n2753), .B(n3636), .C(n2374), .YC(n2373), .YS(product[25]) );
  FAX1 U358 ( .A(n2769), .B(n3637), .C(n2375), .YC(n2374), .YS(product[24]) );
  FAX1 U359 ( .A(n2785), .B(n3638), .C(n2376), .YC(n2375), .YS(product[23]) );
  FAX1 U360 ( .A(n2799), .B(n3639), .C(n2377), .YC(n2376), .YS(product[22]) );
  FAX1 U361 ( .A(n2813), .B(n3640), .C(n2378), .YC(n2377), .YS(product[21]) );
  FAX1 U362 ( .A(n2827), .B(n3641), .C(n2379), .YC(n2378), .YS(product[20]) );
  FAX1 U363 ( .A(n2839), .B(n3642), .C(n2380), .YC(n2379), .YS(product[19]) );
  FAX1 U364 ( .A(n2851), .B(n3643), .C(n2381), .YC(n2380), .YS(product[18]) );
  FAX1 U365 ( .A(n2863), .B(n3644), .C(n2382), .YC(n2381), .YS(product[17]) );
  FAX1 U366 ( .A(n2873), .B(n3645), .C(n2383), .YC(n2382), .YS(product[16]) );
  FAX1 U367 ( .A(n2883), .B(n3646), .C(n2384), .YC(n2383), .YS(product[15]) );
  FAX1 U368 ( .A(n2893), .B(n3647), .C(n2385), .YC(n2384), .YS(product[14]) );
  FAX1 U369 ( .A(n2901), .B(n3648), .C(n2386), .YC(n2385), .YS(product[13]) );
  FAX1 U370 ( .A(n2909), .B(n3649), .C(n2387), .YC(n2386), .YS(product[12]) );
  FAX1 U371 ( .A(n2917), .B(n3650), .C(n2388), .YC(n2387), .YS(product[11]) );
  FAX1 U372 ( .A(n2923), .B(n3651), .C(n2389), .YC(n2388), .YS(product[10]) );
  FAX1 U373 ( .A(n2929), .B(n3652), .C(n2390), .YC(n2389), .YS(product[9]) );
  FAX1 U374 ( .A(n2935), .B(n3653), .C(n2391), .YC(n2390), .YS(product[8]) );
  FAX1 U375 ( .A(n2939), .B(n3654), .C(n2392), .YC(n2391), .YS(product[7]) );
  FAX1 U376 ( .A(n2943), .B(n3655), .C(n2393), .YC(n2392), .YS(product[6]) );
  FAX1 U377 ( .A(n2947), .B(n3656), .C(n2394), .YC(n2393), .YS(product[5]) );
  FAX1 U378 ( .A(n3657), .B(n2949), .C(n2395), .YC(n2394), .YS(product[4]) );
  FAX1 U379 ( .A(n2951), .B(n3658), .C(n2396), .YC(n2395), .YS(product[3]) );
  HAX1 U380 ( .A(n3659), .B(n2397), .YC(n2396), .YS(product[2]) );
  HAX1 U381 ( .A(n2398), .B(n3660), .YC(n2397), .YS(product[1]) );
  HAX1 U382 ( .A(n2132), .B(n3661), .YC(n2398), .YS(product[0]) );
  FAX1 U384 ( .A(n2408), .B(n3455), .C(n2419), .YC(n2405), .YS(n2406) );
  FAX1 U385 ( .A(n2410), .B(n2421), .C(n3425), .YC(n2407), .YS(n2408) );
  FAX1 U386 ( .A(n2412), .B(n3398), .C(n2423), .YC(n2409), .YS(n2410) );
  FAX1 U387 ( .A(n2414), .B(n2425), .C(n3374), .YC(n2411), .YS(n2412) );
  FAX1 U388 ( .A(n2416), .B(n3353), .C(n2427), .YC(n2413), .YS(n2414) );
  FAX1 U389 ( .A(n4781), .B(n2429), .C(n3336), .YC(n2415), .YS(n2416) );
  FAX1 U390 ( .A(n3456), .B(n2420), .C(n3488), .YC(n2417), .YS(n2418) );
  FAX1 U391 ( .A(n2435), .B(n2422), .C(n2433), .YC(n2419), .YS(n2420) );
  FAX1 U392 ( .A(n3399), .B(n2424), .C(n3426), .YC(n2421), .YS(n2422) );
  FAX1 U393 ( .A(n2439), .B(n2426), .C(n2437), .YC(n2423), .YS(n2424) );
  FAX1 U394 ( .A(n2441), .B(n2428), .C(n3375), .YC(n2425), .YS(n2426) );
  FAX1 U395 ( .A(n4747), .B(n3337), .C(n3354), .YC(n2427), .YS(n2428) );
  FAX1 U397 ( .A(n2446), .B(n2434), .C(n3489), .YC(n2431), .YS(n2432) );
  FAX1 U398 ( .A(n2448), .B(n2436), .C(n3457), .YC(n2433), .YS(n2434) );
  FAX1 U399 ( .A(n2450), .B(n2438), .C(n3427), .YC(n2435), .YS(n2436) );
  FAX1 U400 ( .A(n2452), .B(n2440), .C(n3400), .YC(n2437), .YS(n2438) );
  FAX1 U401 ( .A(n2454), .B(n2442), .C(n3376), .YC(n2439), .YS(n2440) );
  FAX1 U402 ( .A(n2456), .B(n4747), .C(n3355), .YC(n2441), .YS(n2442) );
  FAX1 U404 ( .A(n2447), .B(n3490), .C(n2460), .YC(n2444), .YS(n2445) );
  FAX1 U405 ( .A(n2449), .B(n2462), .C(n3458), .YC(n2446), .YS(n2447) );
  FAX1 U406 ( .A(n2451), .B(n3428), .C(n2464), .YC(n2448), .YS(n2449) );
  FAX1 U407 ( .A(n2453), .B(n2466), .C(n3401), .YC(n2450), .YS(n2451) );
  FAX1 U408 ( .A(n2455), .B(n3377), .C(n2468), .YC(n2452), .YS(n2453) );
  FAX1 U409 ( .A(n2457), .B(n3356), .C(n2470), .YC(n2454), .YS(n2455) );
  FAX1 U410 ( .A(n4783), .B(n2472), .C(n3338), .YC(n2456), .YS(n2457) );
  FAX1 U411 ( .A(n3491), .B(n2461), .C(n3523), .YC(n2458), .YS(n2459) );
  FAX1 U412 ( .A(n2478), .B(n2463), .C(n2476), .YC(n2460), .YS(n2461) );
  FAX1 U413 ( .A(n3429), .B(n2465), .C(n3459), .YC(n2462), .YS(n2463) );
  FAX1 U414 ( .A(n2482), .B(n2467), .C(n2480), .YC(n2464), .YS(n2465) );
  FAX1 U415 ( .A(n2484), .B(n2469), .C(n3402), .YC(n2466), .YS(n2467) );
  FAX1 U416 ( .A(n2486), .B(n2471), .C(n3378), .YC(n2468), .YS(n2469) );
  FAX1 U417 ( .A(n4752), .B(n3339), .C(n3357), .YC(n2470), .YS(n2471) );
  FAX1 U419 ( .A(n2491), .B(n2477), .C(n3524), .YC(n2474), .YS(n2475) );
  FAX1 U420 ( .A(n2493), .B(n2479), .C(n3492), .YC(n2476), .YS(n2477) );
  FAX1 U421 ( .A(n2495), .B(n2481), .C(n3460), .YC(n2478), .YS(n2479) );
  FAX1 U422 ( .A(n2497), .B(n2483), .C(n3430), .YC(n2480), .YS(n2481) );
  FAX1 U423 ( .A(n2499), .B(n2485), .C(n3403), .YC(n2482), .YS(n2483) );
  FAX1 U424 ( .A(n2501), .B(n2487), .C(n3379), .YC(n2484), .YS(n2485) );
  FAX1 U425 ( .A(n3340), .B(n4752), .C(n3358), .YC(n2486), .YS(n2487) );
  FAX1 U427 ( .A(n2492), .B(n3525), .C(n2506), .YC(n2489), .YS(n2490) );
  FAX1 U428 ( .A(n2494), .B(n2508), .C(n3493), .YC(n2491), .YS(n2492) );
  FAX1 U429 ( .A(n2496), .B(n3461), .C(n2510), .YC(n2493), .YS(n2494) );
  FAX1 U430 ( .A(n2498), .B(n2512), .C(n3431), .YC(n2495), .YS(n2496) );
  FAX1 U431 ( .A(n2500), .B(n3404), .C(n2514), .YC(n2497), .YS(n2498) );
  FAX1 U432 ( .A(n2502), .B(n3380), .C(n2516), .YC(n2499), .YS(n2500) );
  FAX1 U433 ( .A(n2503), .B(n2518), .C(n3359), .YC(n2501), .YS(n2502) );
  FAX1 U434 ( .A(n4785), .B(n2520), .C(n3341), .YC(n2472), .YS(n2503) );
  FAX1 U435 ( .A(n3526), .B(n2507), .C(n3558), .YC(n2504), .YS(n2505) );
  FAX1 U436 ( .A(n2526), .B(n2509), .C(n2524), .YC(n2506), .YS(n2507) );
  FAX1 U437 ( .A(n3462), .B(n2511), .C(n3494), .YC(n2508), .YS(n2509) );
  FAX1 U438 ( .A(n2530), .B(n2513), .C(n2528), .YC(n2510), .YS(n2511) );
  FAX1 U439 ( .A(n2532), .B(n2515), .C(n3432), .YC(n2512), .YS(n2513) );
  FAX1 U440 ( .A(n2534), .B(n2517), .C(n3405), .YC(n2514), .YS(n2515) );
  FAX1 U441 ( .A(n3360), .B(n2519), .C(n3381), .YC(n2516), .YS(n2517) );
  FAX1 U442 ( .A(n4756), .B(n3342), .C(n2536), .YC(n2518), .YS(n2519) );
  FAX1 U444 ( .A(n2541), .B(n2525), .C(n3559), .YC(n2522), .YS(n2523) );
  FAX1 U445 ( .A(n2543), .B(n2527), .C(n3527), .YC(n2524), .YS(n2525) );
  FAX1 U446 ( .A(n2545), .B(n2529), .C(n3495), .YC(n2526), .YS(n2527) );
  FAX1 U447 ( .A(n2547), .B(n2531), .C(n3463), .YC(n2528), .YS(n2529) );
  FAX1 U448 ( .A(n2549), .B(n2533), .C(n3433), .YC(n2530), .YS(n2531) );
  FAX1 U449 ( .A(n2551), .B(n2535), .C(n3406), .YC(n2532), .YS(n2533) );
  FAX1 U450 ( .A(n2553), .B(n2537), .C(n3382), .YC(n2534), .YS(n2535) );
  FAX1 U451 ( .A(n3343), .B(n4756), .C(n3361), .YC(n2536), .YS(n2537) );
  FAX1 U453 ( .A(n2542), .B(n3560), .C(n2558), .YC(n2539), .YS(n2540) );
  FAX1 U454 ( .A(n2544), .B(n2560), .C(n3528), .YC(n2541), .YS(n2542) );
  FAX1 U455 ( .A(n2546), .B(n3496), .C(n2562), .YC(n2543), .YS(n2544) );
  FAX1 U456 ( .A(n2548), .B(n2564), .C(n3464), .YC(n2545), .YS(n2546) );
  FAX1 U457 ( .A(n2550), .B(n3434), .C(n2566), .YC(n2547), .YS(n2548) );
  FAX1 U458 ( .A(n2552), .B(n3407), .C(n2568), .YC(n2549), .YS(n2550) );
  FAX1 U459 ( .A(n2554), .B(n2570), .C(n3383), .YC(n2551), .YS(n2552) );
  FAX1 U460 ( .A(n2555), .B(n2572), .C(n3362), .YC(n2553), .YS(n2554) );
  FAX1 U461 ( .A(n4595), .B(n4787), .C(n3344), .YC(n2520), .YS(n2555) );
  FAX1 U462 ( .A(n3561), .B(n2559), .C(n3593), .YC(n2556), .YS(n2557) );
  FAX1 U463 ( .A(n2578), .B(n2561), .C(n2576), .YC(n2558), .YS(n2559) );
  FAX1 U464 ( .A(n3497), .B(n2563), .C(n3529), .YC(n2560), .YS(n2561) );
  FAX1 U465 ( .A(n2582), .B(n2565), .C(n2580), .YC(n2562), .YS(n2563) );
  FAX1 U466 ( .A(n2584), .B(n2567), .C(n3465), .YC(n2564), .YS(n2565) );
  FAX1 U467 ( .A(n2586), .B(n2569), .C(n3435), .YC(n2566), .YS(n2567) );
  FAX1 U468 ( .A(n3384), .B(n2571), .C(n3408), .YC(n2568), .YS(n2569) );
  FAX1 U469 ( .A(n3363), .B(n2573), .C(n2588), .YC(n2570), .YS(n2571) );
  FAX1 U470 ( .A(n2132), .B(n3345), .C(n2590), .YC(n2572), .YS(n2573) );
  FAX1 U471 ( .A(n2594), .B(n2577), .C(n3594), .YC(n2574), .YS(n2575) );
  FAX1 U472 ( .A(n3530), .B(n2579), .C(n3562), .YC(n2576), .YS(n2577) );
  FAX1 U473 ( .A(n2598), .B(n2581), .C(n2596), .YC(n2578), .YS(n2579) );
  FAX1 U474 ( .A(n3466), .B(n2583), .C(n3498), .YC(n2580), .YS(n2581) );
  FAX1 U475 ( .A(n3436), .B(n2585), .C(n2600), .YC(n2582), .YS(n2583) );
  FAX1 U476 ( .A(n2604), .B(n2587), .C(n2602), .YC(n2584), .YS(n2585) );
  FAX1 U477 ( .A(n3385), .B(n2589), .C(n3409), .YC(n2586), .YS(n2587) );
  FAX1 U478 ( .A(n3364), .B(n2591), .C(n2606), .YC(n2588), .YS(n2589) );
  FAX1 U479 ( .A(n2132), .B(n3346), .C(n2608), .YC(n2590), .YS(n2591) );
  FAX1 U480 ( .A(n2595), .B(n2612), .C(n3595), .YC(n2592), .YS(n2593) );
  FAX1 U481 ( .A(n2597), .B(n2614), .C(n3563), .YC(n2594), .YS(n2595) );
  FAX1 U482 ( .A(n2599), .B(n2616), .C(n3531), .YC(n2596), .YS(n2597) );
  FAX1 U483 ( .A(n2601), .B(n2618), .C(n3499), .YC(n2598), .YS(n2599) );
  FAX1 U484 ( .A(n2603), .B(n2620), .C(n3467), .YC(n2600), .YS(n2601) );
  FAX1 U485 ( .A(n2605), .B(n2622), .C(n3437), .YC(n2602), .YS(n2603) );
  FAX1 U486 ( .A(n2607), .B(n2624), .C(n3410), .YC(n2604), .YS(n2605) );
  FAX1 U487 ( .A(n2609), .B(n2626), .C(n3386), .YC(n2606), .YS(n2607) );
  FAX1 U488 ( .A(n2132), .B(n3347), .C(n3365), .YC(n2608), .YS(n2609) );
  FAX1 U489 ( .A(n2613), .B(n3596), .C(n3628), .YC(n2610), .YS(n2611) );
  FAX1 U490 ( .A(n2615), .B(n3564), .C(n2630), .YC(n2612), .YS(n2613) );
  FAX1 U491 ( .A(n2617), .B(n3532), .C(n2632), .YC(n2614), .YS(n2615) );
  FAX1 U492 ( .A(n2619), .B(n3500), .C(n2634), .YC(n2616), .YS(n2617) );
  FAX1 U493 ( .A(n2621), .B(n3468), .C(n2636), .YC(n2618), .YS(n2619) );
  FAX1 U494 ( .A(n2623), .B(n3438), .C(n2638), .YC(n2620), .YS(n2621) );
  FAX1 U495 ( .A(n2625), .B(n3411), .C(n2640), .YC(n2622), .YS(n2623) );
  FAX1 U496 ( .A(n2627), .B(n3387), .C(n2642), .YC(n2624), .YS(n2625) );
  FAX1 U497 ( .A(n3348), .B(n3366), .C(n2644), .YC(n2626), .YS(n2627) );
  FAX1 U498 ( .A(n2631), .B(n3597), .C(n2646), .YC(n2628), .YS(n2629) );
  FAX1 U499 ( .A(n2633), .B(n3565), .C(n2648), .YC(n2630), .YS(n2631) );
  FAX1 U500 ( .A(n2635), .B(n3533), .C(n2650), .YC(n2632), .YS(n2633) );
  FAX1 U501 ( .A(n2637), .B(n3501), .C(n2652), .YC(n2634), .YS(n2635) );
  FAX1 U502 ( .A(n2639), .B(n3469), .C(n2654), .YC(n2636), .YS(n2637) );
  FAX1 U503 ( .A(n2641), .B(n3439), .C(n2656), .YC(n2638), .YS(n2639) );
  FAX1 U504 ( .A(n2643), .B(n3412), .C(n2658), .YC(n2640), .YS(n2641) );
  FAX1 U505 ( .A(n2645), .B(n3388), .C(n2660), .YC(n2642), .YS(n2643) );
  FAX1 U506 ( .A(n3349), .B(n3367), .C(n2662), .YC(n2644), .YS(n2645) );
  FAX1 U507 ( .A(n2649), .B(n3598), .C(n2664), .YC(n2646), .YS(n2647) );
  FAX1 U508 ( .A(n2651), .B(n3566), .C(n2666), .YC(n2648), .YS(n2649) );
  FAX1 U509 ( .A(n2653), .B(n3534), .C(n2668), .YC(n2650), .YS(n2651) );
  FAX1 U510 ( .A(n2655), .B(n3502), .C(n2670), .YC(n2652), .YS(n2653) );
  FAX1 U511 ( .A(n2657), .B(n3470), .C(n2672), .YC(n2654), .YS(n2655) );
  FAX1 U512 ( .A(n2659), .B(n3440), .C(n2674), .YC(n2656), .YS(n2657) );
  FAX1 U513 ( .A(n2661), .B(n3413), .C(n2676), .YC(n2658), .YS(n2659) );
  FAX1 U514 ( .A(n2663), .B(n3389), .C(n2678), .YC(n2660), .YS(n2661) );
  FAX1 U515 ( .A(n3350), .B(n3368), .C(n2680), .YC(n2662), .YS(n2663) );
  FAX1 U516 ( .A(n2667), .B(n3599), .C(n2682), .YC(n2664), .YS(n2665) );
  FAX1 U517 ( .A(n2669), .B(n3567), .C(n2684), .YC(n2666), .YS(n2667) );
  FAX1 U518 ( .A(n2671), .B(n3535), .C(n2686), .YC(n2668), .YS(n2669) );
  FAX1 U519 ( .A(n2673), .B(n3503), .C(n2688), .YC(n2670), .YS(n2671) );
  FAX1 U520 ( .A(n2675), .B(n3471), .C(n2690), .YC(n2672), .YS(n2673) );
  FAX1 U521 ( .A(n2677), .B(n3441), .C(n2692), .YC(n2674), .YS(n2675) );
  FAX1 U522 ( .A(n2679), .B(n3414), .C(n2694), .YC(n2676), .YS(n2677) );
  FAX1 U523 ( .A(n2681), .B(n3390), .C(n2696), .YC(n2678), .YS(n2679) );
  FAX1 U524 ( .A(n3351), .B(n3369), .C(n2698), .YC(n2680), .YS(n2681) );
  FAX1 U525 ( .A(n2685), .B(n3600), .C(n2700), .YC(n2682), .YS(n2683) );
  FAX1 U526 ( .A(n2687), .B(n3568), .C(n2702), .YC(n2684), .YS(n2685) );
  FAX1 U527 ( .A(n2689), .B(n3536), .C(n2704), .YC(n2686), .YS(n2687) );
  FAX1 U528 ( .A(n2691), .B(n3504), .C(n2706), .YC(n2688), .YS(n2689) );
  FAX1 U529 ( .A(n2693), .B(n3472), .C(n2708), .YC(n2690), .YS(n2691) );
  FAX1 U530 ( .A(n2695), .B(n3442), .C(n2710), .YC(n2692), .YS(n2693) );
  FAX1 U531 ( .A(n2697), .B(n3415), .C(n2712), .YC(n2694), .YS(n2695) );
  FAX1 U532 ( .A(n2699), .B(n3391), .C(n2714), .YC(n2696), .YS(n2697) );
  HAX1 U533 ( .A(n3370), .B(n2716), .YC(n2698), .YS(n2699) );
  FAX1 U534 ( .A(n2703), .B(n3601), .C(n2718), .YC(n2700), .YS(n2701) );
  FAX1 U535 ( .A(n2705), .B(n3569), .C(n2720), .YC(n2702), .YS(n2703) );
  FAX1 U536 ( .A(n2707), .B(n3537), .C(n2722), .YC(n2704), .YS(n2705) );
  FAX1 U537 ( .A(n2709), .B(n3505), .C(n2724), .YC(n2706), .YS(n2707) );
  FAX1 U538 ( .A(n2711), .B(n3473), .C(n2726), .YC(n2708), .YS(n2709) );
  FAX1 U539 ( .A(n2713), .B(n3443), .C(n2728), .YC(n2710), .YS(n2711) );
  FAX1 U540 ( .A(n2715), .B(n3416), .C(n2730), .YC(n2712), .YS(n2713) );
  FAX1 U541 ( .A(n3392), .B(n2717), .C(n2732), .YC(n2714), .YS(n2715) );
  HAX1 U542 ( .A(n2734), .B(n3371), .YC(n2716), .YS(n2717) );
  FAX1 U543 ( .A(n2721), .B(n3602), .C(n2736), .YC(n2718), .YS(n2719) );
  FAX1 U544 ( .A(n2723), .B(n3570), .C(n2738), .YC(n2720), .YS(n2721) );
  FAX1 U545 ( .A(n2725), .B(n3538), .C(n2740), .YC(n2722), .YS(n2723) );
  FAX1 U546 ( .A(n2727), .B(n3506), .C(n2742), .YC(n2724), .YS(n2725) );
  FAX1 U547 ( .A(n2729), .B(n3474), .C(n2744), .YC(n2726), .YS(n2727) );
  FAX1 U548 ( .A(n2731), .B(n3444), .C(n2746), .YC(n2728), .YS(n2729) );
  FAX1 U549 ( .A(n2733), .B(n3417), .C(n2748), .YC(n2730), .YS(n2731) );
  FAX1 U550 ( .A(n2735), .B(n3393), .C(n2750), .YC(n2732), .YS(n2733) );
  HAX1 U551 ( .A(n2159), .B(n3372), .YC(n2734), .YS(n2735) );
  FAX1 U552 ( .A(n2739), .B(n3603), .C(n2752), .YC(n2736), .YS(n2737) );
  FAX1 U553 ( .A(n2741), .B(n3571), .C(n2754), .YC(n2738), .YS(n2739) );
  FAX1 U554 ( .A(n2743), .B(n3539), .C(n2756), .YC(n2740), .YS(n2741) );
  FAX1 U555 ( .A(n2745), .B(n3507), .C(n2758), .YC(n2742), .YS(n2743) );
  FAX1 U556 ( .A(n2747), .B(n3475), .C(n2760), .YC(n2744), .YS(n2745) );
  FAX1 U557 ( .A(n2749), .B(n3445), .C(n2762), .YC(n2746), .YS(n2747) );
  FAX1 U558 ( .A(n2751), .B(n3418), .C(n2764), .YC(n2748), .YS(n2749) );
  HAX1 U559 ( .A(n3394), .B(n2766), .YC(n2750), .YS(n2751) );
  FAX1 U560 ( .A(n2755), .B(n3604), .C(n2768), .YC(n2752), .YS(n2753) );
  FAX1 U561 ( .A(n2757), .B(n3572), .C(n2770), .YC(n2754), .YS(n2755) );
  FAX1 U562 ( .A(n2759), .B(n3540), .C(n2772), .YC(n2756), .YS(n2757) );
  FAX1 U563 ( .A(n2761), .B(n3508), .C(n2774), .YC(n2758), .YS(n2759) );
  FAX1 U564 ( .A(n2763), .B(n3476), .C(n2776), .YC(n2760), .YS(n2761) );
  FAX1 U565 ( .A(n2765), .B(n3446), .C(n2778), .YC(n2762), .YS(n2763) );
  FAX1 U566 ( .A(n3419), .B(n2767), .C(n2780), .YC(n2764), .YS(n2765) );
  HAX1 U567 ( .A(n2782), .B(n3395), .YC(n2766), .YS(n2767) );
  FAX1 U568 ( .A(n2771), .B(n3605), .C(n2784), .YC(n2768), .YS(n2769) );
  FAX1 U569 ( .A(n2773), .B(n3573), .C(n2786), .YC(n2770), .YS(n2771) );
  FAX1 U570 ( .A(n2775), .B(n3541), .C(n2788), .YC(n2772), .YS(n2773) );
  FAX1 U571 ( .A(n2777), .B(n3509), .C(n2790), .YC(n2774), .YS(n2775) );
  FAX1 U572 ( .A(n2779), .B(n3477), .C(n2792), .YC(n2776), .YS(n2777) );
  FAX1 U573 ( .A(n2781), .B(n3447), .C(n2794), .YC(n2778), .YS(n2779) );
  FAX1 U574 ( .A(n2783), .B(n3420), .C(n2796), .YC(n2780), .YS(n2781) );
  HAX1 U575 ( .A(n2156), .B(n3396), .YC(n2782), .YS(n2783) );
  FAX1 U576 ( .A(n2787), .B(n3606), .C(n2798), .YC(n2784), .YS(n2785) );
  FAX1 U577 ( .A(n2789), .B(n3574), .C(n2800), .YC(n2786), .YS(n2787) );
  FAX1 U578 ( .A(n2791), .B(n3542), .C(n2802), .YC(n2788), .YS(n2789) );
  FAX1 U579 ( .A(n2793), .B(n3510), .C(n2804), .YC(n2790), .YS(n2791) );
  FAX1 U580 ( .A(n2795), .B(n3478), .C(n2806), .YC(n2792), .YS(n2793) );
  FAX1 U581 ( .A(n2797), .B(n3448), .C(n2808), .YC(n2794), .YS(n2795) );
  HAX1 U582 ( .A(n3421), .B(n2810), .YC(n2796), .YS(n2797) );
  FAX1 U583 ( .A(n2801), .B(n3607), .C(n2812), .YC(n2798), .YS(n2799) );
  FAX1 U584 ( .A(n2803), .B(n3575), .C(n2814), .YC(n2800), .YS(n2801) );
  FAX1 U585 ( .A(n2805), .B(n3543), .C(n2816), .YC(n2802), .YS(n2803) );
  FAX1 U586 ( .A(n2807), .B(n3511), .C(n2818), .YC(n2804), .YS(n2805) );
  FAX1 U587 ( .A(n2809), .B(n3479), .C(n2820), .YC(n2806), .YS(n2807) );
  FAX1 U588 ( .A(n3449), .B(n2811), .C(n2822), .YC(n2808), .YS(n2809) );
  HAX1 U589 ( .A(n2824), .B(n3422), .YC(n2810), .YS(n2811) );
  FAX1 U590 ( .A(n2815), .B(n3608), .C(n2826), .YC(n2812), .YS(n2813) );
  FAX1 U591 ( .A(n2817), .B(n3576), .C(n2828), .YC(n2814), .YS(n2815) );
  FAX1 U592 ( .A(n2819), .B(n3544), .C(n2830), .YC(n2816), .YS(n2817) );
  FAX1 U593 ( .A(n2821), .B(n3512), .C(n2832), .YC(n2818), .YS(n2819) );
  FAX1 U594 ( .A(n2823), .B(n3480), .C(n2834), .YC(n2820), .YS(n2821) );
  FAX1 U595 ( .A(n2825), .B(n3450), .C(n2836), .YC(n2822), .YS(n2823) );
  HAX1 U596 ( .A(n2153), .B(n3423), .YC(n2824), .YS(n2825) );
  FAX1 U597 ( .A(n2829), .B(n3609), .C(n2838), .YC(n2826), .YS(n2827) );
  FAX1 U598 ( .A(n2831), .B(n3577), .C(n2840), .YC(n2828), .YS(n2829) );
  FAX1 U599 ( .A(n2833), .B(n3545), .C(n2842), .YC(n2830), .YS(n2831) );
  FAX1 U600 ( .A(n2835), .B(n3513), .C(n2844), .YC(n2832), .YS(n2833) );
  FAX1 U601 ( .A(n2837), .B(n3481), .C(n2846), .YC(n2834), .YS(n2835) );
  HAX1 U602 ( .A(n3451), .B(n2848), .YC(n2836), .YS(n2837) );
  FAX1 U603 ( .A(n2841), .B(n3610), .C(n2850), .YC(n2838), .YS(n2839) );
  FAX1 U604 ( .A(n2843), .B(n3578), .C(n2852), .YC(n2840), .YS(n2841) );
  FAX1 U605 ( .A(n2845), .B(n3546), .C(n2854), .YC(n2842), .YS(n2843) );
  FAX1 U606 ( .A(n2847), .B(n3514), .C(n2856), .YC(n2844), .YS(n2845) );
  FAX1 U607 ( .A(n3482), .B(n2849), .C(n2858), .YC(n2846), .YS(n2847) );
  HAX1 U608 ( .A(n2860), .B(n3452), .YC(n2848), .YS(n2849) );
  FAX1 U609 ( .A(n2853), .B(n3611), .C(n2862), .YC(n2850), .YS(n2851) );
  FAX1 U610 ( .A(n2855), .B(n3579), .C(n2864), .YC(n2852), .YS(n2853) );
  FAX1 U611 ( .A(n2857), .B(n3547), .C(n2866), .YC(n2854), .YS(n2855) );
  FAX1 U612 ( .A(n2859), .B(n3515), .C(n2868), .YC(n2856), .YS(n2857) );
  FAX1 U613 ( .A(n2861), .B(n3483), .C(n2870), .YC(n2858), .YS(n2859) );
  HAX1 U614 ( .A(n4719), .B(n3453), .YC(n2860), .YS(n2861) );
  FAX1 U615 ( .A(n2865), .B(n3612), .C(n2872), .YC(n2862), .YS(n2863) );
  FAX1 U616 ( .A(n2867), .B(n3580), .C(n2874), .YC(n2864), .YS(n2865) );
  FAX1 U617 ( .A(n2869), .B(n3548), .C(n2876), .YC(n2866), .YS(n2867) );
  FAX1 U618 ( .A(n2871), .B(n3516), .C(n2878), .YC(n2868), .YS(n2869) );
  HAX1 U619 ( .A(n3484), .B(n2880), .YC(n2870), .YS(n2871) );
  FAX1 U620 ( .A(n2875), .B(n3613), .C(n2882), .YC(n2872), .YS(n2873) );
  FAX1 U621 ( .A(n2877), .B(n3581), .C(n2884), .YC(n2874), .YS(n2875) );
  FAX1 U622 ( .A(n2879), .B(n3549), .C(n2886), .YC(n2876), .YS(n2877) );
  FAX1 U623 ( .A(n3517), .B(n2881), .C(n2888), .YC(n2878), .YS(n2879) );
  HAX1 U624 ( .A(n2890), .B(n3485), .YC(n2880), .YS(n2881) );
  FAX1 U625 ( .A(n2885), .B(n3614), .C(n2892), .YC(n2882), .YS(n2883) );
  FAX1 U626 ( .A(n2887), .B(n3582), .C(n2894), .YC(n2884), .YS(n2885) );
  FAX1 U627 ( .A(n2889), .B(n3550), .C(n2896), .YC(n2886), .YS(n2887) );
  FAX1 U628 ( .A(n2891), .B(n3518), .C(n2898), .YC(n2888), .YS(n2889) );
  HAX1 U629 ( .A(n2147), .B(n3486), .YC(n2890), .YS(n2891) );
  FAX1 U630 ( .A(n2895), .B(n3615), .C(n2900), .YC(n2892), .YS(n2893) );
  FAX1 U631 ( .A(n2897), .B(n3583), .C(n2902), .YC(n2894), .YS(n2895) );
  FAX1 U632 ( .A(n2899), .B(n3551), .C(n2904), .YC(n2896), .YS(n2897) );
  HAX1 U633 ( .A(n3519), .B(n2906), .YC(n2898), .YS(n2899) );
  FAX1 U634 ( .A(n2903), .B(n3616), .C(n2908), .YC(n2900), .YS(n2901) );
  FAX1 U635 ( .A(n2905), .B(n3584), .C(n2910), .YC(n2902), .YS(n2903) );
  FAX1 U636 ( .A(n3552), .B(n2907), .C(n2912), .YC(n2904), .YS(n2905) );
  HAX1 U637 ( .A(n2914), .B(n3520), .YC(n2906), .YS(n2907) );
  FAX1 U638 ( .A(n2911), .B(n3617), .C(n2916), .YC(n2908), .YS(n2909) );
  FAX1 U639 ( .A(n2913), .B(n3585), .C(n2918), .YC(n2910), .YS(n2911) );
  FAX1 U640 ( .A(n2915), .B(n3553), .C(n2920), .YC(n2912), .YS(n2913) );
  HAX1 U641 ( .A(n2144), .B(n3521), .YC(n2914), .YS(n2915) );
  FAX1 U642 ( .A(n2919), .B(n3618), .C(n2922), .YC(n2916), .YS(n2917) );
  FAX1 U643 ( .A(n2921), .B(n3586), .C(n2924), .YC(n2918), .YS(n2919) );
  HAX1 U644 ( .A(n3554), .B(n2926), .YC(n2920), .YS(n2921) );
  FAX1 U645 ( .A(n2925), .B(n3619), .C(n2928), .YC(n2922), .YS(n2923) );
  FAX1 U646 ( .A(n3587), .B(n2927), .C(n2930), .YC(n2924), .YS(n2925) );
  HAX1 U647 ( .A(n2932), .B(n3555), .YC(n2926), .YS(n2927) );
  FAX1 U648 ( .A(n2931), .B(n3620), .C(n2934), .YC(n2928), .YS(n2929) );
  FAX1 U649 ( .A(n2933), .B(n3588), .C(n2936), .YC(n2930), .YS(n2931) );
  HAX1 U650 ( .A(n2141), .B(n3556), .YC(n2932), .YS(n2933) );
  FAX1 U651 ( .A(n2937), .B(n3621), .C(n2938), .YC(n2934), .YS(n2935) );
  HAX1 U652 ( .A(n3589), .B(n2940), .YC(n2936), .YS(n2937) );
  FAX1 U653 ( .A(n3622), .B(n2941), .C(n2942), .YC(n2938), .YS(n2939) );
  HAX1 U654 ( .A(n2944), .B(n3590), .YC(n2940), .YS(n2941) );
  FAX1 U655 ( .A(n2945), .B(n3623), .C(n2946), .YC(n2942), .YS(n2943) );
  HAX1 U656 ( .A(n2138), .B(n3591), .YC(n2944), .YS(n2945) );
  HAX1 U657 ( .A(n3624), .B(n2948), .YC(n2946), .YS(n2947) );
  HAX1 U658 ( .A(n2950), .B(n3625), .YC(n2948), .YS(n2949) );
  HAX1 U659 ( .A(n2135), .B(n3626), .YC(n2950), .YS(n2951) );
  HAX1 U1990 ( .A(b[31]), .B(n3270), .YC(n3301), .YS(n3302) );
  FAX1 U1991 ( .A(b[31]), .B(b[30]), .C(n3271), .YC(n3270), .YS(n3303) );
  FAX1 U1992 ( .A(b[30]), .B(b[29]), .C(n3272), .YC(n3271), .YS(n3304) );
  FAX1 U1993 ( .A(b[29]), .B(b[28]), .C(n3273), .YC(n3272), .YS(n3305) );
  FAX1 U1994 ( .A(b[28]), .B(b[27]), .C(n3274), .YC(n3273), .YS(n3306) );
  FAX1 U1995 ( .A(b[27]), .B(b[26]), .C(n3275), .YC(n3274), .YS(n3307) );
  FAX1 U1996 ( .A(b[26]), .B(b[25]), .C(n3276), .YC(n3275), .YS(n3308) );
  FAX1 U1997 ( .A(b[25]), .B(n4569), .C(n3277), .YC(n3276), .YS(n3309) );
  FAX1 U1998 ( .A(n4569), .B(n4710), .C(n3278), .YC(n3277), .YS(n3310) );
  FAX1 U1999 ( .A(n4711), .B(n4707), .C(n3279), .YC(n3278), .YS(n3311) );
  FAX1 U2000 ( .A(n4706), .B(n4703), .C(n3280), .YC(n3279), .YS(n3312) );
  FAX1 U2001 ( .A(n4703), .B(n4699), .C(n3281), .YC(n3280), .YS(n3313) );
  FAX1 U2002 ( .A(n4699), .B(n4695), .C(n3282), .YC(n3281), .YS(n3314) );
  FAX1 U2003 ( .A(n4695), .B(n4690), .C(n3283), .YC(n3282), .YS(n3315) );
  FAX1 U2004 ( .A(n4689), .B(n4685), .C(n3284), .YC(n3283), .YS(n3316) );
  FAX1 U2005 ( .A(n4684), .B(n4680), .C(n3285), .YC(n3284), .YS(n3317) );
  FAX1 U2006 ( .A(n4679), .B(n4675), .C(n3286), .YC(n3285), .YS(n3318) );
  FAX1 U2007 ( .A(n4674), .B(n4670), .C(n3287), .YC(n3286), .YS(n3319) );
  FAX1 U2008 ( .A(n4669), .B(n4665), .C(n3288), .YC(n3287), .YS(n3320) );
  FAX1 U2009 ( .A(n4667), .B(n4661), .C(n3289), .YC(n3288), .YS(n3321) );
  FAX1 U2010 ( .A(n4660), .B(n4656), .C(n3290), .YC(n3289), .YS(n3322) );
  FAX1 U2011 ( .A(n4655), .B(n4651), .C(n3291), .YC(n3290), .YS(n3323) );
  FAX1 U2012 ( .A(n4650), .B(n4646), .C(n3292), .YC(n3291), .YS(n3324) );
  FAX1 U2013 ( .A(n4648), .B(n4642), .C(n3293), .YC(n3292), .YS(n3325) );
  FAX1 U2014 ( .A(n4641), .B(n4637), .C(n3294), .YC(n3293), .YS(n3326) );
  FAX1 U2015 ( .A(n4636), .B(n4632), .C(n3295), .YC(n3294), .YS(n3327) );
  FAX1 U2016 ( .A(n4631), .B(n4627), .C(n3296), .YC(n3295), .YS(n3328) );
  FAX1 U2017 ( .A(n4629), .B(n4623), .C(n3297), .YC(n3296), .YS(n3329) );
  FAX1 U2018 ( .A(n4622), .B(n4618), .C(n3298), .YC(n3297), .YS(n3330) );
  FAX1 U2019 ( .A(n4617), .B(n4613), .C(n3299), .YC(n3298), .YS(n3331) );
  FAX1 U2020 ( .A(n4612), .B(n4610), .C(n3300), .YC(n3299), .YS(n3332) );
  HAX1 U2021 ( .A(n4610), .B(n4605), .YC(n3300), .YS(n3333) );
  OR2X2 U2024 ( .A(n5431), .B(n5432), .Y(n4552) );
  OR2X2 U2025 ( .A(n4918), .B(n4790), .Y(n4553) );
  OR2X2 U2026 ( .A(n4780), .B(n5430), .Y(n4554) );
  NAND2X1 U2027 ( .A(n5603), .B(n5601), .Y(n4555) );
  NAND2X1 U2028 ( .A(n4776), .B(n5674), .Y(n4556) );
  NAND2X1 U2029 ( .A(n4773), .B(n5737), .Y(n4557) );
  NAND2X1 U2030 ( .A(a[31]), .B(n4769), .Y(n4558) );
  INVX1 U2031 ( .A(b[29]), .Y(n4727) );
  INVX2 U2032 ( .A(n3329), .Y(n4759) );
  INVX2 U2033 ( .A(n3328), .Y(n4758) );
  INVX2 U2034 ( .A(n3327), .Y(n4757) );
  INVX2 U2035 ( .A(n3325), .Y(n4754) );
  INVX2 U2036 ( .A(n3324), .Y(n4753) );
  INVX2 U2037 ( .A(n3320), .Y(n4748) );
  INVX2 U2038 ( .A(n3326), .Y(n4755) );
  INVX2 U2039 ( .A(n3321), .Y(n4749) );
  INVX2 U2040 ( .A(n3323), .Y(n4751) );
  INVX2 U2041 ( .A(n3318), .Y(n4745) );
  INVX2 U2042 ( .A(n3322), .Y(n4750) );
  INVX2 U2043 ( .A(n3319), .Y(n4746) );
  INVX2 U2044 ( .A(n3317), .Y(n4744) );
  INVX2 U2045 ( .A(n3316), .Y(n4743) );
  INVX2 U2046 ( .A(n3315), .Y(n4742) );
  INVX2 U2047 ( .A(n3314), .Y(n4741) );
  INVX2 U2048 ( .A(n3313), .Y(n4740) );
  INVX2 U2049 ( .A(n3312), .Y(n4739) );
  INVX2 U2050 ( .A(n3311), .Y(n4738) );
  INVX2 U2051 ( .A(n3333), .Y(n4765) );
  INVX2 U2052 ( .A(n4611), .Y(n4610) );
  INVX2 U2053 ( .A(n3332), .Y(n4762) );
  INVX2 U2054 ( .A(n3331), .Y(n4761) );
  INVX2 U2055 ( .A(n3330), .Y(n4760) );
  INVX2 U2056 ( .A(n4605), .Y(n4609) );
  INVX2 U2057 ( .A(n4627), .Y(n4630) );
  INVX2 U2058 ( .A(n4632), .Y(n4635) );
  INVX2 U2059 ( .A(n4637), .Y(n4640) );
  INVX2 U2060 ( .A(n4642), .Y(n4645) );
  INVX2 U2061 ( .A(n4646), .Y(n4649) );
  INVX2 U2062 ( .A(n4622), .Y(n4626) );
  INVX2 U2063 ( .A(n4670), .Y(n4673) );
  INVX2 U2064 ( .A(n4656), .Y(n4659) );
  INVX2 U2065 ( .A(n4651), .Y(n4654) );
  INVX2 U2066 ( .A(n4661), .Y(n4664) );
  INVX2 U2067 ( .A(n4665), .Y(n4668) );
  INVX2 U2068 ( .A(n4680), .Y(n4683) );
  INVX2 U2069 ( .A(n4690), .Y(n4693) );
  INVX2 U2070 ( .A(n4675), .Y(n4678) );
  INVX2 U2071 ( .A(n4694), .Y(n4697) );
  INVX2 U2072 ( .A(n4685), .Y(n4688) );
  INVX2 U2073 ( .A(n4707), .Y(n4709) );
  INVX2 U2074 ( .A(n4702), .Y(n4705) );
  INVX2 U2075 ( .A(n4710), .Y(n4712) );
  INVX2 U2076 ( .A(n4698), .Y(n4701) );
  INVX1 U2077 ( .A(b[1]), .Y(n4611) );
  BUFX2 U2078 ( .A(b[4]), .Y(n4622) );
  BUFX2 U2079 ( .A(b[4]), .Y(n4623) );
  INVX2 U2080 ( .A(n4613), .Y(n4616) );
  INVX2 U2081 ( .A(n4618), .Y(n4621) );
  BUFX2 U2082 ( .A(b[5]), .Y(n4628) );
  BUFX2 U2083 ( .A(b[4]), .Y(n4624) );
  BUFX2 U2084 ( .A(b[6]), .Y(n4631) );
  BUFX2 U2085 ( .A(b[7]), .Y(n4636) );
  BUFX2 U2086 ( .A(b[8]), .Y(n4641) );
  BUFX2 U2087 ( .A(b[10]), .Y(n4650) );
  BUFX2 U2088 ( .A(b[5]), .Y(n4627) );
  BUFX2 U2089 ( .A(b[9]), .Y(n4646) );
  BUFX2 U2090 ( .A(b[6]), .Y(n4632) );
  BUFX2 U2091 ( .A(b[7]), .Y(n4637) );
  BUFX2 U2092 ( .A(b[8]), .Y(n4642) );
  BUFX2 U2093 ( .A(b[5]), .Y(n4629) );
  BUFX2 U2094 ( .A(b[4]), .Y(n4625) );
  BUFX2 U2095 ( .A(b[6]), .Y(n4634) );
  BUFX2 U2096 ( .A(b[9]), .Y(n4647) );
  BUFX2 U2097 ( .A(b[6]), .Y(n4633) );
  BUFX2 U2098 ( .A(b[7]), .Y(n4638) );
  BUFX2 U2099 ( .A(b[8]), .Y(n4643) );
  BUFX2 U2100 ( .A(b[12]), .Y(n4660) );
  BUFX2 U2101 ( .A(b[15]), .Y(n4674) );
  BUFX2 U2102 ( .A(b[11]), .Y(n4655) );
  BUFX2 U2103 ( .A(b[14]), .Y(n4669) );
  BUFX2 U2104 ( .A(b[12]), .Y(n4661) );
  BUFX2 U2105 ( .A(b[14]), .Y(n4670) );
  BUFX2 U2106 ( .A(b[10]), .Y(n4651) );
  BUFX2 U2107 ( .A(b[11]), .Y(n4656) );
  BUFX2 U2108 ( .A(b[13]), .Y(n4665) );
  BUFX2 U2109 ( .A(b[9]), .Y(n4648) );
  BUFX2 U2110 ( .A(b[7]), .Y(n4639) );
  BUFX2 U2111 ( .A(b[8]), .Y(n4644) );
  BUFX2 U2112 ( .A(b[10]), .Y(n4653) );
  BUFX2 U2113 ( .A(b[11]), .Y(n4658) );
  BUFX2 U2114 ( .A(b[19]), .Y(n4694) );
  BUFX2 U2115 ( .A(b[12]), .Y(n4662) );
  BUFX2 U2116 ( .A(b[15]), .Y(n4676) );
  BUFX2 U2117 ( .A(b[10]), .Y(n4652) );
  BUFX2 U2118 ( .A(b[13]), .Y(n4666) );
  BUFX2 U2119 ( .A(b[11]), .Y(n4657) );
  BUFX2 U2120 ( .A(b[14]), .Y(n4671) );
  BUFX2 U2121 ( .A(b[17]), .Y(n4684) );
  BUFX2 U2122 ( .A(b[18]), .Y(n4689) );
  BUFX2 U2123 ( .A(b[15]), .Y(n4675) );
  BUFX2 U2124 ( .A(b[17]), .Y(n4685) );
  BUFX2 U2125 ( .A(b[18]), .Y(n4690) );
  BUFX2 U2126 ( .A(b[19]), .Y(n4695) );
  BUFX2 U2127 ( .A(b[20]), .Y(n4699) );
  BUFX2 U2128 ( .A(b[12]), .Y(n4663) );
  BUFX2 U2129 ( .A(b[14]), .Y(n4672) );
  BUFX2 U2130 ( .A(b[13]), .Y(n4667) );
  INVX2 U2131 ( .A(n4568), .Y(n4569) );
  INVX1 U2132 ( .A(b[24]), .Y(n4568) );
  BUFX2 U2133 ( .A(b[20]), .Y(n4698) );
  BUFX2 U2134 ( .A(b[21]), .Y(n4702) );
  BUFX2 U2135 ( .A(b[17]), .Y(n4686) );
  BUFX2 U2136 ( .A(b[18]), .Y(n4691) );
  BUFX2 U2137 ( .A(b[22]), .Y(n4706) );
  BUFX2 U2138 ( .A(b[19]), .Y(n4696) );
  BUFX2 U2139 ( .A(b[21]), .Y(n4704) );
  BUFX2 U2140 ( .A(b[20]), .Y(n4700) );
  BUFX2 U2141 ( .A(b[22]), .Y(n4707) );
  BUFX2 U2142 ( .A(b[23]), .Y(n4710) );
  BUFX2 U2143 ( .A(b[21]), .Y(n4703) );
  BUFX2 U2144 ( .A(b[22]), .Y(n4708) );
  BUFX2 U2145 ( .A(b[23]), .Y(n4711) );
  BUFX2 U2146 ( .A(b[15]), .Y(n4677) );
  BUFX2 U2147 ( .A(b[18]), .Y(n4692) );
  BUFX2 U2148 ( .A(b[17]), .Y(n4687) );
  BUFX2 U2149 ( .A(b[2]), .Y(n4612) );
  BUFX2 U2150 ( .A(b[3]), .Y(n4617) );
  BUFX2 U2151 ( .A(b[2]), .Y(n4613) );
  BUFX2 U2152 ( .A(b[3]), .Y(n4618) );
  BUFX2 U2153 ( .A(b[2]), .Y(n4614) );
  BUFX2 U2154 ( .A(b[3]), .Y(n4619) );
  BUFX2 U2155 ( .A(b[2]), .Y(n4615) );
  BUFX2 U2156 ( .A(b[3]), .Y(n4620) );
  INVX2 U2157 ( .A(n5526), .Y(n4570) );
  INVX2 U2158 ( .A(n5436), .Y(n4573) );
  INVX2 U2159 ( .A(n5437), .Y(n4575) );
  INVX2 U2160 ( .A(n4927), .Y(n4593) );
  INVX2 U2161 ( .A(n5030), .Y(n4589) );
  INVX2 U2162 ( .A(n5133), .Y(n4585) );
  INVX2 U2163 ( .A(n5236), .Y(n4581) );
  INVX2 U2164 ( .A(n5527), .Y(n4572) );
  INVX2 U2165 ( .A(n5024), .Y(n4590) );
  INVX2 U2166 ( .A(n5127), .Y(n4586) );
  INVX2 U2167 ( .A(n5230), .Y(n4582) );
  INVX2 U2168 ( .A(n5333), .Y(n4578) );
  INVX2 U2169 ( .A(n5134), .Y(n4583) );
  INVX2 U2170 ( .A(n5237), .Y(n4579) );
  INVX2 U2171 ( .A(n4928), .Y(n4591) );
  INVX2 U2172 ( .A(n5031), .Y(n4587) );
  INVX2 U2173 ( .A(n5679), .Y(n4770) );
  INVX2 U2174 ( .A(n5607), .Y(n4774) );
  INVX2 U2175 ( .A(n4559), .Y(n4597) );
  INVX2 U2176 ( .A(n4560), .Y(n4598) );
  INVX2 U2177 ( .A(n5608), .Y(n4775) );
  INVX2 U2178 ( .A(n5680), .Y(n4772) );
  INVX2 U2179 ( .A(n5740), .Y(n4767) );
  INVX2 U2180 ( .A(n5741), .Y(n4768) );
  INVX2 U2181 ( .A(n4561), .Y(n4601) );
  INVX2 U2182 ( .A(n4562), .Y(n4602) );
  INVX2 U2183 ( .A(n4563), .Y(n4603) );
  INVX2 U2184 ( .A(n4564), .Y(n4604) );
  INVX2 U2185 ( .A(n5600), .Y(n4571) );
  INVX2 U2186 ( .A(n5519), .Y(n4574) );
  INVX2 U2187 ( .A(n5672), .Y(n4567) );
  INVX2 U2188 ( .A(n4922), .Y(n4594) );
  INVX2 U2189 ( .A(n5429), .Y(n4576) );
  INVX2 U2190 ( .A(n2147), .Y(n4577) );
  AND2X1 U2191 ( .A(n4780), .B(n5431), .Y(n4559) );
  AND2X1 U2192 ( .A(n4778), .B(n5521), .Y(n4560) );
  INVX2 U2193 ( .A(n2132), .Y(n4595) );
  INVX2 U2194 ( .A(n5735), .Y(n4771) );
  AND2X1 U2195 ( .A(n4788), .B(n5019), .Y(n4561) );
  INVX2 U2196 ( .A(n2135), .Y(n4592) );
  INVX2 U2197 ( .A(n5772), .Y(n4766) );
  INVX2 U2198 ( .A(n2132), .Y(n4596) );
  INVX2 U2199 ( .A(n2138), .Y(n4588) );
  INVX2 U2200 ( .A(n2141), .Y(n4584) );
  INVX2 U2201 ( .A(n2144), .Y(n4580) );
  AND2X1 U2202 ( .A(n4786), .B(n5122), .Y(n4562) );
  AND2X1 U2203 ( .A(n4784), .B(n5225), .Y(n4563) );
  AND2X1 U2204 ( .A(n4782), .B(n5328), .Y(n4564) );
  INVX2 U2205 ( .A(n4565), .Y(n4600) );
  INVX2 U2206 ( .A(n4718), .Y(n4717) );
  INVX2 U2207 ( .A(n4716), .Y(n4715) );
  INVX2 U2208 ( .A(n4714), .Y(n4713) );
  INVX2 U2209 ( .A(n4720), .Y(n4719) );
  INVX2 U2210 ( .A(n4566), .Y(n4599) );
  AND2X1 U2211 ( .A(a[1]), .B(n4790), .Y(n4565) );
  INVX2 U2212 ( .A(n2150), .Y(n4720) );
  INVX2 U2213 ( .A(n2153), .Y(n4718) );
  INVX2 U2214 ( .A(n2156), .Y(n4716) );
  INVX2 U2215 ( .A(n2159), .Y(n4714) );
  AND2X1 U2216 ( .A(a[0]), .B(n4918), .Y(n4566) );
  BUFX2 U2217 ( .A(b[16]), .Y(n4679) );
  BUFX2 U2218 ( .A(b[16]), .Y(n4680) );
  BUFX2 U2219 ( .A(b[16]), .Y(n4681) );
  BUFX2 U2220 ( .A(b[16]), .Y(n4682) );
  INVX1 U2221 ( .A(b[26]), .Y(n4733) );
  INVX1 U2222 ( .A(b[28]), .Y(n4729) );
  BUFX2 U2223 ( .A(b[0]), .Y(n4608) );
  BUFX2 U2224 ( .A(b[0]), .Y(n4607) );
  BUFX2 U2225 ( .A(b[0]), .Y(n4606) );
  BUFX2 U2226 ( .A(b[0]), .Y(n4605) );
  INVX1 U2227 ( .A(b[27]), .Y(n4731) );
  INVX1 U2228 ( .A(b[25]), .Y(n4735) );
  INVX1 U2229 ( .A(b[31]), .Y(n4721) );
  INVX1 U2230 ( .A(b[30]), .Y(n4725) );
  INVX2 U2231 ( .A(n3301), .Y(n4722) );
  INVX2 U2232 ( .A(n3302), .Y(n4723) );
  INVX2 U2233 ( .A(n3303), .Y(n4724) );
  INVX2 U2234 ( .A(n3304), .Y(n4726) );
  INVX2 U2235 ( .A(n3305), .Y(n4728) );
  INVX2 U2236 ( .A(n3306), .Y(n4730) );
  INVX2 U2237 ( .A(n3307), .Y(n4732) );
  INVX2 U2238 ( .A(n3308), .Y(n4734) );
  INVX2 U2239 ( .A(n3309), .Y(n4736) );
  INVX2 U2240 ( .A(n3310), .Y(n4737) );
  INVX2 U2241 ( .A(n2429), .Y(n4747) );
  INVX2 U2242 ( .A(n2472), .Y(n4752) );
  INVX2 U2243 ( .A(n2520), .Y(n4756) );
  INVX2 U2244 ( .A(n5338), .Y(n4763) );
  INVX2 U2245 ( .A(n4827), .Y(n4764) );
  INVX2 U2246 ( .A(n5773), .Y(n4769) );
  INVX2 U2247 ( .A(n5736), .Y(n4773) );
  INVX2 U2248 ( .A(n5673), .Y(n4776) );
  INVX2 U2249 ( .A(n5603), .Y(n4777) );
  INVX2 U2250 ( .A(n5520), .Y(n4778) );
  INVX2 U2251 ( .A(n2147), .Y(n4779) );
  INVX2 U2252 ( .A(n5432), .Y(n4780) );
  INVX2 U2253 ( .A(n2144), .Y(n4781) );
  INVX2 U2254 ( .A(n5329), .Y(n4782) );
  INVX2 U2255 ( .A(n2141), .Y(n4783) );
  INVX2 U2256 ( .A(n5226), .Y(n4784) );
  INVX2 U2257 ( .A(n2138), .Y(n4785) );
  INVX2 U2258 ( .A(n5123), .Y(n4786) );
  INVX2 U2259 ( .A(n2135), .Y(n4787) );
  INVX2 U2260 ( .A(n5020), .Y(n4788) );
  INVX2 U2261 ( .A(a[1]), .Y(n4789) );
  INVX2 U2262 ( .A(a[0]), .Y(n4790) );
  XOR2X1 U2263 ( .A(n4791), .B(n4792), .Y(product[47]) );
  XOR2X1 U2264 ( .A(n4793), .B(n4794), .Y(n4792) );
  XOR2X1 U2265 ( .A(n2405), .B(n2352), .Y(n4794) );
  XOR2X1 U2266 ( .A(n2409), .B(n2407), .Y(n4793) );
  XOR2X1 U2267 ( .A(n4795), .B(n4796), .Y(n4791) );
  XOR2X1 U2268 ( .A(n4717), .B(n4719), .Y(n4796) );
  XOR2X1 U2269 ( .A(n4797), .B(n4798), .Y(n4795) );
  XOR2X1 U2270 ( .A(n4799), .B(n4800), .Y(n4798) );
  XOR2X1 U2271 ( .A(n4801), .B(n4802), .Y(n4800) );
  XOR2X1 U2272 ( .A(n4803), .B(n4804), .Y(n4802) );
  XOR2X1 U2273 ( .A(n2411), .B(n2159), .Y(n4804) );
  XOR2X1 U2274 ( .A(n2415), .B(n2413), .Y(n4803) );
  XOR2X1 U2275 ( .A(n4805), .B(n4806), .Y(n4801) );
  XOR2X1 U2276 ( .A(n4807), .B(n4808), .Y(n4806) );
  OAI21X1 U2277 ( .A(n4558), .B(n4744), .C(n4809), .Y(n4808) );
  OAI22X1 U2278 ( .A(n4677), .B(n4810), .C(n4766), .D(n4810), .Y(n4809) );
  OAI22X1 U2279 ( .A(n4767), .B(n4688), .C(n4768), .D(n4683), .Y(n4810) );
  OAI21X1 U2280 ( .A(n4557), .B(n4741), .C(n4811), .Y(n4807) );
  OAI22X1 U2281 ( .A(n4691), .B(n4812), .C(n4771), .D(n4812), .Y(n4811) );
  OAI22X1 U2282 ( .A(n4770), .B(n4701), .C(n4772), .D(n4697), .Y(n4812) );
  XOR2X1 U2283 ( .A(n4813), .B(n2156), .Y(n4805) );
  OAI21X1 U2284 ( .A(n4556), .B(n4738), .C(n4814), .Y(n4813) );
  OAI22X1 U2285 ( .A(n4704), .B(n4815), .C(n4567), .D(n4815), .Y(n4814) );
  OAI22X1 U2286 ( .A(n4774), .B(n4712), .C(n4775), .D(n4709), .Y(n4815) );
  OAI21X1 U2287 ( .A(n4555), .B(n4734), .C(n4816), .Y(n4799) );
  OAI22X1 U2288 ( .A(n4569), .B(n4817), .C(n4571), .D(n4817), .Y(n4816) );
  OAI22X1 U2289 ( .A(n4570), .B(n4733), .C(n4572), .D(n4735), .Y(n4817) );
  XOR2X1 U2290 ( .A(n4818), .B(n4819), .Y(n4797) );
  XNOR2X1 U2291 ( .A(n2147), .B(n4820), .Y(n4819) );
  OAI21X1 U2292 ( .A(n4597), .B(n4723), .C(n4821), .Y(n4820) );
  OAI22X1 U2293 ( .A(b[30]), .B(n4822), .C(n4576), .D(n4822), .Y(n4821) );
  NOR2X1 U2294 ( .A(n4721), .B(n4554), .Y(n4822) );
  OAI21X1 U2295 ( .A(n4598), .B(n4728), .C(n4823), .Y(n4818) );
  OAI22X1 U2296 ( .A(b[27]), .B(n4824), .C(n4574), .D(n4824), .Y(n4823) );
  OAI22X1 U2297 ( .A(n4573), .B(n4727), .C(n4575), .D(n4729), .Y(n4824) );
  XNOR2X1 U2298 ( .A(n4825), .B(n4595), .Y(n3661) );
  OAI22X1 U2299 ( .A(n4609), .B(n4553), .C(n4599), .D(n4609), .Y(n4825) );
  XNOR2X1 U2300 ( .A(n4826), .B(n4595), .Y(n3660) );
  OAI21X1 U2301 ( .A(n4599), .B(n4765), .C(n4764), .Y(n4826) );
  OAI22X1 U2302 ( .A(n4600), .B(n4609), .C(n4611), .D(n4553), .Y(n4827) );
  XNOR2X1 U2303 ( .A(n4828), .B(n4595), .Y(n3659) );
  OAI21X1 U2304 ( .A(n4599), .B(n4762), .C(n4829), .Y(n4828) );
  OAI22X1 U2305 ( .A(n4607), .B(n4830), .C(n4594), .D(n4830), .Y(n4829) );
  OAI22X1 U2306 ( .A(n4600), .B(n4611), .C(n4553), .D(n4616), .Y(n4830) );
  XNOR2X1 U2307 ( .A(n4831), .B(n4595), .Y(n3658) );
  OAI21X1 U2308 ( .A(n4599), .B(n4761), .C(n4832), .Y(n4831) );
  OAI22X1 U2309 ( .A(n4610), .B(n4833), .C(n4594), .D(n4833), .Y(n4832) );
  OAI22X1 U2310 ( .A(n4600), .B(n4616), .C(n4553), .D(n4621), .Y(n4833) );
  XNOR2X1 U2311 ( .A(n4834), .B(n4595), .Y(n3657) );
  OAI21X1 U2312 ( .A(n4599), .B(n4760), .C(n4835), .Y(n4834) );
  OAI22X1 U2313 ( .A(n4615), .B(n4836), .C(n4594), .D(n4836), .Y(n4835) );
  OAI22X1 U2314 ( .A(n4600), .B(n4621), .C(n4553), .D(n4626), .Y(n4836) );
  XNOR2X1 U2315 ( .A(n4837), .B(n4595), .Y(n3656) );
  OAI21X1 U2316 ( .A(n4599), .B(n4759), .C(n4838), .Y(n4837) );
  OAI22X1 U2317 ( .A(n4620), .B(n4839), .C(n4594), .D(n4839), .Y(n4838) );
  OAI22X1 U2318 ( .A(n4600), .B(n4626), .C(n4553), .D(n4630), .Y(n4839) );
  XNOR2X1 U2319 ( .A(n4840), .B(n4595), .Y(n3655) );
  OAI21X1 U2320 ( .A(n4599), .B(n4758), .C(n4841), .Y(n4840) );
  OAI22X1 U2321 ( .A(n4625), .B(n4842), .C(n4594), .D(n4842), .Y(n4841) );
  OAI22X1 U2322 ( .A(n4600), .B(n4630), .C(n4553), .D(n4635), .Y(n4842) );
  XNOR2X1 U2323 ( .A(n4843), .B(n4595), .Y(n3654) );
  OAI21X1 U2324 ( .A(n4599), .B(n4757), .C(n4844), .Y(n4843) );
  OAI22X1 U2325 ( .A(n4629), .B(n4845), .C(n4594), .D(n4845), .Y(n4844) );
  OAI22X1 U2326 ( .A(n4600), .B(n4635), .C(n4553), .D(n4640), .Y(n4845) );
  XNOR2X1 U2327 ( .A(n4846), .B(n4595), .Y(n3653) );
  OAI21X1 U2328 ( .A(n4599), .B(n4755), .C(n4847), .Y(n4846) );
  OAI22X1 U2329 ( .A(n4634), .B(n4848), .C(n4594), .D(n4848), .Y(n4847) );
  OAI22X1 U2330 ( .A(n4600), .B(n4640), .C(n4553), .D(n4645), .Y(n4848) );
  XNOR2X1 U2331 ( .A(n4849), .B(n4595), .Y(n3652) );
  OAI21X1 U2332 ( .A(n4599), .B(n4754), .C(n4850), .Y(n4849) );
  OAI22X1 U2333 ( .A(n4639), .B(n4851), .C(n4594), .D(n4851), .Y(n4850) );
  OAI22X1 U2334 ( .A(n4600), .B(n4645), .C(n4553), .D(n4649), .Y(n4851) );
  XNOR2X1 U2335 ( .A(n4852), .B(n4595), .Y(n3651) );
  OAI21X1 U2336 ( .A(n4599), .B(n4753), .C(n4853), .Y(n4852) );
  OAI22X1 U2337 ( .A(n4644), .B(n4854), .C(n4594), .D(n4854), .Y(n4853) );
  OAI22X1 U2338 ( .A(n4600), .B(n4649), .C(n4553), .D(n4654), .Y(n4854) );
  XNOR2X1 U2339 ( .A(n4855), .B(n4595), .Y(n3650) );
  OAI21X1 U2340 ( .A(n4599), .B(n4751), .C(n4856), .Y(n4855) );
  OAI22X1 U2341 ( .A(n4648), .B(n4857), .C(n4594), .D(n4857), .Y(n4856) );
  OAI22X1 U2342 ( .A(n4600), .B(n4654), .C(n4553), .D(n4659), .Y(n4857) );
  XNOR2X1 U2343 ( .A(n4858), .B(n4595), .Y(n3649) );
  OAI21X1 U2344 ( .A(n4599), .B(n4750), .C(n4859), .Y(n4858) );
  OAI22X1 U2345 ( .A(n4653), .B(n4860), .C(n4594), .D(n4860), .Y(n4859) );
  OAI22X1 U2346 ( .A(n4600), .B(n4659), .C(n4553), .D(n4664), .Y(n4860) );
  XNOR2X1 U2347 ( .A(n4861), .B(n4595), .Y(n3648) );
  OAI21X1 U2348 ( .A(n4599), .B(n4749), .C(n4862), .Y(n4861) );
  OAI22X1 U2349 ( .A(n4658), .B(n4863), .C(n4594), .D(n4863), .Y(n4862) );
  OAI22X1 U2350 ( .A(n4600), .B(n4664), .C(n4553), .D(n4668), .Y(n4863) );
  XNOR2X1 U2351 ( .A(n4864), .B(n4595), .Y(n3647) );
  OAI21X1 U2352 ( .A(n4599), .B(n4748), .C(n4865), .Y(n4864) );
  OAI22X1 U2353 ( .A(n4663), .B(n4866), .C(n4594), .D(n4866), .Y(n4865) );
  OAI22X1 U2354 ( .A(n4600), .B(n4668), .C(n4553), .D(n4673), .Y(n4866) );
  XNOR2X1 U2355 ( .A(n4867), .B(n4595), .Y(n3646) );
  OAI21X1 U2356 ( .A(n4599), .B(n4746), .C(n4868), .Y(n4867) );
  OAI22X1 U2357 ( .A(n4667), .B(n4869), .C(n4594), .D(n4869), .Y(n4868) );
  OAI22X1 U2358 ( .A(n4600), .B(n4673), .C(n4553), .D(n4678), .Y(n4869) );
  XNOR2X1 U2359 ( .A(n4870), .B(n4595), .Y(n3645) );
  OAI21X1 U2360 ( .A(n4599), .B(n4745), .C(n4871), .Y(n4870) );
  OAI22X1 U2361 ( .A(n4672), .B(n4872), .C(n4594), .D(n4872), .Y(n4871) );
  OAI22X1 U2362 ( .A(n4600), .B(n4678), .C(n4683), .D(n4553), .Y(n4872) );
  XNOR2X1 U2363 ( .A(n4873), .B(n4595), .Y(n3644) );
  OAI21X1 U2364 ( .A(n4744), .B(n4599), .C(n4874), .Y(n4873) );
  OAI22X1 U2365 ( .A(n4676), .B(n4875), .C(n4594), .D(n4875), .Y(n4874) );
  OAI22X1 U2366 ( .A(n4683), .B(n4600), .C(n4688), .D(n4553), .Y(n4875) );
  XNOR2X1 U2367 ( .A(n4876), .B(n4595), .Y(n3643) );
  OAI21X1 U2368 ( .A(n4599), .B(n4743), .C(n4877), .Y(n4876) );
  OAI22X1 U2369 ( .A(n4681), .B(n4878), .C(n4594), .D(n4878), .Y(n4877) );
  OAI22X1 U2370 ( .A(n4688), .B(n4600), .C(n4553), .D(n4693), .Y(n4878) );
  XNOR2X1 U2371 ( .A(n4879), .B(n4595), .Y(n3642) );
  OAI21X1 U2372 ( .A(n4599), .B(n4742), .C(n4880), .Y(n4879) );
  OAI22X1 U2373 ( .A(n4686), .B(n4881), .C(n4594), .D(n4881), .Y(n4880) );
  OAI22X1 U2374 ( .A(n4600), .B(n4693), .C(n4697), .D(n4553), .Y(n4881) );
  XNOR2X1 U2375 ( .A(n4882), .B(n4596), .Y(n3641) );
  OAI21X1 U2376 ( .A(n4741), .B(n4599), .C(n4883), .Y(n4882) );
  OAI22X1 U2377 ( .A(n4691), .B(n4884), .C(n4594), .D(n4884), .Y(n4883) );
  OAI22X1 U2378 ( .A(n4697), .B(n4600), .C(n4701), .D(n4553), .Y(n4884) );
  XNOR2X1 U2379 ( .A(n4885), .B(n4596), .Y(n3640) );
  OAI21X1 U2380 ( .A(n4599), .B(n4740), .C(n4886), .Y(n4885) );
  OAI22X1 U2381 ( .A(n4696), .B(n4887), .C(n4594), .D(n4887), .Y(n4886) );
  OAI22X1 U2382 ( .A(n4701), .B(n4600), .C(n4553), .D(n4705), .Y(n4887) );
  XNOR2X1 U2383 ( .A(n4888), .B(n4596), .Y(n3639) );
  OAI21X1 U2384 ( .A(n4599), .B(n4739), .C(n4889), .Y(n4888) );
  OAI22X1 U2385 ( .A(n4700), .B(n4890), .C(n4594), .D(n4890), .Y(n4889) );
  OAI22X1 U2386 ( .A(n4600), .B(n4705), .C(n4709), .D(n4553), .Y(n4890) );
  XNOR2X1 U2387 ( .A(n4891), .B(n4596), .Y(n3638) );
  OAI21X1 U2388 ( .A(n4738), .B(n4599), .C(n4892), .Y(n4891) );
  OAI22X1 U2389 ( .A(n4704), .B(n4893), .C(n4594), .D(n4893), .Y(n4892) );
  OAI22X1 U2390 ( .A(n4709), .B(n4600), .C(n4712), .D(n4553), .Y(n4893) );
  XNOR2X1 U2391 ( .A(n4894), .B(n4596), .Y(n3637) );
  OAI21X1 U2392 ( .A(n4599), .B(n4737), .C(n4895), .Y(n4894) );
  OAI22X1 U2393 ( .A(n4708), .B(n4896), .C(n4594), .D(n4896), .Y(n4895) );
  OAI22X1 U2394 ( .A(n4712), .B(n4600), .C(n4553), .D(n4568), .Y(n4896) );
  XNOR2X1 U2395 ( .A(n4897), .B(n4596), .Y(n3636) );
  OAI21X1 U2396 ( .A(n4599), .B(n4736), .C(n4898), .Y(n4897) );
  OAI22X1 U2397 ( .A(n4711), .B(n4899), .C(n4594), .D(n4899), .Y(n4898) );
  OAI22X1 U2398 ( .A(n4600), .B(n4568), .C(n4735), .D(n4553), .Y(n4899) );
  XNOR2X1 U2399 ( .A(n4900), .B(n4596), .Y(n3635) );
  OAI21X1 U2400 ( .A(n4734), .B(n4599), .C(n4901), .Y(n4900) );
  OAI22X1 U2401 ( .A(n4569), .B(n4902), .C(n4594), .D(n4902), .Y(n4901) );
  OAI22X1 U2402 ( .A(n4735), .B(n4600), .C(n4733), .D(n4553), .Y(n4902) );
  XNOR2X1 U2403 ( .A(n4903), .B(n4596), .Y(n3634) );
  OAI21X1 U2404 ( .A(n4599), .B(n4732), .C(n4904), .Y(n4903) );
  OAI22X1 U2405 ( .A(b[25]), .B(n4905), .C(n4594), .D(n4905), .Y(n4904) );
  OAI22X1 U2406 ( .A(n4733), .B(n4600), .C(n4553), .D(n4731), .Y(n4905) );
  XNOR2X1 U2407 ( .A(n4906), .B(n4596), .Y(n3633) );
  OAI21X1 U2408 ( .A(n4599), .B(n4730), .C(n4907), .Y(n4906) );
  OAI22X1 U2409 ( .A(b[26]), .B(n4908), .C(n4594), .D(n4908), .Y(n4907) );
  OAI22X1 U2410 ( .A(n4600), .B(n4731), .C(n4729), .D(n4553), .Y(n4908) );
  XNOR2X1 U2411 ( .A(n4909), .B(n4596), .Y(n3632) );
  OAI21X1 U2412 ( .A(n4728), .B(n4599), .C(n4910), .Y(n4909) );
  OAI22X1 U2413 ( .A(b[27]), .B(n4911), .C(n4594), .D(n4911), .Y(n4910) );
  OAI22X1 U2414 ( .A(n4729), .B(n4600), .C(n4727), .D(n4553), .Y(n4911) );
  XNOR2X1 U2415 ( .A(n4912), .B(n4596), .Y(n3631) );
  OAI21X1 U2416 ( .A(n4599), .B(n4726), .C(n4913), .Y(n4912) );
  OAI22X1 U2417 ( .A(b[28]), .B(n4914), .C(n4594), .D(n4914), .Y(n4913) );
  OAI22X1 U2418 ( .A(n4727), .B(n4600), .C(n4553), .D(n4725), .Y(n4914) );
  XNOR2X1 U2419 ( .A(n4915), .B(n4596), .Y(n3630) );
  OAI21X1 U2420 ( .A(n4599), .B(n4724), .C(n4916), .Y(n4915) );
  OAI22X1 U2421 ( .A(b[29]), .B(n4917), .C(n4594), .D(n4917), .Y(n4916) );
  OAI22X1 U2422 ( .A(n4600), .B(n4725), .C(n4721), .D(n4553), .Y(n4917) );
  XNOR2X1 U2423 ( .A(n4919), .B(n4596), .Y(n3629) );
  OAI21X1 U2424 ( .A(n4723), .B(n4599), .C(n4920), .Y(n4919) );
  OAI22X1 U2425 ( .A(b[30]), .B(n4921), .C(n4594), .D(n4921), .Y(n4920) );
  NOR2X1 U2426 ( .A(n4600), .B(n4721), .Y(n4921) );
  XNOR2X1 U2427 ( .A(n4923), .B(n4596), .Y(n3628) );
  OAI22X1 U2428 ( .A(n4721), .B(n4922), .C(n4599), .D(n4722), .Y(n4923) );
  NAND3X1 U2429 ( .A(n4918), .B(n4790), .C(n4789), .Y(n4922) );
  XNOR2X1 U2430 ( .A(a[1]), .B(n4596), .Y(n4918) );
  XNOR2X1 U2431 ( .A(n4924), .B(n4592), .Y(n3626) );
  OAI22X1 U2432 ( .A(n4609), .B(n4591), .C(n4609), .D(n4601), .Y(n4924) );
  XNOR2X1 U2433 ( .A(n4925), .B(n4787), .Y(n3625) );
  OAI21X1 U2434 ( .A(n4765), .B(n4601), .C(n4926), .Y(n4925) );
  AOI22X1 U2435 ( .A(n4927), .B(n4607), .C(n4928), .D(n4610), .Y(n4926) );
  XNOR2X1 U2436 ( .A(n4929), .B(n4787), .Y(n3624) );
  OAI21X1 U2437 ( .A(n4762), .B(n4601), .C(n4930), .Y(n4929) );
  OAI22X1 U2438 ( .A(n4607), .B(n4931), .C(n4590), .D(n4931), .Y(n4930) );
  OAI22X1 U2439 ( .A(n4611), .B(n4593), .C(n4616), .D(n4591), .Y(n4931) );
  XNOR2X1 U2440 ( .A(n4932), .B(n4787), .Y(n3623) );
  OAI21X1 U2441 ( .A(n4761), .B(n4601), .C(n4933), .Y(n4932) );
  OAI22X1 U2442 ( .A(n4610), .B(n4934), .C(n4590), .D(n4934), .Y(n4933) );
  OAI22X1 U2443 ( .A(n4616), .B(n4593), .C(n4621), .D(n4591), .Y(n4934) );
  XNOR2X1 U2444 ( .A(n4935), .B(n4787), .Y(n3622) );
  OAI21X1 U2445 ( .A(n4760), .B(n4601), .C(n4936), .Y(n4935) );
  OAI22X1 U2446 ( .A(n4614), .B(n4937), .C(n4590), .D(n4937), .Y(n4936) );
  OAI22X1 U2447 ( .A(n4621), .B(n4593), .C(n4626), .D(n4591), .Y(n4937) );
  XNOR2X1 U2448 ( .A(n4938), .B(n4787), .Y(n3621) );
  OAI21X1 U2449 ( .A(n4759), .B(n4601), .C(n4939), .Y(n4938) );
  OAI22X1 U2450 ( .A(n4619), .B(n4940), .C(n4590), .D(n4940), .Y(n4939) );
  OAI22X1 U2451 ( .A(n4626), .B(n4593), .C(n4630), .D(n4591), .Y(n4940) );
  XNOR2X1 U2452 ( .A(n4941), .B(n4787), .Y(n3620) );
  OAI21X1 U2453 ( .A(n4758), .B(n4601), .C(n4942), .Y(n4941) );
  OAI22X1 U2454 ( .A(n4624), .B(n4943), .C(n4590), .D(n4943), .Y(n4942) );
  OAI22X1 U2455 ( .A(n4630), .B(n4593), .C(n4635), .D(n4591), .Y(n4943) );
  XNOR2X1 U2456 ( .A(n4944), .B(n4787), .Y(n3619) );
  OAI21X1 U2457 ( .A(n4757), .B(n4601), .C(n4945), .Y(n4944) );
  OAI22X1 U2458 ( .A(n4628), .B(n4946), .C(n4590), .D(n4946), .Y(n4945) );
  OAI22X1 U2459 ( .A(n4635), .B(n4593), .C(n4640), .D(n4591), .Y(n4946) );
  XNOR2X1 U2460 ( .A(n4947), .B(n4787), .Y(n3618) );
  OAI21X1 U2461 ( .A(n4755), .B(n4601), .C(n4948), .Y(n4947) );
  OAI22X1 U2462 ( .A(n4633), .B(n4949), .C(n4590), .D(n4949), .Y(n4948) );
  OAI22X1 U2463 ( .A(n4640), .B(n4593), .C(n4645), .D(n4591), .Y(n4949) );
  XNOR2X1 U2464 ( .A(n4950), .B(n4787), .Y(n3617) );
  OAI21X1 U2465 ( .A(n4754), .B(n4601), .C(n4951), .Y(n4950) );
  OAI22X1 U2466 ( .A(n4638), .B(n4952), .C(n4590), .D(n4952), .Y(n4951) );
  OAI22X1 U2467 ( .A(n4645), .B(n4593), .C(n4649), .D(n4591), .Y(n4952) );
  XNOR2X1 U2468 ( .A(n4953), .B(n4787), .Y(n3616) );
  OAI21X1 U2469 ( .A(n4753), .B(n4601), .C(n4954), .Y(n4953) );
  OAI22X1 U2470 ( .A(n4643), .B(n4955), .C(n4590), .D(n4955), .Y(n4954) );
  OAI22X1 U2471 ( .A(n4649), .B(n4593), .C(n4654), .D(n4591), .Y(n4955) );
  XNOR2X1 U2472 ( .A(n4956), .B(n4787), .Y(n3615) );
  OAI21X1 U2473 ( .A(n4751), .B(n4601), .C(n4957), .Y(n4956) );
  OAI22X1 U2474 ( .A(n4647), .B(n4958), .C(n4590), .D(n4958), .Y(n4957) );
  OAI22X1 U2475 ( .A(n4654), .B(n4593), .C(n4659), .D(n4591), .Y(n4958) );
  XNOR2X1 U2476 ( .A(n4959), .B(n4787), .Y(n3614) );
  OAI21X1 U2477 ( .A(n4750), .B(n4601), .C(n4960), .Y(n4959) );
  OAI22X1 U2478 ( .A(n4652), .B(n4961), .C(n4590), .D(n4961), .Y(n4960) );
  OAI22X1 U2479 ( .A(n4659), .B(n4593), .C(n4664), .D(n4591), .Y(n4961) );
  XNOR2X1 U2480 ( .A(n4962), .B(n4787), .Y(n3613) );
  OAI21X1 U2481 ( .A(n4749), .B(n4601), .C(n4963), .Y(n4962) );
  OAI22X1 U2482 ( .A(n4657), .B(n4964), .C(n4590), .D(n4964), .Y(n4963) );
  OAI22X1 U2483 ( .A(n4664), .B(n4593), .C(n4668), .D(n4591), .Y(n4964) );
  XNOR2X1 U2484 ( .A(n4965), .B(n4787), .Y(n3612) );
  OAI21X1 U2485 ( .A(n4748), .B(n4601), .C(n4966), .Y(n4965) );
  OAI22X1 U2486 ( .A(n4662), .B(n4967), .C(n4590), .D(n4967), .Y(n4966) );
  OAI22X1 U2487 ( .A(n4668), .B(n4593), .C(n4673), .D(n4591), .Y(n4967) );
  XNOR2X1 U2488 ( .A(n4968), .B(n4787), .Y(n3611) );
  OAI21X1 U2489 ( .A(n4746), .B(n4601), .C(n4969), .Y(n4968) );
  OAI22X1 U2490 ( .A(n4666), .B(n4970), .C(n4590), .D(n4970), .Y(n4969) );
  OAI22X1 U2491 ( .A(n4673), .B(n4593), .C(n4678), .D(n4591), .Y(n4970) );
  XNOR2X1 U2492 ( .A(n4971), .B(n4787), .Y(n3610) );
  OAI21X1 U2493 ( .A(n4745), .B(n4601), .C(n4972), .Y(n4971) );
  OAI22X1 U2494 ( .A(n4671), .B(n4973), .C(n4590), .D(n4973), .Y(n4972) );
  OAI22X1 U2495 ( .A(n4678), .B(n4593), .C(n4683), .D(n4591), .Y(n4973) );
  XNOR2X1 U2496 ( .A(n4974), .B(n4787), .Y(n3609) );
  OAI21X1 U2497 ( .A(n4744), .B(n4601), .C(n4975), .Y(n4974) );
  OAI22X1 U2498 ( .A(n4676), .B(n4976), .C(n4590), .D(n4976), .Y(n4975) );
  OAI22X1 U2499 ( .A(n4683), .B(n4593), .C(n4688), .D(n4591), .Y(n4976) );
  XNOR2X1 U2500 ( .A(n4977), .B(n4787), .Y(n3608) );
  OAI21X1 U2501 ( .A(n4743), .B(n4601), .C(n4978), .Y(n4977) );
  OAI22X1 U2502 ( .A(n4681), .B(n4979), .C(n4590), .D(n4979), .Y(n4978) );
  OAI22X1 U2503 ( .A(n4688), .B(n4593), .C(n4693), .D(n4591), .Y(n4979) );
  XNOR2X1 U2504 ( .A(n4980), .B(n4592), .Y(n3607) );
  OAI21X1 U2505 ( .A(n4742), .B(n4601), .C(n4981), .Y(n4980) );
  OAI22X1 U2506 ( .A(n4686), .B(n4982), .C(n4590), .D(n4982), .Y(n4981) );
  OAI22X1 U2507 ( .A(n4693), .B(n4593), .C(n4697), .D(n4591), .Y(n4982) );
  XNOR2X1 U2508 ( .A(n4983), .B(n4592), .Y(n3606) );
  OAI21X1 U2509 ( .A(n4741), .B(n4601), .C(n4984), .Y(n4983) );
  OAI22X1 U2510 ( .A(n4691), .B(n4985), .C(n4590), .D(n4985), .Y(n4984) );
  OAI22X1 U2511 ( .A(n4697), .B(n4593), .C(n4701), .D(n4591), .Y(n4985) );
  XNOR2X1 U2512 ( .A(n4986), .B(n4592), .Y(n3605) );
  OAI21X1 U2513 ( .A(n4740), .B(n4601), .C(n4987), .Y(n4986) );
  OAI22X1 U2514 ( .A(n4696), .B(n4988), .C(n4590), .D(n4988), .Y(n4987) );
  OAI22X1 U2515 ( .A(n4701), .B(n4593), .C(n4705), .D(n4591), .Y(n4988) );
  XNOR2X1 U2516 ( .A(n4989), .B(n4592), .Y(n3604) );
  OAI21X1 U2517 ( .A(n4739), .B(n4601), .C(n4990), .Y(n4989) );
  OAI22X1 U2518 ( .A(n4700), .B(n4991), .C(n4590), .D(n4991), .Y(n4990) );
  OAI22X1 U2519 ( .A(n4705), .B(n4593), .C(n4709), .D(n4591), .Y(n4991) );
  XNOR2X1 U2520 ( .A(n4992), .B(n4592), .Y(n3603) );
  OAI21X1 U2521 ( .A(n4738), .B(n4601), .C(n4993), .Y(n4992) );
  OAI22X1 U2522 ( .A(n4704), .B(n4994), .C(n4590), .D(n4994), .Y(n4993) );
  OAI22X1 U2523 ( .A(n4709), .B(n4593), .C(n4712), .D(n4591), .Y(n4994) );
  XNOR2X1 U2524 ( .A(n4995), .B(n4592), .Y(n3602) );
  OAI21X1 U2525 ( .A(n4737), .B(n4601), .C(n4996), .Y(n4995) );
  OAI22X1 U2526 ( .A(n4708), .B(n4997), .C(n4590), .D(n4997), .Y(n4996) );
  OAI22X1 U2527 ( .A(n4712), .B(n4593), .C(n4568), .D(n4591), .Y(n4997) );
  XNOR2X1 U2528 ( .A(n4998), .B(n4592), .Y(n3601) );
  OAI21X1 U2529 ( .A(n4736), .B(n4601), .C(n4999), .Y(n4998) );
  OAI22X1 U2530 ( .A(n4711), .B(n5000), .C(n4590), .D(n5000), .Y(n4999) );
  OAI22X1 U2531 ( .A(n4568), .B(n4593), .C(n4735), .D(n4591), .Y(n5000) );
  XNOR2X1 U2532 ( .A(n5001), .B(n4592), .Y(n3600) );
  OAI21X1 U2533 ( .A(n4734), .B(n4601), .C(n5002), .Y(n5001) );
  OAI22X1 U2534 ( .A(n4569), .B(n5003), .C(n4590), .D(n5003), .Y(n5002) );
  OAI22X1 U2535 ( .A(n4735), .B(n4593), .C(n4733), .D(n4591), .Y(n5003) );
  XNOR2X1 U2536 ( .A(n5004), .B(n4592), .Y(n3599) );
  OAI21X1 U2537 ( .A(n4732), .B(n4601), .C(n5005), .Y(n5004) );
  OAI22X1 U2538 ( .A(b[25]), .B(n5006), .C(n4590), .D(n5006), .Y(n5005) );
  OAI22X1 U2539 ( .A(n4733), .B(n4593), .C(n4731), .D(n4591), .Y(n5006) );
  XNOR2X1 U2540 ( .A(n5007), .B(n4592), .Y(n3598) );
  OAI21X1 U2541 ( .A(n4730), .B(n4601), .C(n5008), .Y(n5007) );
  OAI22X1 U2542 ( .A(b[26]), .B(n5009), .C(n4590), .D(n5009), .Y(n5008) );
  OAI22X1 U2543 ( .A(n4731), .B(n4593), .C(n4729), .D(n4591), .Y(n5009) );
  XNOR2X1 U2544 ( .A(n5010), .B(n4592), .Y(n3597) );
  OAI21X1 U2545 ( .A(n4728), .B(n4601), .C(n5011), .Y(n5010) );
  OAI22X1 U2546 ( .A(b[27]), .B(n5012), .C(n4590), .D(n5012), .Y(n5011) );
  OAI22X1 U2547 ( .A(n4729), .B(n4593), .C(n4727), .D(n4591), .Y(n5012) );
  XNOR2X1 U2548 ( .A(n5013), .B(n4592), .Y(n3596) );
  OAI21X1 U2549 ( .A(n4726), .B(n4601), .C(n5014), .Y(n5013) );
  OAI22X1 U2550 ( .A(b[28]), .B(n5015), .C(n4590), .D(n5015), .Y(n5014) );
  OAI22X1 U2551 ( .A(n4727), .B(n4593), .C(n4725), .D(n4591), .Y(n5015) );
  XNOR2X1 U2552 ( .A(n5016), .B(n4592), .Y(n3595) );
  OAI21X1 U2553 ( .A(n4724), .B(n4601), .C(n5017), .Y(n5016) );
  OAI22X1 U2554 ( .A(b[29]), .B(n5018), .C(n4590), .D(n5018), .Y(n5017) );
  OAI22X1 U2555 ( .A(n4725), .B(n4593), .C(n4721), .D(n4591), .Y(n5018) );
  NOR2X1 U2556 ( .A(n5019), .B(n5020), .Y(n4928) );
  XNOR2X1 U2557 ( .A(n5021), .B(n4592), .Y(n3594) );
  OAI21X1 U2558 ( .A(n4723), .B(n4601), .C(n5022), .Y(n5021) );
  OAI22X1 U2559 ( .A(b[30]), .B(n5023), .C(n4590), .D(n5023), .Y(n5022) );
  NOR2X1 U2560 ( .A(n4593), .B(n4721), .Y(n5023) );
  NOR2X1 U2561 ( .A(n4788), .B(n5025), .Y(n4927) );
  XNOR2X1 U2562 ( .A(n5026), .B(n4592), .Y(n3593) );
  OAI22X1 U2563 ( .A(n4721), .B(n5024), .C(n4722), .D(n4601), .Y(n5026) );
  NAND3X1 U2564 ( .A(n5020), .B(n5019), .C(n5025), .Y(n5024) );
  XNOR2X1 U2565 ( .A(a[3]), .B(a[4]), .Y(n5025) );
  XNOR2X1 U2566 ( .A(a[4]), .B(n4592), .Y(n5019) );
  XOR2X1 U2567 ( .A(a[3]), .B(n4596), .Y(n5020) );
  XNOR2X1 U2568 ( .A(n5027), .B(n4588), .Y(n3591) );
  OAI22X1 U2569 ( .A(n4609), .B(n4587), .C(n4609), .D(n4602), .Y(n5027) );
  XNOR2X1 U2570 ( .A(n5028), .B(n4785), .Y(n3590) );
  OAI21X1 U2571 ( .A(n4765), .B(n4602), .C(n5029), .Y(n5028) );
  AOI22X1 U2572 ( .A(n5030), .B(n4607), .C(n5031), .D(n4610), .Y(n5029) );
  XNOR2X1 U2573 ( .A(n5032), .B(n4785), .Y(n3589) );
  OAI21X1 U2574 ( .A(n4762), .B(n4602), .C(n5033), .Y(n5032) );
  OAI22X1 U2575 ( .A(n4607), .B(n5034), .C(n4586), .D(n5034), .Y(n5033) );
  OAI22X1 U2576 ( .A(n4611), .B(n4589), .C(n4616), .D(n4587), .Y(n5034) );
  XNOR2X1 U2577 ( .A(n5035), .B(n4785), .Y(n3588) );
  OAI21X1 U2578 ( .A(n4761), .B(n4602), .C(n5036), .Y(n5035) );
  OAI22X1 U2579 ( .A(n4610), .B(n5037), .C(n4586), .D(n5037), .Y(n5036) );
  OAI22X1 U2580 ( .A(n4616), .B(n4589), .C(n4621), .D(n4587), .Y(n5037) );
  XNOR2X1 U2581 ( .A(n5038), .B(n4785), .Y(n3587) );
  OAI21X1 U2582 ( .A(n4760), .B(n4602), .C(n5039), .Y(n5038) );
  OAI22X1 U2583 ( .A(n4614), .B(n5040), .C(n4586), .D(n5040), .Y(n5039) );
  OAI22X1 U2584 ( .A(n4621), .B(n4589), .C(n4626), .D(n4587), .Y(n5040) );
  XNOR2X1 U2585 ( .A(n5041), .B(n4785), .Y(n3586) );
  OAI21X1 U2586 ( .A(n4759), .B(n4602), .C(n5042), .Y(n5041) );
  OAI22X1 U2587 ( .A(n4619), .B(n5043), .C(n4586), .D(n5043), .Y(n5042) );
  OAI22X1 U2588 ( .A(n4626), .B(n4589), .C(n4630), .D(n4587), .Y(n5043) );
  XNOR2X1 U2589 ( .A(n5044), .B(n4785), .Y(n3585) );
  OAI21X1 U2590 ( .A(n4758), .B(n4602), .C(n5045), .Y(n5044) );
  OAI22X1 U2591 ( .A(n4624), .B(n5046), .C(n4586), .D(n5046), .Y(n5045) );
  OAI22X1 U2592 ( .A(n4630), .B(n4589), .C(n4635), .D(n4587), .Y(n5046) );
  XNOR2X1 U2593 ( .A(n5047), .B(n4785), .Y(n3584) );
  OAI21X1 U2594 ( .A(n4757), .B(n4602), .C(n5048), .Y(n5047) );
  OAI22X1 U2595 ( .A(n4628), .B(n5049), .C(n4586), .D(n5049), .Y(n5048) );
  OAI22X1 U2596 ( .A(n4635), .B(n4589), .C(n4640), .D(n4587), .Y(n5049) );
  XNOR2X1 U2597 ( .A(n5050), .B(n4785), .Y(n3583) );
  OAI21X1 U2598 ( .A(n4755), .B(n4602), .C(n5051), .Y(n5050) );
  OAI22X1 U2599 ( .A(n4633), .B(n5052), .C(n4586), .D(n5052), .Y(n5051) );
  OAI22X1 U2600 ( .A(n4640), .B(n4589), .C(n4645), .D(n4587), .Y(n5052) );
  XNOR2X1 U2601 ( .A(n5053), .B(n4785), .Y(n3582) );
  OAI21X1 U2602 ( .A(n4754), .B(n4602), .C(n5054), .Y(n5053) );
  OAI22X1 U2603 ( .A(n4638), .B(n5055), .C(n4586), .D(n5055), .Y(n5054) );
  OAI22X1 U2604 ( .A(n4645), .B(n4589), .C(n4649), .D(n4587), .Y(n5055) );
  XNOR2X1 U2605 ( .A(n5056), .B(n4785), .Y(n3581) );
  OAI21X1 U2606 ( .A(n4753), .B(n4602), .C(n5057), .Y(n5056) );
  OAI22X1 U2607 ( .A(n4643), .B(n5058), .C(n4586), .D(n5058), .Y(n5057) );
  OAI22X1 U2608 ( .A(n4649), .B(n4589), .C(n4654), .D(n4587), .Y(n5058) );
  XNOR2X1 U2609 ( .A(n5059), .B(n4785), .Y(n3580) );
  OAI21X1 U2610 ( .A(n4751), .B(n4602), .C(n5060), .Y(n5059) );
  OAI22X1 U2611 ( .A(n4647), .B(n5061), .C(n4586), .D(n5061), .Y(n5060) );
  OAI22X1 U2612 ( .A(n4654), .B(n4589), .C(n4659), .D(n4587), .Y(n5061) );
  XNOR2X1 U2613 ( .A(n5062), .B(n4785), .Y(n3579) );
  OAI21X1 U2614 ( .A(n4750), .B(n4602), .C(n5063), .Y(n5062) );
  OAI22X1 U2615 ( .A(n4652), .B(n5064), .C(n4586), .D(n5064), .Y(n5063) );
  OAI22X1 U2616 ( .A(n4659), .B(n4589), .C(n4664), .D(n4587), .Y(n5064) );
  XNOR2X1 U2617 ( .A(n5065), .B(n4785), .Y(n3578) );
  OAI21X1 U2618 ( .A(n4749), .B(n4602), .C(n5066), .Y(n5065) );
  OAI22X1 U2619 ( .A(n4657), .B(n5067), .C(n4586), .D(n5067), .Y(n5066) );
  OAI22X1 U2620 ( .A(n4664), .B(n4589), .C(n4668), .D(n4587), .Y(n5067) );
  XNOR2X1 U2621 ( .A(n5068), .B(n4785), .Y(n3577) );
  OAI21X1 U2622 ( .A(n4748), .B(n4602), .C(n5069), .Y(n5068) );
  OAI22X1 U2623 ( .A(n4662), .B(n5070), .C(n4586), .D(n5070), .Y(n5069) );
  OAI22X1 U2624 ( .A(n4668), .B(n4589), .C(n4673), .D(n4587), .Y(n5070) );
  XNOR2X1 U2625 ( .A(n5071), .B(n4785), .Y(n3576) );
  OAI21X1 U2626 ( .A(n4746), .B(n4602), .C(n5072), .Y(n5071) );
  OAI22X1 U2627 ( .A(n4666), .B(n5073), .C(n4586), .D(n5073), .Y(n5072) );
  OAI22X1 U2628 ( .A(n4673), .B(n4589), .C(n4678), .D(n4587), .Y(n5073) );
  XNOR2X1 U2629 ( .A(n5074), .B(n4785), .Y(n3575) );
  OAI21X1 U2630 ( .A(n4745), .B(n4602), .C(n5075), .Y(n5074) );
  OAI22X1 U2631 ( .A(n4671), .B(n5076), .C(n4586), .D(n5076), .Y(n5075) );
  OAI22X1 U2632 ( .A(n4678), .B(n4589), .C(n4683), .D(n4587), .Y(n5076) );
  XNOR2X1 U2633 ( .A(n5077), .B(n4785), .Y(n3574) );
  OAI21X1 U2634 ( .A(n4744), .B(n4602), .C(n5078), .Y(n5077) );
  OAI22X1 U2635 ( .A(n4676), .B(n5079), .C(n4586), .D(n5079), .Y(n5078) );
  OAI22X1 U2636 ( .A(n4683), .B(n4589), .C(n4688), .D(n4587), .Y(n5079) );
  XNOR2X1 U2637 ( .A(n5080), .B(n4785), .Y(n3573) );
  OAI21X1 U2638 ( .A(n4743), .B(n4602), .C(n5081), .Y(n5080) );
  OAI22X1 U2639 ( .A(n4681), .B(n5082), .C(n4586), .D(n5082), .Y(n5081) );
  OAI22X1 U2640 ( .A(n4688), .B(n4589), .C(n4693), .D(n4587), .Y(n5082) );
  XNOR2X1 U2641 ( .A(n5083), .B(n4785), .Y(n3572) );
  OAI21X1 U2642 ( .A(n4742), .B(n4602), .C(n5084), .Y(n5083) );
  OAI22X1 U2643 ( .A(n4686), .B(n5085), .C(n4586), .D(n5085), .Y(n5084) );
  OAI22X1 U2644 ( .A(n4693), .B(n4589), .C(n4697), .D(n4587), .Y(n5085) );
  XNOR2X1 U2645 ( .A(n5086), .B(n4588), .Y(n3571) );
  OAI21X1 U2646 ( .A(n4741), .B(n4602), .C(n5087), .Y(n5086) );
  OAI22X1 U2647 ( .A(n4691), .B(n5088), .C(n4586), .D(n5088), .Y(n5087) );
  OAI22X1 U2648 ( .A(n4697), .B(n4589), .C(n4701), .D(n4587), .Y(n5088) );
  XNOR2X1 U2649 ( .A(n5089), .B(n4588), .Y(n3570) );
  OAI21X1 U2650 ( .A(n4740), .B(n4602), .C(n5090), .Y(n5089) );
  OAI22X1 U2651 ( .A(n4696), .B(n5091), .C(n4586), .D(n5091), .Y(n5090) );
  OAI22X1 U2652 ( .A(n4701), .B(n4589), .C(n4705), .D(n4587), .Y(n5091) );
  XNOR2X1 U2653 ( .A(n5092), .B(n4588), .Y(n3569) );
  OAI21X1 U2654 ( .A(n4739), .B(n4602), .C(n5093), .Y(n5092) );
  OAI22X1 U2655 ( .A(n4700), .B(n5094), .C(n4586), .D(n5094), .Y(n5093) );
  OAI22X1 U2656 ( .A(n4705), .B(n4589), .C(n4709), .D(n4587), .Y(n5094) );
  XNOR2X1 U2657 ( .A(n5095), .B(n4588), .Y(n3568) );
  OAI21X1 U2658 ( .A(n4738), .B(n4602), .C(n5096), .Y(n5095) );
  OAI22X1 U2659 ( .A(n4704), .B(n5097), .C(n4586), .D(n5097), .Y(n5096) );
  OAI22X1 U2660 ( .A(n4709), .B(n4589), .C(n4712), .D(n4587), .Y(n5097) );
  XNOR2X1 U2661 ( .A(n5098), .B(n4588), .Y(n3567) );
  OAI21X1 U2662 ( .A(n4737), .B(n4602), .C(n5099), .Y(n5098) );
  OAI22X1 U2663 ( .A(n4708), .B(n5100), .C(n4586), .D(n5100), .Y(n5099) );
  OAI22X1 U2664 ( .A(n4712), .B(n4589), .C(n4568), .D(n4587), .Y(n5100) );
  XNOR2X1 U2665 ( .A(n5101), .B(n4588), .Y(n3566) );
  OAI21X1 U2666 ( .A(n4736), .B(n4602), .C(n5102), .Y(n5101) );
  OAI22X1 U2667 ( .A(n4711), .B(n5103), .C(n4586), .D(n5103), .Y(n5102) );
  OAI22X1 U2668 ( .A(n4568), .B(n4589), .C(n4735), .D(n4587), .Y(n5103) );
  XNOR2X1 U2669 ( .A(n5104), .B(n4588), .Y(n3565) );
  OAI21X1 U2670 ( .A(n4734), .B(n4602), .C(n5105), .Y(n5104) );
  OAI22X1 U2671 ( .A(n4569), .B(n5106), .C(n4586), .D(n5106), .Y(n5105) );
  OAI22X1 U2672 ( .A(n4735), .B(n4589), .C(n4733), .D(n4587), .Y(n5106) );
  XNOR2X1 U2673 ( .A(n5107), .B(n4588), .Y(n3564) );
  OAI21X1 U2674 ( .A(n4732), .B(n4602), .C(n5108), .Y(n5107) );
  OAI22X1 U2675 ( .A(b[25]), .B(n5109), .C(n4586), .D(n5109), .Y(n5108) );
  OAI22X1 U2676 ( .A(n4733), .B(n4589), .C(n4731), .D(n4587), .Y(n5109) );
  XNOR2X1 U2677 ( .A(n5110), .B(n4588), .Y(n3563) );
  OAI21X1 U2678 ( .A(n4730), .B(n4602), .C(n5111), .Y(n5110) );
  OAI22X1 U2679 ( .A(b[26]), .B(n5112), .C(n4586), .D(n5112), .Y(n5111) );
  OAI22X1 U2680 ( .A(n4731), .B(n4589), .C(n4729), .D(n4587), .Y(n5112) );
  XNOR2X1 U2681 ( .A(n5113), .B(n4588), .Y(n3562) );
  OAI21X1 U2682 ( .A(n4728), .B(n4602), .C(n5114), .Y(n5113) );
  OAI22X1 U2683 ( .A(b[27]), .B(n5115), .C(n4586), .D(n5115), .Y(n5114) );
  OAI22X1 U2684 ( .A(n4729), .B(n4589), .C(n4727), .D(n4587), .Y(n5115) );
  XNOR2X1 U2685 ( .A(n5116), .B(n4588), .Y(n3561) );
  OAI21X1 U2686 ( .A(n4726), .B(n4602), .C(n5117), .Y(n5116) );
  OAI22X1 U2687 ( .A(b[28]), .B(n5118), .C(n4586), .D(n5118), .Y(n5117) );
  OAI22X1 U2688 ( .A(n4727), .B(n4589), .C(n4725), .D(n4587), .Y(n5118) );
  XNOR2X1 U2689 ( .A(n5119), .B(n4588), .Y(n3560) );
  OAI21X1 U2690 ( .A(n4724), .B(n4602), .C(n5120), .Y(n5119) );
  OAI22X1 U2691 ( .A(b[29]), .B(n5121), .C(n4586), .D(n5121), .Y(n5120) );
  OAI22X1 U2692 ( .A(n4725), .B(n4589), .C(n4721), .D(n4587), .Y(n5121) );
  NOR2X1 U2693 ( .A(n5122), .B(n5123), .Y(n5031) );
  XNOR2X1 U2694 ( .A(n5124), .B(n4588), .Y(n3559) );
  OAI21X1 U2695 ( .A(n4723), .B(n4602), .C(n5125), .Y(n5124) );
  OAI22X1 U2696 ( .A(b[30]), .B(n5126), .C(n4586), .D(n5126), .Y(n5125) );
  NOR2X1 U2697 ( .A(n4589), .B(n4721), .Y(n5126) );
  NOR2X1 U2698 ( .A(n4786), .B(n5128), .Y(n5030) );
  XNOR2X1 U2699 ( .A(n5129), .B(n4588), .Y(n3558) );
  OAI22X1 U2700 ( .A(n4721), .B(n5127), .C(n4722), .D(n4602), .Y(n5129) );
  NAND3X1 U2701 ( .A(n5123), .B(n5122), .C(n5128), .Y(n5127) );
  XNOR2X1 U2702 ( .A(a[6]), .B(a[7]), .Y(n5128) );
  XNOR2X1 U2703 ( .A(a[7]), .B(n4588), .Y(n5122) );
  XOR2X1 U2704 ( .A(a[6]), .B(n4592), .Y(n5123) );
  XNOR2X1 U2705 ( .A(n5130), .B(n4584), .Y(n3556) );
  OAI22X1 U2706 ( .A(n4609), .B(n4583), .C(n4609), .D(n4603), .Y(n5130) );
  XNOR2X1 U2707 ( .A(n5131), .B(n4783), .Y(n3555) );
  OAI21X1 U2708 ( .A(n4765), .B(n4603), .C(n5132), .Y(n5131) );
  AOI22X1 U2709 ( .A(n5133), .B(n4607), .C(n5134), .D(n4610), .Y(n5132) );
  XNOR2X1 U2710 ( .A(n5135), .B(n4783), .Y(n3554) );
  OAI21X1 U2711 ( .A(n4762), .B(n4603), .C(n5136), .Y(n5135) );
  OAI22X1 U2712 ( .A(n4608), .B(n5137), .C(n4582), .D(n5137), .Y(n5136) );
  OAI22X1 U2713 ( .A(n4611), .B(n4585), .C(n4616), .D(n4583), .Y(n5137) );
  XNOR2X1 U2714 ( .A(n5138), .B(n4783), .Y(n3553) );
  OAI21X1 U2715 ( .A(n4761), .B(n4603), .C(n5139), .Y(n5138) );
  OAI22X1 U2716 ( .A(n4610), .B(n5140), .C(n4582), .D(n5140), .Y(n5139) );
  OAI22X1 U2717 ( .A(n4616), .B(n4585), .C(n4621), .D(n4583), .Y(n5140) );
  XNOR2X1 U2718 ( .A(n5141), .B(n4783), .Y(n3552) );
  OAI21X1 U2719 ( .A(n4760), .B(n4603), .C(n5142), .Y(n5141) );
  OAI22X1 U2720 ( .A(n4614), .B(n5143), .C(n4582), .D(n5143), .Y(n5142) );
  OAI22X1 U2721 ( .A(n4621), .B(n4585), .C(n4626), .D(n4583), .Y(n5143) );
  XNOR2X1 U2722 ( .A(n5144), .B(n4783), .Y(n3551) );
  OAI21X1 U2723 ( .A(n4759), .B(n4603), .C(n5145), .Y(n5144) );
  OAI22X1 U2724 ( .A(n4619), .B(n5146), .C(n4582), .D(n5146), .Y(n5145) );
  OAI22X1 U2725 ( .A(n4626), .B(n4585), .C(n4630), .D(n4583), .Y(n5146) );
  XNOR2X1 U2726 ( .A(n5147), .B(n4783), .Y(n3550) );
  OAI21X1 U2727 ( .A(n4758), .B(n4603), .C(n5148), .Y(n5147) );
  OAI22X1 U2728 ( .A(n4624), .B(n5149), .C(n4582), .D(n5149), .Y(n5148) );
  OAI22X1 U2729 ( .A(n4630), .B(n4585), .C(n4635), .D(n4583), .Y(n5149) );
  XNOR2X1 U2730 ( .A(n5150), .B(n4783), .Y(n3549) );
  OAI21X1 U2731 ( .A(n4757), .B(n4603), .C(n5151), .Y(n5150) );
  OAI22X1 U2732 ( .A(n4628), .B(n5152), .C(n4582), .D(n5152), .Y(n5151) );
  OAI22X1 U2733 ( .A(n4635), .B(n4585), .C(n4640), .D(n4583), .Y(n5152) );
  XNOR2X1 U2734 ( .A(n5153), .B(n4783), .Y(n3548) );
  OAI21X1 U2735 ( .A(n4755), .B(n4603), .C(n5154), .Y(n5153) );
  OAI22X1 U2736 ( .A(n4633), .B(n5155), .C(n4582), .D(n5155), .Y(n5154) );
  OAI22X1 U2737 ( .A(n4640), .B(n4585), .C(n4645), .D(n4583), .Y(n5155) );
  XNOR2X1 U2738 ( .A(n5156), .B(n4783), .Y(n3547) );
  OAI21X1 U2739 ( .A(n4754), .B(n4603), .C(n5157), .Y(n5156) );
  OAI22X1 U2740 ( .A(n4638), .B(n5158), .C(n4582), .D(n5158), .Y(n5157) );
  OAI22X1 U2741 ( .A(n4645), .B(n4585), .C(n4649), .D(n4583), .Y(n5158) );
  XNOR2X1 U2742 ( .A(n5159), .B(n4783), .Y(n3546) );
  OAI21X1 U2743 ( .A(n4753), .B(n4603), .C(n5160), .Y(n5159) );
  OAI22X1 U2744 ( .A(n4643), .B(n5161), .C(n4582), .D(n5161), .Y(n5160) );
  OAI22X1 U2745 ( .A(n4649), .B(n4585), .C(n4654), .D(n4583), .Y(n5161) );
  XNOR2X1 U2746 ( .A(n5162), .B(n4783), .Y(n3545) );
  OAI21X1 U2747 ( .A(n4751), .B(n4603), .C(n5163), .Y(n5162) );
  OAI22X1 U2748 ( .A(n4647), .B(n5164), .C(n4582), .D(n5164), .Y(n5163) );
  OAI22X1 U2749 ( .A(n4654), .B(n4585), .C(n4659), .D(n4583), .Y(n5164) );
  XNOR2X1 U2750 ( .A(n5165), .B(n4783), .Y(n3544) );
  OAI21X1 U2751 ( .A(n4750), .B(n4603), .C(n5166), .Y(n5165) );
  OAI22X1 U2752 ( .A(n4652), .B(n5167), .C(n4582), .D(n5167), .Y(n5166) );
  OAI22X1 U2753 ( .A(n4659), .B(n4585), .C(n4664), .D(n4583), .Y(n5167) );
  XNOR2X1 U2754 ( .A(n5168), .B(n4783), .Y(n3543) );
  OAI21X1 U2755 ( .A(n4749), .B(n4603), .C(n5169), .Y(n5168) );
  OAI22X1 U2756 ( .A(n4657), .B(n5170), .C(n4582), .D(n5170), .Y(n5169) );
  OAI22X1 U2757 ( .A(n4664), .B(n4585), .C(n4668), .D(n4583), .Y(n5170) );
  XNOR2X1 U2758 ( .A(n5171), .B(n4783), .Y(n3542) );
  OAI21X1 U2759 ( .A(n4748), .B(n4603), .C(n5172), .Y(n5171) );
  OAI22X1 U2760 ( .A(n4662), .B(n5173), .C(n4582), .D(n5173), .Y(n5172) );
  OAI22X1 U2761 ( .A(n4668), .B(n4585), .C(n4673), .D(n4583), .Y(n5173) );
  XNOR2X1 U2762 ( .A(n5174), .B(n4783), .Y(n3541) );
  OAI21X1 U2763 ( .A(n4746), .B(n4603), .C(n5175), .Y(n5174) );
  OAI22X1 U2764 ( .A(n4666), .B(n5176), .C(n4582), .D(n5176), .Y(n5175) );
  OAI22X1 U2765 ( .A(n4673), .B(n4585), .C(n4678), .D(n4583), .Y(n5176) );
  XNOR2X1 U2766 ( .A(n5177), .B(n4783), .Y(n3540) );
  OAI21X1 U2767 ( .A(n4745), .B(n4603), .C(n5178), .Y(n5177) );
  OAI22X1 U2768 ( .A(n4671), .B(n5179), .C(n4582), .D(n5179), .Y(n5178) );
  OAI22X1 U2769 ( .A(n4678), .B(n4585), .C(n4683), .D(n4583), .Y(n5179) );
  XNOR2X1 U2770 ( .A(n5180), .B(n4783), .Y(n3539) );
  OAI21X1 U2771 ( .A(n4744), .B(n4603), .C(n5181), .Y(n5180) );
  OAI22X1 U2772 ( .A(n4676), .B(n5182), .C(n4582), .D(n5182), .Y(n5181) );
  OAI22X1 U2773 ( .A(n4683), .B(n4585), .C(n4688), .D(n4583), .Y(n5182) );
  XNOR2X1 U2774 ( .A(n5183), .B(n4783), .Y(n3538) );
  OAI21X1 U2775 ( .A(n4743), .B(n4603), .C(n5184), .Y(n5183) );
  OAI22X1 U2776 ( .A(n4681), .B(n5185), .C(n4582), .D(n5185), .Y(n5184) );
  OAI22X1 U2777 ( .A(n4688), .B(n4585), .C(n4693), .D(n4583), .Y(n5185) );
  XNOR2X1 U2778 ( .A(n5186), .B(n4783), .Y(n3537) );
  OAI21X1 U2779 ( .A(n4742), .B(n4603), .C(n5187), .Y(n5186) );
  OAI22X1 U2780 ( .A(n4686), .B(n5188), .C(n4582), .D(n5188), .Y(n5187) );
  OAI22X1 U2781 ( .A(n4693), .B(n4585), .C(n4697), .D(n4583), .Y(n5188) );
  XNOR2X1 U2782 ( .A(n5189), .B(n4584), .Y(n3536) );
  OAI21X1 U2783 ( .A(n4741), .B(n4603), .C(n5190), .Y(n5189) );
  OAI22X1 U2784 ( .A(n4691), .B(n5191), .C(n4582), .D(n5191), .Y(n5190) );
  OAI22X1 U2785 ( .A(n4697), .B(n4585), .C(n4701), .D(n4583), .Y(n5191) );
  XNOR2X1 U2786 ( .A(n5192), .B(n4584), .Y(n3535) );
  OAI21X1 U2787 ( .A(n4740), .B(n4603), .C(n5193), .Y(n5192) );
  OAI22X1 U2788 ( .A(n4696), .B(n5194), .C(n4582), .D(n5194), .Y(n5193) );
  OAI22X1 U2789 ( .A(n4701), .B(n4585), .C(n4705), .D(n4583), .Y(n5194) );
  XNOR2X1 U2790 ( .A(n5195), .B(n4584), .Y(n3534) );
  OAI21X1 U2791 ( .A(n4739), .B(n4603), .C(n5196), .Y(n5195) );
  OAI22X1 U2792 ( .A(n4700), .B(n5197), .C(n4582), .D(n5197), .Y(n5196) );
  OAI22X1 U2793 ( .A(n4705), .B(n4585), .C(n4709), .D(n4583), .Y(n5197) );
  XNOR2X1 U2794 ( .A(n5198), .B(n4584), .Y(n3533) );
  OAI21X1 U2795 ( .A(n4738), .B(n4603), .C(n5199), .Y(n5198) );
  OAI22X1 U2796 ( .A(n4704), .B(n5200), .C(n4582), .D(n5200), .Y(n5199) );
  OAI22X1 U2797 ( .A(n4709), .B(n4585), .C(n4712), .D(n4583), .Y(n5200) );
  XNOR2X1 U2798 ( .A(n5201), .B(n4584), .Y(n3532) );
  OAI21X1 U2799 ( .A(n4737), .B(n4603), .C(n5202), .Y(n5201) );
  OAI22X1 U2800 ( .A(n4708), .B(n5203), .C(n4582), .D(n5203), .Y(n5202) );
  OAI22X1 U2801 ( .A(n4712), .B(n4585), .C(n4568), .D(n4583), .Y(n5203) );
  XNOR2X1 U2802 ( .A(n5204), .B(n4584), .Y(n3531) );
  OAI21X1 U2803 ( .A(n4736), .B(n4603), .C(n5205), .Y(n5204) );
  OAI22X1 U2804 ( .A(n4711), .B(n5206), .C(n4582), .D(n5206), .Y(n5205) );
  OAI22X1 U2805 ( .A(n4568), .B(n4585), .C(n4735), .D(n4583), .Y(n5206) );
  XNOR2X1 U2806 ( .A(n5207), .B(n4584), .Y(n3530) );
  OAI21X1 U2807 ( .A(n4734), .B(n4603), .C(n5208), .Y(n5207) );
  OAI22X1 U2808 ( .A(n4569), .B(n5209), .C(n4582), .D(n5209), .Y(n5208) );
  OAI22X1 U2809 ( .A(n4735), .B(n4585), .C(n4733), .D(n4583), .Y(n5209) );
  XNOR2X1 U2810 ( .A(n5210), .B(n4584), .Y(n3529) );
  OAI21X1 U2811 ( .A(n4732), .B(n4603), .C(n5211), .Y(n5210) );
  OAI22X1 U2812 ( .A(b[25]), .B(n5212), .C(n4582), .D(n5212), .Y(n5211) );
  OAI22X1 U2813 ( .A(n4733), .B(n4585), .C(n4731), .D(n4583), .Y(n5212) );
  XNOR2X1 U2814 ( .A(n5213), .B(n4584), .Y(n3528) );
  OAI21X1 U2815 ( .A(n4730), .B(n4603), .C(n5214), .Y(n5213) );
  OAI22X1 U2816 ( .A(b[26]), .B(n5215), .C(n4582), .D(n5215), .Y(n5214) );
  OAI22X1 U2817 ( .A(n4731), .B(n4585), .C(n4729), .D(n4583), .Y(n5215) );
  XNOR2X1 U2818 ( .A(n5216), .B(n4584), .Y(n3527) );
  OAI21X1 U2819 ( .A(n4728), .B(n4603), .C(n5217), .Y(n5216) );
  OAI22X1 U2820 ( .A(b[27]), .B(n5218), .C(n4582), .D(n5218), .Y(n5217) );
  OAI22X1 U2821 ( .A(n4729), .B(n4585), .C(n4727), .D(n4583), .Y(n5218) );
  XNOR2X1 U2822 ( .A(n5219), .B(n4584), .Y(n3526) );
  OAI21X1 U2823 ( .A(n4726), .B(n4603), .C(n5220), .Y(n5219) );
  OAI22X1 U2824 ( .A(b[28]), .B(n5221), .C(n4582), .D(n5221), .Y(n5220) );
  OAI22X1 U2825 ( .A(n4727), .B(n4585), .C(n4725), .D(n4583), .Y(n5221) );
  XNOR2X1 U2826 ( .A(n5222), .B(n4584), .Y(n3525) );
  OAI21X1 U2827 ( .A(n4724), .B(n4603), .C(n5223), .Y(n5222) );
  OAI22X1 U2828 ( .A(b[29]), .B(n5224), .C(n4582), .D(n5224), .Y(n5223) );
  OAI22X1 U2829 ( .A(n4725), .B(n4585), .C(n4721), .D(n4583), .Y(n5224) );
  NOR2X1 U2830 ( .A(n5225), .B(n5226), .Y(n5134) );
  XNOR2X1 U2831 ( .A(n5227), .B(n4584), .Y(n3524) );
  OAI21X1 U2832 ( .A(n4723), .B(n4603), .C(n5228), .Y(n5227) );
  OAI22X1 U2833 ( .A(b[30]), .B(n5229), .C(n4582), .D(n5229), .Y(n5228) );
  NOR2X1 U2834 ( .A(n4585), .B(n4721), .Y(n5229) );
  NOR2X1 U2835 ( .A(n4784), .B(n5231), .Y(n5133) );
  XNOR2X1 U2836 ( .A(n5232), .B(n4584), .Y(n3523) );
  OAI22X1 U2837 ( .A(n4721), .B(n5230), .C(n4722), .D(n4603), .Y(n5232) );
  NAND3X1 U2838 ( .A(n5226), .B(n5225), .C(n5231), .Y(n5230) );
  XNOR2X1 U2839 ( .A(a[10]), .B(a[9]), .Y(n5231) );
  XNOR2X1 U2840 ( .A(a[10]), .B(n4584), .Y(n5225) );
  XOR2X1 U2841 ( .A(a[9]), .B(n4588), .Y(n5226) );
  XNOR2X1 U2842 ( .A(n5233), .B(n4580), .Y(n3521) );
  OAI22X1 U2843 ( .A(n4609), .B(n4579), .C(n4609), .D(n4604), .Y(n5233) );
  XNOR2X1 U2844 ( .A(n5234), .B(n4781), .Y(n3520) );
  OAI21X1 U2845 ( .A(n4765), .B(n4604), .C(n5235), .Y(n5234) );
  AOI22X1 U2846 ( .A(n5236), .B(n4607), .C(n5237), .D(n4610), .Y(n5235) );
  XNOR2X1 U2847 ( .A(n5238), .B(n4781), .Y(n3519) );
  OAI21X1 U2848 ( .A(n4762), .B(n4604), .C(n5239), .Y(n5238) );
  OAI22X1 U2849 ( .A(n4608), .B(n5240), .C(n4578), .D(n5240), .Y(n5239) );
  OAI22X1 U2850 ( .A(n4611), .B(n4581), .C(n4616), .D(n4579), .Y(n5240) );
  XNOR2X1 U2851 ( .A(n5241), .B(n4781), .Y(n3518) );
  OAI21X1 U2852 ( .A(n4761), .B(n4604), .C(n5242), .Y(n5241) );
  OAI22X1 U2853 ( .A(n4610), .B(n5243), .C(n4578), .D(n5243), .Y(n5242) );
  OAI22X1 U2854 ( .A(n4616), .B(n4581), .C(n4621), .D(n4579), .Y(n5243) );
  XNOR2X1 U2855 ( .A(n5244), .B(n4781), .Y(n3517) );
  OAI21X1 U2856 ( .A(n4760), .B(n4604), .C(n5245), .Y(n5244) );
  OAI22X1 U2857 ( .A(n4614), .B(n5246), .C(n4578), .D(n5246), .Y(n5245) );
  OAI22X1 U2858 ( .A(n4621), .B(n4581), .C(n4626), .D(n4579), .Y(n5246) );
  XNOR2X1 U2859 ( .A(n5247), .B(n4781), .Y(n3516) );
  OAI21X1 U2860 ( .A(n4759), .B(n4604), .C(n5248), .Y(n5247) );
  OAI22X1 U2861 ( .A(n4619), .B(n5249), .C(n4578), .D(n5249), .Y(n5248) );
  OAI22X1 U2862 ( .A(n4626), .B(n4581), .C(n4630), .D(n4579), .Y(n5249) );
  XNOR2X1 U2863 ( .A(n5250), .B(n4781), .Y(n3515) );
  OAI21X1 U2864 ( .A(n4758), .B(n4604), .C(n5251), .Y(n5250) );
  OAI22X1 U2865 ( .A(n4624), .B(n5252), .C(n4578), .D(n5252), .Y(n5251) );
  OAI22X1 U2866 ( .A(n4630), .B(n4581), .C(n4635), .D(n4579), .Y(n5252) );
  XNOR2X1 U2867 ( .A(n5253), .B(n4781), .Y(n3514) );
  OAI21X1 U2868 ( .A(n4757), .B(n4604), .C(n5254), .Y(n5253) );
  OAI22X1 U2869 ( .A(n4628), .B(n5255), .C(n4578), .D(n5255), .Y(n5254) );
  OAI22X1 U2870 ( .A(n4635), .B(n4581), .C(n4640), .D(n4579), .Y(n5255) );
  XNOR2X1 U2871 ( .A(n5256), .B(n4781), .Y(n3513) );
  OAI21X1 U2872 ( .A(n4755), .B(n4604), .C(n5257), .Y(n5256) );
  OAI22X1 U2873 ( .A(n4633), .B(n5258), .C(n4578), .D(n5258), .Y(n5257) );
  OAI22X1 U2874 ( .A(n4640), .B(n4581), .C(n4645), .D(n4579), .Y(n5258) );
  XNOR2X1 U2875 ( .A(n5259), .B(n4781), .Y(n3512) );
  OAI21X1 U2876 ( .A(n4754), .B(n4604), .C(n5260), .Y(n5259) );
  OAI22X1 U2877 ( .A(n4638), .B(n5261), .C(n4578), .D(n5261), .Y(n5260) );
  OAI22X1 U2878 ( .A(n4645), .B(n4581), .C(n4649), .D(n4579), .Y(n5261) );
  XNOR2X1 U2879 ( .A(n5262), .B(n4781), .Y(n3511) );
  OAI21X1 U2880 ( .A(n4753), .B(n4604), .C(n5263), .Y(n5262) );
  OAI22X1 U2881 ( .A(n4643), .B(n5264), .C(n4578), .D(n5264), .Y(n5263) );
  OAI22X1 U2882 ( .A(n4649), .B(n4581), .C(n4654), .D(n4579), .Y(n5264) );
  XNOR2X1 U2883 ( .A(n5265), .B(n4781), .Y(n3510) );
  OAI21X1 U2884 ( .A(n4751), .B(n4604), .C(n5266), .Y(n5265) );
  OAI22X1 U2885 ( .A(n4647), .B(n5267), .C(n4578), .D(n5267), .Y(n5266) );
  OAI22X1 U2886 ( .A(n4654), .B(n4581), .C(n4659), .D(n4579), .Y(n5267) );
  XNOR2X1 U2887 ( .A(n5268), .B(n4781), .Y(n3509) );
  OAI21X1 U2888 ( .A(n4750), .B(n4604), .C(n5269), .Y(n5268) );
  OAI22X1 U2889 ( .A(n4652), .B(n5270), .C(n4578), .D(n5270), .Y(n5269) );
  OAI22X1 U2890 ( .A(n4659), .B(n4581), .C(n4664), .D(n4579), .Y(n5270) );
  XNOR2X1 U2891 ( .A(n5271), .B(n4781), .Y(n3508) );
  OAI21X1 U2892 ( .A(n4749), .B(n4604), .C(n5272), .Y(n5271) );
  OAI22X1 U2893 ( .A(n4657), .B(n5273), .C(n4578), .D(n5273), .Y(n5272) );
  OAI22X1 U2894 ( .A(n4664), .B(n4581), .C(n4668), .D(n4579), .Y(n5273) );
  XNOR2X1 U2895 ( .A(n5274), .B(n4781), .Y(n3507) );
  OAI21X1 U2896 ( .A(n4748), .B(n4604), .C(n5275), .Y(n5274) );
  OAI22X1 U2897 ( .A(n4662), .B(n5276), .C(n4578), .D(n5276), .Y(n5275) );
  OAI22X1 U2898 ( .A(n4668), .B(n4581), .C(n4673), .D(n4579), .Y(n5276) );
  XNOR2X1 U2899 ( .A(n5277), .B(n4781), .Y(n3506) );
  OAI21X1 U2900 ( .A(n4746), .B(n4604), .C(n5278), .Y(n5277) );
  OAI22X1 U2901 ( .A(n4666), .B(n5279), .C(n4578), .D(n5279), .Y(n5278) );
  OAI22X1 U2902 ( .A(n4673), .B(n4581), .C(n4678), .D(n4579), .Y(n5279) );
  XNOR2X1 U2903 ( .A(n5280), .B(n4781), .Y(n3505) );
  OAI21X1 U2904 ( .A(n4745), .B(n4604), .C(n5281), .Y(n5280) );
  OAI22X1 U2905 ( .A(n4671), .B(n5282), .C(n4578), .D(n5282), .Y(n5281) );
  OAI22X1 U2906 ( .A(n4678), .B(n4581), .C(n4683), .D(n4579), .Y(n5282) );
  XNOR2X1 U2907 ( .A(n5283), .B(n4781), .Y(n3504) );
  OAI21X1 U2908 ( .A(n4744), .B(n4604), .C(n5284), .Y(n5283) );
  OAI22X1 U2909 ( .A(n4676), .B(n5285), .C(n4578), .D(n5285), .Y(n5284) );
  OAI22X1 U2910 ( .A(n4683), .B(n4581), .C(n4688), .D(n4579), .Y(n5285) );
  XNOR2X1 U2911 ( .A(n5286), .B(n4781), .Y(n3503) );
  OAI21X1 U2912 ( .A(n4743), .B(n4604), .C(n5287), .Y(n5286) );
  OAI22X1 U2913 ( .A(n4681), .B(n5288), .C(n4578), .D(n5288), .Y(n5287) );
  OAI22X1 U2914 ( .A(n4688), .B(n4581), .C(n4693), .D(n4579), .Y(n5288) );
  XNOR2X1 U2915 ( .A(n5289), .B(n4781), .Y(n3502) );
  OAI21X1 U2916 ( .A(n4742), .B(n4604), .C(n5290), .Y(n5289) );
  OAI22X1 U2917 ( .A(n4686), .B(n5291), .C(n4578), .D(n5291), .Y(n5290) );
  OAI22X1 U2918 ( .A(n4693), .B(n4581), .C(n4697), .D(n4579), .Y(n5291) );
  XNOR2X1 U2919 ( .A(n5292), .B(n4580), .Y(n3501) );
  OAI21X1 U2920 ( .A(n4741), .B(n4604), .C(n5293), .Y(n5292) );
  OAI22X1 U2921 ( .A(n4691), .B(n5294), .C(n4578), .D(n5294), .Y(n5293) );
  OAI22X1 U2922 ( .A(n4697), .B(n4581), .C(n4701), .D(n4579), .Y(n5294) );
  XNOR2X1 U2923 ( .A(n5295), .B(n4580), .Y(n3500) );
  OAI21X1 U2924 ( .A(n4740), .B(n4604), .C(n5296), .Y(n5295) );
  OAI22X1 U2925 ( .A(n4696), .B(n5297), .C(n4578), .D(n5297), .Y(n5296) );
  OAI22X1 U2926 ( .A(n4701), .B(n4581), .C(n4705), .D(n4579), .Y(n5297) );
  XNOR2X1 U2927 ( .A(n5298), .B(n4580), .Y(n3499) );
  OAI21X1 U2928 ( .A(n4739), .B(n4604), .C(n5299), .Y(n5298) );
  OAI22X1 U2929 ( .A(n4700), .B(n5300), .C(n4578), .D(n5300), .Y(n5299) );
  OAI22X1 U2930 ( .A(n4705), .B(n4581), .C(n4709), .D(n4579), .Y(n5300) );
  XNOR2X1 U2931 ( .A(n5301), .B(n4580), .Y(n3498) );
  OAI21X1 U2932 ( .A(n4738), .B(n4604), .C(n5302), .Y(n5301) );
  OAI22X1 U2933 ( .A(n4704), .B(n5303), .C(n4578), .D(n5303), .Y(n5302) );
  OAI22X1 U2934 ( .A(n4709), .B(n4581), .C(n4712), .D(n4579), .Y(n5303) );
  XNOR2X1 U2935 ( .A(n5304), .B(n4580), .Y(n3497) );
  OAI21X1 U2936 ( .A(n4737), .B(n4604), .C(n5305), .Y(n5304) );
  OAI22X1 U2937 ( .A(n4708), .B(n5306), .C(n4578), .D(n5306), .Y(n5305) );
  OAI22X1 U2938 ( .A(n4712), .B(n4581), .C(n4568), .D(n4579), .Y(n5306) );
  XNOR2X1 U2939 ( .A(n5307), .B(n4580), .Y(n3496) );
  OAI21X1 U2940 ( .A(n4736), .B(n4604), .C(n5308), .Y(n5307) );
  OAI22X1 U2941 ( .A(n4711), .B(n5309), .C(n4578), .D(n5309), .Y(n5308) );
  OAI22X1 U2942 ( .A(n4568), .B(n4581), .C(n4735), .D(n4579), .Y(n5309) );
  XNOR2X1 U2943 ( .A(n5310), .B(n4580), .Y(n3495) );
  OAI21X1 U2944 ( .A(n4734), .B(n4604), .C(n5311), .Y(n5310) );
  OAI22X1 U2945 ( .A(n4569), .B(n5312), .C(n4578), .D(n5312), .Y(n5311) );
  OAI22X1 U2946 ( .A(n4735), .B(n4581), .C(n4733), .D(n4579), .Y(n5312) );
  XNOR2X1 U2947 ( .A(n5313), .B(n4580), .Y(n3494) );
  OAI21X1 U2948 ( .A(n4732), .B(n4604), .C(n5314), .Y(n5313) );
  OAI22X1 U2949 ( .A(b[25]), .B(n5315), .C(n4578), .D(n5315), .Y(n5314) );
  OAI22X1 U2950 ( .A(n4733), .B(n4581), .C(n4731), .D(n4579), .Y(n5315) );
  XNOR2X1 U2951 ( .A(n5316), .B(n4580), .Y(n3493) );
  OAI21X1 U2952 ( .A(n4730), .B(n4604), .C(n5317), .Y(n5316) );
  OAI22X1 U2953 ( .A(b[26]), .B(n5318), .C(n4578), .D(n5318), .Y(n5317) );
  OAI22X1 U2954 ( .A(n4731), .B(n4581), .C(n4729), .D(n4579), .Y(n5318) );
  XNOR2X1 U2955 ( .A(n5319), .B(n4580), .Y(n3492) );
  OAI21X1 U2956 ( .A(n4728), .B(n4604), .C(n5320), .Y(n5319) );
  OAI22X1 U2957 ( .A(b[27]), .B(n5321), .C(n4578), .D(n5321), .Y(n5320) );
  OAI22X1 U2958 ( .A(n4729), .B(n4581), .C(n4727), .D(n4579), .Y(n5321) );
  XNOR2X1 U2959 ( .A(n5322), .B(n4580), .Y(n3491) );
  OAI21X1 U2960 ( .A(n4726), .B(n4604), .C(n5323), .Y(n5322) );
  OAI22X1 U2961 ( .A(b[28]), .B(n5324), .C(n4578), .D(n5324), .Y(n5323) );
  OAI22X1 U2962 ( .A(n4727), .B(n4581), .C(n4725), .D(n4579), .Y(n5324) );
  XNOR2X1 U2963 ( .A(n5325), .B(n4580), .Y(n3490) );
  OAI21X1 U2964 ( .A(n4724), .B(n4604), .C(n5326), .Y(n5325) );
  OAI22X1 U2965 ( .A(b[29]), .B(n5327), .C(n4578), .D(n5327), .Y(n5326) );
  OAI22X1 U2966 ( .A(n4725), .B(n4581), .C(n4721), .D(n4579), .Y(n5327) );
  NOR2X1 U2967 ( .A(n5328), .B(n5329), .Y(n5237) );
  XNOR2X1 U2968 ( .A(n5330), .B(n4580), .Y(n3489) );
  OAI21X1 U2969 ( .A(n4723), .B(n4604), .C(n5331), .Y(n5330) );
  OAI22X1 U2970 ( .A(b[30]), .B(n5332), .C(n4578), .D(n5332), .Y(n5331) );
  NOR2X1 U2971 ( .A(n4581), .B(n4721), .Y(n5332) );
  NOR2X1 U2972 ( .A(n4782), .B(n5334), .Y(n5236) );
  XNOR2X1 U2973 ( .A(n5335), .B(n4580), .Y(n3488) );
  OAI22X1 U2974 ( .A(n4721), .B(n5333), .C(n4722), .D(n4604), .Y(n5335) );
  NAND3X1 U2975 ( .A(n5329), .B(n5328), .C(n5334), .Y(n5333) );
  XNOR2X1 U2976 ( .A(a[12]), .B(a[13]), .Y(n5334) );
  XNOR2X1 U2977 ( .A(a[13]), .B(n4580), .Y(n5328) );
  XOR2X1 U2978 ( .A(a[12]), .B(n4584), .Y(n5329) );
  XNOR2X1 U2979 ( .A(n5336), .B(n4577), .Y(n3486) );
  OAI22X1 U2980 ( .A(n4609), .B(n4552), .C(n4597), .D(n4609), .Y(n5336) );
  XNOR2X1 U2981 ( .A(n5337), .B(n4779), .Y(n3485) );
  OAI21X1 U2982 ( .A(n4597), .B(n4765), .C(n4763), .Y(n5337) );
  OAI22X1 U2983 ( .A(n4609), .B(n4554), .C(n4552), .D(n4611), .Y(n5338) );
  XNOR2X1 U2984 ( .A(n5339), .B(n4779), .Y(n3484) );
  OAI21X1 U2985 ( .A(n4597), .B(n4762), .C(n5340), .Y(n5339) );
  OAI22X1 U2986 ( .A(n4608), .B(n5341), .C(n4576), .D(n5341), .Y(n5340) );
  OAI22X1 U2987 ( .A(n4616), .B(n4552), .C(n4554), .D(n4611), .Y(n5341) );
  XNOR2X1 U2988 ( .A(n5342), .B(n4779), .Y(n3483) );
  OAI21X1 U2989 ( .A(n4597), .B(n4761), .C(n5343), .Y(n5342) );
  OAI22X1 U2990 ( .A(n4610), .B(n5344), .C(n4576), .D(n5344), .Y(n5343) );
  OAI22X1 U2991 ( .A(n4621), .B(n4552), .C(n4554), .D(n4616), .Y(n5344) );
  XNOR2X1 U2992 ( .A(n5345), .B(n4779), .Y(n3482) );
  OAI21X1 U2993 ( .A(n4597), .B(n4760), .C(n5346), .Y(n5345) );
  OAI22X1 U2994 ( .A(n4614), .B(n5347), .C(n4576), .D(n5347), .Y(n5346) );
  OAI22X1 U2995 ( .A(n4626), .B(n4552), .C(n4554), .D(n4621), .Y(n5347) );
  XNOR2X1 U2996 ( .A(n5348), .B(n4779), .Y(n3481) );
  OAI21X1 U2997 ( .A(n4597), .B(n4759), .C(n5349), .Y(n5348) );
  OAI22X1 U2998 ( .A(n4619), .B(n5350), .C(n4576), .D(n5350), .Y(n5349) );
  OAI22X1 U2999 ( .A(n4630), .B(n4552), .C(n4554), .D(n4626), .Y(n5350) );
  XNOR2X1 U3000 ( .A(n5351), .B(n4779), .Y(n3480) );
  OAI21X1 U3001 ( .A(n4597), .B(n4758), .C(n5352), .Y(n5351) );
  OAI22X1 U3002 ( .A(n4624), .B(n5353), .C(n4576), .D(n5353), .Y(n5352) );
  OAI22X1 U3003 ( .A(n4635), .B(n4552), .C(n4554), .D(n4630), .Y(n5353) );
  XNOR2X1 U3004 ( .A(n5354), .B(n4779), .Y(n3479) );
  OAI21X1 U3005 ( .A(n4597), .B(n4757), .C(n5355), .Y(n5354) );
  OAI22X1 U3006 ( .A(n4628), .B(n5356), .C(n4576), .D(n5356), .Y(n5355) );
  OAI22X1 U3007 ( .A(n4640), .B(n4552), .C(n4554), .D(n4635), .Y(n5356) );
  XNOR2X1 U3008 ( .A(n5357), .B(n4779), .Y(n3478) );
  OAI21X1 U3009 ( .A(n4597), .B(n4755), .C(n5358), .Y(n5357) );
  OAI22X1 U3010 ( .A(n4633), .B(n5359), .C(n4576), .D(n5359), .Y(n5358) );
  OAI22X1 U3011 ( .A(n4645), .B(n4552), .C(n4554), .D(n4640), .Y(n5359) );
  XNOR2X1 U3012 ( .A(n5360), .B(n4779), .Y(n3477) );
  OAI21X1 U3013 ( .A(n4597), .B(n4754), .C(n5361), .Y(n5360) );
  OAI22X1 U3014 ( .A(n4638), .B(n5362), .C(n4576), .D(n5362), .Y(n5361) );
  OAI22X1 U3015 ( .A(n4649), .B(n4552), .C(n4554), .D(n4645), .Y(n5362) );
  XNOR2X1 U3016 ( .A(n5363), .B(n4779), .Y(n3476) );
  OAI21X1 U3017 ( .A(n4597), .B(n4753), .C(n5364), .Y(n5363) );
  OAI22X1 U3018 ( .A(n4643), .B(n5365), .C(n4576), .D(n5365), .Y(n5364) );
  OAI22X1 U3019 ( .A(n4654), .B(n4552), .C(n4554), .D(n4649), .Y(n5365) );
  XNOR2X1 U3020 ( .A(n5366), .B(n4779), .Y(n3475) );
  OAI21X1 U3021 ( .A(n4597), .B(n4751), .C(n5367), .Y(n5366) );
  OAI22X1 U3022 ( .A(n4647), .B(n5368), .C(n4576), .D(n5368), .Y(n5367) );
  OAI22X1 U3023 ( .A(n4659), .B(n4552), .C(n4554), .D(n4654), .Y(n5368) );
  XNOR2X1 U3024 ( .A(n5369), .B(n4779), .Y(n3474) );
  OAI21X1 U3025 ( .A(n4597), .B(n4750), .C(n5370), .Y(n5369) );
  OAI22X1 U3026 ( .A(n4652), .B(n5371), .C(n4576), .D(n5371), .Y(n5370) );
  OAI22X1 U3027 ( .A(n4664), .B(n4552), .C(n4554), .D(n4659), .Y(n5371) );
  XNOR2X1 U3028 ( .A(n5372), .B(n4779), .Y(n3473) );
  OAI21X1 U3029 ( .A(n4597), .B(n4749), .C(n5373), .Y(n5372) );
  OAI22X1 U3030 ( .A(n4657), .B(n5374), .C(n4576), .D(n5374), .Y(n5373) );
  OAI22X1 U3031 ( .A(n4668), .B(n4552), .C(n4554), .D(n4664), .Y(n5374) );
  XNOR2X1 U3032 ( .A(n5375), .B(n4779), .Y(n3472) );
  OAI21X1 U3033 ( .A(n4597), .B(n4748), .C(n5376), .Y(n5375) );
  OAI22X1 U3034 ( .A(n4662), .B(n5377), .C(n4576), .D(n5377), .Y(n5376) );
  OAI22X1 U3035 ( .A(n4673), .B(n4552), .C(n4554), .D(n4668), .Y(n5377) );
  XNOR2X1 U3036 ( .A(n5378), .B(n4779), .Y(n3471) );
  OAI21X1 U3037 ( .A(n4597), .B(n4746), .C(n5379), .Y(n5378) );
  OAI22X1 U3038 ( .A(n4666), .B(n5380), .C(n4576), .D(n5380), .Y(n5379) );
  OAI22X1 U3039 ( .A(n4678), .B(n4552), .C(n4554), .D(n4673), .Y(n5380) );
  XNOR2X1 U3040 ( .A(n5381), .B(n4779), .Y(n3470) );
  OAI21X1 U3041 ( .A(n4597), .B(n4745), .C(n5382), .Y(n5381) );
  OAI22X1 U3042 ( .A(n4671), .B(n5383), .C(n4576), .D(n5383), .Y(n5382) );
  OAI22X1 U3043 ( .A(n4683), .B(n4552), .C(n4554), .D(n4678), .Y(n5383) );
  XNOR2X1 U3044 ( .A(n5384), .B(n4779), .Y(n3469) );
  OAI21X1 U3045 ( .A(n4744), .B(n4597), .C(n5385), .Y(n5384) );
  OAI22X1 U3046 ( .A(n4676), .B(n5386), .C(n4576), .D(n5386), .Y(n5385) );
  OAI22X1 U3047 ( .A(n4688), .B(n4552), .C(n4683), .D(n4554), .Y(n5386) );
  XNOR2X1 U3048 ( .A(n5387), .B(n4779), .Y(n3468) );
  OAI21X1 U3049 ( .A(n4597), .B(n4743), .C(n5388), .Y(n5387) );
  OAI22X1 U3050 ( .A(n4681), .B(n5389), .C(n4576), .D(n5389), .Y(n5388) );
  OAI22X1 U3051 ( .A(n4693), .B(n4552), .C(n4688), .D(n4554), .Y(n5389) );
  XNOR2X1 U3052 ( .A(n5390), .B(n4779), .Y(n3467) );
  OAI21X1 U3053 ( .A(n4597), .B(n4742), .C(n5391), .Y(n5390) );
  OAI22X1 U3054 ( .A(n4686), .B(n5392), .C(n4576), .D(n5392), .Y(n5391) );
  OAI22X1 U3055 ( .A(n4697), .B(n4552), .C(n4554), .D(n4693), .Y(n5392) );
  XNOR2X1 U3056 ( .A(n5393), .B(n4779), .Y(n3466) );
  OAI21X1 U3057 ( .A(n4741), .B(n4597), .C(n5394), .Y(n5393) );
  OAI22X1 U3058 ( .A(n4691), .B(n5395), .C(n4576), .D(n5395), .Y(n5394) );
  OAI22X1 U3059 ( .A(n4701), .B(n4552), .C(n4697), .D(n4554), .Y(n5395) );
  XNOR2X1 U3060 ( .A(n5396), .B(n4779), .Y(n3465) );
  OAI21X1 U3061 ( .A(n4597), .B(n4740), .C(n5397), .Y(n5396) );
  OAI22X1 U3062 ( .A(n4696), .B(n5398), .C(n4576), .D(n5398), .Y(n5397) );
  OAI22X1 U3063 ( .A(n4705), .B(n4552), .C(n4701), .D(n4554), .Y(n5398) );
  XNOR2X1 U3064 ( .A(n5399), .B(n4779), .Y(n3464) );
  OAI21X1 U3065 ( .A(n4597), .B(n4739), .C(n5400), .Y(n5399) );
  OAI22X1 U3066 ( .A(n4700), .B(n5401), .C(n4576), .D(n5401), .Y(n5400) );
  OAI22X1 U3067 ( .A(n4709), .B(n4552), .C(n4554), .D(n4705), .Y(n5401) );
  XNOR2X1 U3068 ( .A(n5402), .B(n4779), .Y(n3463) );
  OAI21X1 U3069 ( .A(n4738), .B(n4597), .C(n5403), .Y(n5402) );
  OAI22X1 U3070 ( .A(n4703), .B(n5404), .C(n4576), .D(n5404), .Y(n5403) );
  OAI22X1 U3071 ( .A(n4712), .B(n4552), .C(n4709), .D(n4554), .Y(n5404) );
  XNOR2X1 U3072 ( .A(n5405), .B(n4577), .Y(n3462) );
  OAI21X1 U3073 ( .A(n4597), .B(n4737), .C(n5406), .Y(n5405) );
  OAI22X1 U3074 ( .A(n4708), .B(n5407), .C(n4576), .D(n5407), .Y(n5406) );
  OAI22X1 U3075 ( .A(n4568), .B(n4552), .C(n4712), .D(n4554), .Y(n5407) );
  XNOR2X1 U3076 ( .A(n5408), .B(n4577), .Y(n3461) );
  OAI21X1 U3077 ( .A(n4597), .B(n4736), .C(n5409), .Y(n5408) );
  OAI22X1 U3078 ( .A(n4711), .B(n5410), .C(n4576), .D(n5410), .Y(n5409) );
  OAI22X1 U3079 ( .A(n4735), .B(n4552), .C(n4554), .D(n4568), .Y(n5410) );
  XNOR2X1 U3080 ( .A(n5411), .B(n4577), .Y(n3460) );
  OAI21X1 U3081 ( .A(n4734), .B(n4597), .C(n5412), .Y(n5411) );
  OAI22X1 U3082 ( .A(n4569), .B(n5413), .C(n4576), .D(n5413), .Y(n5412) );
  OAI22X1 U3083 ( .A(n4733), .B(n4552), .C(n4735), .D(n4554), .Y(n5413) );
  XNOR2X1 U3084 ( .A(n5414), .B(n4577), .Y(n3459) );
  OAI21X1 U3085 ( .A(n4597), .B(n4732), .C(n5415), .Y(n5414) );
  OAI22X1 U3086 ( .A(b[25]), .B(n5416), .C(n4576), .D(n5416), .Y(n5415) );
  OAI22X1 U3087 ( .A(n4731), .B(n4552), .C(n4733), .D(n4554), .Y(n5416) );
  XNOR2X1 U3088 ( .A(n5417), .B(n4577), .Y(n3458) );
  OAI21X1 U3089 ( .A(n4597), .B(n4730), .C(n5418), .Y(n5417) );
  OAI22X1 U3090 ( .A(b[26]), .B(n5419), .C(n4576), .D(n5419), .Y(n5418) );
  OAI22X1 U3091 ( .A(n4729), .B(n4552), .C(n4554), .D(n4731), .Y(n5419) );
  XNOR2X1 U3092 ( .A(n5420), .B(n4577), .Y(n3457) );
  OAI21X1 U3093 ( .A(n4728), .B(n4597), .C(n5421), .Y(n5420) );
  OAI22X1 U3094 ( .A(b[27]), .B(n5422), .C(n4576), .D(n5422), .Y(n5421) );
  OAI22X1 U3095 ( .A(n4727), .B(n4552), .C(n4729), .D(n4554), .Y(n5422) );
  XNOR2X1 U3096 ( .A(n5423), .B(n4577), .Y(n3456) );
  OAI21X1 U3097 ( .A(n4597), .B(n4726), .C(n5424), .Y(n5423) );
  OAI22X1 U3098 ( .A(b[28]), .B(n5425), .C(n4576), .D(n5425), .Y(n5424) );
  OAI22X1 U3099 ( .A(n4727), .B(n4554), .C(n4725), .D(n4552), .Y(n5425) );
  XNOR2X1 U3100 ( .A(n5426), .B(n4577), .Y(n3455) );
  OAI21X1 U3101 ( .A(n4597), .B(n4724), .C(n5427), .Y(n5426) );
  OAI22X1 U3102 ( .A(b[29]), .B(n5428), .C(n4576), .D(n5428), .Y(n5427) );
  NAND3X1 U3103 ( .A(n5430), .B(n5431), .C(n5432), .Y(n5429) );
  OAI22X1 U3104 ( .A(n4554), .B(n4725), .C(n4721), .D(n4552), .Y(n5428) );
  XNOR2X1 U3105 ( .A(a[15]), .B(a[16]), .Y(n5430) );
  XNOR2X1 U3106 ( .A(a[16]), .B(n4577), .Y(n5431) );
  XOR2X1 U3107 ( .A(a[15]), .B(n4580), .Y(n5432) );
  XOR2X1 U3108 ( .A(n5433), .B(n4719), .Y(n3453) );
  OAI22X1 U3109 ( .A(n4573), .B(n4609), .C(n4598), .D(n4609), .Y(n5433) );
  XOR2X1 U3110 ( .A(n5434), .B(n4719), .Y(n3452) );
  OAI21X1 U3111 ( .A(n4598), .B(n4765), .C(n5435), .Y(n5434) );
  AOI22X1 U3112 ( .A(n4610), .B(n5436), .C(n4606), .D(n5437), .Y(n5435) );
  XOR2X1 U3113 ( .A(n5438), .B(n4719), .Y(n3451) );
  OAI21X1 U3114 ( .A(n4598), .B(n4762), .C(n5439), .Y(n5438) );
  OAI22X1 U3115 ( .A(n4608), .B(n5440), .C(n4574), .D(n5440), .Y(n5439) );
  OAI22X1 U3116 ( .A(n4575), .B(n4611), .C(n4573), .D(n4616), .Y(n5440) );
  XOR2X1 U3117 ( .A(n5441), .B(n4719), .Y(n3450) );
  OAI21X1 U3118 ( .A(n4598), .B(n4761), .C(n5442), .Y(n5441) );
  OAI22X1 U3119 ( .A(n4610), .B(n5443), .C(n4574), .D(n5443), .Y(n5442) );
  OAI22X1 U3120 ( .A(n4575), .B(n4616), .C(n4573), .D(n4621), .Y(n5443) );
  XOR2X1 U3121 ( .A(n5444), .B(n4719), .Y(n3449) );
  OAI21X1 U3122 ( .A(n4598), .B(n4760), .C(n5445), .Y(n5444) );
  OAI22X1 U3123 ( .A(n4614), .B(n5446), .C(n4574), .D(n5446), .Y(n5445) );
  OAI22X1 U3124 ( .A(n4575), .B(n4621), .C(n4573), .D(n4626), .Y(n5446) );
  XOR2X1 U3125 ( .A(n5447), .B(n4719), .Y(n3448) );
  OAI21X1 U3126 ( .A(n4598), .B(n4759), .C(n5448), .Y(n5447) );
  OAI22X1 U3127 ( .A(n4619), .B(n5449), .C(n4574), .D(n5449), .Y(n5448) );
  OAI22X1 U3128 ( .A(n4575), .B(n4626), .C(n4573), .D(n4630), .Y(n5449) );
  XOR2X1 U3129 ( .A(n5450), .B(n4719), .Y(n3447) );
  OAI21X1 U3130 ( .A(n4598), .B(n4758), .C(n5451), .Y(n5450) );
  OAI22X1 U3131 ( .A(n4624), .B(n5452), .C(n4574), .D(n5452), .Y(n5451) );
  OAI22X1 U3132 ( .A(n4575), .B(n4630), .C(n4573), .D(n4635), .Y(n5452) );
  XOR2X1 U3133 ( .A(n5453), .B(n4719), .Y(n3446) );
  OAI21X1 U3134 ( .A(n4598), .B(n4757), .C(n5454), .Y(n5453) );
  OAI22X1 U3135 ( .A(n4628), .B(n5455), .C(n4574), .D(n5455), .Y(n5454) );
  OAI22X1 U3136 ( .A(n4575), .B(n4635), .C(n4573), .D(n4640), .Y(n5455) );
  XOR2X1 U3137 ( .A(n5456), .B(n4719), .Y(n3445) );
  OAI21X1 U3138 ( .A(n4598), .B(n4755), .C(n5457), .Y(n5456) );
  OAI22X1 U3139 ( .A(n4633), .B(n5458), .C(n4574), .D(n5458), .Y(n5457) );
  OAI22X1 U3140 ( .A(n4575), .B(n4640), .C(n4573), .D(n4645), .Y(n5458) );
  XOR2X1 U3141 ( .A(n5459), .B(n4719), .Y(n3444) );
  OAI21X1 U3142 ( .A(n4598), .B(n4754), .C(n5460), .Y(n5459) );
  OAI22X1 U3143 ( .A(n4638), .B(n5461), .C(n4574), .D(n5461), .Y(n5460) );
  OAI22X1 U3144 ( .A(n4575), .B(n4645), .C(n4573), .D(n4649), .Y(n5461) );
  XOR2X1 U3145 ( .A(n5462), .B(n4719), .Y(n3443) );
  OAI21X1 U3146 ( .A(n4598), .B(n4753), .C(n5463), .Y(n5462) );
  OAI22X1 U3147 ( .A(n4643), .B(n5464), .C(n4574), .D(n5464), .Y(n5463) );
  OAI22X1 U3148 ( .A(n4575), .B(n4649), .C(n4573), .D(n4654), .Y(n5464) );
  XOR2X1 U3149 ( .A(n5465), .B(n4719), .Y(n3442) );
  OAI21X1 U3150 ( .A(n4598), .B(n4751), .C(n5466), .Y(n5465) );
  OAI22X1 U3151 ( .A(n4647), .B(n5467), .C(n4574), .D(n5467), .Y(n5466) );
  OAI22X1 U3152 ( .A(n4575), .B(n4654), .C(n4573), .D(n4659), .Y(n5467) );
  XOR2X1 U3153 ( .A(n5468), .B(n4719), .Y(n3441) );
  OAI21X1 U3154 ( .A(n4598), .B(n4750), .C(n5469), .Y(n5468) );
  OAI22X1 U3155 ( .A(n4652), .B(n5470), .C(n4574), .D(n5470), .Y(n5469) );
  OAI22X1 U3156 ( .A(n4575), .B(n4659), .C(n4573), .D(n4664), .Y(n5470) );
  XOR2X1 U3157 ( .A(n5471), .B(n4719), .Y(n3440) );
  OAI21X1 U3158 ( .A(n4598), .B(n4749), .C(n5472), .Y(n5471) );
  OAI22X1 U3159 ( .A(n4657), .B(n5473), .C(n4574), .D(n5473), .Y(n5472) );
  OAI22X1 U3160 ( .A(n4575), .B(n4664), .C(n4573), .D(n4668), .Y(n5473) );
  XOR2X1 U3161 ( .A(n5474), .B(n4719), .Y(n3439) );
  OAI21X1 U3162 ( .A(n4598), .B(n4748), .C(n5475), .Y(n5474) );
  OAI22X1 U3163 ( .A(n4662), .B(n5476), .C(n4574), .D(n5476), .Y(n5475) );
  OAI22X1 U3164 ( .A(n4575), .B(n4668), .C(n4573), .D(n4673), .Y(n5476) );
  XOR2X1 U3165 ( .A(n5477), .B(n4719), .Y(n3438) );
  OAI21X1 U3166 ( .A(n4598), .B(n4746), .C(n5478), .Y(n5477) );
  OAI22X1 U3167 ( .A(n4666), .B(n5479), .C(n4574), .D(n5479), .Y(n5478) );
  OAI22X1 U3168 ( .A(n4573), .B(n4678), .C(n4575), .D(n4673), .Y(n5479) );
  XOR2X1 U3169 ( .A(n5480), .B(n4719), .Y(n3437) );
  OAI21X1 U3170 ( .A(n4598), .B(n4745), .C(n5481), .Y(n5480) );
  OAI22X1 U3171 ( .A(n4671), .B(n5482), .C(n4574), .D(n5482), .Y(n5481) );
  OAI22X1 U3172 ( .A(n4575), .B(n4678), .C(n4573), .D(n4683), .Y(n5482) );
  XOR2X1 U3173 ( .A(n5483), .B(n4719), .Y(n3436) );
  OAI21X1 U3174 ( .A(n4598), .B(n4744), .C(n5484), .Y(n5483) );
  OAI22X1 U3175 ( .A(n4676), .B(n5485), .C(n4574), .D(n5485), .Y(n5484) );
  OAI22X1 U3176 ( .A(n4573), .B(n4688), .C(n4575), .D(n4683), .Y(n5485) );
  XOR2X1 U3177 ( .A(n5486), .B(n4719), .Y(n3435) );
  OAI21X1 U3178 ( .A(n4598), .B(n4743), .C(n5487), .Y(n5486) );
  OAI22X1 U3179 ( .A(n4681), .B(n5488), .C(n4574), .D(n5488), .Y(n5487) );
  OAI22X1 U3180 ( .A(n4575), .B(n4688), .C(n4573), .D(n4693), .Y(n5488) );
  XOR2X1 U3181 ( .A(n5489), .B(n4719), .Y(n3434) );
  OAI21X1 U3182 ( .A(n4598), .B(n4742), .C(n5490), .Y(n5489) );
  OAI22X1 U3183 ( .A(n4686), .B(n5491), .C(n4574), .D(n5491), .Y(n5490) );
  OAI22X1 U3184 ( .A(n4575), .B(n4693), .C(n4573), .D(n4697), .Y(n5491) );
  XOR2X1 U3185 ( .A(n5492), .B(n2150), .Y(n3433) );
  OAI21X1 U3186 ( .A(n4598), .B(n4741), .C(n5493), .Y(n5492) );
  OAI22X1 U3187 ( .A(n4691), .B(n5494), .C(n4574), .D(n5494), .Y(n5493) );
  OAI22X1 U3188 ( .A(n4573), .B(n4701), .C(n4575), .D(n4697), .Y(n5494) );
  XOR2X1 U3189 ( .A(n5495), .B(n2150), .Y(n3432) );
  OAI21X1 U3190 ( .A(n4598), .B(n4740), .C(n5496), .Y(n5495) );
  OAI22X1 U3191 ( .A(n4695), .B(n5497), .C(n4574), .D(n5497), .Y(n5496) );
  OAI22X1 U3192 ( .A(n4575), .B(n4701), .C(n4573), .D(n4705), .Y(n5497) );
  XOR2X1 U3193 ( .A(n5498), .B(n2150), .Y(n3431) );
  OAI21X1 U3194 ( .A(n4598), .B(n4739), .C(n5499), .Y(n5498) );
  OAI22X1 U3195 ( .A(n4699), .B(n5500), .C(n4574), .D(n5500), .Y(n5499) );
  OAI22X1 U3196 ( .A(n4575), .B(n4705), .C(n4573), .D(n4709), .Y(n5500) );
  XOR2X1 U3197 ( .A(n5501), .B(n2150), .Y(n3430) );
  OAI21X1 U3198 ( .A(n4598), .B(n4738), .C(n5502), .Y(n5501) );
  OAI22X1 U3199 ( .A(n4704), .B(n5503), .C(n4574), .D(n5503), .Y(n5502) );
  OAI22X1 U3200 ( .A(n4573), .B(n4712), .C(n4575), .D(n4709), .Y(n5503) );
  XOR2X1 U3201 ( .A(n5504), .B(n2150), .Y(n3429) );
  OAI21X1 U3202 ( .A(n4598), .B(n4737), .C(n5505), .Y(n5504) );
  OAI22X1 U3203 ( .A(n4708), .B(n5506), .C(n4574), .D(n5506), .Y(n5505) );
  OAI22X1 U3204 ( .A(n4575), .B(n4712), .C(n4573), .D(n4568), .Y(n5506) );
  XOR2X1 U3205 ( .A(n5507), .B(n2150), .Y(n3428) );
  OAI21X1 U3206 ( .A(n4598), .B(n4736), .C(n5508), .Y(n5507) );
  OAI22X1 U3207 ( .A(n4711), .B(n5509), .C(n4574), .D(n5509), .Y(n5508) );
  OAI22X1 U3208 ( .A(n4575), .B(n4568), .C(n4573), .D(n4735), .Y(n5509) );
  XOR2X1 U3209 ( .A(n5510), .B(n2150), .Y(n3427) );
  OAI21X1 U3210 ( .A(n4598), .B(n4734), .C(n5511), .Y(n5510) );
  OAI22X1 U3211 ( .A(n4569), .B(n5512), .C(n4574), .D(n5512), .Y(n5511) );
  OAI22X1 U3212 ( .A(n4573), .B(n4733), .C(n4575), .D(n4735), .Y(n5512) );
  XOR2X1 U3213 ( .A(n5513), .B(n2150), .Y(n3426) );
  OAI21X1 U3214 ( .A(n4598), .B(n4732), .C(n5514), .Y(n5513) );
  OAI22X1 U3215 ( .A(b[25]), .B(n5515), .C(n4574), .D(n5515), .Y(n5514) );
  OAI22X1 U3216 ( .A(n4575), .B(n4733), .C(n4573), .D(n4731), .Y(n5515) );
  XOR2X1 U3217 ( .A(n5516), .B(n2150), .Y(n3425) );
  OAI21X1 U3218 ( .A(n4598), .B(n4730), .C(n5517), .Y(n5516) );
  OAI22X1 U3219 ( .A(b[26]), .B(n5518), .C(n4574), .D(n5518), .Y(n5517) );
  NAND3X1 U3220 ( .A(n5520), .B(n5521), .C(n5522), .Y(n5519) );
  OAI22X1 U3221 ( .A(n4575), .B(n4731), .C(n4729), .D(n4573), .Y(n5518) );
  NOR2X1 U3222 ( .A(n5521), .B(n5520), .Y(n5436) );
  NOR2X1 U3223 ( .A(n4778), .B(n5522), .Y(n5437) );
  XNOR2X1 U3224 ( .A(a[18]), .B(a[19]), .Y(n5522) );
  XOR2X1 U3225 ( .A(a[19]), .B(n2150), .Y(n5521) );
  XOR2X1 U3226 ( .A(a[18]), .B(n4577), .Y(n5520) );
  XOR2X1 U3227 ( .A(n4717), .B(n5523), .Y(n3423) );
  OAI22X1 U3228 ( .A(n4609), .B(n4555), .C(n4609), .D(n4570), .Y(n5523) );
  XOR2X1 U3229 ( .A(n5524), .B(n2153), .Y(n3422) );
  OAI21X1 U3230 ( .A(n4555), .B(n4765), .C(n5525), .Y(n5524) );
  AOI22X1 U3231 ( .A(n4610), .B(n5526), .C(n4606), .D(n5527), .Y(n5525) );
  XOR2X1 U3232 ( .A(n5528), .B(n2153), .Y(n3421) );
  OAI21X1 U3233 ( .A(n4555), .B(n4762), .C(n5529), .Y(n5528) );
  OAI22X1 U3234 ( .A(n4608), .B(n5530), .C(n4571), .D(n5530), .Y(n5529) );
  OAI22X1 U3235 ( .A(n4572), .B(n4611), .C(n4570), .D(n4616), .Y(n5530) );
  XOR2X1 U3236 ( .A(n5531), .B(n2153), .Y(n3420) );
  OAI21X1 U3237 ( .A(n4555), .B(n4761), .C(n5532), .Y(n5531) );
  OAI22X1 U3238 ( .A(n4610), .B(n5533), .C(n4571), .D(n5533), .Y(n5532) );
  OAI22X1 U3239 ( .A(n4572), .B(n4616), .C(n4570), .D(n4621), .Y(n5533) );
  XOR2X1 U3240 ( .A(n5534), .B(n2153), .Y(n3419) );
  OAI21X1 U3241 ( .A(n4555), .B(n4760), .C(n5535), .Y(n5534) );
  OAI22X1 U3242 ( .A(n4614), .B(n5536), .C(n4571), .D(n5536), .Y(n5535) );
  OAI22X1 U3243 ( .A(n4572), .B(n4621), .C(n4570), .D(n4626), .Y(n5536) );
  XOR2X1 U3244 ( .A(n5537), .B(n2153), .Y(n3418) );
  OAI21X1 U3245 ( .A(n4555), .B(n4759), .C(n5538), .Y(n5537) );
  OAI22X1 U3246 ( .A(n4619), .B(n5539), .C(n4571), .D(n5539), .Y(n5538) );
  OAI22X1 U3247 ( .A(n4572), .B(n4626), .C(n4570), .D(n4630), .Y(n5539) );
  XOR2X1 U3248 ( .A(n5540), .B(n2153), .Y(n3417) );
  OAI21X1 U3249 ( .A(n4555), .B(n4758), .C(n5541), .Y(n5540) );
  OAI22X1 U3250 ( .A(n4624), .B(n5542), .C(n4571), .D(n5542), .Y(n5541) );
  OAI22X1 U3251 ( .A(n4572), .B(n4630), .C(n4570), .D(n4635), .Y(n5542) );
  XOR2X1 U3252 ( .A(n5543), .B(n2153), .Y(n3416) );
  OAI21X1 U3253 ( .A(n4555), .B(n4757), .C(n5544), .Y(n5543) );
  OAI22X1 U3254 ( .A(n4628), .B(n5545), .C(n4571), .D(n5545), .Y(n5544) );
  OAI22X1 U3255 ( .A(n4572), .B(n4635), .C(n4570), .D(n4640), .Y(n5545) );
  XOR2X1 U3256 ( .A(n5546), .B(n2153), .Y(n3415) );
  OAI21X1 U3257 ( .A(n4555), .B(n4755), .C(n5547), .Y(n5546) );
  OAI22X1 U3258 ( .A(n4633), .B(n5548), .C(n4571), .D(n5548), .Y(n5547) );
  OAI22X1 U3259 ( .A(n4572), .B(n4640), .C(n4570), .D(n4645), .Y(n5548) );
  XOR2X1 U3260 ( .A(n5549), .B(n2153), .Y(n3414) );
  OAI21X1 U3261 ( .A(n4555), .B(n4754), .C(n5550), .Y(n5549) );
  OAI22X1 U3262 ( .A(n4638), .B(n5551), .C(n4571), .D(n5551), .Y(n5550) );
  OAI22X1 U3263 ( .A(n4572), .B(n4645), .C(n4570), .D(n4649), .Y(n5551) );
  XOR2X1 U3264 ( .A(n5552), .B(n2153), .Y(n3413) );
  OAI21X1 U3265 ( .A(n4555), .B(n4753), .C(n5553), .Y(n5552) );
  OAI22X1 U3266 ( .A(n4643), .B(n5554), .C(n4571), .D(n5554), .Y(n5553) );
  OAI22X1 U3267 ( .A(n4572), .B(n4649), .C(n4570), .D(n4654), .Y(n5554) );
  XOR2X1 U3268 ( .A(n5555), .B(n2153), .Y(n3412) );
  OAI21X1 U3269 ( .A(n4555), .B(n4751), .C(n5556), .Y(n5555) );
  OAI22X1 U3270 ( .A(n4647), .B(n5557), .C(n4571), .D(n5557), .Y(n5556) );
  OAI22X1 U3271 ( .A(n4572), .B(n4654), .C(n4570), .D(n4659), .Y(n5557) );
  XOR2X1 U3272 ( .A(n5558), .B(n2153), .Y(n3411) );
  OAI21X1 U3273 ( .A(n4555), .B(n4750), .C(n5559), .Y(n5558) );
  OAI22X1 U3274 ( .A(n4652), .B(n5560), .C(n4571), .D(n5560), .Y(n5559) );
  OAI22X1 U3275 ( .A(n4572), .B(n4659), .C(n4570), .D(n4664), .Y(n5560) );
  XOR2X1 U3276 ( .A(n5561), .B(n2153), .Y(n3410) );
  OAI21X1 U3277 ( .A(n4555), .B(n4749), .C(n5562), .Y(n5561) );
  OAI22X1 U3278 ( .A(n4657), .B(n5563), .C(n4571), .D(n5563), .Y(n5562) );
  OAI22X1 U3279 ( .A(n4572), .B(n4664), .C(n4570), .D(n4668), .Y(n5563) );
  XOR2X1 U3280 ( .A(n5564), .B(n4717), .Y(n3409) );
  OAI21X1 U3281 ( .A(n4555), .B(n4748), .C(n5565), .Y(n5564) );
  OAI22X1 U3282 ( .A(n4662), .B(n5566), .C(n4571), .D(n5566), .Y(n5565) );
  OAI22X1 U3283 ( .A(n4572), .B(n4668), .C(n4570), .D(n4673), .Y(n5566) );
  XOR2X1 U3284 ( .A(n5567), .B(n4717), .Y(n3408) );
  OAI21X1 U3285 ( .A(n4555), .B(n4746), .C(n5568), .Y(n5567) );
  OAI22X1 U3286 ( .A(n4666), .B(n5569), .C(n4571), .D(n5569), .Y(n5568) );
  OAI22X1 U3287 ( .A(n4570), .B(n4678), .C(n4572), .D(n4673), .Y(n5569) );
  XOR2X1 U3288 ( .A(n5570), .B(n4717), .Y(n3407) );
  OAI21X1 U3289 ( .A(n4555), .B(n4745), .C(n5571), .Y(n5570) );
  OAI22X1 U3290 ( .A(n4671), .B(n5572), .C(n4571), .D(n5572), .Y(n5571) );
  OAI22X1 U3291 ( .A(n4572), .B(n4678), .C(n4570), .D(n4683), .Y(n5572) );
  XOR2X1 U3292 ( .A(n5573), .B(n4717), .Y(n3406) );
  OAI21X1 U3293 ( .A(n4555), .B(n4744), .C(n5574), .Y(n5573) );
  OAI22X1 U3294 ( .A(n4676), .B(n5575), .C(n4571), .D(n5575), .Y(n5574) );
  OAI22X1 U3295 ( .A(n4570), .B(n4688), .C(n4572), .D(n4683), .Y(n5575) );
  XOR2X1 U3296 ( .A(n5576), .B(n4717), .Y(n3405) );
  OAI21X1 U3297 ( .A(n4555), .B(n4743), .C(n5577), .Y(n5576) );
  OAI22X1 U3298 ( .A(n4681), .B(n5578), .C(n4571), .D(n5578), .Y(n5577) );
  OAI22X1 U3299 ( .A(n4572), .B(n4688), .C(n4570), .D(n4693), .Y(n5578) );
  XOR2X1 U3300 ( .A(n5579), .B(n4717), .Y(n3404) );
  OAI21X1 U3301 ( .A(n4555), .B(n4742), .C(n5580), .Y(n5579) );
  OAI22X1 U3302 ( .A(n4686), .B(n5581), .C(n4571), .D(n5581), .Y(n5580) );
  OAI22X1 U3303 ( .A(n4572), .B(n4693), .C(n4570), .D(n4697), .Y(n5581) );
  XOR2X1 U3304 ( .A(n5582), .B(n4717), .Y(n3403) );
  OAI21X1 U3305 ( .A(n4555), .B(n4741), .C(n5583), .Y(n5582) );
  OAI22X1 U3306 ( .A(n4692), .B(n5584), .C(n4571), .D(n5584), .Y(n5583) );
  OAI22X1 U3307 ( .A(n4570), .B(n4701), .C(n4572), .D(n4697), .Y(n5584) );
  XOR2X1 U3308 ( .A(n5585), .B(n4717), .Y(n3402) );
  OAI21X1 U3309 ( .A(n4555), .B(n4740), .C(n5586), .Y(n5585) );
  OAI22X1 U3310 ( .A(n4696), .B(n5587), .C(n4571), .D(n5587), .Y(n5586) );
  OAI22X1 U3311 ( .A(n4572), .B(n4701), .C(n4570), .D(n4705), .Y(n5587) );
  XOR2X1 U3312 ( .A(n5588), .B(n4717), .Y(n3401) );
  OAI21X1 U3313 ( .A(n4555), .B(n4739), .C(n5589), .Y(n5588) );
  OAI22X1 U3314 ( .A(n4700), .B(n5590), .C(n4571), .D(n5590), .Y(n5589) );
  OAI22X1 U3315 ( .A(n4572), .B(n4705), .C(n4570), .D(n4709), .Y(n5590) );
  XOR2X1 U3316 ( .A(n5591), .B(n4717), .Y(n3400) );
  OAI21X1 U3317 ( .A(n4555), .B(n4738), .C(n5592), .Y(n5591) );
  OAI22X1 U3318 ( .A(n4704), .B(n5593), .C(n4571), .D(n5593), .Y(n5592) );
  OAI22X1 U3319 ( .A(n4570), .B(n4712), .C(n4572), .D(n4709), .Y(n5593) );
  XOR2X1 U3320 ( .A(n5594), .B(n4717), .Y(n3399) );
  OAI21X1 U3321 ( .A(n4555), .B(n4737), .C(n5595), .Y(n5594) );
  OAI22X1 U3322 ( .A(n4708), .B(n5596), .C(n4571), .D(n5596), .Y(n5595) );
  OAI22X1 U3323 ( .A(n4572), .B(n4712), .C(n4570), .D(n4568), .Y(n5596) );
  XOR2X1 U3324 ( .A(n5597), .B(n4717), .Y(n3398) );
  OAI21X1 U3325 ( .A(n4555), .B(n4736), .C(n5598), .Y(n5597) );
  OAI22X1 U3326 ( .A(n4711), .B(n5599), .C(n4571), .D(n5599), .Y(n5598) );
  NAND3X1 U3327 ( .A(n4777), .B(n5601), .C(n5602), .Y(n5600) );
  OAI22X1 U3328 ( .A(n4572), .B(n4568), .C(n4735), .D(n4570), .Y(n5599) );
  NOR2X1 U3329 ( .A(n5601), .B(n4777), .Y(n5526) );
  NOR2X1 U3330 ( .A(n5603), .B(n5602), .Y(n5527) );
  XNOR2X1 U3331 ( .A(a[21]), .B(a[22]), .Y(n5602) );
  XOR2X1 U3332 ( .A(a[22]), .B(n4717), .Y(n5601) );
  XOR2X1 U3333 ( .A(a[21]), .B(n2150), .Y(n5603) );
  XOR2X1 U3334 ( .A(n4715), .B(n5604), .Y(n3396) );
  OAI22X1 U3335 ( .A(n4609), .B(n4556), .C(n4609), .D(n4774), .Y(n5604) );
  XOR2X1 U3336 ( .A(n5605), .B(n2156), .Y(n3395) );
  OAI21X1 U3337 ( .A(n4556), .B(n4765), .C(n5606), .Y(n5605) );
  AOI22X1 U3338 ( .A(n4610), .B(n5607), .C(n4606), .D(n5608), .Y(n5606) );
  XOR2X1 U3339 ( .A(n5609), .B(n2156), .Y(n3394) );
  OAI21X1 U3340 ( .A(n4556), .B(n4762), .C(n5610), .Y(n5609) );
  OAI22X1 U3341 ( .A(n4608), .B(n5611), .C(n4567), .D(n5611), .Y(n5610) );
  OAI22X1 U3342 ( .A(n4775), .B(n4611), .C(n4774), .D(n4616), .Y(n5611) );
  XOR2X1 U3343 ( .A(n5612), .B(n2156), .Y(n3393) );
  OAI21X1 U3344 ( .A(n4556), .B(n4761), .C(n5613), .Y(n5612) );
  OAI22X1 U3345 ( .A(n4610), .B(n5614), .C(n4567), .D(n5614), .Y(n5613) );
  OAI22X1 U3346 ( .A(n4775), .B(n4616), .C(n4774), .D(n4621), .Y(n5614) );
  XOR2X1 U3347 ( .A(n5615), .B(n2156), .Y(n3392) );
  OAI21X1 U3348 ( .A(n4556), .B(n4760), .C(n5616), .Y(n5615) );
  OAI22X1 U3349 ( .A(n4614), .B(n5617), .C(n4567), .D(n5617), .Y(n5616) );
  OAI22X1 U3350 ( .A(n4775), .B(n4621), .C(n4774), .D(n4626), .Y(n5617) );
  XOR2X1 U3351 ( .A(n5618), .B(n2156), .Y(n3391) );
  OAI21X1 U3352 ( .A(n4556), .B(n4759), .C(n5619), .Y(n5618) );
  OAI22X1 U3353 ( .A(n4619), .B(n5620), .C(n4567), .D(n5620), .Y(n5619) );
  OAI22X1 U3354 ( .A(n4775), .B(n4626), .C(n4774), .D(n4630), .Y(n5620) );
  XOR2X1 U3355 ( .A(n5621), .B(n2156), .Y(n3390) );
  OAI21X1 U3356 ( .A(n4556), .B(n4758), .C(n5622), .Y(n5621) );
  OAI22X1 U3357 ( .A(n4624), .B(n5623), .C(n4567), .D(n5623), .Y(n5622) );
  OAI22X1 U3358 ( .A(n4775), .B(n4630), .C(n4774), .D(n4635), .Y(n5623) );
  XOR2X1 U3359 ( .A(n5624), .B(n2156), .Y(n3389) );
  OAI21X1 U3360 ( .A(n4556), .B(n4757), .C(n5625), .Y(n5624) );
  OAI22X1 U3361 ( .A(n4628), .B(n5626), .C(n4567), .D(n5626), .Y(n5625) );
  OAI22X1 U3362 ( .A(n4775), .B(n4635), .C(n4774), .D(n4640), .Y(n5626) );
  XOR2X1 U3363 ( .A(n5627), .B(n2156), .Y(n3388) );
  OAI21X1 U3364 ( .A(n4556), .B(n4755), .C(n5628), .Y(n5627) );
  OAI22X1 U3365 ( .A(n4633), .B(n5629), .C(n4567), .D(n5629), .Y(n5628) );
  OAI22X1 U3366 ( .A(n4775), .B(n4640), .C(n4774), .D(n4645), .Y(n5629) );
  XOR2X1 U3367 ( .A(n5630), .B(n2156), .Y(n3387) );
  OAI21X1 U3368 ( .A(n4556), .B(n4754), .C(n5631), .Y(n5630) );
  OAI22X1 U3369 ( .A(n4638), .B(n5632), .C(n4567), .D(n5632), .Y(n5631) );
  OAI22X1 U3370 ( .A(n4775), .B(n4645), .C(n4774), .D(n4649), .Y(n5632) );
  XOR2X1 U3371 ( .A(n5633), .B(n2156), .Y(n3386) );
  OAI21X1 U3372 ( .A(n4556), .B(n4753), .C(n5634), .Y(n5633) );
  OAI22X1 U3373 ( .A(n4643), .B(n5635), .C(n4567), .D(n5635), .Y(n5634) );
  OAI22X1 U3374 ( .A(n4775), .B(n4649), .C(n4774), .D(n4654), .Y(n5635) );
  XOR2X1 U3375 ( .A(n5636), .B(n4715), .Y(n3385) );
  OAI21X1 U3376 ( .A(n4556), .B(n4751), .C(n5637), .Y(n5636) );
  OAI22X1 U3377 ( .A(n4647), .B(n5638), .C(n4567), .D(n5638), .Y(n5637) );
  OAI22X1 U3378 ( .A(n4775), .B(n4654), .C(n4774), .D(n4659), .Y(n5638) );
  XOR2X1 U3379 ( .A(n5639), .B(n4715), .Y(n3384) );
  OAI21X1 U3380 ( .A(n4556), .B(n4750), .C(n5640), .Y(n5639) );
  OAI22X1 U3381 ( .A(n4652), .B(n5641), .C(n4567), .D(n5641), .Y(n5640) );
  OAI22X1 U3382 ( .A(n4775), .B(n4659), .C(n4774), .D(n4664), .Y(n5641) );
  XOR2X1 U3383 ( .A(n5642), .B(n4715), .Y(n3383) );
  OAI21X1 U3384 ( .A(n4556), .B(n4749), .C(n5643), .Y(n5642) );
  OAI22X1 U3385 ( .A(n4657), .B(n5644), .C(n4567), .D(n5644), .Y(n5643) );
  OAI22X1 U3386 ( .A(n4775), .B(n4664), .C(n4774), .D(n4668), .Y(n5644) );
  XOR2X1 U3387 ( .A(n5645), .B(n4715), .Y(n3382) );
  OAI21X1 U3388 ( .A(n4556), .B(n4748), .C(n5646), .Y(n5645) );
  OAI22X1 U3389 ( .A(n4662), .B(n5647), .C(n4567), .D(n5647), .Y(n5646) );
  OAI22X1 U3390 ( .A(n4775), .B(n4668), .C(n4774), .D(n4673), .Y(n5647) );
  XOR2X1 U3391 ( .A(n5648), .B(n4715), .Y(n3381) );
  OAI21X1 U3392 ( .A(n4556), .B(n4746), .C(n5649), .Y(n5648) );
  OAI22X1 U3393 ( .A(n4666), .B(n5650), .C(n4567), .D(n5650), .Y(n5649) );
  OAI22X1 U3394 ( .A(n4774), .B(n4678), .C(n4775), .D(n4673), .Y(n5650) );
  XOR2X1 U3395 ( .A(n5651), .B(n4715), .Y(n3380) );
  OAI21X1 U3396 ( .A(n4556), .B(n4745), .C(n5652), .Y(n5651) );
  OAI22X1 U3397 ( .A(n4671), .B(n5653), .C(n4567), .D(n5653), .Y(n5652) );
  OAI22X1 U3398 ( .A(n4775), .B(n4678), .C(n4774), .D(n4683), .Y(n5653) );
  XOR2X1 U3399 ( .A(n5654), .B(n4715), .Y(n3379) );
  OAI21X1 U3400 ( .A(n4556), .B(n4744), .C(n5655), .Y(n5654) );
  OAI22X1 U3401 ( .A(n4677), .B(n5656), .C(n4567), .D(n5656), .Y(n5655) );
  OAI22X1 U3402 ( .A(n4774), .B(n4688), .C(n4775), .D(n4683), .Y(n5656) );
  XOR2X1 U3403 ( .A(n5657), .B(n2156), .Y(n3378) );
  OAI21X1 U3404 ( .A(n4556), .B(n4743), .C(n5658), .Y(n5657) );
  OAI22X1 U3405 ( .A(n4682), .B(n5659), .C(n4567), .D(n5659), .Y(n5658) );
  OAI22X1 U3406 ( .A(n4775), .B(n4688), .C(n4774), .D(n4693), .Y(n5659) );
  XOR2X1 U3407 ( .A(n5660), .B(n4715), .Y(n3377) );
  OAI21X1 U3408 ( .A(n4556), .B(n4742), .C(n5661), .Y(n5660) );
  OAI22X1 U3409 ( .A(n4687), .B(n5662), .C(n4567), .D(n5662), .Y(n5661) );
  OAI22X1 U3410 ( .A(n4775), .B(n4693), .C(n4774), .D(n4697), .Y(n5662) );
  XOR2X1 U3411 ( .A(n5663), .B(n4715), .Y(n3376) );
  OAI21X1 U3412 ( .A(n4556), .B(n4741), .C(n5664), .Y(n5663) );
  OAI22X1 U3413 ( .A(n4692), .B(n5665), .C(n4567), .D(n5665), .Y(n5664) );
  OAI22X1 U3414 ( .A(n4774), .B(n4701), .C(n4775), .D(n4697), .Y(n5665) );
  XOR2X1 U3415 ( .A(n5666), .B(n4715), .Y(n3375) );
  OAI21X1 U3416 ( .A(n4556), .B(n4740), .C(n5667), .Y(n5666) );
  OAI22X1 U3417 ( .A(n4696), .B(n5668), .C(n4567), .D(n5668), .Y(n5667) );
  OAI22X1 U3418 ( .A(n4775), .B(n4701), .C(n4774), .D(n4705), .Y(n5668) );
  XOR2X1 U3419 ( .A(n5669), .B(n4715), .Y(n3374) );
  OAI21X1 U3420 ( .A(n4556), .B(n4739), .C(n5670), .Y(n5669) );
  OAI22X1 U3421 ( .A(n4700), .B(n5671), .C(n4567), .D(n5671), .Y(n5670) );
  NAND3X1 U3422 ( .A(n5673), .B(n5674), .C(n5675), .Y(n5672) );
  OAI22X1 U3423 ( .A(n4775), .B(n4705), .C(n4709), .D(n4774), .Y(n5671) );
  NOR2X1 U3424 ( .A(n5674), .B(n5673), .Y(n5607) );
  NOR2X1 U3425 ( .A(n4776), .B(n5675), .Y(n5608) );
  XNOR2X1 U3426 ( .A(a[24]), .B(a[25]), .Y(n5675) );
  XOR2X1 U3427 ( .A(a[25]), .B(n4715), .Y(n5674) );
  XNOR2X1 U3428 ( .A(a[24]), .B(n4717), .Y(n5673) );
  XOR2X1 U3429 ( .A(n4713), .B(n5676), .Y(n3372) );
  OAI22X1 U3430 ( .A(n4609), .B(n4557), .C(n4609), .D(n4770), .Y(n5676) );
  XOR2X1 U3431 ( .A(n5677), .B(n2159), .Y(n3371) );
  OAI21X1 U3432 ( .A(n4557), .B(n4765), .C(n5678), .Y(n5677) );
  AOI22X1 U3433 ( .A(n4610), .B(n5679), .C(n4605), .D(n5680), .Y(n5678) );
  XOR2X1 U3434 ( .A(n5681), .B(n2159), .Y(n3370) );
  OAI21X1 U3435 ( .A(n4557), .B(n4762), .C(n5682), .Y(n5681) );
  OAI22X1 U3436 ( .A(n4608), .B(n5683), .C(n4771), .D(n5683), .Y(n5682) );
  OAI22X1 U3437 ( .A(n4772), .B(n4611), .C(n4770), .D(n4616), .Y(n5683) );
  XOR2X1 U3438 ( .A(n5684), .B(n2159), .Y(n3369) );
  OAI21X1 U3439 ( .A(n4557), .B(n4761), .C(n5685), .Y(n5684) );
  OAI22X1 U3440 ( .A(n4610), .B(n5686), .C(n4771), .D(n5686), .Y(n5685) );
  OAI22X1 U3441 ( .A(n4772), .B(n4616), .C(n4770), .D(n4621), .Y(n5686) );
  XOR2X1 U3442 ( .A(n5687), .B(n2159), .Y(n3368) );
  OAI21X1 U3443 ( .A(n4557), .B(n4760), .C(n5688), .Y(n5687) );
  OAI22X1 U3444 ( .A(n4615), .B(n5689), .C(n4771), .D(n5689), .Y(n5688) );
  OAI22X1 U3445 ( .A(n4772), .B(n4621), .C(n4770), .D(n4626), .Y(n5689) );
  XOR2X1 U3446 ( .A(n5690), .B(n2159), .Y(n3367) );
  OAI21X1 U3447 ( .A(n4557), .B(n4759), .C(n5691), .Y(n5690) );
  OAI22X1 U3448 ( .A(n4620), .B(n5692), .C(n4771), .D(n5692), .Y(n5691) );
  OAI22X1 U3449 ( .A(n4772), .B(n4626), .C(n4770), .D(n4630), .Y(n5692) );
  XOR2X1 U3450 ( .A(n5693), .B(n2159), .Y(n3366) );
  OAI21X1 U3451 ( .A(n4557), .B(n4758), .C(n5694), .Y(n5693) );
  OAI22X1 U3452 ( .A(n4625), .B(n5695), .C(n4771), .D(n5695), .Y(n5694) );
  OAI22X1 U3453 ( .A(n4772), .B(n4630), .C(n4770), .D(n4635), .Y(n5695) );
  XOR2X1 U3454 ( .A(n5696), .B(n2159), .Y(n3365) );
  OAI21X1 U3455 ( .A(n4557), .B(n4757), .C(n5697), .Y(n5696) );
  OAI22X1 U3456 ( .A(n4629), .B(n5698), .C(n4771), .D(n5698), .Y(n5697) );
  OAI22X1 U3457 ( .A(n4772), .B(n4635), .C(n4770), .D(n4640), .Y(n5698) );
  XOR2X1 U3458 ( .A(n5699), .B(n2159), .Y(n3364) );
  OAI21X1 U3459 ( .A(n4557), .B(n4755), .C(n5700), .Y(n5699) );
  OAI22X1 U3460 ( .A(n4634), .B(n5701), .C(n4771), .D(n5701), .Y(n5700) );
  OAI22X1 U3461 ( .A(n4772), .B(n4640), .C(n4770), .D(n4645), .Y(n5701) );
  XOR2X1 U3462 ( .A(n5702), .B(n4713), .Y(n3363) );
  OAI21X1 U3463 ( .A(n4557), .B(n4754), .C(n5703), .Y(n5702) );
  OAI22X1 U3464 ( .A(n4639), .B(n5704), .C(n4771), .D(n5704), .Y(n5703) );
  OAI22X1 U3465 ( .A(n4772), .B(n4645), .C(n4770), .D(n4649), .Y(n5704) );
  XOR2X1 U3466 ( .A(n5705), .B(n4713), .Y(n3362) );
  OAI21X1 U3467 ( .A(n4557), .B(n4753), .C(n5706), .Y(n5705) );
  OAI22X1 U3468 ( .A(n4644), .B(n5707), .C(n4771), .D(n5707), .Y(n5706) );
  OAI22X1 U3469 ( .A(n4772), .B(n4649), .C(n4770), .D(n4654), .Y(n5707) );
  XOR2X1 U3470 ( .A(n5708), .B(n4713), .Y(n3361) );
  OAI21X1 U3471 ( .A(n4557), .B(n4751), .C(n5709), .Y(n5708) );
  OAI22X1 U3472 ( .A(n4648), .B(n5710), .C(n4771), .D(n5710), .Y(n5709) );
  OAI22X1 U3473 ( .A(n4772), .B(n4654), .C(n4770), .D(n4659), .Y(n5710) );
  XOR2X1 U3474 ( .A(n5711), .B(n4713), .Y(n3360) );
  OAI21X1 U3475 ( .A(n4557), .B(n4750), .C(n5712), .Y(n5711) );
  OAI22X1 U3476 ( .A(n4653), .B(n5713), .C(n4771), .D(n5713), .Y(n5712) );
  OAI22X1 U3477 ( .A(n4772), .B(n4659), .C(n4770), .D(n4664), .Y(n5713) );
  XOR2X1 U3478 ( .A(n5714), .B(n4713), .Y(n3359) );
  OAI21X1 U3479 ( .A(n4557), .B(n4749), .C(n5715), .Y(n5714) );
  OAI22X1 U3480 ( .A(n4658), .B(n5716), .C(n4771), .D(n5716), .Y(n5715) );
  OAI22X1 U3481 ( .A(n4772), .B(n4664), .C(n4770), .D(n4668), .Y(n5716) );
  XOR2X1 U3482 ( .A(n5717), .B(n4713), .Y(n3358) );
  OAI21X1 U3483 ( .A(n4557), .B(n4748), .C(n5718), .Y(n5717) );
  OAI22X1 U3484 ( .A(n4663), .B(n5719), .C(n4771), .D(n5719), .Y(n5718) );
  OAI22X1 U3485 ( .A(n4772), .B(n4668), .C(n4770), .D(n4673), .Y(n5719) );
  XOR2X1 U3486 ( .A(n5720), .B(n4713), .Y(n3357) );
  OAI21X1 U3487 ( .A(n4557), .B(n4746), .C(n5721), .Y(n5720) );
  OAI22X1 U3488 ( .A(n4667), .B(n5722), .C(n4771), .D(n5722), .Y(n5721) );
  OAI22X1 U3489 ( .A(n4770), .B(n4678), .C(n4772), .D(n4673), .Y(n5722) );
  XOR2X1 U3490 ( .A(n5723), .B(n4713), .Y(n3356) );
  OAI21X1 U3491 ( .A(n4557), .B(n4745), .C(n5724), .Y(n5723) );
  OAI22X1 U3492 ( .A(n4672), .B(n5725), .C(n4771), .D(n5725), .Y(n5724) );
  OAI22X1 U3493 ( .A(n4772), .B(n4678), .C(n4770), .D(n4683), .Y(n5725) );
  XOR2X1 U3494 ( .A(n5726), .B(n4713), .Y(n3355) );
  OAI21X1 U3495 ( .A(n4557), .B(n4744), .C(n5727), .Y(n5726) );
  OAI22X1 U3496 ( .A(n4677), .B(n5728), .C(n4771), .D(n5728), .Y(n5727) );
  OAI22X1 U3497 ( .A(n4770), .B(n4688), .C(n4772), .D(n4683), .Y(n5728) );
  XOR2X1 U3498 ( .A(n5729), .B(n4713), .Y(n3354) );
  OAI21X1 U3499 ( .A(n4557), .B(n4743), .C(n5730), .Y(n5729) );
  OAI22X1 U3500 ( .A(n4682), .B(n5731), .C(n4771), .D(n5731), .Y(n5730) );
  OAI22X1 U3501 ( .A(n4772), .B(n4688), .C(n4770), .D(n4693), .Y(n5731) );
  XOR2X1 U3502 ( .A(n5732), .B(n4713), .Y(n3353) );
  OAI21X1 U3503 ( .A(n4557), .B(n4742), .C(n5733), .Y(n5732) );
  OAI22X1 U3504 ( .A(n4687), .B(n5734), .C(n4771), .D(n5734), .Y(n5733) );
  NAND3X1 U3505 ( .A(n5736), .B(n5737), .C(n5738), .Y(n5735) );
  OAI22X1 U3506 ( .A(n4772), .B(n4693), .C(n4697), .D(n4770), .Y(n5734) );
  NOR2X1 U3507 ( .A(n5737), .B(n5736), .Y(n5679) );
  NOR2X1 U3508 ( .A(n4773), .B(n5738), .Y(n5680) );
  XNOR2X1 U3509 ( .A(a[27]), .B(a[28]), .Y(n5738) );
  XOR2X1 U3510 ( .A(a[28]), .B(n4713), .Y(n5737) );
  XNOR2X1 U3511 ( .A(a[27]), .B(n4715), .Y(n5736) );
  OAI22X1 U3512 ( .A(n4767), .B(n4609), .C(n4558), .D(n4609), .Y(n3351) );
  OAI21X1 U3513 ( .A(n4558), .B(n4765), .C(n5739), .Y(n3350) );
  AOI22X1 U3514 ( .A(n4610), .B(n5740), .C(n4605), .D(n5741), .Y(n5739) );
  OAI21X1 U3515 ( .A(n4558), .B(n4762), .C(n5742), .Y(n3349) );
  OAI22X1 U3516 ( .A(n4607), .B(n5743), .C(n4766), .D(n5743), .Y(n5742) );
  OAI22X1 U3517 ( .A(n4768), .B(n4611), .C(n4767), .D(n4616), .Y(n5743) );
  OAI21X1 U3518 ( .A(n4558), .B(n4761), .C(n5744), .Y(n3348) );
  OAI22X1 U3519 ( .A(n4610), .B(n5745), .C(n4766), .D(n5745), .Y(n5744) );
  OAI22X1 U3520 ( .A(n4768), .B(n4616), .C(n4767), .D(n4621), .Y(n5745) );
  OAI21X1 U3521 ( .A(n4558), .B(n4760), .C(n5746), .Y(n3347) );
  OAI22X1 U3522 ( .A(n4615), .B(n5747), .C(n4766), .D(n5747), .Y(n5746) );
  OAI22X1 U3523 ( .A(n4768), .B(n4621), .C(n4767), .D(n4626), .Y(n5747) );
  OAI21X1 U3524 ( .A(n4558), .B(n4759), .C(n5748), .Y(n3346) );
  OAI22X1 U3525 ( .A(n4620), .B(n5749), .C(n4766), .D(n5749), .Y(n5748) );
  OAI22X1 U3526 ( .A(n4768), .B(n4626), .C(n4767), .D(n4630), .Y(n5749) );
  OAI21X1 U3527 ( .A(n4558), .B(n4758), .C(n5750), .Y(n3345) );
  OAI22X1 U3528 ( .A(n4625), .B(n5751), .C(n4766), .D(n5751), .Y(n5750) );
  OAI22X1 U3529 ( .A(n4768), .B(n4630), .C(n4767), .D(n4635), .Y(n5751) );
  OAI21X1 U3530 ( .A(n4558), .B(n4757), .C(n5752), .Y(n3344) );
  OAI22X1 U3531 ( .A(n4629), .B(n5753), .C(n4766), .D(n5753), .Y(n5752) );
  OAI22X1 U3532 ( .A(n4768), .B(n4635), .C(n4767), .D(n4640), .Y(n5753) );
  OAI21X1 U3533 ( .A(n4558), .B(n4755), .C(n5754), .Y(n3343) );
  OAI22X1 U3534 ( .A(n4634), .B(n5755), .C(n4766), .D(n5755), .Y(n5754) );
  OAI22X1 U3535 ( .A(n4768), .B(n4640), .C(n4767), .D(n4645), .Y(n5755) );
  OAI21X1 U3536 ( .A(n4558), .B(n4754), .C(n5756), .Y(n3342) );
  OAI22X1 U3537 ( .A(n4639), .B(n5757), .C(n4766), .D(n5757), .Y(n5756) );
  OAI22X1 U3538 ( .A(n4768), .B(n4645), .C(n4767), .D(n4649), .Y(n5757) );
  OAI21X1 U3539 ( .A(n4558), .B(n4753), .C(n5758), .Y(n3341) );
  OAI22X1 U3540 ( .A(n4644), .B(n5759), .C(n4766), .D(n5759), .Y(n5758) );
  OAI22X1 U3541 ( .A(n4768), .B(n4649), .C(n4767), .D(n4654), .Y(n5759) );
  OAI21X1 U3542 ( .A(n4558), .B(n4751), .C(n5760), .Y(n3340) );
  OAI22X1 U3543 ( .A(n4648), .B(n5761), .C(n4766), .D(n5761), .Y(n5760) );
  OAI22X1 U3544 ( .A(n4768), .B(n4654), .C(n4767), .D(n4659), .Y(n5761) );
  OAI21X1 U3545 ( .A(n4558), .B(n4750), .C(n5762), .Y(n3339) );
  OAI22X1 U3546 ( .A(n4653), .B(n5763), .C(n4766), .D(n5763), .Y(n5762) );
  OAI22X1 U3547 ( .A(n4768), .B(n4659), .C(n4767), .D(n4664), .Y(n5763) );
  OAI21X1 U3548 ( .A(n4558), .B(n4749), .C(n5764), .Y(n3338) );
  OAI22X1 U3549 ( .A(n4658), .B(n5765), .C(n4766), .D(n5765), .Y(n5764) );
  OAI22X1 U3550 ( .A(n4768), .B(n4664), .C(n4767), .D(n4668), .Y(n5765) );
  OAI21X1 U3551 ( .A(n4558), .B(n4746), .C(n5766), .Y(n3337) );
  OAI22X1 U3552 ( .A(n4667), .B(n5767), .C(n4766), .D(n5767), .Y(n5766) );
  OAI22X1 U3553 ( .A(n4767), .B(n4678), .C(n4768), .D(n4673), .Y(n5767) );
  OAI21X1 U3554 ( .A(n4558), .B(n4745), .C(n5768), .Y(n3336) );
  OAI22X1 U3555 ( .A(n4672), .B(n5769), .C(n4766), .D(n5769), .Y(n5768) );
  OAI22X1 U3556 ( .A(n4768), .B(n4678), .C(n4683), .D(n4767), .Y(n5769) );
  OAI21X1 U3557 ( .A(n4558), .B(n4748), .C(n5770), .Y(n2429) );
  OAI22X1 U3558 ( .A(n4663), .B(n5771), .C(n4766), .D(n5771), .Y(n5770) );
  NAND3X1 U3559 ( .A(n5773), .B(a[31]), .C(n5774), .Y(n5772) );
  OAI22X1 U3560 ( .A(n4768), .B(n4668), .C(n4767), .D(n4673), .Y(n5771) );
  NOR2X1 U3561 ( .A(n5773), .B(a[31]), .Y(n5740) );
  NOR2X1 U3562 ( .A(n4769), .B(n5774), .Y(n5741) );
  XNOR2X1 U3563 ( .A(a[30]), .B(a[31]), .Y(n5774) );
  XNOR2X1 U3564 ( .A(a[30]), .B(n4713), .Y(n5773) );
endmodule


module poly5_DW_mult_uns_0 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n2132, n2135, n2138, n2141, n2144, n2147, n2150, n2153, n2156, n2159,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748;
  assign n2132 = a[2];
  assign n2135 = a[5];
  assign n2138 = a[8];
  assign n2141 = a[11];
  assign n2144 = a[14];
  assign n2147 = a[17];
  assign n2150 = a[20];
  assign n2153 = a[23];
  assign n2156 = a[26];
  assign n2159 = a[29];

  FAX1 U336 ( .A(n2406), .B(n2417), .C(n2353), .YC(n2352), .YS(product[46]) );
  FAX1 U337 ( .A(n2431), .B(n2418), .C(n2354), .YC(n2353), .YS(product[45]) );
  FAX1 U338 ( .A(n2444), .B(n2432), .C(n2355), .YC(n2354), .YS(product[44]) );
  FAX1 U339 ( .A(n2445), .B(n2458), .C(n2356), .YC(n2355), .YS(product[43]) );
  FAX1 U340 ( .A(n2474), .B(n2459), .C(n2357), .YC(n2356), .YS(product[42]) );
  FAX1 U341 ( .A(n2489), .B(n2475), .C(n2358), .YC(n2357), .YS(product[41]) );
  FAX1 U342 ( .A(n2490), .B(n2504), .C(n2359), .YC(n2358), .YS(product[40]) );
  FAX1 U343 ( .A(n2522), .B(n2505), .C(n2360), .YC(n2359), .YS(product[39]) );
  FAX1 U344 ( .A(n2539), .B(n2523), .C(n2361), .YC(n2360), .YS(product[38]) );
  FAX1 U345 ( .A(n2540), .B(n2556), .C(n2362), .YC(n2361), .YS(product[37]) );
  FAX1 U346 ( .A(n2574), .B(n2557), .C(n2363), .YC(n2362), .YS(product[36]) );
  FAX1 U347 ( .A(n2592), .B(n2575), .C(n2364), .YC(n2363), .YS(product[35]) );
  FAX1 U348 ( .A(n2593), .B(n2610), .C(n2365), .YC(n2364), .YS(product[34]) );
  FAX1 U349 ( .A(n2628), .B(n2611), .C(n2366), .YC(n2365), .YS(product[33]) );
  FAX1 U350 ( .A(n3629), .B(n2629), .C(n2367), .YC(n2366), .YS(product[32]) );
  FAX1 U351 ( .A(n2647), .B(n3630), .C(n2368), .YC(n2367), .YS(product[31]) );
  FAX1 U352 ( .A(n2665), .B(n3631), .C(n2369), .YC(n2368), .YS(product[30]) );
  FAX1 U353 ( .A(n2683), .B(n3632), .C(n2370), .YC(n2369), .YS(product[29]) );
  FAX1 U354 ( .A(n2701), .B(n3633), .C(n2371), .YC(n2370), .YS(product[28]) );
  FAX1 U355 ( .A(n2719), .B(n3634), .C(n2372), .YC(n2371), .YS(product[27]) );
  FAX1 U356 ( .A(n2737), .B(n3635), .C(n2373), .YC(n2372), .YS(product[26]) );
  FAX1 U357 ( .A(n2753), .B(n3636), .C(n2374), .YC(n2373), .YS(product[25]) );
  FAX1 U358 ( .A(n2769), .B(n3637), .C(n2375), .YC(n2374), .YS(product[24]) );
  FAX1 U359 ( .A(n2785), .B(n3638), .C(n2376), .YC(n2375), .YS(product[23]) );
  FAX1 U360 ( .A(n2799), .B(n3639), .C(n2377), .YC(n2376), .YS(product[22]) );
  FAX1 U361 ( .A(n2813), .B(n3640), .C(n2378), .YC(n2377), .YS(product[21]) );
  FAX1 U362 ( .A(n2827), .B(n3641), .C(n2379), .YC(n2378), .YS(product[20]) );
  FAX1 U363 ( .A(n2839), .B(n3642), .C(n2380), .YC(n2379), .YS(product[19]) );
  FAX1 U364 ( .A(n2851), .B(n3643), .C(n2381), .YC(n2380), .YS(product[18]) );
  FAX1 U365 ( .A(n2863), .B(n3644), .C(n2382), .YC(n2381), .YS(product[17]) );
  FAX1 U366 ( .A(n2873), .B(n3645), .C(n2383), .YC(n2382), .YS(product[16]) );
  FAX1 U367 ( .A(n2883), .B(n3646), .C(n2384), .YC(n2383), .YS(product[15]) );
  FAX1 U368 ( .A(n2893), .B(n3647), .C(n2385), .YC(n2384), .YS(product[14]) );
  FAX1 U369 ( .A(n2901), .B(n3648), .C(n2386), .YC(n2385), .YS(product[13]) );
  FAX1 U370 ( .A(n2909), .B(n3649), .C(n2387), .YC(n2386), .YS(product[12]) );
  FAX1 U371 ( .A(n2917), .B(n3650), .C(n2388), .YC(n2387), .YS(product[11]) );
  FAX1 U372 ( .A(n2923), .B(n3651), .C(n2389), .YC(n2388), .YS(product[10]) );
  FAX1 U373 ( .A(n2929), .B(n3652), .C(n2390), .YC(n2389), .YS(product[9]) );
  FAX1 U374 ( .A(n2935), .B(n3653), .C(n2391), .YC(n2390), .YS(product[8]) );
  FAX1 U375 ( .A(n2939), .B(n3654), .C(n2392), .YC(n2391), .YS(product[7]) );
  FAX1 U376 ( .A(n2943), .B(n3655), .C(n2393), .YC(n2392), .YS(product[6]) );
  FAX1 U377 ( .A(n2947), .B(n3656), .C(n2394), .YC(n2393), .YS(product[5]) );
  FAX1 U378 ( .A(n3657), .B(n2949), .C(n2395), .YC(n2394), .YS(product[4]) );
  FAX1 U379 ( .A(n2951), .B(n3658), .C(n2396), .YC(n2395), .YS(product[3]) );
  HAX1 U380 ( .A(n3659), .B(n2397), .YC(n2396), .YS(product[2]) );
  HAX1 U381 ( .A(n2398), .B(n3660), .YC(n2397), .YS(product[1]) );
  HAX1 U382 ( .A(n2132), .B(n3661), .YC(n2398), .YS(product[0]) );
  FAX1 U384 ( .A(n2408), .B(n3455), .C(n2419), .YC(n2405), .YS(n2406) );
  FAX1 U385 ( .A(n2410), .B(n2421), .C(n3425), .YC(n2407), .YS(n2408) );
  FAX1 U386 ( .A(n2412), .B(n3398), .C(n2423), .YC(n2409), .YS(n2410) );
  FAX1 U387 ( .A(n2414), .B(n2425), .C(n3374), .YC(n2411), .YS(n2412) );
  FAX1 U388 ( .A(n2416), .B(n3353), .C(n2427), .YC(n2413), .YS(n2414) );
  FAX1 U389 ( .A(n4603), .B(n2429), .C(n3336), .YC(n2415), .YS(n2416) );
  FAX1 U390 ( .A(n3456), .B(n2420), .C(n3488), .YC(n2417), .YS(n2418) );
  FAX1 U391 ( .A(n2435), .B(n2422), .C(n2433), .YC(n2419), .YS(n2420) );
  FAX1 U392 ( .A(n3399), .B(n2424), .C(n3426), .YC(n2421), .YS(n2422) );
  FAX1 U393 ( .A(n2439), .B(n2426), .C(n2437), .YC(n2423), .YS(n2424) );
  FAX1 U394 ( .A(n2441), .B(n2428), .C(n3375), .YC(n2425), .YS(n2426) );
  FAX1 U395 ( .A(n4723), .B(n3337), .C(n3354), .YC(n2427), .YS(n2428) );
  FAX1 U397 ( .A(n2446), .B(n2434), .C(n3489), .YC(n2431), .YS(n2432) );
  FAX1 U398 ( .A(n2448), .B(n2436), .C(n3457), .YC(n2433), .YS(n2434) );
  FAX1 U399 ( .A(n2450), .B(n2438), .C(n3427), .YC(n2435), .YS(n2436) );
  FAX1 U400 ( .A(n2452), .B(n2440), .C(n3400), .YC(n2437), .YS(n2438) );
  FAX1 U401 ( .A(n2454), .B(n2442), .C(n3376), .YC(n2439), .YS(n2440) );
  FAX1 U402 ( .A(n2456), .B(n4723), .C(n3355), .YC(n2441), .YS(n2442) );
  FAX1 U404 ( .A(n2447), .B(n3490), .C(n2460), .YC(n2444), .YS(n2445) );
  FAX1 U405 ( .A(n2449), .B(n2462), .C(n3458), .YC(n2446), .YS(n2447) );
  FAX1 U406 ( .A(n2451), .B(n3428), .C(n2464), .YC(n2448), .YS(n2449) );
  FAX1 U407 ( .A(n2453), .B(n2466), .C(n3401), .YC(n2450), .YS(n2451) );
  FAX1 U408 ( .A(n2455), .B(n3377), .C(n2468), .YC(n2452), .YS(n2453) );
  FAX1 U409 ( .A(n2457), .B(n3356), .C(n2470), .YC(n2454), .YS(n2455) );
  FAX1 U410 ( .A(n4757), .B(n2472), .C(n3338), .YC(n2456), .YS(n2457) );
  FAX1 U411 ( .A(n3491), .B(n2461), .C(n3523), .YC(n2458), .YS(n2459) );
  FAX1 U412 ( .A(n2478), .B(n2463), .C(n2476), .YC(n2460), .YS(n2461) );
  FAX1 U413 ( .A(n3429), .B(n2465), .C(n3459), .YC(n2462), .YS(n2463) );
  FAX1 U414 ( .A(n2482), .B(n2467), .C(n2480), .YC(n2464), .YS(n2465) );
  FAX1 U415 ( .A(n2484), .B(n2469), .C(n3402), .YC(n2466), .YS(n2467) );
  FAX1 U416 ( .A(n2486), .B(n2471), .C(n3378), .YC(n2468), .YS(n2469) );
  FAX1 U417 ( .A(n4728), .B(n3339), .C(n3357), .YC(n2470), .YS(n2471) );
  FAX1 U419 ( .A(n2491), .B(n2477), .C(n3524), .YC(n2474), .YS(n2475) );
  FAX1 U420 ( .A(n2493), .B(n2479), .C(n3492), .YC(n2476), .YS(n2477) );
  FAX1 U421 ( .A(n2495), .B(n2481), .C(n3460), .YC(n2478), .YS(n2479) );
  FAX1 U422 ( .A(n2497), .B(n2483), .C(n3430), .YC(n2480), .YS(n2481) );
  FAX1 U423 ( .A(n2499), .B(n2485), .C(n3403), .YC(n2482), .YS(n2483) );
  FAX1 U424 ( .A(n2501), .B(n2487), .C(n3379), .YC(n2484), .YS(n2485) );
  FAX1 U425 ( .A(n3340), .B(n4728), .C(n3358), .YC(n2486), .YS(n2487) );
  FAX1 U427 ( .A(n2492), .B(n3525), .C(n2506), .YC(n2489), .YS(n2490) );
  FAX1 U428 ( .A(n2494), .B(n2508), .C(n3493), .YC(n2491), .YS(n2492) );
  FAX1 U429 ( .A(n2496), .B(n3461), .C(n2510), .YC(n2493), .YS(n2494) );
  FAX1 U430 ( .A(n2498), .B(n2512), .C(n3431), .YC(n2495), .YS(n2496) );
  FAX1 U431 ( .A(n2500), .B(n3404), .C(n2514), .YC(n2497), .YS(n2498) );
  FAX1 U432 ( .A(n2502), .B(n3380), .C(n2516), .YC(n2499), .YS(n2500) );
  FAX1 U433 ( .A(n2503), .B(n2518), .C(n3359), .YC(n2501), .YS(n2502) );
  FAX1 U434 ( .A(n4759), .B(n2520), .C(n3341), .YC(n2472), .YS(n2503) );
  FAX1 U435 ( .A(n3526), .B(n2507), .C(n3558), .YC(n2504), .YS(n2505) );
  FAX1 U436 ( .A(n2526), .B(n2509), .C(n2524), .YC(n2506), .YS(n2507) );
  FAX1 U437 ( .A(n3462), .B(n2511), .C(n3494), .YC(n2508), .YS(n2509) );
  FAX1 U438 ( .A(n2530), .B(n2513), .C(n2528), .YC(n2510), .YS(n2511) );
  FAX1 U439 ( .A(n2532), .B(n2515), .C(n3432), .YC(n2512), .YS(n2513) );
  FAX1 U440 ( .A(n2534), .B(n2517), .C(n3405), .YC(n2514), .YS(n2515) );
  FAX1 U441 ( .A(n3360), .B(n2519), .C(n3381), .YC(n2516), .YS(n2517) );
  FAX1 U442 ( .A(n4732), .B(n3342), .C(n2536), .YC(n2518), .YS(n2519) );
  FAX1 U444 ( .A(n2541), .B(n2525), .C(n3559), .YC(n2522), .YS(n2523) );
  FAX1 U445 ( .A(n2543), .B(n2527), .C(n3527), .YC(n2524), .YS(n2525) );
  FAX1 U446 ( .A(n2545), .B(n2529), .C(n3495), .YC(n2526), .YS(n2527) );
  FAX1 U447 ( .A(n2547), .B(n2531), .C(n3463), .YC(n2528), .YS(n2529) );
  FAX1 U448 ( .A(n2549), .B(n2533), .C(n3433), .YC(n2530), .YS(n2531) );
  FAX1 U449 ( .A(n2551), .B(n2535), .C(n3406), .YC(n2532), .YS(n2533) );
  FAX1 U450 ( .A(n2553), .B(n2537), .C(n3382), .YC(n2534), .YS(n2535) );
  FAX1 U451 ( .A(n3343), .B(n4732), .C(n3361), .YC(n2536), .YS(n2537) );
  FAX1 U453 ( .A(n2542), .B(n3560), .C(n2558), .YC(n2539), .YS(n2540) );
  FAX1 U454 ( .A(n2544), .B(n2560), .C(n3528), .YC(n2541), .YS(n2542) );
  FAX1 U455 ( .A(n2546), .B(n3496), .C(n2562), .YC(n2543), .YS(n2544) );
  FAX1 U456 ( .A(n2548), .B(n2564), .C(n3464), .YC(n2545), .YS(n2546) );
  FAX1 U457 ( .A(n2550), .B(n3434), .C(n2566), .YC(n2547), .YS(n2548) );
  FAX1 U458 ( .A(n2552), .B(n3407), .C(n2568), .YC(n2549), .YS(n2550) );
  FAX1 U459 ( .A(n2554), .B(n2570), .C(n3383), .YC(n2551), .YS(n2552) );
  FAX1 U460 ( .A(n2555), .B(n2572), .C(n3362), .YC(n2553), .YS(n2554) );
  FAX1 U461 ( .A(n4619), .B(n4761), .C(n3344), .YC(n2520), .YS(n2555) );
  FAX1 U462 ( .A(n3561), .B(n2559), .C(n3593), .YC(n2556), .YS(n2557) );
  FAX1 U463 ( .A(n2578), .B(n2561), .C(n2576), .YC(n2558), .YS(n2559) );
  FAX1 U464 ( .A(n3497), .B(n2563), .C(n3529), .YC(n2560), .YS(n2561) );
  FAX1 U465 ( .A(n2582), .B(n2565), .C(n2580), .YC(n2562), .YS(n2563) );
  FAX1 U466 ( .A(n2584), .B(n2567), .C(n3465), .YC(n2564), .YS(n2565) );
  FAX1 U467 ( .A(n2586), .B(n2569), .C(n3435), .YC(n2566), .YS(n2567) );
  FAX1 U468 ( .A(n3384), .B(n2571), .C(n3408), .YC(n2568), .YS(n2569) );
  FAX1 U469 ( .A(n3363), .B(n2573), .C(n2588), .YC(n2570), .YS(n2571) );
  FAX1 U470 ( .A(n2132), .B(n3345), .C(n2590), .YC(n2572), .YS(n2573) );
  FAX1 U471 ( .A(n2594), .B(n2577), .C(n3594), .YC(n2574), .YS(n2575) );
  FAX1 U472 ( .A(n3530), .B(n2579), .C(n3562), .YC(n2576), .YS(n2577) );
  FAX1 U473 ( .A(n2598), .B(n2581), .C(n2596), .YC(n2578), .YS(n2579) );
  FAX1 U474 ( .A(n3466), .B(n2583), .C(n3498), .YC(n2580), .YS(n2581) );
  FAX1 U475 ( .A(n3436), .B(n2585), .C(n2600), .YC(n2582), .YS(n2583) );
  FAX1 U476 ( .A(n2604), .B(n2587), .C(n2602), .YC(n2584), .YS(n2585) );
  FAX1 U477 ( .A(n3385), .B(n2589), .C(n3409), .YC(n2586), .YS(n2587) );
  FAX1 U478 ( .A(n3364), .B(n2591), .C(n2606), .YC(n2588), .YS(n2589) );
  FAX1 U479 ( .A(n2132), .B(n3346), .C(n2608), .YC(n2590), .YS(n2591) );
  FAX1 U480 ( .A(n2595), .B(n2612), .C(n3595), .YC(n2592), .YS(n2593) );
  FAX1 U481 ( .A(n2597), .B(n2614), .C(n3563), .YC(n2594), .YS(n2595) );
  FAX1 U482 ( .A(n2599), .B(n2616), .C(n3531), .YC(n2596), .YS(n2597) );
  FAX1 U483 ( .A(n2601), .B(n2618), .C(n3499), .YC(n2598), .YS(n2599) );
  FAX1 U484 ( .A(n2603), .B(n2620), .C(n3467), .YC(n2600), .YS(n2601) );
  FAX1 U485 ( .A(n2605), .B(n2622), .C(n3437), .YC(n2602), .YS(n2603) );
  FAX1 U486 ( .A(n2607), .B(n2624), .C(n3410), .YC(n2604), .YS(n2605) );
  FAX1 U487 ( .A(n2609), .B(n2626), .C(n3386), .YC(n2606), .YS(n2607) );
  FAX1 U488 ( .A(n2132), .B(n3347), .C(n3365), .YC(n2608), .YS(n2609) );
  FAX1 U489 ( .A(n2613), .B(n3596), .C(n3628), .YC(n2610), .YS(n2611) );
  FAX1 U490 ( .A(n2615), .B(n3564), .C(n2630), .YC(n2612), .YS(n2613) );
  FAX1 U491 ( .A(n2617), .B(n3532), .C(n2632), .YC(n2614), .YS(n2615) );
  FAX1 U492 ( .A(n2619), .B(n3500), .C(n2634), .YC(n2616), .YS(n2617) );
  FAX1 U493 ( .A(n2621), .B(n3468), .C(n2636), .YC(n2618), .YS(n2619) );
  FAX1 U494 ( .A(n2623), .B(n3438), .C(n2638), .YC(n2620), .YS(n2621) );
  FAX1 U495 ( .A(n2625), .B(n3411), .C(n2640), .YC(n2622), .YS(n2623) );
  FAX1 U496 ( .A(n2627), .B(n3387), .C(n2642), .YC(n2624), .YS(n2625) );
  FAX1 U497 ( .A(n3348), .B(n3366), .C(n2644), .YC(n2626), .YS(n2627) );
  FAX1 U498 ( .A(n2631), .B(n3597), .C(n2646), .YC(n2628), .YS(n2629) );
  FAX1 U499 ( .A(n2633), .B(n3565), .C(n2648), .YC(n2630), .YS(n2631) );
  FAX1 U500 ( .A(n2635), .B(n3533), .C(n2650), .YC(n2632), .YS(n2633) );
  FAX1 U501 ( .A(n2637), .B(n3501), .C(n2652), .YC(n2634), .YS(n2635) );
  FAX1 U502 ( .A(n2639), .B(n3469), .C(n2654), .YC(n2636), .YS(n2637) );
  FAX1 U503 ( .A(n2641), .B(n3439), .C(n2656), .YC(n2638), .YS(n2639) );
  FAX1 U504 ( .A(n2643), .B(n3412), .C(n2658), .YC(n2640), .YS(n2641) );
  FAX1 U505 ( .A(n2645), .B(n3388), .C(n2660), .YC(n2642), .YS(n2643) );
  FAX1 U506 ( .A(n3349), .B(n3367), .C(n2662), .YC(n2644), .YS(n2645) );
  FAX1 U507 ( .A(n2649), .B(n3598), .C(n2664), .YC(n2646), .YS(n2647) );
  FAX1 U508 ( .A(n2651), .B(n3566), .C(n2666), .YC(n2648), .YS(n2649) );
  FAX1 U509 ( .A(n2653), .B(n3534), .C(n2668), .YC(n2650), .YS(n2651) );
  FAX1 U510 ( .A(n2655), .B(n3502), .C(n2670), .YC(n2652), .YS(n2653) );
  FAX1 U511 ( .A(n2657), .B(n3470), .C(n2672), .YC(n2654), .YS(n2655) );
  FAX1 U512 ( .A(n2659), .B(n3440), .C(n2674), .YC(n2656), .YS(n2657) );
  FAX1 U513 ( .A(n2661), .B(n3413), .C(n2676), .YC(n2658), .YS(n2659) );
  FAX1 U514 ( .A(n2663), .B(n3389), .C(n2678), .YC(n2660), .YS(n2661) );
  FAX1 U515 ( .A(n3350), .B(n3368), .C(n2680), .YC(n2662), .YS(n2663) );
  FAX1 U516 ( .A(n2667), .B(n3599), .C(n2682), .YC(n2664), .YS(n2665) );
  FAX1 U517 ( .A(n2669), .B(n3567), .C(n2684), .YC(n2666), .YS(n2667) );
  FAX1 U518 ( .A(n2671), .B(n3535), .C(n2686), .YC(n2668), .YS(n2669) );
  FAX1 U519 ( .A(n2673), .B(n3503), .C(n2688), .YC(n2670), .YS(n2671) );
  FAX1 U520 ( .A(n2675), .B(n3471), .C(n2690), .YC(n2672), .YS(n2673) );
  FAX1 U521 ( .A(n2677), .B(n3441), .C(n2692), .YC(n2674), .YS(n2675) );
  FAX1 U522 ( .A(n2679), .B(n3414), .C(n2694), .YC(n2676), .YS(n2677) );
  FAX1 U523 ( .A(n2681), .B(n3390), .C(n2696), .YC(n2678), .YS(n2679) );
  FAX1 U524 ( .A(n3351), .B(n3369), .C(n2698), .YC(n2680), .YS(n2681) );
  FAX1 U525 ( .A(n2685), .B(n3600), .C(n2700), .YC(n2682), .YS(n2683) );
  FAX1 U526 ( .A(n2687), .B(n3568), .C(n2702), .YC(n2684), .YS(n2685) );
  FAX1 U527 ( .A(n2689), .B(n3536), .C(n2704), .YC(n2686), .YS(n2687) );
  FAX1 U528 ( .A(n2691), .B(n3504), .C(n2706), .YC(n2688), .YS(n2689) );
  FAX1 U529 ( .A(n2693), .B(n3472), .C(n2708), .YC(n2690), .YS(n2691) );
  FAX1 U530 ( .A(n2695), .B(n3442), .C(n2710), .YC(n2692), .YS(n2693) );
  FAX1 U531 ( .A(n2697), .B(n3415), .C(n2712), .YC(n2694), .YS(n2695) );
  FAX1 U532 ( .A(n2699), .B(n3391), .C(n2714), .YC(n2696), .YS(n2697) );
  HAX1 U533 ( .A(n3370), .B(n2716), .YC(n2698), .YS(n2699) );
  FAX1 U534 ( .A(n2703), .B(n3601), .C(n2718), .YC(n2700), .YS(n2701) );
  FAX1 U535 ( .A(n2705), .B(n3569), .C(n2720), .YC(n2702), .YS(n2703) );
  FAX1 U536 ( .A(n2707), .B(n3537), .C(n2722), .YC(n2704), .YS(n2705) );
  FAX1 U537 ( .A(n2709), .B(n3505), .C(n2724), .YC(n2706), .YS(n2707) );
  FAX1 U538 ( .A(n2711), .B(n3473), .C(n2726), .YC(n2708), .YS(n2709) );
  FAX1 U539 ( .A(n2713), .B(n3443), .C(n2728), .YC(n2710), .YS(n2711) );
  FAX1 U540 ( .A(n2715), .B(n3416), .C(n2730), .YC(n2712), .YS(n2713) );
  FAX1 U541 ( .A(n3392), .B(n2717), .C(n2732), .YC(n2714), .YS(n2715) );
  HAX1 U542 ( .A(n2734), .B(n3371), .YC(n2716), .YS(n2717) );
  FAX1 U543 ( .A(n2721), .B(n3602), .C(n2736), .YC(n2718), .YS(n2719) );
  FAX1 U544 ( .A(n2723), .B(n3570), .C(n2738), .YC(n2720), .YS(n2721) );
  FAX1 U545 ( .A(n2725), .B(n3538), .C(n2740), .YC(n2722), .YS(n2723) );
  FAX1 U546 ( .A(n2727), .B(n3506), .C(n2742), .YC(n2724), .YS(n2725) );
  FAX1 U547 ( .A(n2729), .B(n3474), .C(n2744), .YC(n2726), .YS(n2727) );
  FAX1 U548 ( .A(n2731), .B(n3444), .C(n2746), .YC(n2728), .YS(n2729) );
  FAX1 U549 ( .A(n2733), .B(n3417), .C(n2748), .YC(n2730), .YS(n2731) );
  FAX1 U550 ( .A(n2735), .B(n3393), .C(n2750), .YC(n2732), .YS(n2733) );
  HAX1 U551 ( .A(n2159), .B(n3372), .YC(n2734), .YS(n2735) );
  FAX1 U552 ( .A(n2739), .B(n3603), .C(n2752), .YC(n2736), .YS(n2737) );
  FAX1 U553 ( .A(n2741), .B(n3571), .C(n2754), .YC(n2738), .YS(n2739) );
  FAX1 U554 ( .A(n2743), .B(n3539), .C(n2756), .YC(n2740), .YS(n2741) );
  FAX1 U555 ( .A(n2745), .B(n3507), .C(n2758), .YC(n2742), .YS(n2743) );
  FAX1 U556 ( .A(n2747), .B(n3475), .C(n2760), .YC(n2744), .YS(n2745) );
  FAX1 U557 ( .A(n2749), .B(n3445), .C(n2762), .YC(n2746), .YS(n2747) );
  FAX1 U558 ( .A(n2751), .B(n3418), .C(n2764), .YC(n2748), .YS(n2749) );
  HAX1 U559 ( .A(n3394), .B(n2766), .YC(n2750), .YS(n2751) );
  FAX1 U560 ( .A(n2755), .B(n3604), .C(n2768), .YC(n2752), .YS(n2753) );
  FAX1 U561 ( .A(n2757), .B(n3572), .C(n2770), .YC(n2754), .YS(n2755) );
  FAX1 U562 ( .A(n2759), .B(n3540), .C(n2772), .YC(n2756), .YS(n2757) );
  FAX1 U563 ( .A(n2761), .B(n3508), .C(n2774), .YC(n2758), .YS(n2759) );
  FAX1 U564 ( .A(n2763), .B(n3476), .C(n2776), .YC(n2760), .YS(n2761) );
  FAX1 U565 ( .A(n2765), .B(n3446), .C(n2778), .YC(n2762), .YS(n2763) );
  FAX1 U566 ( .A(n3419), .B(n2767), .C(n2780), .YC(n2764), .YS(n2765) );
  HAX1 U567 ( .A(n2782), .B(n3395), .YC(n2766), .YS(n2767) );
  FAX1 U568 ( .A(n2771), .B(n3605), .C(n2784), .YC(n2768), .YS(n2769) );
  FAX1 U569 ( .A(n2773), .B(n3573), .C(n2786), .YC(n2770), .YS(n2771) );
  FAX1 U570 ( .A(n2775), .B(n3541), .C(n2788), .YC(n2772), .YS(n2773) );
  FAX1 U571 ( .A(n2777), .B(n3509), .C(n2790), .YC(n2774), .YS(n2775) );
  FAX1 U572 ( .A(n2779), .B(n3477), .C(n2792), .YC(n2776), .YS(n2777) );
  FAX1 U573 ( .A(n2781), .B(n3447), .C(n2794), .YC(n2778), .YS(n2779) );
  FAX1 U574 ( .A(n2783), .B(n3420), .C(n2796), .YC(n2780), .YS(n2781) );
  HAX1 U575 ( .A(n2156), .B(n3396), .YC(n2782), .YS(n2783) );
  FAX1 U576 ( .A(n2787), .B(n3606), .C(n2798), .YC(n2784), .YS(n2785) );
  FAX1 U577 ( .A(n2789), .B(n3574), .C(n2800), .YC(n2786), .YS(n2787) );
  FAX1 U578 ( .A(n2791), .B(n3542), .C(n2802), .YC(n2788), .YS(n2789) );
  FAX1 U579 ( .A(n2793), .B(n3510), .C(n2804), .YC(n2790), .YS(n2791) );
  FAX1 U580 ( .A(n2795), .B(n3478), .C(n2806), .YC(n2792), .YS(n2793) );
  FAX1 U581 ( .A(n2797), .B(n3448), .C(n2808), .YC(n2794), .YS(n2795) );
  HAX1 U582 ( .A(n3421), .B(n2810), .YC(n2796), .YS(n2797) );
  FAX1 U583 ( .A(n2801), .B(n3607), .C(n2812), .YC(n2798), .YS(n2799) );
  FAX1 U584 ( .A(n2803), .B(n3575), .C(n2814), .YC(n2800), .YS(n2801) );
  FAX1 U585 ( .A(n2805), .B(n3543), .C(n2816), .YC(n2802), .YS(n2803) );
  FAX1 U586 ( .A(n2807), .B(n3511), .C(n2818), .YC(n2804), .YS(n2805) );
  FAX1 U587 ( .A(n2809), .B(n3479), .C(n2820), .YC(n2806), .YS(n2807) );
  FAX1 U588 ( .A(n3449), .B(n2811), .C(n2822), .YC(n2808), .YS(n2809) );
  HAX1 U589 ( .A(n2824), .B(n3422), .YC(n2810), .YS(n2811) );
  FAX1 U590 ( .A(n2815), .B(n3608), .C(n2826), .YC(n2812), .YS(n2813) );
  FAX1 U591 ( .A(n2817), .B(n3576), .C(n2828), .YC(n2814), .YS(n2815) );
  FAX1 U592 ( .A(n2819), .B(n3544), .C(n2830), .YC(n2816), .YS(n2817) );
  FAX1 U593 ( .A(n2821), .B(n3512), .C(n2832), .YC(n2818), .YS(n2819) );
  FAX1 U594 ( .A(n2823), .B(n3480), .C(n2834), .YC(n2820), .YS(n2821) );
  FAX1 U595 ( .A(n2825), .B(n3450), .C(n2836), .YC(n2822), .YS(n2823) );
  HAX1 U596 ( .A(n2153), .B(n3423), .YC(n2824), .YS(n2825) );
  FAX1 U597 ( .A(n2829), .B(n3609), .C(n2838), .YC(n2826), .YS(n2827) );
  FAX1 U598 ( .A(n2831), .B(n3577), .C(n2840), .YC(n2828), .YS(n2829) );
  FAX1 U599 ( .A(n2833), .B(n3545), .C(n2842), .YC(n2830), .YS(n2831) );
  FAX1 U600 ( .A(n2835), .B(n3513), .C(n2844), .YC(n2832), .YS(n2833) );
  FAX1 U601 ( .A(n2837), .B(n3481), .C(n2846), .YC(n2834), .YS(n2835) );
  HAX1 U602 ( .A(n3451), .B(n2848), .YC(n2836), .YS(n2837) );
  FAX1 U603 ( .A(n2841), .B(n3610), .C(n2850), .YC(n2838), .YS(n2839) );
  FAX1 U604 ( .A(n2843), .B(n3578), .C(n2852), .YC(n2840), .YS(n2841) );
  FAX1 U605 ( .A(n2845), .B(n3546), .C(n2854), .YC(n2842), .YS(n2843) );
  FAX1 U606 ( .A(n2847), .B(n3514), .C(n2856), .YC(n2844), .YS(n2845) );
  FAX1 U607 ( .A(n3482), .B(n2849), .C(n2858), .YC(n2846), .YS(n2847) );
  HAX1 U608 ( .A(n2860), .B(n3452), .YC(n2848), .YS(n2849) );
  FAX1 U609 ( .A(n2853), .B(n3611), .C(n2862), .YC(n2850), .YS(n2851) );
  FAX1 U610 ( .A(n2855), .B(n3579), .C(n2864), .YC(n2852), .YS(n2853) );
  FAX1 U611 ( .A(n2857), .B(n3547), .C(n2866), .YC(n2854), .YS(n2855) );
  FAX1 U612 ( .A(n2859), .B(n3515), .C(n2868), .YC(n2856), .YS(n2857) );
  FAX1 U613 ( .A(n2861), .B(n3483), .C(n2870), .YC(n2858), .YS(n2859) );
  HAX1 U614 ( .A(n4639), .B(n3453), .YC(n2860), .YS(n2861) );
  FAX1 U615 ( .A(n2865), .B(n3612), .C(n2872), .YC(n2862), .YS(n2863) );
  FAX1 U616 ( .A(n2867), .B(n3580), .C(n2874), .YC(n2864), .YS(n2865) );
  FAX1 U617 ( .A(n2869), .B(n3548), .C(n2876), .YC(n2866), .YS(n2867) );
  FAX1 U618 ( .A(n2871), .B(n3516), .C(n2878), .YC(n2868), .YS(n2869) );
  HAX1 U619 ( .A(n3484), .B(n2880), .YC(n2870), .YS(n2871) );
  FAX1 U620 ( .A(n2875), .B(n3613), .C(n2882), .YC(n2872), .YS(n2873) );
  FAX1 U621 ( .A(n2877), .B(n3581), .C(n2884), .YC(n2874), .YS(n2875) );
  FAX1 U622 ( .A(n2879), .B(n3549), .C(n2886), .YC(n2876), .YS(n2877) );
  FAX1 U623 ( .A(n3517), .B(n2881), .C(n2888), .YC(n2878), .YS(n2879) );
  HAX1 U624 ( .A(n2890), .B(n3485), .YC(n2880), .YS(n2881) );
  FAX1 U625 ( .A(n2885), .B(n3614), .C(n2892), .YC(n2882), .YS(n2883) );
  FAX1 U626 ( .A(n2887), .B(n3582), .C(n2894), .YC(n2884), .YS(n2885) );
  FAX1 U627 ( .A(n2889), .B(n3550), .C(n2896), .YC(n2886), .YS(n2887) );
  FAX1 U628 ( .A(n2891), .B(n3518), .C(n2898), .YC(n2888), .YS(n2889) );
  HAX1 U629 ( .A(n2147), .B(n3486), .YC(n2890), .YS(n2891) );
  FAX1 U630 ( .A(n2895), .B(n3615), .C(n2900), .YC(n2892), .YS(n2893) );
  FAX1 U631 ( .A(n2897), .B(n3583), .C(n2902), .YC(n2894), .YS(n2895) );
  FAX1 U632 ( .A(n2899), .B(n3551), .C(n2904), .YC(n2896), .YS(n2897) );
  HAX1 U633 ( .A(n3519), .B(n2906), .YC(n2898), .YS(n2899) );
  FAX1 U634 ( .A(n2903), .B(n3616), .C(n2908), .YC(n2900), .YS(n2901) );
  FAX1 U635 ( .A(n2905), .B(n3584), .C(n2910), .YC(n2902), .YS(n2903) );
  FAX1 U636 ( .A(n3552), .B(n2907), .C(n2912), .YC(n2904), .YS(n2905) );
  HAX1 U637 ( .A(n2914), .B(n3520), .YC(n2906), .YS(n2907) );
  FAX1 U638 ( .A(n2911), .B(n3617), .C(n2916), .YC(n2908), .YS(n2909) );
  FAX1 U639 ( .A(n2913), .B(n3585), .C(n2918), .YC(n2910), .YS(n2911) );
  FAX1 U640 ( .A(n2915), .B(n3553), .C(n2920), .YC(n2912), .YS(n2913) );
  HAX1 U641 ( .A(n2144), .B(n3521), .YC(n2914), .YS(n2915) );
  FAX1 U642 ( .A(n2919), .B(n3618), .C(n2922), .YC(n2916), .YS(n2917) );
  FAX1 U643 ( .A(n2921), .B(n3586), .C(n2924), .YC(n2918), .YS(n2919) );
  HAX1 U644 ( .A(n3554), .B(n2926), .YC(n2920), .YS(n2921) );
  FAX1 U645 ( .A(n2925), .B(n3619), .C(n2928), .YC(n2922), .YS(n2923) );
  FAX1 U646 ( .A(n3587), .B(n2927), .C(n2930), .YC(n2924), .YS(n2925) );
  HAX1 U647 ( .A(n2932), .B(n3555), .YC(n2926), .YS(n2927) );
  FAX1 U648 ( .A(n2931), .B(n3620), .C(n2934), .YC(n2928), .YS(n2929) );
  FAX1 U649 ( .A(n2933), .B(n3588), .C(n2936), .YC(n2930), .YS(n2931) );
  HAX1 U650 ( .A(n2141), .B(n3556), .YC(n2932), .YS(n2933) );
  FAX1 U651 ( .A(n2937), .B(n3621), .C(n2938), .YC(n2934), .YS(n2935) );
  HAX1 U652 ( .A(n3589), .B(n2940), .YC(n2936), .YS(n2937) );
  FAX1 U653 ( .A(n3622), .B(n2941), .C(n2942), .YC(n2938), .YS(n2939) );
  HAX1 U654 ( .A(n2944), .B(n3590), .YC(n2940), .YS(n2941) );
  FAX1 U655 ( .A(n2945), .B(n3623), .C(n2946), .YC(n2942), .YS(n2943) );
  HAX1 U656 ( .A(n2138), .B(n3591), .YC(n2944), .YS(n2945) );
  HAX1 U657 ( .A(n3624), .B(n2948), .YC(n2946), .YS(n2947) );
  HAX1 U658 ( .A(n2950), .B(n3625), .YC(n2948), .YS(n2949) );
  HAX1 U659 ( .A(n2135), .B(n3626), .YC(n2950), .YS(n2951) );
  HAX1 U1990 ( .A(n4631), .B(n3270), .YC(n3301), .YS(n3302) );
  FAX1 U1991 ( .A(n4630), .B(b[30]), .C(n3271), .YC(n3270), .YS(n3303) );
  FAX1 U1992 ( .A(b[30]), .B(b[29]), .C(n3272), .YC(n3271), .YS(n3304) );
  FAX1 U1993 ( .A(b[29]), .B(b[28]), .C(n3273), .YC(n3272), .YS(n3305) );
  FAX1 U1994 ( .A(b[28]), .B(n4642), .C(n3274), .YC(n3273), .YS(n3306) );
  FAX1 U1995 ( .A(n4643), .B(b[26]), .C(n3275), .YC(n3274), .YS(n3307) );
  FAX1 U1996 ( .A(b[26]), .B(n4645), .C(n3276), .YC(n3275), .YS(n3308) );
  FAX1 U1997 ( .A(n4646), .B(n4591), .C(n3277), .YC(n3276), .YS(n3309) );
  FAX1 U1998 ( .A(n4591), .B(n4648), .C(n3278), .YC(n3277), .YS(n3310) );
  FAX1 U1999 ( .A(n4649), .B(n4589), .C(n3279), .YC(n3278), .YS(n3311) );
  FAX1 U2000 ( .A(n4589), .B(n4652), .C(n3280), .YC(n3279), .YS(n3312) );
  FAX1 U2001 ( .A(n4652), .B(n4587), .C(n3281), .YC(n3280), .YS(n3313) );
  FAX1 U2002 ( .A(n4587), .B(n4655), .C(n3282), .YC(n3281), .YS(n3314) );
  FAX1 U2003 ( .A(n4655), .B(n4585), .C(n3283), .YC(n3282), .YS(n3315) );
  FAX1 U2004 ( .A(n4585), .B(n4659), .C(n3284), .YC(n3283), .YS(n3316) );
  FAX1 U2005 ( .A(n4658), .B(n4583), .C(n3285), .YC(n3284), .YS(n3317) );
  FAX1 U2006 ( .A(n4583), .B(n4663), .C(n3286), .YC(n3285), .YS(n3318) );
  FAX1 U2007 ( .A(n4665), .B(n4581), .C(n3287), .YC(n3286), .YS(n3319) );
  FAX1 U2008 ( .A(n4581), .B(n4668), .C(n3288), .YC(n3287), .YS(n3320) );
  FAX1 U2009 ( .A(n4667), .B(n4579), .C(n3289), .YC(n3288), .YS(n3321) );
  FAX1 U2010 ( .A(n4579), .B(n4673), .C(n3290), .YC(n3289), .YS(n3322) );
  FAX1 U2011 ( .A(n4672), .B(n4577), .C(n3291), .YC(n3290), .YS(n3323) );
  FAX1 U2012 ( .A(n4577), .B(n4677), .C(n3292), .YC(n3291), .YS(n3324) );
  FAX1 U2013 ( .A(n4679), .B(n4575), .C(n3293), .YC(n3292), .YS(n3325) );
  FAX1 U2014 ( .A(n4575), .B(n4682), .C(n3294), .YC(n3293), .YS(n3326) );
  FAX1 U2015 ( .A(n4681), .B(n4573), .C(n3295), .YC(n3294), .YS(n3327) );
  FAX1 U2016 ( .A(n4573), .B(n4686), .C(n3296), .YC(n3295), .YS(n3328) );
  FAX1 U2017 ( .A(n4688), .B(n4571), .C(n3297), .YC(n3296), .YS(n3329) );
  FAX1 U2018 ( .A(n4571), .B(n4690), .C(n3298), .YC(n3297), .YS(n3330) );
  FAX1 U2019 ( .A(n4692), .B(n4569), .C(n3299), .YC(n3298), .YS(n3331) );
  FAX1 U2020 ( .A(n4569), .B(n4694), .C(n3300), .YC(n3299), .YS(n3332) );
  HAX1 U2021 ( .A(n4694), .B(n4696), .YC(n3300), .YS(n3333) );
  OR2X2 U2024 ( .A(n4892), .B(n4764), .Y(n4552) );
  OR2X2 U2025 ( .A(n4755), .B(n5404), .Y(n4553) );
  NAND2X1 U2026 ( .A(n5577), .B(n5575), .Y(n4554) );
  NAND2X1 U2027 ( .A(n4749), .B(n5711), .Y(n4555) );
  NAND2X1 U2028 ( .A(n4752), .B(n5648), .Y(n4556) );
  NAND2X1 U2029 ( .A(a[31]), .B(n4745), .Y(n4557) );
  INVX2 U2030 ( .A(n5410), .Y(n4595) );
  INVX2 U2031 ( .A(n5500), .Y(n4592) );
  INVX2 U2032 ( .A(n5411), .Y(n4597) );
  INVX2 U2033 ( .A(n4901), .Y(n4617) );
  INVX2 U2034 ( .A(n5004), .Y(n4613) );
  INVX2 U2035 ( .A(n5107), .Y(n4609) );
  INVX2 U2036 ( .A(n5210), .Y(n4605) );
  INVX2 U2037 ( .A(n5501), .Y(n4594) );
  INVX2 U2038 ( .A(n4998), .Y(n4614) );
  INVX2 U2039 ( .A(n5101), .Y(n4610) );
  INVX2 U2040 ( .A(n5204), .Y(n4606) );
  INVX2 U2041 ( .A(n5307), .Y(n4601) );
  INVX2 U2042 ( .A(n4902), .Y(n4615) );
  INVX2 U2043 ( .A(n5005), .Y(n4611) );
  INVX2 U2044 ( .A(n5108), .Y(n4607) );
  INVX2 U2045 ( .A(n5211), .Y(n4602) );
  INVX2 U2046 ( .A(n5653), .Y(n4746) );
  INVX2 U2047 ( .A(n5654), .Y(n4748) );
  INVX2 U2048 ( .A(n5581), .Y(n4750) );
  INVX2 U2049 ( .A(n4560), .Y(n4627) );
  INVX2 U2050 ( .A(n4561), .Y(n4628) );
  INVX2 U2051 ( .A(n4562), .Y(n4629) );
  INVX2 U2052 ( .A(n4558), .Y(n4621) );
  INVX2 U2053 ( .A(n4559), .Y(n4622) );
  INVX2 U2054 ( .A(n5574), .Y(n4593) );
  INVX2 U2055 ( .A(n5646), .Y(n4567) );
  INVX2 U2056 ( .A(n5582), .Y(n4751) );
  INVX2 U2057 ( .A(n5714), .Y(n4743) );
  INVX2 U2058 ( .A(n5715), .Y(n4744) );
  INVX2 U2059 ( .A(n3332), .Y(n4738) );
  INVX2 U2060 ( .A(n3329), .Y(n4735) );
  INVX2 U2061 ( .A(n3333), .Y(n4741) );
  INVX2 U2062 ( .A(n4563), .Y(n4625) );
  INVX2 U2063 ( .A(n4564), .Y(n4626) );
  INVX2 U2064 ( .A(n4896), .Y(n4618) );
  INVX2 U2065 ( .A(n5403), .Y(n4598) );
  INVX2 U2066 ( .A(n5493), .Y(n4596) );
  INVX2 U2067 ( .A(n4631), .Y(n4632) );
  INVX2 U2068 ( .A(n5709), .Y(n4747) );
  AND2X1 U2069 ( .A(n4755), .B(n5405), .Y(n4558) );
  INVX2 U2070 ( .A(n2132), .Y(n4620) );
  INVX2 U2071 ( .A(n2141), .Y(n4608) );
  INVX2 U2072 ( .A(n2144), .Y(n4604) );
  INVX2 U2073 ( .A(n2147), .Y(n4600) );
  AND2X1 U2074 ( .A(n4754), .B(n5495), .Y(n4559) );
  AND2X1 U2075 ( .A(n4758), .B(n5199), .Y(n4560) );
  AND2X1 U2076 ( .A(n4756), .B(n5302), .Y(n4561) );
  NOR2X1 U2077 ( .A(n5405), .B(n5406), .Y(n4562) );
  INVX2 U2078 ( .A(n2132), .Y(n4619) );
  INVX2 U2079 ( .A(n2144), .Y(n4603) );
  AND2X1 U2080 ( .A(n4762), .B(n4993), .Y(n4563) );
  INVX2 U2081 ( .A(n2135), .Y(n4616) );
  INVX2 U2082 ( .A(n5746), .Y(n4742) );
  INVX2 U2083 ( .A(n2138), .Y(n4612) );
  INVX2 U2084 ( .A(n2147), .Y(n4599) );
  INVX2 U2085 ( .A(n3324), .Y(n4729) );
  INVX2 U2086 ( .A(n3326), .Y(n4731) );
  INVX2 U2087 ( .A(n3320), .Y(n4724) );
  INVX2 U2088 ( .A(n3318), .Y(n4721) );
  INVX2 U2089 ( .A(n3322), .Y(n4726) );
  INVX2 U2090 ( .A(n3327), .Y(n4733) );
  INVX2 U2091 ( .A(n3331), .Y(n4737) );
  INVX2 U2092 ( .A(n3325), .Y(n4730) );
  INVX2 U2093 ( .A(n3321), .Y(n4725) );
  INVX2 U2094 ( .A(n3323), .Y(n4727) );
  INVX2 U2095 ( .A(n3319), .Y(n4722) );
  INVX2 U2096 ( .A(n3328), .Y(n4734) );
  INVX2 U2097 ( .A(n3330), .Y(n4736) );
  INVX2 U2098 ( .A(n3317), .Y(n4720) );
  INVX2 U2099 ( .A(n3316), .Y(n4719) );
  INVX2 U2100 ( .A(n3315), .Y(n4718) );
  INVX2 U2101 ( .A(n3314), .Y(n4717) );
  INVX2 U2102 ( .A(n3313), .Y(n4716) );
  INVX2 U2103 ( .A(n3312), .Y(n4715) );
  INVX2 U2104 ( .A(n3311), .Y(n4714) );
  AND2X1 U2105 ( .A(n4760), .B(n5096), .Y(n4564) );
  INVX2 U2106 ( .A(n4565), .Y(n4624) );
  INVX2 U2107 ( .A(n4696), .Y(n4700) );
  INVX2 U2108 ( .A(n4686), .Y(n4689) );
  BUFX2 U2109 ( .A(b[31]), .Y(n4630) );
  BUFX2 U2110 ( .A(b[31]), .Y(n4631) );
  INVX2 U2111 ( .A(n4638), .Y(n4637) );
  INVX2 U2112 ( .A(n4636), .Y(n4635) );
  INVX2 U2113 ( .A(n4634), .Y(n4633) );
  INVX2 U2114 ( .A(n4566), .Y(n4623) );
  INVX2 U2115 ( .A(n4695), .Y(n4694) );
  INVX2 U2116 ( .A(n4570), .Y(n4571) );
  INVX2 U2117 ( .A(n4640), .Y(n4639) );
  BUFX2 U2118 ( .A(b[0]), .Y(n4698) );
  BUFX2 U2119 ( .A(b[0]), .Y(n4696) );
  AND2X1 U2120 ( .A(a[1]), .B(n4764), .Y(n4565) );
  BUFX2 U2121 ( .A(b[0]), .Y(n4697) );
  INVX2 U2122 ( .A(n4690), .Y(n4693) );
  INVX2 U2123 ( .A(n4568), .Y(n4569) );
  INVX1 U2124 ( .A(b[2]), .Y(n4568) );
  INVX2 U2125 ( .A(n4574), .Y(n4575) );
  INVX2 U2126 ( .A(n4677), .Y(n4680) );
  INVX2 U2127 ( .A(n4682), .Y(n4685) );
  BUFX2 U2128 ( .A(b[5]), .Y(n4686) );
  BUFX2 U2129 ( .A(b[0]), .Y(n4699) );
  BUFX2 U2130 ( .A(b[5]), .Y(n4688) );
  BUFX2 U2131 ( .A(b[5]), .Y(n4687) );
  INVX2 U2132 ( .A(n4673), .Y(n4676) );
  INVX2 U2133 ( .A(n4668), .Y(n4671) );
  INVX2 U2134 ( .A(n4580), .Y(n4581) );
  INVX1 U2135 ( .A(b[14]), .Y(n4580) );
  INVX2 U2136 ( .A(b[19]), .Y(n4657) );
  INVX2 U2137 ( .A(n4663), .Y(n4666) );
  INVX2 U2138 ( .A(n4659), .Y(n4662) );
  INVX2 U2139 ( .A(n4651), .Y(n4654) );
  INVX2 U2140 ( .A(n4648), .Y(n4650) );
  INVX2 U2141 ( .A(n4645), .Y(n4647) );
  INVX2 U2142 ( .A(n4642), .Y(n4644) );
  INVX2 U2143 ( .A(n2150), .Y(n4640) );
  INVX2 U2144 ( .A(n2153), .Y(n4638) );
  AND2X1 U2145 ( .A(a[0]), .B(n4892), .Y(n4566) );
  INVX2 U2146 ( .A(n2156), .Y(n4636) );
  INVX2 U2147 ( .A(n2159), .Y(n4634) );
  BUFX2 U2148 ( .A(b[3]), .Y(n4690) );
  INVX1 U2149 ( .A(b[1]), .Y(n4695) );
  INVX2 U2150 ( .A(n4572), .Y(n4573) );
  INVX2 U2151 ( .A(n4576), .Y(n4577) );
  BUFX2 U2152 ( .A(b[3]), .Y(n4691) );
  BUFX2 U2153 ( .A(b[3]), .Y(n4692) );
  INVX2 U2154 ( .A(n4578), .Y(n4579) );
  INVX2 U2155 ( .A(n4582), .Y(n4583) );
  INVX2 U2156 ( .A(n4586), .Y(n4587) );
  INVX2 U2157 ( .A(n4584), .Y(n4585) );
  INVX1 U2158 ( .A(b[18]), .Y(n4584) );
  INVX2 U2159 ( .A(n4590), .Y(n4591) );
  INVX2 U2160 ( .A(n4588), .Y(n4589) );
  INVX1 U2161 ( .A(b[22]), .Y(n4588) );
  BUFX2 U2162 ( .A(b[21]), .Y(n4651) );
  BUFX2 U2163 ( .A(b[23]), .Y(n4648) );
  BUFX2 U2164 ( .A(b[21]), .Y(n4653) );
  BUFX2 U2165 ( .A(b[21]), .Y(n4652) );
  BUFX2 U2166 ( .A(b[23]), .Y(n4649) );
  BUFX2 U2167 ( .A(b[25]), .Y(n4645) );
  BUFX2 U2168 ( .A(b[27]), .Y(n4642) );
  BUFX2 U2169 ( .A(b[25]), .Y(n4646) );
  INVX1 U2170 ( .A(b[29]), .Y(n4641) );
  INVX1 U2171 ( .A(b[30]), .Y(n4704) );
  BUFX2 U2172 ( .A(b[27]), .Y(n4643) );
  INVX1 U2173 ( .A(b[20]), .Y(n4586) );
  BUFX2 U2174 ( .A(b[17]), .Y(n4661) );
  BUFX2 U2175 ( .A(b[17]), .Y(n4660) );
  BUFX2 U2176 ( .A(b[17]), .Y(n4659) );
  BUFX2 U2177 ( .A(b[17]), .Y(n4658) );
  INVX1 U2178 ( .A(b[4]), .Y(n4570) );
  BUFX2 U2179 ( .A(b[7]), .Y(n4683) );
  BUFX2 U2180 ( .A(b[7]), .Y(n4684) );
  BUFX2 U2181 ( .A(b[7]), .Y(n4682) );
  BUFX2 U2182 ( .A(b[7]), .Y(n4681) );
  BUFX2 U2183 ( .A(b[11]), .Y(n4674) );
  BUFX2 U2184 ( .A(b[11]), .Y(n4675) );
  BUFX2 U2185 ( .A(b[11]), .Y(n4673) );
  BUFX2 U2186 ( .A(b[11]), .Y(n4672) );
  BUFX2 U2187 ( .A(b[13]), .Y(n4669) );
  BUFX2 U2188 ( .A(b[13]), .Y(n4670) );
  BUFX2 U2189 ( .A(b[13]), .Y(n4668) );
  BUFX2 U2190 ( .A(b[13]), .Y(n4667) );
  BUFX2 U2191 ( .A(b[9]), .Y(n4678) );
  BUFX2 U2192 ( .A(b[9]), .Y(n4679) );
  BUFX2 U2193 ( .A(b[9]), .Y(n4677) );
  BUFX2 U2194 ( .A(b[15]), .Y(n4665) );
  BUFX2 U2195 ( .A(b[15]), .Y(n4664) );
  BUFX2 U2196 ( .A(b[15]), .Y(n4663) );
  BUFX2 U2197 ( .A(b[19]), .Y(n4656) );
  BUFX2 U2198 ( .A(b[19]), .Y(n4655) );
  INVX1 U2199 ( .A(b[24]), .Y(n4590) );
  INVX1 U2200 ( .A(b[8]), .Y(n4574) );
  INVX1 U2201 ( .A(b[6]), .Y(n4572) );
  INVX1 U2202 ( .A(b[16]), .Y(n4582) );
  INVX1 U2203 ( .A(b[10]), .Y(n4576) );
  INVX1 U2204 ( .A(b[12]), .Y(n4578) );
  INVX1 U2205 ( .A(b[28]), .Y(n4707) );
  INVX1 U2206 ( .A(b[26]), .Y(n4710) );
  INVX2 U2207 ( .A(n3301), .Y(n4701) );
  INVX2 U2208 ( .A(n3302), .Y(n4702) );
  INVX2 U2209 ( .A(n3303), .Y(n4703) );
  INVX2 U2210 ( .A(n3304), .Y(n4705) );
  INVX2 U2211 ( .A(n3305), .Y(n4706) );
  INVX2 U2212 ( .A(n3306), .Y(n4708) );
  INVX2 U2213 ( .A(n3307), .Y(n4709) );
  INVX2 U2214 ( .A(n3308), .Y(n4711) );
  INVX2 U2215 ( .A(n3309), .Y(n4712) );
  INVX2 U2216 ( .A(n3310), .Y(n4713) );
  INVX2 U2217 ( .A(n2429), .Y(n4723) );
  INVX2 U2218 ( .A(n2472), .Y(n4728) );
  INVX2 U2219 ( .A(n2520), .Y(n4732) );
  INVX2 U2220 ( .A(n5312), .Y(n4739) );
  INVX2 U2221 ( .A(n4801), .Y(n4740) );
  INVX2 U2222 ( .A(n5747), .Y(n4745) );
  INVX2 U2223 ( .A(n5710), .Y(n4749) );
  INVX2 U2224 ( .A(n5647), .Y(n4752) );
  INVX2 U2225 ( .A(n5577), .Y(n4753) );
  INVX2 U2226 ( .A(n5494), .Y(n4754) );
  INVX2 U2227 ( .A(n5406), .Y(n4755) );
  INVX2 U2228 ( .A(n5303), .Y(n4756) );
  INVX2 U2229 ( .A(n2141), .Y(n4757) );
  INVX2 U2230 ( .A(n5200), .Y(n4758) );
  INVX2 U2231 ( .A(n2138), .Y(n4759) );
  INVX2 U2232 ( .A(n5097), .Y(n4760) );
  INVX2 U2233 ( .A(n2135), .Y(n4761) );
  INVX2 U2234 ( .A(n4994), .Y(n4762) );
  INVX2 U2235 ( .A(a[1]), .Y(n4763) );
  INVX2 U2236 ( .A(a[0]), .Y(n4764) );
  XOR2X1 U2237 ( .A(n4765), .B(n4766), .Y(product[47]) );
  XOR2X1 U2238 ( .A(n4767), .B(n4768), .Y(n4766) );
  XOR2X1 U2239 ( .A(n2405), .B(n2352), .Y(n4768) );
  XOR2X1 U2240 ( .A(n2409), .B(n2407), .Y(n4767) );
  XOR2X1 U2241 ( .A(n4769), .B(n4770), .Y(n4765) );
  XOR2X1 U2242 ( .A(n4637), .B(n4639), .Y(n4770) );
  XOR2X1 U2243 ( .A(n4771), .B(n4772), .Y(n4769) );
  XOR2X1 U2244 ( .A(n4773), .B(n4774), .Y(n4772) );
  XOR2X1 U2245 ( .A(n4775), .B(n4776), .Y(n4774) );
  XOR2X1 U2246 ( .A(n4777), .B(n4778), .Y(n4776) );
  XOR2X1 U2247 ( .A(n2411), .B(n2159), .Y(n4778) );
  XOR2X1 U2248 ( .A(n2415), .B(n2413), .Y(n4777) );
  XOR2X1 U2249 ( .A(n4779), .B(n4780), .Y(n4775) );
  XOR2X1 U2250 ( .A(n4781), .B(n4782), .Y(n4780) );
  OAI21X1 U2251 ( .A(n4557), .B(n4720), .C(n4783), .Y(n4782) );
  OAI22X1 U2252 ( .A(n4665), .B(n4784), .C(n4742), .D(n4784), .Y(n4783) );
  OAI22X1 U2253 ( .A(n4743), .B(n4662), .C(n4744), .D(n4582), .Y(n4784) );
  OAI21X1 U2254 ( .A(n4555), .B(n4717), .C(n4785), .Y(n4781) );
  OAI22X1 U2255 ( .A(n4585), .B(n4786), .C(n4747), .D(n4786), .Y(n4785) );
  OAI22X1 U2256 ( .A(n4746), .B(n4586), .C(n4748), .D(n4657), .Y(n4786) );
  XOR2X1 U2257 ( .A(n4787), .B(n2156), .Y(n4779) );
  OAI21X1 U2258 ( .A(n4556), .B(n4714), .C(n4788), .Y(n4787) );
  OAI22X1 U2259 ( .A(n4653), .B(n4789), .C(n4567), .D(n4789), .Y(n4788) );
  OAI22X1 U2260 ( .A(n4750), .B(n4650), .C(n4751), .D(n4588), .Y(n4789) );
  OAI21X1 U2261 ( .A(n4554), .B(n4711), .C(n4790), .Y(n4773) );
  OAI22X1 U2262 ( .A(n4591), .B(n4791), .C(n4593), .D(n4791), .Y(n4790) );
  OAI22X1 U2263 ( .A(n4592), .B(n4710), .C(n4594), .D(n4647), .Y(n4791) );
  XOR2X1 U2264 ( .A(n4792), .B(n4793), .Y(n4771) );
  XNOR2X1 U2265 ( .A(n2147), .B(n4794), .Y(n4793) );
  OAI21X1 U2266 ( .A(n4621), .B(n4702), .C(n4795), .Y(n4794) );
  OAI22X1 U2267 ( .A(b[30]), .B(n4796), .C(n4598), .D(n4796), .Y(n4795) );
  NOR2X1 U2268 ( .A(n4632), .B(n4553), .Y(n4796) );
  OAI21X1 U2269 ( .A(n4622), .B(n4706), .C(n4797), .Y(n4792) );
  OAI22X1 U2270 ( .A(n4643), .B(n4798), .C(n4596), .D(n4798), .Y(n4797) );
  OAI22X1 U2271 ( .A(n4595), .B(n4641), .C(n4597), .D(n4707), .Y(n4798) );
  XNOR2X1 U2272 ( .A(n4799), .B(n4619), .Y(n3661) );
  OAI22X1 U2273 ( .A(n4700), .B(n4552), .C(n4623), .D(n4700), .Y(n4799) );
  XNOR2X1 U2274 ( .A(n4800), .B(n4619), .Y(n3660) );
  OAI21X1 U2275 ( .A(n4623), .B(n4741), .C(n4740), .Y(n4800) );
  OAI22X1 U2276 ( .A(n4624), .B(n4700), .C(n4695), .D(n4552), .Y(n4801) );
  XNOR2X1 U2277 ( .A(n4802), .B(n4619), .Y(n3659) );
  OAI21X1 U2278 ( .A(n4623), .B(n4738), .C(n4803), .Y(n4802) );
  OAI22X1 U2279 ( .A(n4698), .B(n4804), .C(n4618), .D(n4804), .Y(n4803) );
  OAI22X1 U2280 ( .A(n4624), .B(n4695), .C(n4552), .D(n4568), .Y(n4804) );
  XNOR2X1 U2281 ( .A(n4805), .B(n4619), .Y(n3658) );
  OAI21X1 U2282 ( .A(n4623), .B(n4737), .C(n4806), .Y(n4805) );
  OAI22X1 U2283 ( .A(n4694), .B(n4807), .C(n4618), .D(n4807), .Y(n4806) );
  OAI22X1 U2284 ( .A(n4624), .B(n4568), .C(n4552), .D(n4693), .Y(n4807) );
  XNOR2X1 U2285 ( .A(n4808), .B(n4619), .Y(n3657) );
  OAI21X1 U2286 ( .A(n4623), .B(n4736), .C(n4809), .Y(n4808) );
  OAI22X1 U2287 ( .A(n4569), .B(n4810), .C(n4618), .D(n4810), .Y(n4809) );
  OAI22X1 U2288 ( .A(n4624), .B(n4693), .C(n4552), .D(n4570), .Y(n4810) );
  XNOR2X1 U2289 ( .A(n4811), .B(n4619), .Y(n3656) );
  OAI21X1 U2290 ( .A(n4623), .B(n4735), .C(n4812), .Y(n4811) );
  OAI22X1 U2291 ( .A(n4692), .B(n4813), .C(n4618), .D(n4813), .Y(n4812) );
  OAI22X1 U2292 ( .A(n4624), .B(n4570), .C(n4552), .D(n4689), .Y(n4813) );
  XNOR2X1 U2293 ( .A(n4814), .B(n4619), .Y(n3655) );
  OAI21X1 U2294 ( .A(n4623), .B(n4734), .C(n4815), .Y(n4814) );
  OAI22X1 U2295 ( .A(n4571), .B(n4816), .C(n4618), .D(n4816), .Y(n4815) );
  OAI22X1 U2296 ( .A(n4624), .B(n4689), .C(n4552), .D(n4572), .Y(n4816) );
  XNOR2X1 U2297 ( .A(n4817), .B(n4619), .Y(n3654) );
  OAI21X1 U2298 ( .A(n4623), .B(n4733), .C(n4818), .Y(n4817) );
  OAI22X1 U2299 ( .A(n4688), .B(n4819), .C(n4618), .D(n4819), .Y(n4818) );
  OAI22X1 U2300 ( .A(n4624), .B(n4572), .C(n4552), .D(n4685), .Y(n4819) );
  XNOR2X1 U2301 ( .A(n4820), .B(n4619), .Y(n3653) );
  OAI21X1 U2302 ( .A(n4623), .B(n4731), .C(n4821), .Y(n4820) );
  OAI22X1 U2303 ( .A(n4573), .B(n4822), .C(n4618), .D(n4822), .Y(n4821) );
  OAI22X1 U2304 ( .A(n4624), .B(n4685), .C(n4552), .D(n4574), .Y(n4822) );
  XNOR2X1 U2305 ( .A(n4823), .B(n4619), .Y(n3652) );
  OAI21X1 U2306 ( .A(n4623), .B(n4730), .C(n4824), .Y(n4823) );
  OAI22X1 U2307 ( .A(n4684), .B(n4825), .C(n4618), .D(n4825), .Y(n4824) );
  OAI22X1 U2308 ( .A(n4624), .B(n4574), .C(n4552), .D(n4680), .Y(n4825) );
  XNOR2X1 U2309 ( .A(n4826), .B(n4619), .Y(n3651) );
  OAI21X1 U2310 ( .A(n4623), .B(n4729), .C(n4827), .Y(n4826) );
  OAI22X1 U2311 ( .A(n4575), .B(n4828), .C(n4618), .D(n4828), .Y(n4827) );
  OAI22X1 U2312 ( .A(n4624), .B(n4680), .C(n4552), .D(n4576), .Y(n4828) );
  XNOR2X1 U2313 ( .A(n4829), .B(n4619), .Y(n3650) );
  OAI21X1 U2314 ( .A(n4623), .B(n4727), .C(n4830), .Y(n4829) );
  OAI22X1 U2315 ( .A(n4679), .B(n4831), .C(n4618), .D(n4831), .Y(n4830) );
  OAI22X1 U2316 ( .A(n4624), .B(n4576), .C(n4552), .D(n4676), .Y(n4831) );
  XNOR2X1 U2317 ( .A(n4832), .B(n4619), .Y(n3649) );
  OAI21X1 U2318 ( .A(n4623), .B(n4726), .C(n4833), .Y(n4832) );
  OAI22X1 U2319 ( .A(n4577), .B(n4834), .C(n4618), .D(n4834), .Y(n4833) );
  OAI22X1 U2320 ( .A(n4624), .B(n4676), .C(n4552), .D(n4578), .Y(n4834) );
  XNOR2X1 U2321 ( .A(n4835), .B(n4619), .Y(n3648) );
  OAI21X1 U2322 ( .A(n4623), .B(n4725), .C(n4836), .Y(n4835) );
  OAI22X1 U2323 ( .A(n4675), .B(n4837), .C(n4618), .D(n4837), .Y(n4836) );
  OAI22X1 U2324 ( .A(n4624), .B(n4578), .C(n4552), .D(n4671), .Y(n4837) );
  XNOR2X1 U2325 ( .A(n4838), .B(n4619), .Y(n3647) );
  OAI21X1 U2326 ( .A(n4623), .B(n4724), .C(n4839), .Y(n4838) );
  OAI22X1 U2327 ( .A(n4579), .B(n4840), .C(n4618), .D(n4840), .Y(n4839) );
  OAI22X1 U2328 ( .A(n4624), .B(n4671), .C(n4552), .D(n4580), .Y(n4840) );
  XNOR2X1 U2329 ( .A(n4841), .B(n4619), .Y(n3646) );
  OAI21X1 U2330 ( .A(n4623), .B(n4722), .C(n4842), .Y(n4841) );
  OAI22X1 U2331 ( .A(n4670), .B(n4843), .C(n4618), .D(n4843), .Y(n4842) );
  OAI22X1 U2332 ( .A(n4624), .B(n4580), .C(n4552), .D(n4666), .Y(n4843) );
  XNOR2X1 U2333 ( .A(n4844), .B(n4619), .Y(n3645) );
  OAI21X1 U2334 ( .A(n4623), .B(n4721), .C(n4845), .Y(n4844) );
  OAI22X1 U2335 ( .A(n4581), .B(n4846), .C(n4618), .D(n4846), .Y(n4845) );
  OAI22X1 U2336 ( .A(n4624), .B(n4666), .C(n4582), .D(n4552), .Y(n4846) );
  XNOR2X1 U2337 ( .A(n4847), .B(n4619), .Y(n3644) );
  OAI21X1 U2338 ( .A(n4720), .B(n4623), .C(n4848), .Y(n4847) );
  OAI22X1 U2339 ( .A(n4664), .B(n4849), .C(n4618), .D(n4849), .Y(n4848) );
  OAI22X1 U2340 ( .A(n4582), .B(n4624), .C(n4662), .D(n4552), .Y(n4849) );
  XNOR2X1 U2341 ( .A(n4850), .B(n4619), .Y(n3643) );
  OAI21X1 U2342 ( .A(n4623), .B(n4719), .C(n4851), .Y(n4850) );
  OAI22X1 U2343 ( .A(n4583), .B(n4852), .C(n4618), .D(n4852), .Y(n4851) );
  OAI22X1 U2344 ( .A(n4662), .B(n4624), .C(n4552), .D(n4584), .Y(n4852) );
  XNOR2X1 U2345 ( .A(n4853), .B(n4619), .Y(n3642) );
  OAI21X1 U2346 ( .A(n4623), .B(n4718), .C(n4854), .Y(n4853) );
  OAI22X1 U2347 ( .A(n4660), .B(n4855), .C(n4618), .D(n4855), .Y(n4854) );
  OAI22X1 U2348 ( .A(n4624), .B(n4584), .C(n4657), .D(n4552), .Y(n4855) );
  XNOR2X1 U2349 ( .A(n4856), .B(n4620), .Y(n3641) );
  OAI21X1 U2350 ( .A(n4717), .B(n4623), .C(n4857), .Y(n4856) );
  OAI22X1 U2351 ( .A(n4585), .B(n4858), .C(n4618), .D(n4858), .Y(n4857) );
  OAI22X1 U2352 ( .A(n4657), .B(n4624), .C(n4586), .D(n4552), .Y(n4858) );
  XNOR2X1 U2353 ( .A(n4859), .B(n4620), .Y(n3640) );
  OAI21X1 U2354 ( .A(n4623), .B(n4716), .C(n4860), .Y(n4859) );
  OAI22X1 U2355 ( .A(n4656), .B(n4861), .C(n4618), .D(n4861), .Y(n4860) );
  OAI22X1 U2356 ( .A(n4586), .B(n4624), .C(n4552), .D(n4654), .Y(n4861) );
  XNOR2X1 U2357 ( .A(n4862), .B(n4620), .Y(n3639) );
  OAI21X1 U2358 ( .A(n4623), .B(n4715), .C(n4863), .Y(n4862) );
  OAI22X1 U2359 ( .A(n4587), .B(n4864), .C(n4618), .D(n4864), .Y(n4863) );
  OAI22X1 U2360 ( .A(n4624), .B(n4654), .C(n4588), .D(n4552), .Y(n4864) );
  XNOR2X1 U2361 ( .A(n4865), .B(n4620), .Y(n3638) );
  OAI21X1 U2362 ( .A(n4714), .B(n4623), .C(n4866), .Y(n4865) );
  OAI22X1 U2363 ( .A(n4653), .B(n4867), .C(n4618), .D(n4867), .Y(n4866) );
  OAI22X1 U2364 ( .A(n4588), .B(n4624), .C(n4650), .D(n4552), .Y(n4867) );
  XNOR2X1 U2365 ( .A(n4868), .B(n4620), .Y(n3637) );
  OAI21X1 U2366 ( .A(n4623), .B(n4713), .C(n4869), .Y(n4868) );
  OAI22X1 U2367 ( .A(n4589), .B(n4870), .C(n4618), .D(n4870), .Y(n4869) );
  OAI22X1 U2368 ( .A(n4650), .B(n4624), .C(n4552), .D(n4590), .Y(n4870) );
  XNOR2X1 U2369 ( .A(n4871), .B(n4620), .Y(n3636) );
  OAI21X1 U2370 ( .A(n4623), .B(n4712), .C(n4872), .Y(n4871) );
  OAI22X1 U2371 ( .A(n4649), .B(n4873), .C(n4618), .D(n4873), .Y(n4872) );
  OAI22X1 U2372 ( .A(n4624), .B(n4590), .C(n4647), .D(n4552), .Y(n4873) );
  XNOR2X1 U2373 ( .A(n4874), .B(n4620), .Y(n3635) );
  OAI21X1 U2374 ( .A(n4711), .B(n4623), .C(n4875), .Y(n4874) );
  OAI22X1 U2375 ( .A(n4591), .B(n4876), .C(n4618), .D(n4876), .Y(n4875) );
  OAI22X1 U2376 ( .A(n4647), .B(n4624), .C(n4710), .D(n4552), .Y(n4876) );
  XNOR2X1 U2377 ( .A(n4877), .B(n4620), .Y(n3634) );
  OAI21X1 U2378 ( .A(n4623), .B(n4709), .C(n4878), .Y(n4877) );
  OAI22X1 U2379 ( .A(n4646), .B(n4879), .C(n4618), .D(n4879), .Y(n4878) );
  OAI22X1 U2380 ( .A(n4710), .B(n4624), .C(n4552), .D(n4644), .Y(n4879) );
  XNOR2X1 U2381 ( .A(n4880), .B(n4620), .Y(n3633) );
  OAI21X1 U2382 ( .A(n4623), .B(n4708), .C(n4881), .Y(n4880) );
  OAI22X1 U2383 ( .A(b[26]), .B(n4882), .C(n4618), .D(n4882), .Y(n4881) );
  OAI22X1 U2384 ( .A(n4624), .B(n4644), .C(n4707), .D(n4552), .Y(n4882) );
  XNOR2X1 U2385 ( .A(n4883), .B(n4620), .Y(n3632) );
  OAI21X1 U2386 ( .A(n4706), .B(n4623), .C(n4884), .Y(n4883) );
  OAI22X1 U2387 ( .A(n4643), .B(n4885), .C(n4618), .D(n4885), .Y(n4884) );
  OAI22X1 U2388 ( .A(n4707), .B(n4624), .C(n4641), .D(n4552), .Y(n4885) );
  XNOR2X1 U2389 ( .A(n4886), .B(n4620), .Y(n3631) );
  OAI21X1 U2390 ( .A(n4623), .B(n4705), .C(n4887), .Y(n4886) );
  OAI22X1 U2391 ( .A(b[28]), .B(n4888), .C(n4618), .D(n4888), .Y(n4887) );
  OAI22X1 U2392 ( .A(n4641), .B(n4624), .C(n4552), .D(n4704), .Y(n4888) );
  XNOR2X1 U2393 ( .A(n4889), .B(n4620), .Y(n3630) );
  OAI21X1 U2394 ( .A(n4623), .B(n4703), .C(n4890), .Y(n4889) );
  OAI22X1 U2395 ( .A(b[29]), .B(n4891), .C(n4618), .D(n4891), .Y(n4890) );
  OAI22X1 U2396 ( .A(n4624), .B(n4704), .C(n4632), .D(n4552), .Y(n4891) );
  XNOR2X1 U2397 ( .A(n4893), .B(n4620), .Y(n3629) );
  OAI21X1 U2398 ( .A(n4702), .B(n4623), .C(n4894), .Y(n4893) );
  OAI22X1 U2399 ( .A(b[30]), .B(n4895), .C(n4618), .D(n4895), .Y(n4894) );
  NOR2X1 U2400 ( .A(n4624), .B(n4632), .Y(n4895) );
  XNOR2X1 U2401 ( .A(n4897), .B(n4620), .Y(n3628) );
  OAI22X1 U2402 ( .A(n4632), .B(n4896), .C(n4623), .D(n4701), .Y(n4897) );
  NAND3X1 U2403 ( .A(n4892), .B(n4764), .C(n4763), .Y(n4896) );
  XNOR2X1 U2404 ( .A(a[1]), .B(n4620), .Y(n4892) );
  XNOR2X1 U2405 ( .A(n4898), .B(n4616), .Y(n3626) );
  OAI22X1 U2406 ( .A(n4700), .B(n4615), .C(n4700), .D(n4625), .Y(n4898) );
  XNOR2X1 U2407 ( .A(n4899), .B(n4761), .Y(n3625) );
  OAI21X1 U2408 ( .A(n4741), .B(n4625), .C(n4900), .Y(n4899) );
  AOI22X1 U2409 ( .A(n4901), .B(n4698), .C(n4902), .D(n4694), .Y(n4900) );
  XNOR2X1 U2410 ( .A(n4903), .B(n4761), .Y(n3624) );
  OAI21X1 U2411 ( .A(n4738), .B(n4625), .C(n4904), .Y(n4903) );
  OAI22X1 U2412 ( .A(n4698), .B(n4905), .C(n4614), .D(n4905), .Y(n4904) );
  OAI22X1 U2413 ( .A(n4695), .B(n4617), .C(n4568), .D(n4615), .Y(n4905) );
  XNOR2X1 U2414 ( .A(n4906), .B(n4761), .Y(n3623) );
  OAI21X1 U2415 ( .A(n4737), .B(n4625), .C(n4907), .Y(n4906) );
  OAI22X1 U2416 ( .A(n4694), .B(n4908), .C(n4614), .D(n4908), .Y(n4907) );
  OAI22X1 U2417 ( .A(n4568), .B(n4617), .C(n4693), .D(n4615), .Y(n4908) );
  XNOR2X1 U2418 ( .A(n4909), .B(n4761), .Y(n3622) );
  OAI21X1 U2419 ( .A(n4736), .B(n4625), .C(n4910), .Y(n4909) );
  OAI22X1 U2420 ( .A(n4569), .B(n4911), .C(n4614), .D(n4911), .Y(n4910) );
  OAI22X1 U2421 ( .A(n4693), .B(n4617), .C(n4570), .D(n4615), .Y(n4911) );
  XNOR2X1 U2422 ( .A(n4912), .B(n4761), .Y(n3621) );
  OAI21X1 U2423 ( .A(n4735), .B(n4625), .C(n4913), .Y(n4912) );
  OAI22X1 U2424 ( .A(n4691), .B(n4914), .C(n4614), .D(n4914), .Y(n4913) );
  OAI22X1 U2425 ( .A(n4570), .B(n4617), .C(n4689), .D(n4615), .Y(n4914) );
  XNOR2X1 U2426 ( .A(n4915), .B(n4761), .Y(n3620) );
  OAI21X1 U2427 ( .A(n4734), .B(n4625), .C(n4916), .Y(n4915) );
  OAI22X1 U2428 ( .A(n4571), .B(n4917), .C(n4614), .D(n4917), .Y(n4916) );
  OAI22X1 U2429 ( .A(n4689), .B(n4617), .C(n4572), .D(n4615), .Y(n4917) );
  XNOR2X1 U2430 ( .A(n4918), .B(n4761), .Y(n3619) );
  OAI21X1 U2431 ( .A(n4733), .B(n4625), .C(n4919), .Y(n4918) );
  OAI22X1 U2432 ( .A(n4687), .B(n4920), .C(n4614), .D(n4920), .Y(n4919) );
  OAI22X1 U2433 ( .A(n4572), .B(n4617), .C(n4685), .D(n4615), .Y(n4920) );
  XNOR2X1 U2434 ( .A(n4921), .B(n4761), .Y(n3618) );
  OAI21X1 U2435 ( .A(n4731), .B(n4625), .C(n4922), .Y(n4921) );
  OAI22X1 U2436 ( .A(n4573), .B(n4923), .C(n4614), .D(n4923), .Y(n4922) );
  OAI22X1 U2437 ( .A(n4685), .B(n4617), .C(n4574), .D(n4615), .Y(n4923) );
  XNOR2X1 U2438 ( .A(n4924), .B(n4761), .Y(n3617) );
  OAI21X1 U2439 ( .A(n4730), .B(n4625), .C(n4925), .Y(n4924) );
  OAI22X1 U2440 ( .A(n4683), .B(n4926), .C(n4614), .D(n4926), .Y(n4925) );
  OAI22X1 U2441 ( .A(n4574), .B(n4617), .C(n4680), .D(n4615), .Y(n4926) );
  XNOR2X1 U2442 ( .A(n4927), .B(n4761), .Y(n3616) );
  OAI21X1 U2443 ( .A(n4729), .B(n4625), .C(n4928), .Y(n4927) );
  OAI22X1 U2444 ( .A(n4575), .B(n4929), .C(n4614), .D(n4929), .Y(n4928) );
  OAI22X1 U2445 ( .A(n4680), .B(n4617), .C(n4576), .D(n4615), .Y(n4929) );
  XNOR2X1 U2446 ( .A(n4930), .B(n4761), .Y(n3615) );
  OAI21X1 U2447 ( .A(n4727), .B(n4625), .C(n4931), .Y(n4930) );
  OAI22X1 U2448 ( .A(n4678), .B(n4932), .C(n4614), .D(n4932), .Y(n4931) );
  OAI22X1 U2449 ( .A(n4576), .B(n4617), .C(n4676), .D(n4615), .Y(n4932) );
  XNOR2X1 U2450 ( .A(n4933), .B(n4761), .Y(n3614) );
  OAI21X1 U2451 ( .A(n4726), .B(n4625), .C(n4934), .Y(n4933) );
  OAI22X1 U2452 ( .A(n4577), .B(n4935), .C(n4614), .D(n4935), .Y(n4934) );
  OAI22X1 U2453 ( .A(n4676), .B(n4617), .C(n4578), .D(n4615), .Y(n4935) );
  XNOR2X1 U2454 ( .A(n4936), .B(n4761), .Y(n3613) );
  OAI21X1 U2455 ( .A(n4725), .B(n4625), .C(n4937), .Y(n4936) );
  OAI22X1 U2456 ( .A(n4674), .B(n4938), .C(n4614), .D(n4938), .Y(n4937) );
  OAI22X1 U2457 ( .A(n4578), .B(n4617), .C(n4671), .D(n4615), .Y(n4938) );
  XNOR2X1 U2458 ( .A(n4939), .B(n4761), .Y(n3612) );
  OAI21X1 U2459 ( .A(n4724), .B(n4625), .C(n4940), .Y(n4939) );
  OAI22X1 U2460 ( .A(n4579), .B(n4941), .C(n4614), .D(n4941), .Y(n4940) );
  OAI22X1 U2461 ( .A(n4671), .B(n4617), .C(n4580), .D(n4615), .Y(n4941) );
  XNOR2X1 U2462 ( .A(n4942), .B(n4761), .Y(n3611) );
  OAI21X1 U2463 ( .A(n4722), .B(n4625), .C(n4943), .Y(n4942) );
  OAI22X1 U2464 ( .A(n4669), .B(n4944), .C(n4614), .D(n4944), .Y(n4943) );
  OAI22X1 U2465 ( .A(n4580), .B(n4617), .C(n4666), .D(n4615), .Y(n4944) );
  XNOR2X1 U2466 ( .A(n4945), .B(n4761), .Y(n3610) );
  OAI21X1 U2467 ( .A(n4721), .B(n4625), .C(n4946), .Y(n4945) );
  OAI22X1 U2468 ( .A(n4581), .B(n4947), .C(n4614), .D(n4947), .Y(n4946) );
  OAI22X1 U2469 ( .A(n4666), .B(n4617), .C(n4582), .D(n4615), .Y(n4947) );
  XNOR2X1 U2470 ( .A(n4948), .B(n4761), .Y(n3609) );
  OAI21X1 U2471 ( .A(n4720), .B(n4625), .C(n4949), .Y(n4948) );
  OAI22X1 U2472 ( .A(n4664), .B(n4950), .C(n4614), .D(n4950), .Y(n4949) );
  OAI22X1 U2473 ( .A(n4582), .B(n4617), .C(n4662), .D(n4615), .Y(n4950) );
  XNOR2X1 U2474 ( .A(n4951), .B(n4761), .Y(n3608) );
  OAI21X1 U2475 ( .A(n4719), .B(n4625), .C(n4952), .Y(n4951) );
  OAI22X1 U2476 ( .A(n4583), .B(n4953), .C(n4614), .D(n4953), .Y(n4952) );
  OAI22X1 U2477 ( .A(n4662), .B(n4617), .C(n4584), .D(n4615), .Y(n4953) );
  XNOR2X1 U2478 ( .A(n4954), .B(n4616), .Y(n3607) );
  OAI21X1 U2479 ( .A(n4718), .B(n4625), .C(n4955), .Y(n4954) );
  OAI22X1 U2480 ( .A(n4660), .B(n4956), .C(n4614), .D(n4956), .Y(n4955) );
  OAI22X1 U2481 ( .A(n4584), .B(n4617), .C(n4657), .D(n4615), .Y(n4956) );
  XNOR2X1 U2482 ( .A(n4957), .B(n4616), .Y(n3606) );
  OAI21X1 U2483 ( .A(n4717), .B(n4625), .C(n4958), .Y(n4957) );
  OAI22X1 U2484 ( .A(n4585), .B(n4959), .C(n4614), .D(n4959), .Y(n4958) );
  OAI22X1 U2485 ( .A(n4657), .B(n4617), .C(n4586), .D(n4615), .Y(n4959) );
  XNOR2X1 U2486 ( .A(n4960), .B(n4616), .Y(n3605) );
  OAI21X1 U2487 ( .A(n4716), .B(n4625), .C(n4961), .Y(n4960) );
  OAI22X1 U2488 ( .A(n4656), .B(n4962), .C(n4614), .D(n4962), .Y(n4961) );
  OAI22X1 U2489 ( .A(n4586), .B(n4617), .C(n4654), .D(n4615), .Y(n4962) );
  XNOR2X1 U2490 ( .A(n4963), .B(n4616), .Y(n3604) );
  OAI21X1 U2491 ( .A(n4715), .B(n4625), .C(n4964), .Y(n4963) );
  OAI22X1 U2492 ( .A(n4587), .B(n4965), .C(n4614), .D(n4965), .Y(n4964) );
  OAI22X1 U2493 ( .A(n4654), .B(n4617), .C(n4588), .D(n4615), .Y(n4965) );
  XNOR2X1 U2494 ( .A(n4966), .B(n4616), .Y(n3603) );
  OAI21X1 U2495 ( .A(n4714), .B(n4625), .C(n4967), .Y(n4966) );
  OAI22X1 U2496 ( .A(n4653), .B(n4968), .C(n4614), .D(n4968), .Y(n4967) );
  OAI22X1 U2497 ( .A(n4588), .B(n4617), .C(n4650), .D(n4615), .Y(n4968) );
  XNOR2X1 U2498 ( .A(n4969), .B(n4616), .Y(n3602) );
  OAI21X1 U2499 ( .A(n4713), .B(n4625), .C(n4970), .Y(n4969) );
  OAI22X1 U2500 ( .A(n4589), .B(n4971), .C(n4614), .D(n4971), .Y(n4970) );
  OAI22X1 U2501 ( .A(n4650), .B(n4617), .C(n4590), .D(n4615), .Y(n4971) );
  XNOR2X1 U2502 ( .A(n4972), .B(n4616), .Y(n3601) );
  OAI21X1 U2503 ( .A(n4712), .B(n4625), .C(n4973), .Y(n4972) );
  OAI22X1 U2504 ( .A(n4649), .B(n4974), .C(n4614), .D(n4974), .Y(n4973) );
  OAI22X1 U2505 ( .A(n4590), .B(n4617), .C(n4647), .D(n4615), .Y(n4974) );
  XNOR2X1 U2506 ( .A(n4975), .B(n4616), .Y(n3600) );
  OAI21X1 U2507 ( .A(n4711), .B(n4625), .C(n4976), .Y(n4975) );
  OAI22X1 U2508 ( .A(n4591), .B(n4977), .C(n4614), .D(n4977), .Y(n4976) );
  OAI22X1 U2509 ( .A(n4647), .B(n4617), .C(n4710), .D(n4615), .Y(n4977) );
  XNOR2X1 U2510 ( .A(n4978), .B(n4616), .Y(n3599) );
  OAI21X1 U2511 ( .A(n4709), .B(n4625), .C(n4979), .Y(n4978) );
  OAI22X1 U2512 ( .A(n4646), .B(n4980), .C(n4614), .D(n4980), .Y(n4979) );
  OAI22X1 U2513 ( .A(n4710), .B(n4617), .C(n4644), .D(n4615), .Y(n4980) );
  XNOR2X1 U2514 ( .A(n4981), .B(n4616), .Y(n3598) );
  OAI21X1 U2515 ( .A(n4708), .B(n4625), .C(n4982), .Y(n4981) );
  OAI22X1 U2516 ( .A(b[26]), .B(n4983), .C(n4614), .D(n4983), .Y(n4982) );
  OAI22X1 U2517 ( .A(n4644), .B(n4617), .C(n4707), .D(n4615), .Y(n4983) );
  XNOR2X1 U2518 ( .A(n4984), .B(n4616), .Y(n3597) );
  OAI21X1 U2519 ( .A(n4706), .B(n4625), .C(n4985), .Y(n4984) );
  OAI22X1 U2520 ( .A(n4643), .B(n4986), .C(n4614), .D(n4986), .Y(n4985) );
  OAI22X1 U2521 ( .A(n4707), .B(n4617), .C(n4641), .D(n4615), .Y(n4986) );
  XNOR2X1 U2522 ( .A(n4987), .B(n4616), .Y(n3596) );
  OAI21X1 U2523 ( .A(n4705), .B(n4625), .C(n4988), .Y(n4987) );
  OAI22X1 U2524 ( .A(b[28]), .B(n4989), .C(n4614), .D(n4989), .Y(n4988) );
  OAI22X1 U2525 ( .A(n4641), .B(n4617), .C(n4704), .D(n4615), .Y(n4989) );
  XNOR2X1 U2526 ( .A(n4990), .B(n4616), .Y(n3595) );
  OAI21X1 U2527 ( .A(n4703), .B(n4625), .C(n4991), .Y(n4990) );
  OAI22X1 U2528 ( .A(b[29]), .B(n4992), .C(n4614), .D(n4992), .Y(n4991) );
  OAI22X1 U2529 ( .A(n4704), .B(n4617), .C(n4632), .D(n4615), .Y(n4992) );
  NOR2X1 U2530 ( .A(n4993), .B(n4994), .Y(n4902) );
  XNOR2X1 U2531 ( .A(n4995), .B(n4616), .Y(n3594) );
  OAI21X1 U2532 ( .A(n4702), .B(n4625), .C(n4996), .Y(n4995) );
  OAI22X1 U2533 ( .A(b[30]), .B(n4997), .C(n4614), .D(n4997), .Y(n4996) );
  NOR2X1 U2534 ( .A(n4617), .B(n4632), .Y(n4997) );
  NOR2X1 U2535 ( .A(n4762), .B(n4999), .Y(n4901) );
  XNOR2X1 U2536 ( .A(n5000), .B(n4616), .Y(n3593) );
  OAI22X1 U2537 ( .A(n4632), .B(n4998), .C(n4701), .D(n4625), .Y(n5000) );
  NAND3X1 U2538 ( .A(n4994), .B(n4993), .C(n4999), .Y(n4998) );
  XNOR2X1 U2539 ( .A(a[3]), .B(a[4]), .Y(n4999) );
  XNOR2X1 U2540 ( .A(a[4]), .B(n4616), .Y(n4993) );
  XOR2X1 U2541 ( .A(a[3]), .B(n4620), .Y(n4994) );
  XNOR2X1 U2542 ( .A(n5001), .B(n4612), .Y(n3591) );
  OAI22X1 U2543 ( .A(n4700), .B(n4611), .C(n4700), .D(n4626), .Y(n5001) );
  XNOR2X1 U2544 ( .A(n5002), .B(n4759), .Y(n3590) );
  OAI21X1 U2545 ( .A(n4741), .B(n4626), .C(n5003), .Y(n5002) );
  AOI22X1 U2546 ( .A(n5004), .B(n4698), .C(n5005), .D(n4694), .Y(n5003) );
  XNOR2X1 U2547 ( .A(n5006), .B(n4759), .Y(n3589) );
  OAI21X1 U2548 ( .A(n4738), .B(n4626), .C(n5007), .Y(n5006) );
  OAI22X1 U2549 ( .A(n4698), .B(n5008), .C(n4610), .D(n5008), .Y(n5007) );
  OAI22X1 U2550 ( .A(n4695), .B(n4613), .C(n4568), .D(n4611), .Y(n5008) );
  XNOR2X1 U2551 ( .A(n5009), .B(n4759), .Y(n3588) );
  OAI21X1 U2552 ( .A(n4737), .B(n4626), .C(n5010), .Y(n5009) );
  OAI22X1 U2553 ( .A(n4694), .B(n5011), .C(n4610), .D(n5011), .Y(n5010) );
  OAI22X1 U2554 ( .A(n4568), .B(n4613), .C(n4693), .D(n4611), .Y(n5011) );
  XNOR2X1 U2555 ( .A(n5012), .B(n4759), .Y(n3587) );
  OAI21X1 U2556 ( .A(n4736), .B(n4626), .C(n5013), .Y(n5012) );
  OAI22X1 U2557 ( .A(n4569), .B(n5014), .C(n4610), .D(n5014), .Y(n5013) );
  OAI22X1 U2558 ( .A(n4693), .B(n4613), .C(n4570), .D(n4611), .Y(n5014) );
  XNOR2X1 U2559 ( .A(n5015), .B(n4759), .Y(n3586) );
  OAI21X1 U2560 ( .A(n4735), .B(n4626), .C(n5016), .Y(n5015) );
  OAI22X1 U2561 ( .A(n4691), .B(n5017), .C(n4610), .D(n5017), .Y(n5016) );
  OAI22X1 U2562 ( .A(n4570), .B(n4613), .C(n4689), .D(n4611), .Y(n5017) );
  XNOR2X1 U2563 ( .A(n5018), .B(n4759), .Y(n3585) );
  OAI21X1 U2564 ( .A(n4734), .B(n4626), .C(n5019), .Y(n5018) );
  OAI22X1 U2565 ( .A(n4571), .B(n5020), .C(n4610), .D(n5020), .Y(n5019) );
  OAI22X1 U2566 ( .A(n4689), .B(n4613), .C(n4572), .D(n4611), .Y(n5020) );
  XNOR2X1 U2567 ( .A(n5021), .B(n4759), .Y(n3584) );
  OAI21X1 U2568 ( .A(n4733), .B(n4626), .C(n5022), .Y(n5021) );
  OAI22X1 U2569 ( .A(n4687), .B(n5023), .C(n4610), .D(n5023), .Y(n5022) );
  OAI22X1 U2570 ( .A(n4572), .B(n4613), .C(n4685), .D(n4611), .Y(n5023) );
  XNOR2X1 U2571 ( .A(n5024), .B(n4759), .Y(n3583) );
  OAI21X1 U2572 ( .A(n4731), .B(n4626), .C(n5025), .Y(n5024) );
  OAI22X1 U2573 ( .A(n4573), .B(n5026), .C(n4610), .D(n5026), .Y(n5025) );
  OAI22X1 U2574 ( .A(n4685), .B(n4613), .C(n4574), .D(n4611), .Y(n5026) );
  XNOR2X1 U2575 ( .A(n5027), .B(n4759), .Y(n3582) );
  OAI21X1 U2576 ( .A(n4730), .B(n4626), .C(n5028), .Y(n5027) );
  OAI22X1 U2577 ( .A(n4683), .B(n5029), .C(n4610), .D(n5029), .Y(n5028) );
  OAI22X1 U2578 ( .A(n4574), .B(n4613), .C(n4680), .D(n4611), .Y(n5029) );
  XNOR2X1 U2579 ( .A(n5030), .B(n4759), .Y(n3581) );
  OAI21X1 U2580 ( .A(n4729), .B(n4626), .C(n5031), .Y(n5030) );
  OAI22X1 U2581 ( .A(n4575), .B(n5032), .C(n4610), .D(n5032), .Y(n5031) );
  OAI22X1 U2582 ( .A(n4680), .B(n4613), .C(n4576), .D(n4611), .Y(n5032) );
  XNOR2X1 U2583 ( .A(n5033), .B(n4759), .Y(n3580) );
  OAI21X1 U2584 ( .A(n4727), .B(n4626), .C(n5034), .Y(n5033) );
  OAI22X1 U2585 ( .A(n4678), .B(n5035), .C(n4610), .D(n5035), .Y(n5034) );
  OAI22X1 U2586 ( .A(n4576), .B(n4613), .C(n4676), .D(n4611), .Y(n5035) );
  XNOR2X1 U2587 ( .A(n5036), .B(n4759), .Y(n3579) );
  OAI21X1 U2588 ( .A(n4726), .B(n4626), .C(n5037), .Y(n5036) );
  OAI22X1 U2589 ( .A(n4577), .B(n5038), .C(n4610), .D(n5038), .Y(n5037) );
  OAI22X1 U2590 ( .A(n4676), .B(n4613), .C(n4578), .D(n4611), .Y(n5038) );
  XNOR2X1 U2591 ( .A(n5039), .B(n4759), .Y(n3578) );
  OAI21X1 U2592 ( .A(n4725), .B(n4626), .C(n5040), .Y(n5039) );
  OAI22X1 U2593 ( .A(n4674), .B(n5041), .C(n4610), .D(n5041), .Y(n5040) );
  OAI22X1 U2594 ( .A(n4578), .B(n4613), .C(n4671), .D(n4611), .Y(n5041) );
  XNOR2X1 U2595 ( .A(n5042), .B(n4759), .Y(n3577) );
  OAI21X1 U2596 ( .A(n4724), .B(n4626), .C(n5043), .Y(n5042) );
  OAI22X1 U2597 ( .A(n4579), .B(n5044), .C(n4610), .D(n5044), .Y(n5043) );
  OAI22X1 U2598 ( .A(n4671), .B(n4613), .C(n4580), .D(n4611), .Y(n5044) );
  XNOR2X1 U2599 ( .A(n5045), .B(n4759), .Y(n3576) );
  OAI21X1 U2600 ( .A(n4722), .B(n4626), .C(n5046), .Y(n5045) );
  OAI22X1 U2601 ( .A(n4669), .B(n5047), .C(n4610), .D(n5047), .Y(n5046) );
  OAI22X1 U2602 ( .A(n4580), .B(n4613), .C(n4666), .D(n4611), .Y(n5047) );
  XNOR2X1 U2603 ( .A(n5048), .B(n4759), .Y(n3575) );
  OAI21X1 U2604 ( .A(n4721), .B(n4626), .C(n5049), .Y(n5048) );
  OAI22X1 U2605 ( .A(n4581), .B(n5050), .C(n4610), .D(n5050), .Y(n5049) );
  OAI22X1 U2606 ( .A(n4666), .B(n4613), .C(n4582), .D(n4611), .Y(n5050) );
  XNOR2X1 U2607 ( .A(n5051), .B(n4759), .Y(n3574) );
  OAI21X1 U2608 ( .A(n4720), .B(n4626), .C(n5052), .Y(n5051) );
  OAI22X1 U2609 ( .A(n4664), .B(n5053), .C(n4610), .D(n5053), .Y(n5052) );
  OAI22X1 U2610 ( .A(n4582), .B(n4613), .C(n4662), .D(n4611), .Y(n5053) );
  XNOR2X1 U2611 ( .A(n5054), .B(n4759), .Y(n3573) );
  OAI21X1 U2612 ( .A(n4719), .B(n4626), .C(n5055), .Y(n5054) );
  OAI22X1 U2613 ( .A(n4583), .B(n5056), .C(n4610), .D(n5056), .Y(n5055) );
  OAI22X1 U2614 ( .A(n4662), .B(n4613), .C(n4584), .D(n4611), .Y(n5056) );
  XNOR2X1 U2615 ( .A(n5057), .B(n4759), .Y(n3572) );
  OAI21X1 U2616 ( .A(n4718), .B(n4626), .C(n5058), .Y(n5057) );
  OAI22X1 U2617 ( .A(n4660), .B(n5059), .C(n4610), .D(n5059), .Y(n5058) );
  OAI22X1 U2618 ( .A(n4584), .B(n4613), .C(n4657), .D(n4611), .Y(n5059) );
  XNOR2X1 U2619 ( .A(n5060), .B(n4612), .Y(n3571) );
  OAI21X1 U2620 ( .A(n4717), .B(n4626), .C(n5061), .Y(n5060) );
  OAI22X1 U2621 ( .A(n4585), .B(n5062), .C(n4610), .D(n5062), .Y(n5061) );
  OAI22X1 U2622 ( .A(n4657), .B(n4613), .C(n4586), .D(n4611), .Y(n5062) );
  XNOR2X1 U2623 ( .A(n5063), .B(n4612), .Y(n3570) );
  OAI21X1 U2624 ( .A(n4716), .B(n4626), .C(n5064), .Y(n5063) );
  OAI22X1 U2625 ( .A(n4656), .B(n5065), .C(n4610), .D(n5065), .Y(n5064) );
  OAI22X1 U2626 ( .A(n4586), .B(n4613), .C(n4654), .D(n4611), .Y(n5065) );
  XNOR2X1 U2627 ( .A(n5066), .B(n4612), .Y(n3569) );
  OAI21X1 U2628 ( .A(n4715), .B(n4626), .C(n5067), .Y(n5066) );
  OAI22X1 U2629 ( .A(n4587), .B(n5068), .C(n4610), .D(n5068), .Y(n5067) );
  OAI22X1 U2630 ( .A(n4654), .B(n4613), .C(n4588), .D(n4611), .Y(n5068) );
  XNOR2X1 U2631 ( .A(n5069), .B(n4612), .Y(n3568) );
  OAI21X1 U2632 ( .A(n4714), .B(n4626), .C(n5070), .Y(n5069) );
  OAI22X1 U2633 ( .A(n4653), .B(n5071), .C(n4610), .D(n5071), .Y(n5070) );
  OAI22X1 U2634 ( .A(n4588), .B(n4613), .C(n4650), .D(n4611), .Y(n5071) );
  XNOR2X1 U2635 ( .A(n5072), .B(n4612), .Y(n3567) );
  OAI21X1 U2636 ( .A(n4713), .B(n4626), .C(n5073), .Y(n5072) );
  OAI22X1 U2637 ( .A(n4589), .B(n5074), .C(n4610), .D(n5074), .Y(n5073) );
  OAI22X1 U2638 ( .A(n4650), .B(n4613), .C(n4590), .D(n4611), .Y(n5074) );
  XNOR2X1 U2639 ( .A(n5075), .B(n4612), .Y(n3566) );
  OAI21X1 U2640 ( .A(n4712), .B(n4626), .C(n5076), .Y(n5075) );
  OAI22X1 U2641 ( .A(n4649), .B(n5077), .C(n4610), .D(n5077), .Y(n5076) );
  OAI22X1 U2642 ( .A(n4590), .B(n4613), .C(n4647), .D(n4611), .Y(n5077) );
  XNOR2X1 U2643 ( .A(n5078), .B(n4612), .Y(n3565) );
  OAI21X1 U2644 ( .A(n4711), .B(n4626), .C(n5079), .Y(n5078) );
  OAI22X1 U2645 ( .A(n4591), .B(n5080), .C(n4610), .D(n5080), .Y(n5079) );
  OAI22X1 U2646 ( .A(n4647), .B(n4613), .C(n4710), .D(n4611), .Y(n5080) );
  XNOR2X1 U2647 ( .A(n5081), .B(n4612), .Y(n3564) );
  OAI21X1 U2648 ( .A(n4709), .B(n4626), .C(n5082), .Y(n5081) );
  OAI22X1 U2649 ( .A(n4646), .B(n5083), .C(n4610), .D(n5083), .Y(n5082) );
  OAI22X1 U2650 ( .A(n4710), .B(n4613), .C(n4644), .D(n4611), .Y(n5083) );
  XNOR2X1 U2651 ( .A(n5084), .B(n4612), .Y(n3563) );
  OAI21X1 U2652 ( .A(n4708), .B(n4626), .C(n5085), .Y(n5084) );
  OAI22X1 U2653 ( .A(b[26]), .B(n5086), .C(n4610), .D(n5086), .Y(n5085) );
  OAI22X1 U2654 ( .A(n4644), .B(n4613), .C(n4707), .D(n4611), .Y(n5086) );
  XNOR2X1 U2655 ( .A(n5087), .B(n4612), .Y(n3562) );
  OAI21X1 U2656 ( .A(n4706), .B(n4626), .C(n5088), .Y(n5087) );
  OAI22X1 U2657 ( .A(n4643), .B(n5089), .C(n4610), .D(n5089), .Y(n5088) );
  OAI22X1 U2658 ( .A(n4707), .B(n4613), .C(n4641), .D(n4611), .Y(n5089) );
  XNOR2X1 U2659 ( .A(n5090), .B(n4612), .Y(n3561) );
  OAI21X1 U2660 ( .A(n4705), .B(n4626), .C(n5091), .Y(n5090) );
  OAI22X1 U2661 ( .A(b[28]), .B(n5092), .C(n4610), .D(n5092), .Y(n5091) );
  OAI22X1 U2662 ( .A(n4641), .B(n4613), .C(n4704), .D(n4611), .Y(n5092) );
  XNOR2X1 U2663 ( .A(n5093), .B(n4612), .Y(n3560) );
  OAI21X1 U2664 ( .A(n4703), .B(n4626), .C(n5094), .Y(n5093) );
  OAI22X1 U2665 ( .A(b[29]), .B(n5095), .C(n4610), .D(n5095), .Y(n5094) );
  OAI22X1 U2666 ( .A(n4704), .B(n4613), .C(n4632), .D(n4611), .Y(n5095) );
  NOR2X1 U2667 ( .A(n5096), .B(n5097), .Y(n5005) );
  XNOR2X1 U2668 ( .A(n5098), .B(n4612), .Y(n3559) );
  OAI21X1 U2669 ( .A(n4702), .B(n4626), .C(n5099), .Y(n5098) );
  OAI22X1 U2670 ( .A(b[30]), .B(n5100), .C(n4610), .D(n5100), .Y(n5099) );
  NOR2X1 U2671 ( .A(n4613), .B(n4632), .Y(n5100) );
  NOR2X1 U2672 ( .A(n4760), .B(n5102), .Y(n5004) );
  XNOR2X1 U2673 ( .A(n5103), .B(n4612), .Y(n3558) );
  OAI22X1 U2674 ( .A(n4632), .B(n5101), .C(n4701), .D(n4626), .Y(n5103) );
  NAND3X1 U2675 ( .A(n5097), .B(n5096), .C(n5102), .Y(n5101) );
  XNOR2X1 U2676 ( .A(a[6]), .B(a[7]), .Y(n5102) );
  XNOR2X1 U2677 ( .A(a[7]), .B(n4612), .Y(n5096) );
  XOR2X1 U2678 ( .A(a[6]), .B(n4616), .Y(n5097) );
  XNOR2X1 U2679 ( .A(n5104), .B(n4608), .Y(n3556) );
  OAI22X1 U2680 ( .A(n4700), .B(n4607), .C(n4700), .D(n4627), .Y(n5104) );
  XNOR2X1 U2681 ( .A(n5105), .B(n4757), .Y(n3555) );
  OAI21X1 U2682 ( .A(n4741), .B(n4627), .C(n5106), .Y(n5105) );
  AOI22X1 U2683 ( .A(n5107), .B(n4698), .C(n5108), .D(n4694), .Y(n5106) );
  XNOR2X1 U2684 ( .A(n5109), .B(n4757), .Y(n3554) );
  OAI21X1 U2685 ( .A(n4738), .B(n4627), .C(n5110), .Y(n5109) );
  OAI22X1 U2686 ( .A(n4699), .B(n5111), .C(n4606), .D(n5111), .Y(n5110) );
  OAI22X1 U2687 ( .A(n4695), .B(n4609), .C(n4568), .D(n4607), .Y(n5111) );
  XNOR2X1 U2688 ( .A(n5112), .B(n4757), .Y(n3553) );
  OAI21X1 U2689 ( .A(n4737), .B(n4627), .C(n5113), .Y(n5112) );
  OAI22X1 U2690 ( .A(n4694), .B(n5114), .C(n4606), .D(n5114), .Y(n5113) );
  OAI22X1 U2691 ( .A(n4568), .B(n4609), .C(n4693), .D(n4607), .Y(n5114) );
  XNOR2X1 U2692 ( .A(n5115), .B(n4757), .Y(n3552) );
  OAI21X1 U2693 ( .A(n4736), .B(n4627), .C(n5116), .Y(n5115) );
  OAI22X1 U2694 ( .A(n4569), .B(n5117), .C(n4606), .D(n5117), .Y(n5116) );
  OAI22X1 U2695 ( .A(n4693), .B(n4609), .C(n4570), .D(n4607), .Y(n5117) );
  XNOR2X1 U2696 ( .A(n5118), .B(n4757), .Y(n3551) );
  OAI21X1 U2697 ( .A(n4735), .B(n4627), .C(n5119), .Y(n5118) );
  OAI22X1 U2698 ( .A(n4691), .B(n5120), .C(n4606), .D(n5120), .Y(n5119) );
  OAI22X1 U2699 ( .A(n4570), .B(n4609), .C(n4689), .D(n4607), .Y(n5120) );
  XNOR2X1 U2700 ( .A(n5121), .B(n4757), .Y(n3550) );
  OAI21X1 U2701 ( .A(n4734), .B(n4627), .C(n5122), .Y(n5121) );
  OAI22X1 U2702 ( .A(n4571), .B(n5123), .C(n4606), .D(n5123), .Y(n5122) );
  OAI22X1 U2703 ( .A(n4689), .B(n4609), .C(n4572), .D(n4607), .Y(n5123) );
  XNOR2X1 U2704 ( .A(n5124), .B(n4757), .Y(n3549) );
  OAI21X1 U2705 ( .A(n4733), .B(n4627), .C(n5125), .Y(n5124) );
  OAI22X1 U2706 ( .A(n4687), .B(n5126), .C(n4606), .D(n5126), .Y(n5125) );
  OAI22X1 U2707 ( .A(n4572), .B(n4609), .C(n4685), .D(n4607), .Y(n5126) );
  XNOR2X1 U2708 ( .A(n5127), .B(n4757), .Y(n3548) );
  OAI21X1 U2709 ( .A(n4731), .B(n4627), .C(n5128), .Y(n5127) );
  OAI22X1 U2710 ( .A(n4573), .B(n5129), .C(n4606), .D(n5129), .Y(n5128) );
  OAI22X1 U2711 ( .A(n4685), .B(n4609), .C(n4574), .D(n4607), .Y(n5129) );
  XNOR2X1 U2712 ( .A(n5130), .B(n4757), .Y(n3547) );
  OAI21X1 U2713 ( .A(n4730), .B(n4627), .C(n5131), .Y(n5130) );
  OAI22X1 U2714 ( .A(n4683), .B(n5132), .C(n4606), .D(n5132), .Y(n5131) );
  OAI22X1 U2715 ( .A(n4574), .B(n4609), .C(n4680), .D(n4607), .Y(n5132) );
  XNOR2X1 U2716 ( .A(n5133), .B(n4757), .Y(n3546) );
  OAI21X1 U2717 ( .A(n4729), .B(n4627), .C(n5134), .Y(n5133) );
  OAI22X1 U2718 ( .A(n4575), .B(n5135), .C(n4606), .D(n5135), .Y(n5134) );
  OAI22X1 U2719 ( .A(n4680), .B(n4609), .C(n4576), .D(n4607), .Y(n5135) );
  XNOR2X1 U2720 ( .A(n5136), .B(n4757), .Y(n3545) );
  OAI21X1 U2721 ( .A(n4727), .B(n4627), .C(n5137), .Y(n5136) );
  OAI22X1 U2722 ( .A(n4678), .B(n5138), .C(n4606), .D(n5138), .Y(n5137) );
  OAI22X1 U2723 ( .A(n4576), .B(n4609), .C(n4676), .D(n4607), .Y(n5138) );
  XNOR2X1 U2724 ( .A(n5139), .B(n4757), .Y(n3544) );
  OAI21X1 U2725 ( .A(n4726), .B(n4627), .C(n5140), .Y(n5139) );
  OAI22X1 U2726 ( .A(n4577), .B(n5141), .C(n4606), .D(n5141), .Y(n5140) );
  OAI22X1 U2727 ( .A(n4676), .B(n4609), .C(n4578), .D(n4607), .Y(n5141) );
  XNOR2X1 U2728 ( .A(n5142), .B(n4757), .Y(n3543) );
  OAI21X1 U2729 ( .A(n4725), .B(n4627), .C(n5143), .Y(n5142) );
  OAI22X1 U2730 ( .A(n4674), .B(n5144), .C(n4606), .D(n5144), .Y(n5143) );
  OAI22X1 U2731 ( .A(n4578), .B(n4609), .C(n4671), .D(n4607), .Y(n5144) );
  XNOR2X1 U2732 ( .A(n5145), .B(n4757), .Y(n3542) );
  OAI21X1 U2733 ( .A(n4724), .B(n4627), .C(n5146), .Y(n5145) );
  OAI22X1 U2734 ( .A(n4579), .B(n5147), .C(n4606), .D(n5147), .Y(n5146) );
  OAI22X1 U2735 ( .A(n4671), .B(n4609), .C(n4580), .D(n4607), .Y(n5147) );
  XNOR2X1 U2736 ( .A(n5148), .B(n4757), .Y(n3541) );
  OAI21X1 U2737 ( .A(n4722), .B(n4627), .C(n5149), .Y(n5148) );
  OAI22X1 U2738 ( .A(n4669), .B(n5150), .C(n4606), .D(n5150), .Y(n5149) );
  OAI22X1 U2739 ( .A(n4580), .B(n4609), .C(n4666), .D(n4607), .Y(n5150) );
  XNOR2X1 U2740 ( .A(n5151), .B(n4757), .Y(n3540) );
  OAI21X1 U2741 ( .A(n4721), .B(n4627), .C(n5152), .Y(n5151) );
  OAI22X1 U2742 ( .A(n4581), .B(n5153), .C(n4606), .D(n5153), .Y(n5152) );
  OAI22X1 U2743 ( .A(n4666), .B(n4609), .C(n4582), .D(n4607), .Y(n5153) );
  XNOR2X1 U2744 ( .A(n5154), .B(n4757), .Y(n3539) );
  OAI21X1 U2745 ( .A(n4720), .B(n4627), .C(n5155), .Y(n5154) );
  OAI22X1 U2746 ( .A(n4664), .B(n5156), .C(n4606), .D(n5156), .Y(n5155) );
  OAI22X1 U2747 ( .A(n4582), .B(n4609), .C(n4662), .D(n4607), .Y(n5156) );
  XNOR2X1 U2748 ( .A(n5157), .B(n4757), .Y(n3538) );
  OAI21X1 U2749 ( .A(n4719), .B(n4627), .C(n5158), .Y(n5157) );
  OAI22X1 U2750 ( .A(n4583), .B(n5159), .C(n4606), .D(n5159), .Y(n5158) );
  OAI22X1 U2751 ( .A(n4662), .B(n4609), .C(n4584), .D(n4607), .Y(n5159) );
  XNOR2X1 U2752 ( .A(n5160), .B(n4757), .Y(n3537) );
  OAI21X1 U2753 ( .A(n4718), .B(n4627), .C(n5161), .Y(n5160) );
  OAI22X1 U2754 ( .A(n4660), .B(n5162), .C(n4606), .D(n5162), .Y(n5161) );
  OAI22X1 U2755 ( .A(n4584), .B(n4609), .C(n4657), .D(n4607), .Y(n5162) );
  XNOR2X1 U2756 ( .A(n5163), .B(n4608), .Y(n3536) );
  OAI21X1 U2757 ( .A(n4717), .B(n4627), .C(n5164), .Y(n5163) );
  OAI22X1 U2758 ( .A(n4585), .B(n5165), .C(n4606), .D(n5165), .Y(n5164) );
  OAI22X1 U2759 ( .A(n4657), .B(n4609), .C(n4586), .D(n4607), .Y(n5165) );
  XNOR2X1 U2760 ( .A(n5166), .B(n4608), .Y(n3535) );
  OAI21X1 U2761 ( .A(n4716), .B(n4627), .C(n5167), .Y(n5166) );
  OAI22X1 U2762 ( .A(n4656), .B(n5168), .C(n4606), .D(n5168), .Y(n5167) );
  OAI22X1 U2763 ( .A(n4586), .B(n4609), .C(n4654), .D(n4607), .Y(n5168) );
  XNOR2X1 U2764 ( .A(n5169), .B(n4608), .Y(n3534) );
  OAI21X1 U2765 ( .A(n4715), .B(n4627), .C(n5170), .Y(n5169) );
  OAI22X1 U2766 ( .A(n4587), .B(n5171), .C(n4606), .D(n5171), .Y(n5170) );
  OAI22X1 U2767 ( .A(n4654), .B(n4609), .C(n4588), .D(n4607), .Y(n5171) );
  XNOR2X1 U2768 ( .A(n5172), .B(n4608), .Y(n3533) );
  OAI21X1 U2769 ( .A(n4714), .B(n4627), .C(n5173), .Y(n5172) );
  OAI22X1 U2770 ( .A(n4653), .B(n5174), .C(n4606), .D(n5174), .Y(n5173) );
  OAI22X1 U2771 ( .A(n4588), .B(n4609), .C(n4650), .D(n4607), .Y(n5174) );
  XNOR2X1 U2772 ( .A(n5175), .B(n4608), .Y(n3532) );
  OAI21X1 U2773 ( .A(n4713), .B(n4627), .C(n5176), .Y(n5175) );
  OAI22X1 U2774 ( .A(n4589), .B(n5177), .C(n4606), .D(n5177), .Y(n5176) );
  OAI22X1 U2775 ( .A(n4650), .B(n4609), .C(n4590), .D(n4607), .Y(n5177) );
  XNOR2X1 U2776 ( .A(n5178), .B(n4608), .Y(n3531) );
  OAI21X1 U2777 ( .A(n4712), .B(n4627), .C(n5179), .Y(n5178) );
  OAI22X1 U2778 ( .A(n4649), .B(n5180), .C(n4606), .D(n5180), .Y(n5179) );
  OAI22X1 U2779 ( .A(n4590), .B(n4609), .C(n4647), .D(n4607), .Y(n5180) );
  XNOR2X1 U2780 ( .A(n5181), .B(n4608), .Y(n3530) );
  OAI21X1 U2781 ( .A(n4711), .B(n4627), .C(n5182), .Y(n5181) );
  OAI22X1 U2782 ( .A(n4591), .B(n5183), .C(n4606), .D(n5183), .Y(n5182) );
  OAI22X1 U2783 ( .A(n4647), .B(n4609), .C(n4710), .D(n4607), .Y(n5183) );
  XNOR2X1 U2784 ( .A(n5184), .B(n4608), .Y(n3529) );
  OAI21X1 U2785 ( .A(n4709), .B(n4627), .C(n5185), .Y(n5184) );
  OAI22X1 U2786 ( .A(n4646), .B(n5186), .C(n4606), .D(n5186), .Y(n5185) );
  OAI22X1 U2787 ( .A(n4710), .B(n4609), .C(n4644), .D(n4607), .Y(n5186) );
  XNOR2X1 U2788 ( .A(n5187), .B(n4608), .Y(n3528) );
  OAI21X1 U2789 ( .A(n4708), .B(n4627), .C(n5188), .Y(n5187) );
  OAI22X1 U2790 ( .A(b[26]), .B(n5189), .C(n4606), .D(n5189), .Y(n5188) );
  OAI22X1 U2791 ( .A(n4644), .B(n4609), .C(n4707), .D(n4607), .Y(n5189) );
  XNOR2X1 U2792 ( .A(n5190), .B(n4608), .Y(n3527) );
  OAI21X1 U2793 ( .A(n4706), .B(n4627), .C(n5191), .Y(n5190) );
  OAI22X1 U2794 ( .A(n4643), .B(n5192), .C(n4606), .D(n5192), .Y(n5191) );
  OAI22X1 U2795 ( .A(n4707), .B(n4609), .C(n4641), .D(n4607), .Y(n5192) );
  XNOR2X1 U2796 ( .A(n5193), .B(n4608), .Y(n3526) );
  OAI21X1 U2797 ( .A(n4705), .B(n4627), .C(n5194), .Y(n5193) );
  OAI22X1 U2798 ( .A(b[28]), .B(n5195), .C(n4606), .D(n5195), .Y(n5194) );
  OAI22X1 U2799 ( .A(n4641), .B(n4609), .C(n4704), .D(n4607), .Y(n5195) );
  XNOR2X1 U2800 ( .A(n5196), .B(n4608), .Y(n3525) );
  OAI21X1 U2801 ( .A(n4703), .B(n4627), .C(n5197), .Y(n5196) );
  OAI22X1 U2802 ( .A(b[29]), .B(n5198), .C(n4606), .D(n5198), .Y(n5197) );
  OAI22X1 U2803 ( .A(n4704), .B(n4609), .C(n4632), .D(n4607), .Y(n5198) );
  NOR2X1 U2804 ( .A(n5199), .B(n5200), .Y(n5108) );
  XNOR2X1 U2805 ( .A(n5201), .B(n4608), .Y(n3524) );
  OAI21X1 U2806 ( .A(n4702), .B(n4627), .C(n5202), .Y(n5201) );
  OAI22X1 U2807 ( .A(b[30]), .B(n5203), .C(n4606), .D(n5203), .Y(n5202) );
  NOR2X1 U2808 ( .A(n4609), .B(n4632), .Y(n5203) );
  NOR2X1 U2809 ( .A(n4758), .B(n5205), .Y(n5107) );
  XNOR2X1 U2810 ( .A(n5206), .B(n4608), .Y(n3523) );
  OAI22X1 U2811 ( .A(n4632), .B(n5204), .C(n4701), .D(n4627), .Y(n5206) );
  NAND3X1 U2812 ( .A(n5200), .B(n5199), .C(n5205), .Y(n5204) );
  XNOR2X1 U2813 ( .A(a[10]), .B(a[9]), .Y(n5205) );
  XNOR2X1 U2814 ( .A(a[10]), .B(n4608), .Y(n5199) );
  XOR2X1 U2815 ( .A(a[9]), .B(n4612), .Y(n5200) );
  XNOR2X1 U2816 ( .A(n5207), .B(n4603), .Y(n3521) );
  OAI22X1 U2817 ( .A(n4700), .B(n4602), .C(n4700), .D(n4628), .Y(n5207) );
  XNOR2X1 U2818 ( .A(n5208), .B(n4603), .Y(n3520) );
  OAI21X1 U2819 ( .A(n4741), .B(n4628), .C(n5209), .Y(n5208) );
  AOI22X1 U2820 ( .A(n5210), .B(n4698), .C(n5211), .D(n4694), .Y(n5209) );
  XNOR2X1 U2821 ( .A(n5212), .B(n4603), .Y(n3519) );
  OAI21X1 U2822 ( .A(n4738), .B(n4628), .C(n5213), .Y(n5212) );
  OAI22X1 U2823 ( .A(n4699), .B(n5214), .C(n4601), .D(n5214), .Y(n5213) );
  OAI22X1 U2824 ( .A(n4695), .B(n4605), .C(n4568), .D(n4602), .Y(n5214) );
  XNOR2X1 U2825 ( .A(n5215), .B(n4603), .Y(n3518) );
  OAI21X1 U2826 ( .A(n4737), .B(n4628), .C(n5216), .Y(n5215) );
  OAI22X1 U2827 ( .A(n4694), .B(n5217), .C(n4601), .D(n5217), .Y(n5216) );
  OAI22X1 U2828 ( .A(n4568), .B(n4605), .C(n4693), .D(n4602), .Y(n5217) );
  XNOR2X1 U2829 ( .A(n5218), .B(n4603), .Y(n3517) );
  OAI21X1 U2830 ( .A(n4736), .B(n4628), .C(n5219), .Y(n5218) );
  OAI22X1 U2831 ( .A(n4569), .B(n5220), .C(n4601), .D(n5220), .Y(n5219) );
  OAI22X1 U2832 ( .A(n4693), .B(n4605), .C(n4570), .D(n4602), .Y(n5220) );
  XNOR2X1 U2833 ( .A(n5221), .B(n4603), .Y(n3516) );
  OAI21X1 U2834 ( .A(n4735), .B(n4628), .C(n5222), .Y(n5221) );
  OAI22X1 U2835 ( .A(n4691), .B(n5223), .C(n4601), .D(n5223), .Y(n5222) );
  OAI22X1 U2836 ( .A(n4570), .B(n4605), .C(n4689), .D(n4602), .Y(n5223) );
  XNOR2X1 U2837 ( .A(n5224), .B(n4603), .Y(n3515) );
  OAI21X1 U2838 ( .A(n4734), .B(n4628), .C(n5225), .Y(n5224) );
  OAI22X1 U2839 ( .A(n4571), .B(n5226), .C(n4601), .D(n5226), .Y(n5225) );
  OAI22X1 U2840 ( .A(n4689), .B(n4605), .C(n4572), .D(n4602), .Y(n5226) );
  XNOR2X1 U2841 ( .A(n5227), .B(n4603), .Y(n3514) );
  OAI21X1 U2842 ( .A(n4733), .B(n4628), .C(n5228), .Y(n5227) );
  OAI22X1 U2843 ( .A(n4687), .B(n5229), .C(n4601), .D(n5229), .Y(n5228) );
  OAI22X1 U2844 ( .A(n4572), .B(n4605), .C(n4685), .D(n4602), .Y(n5229) );
  XNOR2X1 U2845 ( .A(n5230), .B(n4603), .Y(n3513) );
  OAI21X1 U2846 ( .A(n4731), .B(n4628), .C(n5231), .Y(n5230) );
  OAI22X1 U2847 ( .A(n4573), .B(n5232), .C(n4601), .D(n5232), .Y(n5231) );
  OAI22X1 U2848 ( .A(n4685), .B(n4605), .C(n4574), .D(n4602), .Y(n5232) );
  XNOR2X1 U2849 ( .A(n5233), .B(n4603), .Y(n3512) );
  OAI21X1 U2850 ( .A(n4730), .B(n4628), .C(n5234), .Y(n5233) );
  OAI22X1 U2851 ( .A(n4683), .B(n5235), .C(n4601), .D(n5235), .Y(n5234) );
  OAI22X1 U2852 ( .A(n4574), .B(n4605), .C(n4680), .D(n4602), .Y(n5235) );
  XNOR2X1 U2853 ( .A(n5236), .B(n4603), .Y(n3511) );
  OAI21X1 U2854 ( .A(n4729), .B(n4628), .C(n5237), .Y(n5236) );
  OAI22X1 U2855 ( .A(n4575), .B(n5238), .C(n4601), .D(n5238), .Y(n5237) );
  OAI22X1 U2856 ( .A(n4680), .B(n4605), .C(n4576), .D(n4602), .Y(n5238) );
  XNOR2X1 U2857 ( .A(n5239), .B(n4603), .Y(n3510) );
  OAI21X1 U2858 ( .A(n4727), .B(n4628), .C(n5240), .Y(n5239) );
  OAI22X1 U2859 ( .A(n4678), .B(n5241), .C(n4601), .D(n5241), .Y(n5240) );
  OAI22X1 U2860 ( .A(n4576), .B(n4605), .C(n4676), .D(n4602), .Y(n5241) );
  XNOR2X1 U2861 ( .A(n5242), .B(n4603), .Y(n3509) );
  OAI21X1 U2862 ( .A(n4726), .B(n4628), .C(n5243), .Y(n5242) );
  OAI22X1 U2863 ( .A(n4577), .B(n5244), .C(n4601), .D(n5244), .Y(n5243) );
  OAI22X1 U2864 ( .A(n4676), .B(n4605), .C(n4578), .D(n4602), .Y(n5244) );
  XNOR2X1 U2865 ( .A(n5245), .B(n4603), .Y(n3508) );
  OAI21X1 U2866 ( .A(n4725), .B(n4628), .C(n5246), .Y(n5245) );
  OAI22X1 U2867 ( .A(n4674), .B(n5247), .C(n4601), .D(n5247), .Y(n5246) );
  OAI22X1 U2868 ( .A(n4578), .B(n4605), .C(n4671), .D(n4602), .Y(n5247) );
  XNOR2X1 U2869 ( .A(n5248), .B(n4603), .Y(n3507) );
  OAI21X1 U2870 ( .A(n4724), .B(n4628), .C(n5249), .Y(n5248) );
  OAI22X1 U2871 ( .A(n4579), .B(n5250), .C(n4601), .D(n5250), .Y(n5249) );
  OAI22X1 U2872 ( .A(n4671), .B(n4605), .C(n4580), .D(n4602), .Y(n5250) );
  XNOR2X1 U2873 ( .A(n5251), .B(n4603), .Y(n3506) );
  OAI21X1 U2874 ( .A(n4722), .B(n4628), .C(n5252), .Y(n5251) );
  OAI22X1 U2875 ( .A(n4669), .B(n5253), .C(n4601), .D(n5253), .Y(n5252) );
  OAI22X1 U2876 ( .A(n4580), .B(n4605), .C(n4666), .D(n4602), .Y(n5253) );
  XNOR2X1 U2877 ( .A(n5254), .B(n4603), .Y(n3505) );
  OAI21X1 U2878 ( .A(n4721), .B(n4628), .C(n5255), .Y(n5254) );
  OAI22X1 U2879 ( .A(n4581), .B(n5256), .C(n4601), .D(n5256), .Y(n5255) );
  OAI22X1 U2880 ( .A(n4666), .B(n4605), .C(n4582), .D(n4602), .Y(n5256) );
  XNOR2X1 U2881 ( .A(n5257), .B(n4603), .Y(n3504) );
  OAI21X1 U2882 ( .A(n4720), .B(n4628), .C(n5258), .Y(n5257) );
  OAI22X1 U2883 ( .A(n4664), .B(n5259), .C(n4601), .D(n5259), .Y(n5258) );
  OAI22X1 U2884 ( .A(n4582), .B(n4605), .C(n4662), .D(n4602), .Y(n5259) );
  XNOR2X1 U2885 ( .A(n5260), .B(n4603), .Y(n3503) );
  OAI21X1 U2886 ( .A(n4719), .B(n4628), .C(n5261), .Y(n5260) );
  OAI22X1 U2887 ( .A(n4583), .B(n5262), .C(n4601), .D(n5262), .Y(n5261) );
  OAI22X1 U2888 ( .A(n4662), .B(n4605), .C(n4584), .D(n4602), .Y(n5262) );
  XNOR2X1 U2889 ( .A(n5263), .B(n4603), .Y(n3502) );
  OAI21X1 U2890 ( .A(n4718), .B(n4628), .C(n5264), .Y(n5263) );
  OAI22X1 U2891 ( .A(n4660), .B(n5265), .C(n4601), .D(n5265), .Y(n5264) );
  OAI22X1 U2892 ( .A(n4584), .B(n4605), .C(n4657), .D(n4602), .Y(n5265) );
  XNOR2X1 U2893 ( .A(n5266), .B(n4604), .Y(n3501) );
  OAI21X1 U2894 ( .A(n4717), .B(n4628), .C(n5267), .Y(n5266) );
  OAI22X1 U2895 ( .A(n4585), .B(n5268), .C(n4601), .D(n5268), .Y(n5267) );
  OAI22X1 U2896 ( .A(n4657), .B(n4605), .C(n4586), .D(n4602), .Y(n5268) );
  XNOR2X1 U2897 ( .A(n5269), .B(n4604), .Y(n3500) );
  OAI21X1 U2898 ( .A(n4716), .B(n4628), .C(n5270), .Y(n5269) );
  OAI22X1 U2899 ( .A(n4656), .B(n5271), .C(n4601), .D(n5271), .Y(n5270) );
  OAI22X1 U2900 ( .A(n4586), .B(n4605), .C(n4654), .D(n4602), .Y(n5271) );
  XNOR2X1 U2901 ( .A(n5272), .B(n4604), .Y(n3499) );
  OAI21X1 U2902 ( .A(n4715), .B(n4628), .C(n5273), .Y(n5272) );
  OAI22X1 U2903 ( .A(n4587), .B(n5274), .C(n4601), .D(n5274), .Y(n5273) );
  OAI22X1 U2904 ( .A(n4654), .B(n4605), .C(n4588), .D(n4602), .Y(n5274) );
  XNOR2X1 U2905 ( .A(n5275), .B(n4604), .Y(n3498) );
  OAI21X1 U2906 ( .A(n4714), .B(n4628), .C(n5276), .Y(n5275) );
  OAI22X1 U2907 ( .A(n4653), .B(n5277), .C(n4601), .D(n5277), .Y(n5276) );
  OAI22X1 U2908 ( .A(n4588), .B(n4605), .C(n4650), .D(n4602), .Y(n5277) );
  XNOR2X1 U2909 ( .A(n5278), .B(n4604), .Y(n3497) );
  OAI21X1 U2910 ( .A(n4713), .B(n4628), .C(n5279), .Y(n5278) );
  OAI22X1 U2911 ( .A(n4589), .B(n5280), .C(n4601), .D(n5280), .Y(n5279) );
  OAI22X1 U2912 ( .A(n4650), .B(n4605), .C(n4590), .D(n4602), .Y(n5280) );
  XNOR2X1 U2913 ( .A(n5281), .B(n4604), .Y(n3496) );
  OAI21X1 U2914 ( .A(n4712), .B(n4628), .C(n5282), .Y(n5281) );
  OAI22X1 U2915 ( .A(n4649), .B(n5283), .C(n4601), .D(n5283), .Y(n5282) );
  OAI22X1 U2916 ( .A(n4590), .B(n4605), .C(n4647), .D(n4602), .Y(n5283) );
  XNOR2X1 U2917 ( .A(n5284), .B(n4604), .Y(n3495) );
  OAI21X1 U2918 ( .A(n4711), .B(n4628), .C(n5285), .Y(n5284) );
  OAI22X1 U2919 ( .A(n4591), .B(n5286), .C(n4601), .D(n5286), .Y(n5285) );
  OAI22X1 U2920 ( .A(n4647), .B(n4605), .C(n4710), .D(n4602), .Y(n5286) );
  XNOR2X1 U2921 ( .A(n5287), .B(n4604), .Y(n3494) );
  OAI21X1 U2922 ( .A(n4709), .B(n4628), .C(n5288), .Y(n5287) );
  OAI22X1 U2923 ( .A(n4646), .B(n5289), .C(n4601), .D(n5289), .Y(n5288) );
  OAI22X1 U2924 ( .A(n4710), .B(n4605), .C(n4644), .D(n4602), .Y(n5289) );
  XNOR2X1 U2925 ( .A(n5290), .B(n4604), .Y(n3493) );
  OAI21X1 U2926 ( .A(n4708), .B(n4628), .C(n5291), .Y(n5290) );
  OAI22X1 U2927 ( .A(b[26]), .B(n5292), .C(n4601), .D(n5292), .Y(n5291) );
  OAI22X1 U2928 ( .A(n4644), .B(n4605), .C(n4707), .D(n4602), .Y(n5292) );
  XNOR2X1 U2929 ( .A(n5293), .B(n4604), .Y(n3492) );
  OAI21X1 U2930 ( .A(n4706), .B(n4628), .C(n5294), .Y(n5293) );
  OAI22X1 U2931 ( .A(n4643), .B(n5295), .C(n4601), .D(n5295), .Y(n5294) );
  OAI22X1 U2932 ( .A(n4707), .B(n4605), .C(n4641), .D(n4602), .Y(n5295) );
  XNOR2X1 U2933 ( .A(n5296), .B(n4604), .Y(n3491) );
  OAI21X1 U2934 ( .A(n4705), .B(n4628), .C(n5297), .Y(n5296) );
  OAI22X1 U2935 ( .A(b[28]), .B(n5298), .C(n4601), .D(n5298), .Y(n5297) );
  OAI22X1 U2936 ( .A(n4641), .B(n4605), .C(n4704), .D(n4602), .Y(n5298) );
  XNOR2X1 U2937 ( .A(n5299), .B(n4604), .Y(n3490) );
  OAI21X1 U2938 ( .A(n4703), .B(n4628), .C(n5300), .Y(n5299) );
  OAI22X1 U2939 ( .A(b[29]), .B(n5301), .C(n4601), .D(n5301), .Y(n5300) );
  OAI22X1 U2940 ( .A(n4704), .B(n4605), .C(n4632), .D(n4602), .Y(n5301) );
  NOR2X1 U2941 ( .A(n5302), .B(n5303), .Y(n5211) );
  XNOR2X1 U2942 ( .A(n5304), .B(n4604), .Y(n3489) );
  OAI21X1 U2943 ( .A(n4702), .B(n4628), .C(n5305), .Y(n5304) );
  OAI22X1 U2944 ( .A(b[30]), .B(n5306), .C(n4601), .D(n5306), .Y(n5305) );
  NOR2X1 U2945 ( .A(n4605), .B(n4632), .Y(n5306) );
  NOR2X1 U2946 ( .A(n4756), .B(n5308), .Y(n5210) );
  XNOR2X1 U2947 ( .A(n5309), .B(n4604), .Y(n3488) );
  OAI22X1 U2948 ( .A(n4632), .B(n5307), .C(n4701), .D(n4628), .Y(n5309) );
  NAND3X1 U2949 ( .A(n5303), .B(n5302), .C(n5308), .Y(n5307) );
  XNOR2X1 U2950 ( .A(a[12]), .B(a[13]), .Y(n5308) );
  XNOR2X1 U2951 ( .A(a[13]), .B(n4604), .Y(n5302) );
  XOR2X1 U2952 ( .A(a[12]), .B(n4608), .Y(n5303) );
  XNOR2X1 U2953 ( .A(n5310), .B(n4599), .Y(n3486) );
  OAI22X1 U2954 ( .A(n4700), .B(n4629), .C(n4621), .D(n4700), .Y(n5310) );
  XNOR2X1 U2955 ( .A(n5311), .B(n4599), .Y(n3485) );
  OAI21X1 U2956 ( .A(n4621), .B(n4741), .C(n4739), .Y(n5311) );
  OAI22X1 U2957 ( .A(n4700), .B(n4553), .C(n4629), .D(n4695), .Y(n5312) );
  XNOR2X1 U2958 ( .A(n5313), .B(n4599), .Y(n3484) );
  OAI21X1 U2959 ( .A(n4621), .B(n4738), .C(n5314), .Y(n5313) );
  OAI22X1 U2960 ( .A(n4699), .B(n5315), .C(n4598), .D(n5315), .Y(n5314) );
  OAI22X1 U2961 ( .A(n4568), .B(n4629), .C(n4553), .D(n4695), .Y(n5315) );
  XNOR2X1 U2962 ( .A(n5316), .B(n4599), .Y(n3483) );
  OAI21X1 U2963 ( .A(n4621), .B(n4737), .C(n5317), .Y(n5316) );
  OAI22X1 U2964 ( .A(n4694), .B(n5318), .C(n4598), .D(n5318), .Y(n5317) );
  OAI22X1 U2965 ( .A(n4693), .B(n4629), .C(n4553), .D(n4568), .Y(n5318) );
  XNOR2X1 U2966 ( .A(n5319), .B(n4599), .Y(n3482) );
  OAI21X1 U2967 ( .A(n4621), .B(n4736), .C(n5320), .Y(n5319) );
  OAI22X1 U2968 ( .A(n4569), .B(n5321), .C(n4598), .D(n5321), .Y(n5320) );
  OAI22X1 U2969 ( .A(n4570), .B(n4629), .C(n4553), .D(n4693), .Y(n5321) );
  XNOR2X1 U2970 ( .A(n5322), .B(n4599), .Y(n3481) );
  OAI21X1 U2971 ( .A(n4621), .B(n4735), .C(n5323), .Y(n5322) );
  OAI22X1 U2972 ( .A(n4691), .B(n5324), .C(n4598), .D(n5324), .Y(n5323) );
  OAI22X1 U2973 ( .A(n4689), .B(n4629), .C(n4553), .D(n4570), .Y(n5324) );
  XNOR2X1 U2974 ( .A(n5325), .B(n4599), .Y(n3480) );
  OAI21X1 U2975 ( .A(n4621), .B(n4734), .C(n5326), .Y(n5325) );
  OAI22X1 U2976 ( .A(n4571), .B(n5327), .C(n4598), .D(n5327), .Y(n5326) );
  OAI22X1 U2977 ( .A(n4572), .B(n4629), .C(n4553), .D(n4689), .Y(n5327) );
  XNOR2X1 U2978 ( .A(n5328), .B(n4599), .Y(n3479) );
  OAI21X1 U2979 ( .A(n4621), .B(n4733), .C(n5329), .Y(n5328) );
  OAI22X1 U2980 ( .A(n4687), .B(n5330), .C(n4598), .D(n5330), .Y(n5329) );
  OAI22X1 U2981 ( .A(n4685), .B(n4629), .C(n4553), .D(n4572), .Y(n5330) );
  XNOR2X1 U2982 ( .A(n5331), .B(n4599), .Y(n3478) );
  OAI21X1 U2983 ( .A(n4621), .B(n4731), .C(n5332), .Y(n5331) );
  OAI22X1 U2984 ( .A(n4573), .B(n5333), .C(n4598), .D(n5333), .Y(n5332) );
  OAI22X1 U2985 ( .A(n4574), .B(n4629), .C(n4553), .D(n4685), .Y(n5333) );
  XNOR2X1 U2986 ( .A(n5334), .B(n4599), .Y(n3477) );
  OAI21X1 U2987 ( .A(n4621), .B(n4730), .C(n5335), .Y(n5334) );
  OAI22X1 U2988 ( .A(n4683), .B(n5336), .C(n4598), .D(n5336), .Y(n5335) );
  OAI22X1 U2989 ( .A(n4680), .B(n4629), .C(n4553), .D(n4574), .Y(n5336) );
  XNOR2X1 U2990 ( .A(n5337), .B(n4599), .Y(n3476) );
  OAI21X1 U2991 ( .A(n4621), .B(n4729), .C(n5338), .Y(n5337) );
  OAI22X1 U2992 ( .A(n4575), .B(n5339), .C(n4598), .D(n5339), .Y(n5338) );
  OAI22X1 U2993 ( .A(n4576), .B(n4629), .C(n4553), .D(n4680), .Y(n5339) );
  XNOR2X1 U2994 ( .A(n5340), .B(n4599), .Y(n3475) );
  OAI21X1 U2995 ( .A(n4621), .B(n4727), .C(n5341), .Y(n5340) );
  OAI22X1 U2996 ( .A(n4678), .B(n5342), .C(n4598), .D(n5342), .Y(n5341) );
  OAI22X1 U2997 ( .A(n4676), .B(n4629), .C(n4553), .D(n4576), .Y(n5342) );
  XNOR2X1 U2998 ( .A(n5343), .B(n4599), .Y(n3474) );
  OAI21X1 U2999 ( .A(n4621), .B(n4726), .C(n5344), .Y(n5343) );
  OAI22X1 U3000 ( .A(n4577), .B(n5345), .C(n4598), .D(n5345), .Y(n5344) );
  OAI22X1 U3001 ( .A(n4578), .B(n4629), .C(n4553), .D(n4676), .Y(n5345) );
  XNOR2X1 U3002 ( .A(n5346), .B(n4599), .Y(n3473) );
  OAI21X1 U3003 ( .A(n4621), .B(n4725), .C(n5347), .Y(n5346) );
  OAI22X1 U3004 ( .A(n4674), .B(n5348), .C(n4598), .D(n5348), .Y(n5347) );
  OAI22X1 U3005 ( .A(n4671), .B(n4629), .C(n4553), .D(n4578), .Y(n5348) );
  XNOR2X1 U3006 ( .A(n5349), .B(n4599), .Y(n3472) );
  OAI21X1 U3007 ( .A(n4621), .B(n4724), .C(n5350), .Y(n5349) );
  OAI22X1 U3008 ( .A(n4579), .B(n5351), .C(n4598), .D(n5351), .Y(n5350) );
  OAI22X1 U3009 ( .A(n4580), .B(n4629), .C(n4553), .D(n4671), .Y(n5351) );
  XNOR2X1 U3010 ( .A(n5352), .B(n4599), .Y(n3471) );
  OAI21X1 U3011 ( .A(n4621), .B(n4722), .C(n5353), .Y(n5352) );
  OAI22X1 U3012 ( .A(n4669), .B(n5354), .C(n4598), .D(n5354), .Y(n5353) );
  OAI22X1 U3013 ( .A(n4666), .B(n4629), .C(n4553), .D(n4580), .Y(n5354) );
  XNOR2X1 U3014 ( .A(n5355), .B(n4599), .Y(n3470) );
  OAI21X1 U3015 ( .A(n4621), .B(n4721), .C(n5356), .Y(n5355) );
  OAI22X1 U3016 ( .A(n4581), .B(n5357), .C(n4598), .D(n5357), .Y(n5356) );
  OAI22X1 U3017 ( .A(n4582), .B(n4629), .C(n4553), .D(n4666), .Y(n5357) );
  XNOR2X1 U3018 ( .A(n5358), .B(n4599), .Y(n3469) );
  OAI21X1 U3019 ( .A(n4720), .B(n4621), .C(n5359), .Y(n5358) );
  OAI22X1 U3020 ( .A(n4664), .B(n5360), .C(n4598), .D(n5360), .Y(n5359) );
  OAI22X1 U3021 ( .A(n4662), .B(n4629), .C(n4582), .D(n4553), .Y(n5360) );
  XNOR2X1 U3022 ( .A(n5361), .B(n4599), .Y(n3468) );
  OAI21X1 U3023 ( .A(n4621), .B(n4719), .C(n5362), .Y(n5361) );
  OAI22X1 U3024 ( .A(n4583), .B(n5363), .C(n4598), .D(n5363), .Y(n5362) );
  OAI22X1 U3025 ( .A(n4584), .B(n4629), .C(n4662), .D(n4553), .Y(n5363) );
  XNOR2X1 U3026 ( .A(n5364), .B(n4599), .Y(n3467) );
  OAI21X1 U3027 ( .A(n4621), .B(n4718), .C(n5365), .Y(n5364) );
  OAI22X1 U3028 ( .A(n4660), .B(n5366), .C(n4598), .D(n5366), .Y(n5365) );
  OAI22X1 U3029 ( .A(n4657), .B(n4629), .C(n4553), .D(n4584), .Y(n5366) );
  XNOR2X1 U3030 ( .A(n5367), .B(n4599), .Y(n3466) );
  OAI21X1 U3031 ( .A(n4717), .B(n4621), .C(n5368), .Y(n5367) );
  OAI22X1 U3032 ( .A(n4585), .B(n5369), .C(n4598), .D(n5369), .Y(n5368) );
  OAI22X1 U3033 ( .A(n4586), .B(n4629), .C(n4657), .D(n4553), .Y(n5369) );
  XNOR2X1 U3034 ( .A(n5370), .B(n4599), .Y(n3465) );
  OAI21X1 U3035 ( .A(n4621), .B(n4716), .C(n5371), .Y(n5370) );
  OAI22X1 U3036 ( .A(n4656), .B(n5372), .C(n4598), .D(n5372), .Y(n5371) );
  OAI22X1 U3037 ( .A(n4654), .B(n4629), .C(n4586), .D(n4553), .Y(n5372) );
  XNOR2X1 U3038 ( .A(n5373), .B(n4599), .Y(n3464) );
  OAI21X1 U3039 ( .A(n4621), .B(n4715), .C(n5374), .Y(n5373) );
  OAI22X1 U3040 ( .A(n4587), .B(n5375), .C(n4598), .D(n5375), .Y(n5374) );
  OAI22X1 U3041 ( .A(n4588), .B(n4629), .C(n4553), .D(n4654), .Y(n5375) );
  XNOR2X1 U3042 ( .A(n5376), .B(n4599), .Y(n3463) );
  OAI21X1 U3043 ( .A(n4714), .B(n4621), .C(n5377), .Y(n5376) );
  OAI22X1 U3044 ( .A(n4652), .B(n5378), .C(n4598), .D(n5378), .Y(n5377) );
  OAI22X1 U3045 ( .A(n4650), .B(n4629), .C(n4588), .D(n4553), .Y(n5378) );
  XNOR2X1 U3046 ( .A(n5379), .B(n4600), .Y(n3462) );
  OAI21X1 U3047 ( .A(n4621), .B(n4713), .C(n5380), .Y(n5379) );
  OAI22X1 U3048 ( .A(n4589), .B(n5381), .C(n4598), .D(n5381), .Y(n5380) );
  OAI22X1 U3049 ( .A(n4590), .B(n4629), .C(n4650), .D(n4553), .Y(n5381) );
  XNOR2X1 U3050 ( .A(n5382), .B(n4600), .Y(n3461) );
  OAI21X1 U3051 ( .A(n4621), .B(n4712), .C(n5383), .Y(n5382) );
  OAI22X1 U3052 ( .A(n4649), .B(n5384), .C(n4598), .D(n5384), .Y(n5383) );
  OAI22X1 U3053 ( .A(n4647), .B(n4629), .C(n4553), .D(n4590), .Y(n5384) );
  XNOR2X1 U3054 ( .A(n5385), .B(n4600), .Y(n3460) );
  OAI21X1 U3055 ( .A(n4711), .B(n4621), .C(n5386), .Y(n5385) );
  OAI22X1 U3056 ( .A(n4591), .B(n5387), .C(n4598), .D(n5387), .Y(n5386) );
  OAI22X1 U3057 ( .A(n4710), .B(n4629), .C(n4647), .D(n4553), .Y(n5387) );
  XNOR2X1 U3058 ( .A(n5388), .B(n4600), .Y(n3459) );
  OAI21X1 U3059 ( .A(n4621), .B(n4709), .C(n5389), .Y(n5388) );
  OAI22X1 U3060 ( .A(n4646), .B(n5390), .C(n4598), .D(n5390), .Y(n5389) );
  OAI22X1 U3061 ( .A(n4644), .B(n4629), .C(n4710), .D(n4553), .Y(n5390) );
  XNOR2X1 U3062 ( .A(n5391), .B(n4600), .Y(n3458) );
  OAI21X1 U3063 ( .A(n4621), .B(n4708), .C(n5392), .Y(n5391) );
  OAI22X1 U3064 ( .A(b[26]), .B(n5393), .C(n4598), .D(n5393), .Y(n5392) );
  OAI22X1 U3065 ( .A(n4707), .B(n4629), .C(n4553), .D(n4644), .Y(n5393) );
  XNOR2X1 U3066 ( .A(n5394), .B(n4600), .Y(n3457) );
  OAI21X1 U3067 ( .A(n4706), .B(n4621), .C(n5395), .Y(n5394) );
  OAI22X1 U3068 ( .A(n4643), .B(n5396), .C(n4598), .D(n5396), .Y(n5395) );
  OAI22X1 U3069 ( .A(n4641), .B(n4629), .C(n4707), .D(n4553), .Y(n5396) );
  XNOR2X1 U3070 ( .A(n5397), .B(n4600), .Y(n3456) );
  OAI21X1 U3071 ( .A(n4621), .B(n4705), .C(n5398), .Y(n5397) );
  OAI22X1 U3072 ( .A(b[28]), .B(n5399), .C(n4598), .D(n5399), .Y(n5398) );
  OAI22X1 U3073 ( .A(n4641), .B(n4553), .C(n4704), .D(n4629), .Y(n5399) );
  XNOR2X1 U3074 ( .A(n5400), .B(n4600), .Y(n3455) );
  OAI21X1 U3075 ( .A(n4621), .B(n4703), .C(n5401), .Y(n5400) );
  OAI22X1 U3076 ( .A(b[29]), .B(n5402), .C(n4598), .D(n5402), .Y(n5401) );
  NAND3X1 U3077 ( .A(n5404), .B(n5405), .C(n5406), .Y(n5403) );
  OAI22X1 U3078 ( .A(n4553), .B(n4704), .C(n4632), .D(n4629), .Y(n5402) );
  XNOR2X1 U3079 ( .A(a[15]), .B(a[16]), .Y(n5404) );
  XNOR2X1 U3080 ( .A(a[16]), .B(n4600), .Y(n5405) );
  XOR2X1 U3081 ( .A(a[15]), .B(n4604), .Y(n5406) );
  XOR2X1 U3082 ( .A(n5407), .B(n4639), .Y(n3453) );
  OAI22X1 U3083 ( .A(n4595), .B(n4700), .C(n4622), .D(n4700), .Y(n5407) );
  XOR2X1 U3084 ( .A(n5408), .B(n4639), .Y(n3452) );
  OAI21X1 U3085 ( .A(n4622), .B(n4741), .C(n5409), .Y(n5408) );
  AOI22X1 U3086 ( .A(n4694), .B(n5410), .C(n4697), .D(n5411), .Y(n5409) );
  XOR2X1 U3087 ( .A(n5412), .B(n4639), .Y(n3451) );
  OAI21X1 U3088 ( .A(n4622), .B(n4738), .C(n5413), .Y(n5412) );
  OAI22X1 U3089 ( .A(n4699), .B(n5414), .C(n4596), .D(n5414), .Y(n5413) );
  OAI22X1 U3090 ( .A(n4597), .B(n4695), .C(n4595), .D(n4568), .Y(n5414) );
  XOR2X1 U3091 ( .A(n5415), .B(n4639), .Y(n3450) );
  OAI21X1 U3092 ( .A(n4622), .B(n4737), .C(n5416), .Y(n5415) );
  OAI22X1 U3093 ( .A(n4694), .B(n5417), .C(n4596), .D(n5417), .Y(n5416) );
  OAI22X1 U3094 ( .A(n4597), .B(n4568), .C(n4595), .D(n4693), .Y(n5417) );
  XOR2X1 U3095 ( .A(n5418), .B(n4639), .Y(n3449) );
  OAI21X1 U3096 ( .A(n4622), .B(n4736), .C(n5419), .Y(n5418) );
  OAI22X1 U3097 ( .A(n4569), .B(n5420), .C(n4596), .D(n5420), .Y(n5419) );
  OAI22X1 U3098 ( .A(n4597), .B(n4693), .C(n4595), .D(n4570), .Y(n5420) );
  XOR2X1 U3099 ( .A(n5421), .B(n4639), .Y(n3448) );
  OAI21X1 U3100 ( .A(n4622), .B(n4735), .C(n5422), .Y(n5421) );
  OAI22X1 U3101 ( .A(n4691), .B(n5423), .C(n4596), .D(n5423), .Y(n5422) );
  OAI22X1 U3102 ( .A(n4597), .B(n4570), .C(n4595), .D(n4689), .Y(n5423) );
  XOR2X1 U3103 ( .A(n5424), .B(n4639), .Y(n3447) );
  OAI21X1 U3104 ( .A(n4622), .B(n4734), .C(n5425), .Y(n5424) );
  OAI22X1 U3105 ( .A(n4571), .B(n5426), .C(n4596), .D(n5426), .Y(n5425) );
  OAI22X1 U3106 ( .A(n4597), .B(n4689), .C(n4595), .D(n4572), .Y(n5426) );
  XOR2X1 U3107 ( .A(n5427), .B(n4639), .Y(n3446) );
  OAI21X1 U3108 ( .A(n4622), .B(n4733), .C(n5428), .Y(n5427) );
  OAI22X1 U3109 ( .A(n4687), .B(n5429), .C(n4596), .D(n5429), .Y(n5428) );
  OAI22X1 U3110 ( .A(n4597), .B(n4572), .C(n4595), .D(n4685), .Y(n5429) );
  XOR2X1 U3111 ( .A(n5430), .B(n4639), .Y(n3445) );
  OAI21X1 U3112 ( .A(n4622), .B(n4731), .C(n5431), .Y(n5430) );
  OAI22X1 U3113 ( .A(n4573), .B(n5432), .C(n4596), .D(n5432), .Y(n5431) );
  OAI22X1 U3114 ( .A(n4597), .B(n4685), .C(n4595), .D(n4574), .Y(n5432) );
  XOR2X1 U3115 ( .A(n5433), .B(n4639), .Y(n3444) );
  OAI21X1 U3116 ( .A(n4622), .B(n4730), .C(n5434), .Y(n5433) );
  OAI22X1 U3117 ( .A(n4683), .B(n5435), .C(n4596), .D(n5435), .Y(n5434) );
  OAI22X1 U3118 ( .A(n4597), .B(n4574), .C(n4595), .D(n4680), .Y(n5435) );
  XOR2X1 U3119 ( .A(n5436), .B(n4639), .Y(n3443) );
  OAI21X1 U3120 ( .A(n4622), .B(n4729), .C(n5437), .Y(n5436) );
  OAI22X1 U3121 ( .A(n4575), .B(n5438), .C(n4596), .D(n5438), .Y(n5437) );
  OAI22X1 U3122 ( .A(n4597), .B(n4680), .C(n4595), .D(n4576), .Y(n5438) );
  XOR2X1 U3123 ( .A(n5439), .B(n4639), .Y(n3442) );
  OAI21X1 U3124 ( .A(n4622), .B(n4727), .C(n5440), .Y(n5439) );
  OAI22X1 U3125 ( .A(n4678), .B(n5441), .C(n4596), .D(n5441), .Y(n5440) );
  OAI22X1 U3126 ( .A(n4597), .B(n4576), .C(n4595), .D(n4676), .Y(n5441) );
  XOR2X1 U3127 ( .A(n5442), .B(n4639), .Y(n3441) );
  OAI21X1 U3128 ( .A(n4622), .B(n4726), .C(n5443), .Y(n5442) );
  OAI22X1 U3129 ( .A(n4577), .B(n5444), .C(n4596), .D(n5444), .Y(n5443) );
  OAI22X1 U3130 ( .A(n4597), .B(n4676), .C(n4595), .D(n4578), .Y(n5444) );
  XOR2X1 U3131 ( .A(n5445), .B(n4639), .Y(n3440) );
  OAI21X1 U3132 ( .A(n4622), .B(n4725), .C(n5446), .Y(n5445) );
  OAI22X1 U3133 ( .A(n4674), .B(n5447), .C(n4596), .D(n5447), .Y(n5446) );
  OAI22X1 U3134 ( .A(n4597), .B(n4578), .C(n4595), .D(n4671), .Y(n5447) );
  XOR2X1 U3135 ( .A(n5448), .B(n4639), .Y(n3439) );
  OAI21X1 U3136 ( .A(n4622), .B(n4724), .C(n5449), .Y(n5448) );
  OAI22X1 U3137 ( .A(n4579), .B(n5450), .C(n4596), .D(n5450), .Y(n5449) );
  OAI22X1 U3138 ( .A(n4597), .B(n4671), .C(n4595), .D(n4580), .Y(n5450) );
  XOR2X1 U3139 ( .A(n5451), .B(n4639), .Y(n3438) );
  OAI21X1 U3140 ( .A(n4622), .B(n4722), .C(n5452), .Y(n5451) );
  OAI22X1 U3141 ( .A(n4669), .B(n5453), .C(n4596), .D(n5453), .Y(n5452) );
  OAI22X1 U3142 ( .A(n4595), .B(n4666), .C(n4597), .D(n4580), .Y(n5453) );
  XOR2X1 U3143 ( .A(n5454), .B(n4639), .Y(n3437) );
  OAI21X1 U3144 ( .A(n4622), .B(n4721), .C(n5455), .Y(n5454) );
  OAI22X1 U3145 ( .A(n4581), .B(n5456), .C(n4596), .D(n5456), .Y(n5455) );
  OAI22X1 U3146 ( .A(n4597), .B(n4666), .C(n4595), .D(n4582), .Y(n5456) );
  XOR2X1 U3147 ( .A(n5457), .B(n4639), .Y(n3436) );
  OAI21X1 U3148 ( .A(n4622), .B(n4720), .C(n5458), .Y(n5457) );
  OAI22X1 U3149 ( .A(n4664), .B(n5459), .C(n4596), .D(n5459), .Y(n5458) );
  OAI22X1 U3150 ( .A(n4595), .B(n4662), .C(n4597), .D(n4582), .Y(n5459) );
  XOR2X1 U3151 ( .A(n5460), .B(n4639), .Y(n3435) );
  OAI21X1 U3152 ( .A(n4622), .B(n4719), .C(n5461), .Y(n5460) );
  OAI22X1 U3153 ( .A(n4583), .B(n5462), .C(n4596), .D(n5462), .Y(n5461) );
  OAI22X1 U3154 ( .A(n4597), .B(n4662), .C(n4595), .D(n4584), .Y(n5462) );
  XOR2X1 U3155 ( .A(n5463), .B(n4639), .Y(n3434) );
  OAI21X1 U3156 ( .A(n4622), .B(n4718), .C(n5464), .Y(n5463) );
  OAI22X1 U3157 ( .A(n4660), .B(n5465), .C(n4596), .D(n5465), .Y(n5464) );
  OAI22X1 U3158 ( .A(n4597), .B(n4584), .C(n4595), .D(n4657), .Y(n5465) );
  XOR2X1 U3159 ( .A(n5466), .B(n2150), .Y(n3433) );
  OAI21X1 U3160 ( .A(n4622), .B(n4717), .C(n5467), .Y(n5466) );
  OAI22X1 U3161 ( .A(n4585), .B(n5468), .C(n4596), .D(n5468), .Y(n5467) );
  OAI22X1 U3162 ( .A(n4595), .B(n4586), .C(n4597), .D(n4657), .Y(n5468) );
  XOR2X1 U3163 ( .A(n5469), .B(n2150), .Y(n3432) );
  OAI21X1 U3164 ( .A(n4622), .B(n4716), .C(n5470), .Y(n5469) );
  OAI22X1 U3165 ( .A(n4655), .B(n5471), .C(n4596), .D(n5471), .Y(n5470) );
  OAI22X1 U3166 ( .A(n4597), .B(n4586), .C(n4595), .D(n4654), .Y(n5471) );
  XOR2X1 U3167 ( .A(n5472), .B(n2150), .Y(n3431) );
  OAI21X1 U3168 ( .A(n4622), .B(n4715), .C(n5473), .Y(n5472) );
  OAI22X1 U3169 ( .A(n4587), .B(n5474), .C(n4596), .D(n5474), .Y(n5473) );
  OAI22X1 U3170 ( .A(n4597), .B(n4654), .C(n4595), .D(n4588), .Y(n5474) );
  XOR2X1 U3171 ( .A(n5475), .B(n2150), .Y(n3430) );
  OAI21X1 U3172 ( .A(n4622), .B(n4714), .C(n5476), .Y(n5475) );
  OAI22X1 U3173 ( .A(n4653), .B(n5477), .C(n4596), .D(n5477), .Y(n5476) );
  OAI22X1 U3174 ( .A(n4595), .B(n4650), .C(n4597), .D(n4588), .Y(n5477) );
  XOR2X1 U3175 ( .A(n5478), .B(n2150), .Y(n3429) );
  OAI21X1 U3176 ( .A(n4622), .B(n4713), .C(n5479), .Y(n5478) );
  OAI22X1 U3177 ( .A(n4589), .B(n5480), .C(n4596), .D(n5480), .Y(n5479) );
  OAI22X1 U3178 ( .A(n4597), .B(n4650), .C(n4595), .D(n4590), .Y(n5480) );
  XOR2X1 U3179 ( .A(n5481), .B(n2150), .Y(n3428) );
  OAI21X1 U3180 ( .A(n4622), .B(n4712), .C(n5482), .Y(n5481) );
  OAI22X1 U3181 ( .A(n4649), .B(n5483), .C(n4596), .D(n5483), .Y(n5482) );
  OAI22X1 U3182 ( .A(n4597), .B(n4590), .C(n4595), .D(n4647), .Y(n5483) );
  XOR2X1 U3183 ( .A(n5484), .B(n2150), .Y(n3427) );
  OAI21X1 U3184 ( .A(n4622), .B(n4711), .C(n5485), .Y(n5484) );
  OAI22X1 U3185 ( .A(n4591), .B(n5486), .C(n4596), .D(n5486), .Y(n5485) );
  OAI22X1 U3186 ( .A(n4595), .B(n4710), .C(n4597), .D(n4647), .Y(n5486) );
  XOR2X1 U3187 ( .A(n5487), .B(n2150), .Y(n3426) );
  OAI21X1 U3188 ( .A(n4622), .B(n4709), .C(n5488), .Y(n5487) );
  OAI22X1 U3189 ( .A(n4646), .B(n5489), .C(n4596), .D(n5489), .Y(n5488) );
  OAI22X1 U3190 ( .A(n4597), .B(n4710), .C(n4595), .D(n4644), .Y(n5489) );
  XOR2X1 U3191 ( .A(n5490), .B(n2150), .Y(n3425) );
  OAI21X1 U3192 ( .A(n4622), .B(n4708), .C(n5491), .Y(n5490) );
  OAI22X1 U3193 ( .A(b[26]), .B(n5492), .C(n4596), .D(n5492), .Y(n5491) );
  NAND3X1 U3194 ( .A(n5494), .B(n5495), .C(n5496), .Y(n5493) );
  OAI22X1 U3195 ( .A(n4597), .B(n4644), .C(n4707), .D(n4595), .Y(n5492) );
  NOR2X1 U3196 ( .A(n5495), .B(n5494), .Y(n5410) );
  NOR2X1 U3197 ( .A(n4754), .B(n5496), .Y(n5411) );
  XNOR2X1 U3198 ( .A(a[18]), .B(a[19]), .Y(n5496) );
  XOR2X1 U3199 ( .A(a[19]), .B(n2150), .Y(n5495) );
  XOR2X1 U3200 ( .A(a[18]), .B(n4600), .Y(n5494) );
  XOR2X1 U3201 ( .A(n4637), .B(n5497), .Y(n3423) );
  OAI22X1 U3202 ( .A(n4700), .B(n4554), .C(n4700), .D(n4592), .Y(n5497) );
  XOR2X1 U3203 ( .A(n5498), .B(n2153), .Y(n3422) );
  OAI21X1 U3204 ( .A(n4554), .B(n4741), .C(n5499), .Y(n5498) );
  AOI22X1 U3205 ( .A(n4694), .B(n5500), .C(n4697), .D(n5501), .Y(n5499) );
  XOR2X1 U3206 ( .A(n5502), .B(n2153), .Y(n3421) );
  OAI21X1 U3207 ( .A(n4554), .B(n4738), .C(n5503), .Y(n5502) );
  OAI22X1 U3208 ( .A(n4699), .B(n5504), .C(n4593), .D(n5504), .Y(n5503) );
  OAI22X1 U3209 ( .A(n4594), .B(n4695), .C(n4592), .D(n4568), .Y(n5504) );
  XOR2X1 U3210 ( .A(n5505), .B(n2153), .Y(n3420) );
  OAI21X1 U3211 ( .A(n4554), .B(n4737), .C(n5506), .Y(n5505) );
  OAI22X1 U3212 ( .A(n4694), .B(n5507), .C(n4593), .D(n5507), .Y(n5506) );
  OAI22X1 U3213 ( .A(n4594), .B(n4568), .C(n4592), .D(n4693), .Y(n5507) );
  XOR2X1 U3214 ( .A(n5508), .B(n2153), .Y(n3419) );
  OAI21X1 U3215 ( .A(n4554), .B(n4736), .C(n5509), .Y(n5508) );
  OAI22X1 U3216 ( .A(n4569), .B(n5510), .C(n4593), .D(n5510), .Y(n5509) );
  OAI22X1 U3217 ( .A(n4594), .B(n4693), .C(n4592), .D(n4570), .Y(n5510) );
  XOR2X1 U3218 ( .A(n5511), .B(n2153), .Y(n3418) );
  OAI21X1 U3219 ( .A(n4554), .B(n4735), .C(n5512), .Y(n5511) );
  OAI22X1 U3220 ( .A(n4691), .B(n5513), .C(n4593), .D(n5513), .Y(n5512) );
  OAI22X1 U3221 ( .A(n4594), .B(n4570), .C(n4592), .D(n4689), .Y(n5513) );
  XOR2X1 U3222 ( .A(n5514), .B(n2153), .Y(n3417) );
  OAI21X1 U3223 ( .A(n4554), .B(n4734), .C(n5515), .Y(n5514) );
  OAI22X1 U3224 ( .A(n4571), .B(n5516), .C(n4593), .D(n5516), .Y(n5515) );
  OAI22X1 U3225 ( .A(n4594), .B(n4689), .C(n4592), .D(n4572), .Y(n5516) );
  XOR2X1 U3226 ( .A(n5517), .B(n2153), .Y(n3416) );
  OAI21X1 U3227 ( .A(n4554), .B(n4733), .C(n5518), .Y(n5517) );
  OAI22X1 U3228 ( .A(n4687), .B(n5519), .C(n4593), .D(n5519), .Y(n5518) );
  OAI22X1 U3229 ( .A(n4594), .B(n4572), .C(n4592), .D(n4685), .Y(n5519) );
  XOR2X1 U3230 ( .A(n5520), .B(n2153), .Y(n3415) );
  OAI21X1 U3231 ( .A(n4554), .B(n4731), .C(n5521), .Y(n5520) );
  OAI22X1 U3232 ( .A(n4573), .B(n5522), .C(n4593), .D(n5522), .Y(n5521) );
  OAI22X1 U3233 ( .A(n4594), .B(n4685), .C(n4592), .D(n4574), .Y(n5522) );
  XOR2X1 U3234 ( .A(n5523), .B(n2153), .Y(n3414) );
  OAI21X1 U3235 ( .A(n4554), .B(n4730), .C(n5524), .Y(n5523) );
  OAI22X1 U3236 ( .A(n4683), .B(n5525), .C(n4593), .D(n5525), .Y(n5524) );
  OAI22X1 U3237 ( .A(n4594), .B(n4574), .C(n4592), .D(n4680), .Y(n5525) );
  XOR2X1 U3238 ( .A(n5526), .B(n2153), .Y(n3413) );
  OAI21X1 U3239 ( .A(n4554), .B(n4729), .C(n5527), .Y(n5526) );
  OAI22X1 U3240 ( .A(n4575), .B(n5528), .C(n4593), .D(n5528), .Y(n5527) );
  OAI22X1 U3241 ( .A(n4594), .B(n4680), .C(n4592), .D(n4576), .Y(n5528) );
  XOR2X1 U3242 ( .A(n5529), .B(n2153), .Y(n3412) );
  OAI21X1 U3243 ( .A(n4554), .B(n4727), .C(n5530), .Y(n5529) );
  OAI22X1 U3244 ( .A(n4678), .B(n5531), .C(n4593), .D(n5531), .Y(n5530) );
  OAI22X1 U3245 ( .A(n4594), .B(n4576), .C(n4592), .D(n4676), .Y(n5531) );
  XOR2X1 U3246 ( .A(n5532), .B(n2153), .Y(n3411) );
  OAI21X1 U3247 ( .A(n4554), .B(n4726), .C(n5533), .Y(n5532) );
  OAI22X1 U3248 ( .A(n4577), .B(n5534), .C(n4593), .D(n5534), .Y(n5533) );
  OAI22X1 U3249 ( .A(n4594), .B(n4676), .C(n4592), .D(n4578), .Y(n5534) );
  XOR2X1 U3250 ( .A(n5535), .B(n2153), .Y(n3410) );
  OAI21X1 U3251 ( .A(n4554), .B(n4725), .C(n5536), .Y(n5535) );
  OAI22X1 U3252 ( .A(n4674), .B(n5537), .C(n4593), .D(n5537), .Y(n5536) );
  OAI22X1 U3253 ( .A(n4594), .B(n4578), .C(n4592), .D(n4671), .Y(n5537) );
  XOR2X1 U3254 ( .A(n5538), .B(n4637), .Y(n3409) );
  OAI21X1 U3255 ( .A(n4554), .B(n4724), .C(n5539), .Y(n5538) );
  OAI22X1 U3256 ( .A(n4579), .B(n5540), .C(n4593), .D(n5540), .Y(n5539) );
  OAI22X1 U3257 ( .A(n4594), .B(n4671), .C(n4592), .D(n4580), .Y(n5540) );
  XOR2X1 U3258 ( .A(n5541), .B(n4637), .Y(n3408) );
  OAI21X1 U3259 ( .A(n4554), .B(n4722), .C(n5542), .Y(n5541) );
  OAI22X1 U3260 ( .A(n4669), .B(n5543), .C(n4593), .D(n5543), .Y(n5542) );
  OAI22X1 U3261 ( .A(n4592), .B(n4666), .C(n4594), .D(n4580), .Y(n5543) );
  XOR2X1 U3262 ( .A(n5544), .B(n4637), .Y(n3407) );
  OAI21X1 U3263 ( .A(n4554), .B(n4721), .C(n5545), .Y(n5544) );
  OAI22X1 U3264 ( .A(n4581), .B(n5546), .C(n4593), .D(n5546), .Y(n5545) );
  OAI22X1 U3265 ( .A(n4594), .B(n4666), .C(n4592), .D(n4582), .Y(n5546) );
  XOR2X1 U3266 ( .A(n5547), .B(n4637), .Y(n3406) );
  OAI21X1 U3267 ( .A(n4554), .B(n4720), .C(n5548), .Y(n5547) );
  OAI22X1 U3268 ( .A(n4664), .B(n5549), .C(n4593), .D(n5549), .Y(n5548) );
  OAI22X1 U3269 ( .A(n4592), .B(n4662), .C(n4594), .D(n4582), .Y(n5549) );
  XOR2X1 U3270 ( .A(n5550), .B(n4637), .Y(n3405) );
  OAI21X1 U3271 ( .A(n4554), .B(n4719), .C(n5551), .Y(n5550) );
  OAI22X1 U3272 ( .A(n4583), .B(n5552), .C(n4593), .D(n5552), .Y(n5551) );
  OAI22X1 U3273 ( .A(n4594), .B(n4662), .C(n4592), .D(n4584), .Y(n5552) );
  XOR2X1 U3274 ( .A(n5553), .B(n4637), .Y(n3404) );
  OAI21X1 U3275 ( .A(n4554), .B(n4718), .C(n5554), .Y(n5553) );
  OAI22X1 U3276 ( .A(n4660), .B(n5555), .C(n4593), .D(n5555), .Y(n5554) );
  OAI22X1 U3277 ( .A(n4594), .B(n4584), .C(n4592), .D(n4657), .Y(n5555) );
  XOR2X1 U3278 ( .A(n5556), .B(n4637), .Y(n3403) );
  OAI21X1 U3279 ( .A(n4554), .B(n4717), .C(n5557), .Y(n5556) );
  OAI22X1 U3280 ( .A(n4585), .B(n5558), .C(n4593), .D(n5558), .Y(n5557) );
  OAI22X1 U3281 ( .A(n4592), .B(n4586), .C(n4594), .D(n4657), .Y(n5558) );
  XOR2X1 U3282 ( .A(n5559), .B(n4637), .Y(n3402) );
  OAI21X1 U3283 ( .A(n4554), .B(n4716), .C(n5560), .Y(n5559) );
  OAI22X1 U3284 ( .A(n4656), .B(n5561), .C(n4593), .D(n5561), .Y(n5560) );
  OAI22X1 U3285 ( .A(n4594), .B(n4586), .C(n4592), .D(n4654), .Y(n5561) );
  XOR2X1 U3286 ( .A(n5562), .B(n4637), .Y(n3401) );
  OAI21X1 U3287 ( .A(n4554), .B(n4715), .C(n5563), .Y(n5562) );
  OAI22X1 U3288 ( .A(n4587), .B(n5564), .C(n4593), .D(n5564), .Y(n5563) );
  OAI22X1 U3289 ( .A(n4594), .B(n4654), .C(n4592), .D(n4588), .Y(n5564) );
  XOR2X1 U3290 ( .A(n5565), .B(n4637), .Y(n3400) );
  OAI21X1 U3291 ( .A(n4554), .B(n4714), .C(n5566), .Y(n5565) );
  OAI22X1 U3292 ( .A(n4653), .B(n5567), .C(n4593), .D(n5567), .Y(n5566) );
  OAI22X1 U3293 ( .A(n4592), .B(n4650), .C(n4594), .D(n4588), .Y(n5567) );
  XOR2X1 U3294 ( .A(n5568), .B(n4637), .Y(n3399) );
  OAI21X1 U3295 ( .A(n4554), .B(n4713), .C(n5569), .Y(n5568) );
  OAI22X1 U3296 ( .A(n4589), .B(n5570), .C(n4593), .D(n5570), .Y(n5569) );
  OAI22X1 U3297 ( .A(n4594), .B(n4650), .C(n4592), .D(n4590), .Y(n5570) );
  XOR2X1 U3298 ( .A(n5571), .B(n4637), .Y(n3398) );
  OAI21X1 U3299 ( .A(n4554), .B(n4712), .C(n5572), .Y(n5571) );
  OAI22X1 U3300 ( .A(n4649), .B(n5573), .C(n4593), .D(n5573), .Y(n5572) );
  NAND3X1 U3301 ( .A(n4753), .B(n5575), .C(n5576), .Y(n5574) );
  OAI22X1 U3302 ( .A(n4594), .B(n4590), .C(n4647), .D(n4592), .Y(n5573) );
  NOR2X1 U3303 ( .A(n5575), .B(n4753), .Y(n5500) );
  NOR2X1 U3304 ( .A(n5577), .B(n5576), .Y(n5501) );
  XNOR2X1 U3305 ( .A(a[21]), .B(a[22]), .Y(n5576) );
  XOR2X1 U3306 ( .A(a[22]), .B(n4637), .Y(n5575) );
  XOR2X1 U3307 ( .A(a[21]), .B(n2150), .Y(n5577) );
  XOR2X1 U3308 ( .A(n4635), .B(n5578), .Y(n3396) );
  OAI22X1 U3309 ( .A(n4700), .B(n4556), .C(n4700), .D(n4750), .Y(n5578) );
  XOR2X1 U3310 ( .A(n5579), .B(n2156), .Y(n3395) );
  OAI21X1 U3311 ( .A(n4556), .B(n4741), .C(n5580), .Y(n5579) );
  AOI22X1 U3312 ( .A(n4694), .B(n5581), .C(n4697), .D(n5582), .Y(n5580) );
  XOR2X1 U3313 ( .A(n5583), .B(n2156), .Y(n3394) );
  OAI21X1 U3314 ( .A(n4556), .B(n4738), .C(n5584), .Y(n5583) );
  OAI22X1 U3315 ( .A(n4699), .B(n5585), .C(n4567), .D(n5585), .Y(n5584) );
  OAI22X1 U3316 ( .A(n4751), .B(n4695), .C(n4750), .D(n4568), .Y(n5585) );
  XOR2X1 U3317 ( .A(n5586), .B(n2156), .Y(n3393) );
  OAI21X1 U3318 ( .A(n4556), .B(n4737), .C(n5587), .Y(n5586) );
  OAI22X1 U3319 ( .A(n4694), .B(n5588), .C(n4567), .D(n5588), .Y(n5587) );
  OAI22X1 U3320 ( .A(n4751), .B(n4568), .C(n4750), .D(n4693), .Y(n5588) );
  XOR2X1 U3321 ( .A(n5589), .B(n2156), .Y(n3392) );
  OAI21X1 U3322 ( .A(n4556), .B(n4736), .C(n5590), .Y(n5589) );
  OAI22X1 U3323 ( .A(n4569), .B(n5591), .C(n4567), .D(n5591), .Y(n5590) );
  OAI22X1 U3324 ( .A(n4751), .B(n4693), .C(n4750), .D(n4570), .Y(n5591) );
  XOR2X1 U3325 ( .A(n5592), .B(n2156), .Y(n3391) );
  OAI21X1 U3326 ( .A(n4556), .B(n4735), .C(n5593), .Y(n5592) );
  OAI22X1 U3327 ( .A(n4691), .B(n5594), .C(n4567), .D(n5594), .Y(n5593) );
  OAI22X1 U3328 ( .A(n4751), .B(n4570), .C(n4750), .D(n4689), .Y(n5594) );
  XOR2X1 U3329 ( .A(n5595), .B(n2156), .Y(n3390) );
  OAI21X1 U3330 ( .A(n4556), .B(n4734), .C(n5596), .Y(n5595) );
  OAI22X1 U3331 ( .A(n4571), .B(n5597), .C(n4567), .D(n5597), .Y(n5596) );
  OAI22X1 U3332 ( .A(n4751), .B(n4689), .C(n4750), .D(n4572), .Y(n5597) );
  XOR2X1 U3333 ( .A(n5598), .B(n2156), .Y(n3389) );
  OAI21X1 U3334 ( .A(n4556), .B(n4733), .C(n5599), .Y(n5598) );
  OAI22X1 U3335 ( .A(n4687), .B(n5600), .C(n4567), .D(n5600), .Y(n5599) );
  OAI22X1 U3336 ( .A(n4751), .B(n4572), .C(n4750), .D(n4685), .Y(n5600) );
  XOR2X1 U3337 ( .A(n5601), .B(n2156), .Y(n3388) );
  OAI21X1 U3338 ( .A(n4556), .B(n4731), .C(n5602), .Y(n5601) );
  OAI22X1 U3339 ( .A(n4573), .B(n5603), .C(n4567), .D(n5603), .Y(n5602) );
  OAI22X1 U3340 ( .A(n4751), .B(n4685), .C(n4750), .D(n4574), .Y(n5603) );
  XOR2X1 U3341 ( .A(n5604), .B(n2156), .Y(n3387) );
  OAI21X1 U3342 ( .A(n4556), .B(n4730), .C(n5605), .Y(n5604) );
  OAI22X1 U3343 ( .A(n4683), .B(n5606), .C(n4567), .D(n5606), .Y(n5605) );
  OAI22X1 U3344 ( .A(n4751), .B(n4574), .C(n4750), .D(n4680), .Y(n5606) );
  XOR2X1 U3345 ( .A(n5607), .B(n2156), .Y(n3386) );
  OAI21X1 U3346 ( .A(n4556), .B(n4729), .C(n5608), .Y(n5607) );
  OAI22X1 U3347 ( .A(n4575), .B(n5609), .C(n4567), .D(n5609), .Y(n5608) );
  OAI22X1 U3348 ( .A(n4751), .B(n4680), .C(n4750), .D(n4576), .Y(n5609) );
  XOR2X1 U3349 ( .A(n5610), .B(n4635), .Y(n3385) );
  OAI21X1 U3350 ( .A(n4556), .B(n4727), .C(n5611), .Y(n5610) );
  OAI22X1 U3351 ( .A(n4678), .B(n5612), .C(n4567), .D(n5612), .Y(n5611) );
  OAI22X1 U3352 ( .A(n4751), .B(n4576), .C(n4750), .D(n4676), .Y(n5612) );
  XOR2X1 U3353 ( .A(n5613), .B(n4635), .Y(n3384) );
  OAI21X1 U3354 ( .A(n4556), .B(n4726), .C(n5614), .Y(n5613) );
  OAI22X1 U3355 ( .A(n4577), .B(n5615), .C(n4567), .D(n5615), .Y(n5614) );
  OAI22X1 U3356 ( .A(n4751), .B(n4676), .C(n4750), .D(n4578), .Y(n5615) );
  XOR2X1 U3357 ( .A(n5616), .B(n4635), .Y(n3383) );
  OAI21X1 U3358 ( .A(n4556), .B(n4725), .C(n5617), .Y(n5616) );
  OAI22X1 U3359 ( .A(n4674), .B(n5618), .C(n4567), .D(n5618), .Y(n5617) );
  OAI22X1 U3360 ( .A(n4751), .B(n4578), .C(n4750), .D(n4671), .Y(n5618) );
  XOR2X1 U3361 ( .A(n5619), .B(n4635), .Y(n3382) );
  OAI21X1 U3362 ( .A(n4556), .B(n4724), .C(n5620), .Y(n5619) );
  OAI22X1 U3363 ( .A(n4579), .B(n5621), .C(n4567), .D(n5621), .Y(n5620) );
  OAI22X1 U3364 ( .A(n4751), .B(n4671), .C(n4750), .D(n4580), .Y(n5621) );
  XOR2X1 U3365 ( .A(n5622), .B(n4635), .Y(n3381) );
  OAI21X1 U3366 ( .A(n4556), .B(n4722), .C(n5623), .Y(n5622) );
  OAI22X1 U3367 ( .A(n4669), .B(n5624), .C(n4567), .D(n5624), .Y(n5623) );
  OAI22X1 U3368 ( .A(n4750), .B(n4666), .C(n4751), .D(n4580), .Y(n5624) );
  XOR2X1 U3369 ( .A(n5625), .B(n4635), .Y(n3380) );
  OAI21X1 U3370 ( .A(n4556), .B(n4721), .C(n5626), .Y(n5625) );
  OAI22X1 U3371 ( .A(n4581), .B(n5627), .C(n4567), .D(n5627), .Y(n5626) );
  OAI22X1 U3372 ( .A(n4751), .B(n4666), .C(n4750), .D(n4582), .Y(n5627) );
  XOR2X1 U3373 ( .A(n5628), .B(n4635), .Y(n3379) );
  OAI21X1 U3374 ( .A(n4556), .B(n4720), .C(n5629), .Y(n5628) );
  OAI22X1 U3375 ( .A(n4665), .B(n5630), .C(n4567), .D(n5630), .Y(n5629) );
  OAI22X1 U3376 ( .A(n4750), .B(n4662), .C(n4751), .D(n4582), .Y(n5630) );
  XOR2X1 U3377 ( .A(n5631), .B(n2156), .Y(n3378) );
  OAI21X1 U3378 ( .A(n4556), .B(n4719), .C(n5632), .Y(n5631) );
  OAI22X1 U3379 ( .A(n4583), .B(n5633), .C(n4567), .D(n5633), .Y(n5632) );
  OAI22X1 U3380 ( .A(n4751), .B(n4662), .C(n4750), .D(n4584), .Y(n5633) );
  XOR2X1 U3381 ( .A(n5634), .B(n4635), .Y(n3377) );
  OAI21X1 U3382 ( .A(n4556), .B(n4718), .C(n5635), .Y(n5634) );
  OAI22X1 U3383 ( .A(n4661), .B(n5636), .C(n4567), .D(n5636), .Y(n5635) );
  OAI22X1 U3384 ( .A(n4751), .B(n4584), .C(n4750), .D(n4657), .Y(n5636) );
  XOR2X1 U3385 ( .A(n5637), .B(n4635), .Y(n3376) );
  OAI21X1 U3386 ( .A(n4556), .B(n4717), .C(n5638), .Y(n5637) );
  OAI22X1 U3387 ( .A(n4585), .B(n5639), .C(n4567), .D(n5639), .Y(n5638) );
  OAI22X1 U3388 ( .A(n4750), .B(n4586), .C(n4751), .D(n4657), .Y(n5639) );
  XOR2X1 U3389 ( .A(n5640), .B(n4635), .Y(n3375) );
  OAI21X1 U3390 ( .A(n4556), .B(n4716), .C(n5641), .Y(n5640) );
  OAI22X1 U3391 ( .A(n4656), .B(n5642), .C(n4567), .D(n5642), .Y(n5641) );
  OAI22X1 U3392 ( .A(n4751), .B(n4586), .C(n4750), .D(n4654), .Y(n5642) );
  XOR2X1 U3393 ( .A(n5643), .B(n4635), .Y(n3374) );
  OAI21X1 U3394 ( .A(n4556), .B(n4715), .C(n5644), .Y(n5643) );
  OAI22X1 U3395 ( .A(n4587), .B(n5645), .C(n4567), .D(n5645), .Y(n5644) );
  NAND3X1 U3396 ( .A(n5647), .B(n5648), .C(n5649), .Y(n5646) );
  OAI22X1 U3397 ( .A(n4751), .B(n4654), .C(n4588), .D(n4750), .Y(n5645) );
  NOR2X1 U3398 ( .A(n5648), .B(n5647), .Y(n5581) );
  NOR2X1 U3399 ( .A(n4752), .B(n5649), .Y(n5582) );
  XNOR2X1 U3400 ( .A(a[24]), .B(a[25]), .Y(n5649) );
  XOR2X1 U3401 ( .A(a[25]), .B(n4635), .Y(n5648) );
  XNOR2X1 U3402 ( .A(a[24]), .B(n4637), .Y(n5647) );
  XOR2X1 U3403 ( .A(n4633), .B(n5650), .Y(n3372) );
  OAI22X1 U3404 ( .A(n4700), .B(n4555), .C(n4700), .D(n4746), .Y(n5650) );
  XOR2X1 U3405 ( .A(n5651), .B(n2159), .Y(n3371) );
  OAI21X1 U3406 ( .A(n4555), .B(n4741), .C(n5652), .Y(n5651) );
  AOI22X1 U3407 ( .A(n4694), .B(n5653), .C(n4696), .D(n5654), .Y(n5652) );
  XOR2X1 U3408 ( .A(n5655), .B(n2159), .Y(n3370) );
  OAI21X1 U3409 ( .A(n4555), .B(n4738), .C(n5656), .Y(n5655) );
  OAI22X1 U3410 ( .A(n4699), .B(n5657), .C(n4747), .D(n5657), .Y(n5656) );
  OAI22X1 U3411 ( .A(n4748), .B(n4695), .C(n4746), .D(n4568), .Y(n5657) );
  XOR2X1 U3412 ( .A(n5658), .B(n2159), .Y(n3369) );
  OAI21X1 U3413 ( .A(n4555), .B(n4737), .C(n5659), .Y(n5658) );
  OAI22X1 U3414 ( .A(n4694), .B(n5660), .C(n4747), .D(n5660), .Y(n5659) );
  OAI22X1 U3415 ( .A(n4748), .B(n4568), .C(n4746), .D(n4693), .Y(n5660) );
  XOR2X1 U3416 ( .A(n5661), .B(n2159), .Y(n3368) );
  OAI21X1 U3417 ( .A(n4555), .B(n4736), .C(n5662), .Y(n5661) );
  OAI22X1 U3418 ( .A(n4569), .B(n5663), .C(n4747), .D(n5663), .Y(n5662) );
  OAI22X1 U3419 ( .A(n4748), .B(n4693), .C(n4746), .D(n4570), .Y(n5663) );
  XOR2X1 U3420 ( .A(n5664), .B(n2159), .Y(n3367) );
  OAI21X1 U3421 ( .A(n4555), .B(n4735), .C(n5665), .Y(n5664) );
  OAI22X1 U3422 ( .A(n4692), .B(n5666), .C(n4747), .D(n5666), .Y(n5665) );
  OAI22X1 U3423 ( .A(n4748), .B(n4570), .C(n4746), .D(n4689), .Y(n5666) );
  XOR2X1 U3424 ( .A(n5667), .B(n2159), .Y(n3366) );
  OAI21X1 U3425 ( .A(n4555), .B(n4734), .C(n5668), .Y(n5667) );
  OAI22X1 U3426 ( .A(n4571), .B(n5669), .C(n4747), .D(n5669), .Y(n5668) );
  OAI22X1 U3427 ( .A(n4748), .B(n4689), .C(n4746), .D(n4572), .Y(n5669) );
  XOR2X1 U3428 ( .A(n5670), .B(n2159), .Y(n3365) );
  OAI21X1 U3429 ( .A(n4555), .B(n4733), .C(n5671), .Y(n5670) );
  OAI22X1 U3430 ( .A(n4688), .B(n5672), .C(n4747), .D(n5672), .Y(n5671) );
  OAI22X1 U3431 ( .A(n4748), .B(n4572), .C(n4746), .D(n4685), .Y(n5672) );
  XOR2X1 U3432 ( .A(n5673), .B(n2159), .Y(n3364) );
  OAI21X1 U3433 ( .A(n4555), .B(n4731), .C(n5674), .Y(n5673) );
  OAI22X1 U3434 ( .A(n4573), .B(n5675), .C(n4747), .D(n5675), .Y(n5674) );
  OAI22X1 U3435 ( .A(n4748), .B(n4685), .C(n4746), .D(n4574), .Y(n5675) );
  XOR2X1 U3436 ( .A(n5676), .B(n4633), .Y(n3363) );
  OAI21X1 U3437 ( .A(n4555), .B(n4730), .C(n5677), .Y(n5676) );
  OAI22X1 U3438 ( .A(n4684), .B(n5678), .C(n4747), .D(n5678), .Y(n5677) );
  OAI22X1 U3439 ( .A(n4748), .B(n4574), .C(n4746), .D(n4680), .Y(n5678) );
  XOR2X1 U3440 ( .A(n5679), .B(n4633), .Y(n3362) );
  OAI21X1 U3441 ( .A(n4555), .B(n4729), .C(n5680), .Y(n5679) );
  OAI22X1 U3442 ( .A(n4575), .B(n5681), .C(n4747), .D(n5681), .Y(n5680) );
  OAI22X1 U3443 ( .A(n4748), .B(n4680), .C(n4746), .D(n4576), .Y(n5681) );
  XOR2X1 U3444 ( .A(n5682), .B(n4633), .Y(n3361) );
  OAI21X1 U3445 ( .A(n4555), .B(n4727), .C(n5683), .Y(n5682) );
  OAI22X1 U3446 ( .A(n4679), .B(n5684), .C(n4747), .D(n5684), .Y(n5683) );
  OAI22X1 U3447 ( .A(n4748), .B(n4576), .C(n4746), .D(n4676), .Y(n5684) );
  XOR2X1 U3448 ( .A(n5685), .B(n4633), .Y(n3360) );
  OAI21X1 U3449 ( .A(n4555), .B(n4726), .C(n5686), .Y(n5685) );
  OAI22X1 U3450 ( .A(n4577), .B(n5687), .C(n4747), .D(n5687), .Y(n5686) );
  OAI22X1 U3451 ( .A(n4748), .B(n4676), .C(n4746), .D(n4578), .Y(n5687) );
  XOR2X1 U3452 ( .A(n5688), .B(n4633), .Y(n3359) );
  OAI21X1 U3453 ( .A(n4555), .B(n4725), .C(n5689), .Y(n5688) );
  OAI22X1 U3454 ( .A(n4675), .B(n5690), .C(n4747), .D(n5690), .Y(n5689) );
  OAI22X1 U3455 ( .A(n4748), .B(n4578), .C(n4746), .D(n4671), .Y(n5690) );
  XOR2X1 U3456 ( .A(n5691), .B(n4633), .Y(n3358) );
  OAI21X1 U3457 ( .A(n4555), .B(n4724), .C(n5692), .Y(n5691) );
  OAI22X1 U3458 ( .A(n4579), .B(n5693), .C(n4747), .D(n5693), .Y(n5692) );
  OAI22X1 U3459 ( .A(n4748), .B(n4671), .C(n4746), .D(n4580), .Y(n5693) );
  XOR2X1 U3460 ( .A(n5694), .B(n4633), .Y(n3357) );
  OAI21X1 U3461 ( .A(n4555), .B(n4722), .C(n5695), .Y(n5694) );
  OAI22X1 U3462 ( .A(n4670), .B(n5696), .C(n4747), .D(n5696), .Y(n5695) );
  OAI22X1 U3463 ( .A(n4746), .B(n4666), .C(n4748), .D(n4580), .Y(n5696) );
  XOR2X1 U3464 ( .A(n5697), .B(n4633), .Y(n3356) );
  OAI21X1 U3465 ( .A(n4555), .B(n4721), .C(n5698), .Y(n5697) );
  OAI22X1 U3466 ( .A(n4581), .B(n5699), .C(n4747), .D(n5699), .Y(n5698) );
  OAI22X1 U3467 ( .A(n4748), .B(n4666), .C(n4746), .D(n4582), .Y(n5699) );
  XOR2X1 U3468 ( .A(n5700), .B(n4633), .Y(n3355) );
  OAI21X1 U3469 ( .A(n4555), .B(n4720), .C(n5701), .Y(n5700) );
  OAI22X1 U3470 ( .A(n4665), .B(n5702), .C(n4747), .D(n5702), .Y(n5701) );
  OAI22X1 U3471 ( .A(n4746), .B(n4662), .C(n4748), .D(n4582), .Y(n5702) );
  XOR2X1 U3472 ( .A(n5703), .B(n4633), .Y(n3354) );
  OAI21X1 U3473 ( .A(n4555), .B(n4719), .C(n5704), .Y(n5703) );
  OAI22X1 U3474 ( .A(n4583), .B(n5705), .C(n4747), .D(n5705), .Y(n5704) );
  OAI22X1 U3475 ( .A(n4748), .B(n4662), .C(n4746), .D(n4584), .Y(n5705) );
  XOR2X1 U3476 ( .A(n5706), .B(n4633), .Y(n3353) );
  OAI21X1 U3477 ( .A(n4555), .B(n4718), .C(n5707), .Y(n5706) );
  OAI22X1 U3478 ( .A(n4661), .B(n5708), .C(n4747), .D(n5708), .Y(n5707) );
  NAND3X1 U3479 ( .A(n5710), .B(n5711), .C(n5712), .Y(n5709) );
  OAI22X1 U3480 ( .A(n4748), .B(n4584), .C(n4657), .D(n4746), .Y(n5708) );
  NOR2X1 U3481 ( .A(n5711), .B(n5710), .Y(n5653) );
  NOR2X1 U3482 ( .A(n4749), .B(n5712), .Y(n5654) );
  XNOR2X1 U3483 ( .A(a[27]), .B(a[28]), .Y(n5712) );
  XOR2X1 U3484 ( .A(a[28]), .B(n4633), .Y(n5711) );
  XNOR2X1 U3485 ( .A(a[27]), .B(n4635), .Y(n5710) );
  OAI22X1 U3486 ( .A(n4743), .B(n4700), .C(n4557), .D(n4700), .Y(n3351) );
  OAI21X1 U3487 ( .A(n4557), .B(n4741), .C(n5713), .Y(n3350) );
  AOI22X1 U3488 ( .A(n4694), .B(n5714), .C(n4696), .D(n5715), .Y(n5713) );
  OAI21X1 U3489 ( .A(n4557), .B(n4738), .C(n5716), .Y(n3349) );
  OAI22X1 U3490 ( .A(n4698), .B(n5717), .C(n4742), .D(n5717), .Y(n5716) );
  OAI22X1 U3491 ( .A(n4744), .B(n4695), .C(n4743), .D(n4568), .Y(n5717) );
  OAI21X1 U3492 ( .A(n4557), .B(n4737), .C(n5718), .Y(n3348) );
  OAI22X1 U3493 ( .A(n4694), .B(n5719), .C(n4742), .D(n5719), .Y(n5718) );
  OAI22X1 U3494 ( .A(n4744), .B(n4568), .C(n4743), .D(n4693), .Y(n5719) );
  OAI21X1 U3495 ( .A(n4557), .B(n4736), .C(n5720), .Y(n3347) );
  OAI22X1 U3496 ( .A(n4569), .B(n5721), .C(n4742), .D(n5721), .Y(n5720) );
  OAI22X1 U3497 ( .A(n4744), .B(n4693), .C(n4743), .D(n4570), .Y(n5721) );
  OAI21X1 U3498 ( .A(n4557), .B(n4735), .C(n5722), .Y(n3346) );
  OAI22X1 U3499 ( .A(n4692), .B(n5723), .C(n4742), .D(n5723), .Y(n5722) );
  OAI22X1 U3500 ( .A(n4744), .B(n4570), .C(n4743), .D(n4689), .Y(n5723) );
  OAI21X1 U3501 ( .A(n4557), .B(n4734), .C(n5724), .Y(n3345) );
  OAI22X1 U3502 ( .A(n4571), .B(n5725), .C(n4742), .D(n5725), .Y(n5724) );
  OAI22X1 U3503 ( .A(n4744), .B(n4689), .C(n4743), .D(n4572), .Y(n5725) );
  OAI21X1 U3504 ( .A(n4557), .B(n4733), .C(n5726), .Y(n3344) );
  OAI22X1 U3505 ( .A(n4688), .B(n5727), .C(n4742), .D(n5727), .Y(n5726) );
  OAI22X1 U3506 ( .A(n4744), .B(n4572), .C(n4743), .D(n4685), .Y(n5727) );
  OAI21X1 U3507 ( .A(n4557), .B(n4731), .C(n5728), .Y(n3343) );
  OAI22X1 U3508 ( .A(n4573), .B(n5729), .C(n4742), .D(n5729), .Y(n5728) );
  OAI22X1 U3509 ( .A(n4744), .B(n4685), .C(n4743), .D(n4574), .Y(n5729) );
  OAI21X1 U3510 ( .A(n4557), .B(n4730), .C(n5730), .Y(n3342) );
  OAI22X1 U3511 ( .A(n4684), .B(n5731), .C(n4742), .D(n5731), .Y(n5730) );
  OAI22X1 U3512 ( .A(n4744), .B(n4574), .C(n4743), .D(n4680), .Y(n5731) );
  OAI21X1 U3513 ( .A(n4557), .B(n4729), .C(n5732), .Y(n3341) );
  OAI22X1 U3514 ( .A(n4575), .B(n5733), .C(n4742), .D(n5733), .Y(n5732) );
  OAI22X1 U3515 ( .A(n4744), .B(n4680), .C(n4743), .D(n4576), .Y(n5733) );
  OAI21X1 U3516 ( .A(n4557), .B(n4727), .C(n5734), .Y(n3340) );
  OAI22X1 U3517 ( .A(n4679), .B(n5735), .C(n4742), .D(n5735), .Y(n5734) );
  OAI22X1 U3518 ( .A(n4744), .B(n4576), .C(n4743), .D(n4676), .Y(n5735) );
  OAI21X1 U3519 ( .A(n4557), .B(n4726), .C(n5736), .Y(n3339) );
  OAI22X1 U3520 ( .A(n4577), .B(n5737), .C(n4742), .D(n5737), .Y(n5736) );
  OAI22X1 U3521 ( .A(n4744), .B(n4676), .C(n4743), .D(n4578), .Y(n5737) );
  OAI21X1 U3522 ( .A(n4557), .B(n4725), .C(n5738), .Y(n3338) );
  OAI22X1 U3523 ( .A(n4675), .B(n5739), .C(n4742), .D(n5739), .Y(n5738) );
  OAI22X1 U3524 ( .A(n4744), .B(n4578), .C(n4743), .D(n4671), .Y(n5739) );
  OAI21X1 U3525 ( .A(n4557), .B(n4722), .C(n5740), .Y(n3337) );
  OAI22X1 U3526 ( .A(n4670), .B(n5741), .C(n4742), .D(n5741), .Y(n5740) );
  OAI22X1 U3527 ( .A(n4743), .B(n4666), .C(n4744), .D(n4580), .Y(n5741) );
  OAI21X1 U3528 ( .A(n4557), .B(n4721), .C(n5742), .Y(n3336) );
  OAI22X1 U3529 ( .A(n4581), .B(n5743), .C(n4742), .D(n5743), .Y(n5742) );
  OAI22X1 U3530 ( .A(n4744), .B(n4666), .C(n4582), .D(n4743), .Y(n5743) );
  OAI21X1 U3531 ( .A(n4557), .B(n4724), .C(n5744), .Y(n2429) );
  OAI22X1 U3532 ( .A(n4579), .B(n5745), .C(n4742), .D(n5745), .Y(n5744) );
  NAND3X1 U3533 ( .A(n5747), .B(a[31]), .C(n5748), .Y(n5746) );
  OAI22X1 U3534 ( .A(n4744), .B(n4671), .C(n4743), .D(n4580), .Y(n5745) );
  NOR2X1 U3535 ( .A(n5747), .B(a[31]), .Y(n5714) );
  NOR2X1 U3536 ( .A(n4745), .B(n5748), .Y(n5715) );
  XNOR2X1 U3537 ( .A(a[30]), .B(a[31]), .Y(n5748) );
  XNOR2X1 U3538 ( .A(a[30]), .B(n4633), .Y(n5747) );
endmodule


module poly5_DW01_sub_22 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31, n32,
         n33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n46, n47, n48,
         n49, n50, n51, n53, n54, n55, n56, n57, n58, n59, n62, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79, n80, n82,
         n83, n84, n85, n86, n88, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n102, n103, n104, n105, n106, n107, n108, n109, \B[0] , n212,
         n213, n214, n215, n216, n217, n218, n219, n220;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2X1 U4 ( .A(n5), .B(B[31]), .Y(DIFF[31]) );
  XNOR2X1 U5 ( .A(n10), .B(B[30]), .Y(DIFF[30]) );
  NOR2X1 U6 ( .A(n220), .B(n6), .Y(n5) );
  NAND2X1 U7 ( .A(n7), .B(n215), .Y(n6) );
  NOR2X1 U8 ( .A(n8), .B(n4), .Y(n7) );
  NAND2X1 U9 ( .A(n9), .B(n14), .Y(n8) );
  XNOR2X1 U11 ( .A(n15), .B(B[29]), .Y(DIFF[29]) );
  NOR2X1 U12 ( .A(n220), .B(n11), .Y(n10) );
  NAND2X1 U13 ( .A(n12), .B(n3), .Y(n11) );
  NOR2X1 U14 ( .A(n13), .B(n4), .Y(n12) );
  NOR2X1 U16 ( .A(B[29]), .B(B[28]), .Y(n14) );
  XNOR2X1 U17 ( .A(n18), .B(B[28]), .Y(DIFF[28]) );
  NOR2X1 U18 ( .A(n220), .B(n16), .Y(n15) );
  NAND2X1 U19 ( .A(n17), .B(n215), .Y(n16) );
  NOR2X1 U20 ( .A(B[28]), .B(n4), .Y(n17) );
  XNOR2X1 U21 ( .A(n22), .B(B[27]), .Y(DIFF[27]) );
  NOR2X1 U22 ( .A(n220), .B(n19), .Y(n18) );
  NAND2X1 U23 ( .A(n20), .B(n3), .Y(n19) );
  NAND2X1 U25 ( .A(n21), .B(n27), .Y(n4) );
  NOR2X1 U26 ( .A(B[27]), .B(B[26]), .Y(n21) );
  XNOR2X1 U27 ( .A(n25), .B(B[26]), .Y(DIFF[26]) );
  NOR2X1 U28 ( .A(n220), .B(n23), .Y(n22) );
  NAND2X1 U29 ( .A(n24), .B(n215), .Y(n23) );
  NOR2X1 U30 ( .A(B[26]), .B(n28), .Y(n24) );
  XNOR2X1 U31 ( .A(n30), .B(B[25]), .Y(DIFF[25]) );
  NOR2X1 U32 ( .A(n220), .B(n26), .Y(n25) );
  NAND2X1 U33 ( .A(n27), .B(n215), .Y(n26) );
  NOR2X1 U36 ( .A(B[25]), .B(B[24]), .Y(n27) );
  XNOR2X1 U37 ( .A(n33), .B(B[24]), .Y(DIFF[24]) );
  NOR2X1 U38 ( .A(n220), .B(n31), .Y(n30) );
  NAND2X1 U39 ( .A(n32), .B(n215), .Y(n31) );
  XNOR2X1 U41 ( .A(n38), .B(B[23]), .Y(DIFF[23]) );
  NOR2X1 U42 ( .A(n34), .B(n220), .Y(n33) );
  NOR2X1 U44 ( .A(n36), .B(n50), .Y(n3) );
  NAND2X1 U45 ( .A(n37), .B(n43), .Y(n36) );
  NOR2X1 U46 ( .A(B[23]), .B(B[22]), .Y(n37) );
  XNOR2X1 U47 ( .A(n41), .B(B[22]), .Y(DIFF[22]) );
  NOR2X1 U48 ( .A(n39), .B(n220), .Y(n38) );
  NAND2X1 U49 ( .A(n51), .B(n40), .Y(n39) );
  NOR2X1 U50 ( .A(B[22]), .B(n44), .Y(n40) );
  XNOR2X1 U51 ( .A(n46), .B(B[21]), .Y(DIFF[21]) );
  NOR2X1 U52 ( .A(n42), .B(n220), .Y(n41) );
  NAND2X1 U53 ( .A(n43), .B(n51), .Y(n42) );
  NOR2X1 U56 ( .A(B[21]), .B(B[20]), .Y(n43) );
  NOR2X1 U58 ( .A(n47), .B(n220), .Y(n46) );
  NAND2X1 U59 ( .A(n48), .B(n51), .Y(n47) );
  XNOR2X1 U61 ( .A(n54), .B(B[19]), .Y(DIFF[19]) );
  NOR2X1 U62 ( .A(n50), .B(n220), .Y(n49) );
  NAND2X1 U65 ( .A(n53), .B(n59), .Y(n50) );
  NOR2X1 U66 ( .A(B[19]), .B(B[18]), .Y(n53) );
  XNOR2X1 U67 ( .A(n57), .B(B[18]), .Y(DIFF[18]) );
  NOR2X1 U68 ( .A(n55), .B(n220), .Y(n54) );
  NAND2X1 U69 ( .A(n56), .B(n59), .Y(n55) );
  XNOR2X1 U71 ( .A(n62), .B(B[17]), .Y(DIFF[17]) );
  NOR2X1 U72 ( .A(n58), .B(n220), .Y(n57) );
  NOR2X1 U76 ( .A(B[17]), .B(B[16]), .Y(n59) );
  XOR2X1 U77 ( .A(n220), .B(B[16]), .Y(DIFF[16]) );
  NOR2X1 U78 ( .A(B[16]), .B(n220), .Y(n62) );
  XNOR2X1 U79 ( .A(n67), .B(B[15]), .Y(DIFF[15]) );
  NOR2X1 U81 ( .A(n65), .B(n79), .Y(n64) );
  NAND2X1 U82 ( .A(n66), .B(n72), .Y(n65) );
  NOR2X1 U83 ( .A(B[15]), .B(B[14]), .Y(n66) );
  XNOR2X1 U84 ( .A(n70), .B(B[14]), .Y(DIFF[14]) );
  NOR2X1 U85 ( .A(n218), .B(n68), .Y(n67) );
  NAND2X1 U86 ( .A(n80), .B(n69), .Y(n68) );
  NOR2X1 U87 ( .A(B[14]), .B(n73), .Y(n69) );
  XNOR2X1 U88 ( .A(n75), .B(B[13]), .Y(DIFF[13]) );
  NOR2X1 U89 ( .A(n218), .B(n71), .Y(n70) );
  NAND2X1 U90 ( .A(n212), .B(n80), .Y(n71) );
  NOR2X1 U93 ( .A(B[13]), .B(B[12]), .Y(n72) );
  XNOR2X1 U94 ( .A(n78), .B(B[12]), .Y(DIFF[12]) );
  NOR2X1 U95 ( .A(n217), .B(n76), .Y(n75) );
  NAND2X1 U96 ( .A(n77), .B(n80), .Y(n76) );
  XNOR2X1 U98 ( .A(n83), .B(B[11]), .Y(DIFF[11]) );
  NOR2X1 U99 ( .A(n216), .B(n217), .Y(n78) );
  NAND2X1 U102 ( .A(n82), .B(n88), .Y(n79) );
  NOR2X1 U103 ( .A(B[11]), .B(B[10]), .Y(n82) );
  XNOR2X1 U104 ( .A(n86), .B(B[10]), .Y(DIFF[10]) );
  NOR2X1 U105 ( .A(n84), .B(n218), .Y(n83) );
  NAND2X1 U106 ( .A(n85), .B(n214), .Y(n84) );
  NOR2X1 U109 ( .A(n213), .B(n218), .Y(n86) );
  NOR2X1 U113 ( .A(B[9]), .B(B[8]), .Y(n88) );
  XOR2X1 U114 ( .A(n218), .B(B[8]), .Y(DIFF[8]) );
  NOR2X1 U115 ( .A(B[8]), .B(n217), .Y(n91) );
  XOR2X1 U116 ( .A(n96), .B(B[7]), .Y(DIFF[7]) );
  NOR2X1 U118 ( .A(n94), .B(n105), .Y(n93) );
  NAND2X1 U119 ( .A(n95), .B(n99), .Y(n94) );
  NOR2X1 U120 ( .A(B[7]), .B(B[6]), .Y(n95) );
  XOR2X1 U121 ( .A(n98), .B(B[6]), .Y(DIFF[6]) );
  NAND2X1 U122 ( .A(n104), .B(n97), .Y(n96) );
  NOR2X1 U123 ( .A(B[6]), .B(n100), .Y(n97) );
  XOR2X1 U124 ( .A(n102), .B(B[5]), .Y(DIFF[5]) );
  NAND2X1 U125 ( .A(n99), .B(n104), .Y(n98) );
  NOR2X1 U128 ( .A(B[5]), .B(B[4]), .Y(n99) );
  XNOR2X1 U129 ( .A(n104), .B(B[4]), .Y(DIFF[4]) );
  NAND2X1 U130 ( .A(n103), .B(n104), .Y(n102) );
  XNOR2X1 U132 ( .A(n107), .B(B[3]), .Y(DIFF[3]) );
  NAND2X1 U134 ( .A(n109), .B(n106), .Y(n105) );
  NOR2X1 U135 ( .A(B[3]), .B(B[2]), .Y(n106) );
  XOR2X1 U136 ( .A(n108), .B(B[2]), .Y(DIFF[2]) );
  NOR2X1 U137 ( .A(B[2]), .B(n108), .Y(n107) );
  XOR2X1 U138 ( .A(B[1]), .B(\B[0] ), .Y(DIFF[1]) );
  NOR2X1 U140 ( .A(\B[0] ), .B(B[1]), .Y(n109) );
  BUFX4 U144 ( .A(n92), .Y(n218) );
  XOR2X1 U145 ( .A(n49), .B(n48), .Y(DIFF[20]) );
  INVX1 U146 ( .A(n73), .Y(n212) );
  INVX1 U147 ( .A(n88), .Y(n213) );
  INVX1 U148 ( .A(n213), .Y(n214) );
  NOR2X1 U149 ( .A(n36), .B(n50), .Y(n215) );
  INVX1 U150 ( .A(n80), .Y(n216) );
  XNOR2X1 U151 ( .A(n91), .B(B[9]), .Y(DIFF[9]) );
  BUFX2 U152 ( .A(n92), .Y(n217) );
  INVX1 U153 ( .A(n79), .Y(n80) );
  INVX1 U154 ( .A(n99), .Y(n100) );
  INVX1 U155 ( .A(B[10]), .Y(n85) );
  INVX1 U156 ( .A(B[12]), .Y(n77) );
  INVX1 U157 ( .A(n72), .Y(n73) );
  INVX1 U158 ( .A(n93), .Y(n92) );
  INVX1 U159 ( .A(n59), .Y(n58) );
  INVX1 U160 ( .A(n50), .Y(n51) );
  AND2X2 U161 ( .A(n93), .B(n64), .Y(n219) );
  INVX1 U162 ( .A(n3), .Y(n34) );
  INVX1 U163 ( .A(n109), .Y(n108) );
  INVX1 U164 ( .A(n105), .Y(n104) );
  INVX8 U165 ( .A(n219), .Y(n220) );
  INVX2 U166 ( .A(B[30]), .Y(n9) );
  INVX2 U167 ( .A(B[18]), .Y(n56) );
  INVX2 U168 ( .A(B[20]), .Y(n48) );
  INVX2 U169 ( .A(n43), .Y(n44) );
  INVX2 U170 ( .A(B[24]), .Y(n32) );
  INVX2 U171 ( .A(n27), .Y(n28) );
  INVX2 U172 ( .A(n4), .Y(n20) );
  INVX2 U173 ( .A(n14), .Y(n13) );
  INVX2 U174 ( .A(B[4]), .Y(n103) );
endmodule


module poly5_DW01_sub_39 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n45,
         n46, n47, n48, n49, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n70, n71, n72, n73, n74, n75,
         n76, n77, n79, n80, n81, n82, n83, n84, n86, n87, n90, n91, n92, n93,
         n94, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n108, n110, n111, n112, n113, n114, n115, n116, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n273, n274, n275, n276, n277,
         n278;

  XOR2X1 U3 ( .A(n3), .B(B[47]), .Y(DIFF[47]) );
  XOR2X1 U4 ( .A(n9), .B(B[46]), .Y(DIFF[46]) );
  NAND2X1 U5 ( .A(n2), .B(n4), .Y(n3) );
  NAND2X1 U7 ( .A(n32), .B(n6), .Y(n5) );
  NOR2X1 U8 ( .A(n7), .B(n19), .Y(n6) );
  NAND2X1 U9 ( .A(n8), .B(n12), .Y(n7) );
  XOR2X1 U11 ( .A(n13), .B(B[45]), .Y(DIFF[45]) );
  NAND2X1 U12 ( .A(n2), .B(n10), .Y(n9) );
  NOR2X1 U13 ( .A(n11), .B(n17), .Y(n10) );
  NOR2X1 U15 ( .A(B[45]), .B(B[44]), .Y(n12) );
  XOR2X1 U16 ( .A(n15), .B(B[44]), .Y(DIFF[44]) );
  NAND2X1 U17 ( .A(n2), .B(n14), .Y(n13) );
  NOR2X1 U18 ( .A(B[44]), .B(n17), .Y(n14) );
  XOR2X1 U19 ( .A(n21), .B(B[43]), .Y(DIFF[43]) );
  NAND2X1 U20 ( .A(n16), .B(n2), .Y(n15) );
  NAND2X1 U22 ( .A(n18), .B(n32), .Y(n17) );
  NAND2X1 U24 ( .A(n20), .B(n26), .Y(n19) );
  NOR2X1 U25 ( .A(B[43]), .B(B[42]), .Y(n20) );
  XOR2X1 U26 ( .A(n23), .B(B[42]), .Y(DIFF[42]) );
  NAND2X1 U27 ( .A(n2), .B(n22), .Y(n21) );
  NOR2X1 U28 ( .A(B[42]), .B(n25), .Y(n22) );
  XOR2X1 U29 ( .A(n27), .B(B[41]), .Y(DIFF[41]) );
  NAND2X1 U30 ( .A(n24), .B(n2), .Y(n23) );
  NAND2X1 U32 ( .A(n26), .B(n32), .Y(n25) );
  NOR2X1 U33 ( .A(B[41]), .B(B[40]), .Y(n26) );
  XOR2X1 U34 ( .A(n29), .B(B[40]), .Y(DIFF[40]) );
  NAND2X1 U35 ( .A(n28), .B(n2), .Y(n27) );
  NOR2X1 U36 ( .A(B[40]), .B(n31), .Y(n28) );
  XOR2X1 U37 ( .A(n35), .B(B[39]), .Y(DIFF[39]) );
  NAND2X1 U38 ( .A(n30), .B(n2), .Y(n29) );
  NOR2X1 U41 ( .A(n33), .B(n47), .Y(n32) );
  NAND2X1 U42 ( .A(n34), .B(n40), .Y(n33) );
  NOR2X1 U43 ( .A(B[39]), .B(B[38]), .Y(n34) );
  XOR2X1 U44 ( .A(n37), .B(B[38]), .Y(DIFF[38]) );
  NAND2X1 U45 ( .A(n36), .B(n1), .Y(n35) );
  NOR2X1 U46 ( .A(B[38]), .B(n39), .Y(n36) );
  XOR2X1 U47 ( .A(n41), .B(B[37]), .Y(DIFF[37]) );
  NAND2X1 U48 ( .A(n38), .B(n1), .Y(n37) );
  NAND2X1 U50 ( .A(n40), .B(n46), .Y(n39) );
  NOR2X1 U51 ( .A(B[37]), .B(B[36]), .Y(n40) );
  XOR2X1 U52 ( .A(n43), .B(B[36]), .Y(DIFF[36]) );
  NAND2X1 U53 ( .A(n42), .B(n1), .Y(n41) );
  NOR2X1 U54 ( .A(B[36]), .B(n45), .Y(n42) );
  XOR2X1 U55 ( .A(n49), .B(B[35]), .Y(DIFF[35]) );
  NAND2X1 U56 ( .A(n46), .B(n1), .Y(n43) );
  NAND2X1 U60 ( .A(n48), .B(n54), .Y(n47) );
  NOR2X1 U61 ( .A(B[35]), .B(B[34]), .Y(n48) );
  XOR2X1 U62 ( .A(n51), .B(B[34]), .Y(DIFF[34]) );
  NAND2X1 U63 ( .A(n50), .B(n1), .Y(n49) );
  NOR2X1 U64 ( .A(B[34]), .B(n53), .Y(n50) );
  XOR2X1 U65 ( .A(n55), .B(B[33]), .Y(DIFF[33]) );
  NAND2X1 U66 ( .A(n54), .B(n1), .Y(n51) );
  NOR2X1 U69 ( .A(B[33]), .B(B[32]), .Y(n54) );
  XNOR2X1 U70 ( .A(n1), .B(B[32]), .Y(DIFF[32]) );
  NAND2X1 U71 ( .A(n56), .B(n1), .Y(n55) );
  XOR2X1 U73 ( .A(n62), .B(B[31]), .Y(DIFF[31]) );
  NOR2X1 U74 ( .A(n123), .B(n58), .Y(n57) );
  NAND2X1 U75 ( .A(n59), .B(n97), .Y(n58) );
  NOR2X1 U76 ( .A(n60), .B(n80), .Y(n59) );
  NAND2X1 U77 ( .A(n61), .B(n71), .Y(n60) );
  NOR2X1 U78 ( .A(B[31]), .B(B[30]), .Y(n61) );
  XOR2X1 U79 ( .A(n66), .B(B[30]), .Y(DIFF[30]) );
  NAND2X1 U80 ( .A(n122), .B(n63), .Y(n62) );
  NOR2X1 U81 ( .A(n64), .B(n96), .Y(n63) );
  NAND2X1 U82 ( .A(n79), .B(n65), .Y(n64) );
  NOR2X1 U83 ( .A(B[30]), .B(n70), .Y(n65) );
  XOR2X1 U84 ( .A(n72), .B(n273), .Y(DIFF[29]) );
  NAND2X1 U85 ( .A(n122), .B(n67), .Y(n66) );
  NOR2X1 U86 ( .A(n68), .B(n96), .Y(n67) );
  NAND2X1 U87 ( .A(n71), .B(n79), .Y(n68) );
  NOR2X1 U90 ( .A(B[29]), .B(B[28]), .Y(n71) );
  XOR2X1 U91 ( .A(n76), .B(B[28]), .Y(DIFF[28]) );
  NAND2X1 U92 ( .A(n122), .B(n73), .Y(n72) );
  NOR2X1 U93 ( .A(n74), .B(n96), .Y(n73) );
  NAND2X1 U94 ( .A(n75), .B(n79), .Y(n74) );
  XOR2X1 U96 ( .A(n82), .B(B[27]), .Y(DIFF[27]) );
  NAND2X1 U97 ( .A(n122), .B(n77), .Y(n76) );
  NOR2X1 U98 ( .A(n80), .B(n96), .Y(n77) );
  NAND2X1 U101 ( .A(n81), .B(n91), .Y(n80) );
  NOR2X1 U102 ( .A(B[27]), .B(B[26]), .Y(n81) );
  XOR2X1 U103 ( .A(n86), .B(B[26]), .Y(DIFF[26]) );
  NAND2X1 U104 ( .A(n122), .B(n83), .Y(n82) );
  NOR2X1 U105 ( .A(n96), .B(n84), .Y(n83) );
  XOR2X1 U108 ( .A(n92), .B(B[25]), .Y(DIFF[25]) );
  NAND2X1 U109 ( .A(n122), .B(n87), .Y(n86) );
  NOR2X1 U110 ( .A(n90), .B(n96), .Y(n87) );
  NOR2X1 U114 ( .A(B[25]), .B(B[24]), .Y(n91) );
  XOR2X1 U115 ( .A(n94), .B(B[24]), .Y(DIFF[24]) );
  NAND2X1 U116 ( .A(n122), .B(n93), .Y(n92) );
  NOR2X1 U117 ( .A(B[24]), .B(n96), .Y(n93) );
  XOR2X1 U118 ( .A(n100), .B(B[23]), .Y(DIFF[23]) );
  NAND2X1 U119 ( .A(n97), .B(n122), .Y(n94) );
  NOR2X1 U122 ( .A(n98), .B(n112), .Y(n97) );
  NAND2X1 U123 ( .A(n99), .B(n105), .Y(n98) );
  NOR2X1 U124 ( .A(B[23]), .B(B[22]), .Y(n99) );
  XOR2X1 U125 ( .A(n102), .B(B[22]), .Y(DIFF[22]) );
  NAND2X1 U126 ( .A(n122), .B(n101), .Y(n100) );
  NOR2X1 U127 ( .A(B[22]), .B(n104), .Y(n101) );
  NAND2X1 U129 ( .A(n103), .B(n122), .Y(n102) );
  NAND2X1 U131 ( .A(n105), .B(n111), .Y(n104) );
  NOR2X1 U132 ( .A(B[21]), .B(B[20]), .Y(n105) );
  XOR2X1 U133 ( .A(n108), .B(B[20]), .Y(DIFF[20]) );
  XOR2X1 U136 ( .A(n114), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U141 ( .A(n119), .B(n113), .Y(n112) );
  NOR2X1 U142 ( .A(B[19]), .B(B[18]), .Y(n113) );
  XOR2X1 U143 ( .A(n116), .B(B[18]), .Y(DIFF[18]) );
  NAND2X1 U144 ( .A(n115), .B(n122), .Y(n114) );
  NOR2X1 U145 ( .A(B[18]), .B(n118), .Y(n115) );
  XOR2X1 U146 ( .A(n120), .B(B[17]), .Y(DIFF[17]) );
  NAND2X1 U147 ( .A(n119), .B(n122), .Y(n116) );
  NOR2X1 U150 ( .A(B[17]), .B(B[16]), .Y(n119) );
  XNOR2X1 U151 ( .A(n122), .B(B[16]), .Y(DIFF[16]) );
  NAND2X1 U152 ( .A(n121), .B(n122), .Y(n120) );
  INVX4 U154 ( .A(n123), .Y(n122) );
  NAND2X1 U155 ( .A(n131), .B(n124), .Y(n123) );
  NOR2X1 U156 ( .A(n125), .B(n128), .Y(n124) );
  NAND2X1 U157 ( .A(n126), .B(n127), .Y(n125) );
  NOR2X1 U158 ( .A(B[15]), .B(B[14]), .Y(n126) );
  NOR2X1 U159 ( .A(B[13]), .B(B[12]), .Y(n127) );
  NAND2X1 U160 ( .A(n129), .B(n130), .Y(n128) );
  NOR2X1 U161 ( .A(B[11]), .B(B[10]), .Y(n129) );
  NOR2X1 U162 ( .A(B[9]), .B(B[8]), .Y(n130) );
  NOR2X1 U163 ( .A(n135), .B(n132), .Y(n131) );
  NAND2X1 U164 ( .A(n133), .B(n134), .Y(n132) );
  NOR2X1 U165 ( .A(B[7]), .B(B[6]), .Y(n133) );
  NOR2X1 U166 ( .A(B[5]), .B(B[4]), .Y(n134) );
  NAND2X1 U167 ( .A(n137), .B(n136), .Y(n135) );
  NOR2X1 U168 ( .A(B[3]), .B(B[2]), .Y(n136) );
  NOR2X1 U169 ( .A(B[0]), .B(B[1]), .Y(n137) );
  BUFX4 U173 ( .A(n57), .Y(n1) );
  INVX4 U174 ( .A(n97), .Y(n96) );
  OR2X2 U175 ( .A(n110), .B(n123), .Y(n108) );
  INVX1 U176 ( .A(n111), .Y(n110) );
  INVX1 U177 ( .A(n47), .Y(n46) );
  BUFX2 U178 ( .A(B[29]), .Y(n273) );
  INVX1 U179 ( .A(n39), .Y(n38) );
  INVX1 U180 ( .A(n25), .Y(n24) );
  INVX2 U181 ( .A(n46), .Y(n45) );
  INVX1 U182 ( .A(n31), .Y(n30) );
  INVX1 U183 ( .A(n19), .Y(n18) );
  INVX2 U184 ( .A(n80), .Y(n79) );
  INVX1 U185 ( .A(B[32]), .Y(n56) );
  INVX1 U186 ( .A(n104), .Y(n103) );
  INVX1 U187 ( .A(n119), .Y(n118) );
  INVX1 U188 ( .A(B[46]), .Y(n8) );
  INVX1 U189 ( .A(B[28]), .Y(n75) );
  INVX2 U190 ( .A(B[16]), .Y(n121) );
  BUFX2 U191 ( .A(n57), .Y(n2) );
  INVX2 U192 ( .A(n54), .Y(n53) );
  INVX1 U193 ( .A(n5), .Y(n4) );
  OR2X2 U194 ( .A(B[26]), .B(n90), .Y(n84) );
  NAND2X1 U195 ( .A(n106), .B(n275), .Y(n276) );
  NAND2X1 U196 ( .A(n274), .B(B[21]), .Y(n277) );
  NAND2X1 U197 ( .A(n276), .B(n277), .Y(DIFF[21]) );
  INVX1 U198 ( .A(n106), .Y(n274) );
  INVX1 U199 ( .A(B[21]), .Y(n275) );
  OR2X2 U200 ( .A(B[20]), .B(n278), .Y(n106) );
  NAND2X1 U201 ( .A(n111), .B(n122), .Y(n278) );
  INVX1 U202 ( .A(n17), .Y(n16) );
  INVX2 U203 ( .A(n91), .Y(n90) );
  INVX2 U204 ( .A(n112), .Y(n111) );
  INVX2 U205 ( .A(n32), .Y(n31) );
  INVX2 U206 ( .A(n71), .Y(n70) );
  INVX1 U207 ( .A(n12), .Y(n11) );
endmodule


module poly5_DW01_sub_43 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n57, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, \B[0] ;
  assign n57 = B[10];
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2X1 U1 ( .A(n1), .B(B[31]), .Y(DIFF[31]) );
  XOR2X1 U2 ( .A(n2), .B(B[30]), .Y(DIFF[30]) );
  NOR2X1 U3 ( .A(B[30]), .B(n2), .Y(n1) );
  XNOR2X1 U4 ( .A(n6), .B(B[29]), .Y(DIFF[29]) );
  NAND2X1 U5 ( .A(n24), .B(n3), .Y(n2) );
  NOR2X1 U6 ( .A(n10), .B(n4), .Y(n3) );
  NAND2X1 U7 ( .A(n8), .B(n5), .Y(n4) );
  XNOR2X1 U9 ( .A(n9), .B(B[28]), .Y(DIFF[28]) );
  NOR2X1 U10 ( .A(n23), .B(n7), .Y(n6) );
  NAND2X1 U11 ( .A(n8), .B(n11), .Y(n7) );
  XNOR2X1 U13 ( .A(n14), .B(B[27]), .Y(DIFF[27]) );
  NOR2X1 U14 ( .A(n10), .B(n23), .Y(n9) );
  NAND2X1 U17 ( .A(n19), .B(n13), .Y(n10) );
  NOR2X1 U18 ( .A(B[26]), .B(B[27]), .Y(n13) );
  XNOR2X1 U19 ( .A(n17), .B(B[26]), .Y(DIFF[26]) );
  NOR2X1 U20 ( .A(n15), .B(n23), .Y(n14) );
  NAND2X1 U21 ( .A(n16), .B(n19), .Y(n15) );
  XNOR2X1 U23 ( .A(n22), .B(B[25]), .Y(DIFF[25]) );
  NOR2X1 U24 ( .A(n18), .B(n23), .Y(n17) );
  NOR2X1 U28 ( .A(B[25]), .B(B[24]), .Y(n19) );
  XOR2X1 U29 ( .A(n23), .B(B[24]), .Y(DIFF[24]) );
  NOR2X1 U30 ( .A(B[24]), .B(n23), .Y(n22) );
  XOR2X1 U31 ( .A(n27), .B(B[23]), .Y(DIFF[23]) );
  NOR2X1 U33 ( .A(n36), .B(n25), .Y(n24) );
  NAND2X1 U34 ( .A(n26), .B(n30), .Y(n25) );
  NOR2X1 U35 ( .A(B[23]), .B(B[22]), .Y(n26) );
  XOR2X1 U36 ( .A(n29), .B(B[22]), .Y(DIFF[22]) );
  NAND2X1 U37 ( .A(n35), .B(n28), .Y(n27) );
  NOR2X1 U38 ( .A(B[22]), .B(n31), .Y(n28) );
  XOR2X1 U39 ( .A(n33), .B(B[21]), .Y(DIFF[21]) );
  NAND2X1 U40 ( .A(n30), .B(n35), .Y(n29) );
  NOR2X1 U43 ( .A(B[21]), .B(B[20]), .Y(n30) );
  XNOR2X1 U44 ( .A(n35), .B(B[20]), .Y(DIFF[20]) );
  NAND2X1 U45 ( .A(n34), .B(n35), .Y(n33) );
  XNOR2X1 U47 ( .A(n38), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U49 ( .A(n40), .B(n37), .Y(n36) );
  NOR2X1 U50 ( .A(B[19]), .B(B[18]), .Y(n37) );
  XOR2X1 U51 ( .A(n39), .B(B[18]), .Y(DIFF[18]) );
  NOR2X1 U52 ( .A(B[18]), .B(n39), .Y(n38) );
  XOR2X1 U53 ( .A(B[17]), .B(n41), .Y(DIFF[17]) );
  NOR2X1 U55 ( .A(B[17]), .B(n41), .Y(n40) );
  XNOR2X1 U56 ( .A(B[16]), .B(n43), .Y(DIFF[16]) );
  NAND2X1 U57 ( .A(n43), .B(n42), .Y(n41) );
  XOR2X1 U59 ( .A(n46), .B(B[15]), .Y(DIFF[15]) );
  NOR2X1 U60 ( .A(n51), .B(n44), .Y(n43) );
  NAND2X1 U61 ( .A(n45), .B(n47), .Y(n44) );
  XOR2X1 U63 ( .A(n48), .B(B[14]), .Y(DIFF[14]) );
  NAND2X1 U64 ( .A(n47), .B(n50), .Y(n46) );
  NOR2X1 U65 ( .A(B[13]), .B(B[14]), .Y(n47) );
  XNOR2X1 U66 ( .A(n50), .B(B[13]), .Y(DIFF[13]) );
  NAND2X1 U67 ( .A(n49), .B(n50), .Y(n48) );
  XNOR2X1 U69 ( .A(n53), .B(B[12]), .Y(DIFF[12]) );
  NAND2X1 U71 ( .A(n60), .B(n52), .Y(n51) );
  NOR2X1 U72 ( .A(B[12]), .B(n54), .Y(n52) );
  XNOR2X1 U73 ( .A(n56), .B(B[11]), .Y(DIFF[11]) );
  NOR2X1 U74 ( .A(n54), .B(n59), .Y(n53) );
  XOR2X1 U77 ( .A(n59), .B(n57), .Y(DIFF[10]) );
  NOR2X1 U78 ( .A(n57), .B(n59), .Y(n56) );
  XOR2X1 U81 ( .A(B[9]), .B(n63), .Y(DIFF[9]) );
  NOR2X1 U83 ( .A(n66), .B(n61), .Y(n60) );
  NAND2X1 U84 ( .A(n64), .B(n62), .Y(n61) );
  XNOR2X1 U86 ( .A(B[8]), .B(n65), .Y(DIFF[8]) );
  NAND2X1 U87 ( .A(n64), .B(n65), .Y(n63) );
  XNOR2X1 U89 ( .A(n68), .B(B[7]), .Y(DIFF[7]) );
  NAND2X1 U91 ( .A(n67), .B(n70), .Y(n66) );
  NOR2X1 U92 ( .A(B[6]), .B(B[7]), .Y(n67) );
  XOR2X1 U93 ( .A(n69), .B(B[6]), .Y(DIFF[6]) );
  NOR2X1 U94 ( .A(B[6]), .B(n69), .Y(n68) );
  XOR2X1 U95 ( .A(n73), .B(B[5]), .Y(DIFF[5]) );
  NOR2X1 U97 ( .A(n76), .B(n71), .Y(n70) );
  NAND2X1 U98 ( .A(n74), .B(n72), .Y(n71) );
  XNOR2X1 U100 ( .A(n75), .B(B[4]), .Y(DIFF[4]) );
  NAND2X1 U101 ( .A(n74), .B(n75), .Y(n73) );
  XNOR2X1 U103 ( .A(n78), .B(B[3]), .Y(DIFF[3]) );
  NAND2X1 U105 ( .A(n80), .B(n77), .Y(n76) );
  NOR2X1 U106 ( .A(B[3]), .B(B[2]), .Y(n77) );
  XOR2X1 U107 ( .A(n79), .B(B[2]), .Y(DIFF[2]) );
  NOR2X1 U108 ( .A(B[2]), .B(n79), .Y(n78) );
  XOR2X1 U109 ( .A(B[1]), .B(\B[0] ), .Y(DIFF[1]) );
  NOR2X1 U111 ( .A(\B[0] ), .B(B[1]), .Y(n80) );
  INVX2 U115 ( .A(B[4]), .Y(n74) );
  INVX2 U116 ( .A(B[8]), .Y(n64) );
  INVX2 U117 ( .A(B[28]), .Y(n8) );
  OR2X2 U118 ( .A(B[11]), .B(n57), .Y(n54) );
  INVX1 U119 ( .A(n51), .Y(n50) );
  INVX4 U120 ( .A(n24), .Y(n23) );
  INVX1 U121 ( .A(n19), .Y(n18) );
  INVX1 U122 ( .A(n60), .Y(n59) );
  INVX1 U123 ( .A(n40), .Y(n39) );
  INVX1 U124 ( .A(n10), .Y(n11) );
  INVX1 U125 ( .A(n36), .Y(n35) );
  INVX2 U126 ( .A(n80), .Y(n79) );
  INVX2 U127 ( .A(n76), .Y(n75) );
  INVX2 U128 ( .A(B[5]), .Y(n72) );
  INVX2 U129 ( .A(n70), .Y(n69) );
  INVX2 U130 ( .A(n66), .Y(n65) );
  INVX2 U131 ( .A(B[9]), .Y(n62) );
  INVX2 U132 ( .A(B[29]), .Y(n5) );
  INVX2 U133 ( .A(B[13]), .Y(n49) );
  INVX2 U134 ( .A(B[15]), .Y(n45) );
  INVX2 U135 ( .A(B[16]), .Y(n42) );
  INVX2 U136 ( .A(B[20]), .Y(n34) );
  INVX2 U137 ( .A(n30), .Y(n31) );
  INVX2 U138 ( .A(B[26]), .Y(n16) );
endmodule


module poly5_DW_mult_uns_35 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n8, n13, n18, n23, n28, n33, n38, n68, n80, n84, n89, n98, n107, n116,
         n125, n134, n143, n152, n163, n164, n168, n179, n184, n194, n195,
         n210, n211, n227, n228, n232, n242, n243, n258, n259, n275, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n333, n334, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n439, n443, n447, n451, n455, n459,
         n463, n467, n471, n475, n479, n483, n487, n491, n495, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n548, n549, n551, n553, n554, n555, n557, n559, n560, n561, n562,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n596, n599, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n709, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n723, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n764, n766, n767, n768,
         n769, n770, n772, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n804,
         n806, n807, n808, n810, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n830,
         n832, n833, n834, n835, n836, n838, n840, n841, n843, n846, n848,
         n850, n851, n852, n854, n856, n858, n859, n860, n861, n862, n868,
         n869, n870, n872, n876, n878, n879, n883, n884, n885, n886, n888,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2240, n2242, n2244, n2246, n2248, n2250, n2252, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020;

  NAND2X1 OR_NOTi ( .A(n3013), .B(n3015), .Y(n2725) );
  INVX2 U21 ( .A(n387), .Y(n275) );
  OAI21X1 AO21i ( .A(a[0]), .B(n275), .C(n3015), .Y(n2206) );
  NAND2X1 OR_NOTi1 ( .A(n3013), .B(n292), .Y(n2692) );
  INVX2 U15 ( .A(n340), .Y(n258) );
  OAI21X1 AO21i1 ( .A(n258), .B(n259), .C(n292), .Y(n2172) );
  NAND2X1 OR_NOTi2 ( .A(n3013), .B(n295), .Y(n2659) );
  INVX2 U25 ( .A(n393), .Y(n243) );
  INVX2 U18 ( .A(n343), .Y(n242) );
  OAI21X1 AO21i2 ( .A(n242), .B(n243), .C(n295), .Y(n2138) );
  NAND2X1 OR_NOTi3 ( .A(n3013), .B(n297), .Y(n2626) );
  INVX2 U33 ( .A(n2808), .Y(n228) );
  INVX2 U27 ( .A(n396), .Y(n227) );
  OAI21X1 AO21i3 ( .A(n232), .B(n227), .C(n228), .Y(n2104) );
  NAND2X1 OR_NOTi4 ( .A(n3013), .B(n301), .Y(n2593) );
  INVX2 U29 ( .A(n399), .Y(n211) );
  INVX2 U114 ( .A(n349), .Y(n210) );
  OAI21X1 AO21i4 ( .A(n210), .B(n211), .C(n301), .Y(n2070) );
  NAND2X1 OR_NOTi5 ( .A(n3013), .B(n304), .Y(n2560) );
  INVX2 U211 ( .A(n402), .Y(n195) );
  INVX2 U117 ( .A(n352), .Y(n194) );
  OAI21X1 AO21i5 ( .A(n194), .B(n195), .C(n303), .Y(n2036) );
  NAND2X1 OR_NOTi6 ( .A(n3013), .B(n307), .Y(n2527) );
  OAI21X1 AO21i6 ( .A(n184), .B(n179), .C(n307), .Y(n2002) );
  NAND2X1 OR_NOTi7 ( .A(n3013), .B(n310), .Y(n2494) );
  INVX2 U122 ( .A(n358), .Y(n168) );
  INVX2 U37 ( .A(n2804), .Y(n164) );
  INVX2 U215 ( .A(n408), .Y(n163) );
  OAI21X1 AO21i7 ( .A(n168), .B(n163), .C(n164), .Y(n1968) );
  NAND2X1 OR_NOTi8 ( .A(n3013), .B(n313), .Y(n2461) );
  INVX2 U125 ( .A(n361), .Y(n152) );
  NAND2X1 OR_NOTi9 ( .A(n3013), .B(n316), .Y(n2428) );
  NAND2X1 OR_NOTi10 ( .A(n3013), .B(n319), .Y(n2397) );
  INVX2 U129 ( .A(n367), .Y(n134) );
  NAND2X1 OR_NOTi11 ( .A(n3013), .B(n322), .Y(n2368) );
  INVX2 U131 ( .A(n370), .Y(n125) );
  NAND2X1 OR_NOTi12 ( .A(n3013), .B(n323), .Y(n2341) );
  NAND2X1 OR_NOTi13 ( .A(n3013), .B(n328), .Y(n2316) );
  INVX2 U135 ( .A(n376), .Y(n107) );
  NAND2X1 OR_NOTi14 ( .A(n3013), .B(n331), .Y(n2293) );
  INVX2 U137 ( .A(n379), .Y(n98) );
  NAND2X1 OR_NOTi15 ( .A(n3013), .B(n334), .Y(n2272) );
  XOR2X1 U225 ( .A(n1759), .B(n918), .Y(n80) );
  XOR2X1 U141 ( .A(n1852), .B(n80), .Y(n899) );
  XOR2X1 U226 ( .A(n1768), .B(n1828), .Y(n68) );
  XOR2X1 U142 ( .A(n1786), .B(n68), .Y(n898) );
  XOR2X1 U227 ( .A(n1906), .B(n1806), .Y(n38) );
  XOR2X1 U143 ( .A(n1878), .B(n38), .Y(n897) );
  XOR2X1 U228 ( .A(n1968), .B(n1936), .Y(n33) );
  XOR2X1 U144 ( .A(n899), .B(n33), .Y(n896) );
  XOR2X1 U229 ( .A(n914), .B(n916), .Y(n28) );
  XOR2X1 U145 ( .A(n912), .B(n28), .Y(n895) );
  XOR2X1 U230 ( .A(n898), .B(n897), .Y(n23) );
  XOR2X1 U146 ( .A(n910), .B(n23), .Y(n894) );
  XOR2X1 U231 ( .A(n908), .B(n896), .Y(n18) );
  XOR2X1 U147 ( .A(n895), .B(n18), .Y(n893) );
  XOR2X1 U232 ( .A(n894), .B(n906), .Y(n13) );
  XOR2X1 U148 ( .A(n904), .B(n13), .Y(n892) );
  XOR2X1 U233 ( .A(n902), .B(n893), .Y(n8) );
  XOR2X1 U149 ( .A(n892), .B(n8), .Y(n891) );
  NAND2X1 U293 ( .A(n548), .B(n2935), .Y(n500) );
  NAND2X1 U296 ( .A(n900), .B(n891), .Y(n548) );
  XNOR2X1 U297 ( .A(n560), .B(n501), .Y(product[46]) );
  OAI21X1 U298 ( .A(n2945), .B(n499), .C(n551), .Y(n549) );
  OAI21X1 U302 ( .A(n554), .B(n582), .C(n555), .Y(n553) );
  NAND2X1 U303 ( .A(n2924), .B(n565), .Y(n554) );
  AOI21X1 U304 ( .A(n2924), .B(n566), .C(n557), .Y(n555) );
  NAND2X1 U307 ( .A(n559), .B(n2924), .Y(n501) );
  NAND2X1 U310 ( .A(n920), .B(n901), .Y(n559) );
  XNOR2X1 U311 ( .A(n569), .B(n502), .Y(product[45]) );
  OAI21X1 U312 ( .A(n561), .B(n499), .C(n562), .Y(n560) );
  NAND2X1 U313 ( .A(n565), .B(n579), .Y(n561) );
  AOI21X1 U314 ( .A(n565), .B(n580), .C(n566), .Y(n562) );
  NOR2X1 U317 ( .A(n567), .B(n574), .Y(n565) );
  OAI21X1 U318 ( .A(n567), .B(n575), .C(n568), .Y(n566) );
  NAND2X1 U319 ( .A(n568), .B(n846), .Y(n502) );
  INVX2 U320 ( .A(n567), .Y(n846) );
  NOR2X1 U321 ( .A(n921), .B(n940), .Y(n567) );
  NAND2X1 U322 ( .A(n921), .B(n940), .Y(n568) );
  XNOR2X1 U323 ( .A(n576), .B(n503), .Y(product[44]) );
  OAI21X1 U324 ( .A(n570), .B(n499), .C(n571), .Y(n569) );
  NAND2X1 U325 ( .A(n572), .B(n579), .Y(n570) );
  AOI21X1 U326 ( .A(n572), .B(n580), .C(n573), .Y(n571) );
  NAND2X1 U329 ( .A(n575), .B(n572), .Y(n503) );
  NOR2X1 U331 ( .A(n962), .B(n941), .Y(n574) );
  NAND2X1 U332 ( .A(n962), .B(n941), .Y(n575) );
  XNOR2X1 U333 ( .A(n587), .B(n504), .Y(product[43]) );
  OAI21X1 U334 ( .A(n581), .B(n499), .C(n582), .Y(n576) );
  NAND2X1 U339 ( .A(n583), .B(n601), .Y(n581) );
  AOI21X1 U340 ( .A(n583), .B(n602), .C(n584), .Y(n582) );
  NOR2X1 U341 ( .A(n585), .B(n592), .Y(n583) );
  OAI21X1 U342 ( .A(n593), .B(n585), .C(n586), .Y(n584) );
  NAND2X1 U343 ( .A(n586), .B(n848), .Y(n504) );
  INVX2 U344 ( .A(n585), .Y(n848) );
  NOR2X1 U345 ( .A(n984), .B(n963), .Y(n585) );
  NAND2X1 U346 ( .A(n984), .B(n963), .Y(n586) );
  XNOR2X1 U347 ( .A(n594), .B(n505), .Y(product[42]) );
  OAI21X1 U348 ( .A(n588), .B(n499), .C(n589), .Y(n587) );
  NAND2X1 U349 ( .A(n590), .B(n601), .Y(n588) );
  AOI21X1 U350 ( .A(n590), .B(n602), .C(n591), .Y(n589) );
  NAND2X1 U353 ( .A(n593), .B(n590), .Y(n505) );
  NOR2X1 U355 ( .A(n1008), .B(n985), .Y(n592) );
  NAND2X1 U356 ( .A(n1008), .B(n985), .Y(n593) );
  XNOR2X1 U357 ( .A(n605), .B(n506), .Y(product[41]) );
  OAI21X1 U358 ( .A(n599), .B(n499), .C(n596), .Y(n594) );
  NOR2X1 U365 ( .A(n603), .B(n606), .Y(n601) );
  OAI21X1 U366 ( .A(n607), .B(n603), .C(n604), .Y(n602) );
  NAND2X1 U367 ( .A(n604), .B(n850), .Y(n506) );
  INVX2 U368 ( .A(n603), .Y(n850) );
  NOR2X1 U369 ( .A(n1032), .B(n1009), .Y(n603) );
  NAND2X1 U370 ( .A(n1032), .B(n1009), .Y(n604) );
  XOR2X1 U371 ( .A(n499), .B(n507), .Y(product[40]) );
  OAI21X1 U372 ( .A(n606), .B(n499), .C(n607), .Y(n605) );
  NAND2X1 U373 ( .A(n607), .B(n851), .Y(n507) );
  INVX2 U374 ( .A(n606), .Y(n851) );
  NOR2X1 U375 ( .A(n1058), .B(n1033), .Y(n606) );
  NAND2X1 U376 ( .A(n1058), .B(n1033), .Y(n607) );
  XNOR2X1 U377 ( .A(n617), .B(n508), .Y(product[39]) );
  AOI21X1 U378 ( .A(n677), .B(n609), .C(n610), .Y(n608) );
  NOR2X1 U379 ( .A(n649), .B(n611), .Y(n609) );
  OAI21X1 U380 ( .A(n611), .B(n650), .C(n612), .Y(n610) );
  NAND2X1 U381 ( .A(n613), .B(n633), .Y(n611) );
  AOI21X1 U382 ( .A(n634), .B(n613), .C(n614), .Y(n612) );
  NOR2X1 U383 ( .A(n615), .B(n624), .Y(n613) );
  OAI21X1 U384 ( .A(n625), .B(n615), .C(n616), .Y(n614) );
  NAND2X1 U385 ( .A(n616), .B(n852), .Y(n508) );
  NOR2X1 U387 ( .A(n1084), .B(n1059), .Y(n615) );
  NAND2X1 U388 ( .A(n1084), .B(n1059), .Y(n616) );
  XNOR2X1 U389 ( .A(n626), .B(n509), .Y(product[38]) );
  OAI21X1 U390 ( .A(n676), .B(n618), .C(n619), .Y(n617) );
  NAND2X1 U391 ( .A(n647), .B(n620), .Y(n618) );
  AOI21X1 U392 ( .A(n648), .B(n620), .C(n621), .Y(n619) );
  NOR2X1 U393 ( .A(n622), .B(n631), .Y(n620) );
  OAI21X1 U394 ( .A(n622), .B(n632), .C(n625), .Y(n621) );
  NAND2X1 U397 ( .A(n625), .B(n623), .Y(n509) );
  NOR2X1 U399 ( .A(n1112), .B(n1085), .Y(n624) );
  NAND2X1 U400 ( .A(n1112), .B(n1085), .Y(n625) );
  XNOR2X1 U401 ( .A(n637), .B(n510), .Y(product[37]) );
  OAI21X1 U402 ( .A(n676), .B(n627), .C(n628), .Y(n626) );
  NAND2X1 U403 ( .A(n629), .B(n647), .Y(n627) );
  AOI21X1 U404 ( .A(n629), .B(n648), .C(n630), .Y(n628) );
  NOR2X1 U409 ( .A(n635), .B(n642), .Y(n633) );
  OAI21X1 U410 ( .A(n643), .B(n635), .C(n636), .Y(n634) );
  NAND2X1 U411 ( .A(n636), .B(n854), .Y(n510) );
  INVX2 U412 ( .A(n635), .Y(n854) );
  NOR2X1 U413 ( .A(n1140), .B(n1113), .Y(n635) );
  NAND2X1 U414 ( .A(n1140), .B(n1113), .Y(n636) );
  XNOR2X1 U415 ( .A(n644), .B(n511), .Y(product[36]) );
  OAI21X1 U416 ( .A(n676), .B(n638), .C(n639), .Y(n637) );
  NAND2X1 U417 ( .A(n640), .B(n647), .Y(n638) );
  AOI21X1 U418 ( .A(n640), .B(n648), .C(n641), .Y(n639) );
  NAND2X1 U421 ( .A(n643), .B(n640), .Y(n511) );
  NOR2X1 U423 ( .A(n1170), .B(n1141), .Y(n642) );
  NAND2X1 U424 ( .A(n1170), .B(n1141), .Y(n643) );
  XNOR2X1 U425 ( .A(n655), .B(n512), .Y(product[35]) );
  OAI21X1 U426 ( .A(n649), .B(n676), .C(n646), .Y(n644) );
  NAND2X1 U431 ( .A(n669), .B(n651), .Y(n649) );
  AOI21X1 U432 ( .A(n670), .B(n651), .C(n652), .Y(n650) );
  NOR2X1 U433 ( .A(n653), .B(n660), .Y(n651) );
  OAI21X1 U434 ( .A(n661), .B(n653), .C(n654), .Y(n652) );
  NAND2X1 U435 ( .A(n654), .B(n856), .Y(n512) );
  NOR2X1 U437 ( .A(n1200), .B(n1171), .Y(n653) );
  NAND2X1 U438 ( .A(n1200), .B(n1171), .Y(n654) );
  XNOR2X1 U439 ( .A(n662), .B(n513), .Y(product[34]) );
  OAI21X1 U440 ( .A(n656), .B(n676), .C(n657), .Y(n655) );
  NAND2X1 U441 ( .A(n658), .B(n665), .Y(n656) );
  AOI21X1 U442 ( .A(n658), .B(n666), .C(n659), .Y(n657) );
  NAND2X1 U445 ( .A(n661), .B(n658), .Y(n513) );
  NOR2X1 U447 ( .A(n1232), .B(n1201), .Y(n660) );
  NAND2X1 U448 ( .A(n1232), .B(n1201), .Y(n661) );
  XNOR2X1 U449 ( .A(n673), .B(n514), .Y(product[33]) );
  OAI21X1 U450 ( .A(n667), .B(n676), .C(n668), .Y(n662) );
  NOR2X1 U457 ( .A(n674), .B(n671), .Y(n669) );
  OAI21X1 U458 ( .A(n675), .B(n671), .C(n672), .Y(n670) );
  NAND2X1 U459 ( .A(n672), .B(n858), .Y(n514) );
  NOR2X1 U461 ( .A(n1263), .B(n1233), .Y(n671) );
  NAND2X1 U462 ( .A(n1263), .B(n1233), .Y(n672) );
  XOR2X1 U463 ( .A(n676), .B(n515), .Y(product[32]) );
  OAI21X1 U464 ( .A(n674), .B(n676), .C(n675), .Y(n673) );
  NAND2X1 U465 ( .A(n675), .B(n859), .Y(n515) );
  INVX2 U466 ( .A(n674), .Y(n859) );
  NOR2X1 U467 ( .A(n1293), .B(n1264), .Y(n674) );
  NAND2X1 U468 ( .A(n1293), .B(n1264), .Y(n675) );
  XNOR2X1 U469 ( .A(n684), .B(n516), .Y(product[31]) );
  INVX4 U470 ( .A(n677), .Y(n676) );
  OAI21X1 U471 ( .A(n698), .B(n678), .C(n679), .Y(n677) );
  NAND2X1 U472 ( .A(n688), .B(n680), .Y(n678) );
  AOI21X1 U473 ( .A(n689), .B(n680), .C(n681), .Y(n679) );
  NOR2X1 U474 ( .A(n685), .B(n682), .Y(n680) );
  OAI21X1 U475 ( .A(n686), .B(n682), .C(n683), .Y(n681) );
  NAND2X1 U476 ( .A(n683), .B(n860), .Y(n516) );
  NOR2X1 U478 ( .A(n1323), .B(n1294), .Y(n682) );
  NAND2X1 U479 ( .A(n1323), .B(n1294), .Y(n683) );
  XOR2X1 U480 ( .A(n687), .B(n517), .Y(product[30]) );
  OAI21X1 U481 ( .A(n685), .B(n687), .C(n686), .Y(n684) );
  NAND2X1 U482 ( .A(n686), .B(n861), .Y(n517) );
  INVX2 U483 ( .A(n685), .Y(n861) );
  NOR2X1 U484 ( .A(n1351), .B(n1324), .Y(n685) );
  NAND2X1 U485 ( .A(n1351), .B(n1324), .Y(n686) );
  XOR2X1 U486 ( .A(n692), .B(n518), .Y(product[29]) );
  AOI21X1 U487 ( .A(n688), .B(n697), .C(n689), .Y(n687) );
  NOR2X1 U488 ( .A(n695), .B(n690), .Y(n688) );
  OAI21X1 U489 ( .A(n696), .B(n690), .C(n691), .Y(n689) );
  NAND2X1 U490 ( .A(n691), .B(n862), .Y(n518) );
  INVX2 U491 ( .A(n690), .Y(n862) );
  NOR2X1 U492 ( .A(n1379), .B(n1352), .Y(n690) );
  NAND2X1 U493 ( .A(n1379), .B(n1352), .Y(n691) );
  XNOR2X1 U494 ( .A(n697), .B(n519), .Y(product[28]) );
  AOI21X1 U495 ( .A(n693), .B(n697), .C(n694), .Y(n692) );
  NAND2X1 U498 ( .A(n696), .B(n693), .Y(n519) );
  NOR2X1 U500 ( .A(n1405), .B(n1380), .Y(n695) );
  NAND2X1 U501 ( .A(n1405), .B(n1380), .Y(n696) );
  AOI21X1 U504 ( .A(n699), .B(n727), .C(n700), .Y(n698) );
  NOR2X1 U505 ( .A(n713), .B(n701), .Y(n699) );
  OAI21X1 U506 ( .A(n714), .B(n701), .C(n702), .Y(n700) );
  NAND2X1 U507 ( .A(n2923), .B(n703), .Y(n701) );
  AOI21X1 U508 ( .A(n709), .B(n703), .C(n704), .Y(n702) );
  NOR2X1 U513 ( .A(n1431), .B(n1406), .Y(n705) );
  NAND2X1 U514 ( .A(n1431), .B(n1406), .Y(n706) );
  XNOR2X1 U515 ( .A(n712), .B(n521), .Y(product[26]) );
  AOI21X1 U516 ( .A(n2923), .B(n712), .C(n709), .Y(n707) );
  NAND2X1 U519 ( .A(n711), .B(n2923), .Y(n521) );
  NAND2X1 U522 ( .A(n1455), .B(n1432), .Y(n711) );
  XNOR2X1 U523 ( .A(n719), .B(n522), .Y(product[25]) );
  OAI21X1 U524 ( .A(n713), .B(n726), .C(n714), .Y(n712) );
  NAND2X1 U525 ( .A(n2926), .B(n715), .Y(n713) );
  AOI21X1 U526 ( .A(n723), .B(n715), .C(n716), .Y(n714) );
  NAND2X1 U529 ( .A(n718), .B(n715), .Y(n522) );
  NOR2X1 U531 ( .A(n1479), .B(n1456), .Y(n717) );
  NAND2X1 U532 ( .A(n1479), .B(n1456), .Y(n718) );
  XOR2X1 U533 ( .A(n726), .B(n523), .Y(product[24]) );
  OAI21X1 U534 ( .A(n720), .B(n726), .C(n725), .Y(n719) );
  NAND2X1 U539 ( .A(n725), .B(n2926), .Y(n523) );
  NAND2X1 U542 ( .A(n1501), .B(n1480), .Y(n725) );
  XNOR2X1 U543 ( .A(n734), .B(n524), .Y(product[23]) );
  OAI21X1 U545 ( .A(n748), .B(n728), .C(n729), .Y(n727) );
  NAND2X1 U546 ( .A(n738), .B(n730), .Y(n728) );
  AOI21X1 U547 ( .A(n739), .B(n730), .C(n731), .Y(n729) );
  NOR2X1 U548 ( .A(n735), .B(n732), .Y(n730) );
  OAI21X1 U549 ( .A(n736), .B(n732), .C(n733), .Y(n731) );
  NAND2X1 U550 ( .A(n733), .B(n868), .Y(n524) );
  INVX2 U551 ( .A(n732), .Y(n868) );
  NOR2X1 U552 ( .A(n1523), .B(n1502), .Y(n732) );
  NAND2X1 U553 ( .A(n1523), .B(n1502), .Y(n733) );
  XOR2X1 U554 ( .A(n737), .B(n525), .Y(product[22]) );
  OAI21X1 U555 ( .A(n735), .B(n737), .C(n736), .Y(n734) );
  NAND2X1 U556 ( .A(n736), .B(n869), .Y(n525) );
  INVX2 U557 ( .A(n735), .Y(n869) );
  NOR2X1 U558 ( .A(n1543), .B(n1524), .Y(n735) );
  NAND2X1 U559 ( .A(n1543), .B(n1524), .Y(n736) );
  XOR2X1 U560 ( .A(n742), .B(n526), .Y(product[21]) );
  AOI21X1 U561 ( .A(n738), .B(n747), .C(n739), .Y(n737) );
  NOR2X1 U562 ( .A(n745), .B(n740), .Y(n738) );
  OAI21X1 U563 ( .A(n746), .B(n740), .C(n741), .Y(n739) );
  NAND2X1 U564 ( .A(n741), .B(n870), .Y(n526) );
  INVX2 U565 ( .A(n740), .Y(n870) );
  NOR2X1 U566 ( .A(n1563), .B(n1544), .Y(n740) );
  NAND2X1 U567 ( .A(n1563), .B(n1544), .Y(n741) );
  XNOR2X1 U568 ( .A(n747), .B(n527), .Y(product[20]) );
  AOI21X1 U569 ( .A(n743), .B(n747), .C(n744), .Y(n742) );
  NAND2X1 U572 ( .A(n746), .B(n743), .Y(n527) );
  NOR2X1 U574 ( .A(n1581), .B(n1564), .Y(n745) );
  NAND2X1 U575 ( .A(n1581), .B(n1564), .Y(n746) );
  XNOR2X1 U576 ( .A(n753), .B(n528), .Y(product[19]) );
  AOI21X1 U578 ( .A(n749), .B(n768), .C(n750), .Y(n748) );
  NOR2X1 U579 ( .A(n751), .B(n754), .Y(n749) );
  OAI21X1 U580 ( .A(n751), .B(n755), .C(n752), .Y(n750) );
  NAND2X1 U581 ( .A(n752), .B(n872), .Y(n528) );
  INVX2 U582 ( .A(n751), .Y(n872) );
  NOR2X1 U583 ( .A(n1599), .B(n1582), .Y(n751) );
  NAND2X1 U584 ( .A(n1599), .B(n1582), .Y(n752) );
  XNOR2X1 U585 ( .A(n760), .B(n529), .Y(product[18]) );
  OAI21X1 U586 ( .A(n754), .B(n767), .C(n755), .Y(n753) );
  NAND2X1 U587 ( .A(n2925), .B(n756), .Y(n754) );
  AOI21X1 U588 ( .A(n764), .B(n756), .C(n757), .Y(n755) );
  NAND2X1 U591 ( .A(n759), .B(n756), .Y(n529) );
  NOR2X1 U593 ( .A(n1615), .B(n1600), .Y(n758) );
  NAND2X1 U594 ( .A(n1615), .B(n1600), .Y(n759) );
  XOR2X1 U595 ( .A(n767), .B(n530), .Y(product[17]) );
  OAI21X1 U596 ( .A(n761), .B(n767), .C(n766), .Y(n760) );
  NAND2X1 U601 ( .A(n766), .B(n2925), .Y(n530) );
  NAND2X1 U604 ( .A(n1631), .B(n1616), .Y(n766) );
  XOR2X1 U605 ( .A(n775), .B(n531), .Y(product[16]) );
  OAI21X1 U607 ( .A(n786), .B(n769), .C(n770), .Y(n768) );
  NAND2X1 U608 ( .A(n2922), .B(n776), .Y(n769) );
  AOI21X1 U609 ( .A(n2922), .B(n777), .C(n772), .Y(n770) );
  NAND2X1 U612 ( .A(n774), .B(n2922), .Y(n531) );
  NAND2X1 U615 ( .A(n1645), .B(n1632), .Y(n774) );
  XOR2X1 U616 ( .A(n780), .B(n532), .Y(product[15]) );
  AOI21X1 U617 ( .A(n776), .B(n785), .C(n777), .Y(n775) );
  NOR2X1 U618 ( .A(n783), .B(n778), .Y(n776) );
  OAI21X1 U619 ( .A(n784), .B(n778), .C(n779), .Y(n777) );
  NAND2X1 U620 ( .A(n779), .B(n876), .Y(n532) );
  INVX2 U621 ( .A(n778), .Y(n876) );
  NOR2X1 U622 ( .A(n1659), .B(n1646), .Y(n778) );
  NAND2X1 U623 ( .A(n1659), .B(n1646), .Y(n779) );
  XNOR2X1 U624 ( .A(n785), .B(n533), .Y(product[14]) );
  AOI21X1 U625 ( .A(n781), .B(n785), .C(n782), .Y(n780) );
  NAND2X1 U628 ( .A(n784), .B(n781), .Y(n533) );
  NOR2X1 U630 ( .A(n1671), .B(n1660), .Y(n783) );
  NAND2X1 U631 ( .A(n1671), .B(n1660), .Y(n784) );
  XNOR2X1 U632 ( .A(n791), .B(n534), .Y(product[13]) );
  AOI21X1 U634 ( .A(n787), .B(n795), .C(n788), .Y(n786) );
  NOR2X1 U635 ( .A(n792), .B(n789), .Y(n787) );
  OAI21X1 U636 ( .A(n793), .B(n789), .C(n790), .Y(n788) );
  NAND2X1 U637 ( .A(n790), .B(n878), .Y(n534) );
  INVX2 U638 ( .A(n789), .Y(n878) );
  NOR2X1 U639 ( .A(n1683), .B(n1672), .Y(n789) );
  NAND2X1 U640 ( .A(n1683), .B(n1672), .Y(n790) );
  XOR2X1 U641 ( .A(n794), .B(n535), .Y(product[12]) );
  OAI21X1 U642 ( .A(n792), .B(n794), .C(n793), .Y(n791) );
  NAND2X1 U643 ( .A(n793), .B(n879), .Y(n535) );
  INVX2 U644 ( .A(n792), .Y(n879) );
  NOR2X1 U645 ( .A(n1693), .B(n1684), .Y(n792) );
  NAND2X1 U646 ( .A(n1693), .B(n1684), .Y(n793) );
  XOR2X1 U647 ( .A(n802), .B(n536), .Y(product[11]) );
  OAI21X1 U649 ( .A(n796), .B(n808), .C(n797), .Y(n795) );
  NAND2X1 U650 ( .A(n2921), .B(n798), .Y(n796) );
  AOI21X1 U651 ( .A(n804), .B(n798), .C(n799), .Y(n797) );
  NAND2X1 U654 ( .A(n801), .B(n798), .Y(n536) );
  NOR2X1 U656 ( .A(n1703), .B(n1694), .Y(n800) );
  NAND2X1 U657 ( .A(n1703), .B(n1694), .Y(n801) );
  XNOR2X1 U658 ( .A(n807), .B(n537), .Y(product[10]) );
  AOI21X1 U659 ( .A(n2921), .B(n807), .C(n804), .Y(n802) );
  NAND2X1 U662 ( .A(n806), .B(n2921), .Y(n537) );
  NAND2X1 U665 ( .A(n1711), .B(n1704), .Y(n806) );
  XNOR2X1 U666 ( .A(n813), .B(n538), .Y(product[9]) );
  AOI21X1 U668 ( .A(n2920), .B(n813), .C(n810), .Y(n808) );
  NAND2X1 U671 ( .A(n812), .B(n2920), .Y(n538) );
  NAND2X1 U674 ( .A(n1719), .B(n1712), .Y(n812) );
  XOR2X1 U675 ( .A(n816), .B(n539), .Y(product[8]) );
  OAI21X1 U676 ( .A(n814), .B(n816), .C(n815), .Y(n813) );
  NAND2X1 U677 ( .A(n815), .B(n883), .Y(n539) );
  INVX2 U678 ( .A(n814), .Y(n883) );
  NOR2X1 U679 ( .A(n1725), .B(n1720), .Y(n814) );
  NAND2X1 U680 ( .A(n1725), .B(n1720), .Y(n815) );
  XNOR2X1 U681 ( .A(n821), .B(n540), .Y(product[7]) );
  AOI21X1 U682 ( .A(n825), .B(n817), .C(n818), .Y(n816) );
  NOR2X1 U683 ( .A(n822), .B(n819), .Y(n817) );
  OAI21X1 U684 ( .A(n823), .B(n819), .C(n820), .Y(n818) );
  NAND2X1 U685 ( .A(n820), .B(n884), .Y(n540) );
  INVX2 U686 ( .A(n819), .Y(n884) );
  NOR2X1 U687 ( .A(n1731), .B(n1726), .Y(n819) );
  NAND2X1 U688 ( .A(n1731), .B(n1726), .Y(n820) );
  XOR2X1 U689 ( .A(n541), .B(n824), .Y(product[6]) );
  OAI21X1 U690 ( .A(n822), .B(n824), .C(n823), .Y(n821) );
  NAND2X1 U691 ( .A(n823), .B(n885), .Y(n541) );
  INVX2 U692 ( .A(n822), .Y(n885) );
  NOR2X1 U693 ( .A(n1735), .B(n1732), .Y(n822) );
  NAND2X1 U694 ( .A(n1735), .B(n1732), .Y(n823) );
  XOR2X1 U695 ( .A(n542), .B(n828), .Y(product[5]) );
  OAI21X1 U697 ( .A(n826), .B(n828), .C(n827), .Y(n825) );
  NAND2X1 U698 ( .A(n827), .B(n886), .Y(n542) );
  INVX2 U699 ( .A(n826), .Y(n886) );
  NOR2X1 U700 ( .A(n1739), .B(n1736), .Y(n826) );
  NAND2X1 U701 ( .A(n1739), .B(n1736), .Y(n827) );
  XNOR2X1 U702 ( .A(n543), .B(n833), .Y(product[4]) );
  AOI21X1 U703 ( .A(n833), .B(n2919), .C(n830), .Y(n828) );
  NAND2X1 U706 ( .A(n832), .B(n2919), .Y(n543) );
  NAND2X1 U709 ( .A(n1741), .B(n1740), .Y(n832) );
  XOR2X1 U710 ( .A(n544), .B(n836), .Y(product[3]) );
  OAI21X1 U711 ( .A(n834), .B(n836), .C(n835), .Y(n833) );
  NAND2X1 U712 ( .A(n835), .B(n888), .Y(n544) );
  INVX2 U713 ( .A(n834), .Y(n888) );
  NOR2X1 U714 ( .A(n1757), .B(n1742), .Y(n834) );
  NAND2X1 U715 ( .A(n1757), .B(n1742), .Y(n835) );
  XNOR2X1 U716 ( .A(n545), .B(n841), .Y(product[2]) );
  AOI21X1 U717 ( .A(n841), .B(n2927), .C(n838), .Y(n836) );
  NAND2X1 U720 ( .A(n840), .B(n2927), .Y(n545) );
  NAND2X1 U723 ( .A(n2237), .B(n2953), .Y(n840) );
  NAND2X1 U729 ( .A(n1758), .B(n2238), .Y(n843) );
  FAX1 U730 ( .A(n905), .B(n922), .C(n903), .YC(n900), .YS(n901) );
  FAX1 U731 ( .A(n926), .B(n907), .C(n924), .YC(n902), .YS(n903) );
  FAX1 U732 ( .A(n911), .B(n928), .C(n909), .YC(n904), .YS(n905) );
  FAX1 U733 ( .A(n915), .B(n932), .C(n930), .YC(n906), .YS(n907) );
  FAX1 U734 ( .A(n934), .B(n917), .C(n913), .YC(n908), .YS(n909) );
  FAX1 U735 ( .A(n1829), .B(n938), .C(n936), .YC(n910), .YS(n911) );
  FAX1 U736 ( .A(n1853), .B(n1787), .C(n1807), .YC(n912), .YS(n913) );
  FAX1 U737 ( .A(n1907), .B(n1769), .C(n1879), .YC(n914), .YS(n915) );
  FAX1 U738 ( .A(n919), .B(n1969), .C(n1937), .YC(n916), .YS(n917) );
  INVX2 U739 ( .A(n918), .Y(n919) );
  FAX1 U740 ( .A(n925), .B(n942), .C(n923), .YC(n920), .YS(n921) );
  FAX1 U741 ( .A(n946), .B(n927), .C(n944), .YC(n922), .YS(n923) );
  FAX1 U742 ( .A(n948), .B(n931), .C(n929), .YC(n924), .YS(n925) );
  FAX1 U743 ( .A(n933), .B(n952), .C(n950), .YC(n926), .YS(n927) );
  FAX1 U744 ( .A(n954), .B(n935), .C(n937), .YC(n928), .YS(n929) );
  FAX1 U745 ( .A(n958), .B(n956), .C(n939), .YC(n930), .YS(n931) );
  FAX1 U746 ( .A(n1970), .B(n1938), .C(n2002), .YC(n932), .YS(n933) );
  FAX1 U747 ( .A(n1788), .B(n1908), .C(n1830), .YC(n934), .YS(n935) );
  FAX1 U748 ( .A(n1854), .B(n1770), .C(n1808), .YC(n936), .YS(n937) );
  FAX1 U749 ( .A(n960), .B(n1760), .C(n1880), .YC(n938), .YS(n939) );
  FAX1 U750 ( .A(n945), .B(n964), .C(n943), .YC(n940), .YS(n941) );
  FAX1 U751 ( .A(n968), .B(n947), .C(n966), .YC(n942), .YS(n943) );
  FAX1 U752 ( .A(n970), .B(n951), .C(n949), .YC(n944), .YS(n945) );
  FAX1 U753 ( .A(n953), .B(n974), .C(n972), .YC(n946), .YS(n947) );
  FAX1 U754 ( .A(n959), .B(n955), .C(n957), .YC(n948), .YS(n949) );
  FAX1 U755 ( .A(n980), .B(n976), .C(n978), .YC(n950), .YS(n951) );
  FAX1 U756 ( .A(n1909), .B(n1881), .C(n982), .YC(n952), .YS(n953) );
  FAX1 U757 ( .A(n1855), .B(n1809), .C(n1831), .YC(n954), .YS(n955) );
  FAX1 U758 ( .A(n1939), .B(n1771), .C(n1789), .YC(n956), .YS(n957) );
  FAX1 U759 ( .A(n961), .B(n2003), .C(n1971), .YC(n958), .YS(n959) );
  INVX2 U760 ( .A(n960), .Y(n961) );
  FAX1 U761 ( .A(n988), .B(n986), .C(n965), .YC(n962), .YS(n963) );
  FAX1 U762 ( .A(n990), .B(n969), .C(n967), .YC(n964), .YS(n965) );
  FAX1 U763 ( .A(n973), .B(n971), .C(n992), .YC(n966), .YS(n967) );
  FAX1 U764 ( .A(n996), .B(n994), .C(n975), .YC(n968), .YS(n969) );
  FAX1 U765 ( .A(n977), .B(n981), .C(n979), .YC(n970), .YS(n971) );
  FAX1 U766 ( .A(n1000), .B(n998), .C(n983), .YC(n972), .YS(n973) );
  FAX1 U767 ( .A(n2036), .B(n1004), .C(n1002), .YC(n974), .YS(n975) );
  FAX1 U768 ( .A(n2004), .B(n1832), .C(n1972), .YC(n976), .YS(n977) );
  FAX1 U769 ( .A(n1910), .B(n1810), .C(n1940), .YC(n978), .YS(n979) );
  FAX1 U770 ( .A(n1856), .B(n1772), .C(n1790), .YC(n980), .YS(n981) );
  FAX1 U771 ( .A(n1006), .B(n1761), .C(n1882), .YC(n982), .YS(n983) );
  FAX1 U772 ( .A(n989), .B(n1010), .C(n987), .YC(n984), .YS(n985) );
  FAX1 U773 ( .A(n1014), .B(n991), .C(n1012), .YC(n986), .YS(n987) );
  FAX1 U774 ( .A(n995), .B(n1016), .C(n993), .YC(n988), .YS(n989) );
  FAX1 U775 ( .A(n1020), .B(n1018), .C(n997), .YC(n990), .YS(n991) );
  FAX1 U776 ( .A(n1003), .B(n1001), .C(n1022), .YC(n992), .YS(n993) );
  FAX1 U777 ( .A(n1024), .B(n1005), .C(n999), .YC(n994), .YS(n995) );
  FAX1 U778 ( .A(n1030), .B(n1028), .C(n1026), .YC(n996), .YS(n997) );
  FAX1 U779 ( .A(n1911), .B(n1857), .C(n1883), .YC(n998), .YS(n999) );
  FAX1 U780 ( .A(n1811), .B(n1941), .C(n1833), .YC(n1000), .YS(n1001) );
  FAX1 U781 ( .A(n1973), .B(n1773), .C(n1791), .YC(n1002), .YS(n1003) );
  FAX1 U782 ( .A(n1007), .B(n2037), .C(n2005), .YC(n1004), .YS(n1005) );
  INVX2 U783 ( .A(n1006), .Y(n1007) );
  FAX1 U784 ( .A(n1013), .B(n1034), .C(n1011), .YC(n1008), .YS(n1009) );
  FAX1 U785 ( .A(n1038), .B(n1015), .C(n1036), .YC(n1010), .YS(n1011) );
  FAX1 U786 ( .A(n1019), .B(n1040), .C(n1017), .YC(n1012), .YS(n1013) );
  FAX1 U787 ( .A(n1023), .B(n1042), .C(n1021), .YC(n1014), .YS(n1015) );
  FAX1 U788 ( .A(n1029), .B(n1046), .C(n1044), .YC(n1016), .YS(n1017) );
  FAX1 U789 ( .A(n1050), .B(n1025), .C(n1027), .YC(n1018), .YS(n1019) );
  FAX1 U790 ( .A(n1052), .B(n1048), .C(n1031), .YC(n1020), .YS(n1021) );
  FAX1 U791 ( .A(n2038), .B(n2070), .C(n1054), .YC(n1022), .YS(n1023) );
  FAX1 U792 ( .A(n2006), .B(n1834), .C(n1974), .YC(n1024), .YS(n1025) );
  FAX1 U793 ( .A(n1942), .B(n1774), .C(n1858), .YC(n1026), .YS(n1027) );
  FAX1 U794 ( .A(n1884), .B(n1792), .C(n1812), .YC(n1028), .YS(n1029) );
  FAX1 U795 ( .A(n1056), .B(n1762), .C(n1912), .YC(n1030), .YS(n1031) );
  FAX1 U796 ( .A(n1037), .B(n1060), .C(n1035), .YC(n1032), .YS(n1033) );
  FAX1 U797 ( .A(n1064), .B(n1039), .C(n1062), .YC(n1034), .YS(n1035) );
  FAX1 U798 ( .A(n1043), .B(n1066), .C(n1041), .YC(n1036), .YS(n1037) );
  FAX1 U799 ( .A(n1047), .B(n1045), .C(n1068), .YC(n1038), .YS(n1039) );
  FAX1 U800 ( .A(n1053), .B(n1072), .C(n1070), .YC(n1040), .YS(n1041) );
  FAX1 U801 ( .A(n1051), .B(n1049), .C(n1074), .YC(n1042), .YS(n1043) );
  FAX1 U802 ( .A(n1078), .B(n1076), .C(n1055), .YC(n1044), .YS(n1045) );
  FAX1 U803 ( .A(n1943), .B(n1082), .C(n1080), .YC(n1046), .YS(n1047) );
  FAX1 U804 ( .A(n1975), .B(n1859), .C(n1913), .YC(n1048), .YS(n1049) );
  FAX1 U805 ( .A(n1835), .B(n2007), .C(n1813), .YC(n1050), .YS(n1051) );
  FAX1 U806 ( .A(n2039), .B(n1775), .C(n1793), .YC(n1052), .YS(n1053) );
  FAX1 U807 ( .A(n1057), .B(n2071), .C(n1885), .YC(n1054), .YS(n1055) );
  INVX2 U808 ( .A(n1056), .Y(n1057) );
  FAX1 U809 ( .A(n1063), .B(n1086), .C(n1061), .YC(n1058), .YS(n1059) );
  FAX1 U810 ( .A(n1090), .B(n1065), .C(n1088), .YC(n1060), .YS(n1061) );
  FAX1 U811 ( .A(n1094), .B(n1092), .C(n1067), .YC(n1062), .YS(n1063) );
  FAX1 U812 ( .A(n1073), .B(n1071), .C(n1069), .YC(n1064), .YS(n1065) );
  FAX1 U813 ( .A(n1100), .B(n1098), .C(n1096), .YC(n1066), .YS(n1067) );
  FAX1 U814 ( .A(n1079), .B(n1081), .C(n1075), .YC(n1068), .YS(n1069) );
  FAX1 U815 ( .A(n1104), .B(n1102), .C(n1077), .YC(n1070), .YS(n1071) );
  FAX1 U816 ( .A(n1108), .B(n1106), .C(n1083), .YC(n1072), .YS(n1073) );
  FAX1 U817 ( .A(n2072), .B(n2040), .C(n2104), .YC(n1074), .YS(n1075) );
  FAX1 U818 ( .A(n1860), .B(n2008), .C(n1976), .YC(n1076), .YS(n1077) );
  FAX1 U819 ( .A(n1776), .B(n1914), .C(n1836), .YC(n1078), .YS(n1079) );
  FAX1 U820 ( .A(n1886), .B(n1794), .C(n1814), .YC(n1080), .YS(n1081) );
  FAX1 U821 ( .A(n1110), .B(n1763), .C(n1944), .YC(n1082), .YS(n1083) );
  FAX1 U822 ( .A(n1089), .B(n1114), .C(n1087), .YC(n1084), .YS(n1085) );
  FAX1 U823 ( .A(n1118), .B(n1091), .C(n1116), .YC(n1086), .YS(n1087) );
  FAX1 U824 ( .A(n1095), .B(n1120), .C(n1093), .YC(n1088), .YS(n1089) );
  FAX1 U825 ( .A(n1099), .B(n1097), .C(n1122), .YC(n1090), .YS(n1091) );
  FAX1 U826 ( .A(n1128), .B(n1126), .C(n1124), .YC(n1092), .YS(n1093) );
  FAX1 U827 ( .A(n1105), .B(n1107), .C(n1101), .YC(n1094), .YS(n1095) );
  FAX1 U828 ( .A(n1132), .B(n1109), .C(n1103), .YC(n1096), .YS(n1097) );
  FAX1 U829 ( .A(n1136), .B(n1130), .C(n1134), .YC(n1098), .YS(n1099) );
  FAX1 U830 ( .A(n1915), .B(n1861), .C(n1138), .YC(n1100), .YS(n1101) );
  FAX1 U831 ( .A(n1945), .B(n1815), .C(n1837), .YC(n1102), .YS(n1103) );
  FAX1 U832 ( .A(n2009), .B(n1795), .C(n1977), .YC(n1104), .YS(n1105) );
  FAX1 U833 ( .A(n1887), .B(n2041), .C(n1777), .YC(n1106), .YS(n1107) );
  FAX1 U834 ( .A(n1111), .B(n2105), .C(n2073), .YC(n1108), .YS(n1109) );
  INVX2 U835 ( .A(n1110), .Y(n1111) );
  FAX1 U836 ( .A(n1117), .B(n1142), .C(n1115), .YC(n1112), .YS(n1113) );
  FAX1 U837 ( .A(n1146), .B(n1119), .C(n1144), .YC(n1114), .YS(n1115) );
  FAX1 U838 ( .A(n1123), .B(n1148), .C(n1121), .YC(n1116), .YS(n1117) );
  FAX1 U839 ( .A(n1127), .B(n1125), .C(n1150), .YC(n1118), .YS(n1119) );
  FAX1 U840 ( .A(n1154), .B(n1129), .C(n1152), .YC(n1120), .YS(n1121) );
  FAX1 U841 ( .A(n1137), .B(n1135), .C(n1156), .YC(n1122), .YS(n1123) );
  FAX1 U842 ( .A(n1162), .B(n1131), .C(n1133), .YC(n1124), .YS(n1125) );
  FAX1 U843 ( .A(n1160), .B(n1164), .C(n1139), .YC(n1126), .YS(n1127) );
  FAX1 U844 ( .A(n2138), .B(n1166), .C(n1158), .YC(n1128), .YS(n1129) );
  FAX1 U845 ( .A(n2074), .B(n2106), .C(n1888), .YC(n1130), .YS(n1131) );
  FAX1 U846 ( .A(n1862), .B(n2010), .C(n2042), .YC(n1132), .YS(n1133) );
  FAX1 U847 ( .A(n1978), .B(n1796), .C(n1838), .YC(n1134), .YS(n1135) );
  FAX1 U848 ( .A(n1916), .B(n1778), .C(n1816), .YC(n1136), .YS(n1137) );
  FAX1 U849 ( .A(n1168), .B(n1764), .C(n1946), .YC(n1138), .YS(n1139) );
  FAX1 U850 ( .A(n1145), .B(n1172), .C(n1143), .YC(n1140), .YS(n1141) );
  FAX1 U851 ( .A(n1176), .B(n1147), .C(n1174), .YC(n1142), .YS(n1143) );
  FAX1 U852 ( .A(n1151), .B(n1178), .C(n1149), .YC(n1144), .YS(n1145) );
  FAX1 U853 ( .A(n1155), .B(n1153), .C(n1180), .YC(n1146), .YS(n1147) );
  FAX1 U854 ( .A(n1184), .B(n1157), .C(n1182), .YC(n1148), .YS(n1149) );
  FAX1 U855 ( .A(n1163), .B(n1188), .C(n1186), .YC(n1150), .YS(n1151) );
  FAX1 U856 ( .A(n1159), .B(n1165), .C(n1161), .YC(n1152), .YS(n1153) );
  FAX1 U857 ( .A(n1194), .B(n1196), .C(n1167), .YC(n1154), .YS(n1155) );
  FAX1 U858 ( .A(n1198), .B(n1190), .C(n1192), .YC(n1156), .YS(n1157) );
  FAX1 U859 ( .A(n1947), .B(n1863), .C(n1917), .YC(n1158), .YS(n1159) );
  FAX1 U860 ( .A(n1979), .B(n1817), .C(n1839), .YC(n1160), .YS(n1161) );
  FAX1 U861 ( .A(n2043), .B(n1797), .C(n2011), .YC(n1162), .YS(n1163) );
  FAX1 U862 ( .A(n1889), .B(n2075), .C(n1779), .YC(n1164), .YS(n1165) );
  FAX1 U863 ( .A(n1169), .B(n2139), .C(n2107), .YC(n1166), .YS(n1167) );
  INVX2 U864 ( .A(n1168), .Y(n1169) );
  FAX1 U865 ( .A(n1175), .B(n1202), .C(n1173), .YC(n1170), .YS(n1171) );
  FAX1 U866 ( .A(n1206), .B(n1177), .C(n1204), .YC(n1172), .YS(n1173) );
  FAX1 U867 ( .A(n1181), .B(n1208), .C(n1179), .YC(n1174), .YS(n1175) );
  FAX1 U868 ( .A(n1185), .B(n1183), .C(n1210), .YC(n1176), .YS(n1177) );
  FAX1 U869 ( .A(n1214), .B(n1212), .C(n1187), .YC(n1178), .YS(n1179) );
  FAX1 U870 ( .A(n1218), .B(n1189), .C(n1216), .YC(n1180), .YS(n1181) );
  FAX1 U871 ( .A(n1195), .B(n1197), .C(n1193), .YC(n1182), .YS(n1183) );
  FAX1 U872 ( .A(n1224), .B(n1222), .C(n1191), .YC(n1184), .YS(n1185) );
  FAX1 U873 ( .A(n1220), .B(n1226), .C(n1199), .YC(n1186), .YS(n1187) );
  FAX1 U874 ( .A(n2076), .B(n2172), .C(n1228), .YC(n1188), .YS(n1189) );
  FAX1 U875 ( .A(n2108), .B(n2044), .C(n2140), .YC(n1190), .YS(n1191) );
  FAX1 U876 ( .A(n1864), .B(n1948), .C(n1890), .YC(n1192), .YS(n1193) );
  FAX1 U877 ( .A(n2012), .B(n1840), .C(n1818), .YC(n1194), .YS(n1195) );
  FAX1 U878 ( .A(n1918), .B(n1780), .C(n1798), .YC(n1196), .YS(n1197) );
  FAX1 U879 ( .A(n2918), .B(n1765), .C(n1980), .YC(n1198), .YS(n1199) );
  FAX1 U880 ( .A(n1205), .B(n1234), .C(n1203), .YC(n1200), .YS(n1201) );
  FAX1 U881 ( .A(n1238), .B(n1207), .C(n1236), .YC(n1202), .YS(n1203) );
  FAX1 U882 ( .A(n1240), .B(n1211), .C(n1209), .YC(n1204), .YS(n1205) );
  FAX1 U883 ( .A(n1217), .B(n1213), .C(n1242), .YC(n1206), .YS(n1207) );
  FAX1 U884 ( .A(n1246), .B(n1244), .C(n1215), .YC(n1208), .YS(n1209) );
  FAX1 U885 ( .A(n1250), .B(n1248), .C(n1219), .YC(n1210), .YS(n1211) );
  FAX1 U886 ( .A(n1225), .B(n1227), .C(n1223), .YC(n1212), .YS(n1213) );
  FAX1 U887 ( .A(n1256), .B(n1254), .C(n1221), .YC(n1214), .YS(n1215) );
  FAX1 U888 ( .A(n1252), .B(n1258), .C(n1229), .YC(n1216), .YS(n1217) );
  FAX1 U889 ( .A(n1981), .B(n2013), .C(n1260), .YC(n1218), .YS(n1219) );
  FAX1 U890 ( .A(n2045), .B(n1919), .C(n1949), .YC(n1220), .YS(n1221) );
  FAX1 U891 ( .A(n1865), .B(n2077), .C(n1891), .YC(n1222), .YS(n1223) );
  FAX1 U892 ( .A(n2109), .B(n1819), .C(n1841), .YC(n1224), .YS(n1225) );
  FAX1 U893 ( .A(n2141), .B(n1781), .C(n1799), .YC(n1226), .YS(n1227) );
  FAX1 U894 ( .A(n1766), .B(n1231), .C(n2173), .YC(n1228), .YS(n1229) );
  FAX1 U896 ( .A(n1237), .B(n1265), .C(n1235), .YC(n1232), .YS(n1233) );
  FAX1 U897 ( .A(n1269), .B(n1239), .C(n1267), .YC(n1234), .YS(n1235) );
  FAX1 U898 ( .A(n1271), .B(n1243), .C(n1241), .YC(n1236), .YS(n1237) );
  FAX1 U899 ( .A(n1247), .B(n1245), .C(n1273), .YC(n1238), .YS(n1239) );
  FAX1 U900 ( .A(n1251), .B(n1275), .C(n1249), .YC(n1240), .YS(n1241) );
  FAX1 U901 ( .A(n1255), .B(n1279), .C(n1277), .YC(n1242), .YS(n1243) );
  FAX1 U902 ( .A(n1257), .B(n1259), .C(n1281), .YC(n1244), .YS(n1245) );
  FAX1 U903 ( .A(n1285), .B(n1261), .C(n1253), .YC(n1246), .YS(n1247) );
  FAX1 U904 ( .A(n1283), .B(n1289), .C(n1287), .YC(n1248), .YS(n1249) );
  FAX1 U905 ( .A(n2110), .B(n2206), .C(n1291), .YC(n1250), .YS(n1251) );
  FAX1 U906 ( .A(n2142), .B(n2078), .C(n2174), .YC(n1252), .YS(n1253) );
  FAX1 U907 ( .A(n1892), .B(n1982), .C(n1920), .YC(n1254), .YS(n1255) );
  FAX1 U908 ( .A(n2046), .B(n1866), .C(n1842), .YC(n1256), .YS(n1257) );
  FAX1 U909 ( .A(n1950), .B(n1782), .C(n1820), .YC(n1258), .YS(n1259) );
  FAX1 U910 ( .A(n1262), .B(n2014), .C(n1800), .YC(n1260), .YS(n1261) );
  INVX2 U911 ( .A(n2918), .Y(n1262) );
  FAX1 U912 ( .A(n1268), .B(n1295), .C(n1266), .YC(n1263), .YS(n1264) );
  FAX1 U913 ( .A(n1272), .B(n1270), .C(n1297), .YC(n1265), .YS(n1266) );
  FAX1 U914 ( .A(n1274), .B(n1301), .C(n1299), .YC(n1267), .YS(n1268) );
  FAX1 U915 ( .A(n1278), .B(n1276), .C(n1303), .YC(n1269), .YS(n1270) );
  FAX1 U916 ( .A(n1307), .B(n1305), .C(n1280), .YC(n1271), .YS(n1272) );
  FAX1 U917 ( .A(n1288), .B(n1282), .C(n1309), .YC(n1273), .YS(n1274) );
  FAX1 U918 ( .A(n1284), .B(n1290), .C(n1286), .YC(n1275), .YS(n1276) );
  FAX1 U919 ( .A(n1311), .B(n1315), .C(n1292), .YC(n1277), .YS(n1278) );
  FAX1 U920 ( .A(n1313), .B(n1319), .C(n1317), .YC(n1279), .YS(n1280) );
  FAX1 U921 ( .A(n2015), .B(n2047), .C(n1321), .YC(n1281), .YS(n1282) );
  FAX1 U922 ( .A(n2079), .B(n1921), .C(n1951), .YC(n1283), .YS(n1284) );
  FAX1 U923 ( .A(n2111), .B(n1867), .C(n1893), .YC(n1285), .YS(n1286) );
  FAX1 U924 ( .A(n1983), .B(n2143), .C(n1843), .YC(n1287), .YS(n1288) );
  FAX1 U925 ( .A(n2175), .B(n1801), .C(n1821), .YC(n1289), .YS(n1290) );
  FAX1 U926 ( .A(n2928), .B(n2207), .C(n1783), .YC(n1291), .YS(n1292) );
  FAX1 U927 ( .A(n1298), .B(n1325), .C(n1296), .YC(n1293), .YS(n1294) );
  FAX1 U928 ( .A(n1302), .B(n1300), .C(n1327), .YC(n1295), .YS(n1296) );
  FAX1 U929 ( .A(n1304), .B(n1331), .C(n1329), .YC(n1297), .YS(n1298) );
  FAX1 U930 ( .A(n1308), .B(n1333), .C(n1306), .YC(n1299), .YS(n1300) );
  FAX1 U931 ( .A(n1337), .B(n1310), .C(n1335), .YC(n1301), .YS(n1302) );
  FAX1 U932 ( .A(n1314), .B(n1316), .C(n1339), .YC(n1303), .YS(n1304) );
  FAX1 U933 ( .A(n1312), .B(n1320), .C(n1318), .YC(n1305), .YS(n1306) );
  FAX1 U934 ( .A(n1341), .B(n1345), .C(n1343), .YC(n1307), .YS(n1308) );
  FAX1 U935 ( .A(n1322), .B(n1349), .C(n1347), .YC(n1309), .YS(n1310) );
  FAX1 U936 ( .A(n1868), .B(n2016), .C(n1922), .YC(n1311), .YS(n1312) );
  FAX1 U937 ( .A(n2048), .B(n1822), .C(n1844), .YC(n1313), .YS(n1314) );
  FAX1 U938 ( .A(n1894), .B(n2112), .C(n2080), .YC(n1315), .YS(n1316) );
  FAX1 U939 ( .A(n1984), .B(n2176), .C(n2144), .YC(n1317), .YS(n1318) );
  FAX1 U940 ( .A(n1952), .B(n1784), .C(n1802), .YC(n1319), .YS(n1320) );
  HAX1 U941 ( .A(n2208), .B(n1743), .YC(n1321), .YS(n1322) );
  FAX1 U942 ( .A(n1328), .B(n1353), .C(n1326), .YC(n1323), .YS(n1324) );
  FAX1 U943 ( .A(n1332), .B(n1330), .C(n1355), .YC(n1325), .YS(n1326) );
  FAX1 U944 ( .A(n1334), .B(n1359), .C(n1357), .YC(n1327), .YS(n1328) );
  FAX1 U945 ( .A(n1361), .B(n1338), .C(n1336), .YC(n1329), .YS(n1330) );
  FAX1 U946 ( .A(n1365), .B(n1340), .C(n1363), .YC(n1331), .YS(n1332) );
  FAX1 U947 ( .A(n1344), .B(n1346), .C(n1367), .YC(n1333), .YS(n1334) );
  FAX1 U948 ( .A(n1350), .B(n1342), .C(n1348), .YC(n1335), .YS(n1336) );
  FAX1 U949 ( .A(n1371), .B(n1375), .C(n1373), .YC(n1337), .YS(n1338) );
  FAX1 U950 ( .A(n2948), .B(n1377), .C(n1369), .YC(n1339), .YS(n1340) );
  FAX1 U951 ( .A(n2017), .B(n1953), .C(n1985), .YC(n1341), .YS(n1342) );
  FAX1 U952 ( .A(n2049), .B(n1895), .C(n1923), .YC(n1343), .YS(n1344) );
  FAX1 U953 ( .A(n2081), .B(n1845), .C(n1869), .YC(n1345), .YS(n1346) );
  FAX1 U954 ( .A(n2145), .B(n1823), .C(n2113), .YC(n1347), .YS(n1348) );
  FAX1 U955 ( .A(n2209), .B(n2177), .C(n1803), .YC(n1349), .YS(n1350) );
  FAX1 U956 ( .A(n1356), .B(n1381), .C(n1354), .YC(n1351), .YS(n1352) );
  FAX1 U957 ( .A(n1385), .B(n1358), .C(n1383), .YC(n1353), .YS(n1354) );
  FAX1 U958 ( .A(n1362), .B(n1387), .C(n1360), .YC(n1355), .YS(n1356) );
  FAX1 U959 ( .A(n1366), .B(n1389), .C(n1364), .YC(n1357), .YS(n1358) );
  FAX1 U960 ( .A(n1368), .B(n1393), .C(n1391), .YC(n1359), .YS(n1360) );
  FAX1 U961 ( .A(n1374), .B(n1376), .C(n1395), .YC(n1361), .YS(n1362) );
  FAX1 U962 ( .A(n1401), .B(n1370), .C(n1372), .YC(n1363), .YS(n1364) );
  FAX1 U963 ( .A(n1403), .B(n1397), .C(n1399), .YC(n1365), .YS(n1366) );
  FAX1 U964 ( .A(n2018), .B(n2050), .C(n1378), .YC(n1367), .YS(n1368) );
  FAX1 U965 ( .A(n2082), .B(n1924), .C(n1954), .YC(n1369), .YS(n1370) );
  FAX1 U966 ( .A(n1846), .B(n1870), .C(n1824), .YC(n1371), .YS(n1372) );
  FAX1 U967 ( .A(n1896), .B(n2114), .C(n1804), .YC(n1373), .YS(n1374) );
  FAX1 U968 ( .A(n1986), .B(n2178), .C(n2146), .YC(n1375), .YS(n1376) );
  HAX1 U969 ( .A(n2210), .B(n1744), .YC(n1377), .YS(n1378) );
  FAX1 U970 ( .A(n1384), .B(n1407), .C(n1382), .YC(n1379), .YS(n1380) );
  FAX1 U971 ( .A(n1411), .B(n1386), .C(n1409), .YC(n1381), .YS(n1382) );
  FAX1 U972 ( .A(n1390), .B(n1413), .C(n1388), .YC(n1383), .YS(n1384) );
  FAX1 U973 ( .A(n1394), .B(n1415), .C(n1392), .YC(n1385), .YS(n1386) );
  FAX1 U974 ( .A(n1396), .B(n1419), .C(n1417), .YC(n1387), .YS(n1388) );
  FAX1 U975 ( .A(n1400), .B(n1398), .C(n1402), .YC(n1389), .YS(n1390) );
  FAX1 U976 ( .A(n1421), .B(n1423), .C(n1404), .YC(n1391), .YS(n1392) );
  FAX1 U977 ( .A(n1429), .B(n1427), .C(n1425), .YC(n1393), .YS(n1394) );
  FAX1 U978 ( .A(n2019), .B(n1987), .C(n2933), .YC(n1395), .YS(n1396) );
  FAX1 U979 ( .A(n2051), .B(n1925), .C(n1955), .YC(n1397), .YS(n1398) );
  FAX1 U980 ( .A(n2083), .B(n1871), .C(n1897), .YC(n1399), .YS(n1400) );
  FAX1 U981 ( .A(n2147), .B(n1847), .C(n2115), .YC(n1401), .YS(n1402) );
  FAX1 U982 ( .A(n2211), .B(n2179), .C(n1825), .YC(n1403), .YS(n1404) );
  FAX1 U983 ( .A(n1410), .B(n1433), .C(n1408), .YC(n1405), .YS(n1406) );
  FAX1 U984 ( .A(n1414), .B(n1412), .C(n1435), .YC(n1407), .YS(n1408) );
  FAX1 U985 ( .A(n1416), .B(n1439), .C(n1437), .YC(n1409), .YS(n1410) );
  FAX1 U986 ( .A(n1420), .B(n1441), .C(n1418), .YC(n1411), .YS(n1412) );
  FAX1 U987 ( .A(n1424), .B(n1445), .C(n1443), .YC(n1413), .YS(n1414) );
  FAX1 U988 ( .A(n1422), .B(n1428), .C(n1426), .YC(n1415), .YS(n1416) );
  FAX1 U989 ( .A(n1447), .B(n1449), .C(n1451), .YC(n1417), .YS(n1418) );
  FAX1 U990 ( .A(n2084), .B(n1430), .C(n1453), .YC(n1419), .YS(n1420) );
  FAX1 U991 ( .A(n2116), .B(n1956), .C(n2052), .YC(n1421), .YS(n1422) );
  FAX1 U992 ( .A(n2148), .B(n1898), .C(n1926), .YC(n1423), .YS(n1424) );
  FAX1 U993 ( .A(n2020), .B(n1872), .C(n2180), .YC(n1425), .YS(n1426) );
  FAX1 U994 ( .A(n1988), .B(n1848), .C(n1826), .YC(n1427), .YS(n1428) );
  HAX1 U995 ( .A(n2212), .B(n1745), .YC(n1429), .YS(n1430) );
  FAX1 U996 ( .A(n1436), .B(n1457), .C(n1434), .YC(n1431), .YS(n1432) );
  FAX1 U997 ( .A(n1461), .B(n1459), .C(n1438), .YC(n1433), .YS(n1434) );
  FAX1 U998 ( .A(n1444), .B(n1442), .C(n1440), .YC(n1435), .YS(n1436) );
  FAX1 U999 ( .A(n1467), .B(n1465), .C(n1463), .YC(n1437), .YS(n1438) );
  FAX1 U1000 ( .A(n1452), .B(n1450), .C(n1446), .YC(n1439), .YS(n1440) );
  FAX1 U1001 ( .A(n1473), .B(n1454), .C(n1448), .YC(n1441), .YS(n1442) );
  FAX1 U1002 ( .A(n1475), .B(n1469), .C(n1471), .YC(n1443), .YS(n1444) );
  FAX1 U1003 ( .A(n2053), .B(n2957), .C(n1477), .YC(n1445), .YS(n1446) );
  FAX1 U1004 ( .A(n2085), .B(n1989), .C(n2021), .YC(n1447), .YS(n1448) );
  FAX1 U1005 ( .A(n2117), .B(n1927), .C(n1957), .YC(n1449), .YS(n1450) );
  FAX1 U1006 ( .A(n2149), .B(n1873), .C(n1899), .YC(n1451), .YS(n1452) );
  FAX1 U1007 ( .A(n2213), .B(n2181), .C(n1849), .YC(n1453), .YS(n1454) );
  FAX1 U1008 ( .A(n1460), .B(n1481), .C(n1458), .YC(n1455), .YS(n1456) );
  FAX1 U1009 ( .A(n1485), .B(n1483), .C(n1462), .YC(n1457), .YS(n1458) );
  FAX1 U1010 ( .A(n1487), .B(n1466), .C(n1464), .YC(n1459), .YS(n1460) );
  FAX1 U1011 ( .A(n1491), .B(n1489), .C(n1468), .YC(n1461), .YS(n1462) );
  FAX1 U1012 ( .A(n1472), .B(n1476), .C(n1474), .YC(n1463), .YS(n1464) );
  FAX1 U1013 ( .A(n1495), .B(n1493), .C(n1470), .YC(n1465), .YS(n1466) );
  FAX1 U1014 ( .A(n1478), .B(n1499), .C(n1497), .YC(n1467), .YS(n1468) );
  FAX1 U1015 ( .A(n2086), .B(n1990), .C(n2054), .YC(n1469), .YS(n1470) );
  FAX1 U1016 ( .A(n2118), .B(n1900), .C(n1958), .YC(n1471), .YS(n1472) );
  FAX1 U1017 ( .A(n1928), .B(n1850), .C(n1874), .YC(n1473), .YS(n1474) );
  FAX1 U1018 ( .A(n2022), .B(n2182), .C(n2150), .YC(n1475), .YS(n1476) );
  HAX1 U1019 ( .A(n2214), .B(n1746), .YC(n1477), .YS(n1478) );
  FAX1 U1020 ( .A(n1484), .B(n1503), .C(n1482), .YC(n1479), .YS(n1480) );
  FAX1 U1021 ( .A(n1507), .B(n1486), .C(n1505), .YC(n1481), .YS(n1482) );
  FAX1 U1022 ( .A(n1509), .B(n1490), .C(n1488), .YC(n1483), .YS(n1484) );
  FAX1 U1023 ( .A(n1513), .B(n1511), .C(n1492), .YC(n1485), .YS(n1486) );
  FAX1 U1024 ( .A(n1494), .B(n1498), .C(n1496), .YC(n1487), .YS(n1488) );
  FAX1 U1025 ( .A(n1517), .B(n1515), .C(n1500), .YC(n1489), .YS(n1490) );
  FAX1 U1026 ( .A(n2951), .B(n1521), .C(n1519), .YC(n1491), .YS(n1492) );
  FAX1 U1027 ( .A(n2087), .B(n2023), .C(n2055), .YC(n1493), .YS(n1494) );
  FAX1 U1028 ( .A(n2119), .B(n1959), .C(n1991), .YC(n1495), .YS(n1496) );
  FAX1 U1029 ( .A(n2151), .B(n1901), .C(n1929), .YC(n1497), .YS(n1498) );
  FAX1 U1030 ( .A(n2215), .B(n2183), .C(n1875), .YC(n1499), .YS(n1500) );
  FAX1 U1031 ( .A(n1506), .B(n1525), .C(n1504), .YC(n1501), .YS(n1502) );
  FAX1 U1032 ( .A(n1529), .B(n1508), .C(n1527), .YC(n1503), .YS(n1504) );
  FAX1 U1033 ( .A(n1531), .B(n1512), .C(n1510), .YC(n1505), .YS(n1506) );
  FAX1 U1034 ( .A(n1518), .B(n1514), .C(n1533), .YC(n1507), .YS(n1508) );
  FAX1 U1035 ( .A(n1516), .B(n1520), .C(n1535), .YC(n1509), .YS(n1510) );
  FAX1 U1036 ( .A(n1541), .B(n1539), .C(n1537), .YC(n1511), .YS(n1512) );
  FAX1 U1037 ( .A(n2088), .B(n1992), .C(n1522), .YC(n1513), .YS(n1514) );
  FAX1 U1038 ( .A(n2120), .B(n1930), .C(n1960), .YC(n1515), .YS(n1516) );
  FAX1 U1039 ( .A(n2056), .B(n2184), .C(n2152), .YC(n1517), .YS(n1518) );
  FAX1 U1040 ( .A(n2024), .B(n1876), .C(n1902), .YC(n1519), .YS(n1520) );
  HAX1 U1041 ( .A(n2216), .B(n1747), .YC(n1521), .YS(n1522) );
  FAX1 U1042 ( .A(n1528), .B(n1545), .C(n1526), .YC(n1523), .YS(n1524) );
  FAX1 U1043 ( .A(n1532), .B(n1530), .C(n1547), .YC(n1525), .YS(n1526) );
  FAX1 U1044 ( .A(n1551), .B(n1534), .C(n1549), .YC(n1527), .YS(n1528) );
  FAX1 U1045 ( .A(n1540), .B(n1536), .C(n1553), .YC(n1529), .YS(n1530) );
  FAX1 U1046 ( .A(n1555), .B(n1542), .C(n1538), .YC(n1531), .YS(n1532) );
  FAX1 U1047 ( .A(n1561), .B(n1559), .C(n1557), .YC(n1533), .YS(n1534) );
  FAX1 U1048 ( .A(n2089), .B(n2057), .C(n2932), .YC(n1535), .YS(n1536) );
  FAX1 U1049 ( .A(n2121), .B(n1993), .C(n2025), .YC(n1537), .YS(n1538) );
  FAX1 U1050 ( .A(n2153), .B(n1931), .C(n1961), .YC(n1539), .YS(n1540) );
  FAX1 U1051 ( .A(n2217), .B(n2185), .C(n1903), .YC(n1541), .YS(n1542) );
  FAX1 U1052 ( .A(n1548), .B(n1565), .C(n1546), .YC(n1543), .YS(n1544) );
  FAX1 U1053 ( .A(n1552), .B(n1550), .C(n1567), .YC(n1545), .YS(n1546) );
  FAX1 U1054 ( .A(n1571), .B(n1554), .C(n1569), .YC(n1547), .YS(n1548) );
  FAX1 U1055 ( .A(n1558), .B(n1560), .C(n1573), .YC(n1549), .YS(n1550) );
  FAX1 U1056 ( .A(n1577), .B(n1575), .C(n1556), .YC(n1551), .YS(n1552) );
  FAX1 U1057 ( .A(n1994), .B(n1562), .C(n1579), .YC(n1553), .YS(n1554) );
  FAX1 U1058 ( .A(n2058), .B(n1932), .C(n1904), .YC(n1555), .YS(n1556) );
  FAX1 U1059 ( .A(n1962), .B(n2122), .C(n2090), .YC(n1557), .YS(n1558) );
  FAX1 U1060 ( .A(n2026), .B(n2186), .C(n2154), .YC(n1559), .YS(n1560) );
  HAX1 U1061 ( .A(n2218), .B(n1748), .YC(n1561), .YS(n1562) );
  FAX1 U1062 ( .A(n1568), .B(n1583), .C(n1566), .YC(n1563), .YS(n1564) );
  FAX1 U1063 ( .A(n1572), .B(n1570), .C(n1585), .YC(n1565), .YS(n1566) );
  FAX1 U1064 ( .A(n1574), .B(n1589), .C(n1587), .YC(n1567), .YS(n1568) );
  FAX1 U1065 ( .A(n1580), .B(n1576), .C(n1578), .YC(n1569), .YS(n1570) );
  FAX1 U1066 ( .A(n1595), .B(n1591), .C(n1593), .YC(n1571), .YS(n1572) );
  FAX1 U1067 ( .A(n2091), .B(n2956), .C(n1597), .YC(n1573), .YS(n1574) );
  FAX1 U1068 ( .A(n2123), .B(n2027), .C(n2059), .YC(n1575), .YS(n1576) );
  FAX1 U1069 ( .A(n2155), .B(n1963), .C(n1995), .YC(n1577), .YS(n1578) );
  FAX1 U1070 ( .A(n2219), .B(n2187), .C(n1933), .YC(n1579), .YS(n1580) );
  FAX1 U1071 ( .A(n1586), .B(n1601), .C(n1584), .YC(n1581), .YS(n1582) );
  FAX1 U1072 ( .A(n1590), .B(n1588), .C(n1603), .YC(n1583), .YS(n1584) );
  FAX1 U1073 ( .A(n1596), .B(n1607), .C(n1605), .YC(n1585), .YS(n1586) );
  FAX1 U1074 ( .A(n1609), .B(n1592), .C(n1594), .YC(n1587), .YS(n1588) );
  FAX1 U1075 ( .A(n1598), .B(n1613), .C(n1611), .YC(n1589), .YS(n1590) );
  FAX1 U1076 ( .A(n2156), .B(n2028), .C(n2124), .YC(n1591), .YS(n1592) );
  FAX1 U1077 ( .A(n2092), .B(n2188), .C(n1996), .YC(n1593), .YS(n1594) );
  FAX1 U1078 ( .A(n2060), .B(n1934), .C(n1964), .YC(n1595), .YS(n1596) );
  HAX1 U1079 ( .A(n2220), .B(n1749), .YC(n1597), .YS(n1598) );
  FAX1 U1080 ( .A(n1604), .B(n1617), .C(n1602), .YC(n1599), .YS(n1600) );
  FAX1 U1081 ( .A(n1608), .B(n1606), .C(n1619), .YC(n1601), .YS(n1602) );
  FAX1 U1082 ( .A(n1612), .B(n1623), .C(n1621), .YC(n1603), .YS(n1604) );
  FAX1 U1083 ( .A(n1625), .B(n1614), .C(n1610), .YC(n1605), .YS(n1606) );
  FAX1 U1084 ( .A(n2946), .B(n1629), .C(n1627), .YC(n1607), .YS(n1608) );
  FAX1 U1085 ( .A(n2125), .B(n2061), .C(n2093), .YC(n1609), .YS(n1610) );
  FAX1 U1086 ( .A(n2157), .B(n1997), .C(n2029), .YC(n1611), .YS(n1612) );
  FAX1 U1087 ( .A(n2221), .B(n2189), .C(n1965), .YC(n1613), .YS(n1614) );
  FAX1 U1088 ( .A(n1620), .B(n1633), .C(n1618), .YC(n1615), .YS(n1616) );
  FAX1 U1089 ( .A(n1637), .B(n1622), .C(n1635), .YC(n1617), .YS(n1618) );
  FAX1 U1090 ( .A(n1628), .B(n1639), .C(n1624), .YC(n1619), .YS(n1620) );
  FAX1 U1091 ( .A(n1643), .B(n1641), .C(n1626), .YC(n1621), .YS(n1622) );
  FAX1 U1092 ( .A(n2094), .B(n2030), .C(n1630), .YC(n1623), .YS(n1624) );
  FAX1 U1093 ( .A(n2126), .B(n1966), .C(n1998), .YC(n1625), .YS(n1626) );
  FAX1 U1094 ( .A(n2062), .B(n2190), .C(n2158), .YC(n1627), .YS(n1628) );
  HAX1 U1095 ( .A(n2222), .B(n1750), .YC(n1629), .YS(n1630) );
  FAX1 U1096 ( .A(n1636), .B(n1647), .C(n1634), .YC(n1631), .YS(n1632) );
  FAX1 U1097 ( .A(n1651), .B(n1649), .C(n1638), .YC(n1633), .YS(n1634) );
  FAX1 U1098 ( .A(n1644), .B(n1642), .C(n1640), .YC(n1635), .YS(n1636) );
  FAX1 U1099 ( .A(n1657), .B(n1655), .C(n1653), .YC(n1637), .YS(n1638) );
  FAX1 U1100 ( .A(n2127), .B(n2095), .C(n2931), .YC(n1639), .YS(n1640) );
  FAX1 U1101 ( .A(n2159), .B(n2031), .C(n2063), .YC(n1641), .YS(n1642) );
  FAX1 U1102 ( .A(n2223), .B(n2191), .C(n1999), .YC(n1643), .YS(n1644) );
  FAX1 U1103 ( .A(n1650), .B(n1661), .C(n1648), .YC(n1645), .YS(n1646) );
  FAX1 U1104 ( .A(n1665), .B(n1663), .C(n1652), .YC(n1647), .YS(n1648) );
  FAX1 U1105 ( .A(n1667), .B(n1654), .C(n1656), .YC(n1649), .YS(n1650) );
  FAX1 U1106 ( .A(n2160), .B(n1658), .C(n1669), .YC(n1651), .YS(n1652) );
  FAX1 U1107 ( .A(n2192), .B(n2064), .C(n2128), .YC(n1653), .YS(n1654) );
  FAX1 U1108 ( .A(n2096), .B(n2000), .C(n2032), .YC(n1655), .YS(n1656) );
  HAX1 U1109 ( .A(n2224), .B(n1751), .YC(n1657), .YS(n1658) );
  FAX1 U1110 ( .A(n1664), .B(n1673), .C(n1662), .YC(n1659), .YS(n1660) );
  FAX1 U1111 ( .A(n1668), .B(n1666), .C(n1675), .YC(n1661), .YS(n1662) );
  FAX1 U1112 ( .A(n1679), .B(n1677), .C(n1670), .YC(n1663), .YS(n1664) );
  FAX1 U1113 ( .A(n2129), .B(n2947), .C(n1681), .YC(n1665), .YS(n1666) );
  FAX1 U1114 ( .A(n2161), .B(n2065), .C(n2097), .YC(n1667), .YS(n1668) );
  FAX1 U1115 ( .A(n2225), .B(n2193), .C(n2033), .YC(n1669), .YS(n1670) );
  FAX1 U1116 ( .A(n1676), .B(n1685), .C(n1674), .YC(n1671), .YS(n1672) );
  FAX1 U1117 ( .A(n1678), .B(n1680), .C(n1687), .YC(n1673), .YS(n1674) );
  FAX1 U1118 ( .A(n1682), .B(n1691), .C(n1689), .YC(n1675), .YS(n1676) );
  FAX1 U1119 ( .A(n2130), .B(n2034), .C(n2066), .YC(n1677), .YS(n1678) );
  FAX1 U1120 ( .A(n2098), .B(n2194), .C(n2162), .YC(n1679), .YS(n1680) );
  HAX1 U1121 ( .A(n2226), .B(n1752), .YC(n1681), .YS(n1682) );
  FAX1 U1122 ( .A(n1688), .B(n1695), .C(n1686), .YC(n1683), .YS(n1684) );
  FAX1 U1123 ( .A(n1692), .B(n1690), .C(n1697), .YC(n1685), .YS(n1686) );
  FAX1 U1124 ( .A(n2949), .B(n1701), .C(n1699), .YC(n1687), .YS(n1688) );
  FAX1 U1125 ( .A(n2163), .B(n2099), .C(n2131), .YC(n1689), .YS(n1690) );
  FAX1 U1126 ( .A(n2227), .B(n2195), .C(n2067), .YC(n1691), .YS(n1692) );
  FAX1 U1127 ( .A(n1698), .B(n1705), .C(n1696), .YC(n1693), .YS(n1694) );
  FAX1 U1128 ( .A(n1709), .B(n1700), .C(n1707), .YC(n1695), .YS(n1696) );
  FAX1 U1129 ( .A(n2164), .B(n2100), .C(n1702), .YC(n1697), .YS(n1698) );
  FAX1 U1130 ( .A(n2132), .B(n2068), .C(n2196), .YC(n1699), .YS(n1700) );
  HAX1 U1131 ( .A(n2228), .B(n1753), .YC(n1701), .YS(n1702) );
  FAX1 U1132 ( .A(n1708), .B(n1713), .C(n1706), .YC(n1703), .YS(n1704) );
  FAX1 U1133 ( .A(n1717), .B(n1715), .C(n1710), .YC(n1705), .YS(n1706) );
  FAX1 U1134 ( .A(n2165), .B(n2133), .C(n2930), .YC(n1707), .YS(n1708) );
  FAX1 U1135 ( .A(n2229), .B(n2197), .C(n2101), .YC(n1709), .YS(n1710) );
  FAX1 U1136 ( .A(n1716), .B(n1721), .C(n1714), .YC(n1711), .YS(n1712) );
  FAX1 U1137 ( .A(n2198), .B(n1718), .C(n1723), .YC(n1713), .YS(n1714) );
  FAX1 U1138 ( .A(n2134), .B(n2102), .C(n2166), .YC(n1715), .YS(n1716) );
  HAX1 U1139 ( .A(n2230), .B(n1754), .YC(n1717), .YS(n1718) );
  FAX1 U1140 ( .A(n1727), .B(n1724), .C(n1722), .YC(n1719), .YS(n1720) );
  FAX1 U1141 ( .A(n2167), .B(n2950), .C(n1729), .YC(n1721), .YS(n1722) );
  FAX1 U1142 ( .A(n2231), .B(n2199), .C(n2135), .YC(n1723), .YS(n1724) );
  FAX1 U1143 ( .A(n1730), .B(n1733), .C(n1728), .YC(n1725), .YS(n1726) );
  FAX1 U1144 ( .A(n2200), .B(n2136), .C(n2168), .YC(n1727), .YS(n1728) );
  HAX1 U1145 ( .A(n2232), .B(n1755), .YC(n1729), .YS(n1730) );
  FAX1 U1146 ( .A(n2952), .B(n1737), .C(n1734), .YC(n1731), .YS(n1732) );
  FAX1 U1147 ( .A(n2233), .B(n2201), .C(n2169), .YC(n1733), .YS(n1734) );
  FAX1 U1148 ( .A(n2202), .B(n2170), .C(n1738), .YC(n1735), .YS(n1736) );
  HAX1 U1149 ( .A(n2234), .B(n1756), .YC(n1737), .YS(n1738) );
  FAX1 U1150 ( .A(n2235), .B(n2203), .C(n2929), .YC(n1739), .YS(n1740) );
  HAX1 U1151 ( .A(n2236), .B(n2204), .YC(n1741), .YS(n1742) );
  NOR2X1 U1152 ( .A(n2990), .B(n383), .Y(n1759) );
  NOR2X1 U1153 ( .A(n2240), .B(n383), .Y(n918) );
  NOR2X1 U1154 ( .A(n2993), .B(n383), .Y(n1760) );
  NOR2X1 U1155 ( .A(n2242), .B(n383), .Y(n960) );
  NOR2X1 U1156 ( .A(n2996), .B(n383), .Y(n1761) );
  NOR2X1 U1157 ( .A(n2244), .B(n383), .Y(n1006) );
  NOR2X1 U1158 ( .A(n2999), .B(n383), .Y(n1762) );
  NOR2X1 U1159 ( .A(n2246), .B(n383), .Y(n1056) );
  NOR2X1 U1160 ( .A(n3002), .B(n383), .Y(n1763) );
  NOR2X1 U1161 ( .A(n2248), .B(n383), .Y(n1110) );
  NOR2X1 U1162 ( .A(n3005), .B(n383), .Y(n1764) );
  NOR2X1 U1163 ( .A(n2250), .B(n383), .Y(n1168) );
  NOR2X1 U1164 ( .A(n3008), .B(n383), .Y(n1765) );
  NOR2X1 U1165 ( .A(n2252), .B(n383), .Y(n1766) );
  NOR2X1 U1166 ( .A(n3010), .B(n383), .Y(n1230) );
  INVX2 U1168 ( .A(n463), .Y(n2240) );
  INVX2 U1170 ( .A(n459), .Y(n2242) );
  INVX2 U1172 ( .A(n455), .Y(n2244) );
  INVX2 U1174 ( .A(n451), .Y(n2246) );
  INVX2 U1176 ( .A(n447), .Y(n2248) );
  INVX2 U1178 ( .A(n443), .Y(n2250) );
  INVX2 U1180 ( .A(n439), .Y(n2252) );
  OAI22X1 U1182 ( .A(n382), .B(n2272), .C(n2796), .D(n432), .Y(n1743) );
  OAI22X1 U1183 ( .A(n2254), .B(n381), .C(n2255), .D(n431), .Y(n1768) );
  OAI22X1 U1184 ( .A(n2255), .B(n381), .C(n2256), .D(n431), .Y(n1769) );
  OAI22X1 U1185 ( .A(n2256), .B(n381), .C(n2257), .D(n431), .Y(n1770) );
  OAI22X1 U1186 ( .A(n2257), .B(n381), .C(n2258), .D(n431), .Y(n1771) );
  OAI22X1 U1187 ( .A(n2258), .B(n381), .C(n2259), .D(n431), .Y(n1772) );
  OAI22X1 U1188 ( .A(n2259), .B(n381), .C(n2260), .D(n431), .Y(n1773) );
  OAI22X1 U1189 ( .A(n2260), .B(n380), .C(n2261), .D(n431), .Y(n1774) );
  OAI22X1 U1190 ( .A(n2261), .B(n380), .C(n2262), .D(n431), .Y(n1775) );
  OAI22X1 U1191 ( .A(n2262), .B(n380), .C(n2263), .D(n430), .Y(n1776) );
  OAI22X1 U1192 ( .A(n2263), .B(n380), .C(n2264), .D(n431), .Y(n1777) );
  OAI22X1 U1193 ( .A(n2264), .B(n380), .C(n2265), .D(n430), .Y(n1778) );
  OAI22X1 U1194 ( .A(n2265), .B(n380), .C(n2266), .D(n430), .Y(n1779) );
  OAI22X1 U1195 ( .A(n2266), .B(n380), .C(n2267), .D(n430), .Y(n1780) );
  OAI22X1 U1196 ( .A(n2267), .B(n380), .C(n2268), .D(n430), .Y(n1781) );
  OAI22X1 U1197 ( .A(n2268), .B(n380), .C(n2269), .D(n430), .Y(n1782) );
  OAI22X1 U1198 ( .A(n2269), .B(n380), .C(n2270), .D(n430), .Y(n1783) );
  OAI22X1 U1199 ( .A(n2270), .B(n380), .C(n2271), .D(n430), .Y(n1784) );
  XNOR2X1 U1200 ( .A(n333), .B(n2986), .Y(n2254) );
  XNOR2X1 U1201 ( .A(n333), .B(n467), .Y(n2255) );
  XNOR2X1 U1202 ( .A(n333), .B(n2988), .Y(n2256) );
  XNOR2X1 U1203 ( .A(n333), .B(n463), .Y(n2257) );
  XNOR2X1 U1204 ( .A(n333), .B(n2991), .Y(n2258) );
  XNOR2X1 U1205 ( .A(n333), .B(n459), .Y(n2259) );
  XNOR2X1 U1206 ( .A(n333), .B(n2994), .Y(n2260) );
  XNOR2X1 U1207 ( .A(n333), .B(n455), .Y(n2261) );
  XNOR2X1 U1208 ( .A(n333), .B(n2997), .Y(n2262) );
  XNOR2X1 U1209 ( .A(n2968), .B(n451), .Y(n2263) );
  XNOR2X1 U1210 ( .A(n334), .B(n3000), .Y(n2264) );
  XNOR2X1 U1211 ( .A(n2968), .B(n447), .Y(n2265) );
  XNOR2X1 U1212 ( .A(n2968), .B(n3003), .Y(n2266) );
  XNOR2X1 U1213 ( .A(n2967), .B(n443), .Y(n2267) );
  XNOR2X1 U1214 ( .A(n2967), .B(n3006), .Y(n2268) );
  XNOR2X1 U1215 ( .A(n2968), .B(n439), .Y(n2269) );
  XNOR2X1 U1216 ( .A(n2967), .B(n3009), .Y(n2270) );
  XNOR2X1 U1217 ( .A(n334), .B(n3012), .Y(n2271) );
  OAI22X1 U1218 ( .A(n379), .B(n2293), .C(n2797), .D(n429), .Y(n1744) );
  OAI22X1 U1219 ( .A(n2273), .B(n378), .C(n2274), .D(n428), .Y(n1786) );
  OAI22X1 U1220 ( .A(n2274), .B(n378), .C(n2275), .D(n428), .Y(n1787) );
  OAI22X1 U1221 ( .A(n2275), .B(n378), .C(n2276), .D(n428), .Y(n1788) );
  OAI22X1 U1222 ( .A(n2276), .B(n378), .C(n2277), .D(n428), .Y(n1789) );
  OAI22X1 U1223 ( .A(n2277), .B(n378), .C(n2278), .D(n428), .Y(n1790) );
  OAI22X1 U1224 ( .A(n2278), .B(n378), .C(n2279), .D(n428), .Y(n1791) );
  OAI22X1 U1225 ( .A(n2279), .B(n378), .C(n2280), .D(n428), .Y(n1792) );
  OAI22X1 U1226 ( .A(n2280), .B(n378), .C(n2281), .D(n428), .Y(n1793) );
  OAI22X1 U1227 ( .A(n2281), .B(n377), .C(n2282), .D(n428), .Y(n1794) );
  OAI22X1 U1228 ( .A(n2282), .B(n377), .C(n2283), .D(n427), .Y(n1795) );
  OAI22X1 U1229 ( .A(n2283), .B(n377), .C(n2284), .D(n427), .Y(n1796) );
  OAI22X1 U1230 ( .A(n2284), .B(n377), .C(n2285), .D(n427), .Y(n1797) );
  OAI22X1 U1231 ( .A(n2285), .B(n377), .C(n2286), .D(n427), .Y(n1798) );
  OAI22X1 U1232 ( .A(n2286), .B(n377), .C(n2287), .D(n427), .Y(n1799) );
  OAI22X1 U1233 ( .A(n2287), .B(n377), .C(n2288), .D(n427), .Y(n1800) );
  OAI22X1 U1234 ( .A(n2288), .B(n377), .C(n2289), .D(n427), .Y(n1801) );
  OAI22X1 U1235 ( .A(n2289), .B(n377), .C(n2290), .D(n427), .Y(n1802) );
  OAI22X1 U1236 ( .A(n2290), .B(n377), .C(n2291), .D(n427), .Y(n1803) );
  OAI22X1 U1237 ( .A(n2291), .B(n377), .C(n2292), .D(n427), .Y(n1804) );
  XNOR2X1 U1238 ( .A(n2914), .B(b[19]), .Y(n2273) );
  XNOR2X1 U1239 ( .A(n2914), .B(n471), .Y(n2274) );
  XNOR2X1 U1240 ( .A(n2914), .B(n2986), .Y(n2275) );
  XNOR2X1 U1241 ( .A(n2914), .B(n467), .Y(n2276) );
  XNOR2X1 U1242 ( .A(n2914), .B(n2988), .Y(n2277) );
  XNOR2X1 U1243 ( .A(n2914), .B(n463), .Y(n2278) );
  XNOR2X1 U1244 ( .A(n2914), .B(n2991), .Y(n2279) );
  XNOR2X1 U1245 ( .A(n2914), .B(n459), .Y(n2280) );
  XNOR2X1 U1246 ( .A(n2913), .B(n2994), .Y(n2281) );
  XNOR2X1 U1247 ( .A(n2913), .B(n455), .Y(n2282) );
  XNOR2X1 U1248 ( .A(n2913), .B(n2997), .Y(n2283) );
  XNOR2X1 U1249 ( .A(n2959), .B(n451), .Y(n2284) );
  XNOR2X1 U1250 ( .A(n2960), .B(n3000), .Y(n2285) );
  XNOR2X1 U1251 ( .A(n2960), .B(n447), .Y(n2286) );
  XNOR2X1 U1252 ( .A(n2958), .B(n3003), .Y(n2287) );
  XNOR2X1 U1253 ( .A(n2958), .B(n443), .Y(n2288) );
  XNOR2X1 U1254 ( .A(n2959), .B(n3006), .Y(n2289) );
  XNOR2X1 U1255 ( .A(n2959), .B(n439), .Y(n2290) );
  XNOR2X1 U1256 ( .A(n2960), .B(n3009), .Y(n2291) );
  XNOR2X1 U1257 ( .A(n2960), .B(n3011), .Y(n2292) );
  OAI22X1 U1258 ( .A(n376), .B(n2316), .C(n2798), .D(n426), .Y(n1745) );
  OAI22X1 U1259 ( .A(n2294), .B(n375), .C(n2295), .D(n425), .Y(n1806) );
  OAI22X1 U1260 ( .A(n2295), .B(n375), .C(n2296), .D(n425), .Y(n1807) );
  OAI22X1 U1261 ( .A(n2296), .B(n375), .C(n2297), .D(n425), .Y(n1808) );
  OAI22X1 U1262 ( .A(n2297), .B(n375), .C(n2298), .D(n425), .Y(n1809) );
  OAI22X1 U1263 ( .A(n2298), .B(n375), .C(n2299), .D(n425), .Y(n1810) );
  OAI22X1 U1264 ( .A(n2299), .B(n375), .C(n2300), .D(n425), .Y(n1811) );
  OAI22X1 U1265 ( .A(n2300), .B(n375), .C(n2301), .D(n425), .Y(n1812) );
  OAI22X1 U1266 ( .A(n2301), .B(n375), .C(n2302), .D(n425), .Y(n1813) );
  OAI22X1 U1267 ( .A(n2302), .B(n375), .C(n2303), .D(n425), .Y(n1814) );
  OAI22X1 U1268 ( .A(n2303), .B(n375), .C(n2304), .D(n425), .Y(n1815) );
  OAI22X1 U1269 ( .A(n2304), .B(n374), .C(n2305), .D(n425), .Y(n1816) );
  OAI22X1 U1270 ( .A(n2305), .B(n374), .C(n2306), .D(n424), .Y(n1817) );
  OAI22X1 U1271 ( .A(n2306), .B(n374), .C(n2307), .D(n424), .Y(n1818) );
  OAI22X1 U1272 ( .A(n2307), .B(n374), .C(n2308), .D(n424), .Y(n1819) );
  OAI22X1 U1273 ( .A(n2308), .B(n374), .C(n2309), .D(n424), .Y(n1820) );
  OAI22X1 U1274 ( .A(n2309), .B(n374), .C(n2310), .D(n424), .Y(n1821) );
  OAI22X1 U1275 ( .A(n2310), .B(n374), .C(n2311), .D(n424), .Y(n1822) );
  OAI22X1 U1276 ( .A(n2311), .B(n374), .C(n2312), .D(n424), .Y(n1823) );
  OAI22X1 U1277 ( .A(n2312), .B(n374), .C(n2313), .D(n424), .Y(n1824) );
  OAI22X1 U1278 ( .A(n2313), .B(n374), .C(n2314), .D(n424), .Y(n1825) );
  OAI22X1 U1279 ( .A(n2314), .B(n374), .C(n2315), .D(n424), .Y(n1826) );
  XNOR2X1 U1280 ( .A(n328), .B(n2981), .Y(n2294) );
  XNOR2X1 U1281 ( .A(n2941), .B(n475), .Y(n2295) );
  XNOR2X1 U1282 ( .A(n2942), .B(b[19]), .Y(n2296) );
  XNOR2X1 U1283 ( .A(n2941), .B(n471), .Y(n2297) );
  XNOR2X1 U1284 ( .A(n2941), .B(n2986), .Y(n2298) );
  XNOR2X1 U1285 ( .A(n2942), .B(n467), .Y(n2299) );
  XNOR2X1 U1286 ( .A(n2942), .B(n2988), .Y(n2300) );
  XNOR2X1 U1287 ( .A(n2941), .B(n463), .Y(n2301) );
  XNOR2X1 U1288 ( .A(n2942), .B(n2991), .Y(n2302) );
  XNOR2X1 U1289 ( .A(n2942), .B(n459), .Y(n2303) );
  XNOR2X1 U1290 ( .A(n2941), .B(n2994), .Y(n2304) );
  XNOR2X1 U1291 ( .A(n2940), .B(n455), .Y(n2305) );
  XNOR2X1 U1292 ( .A(n2940), .B(n2997), .Y(n2306) );
  XNOR2X1 U1293 ( .A(n2964), .B(n451), .Y(n2307) );
  XNOR2X1 U1294 ( .A(n2964), .B(n3000), .Y(n2308) );
  XNOR2X1 U1295 ( .A(n2966), .B(n447), .Y(n2309) );
  XNOR2X1 U1296 ( .A(n2965), .B(n3003), .Y(n2310) );
  XNOR2X1 U1297 ( .A(n2966), .B(n443), .Y(n2311) );
  XNOR2X1 U1298 ( .A(n2965), .B(n3006), .Y(n2312) );
  XNOR2X1 U1299 ( .A(n2965), .B(n439), .Y(n2313) );
  XNOR2X1 U1300 ( .A(n2966), .B(n3009), .Y(n2314) );
  XNOR2X1 U1301 ( .A(n2966), .B(n3012), .Y(n2315) );
  OAI22X1 U1302 ( .A(n373), .B(n2341), .C(n2799), .D(n423), .Y(n1746) );
  OAI22X1 U1303 ( .A(n2317), .B(n372), .C(n2318), .D(n423), .Y(n1828) );
  OAI22X1 U1304 ( .A(n2318), .B(n372), .C(n2319), .D(n422), .Y(n1829) );
  OAI22X1 U1305 ( .A(n2319), .B(n372), .C(n2320), .D(n422), .Y(n1830) );
  OAI22X1 U1306 ( .A(n2320), .B(n372), .C(n2321), .D(n422), .Y(n1831) );
  OAI22X1 U1307 ( .A(n2321), .B(n372), .C(n2322), .D(n422), .Y(n1832) );
  OAI22X1 U1308 ( .A(n2322), .B(n372), .C(n2323), .D(n422), .Y(n1833) );
  OAI22X1 U1309 ( .A(n2323), .B(n372), .C(n2324), .D(n422), .Y(n1834) );
  OAI22X1 U1310 ( .A(n2324), .B(n372), .C(n2325), .D(n422), .Y(n1835) );
  OAI22X1 U1311 ( .A(n2325), .B(n372), .C(n2326), .D(n422), .Y(n1836) );
  OAI22X1 U1312 ( .A(n2326), .B(n372), .C(n2327), .D(n422), .Y(n1837) );
  OAI22X1 U1313 ( .A(n2327), .B(n372), .C(n2328), .D(n422), .Y(n1838) );
  OAI22X1 U1314 ( .A(n2328), .B(n372), .C(n2329), .D(n422), .Y(n1839) );
  OAI22X1 U1315 ( .A(n2329), .B(n371), .C(n2330), .D(n422), .Y(n1840) );
  OAI22X1 U1316 ( .A(n2330), .B(n371), .C(n2331), .D(n421), .Y(n1841) );
  OAI22X1 U1317 ( .A(n2331), .B(n371), .C(n2332), .D(n421), .Y(n1842) );
  OAI22X1 U1318 ( .A(n2332), .B(n371), .C(n2333), .D(n421), .Y(n1843) );
  OAI22X1 U1319 ( .A(n2333), .B(n371), .C(n2334), .D(n421), .Y(n1844) );
  OAI22X1 U1320 ( .A(n2334), .B(n371), .C(n2335), .D(n421), .Y(n1845) );
  OAI22X1 U1321 ( .A(n2335), .B(n371), .C(n2336), .D(n421), .Y(n1846) );
  OAI22X1 U1322 ( .A(n2336), .B(n371), .C(n2337), .D(n421), .Y(n1847) );
  OAI22X1 U1323 ( .A(n2337), .B(n371), .C(n2338), .D(n421), .Y(n1848) );
  OAI22X1 U1324 ( .A(n2338), .B(n371), .C(n2339), .D(n421), .Y(n1849) );
  OAI22X1 U1325 ( .A(n2339), .B(n371), .C(n2340), .D(n421), .Y(n1850) );
  XNOR2X1 U1326 ( .A(n323), .B(n2978), .Y(n2317) );
  XNOR2X1 U1327 ( .A(n2937), .B(n479), .Y(n2318) );
  XNOR2X1 U1328 ( .A(n2936), .B(n2981), .Y(n2319) );
  XNOR2X1 U1329 ( .A(n2962), .B(n475), .Y(n2320) );
  XNOR2X1 U1330 ( .A(n2963), .B(n2983), .Y(n2321) );
  XNOR2X1 U1331 ( .A(n2963), .B(n471), .Y(n2322) );
  XNOR2X1 U1332 ( .A(n2962), .B(n2986), .Y(n2323) );
  XNOR2X1 U1333 ( .A(n2962), .B(n467), .Y(n2324) );
  XNOR2X1 U1334 ( .A(n2963), .B(n2988), .Y(n2325) );
  XNOR2X1 U1335 ( .A(n2963), .B(n463), .Y(n2326) );
  XNOR2X1 U1336 ( .A(n2962), .B(n2991), .Y(n2327) );
  XNOR2X1 U1337 ( .A(n2962), .B(n459), .Y(n2328) );
  XNOR2X1 U1338 ( .A(n2961), .B(n2994), .Y(n2329) );
  XNOR2X1 U1339 ( .A(n2961), .B(n455), .Y(n2330) );
  XNOR2X1 U1340 ( .A(n2961), .B(n2997), .Y(n2331) );
  XNOR2X1 U1341 ( .A(n2936), .B(n451), .Y(n2332) );
  XNOR2X1 U1342 ( .A(n2936), .B(n3000), .Y(n2333) );
  XNOR2X1 U1343 ( .A(n2937), .B(n447), .Y(n2334) );
  XNOR2X1 U1344 ( .A(n323), .B(n3003), .Y(n2335) );
  XNOR2X1 U1345 ( .A(n323), .B(n443), .Y(n2336) );
  XNOR2X1 U1346 ( .A(n325), .B(n3006), .Y(n2337) );
  XNOR2X1 U1347 ( .A(n2937), .B(n439), .Y(n2338) );
  XNOR2X1 U1348 ( .A(n2936), .B(n3009), .Y(n2339) );
  XNOR2X1 U1349 ( .A(n2937), .B(n3012), .Y(n2340) );
  OAI22X1 U1350 ( .A(n370), .B(n2368), .C(n2800), .D(n420), .Y(n1747) );
  OAI22X1 U1351 ( .A(n2342), .B(n370), .C(n2343), .D(n420), .Y(n1852) );
  OAI22X1 U1352 ( .A(n2343), .B(n370), .C(n2344), .D(n420), .Y(n1853) );
  OAI22X1 U1353 ( .A(n2344), .B(n369), .C(n2345), .D(n420), .Y(n1854) );
  OAI22X1 U1354 ( .A(n2345), .B(n369), .C(n2346), .D(n419), .Y(n1855) );
  OAI22X1 U1355 ( .A(n2346), .B(n369), .C(n2347), .D(n419), .Y(n1856) );
  OAI22X1 U1356 ( .A(n2347), .B(n369), .C(n2348), .D(n419), .Y(n1857) );
  OAI22X1 U1357 ( .A(n2348), .B(n369), .C(n2349), .D(n419), .Y(n1858) );
  OAI22X1 U1358 ( .A(n2349), .B(n369), .C(n2350), .D(n419), .Y(n1859) );
  OAI22X1 U1359 ( .A(n2350), .B(n369), .C(n2351), .D(n419), .Y(n1860) );
  OAI22X1 U1360 ( .A(n2351), .B(n369), .C(n2352), .D(n419), .Y(n1861) );
  OAI22X1 U1361 ( .A(n2352), .B(n369), .C(n2353), .D(n419), .Y(n1862) );
  OAI22X1 U1362 ( .A(n2353), .B(n369), .C(n2354), .D(n419), .Y(n1863) );
  OAI22X1 U1363 ( .A(n2354), .B(n369), .C(n2355), .D(n419), .Y(n1864) );
  OAI22X1 U1364 ( .A(n2355), .B(n369), .C(n2356), .D(n419), .Y(n1865) );
  OAI22X1 U1365 ( .A(n2356), .B(n368), .C(n2357), .D(n419), .Y(n1866) );
  OAI22X1 U1366 ( .A(n2357), .B(n368), .C(n2358), .D(n418), .Y(n1867) );
  OAI22X1 U1367 ( .A(n2358), .B(n368), .C(n2359), .D(n418), .Y(n1868) );
  OAI22X1 U1368 ( .A(n2359), .B(n368), .C(n2360), .D(n418), .Y(n1869) );
  OAI22X1 U1369 ( .A(n2360), .B(n368), .C(n2361), .D(n418), .Y(n1870) );
  OAI22X1 U1370 ( .A(n2361), .B(n368), .C(n2362), .D(n418), .Y(n1871) );
  OAI22X1 U1371 ( .A(n2362), .B(n368), .C(n2363), .D(n418), .Y(n1872) );
  OAI22X1 U1372 ( .A(n2363), .B(n368), .C(n2364), .D(n418), .Y(n1873) );
  OAI22X1 U1373 ( .A(n2364), .B(n368), .C(n2365), .D(n418), .Y(n1874) );
  OAI22X1 U1374 ( .A(n2365), .B(n368), .C(n2366), .D(n418), .Y(n1875) );
  OAI22X1 U1375 ( .A(n2366), .B(n368), .C(n2367), .D(n418), .Y(n1876) );
  XNOR2X1 U1376 ( .A(n320), .B(n2975), .Y(n2342) );
  XNOR2X1 U1377 ( .A(n322), .B(n483), .Y(n2343) );
  XNOR2X1 U1378 ( .A(n2939), .B(n2977), .Y(n2344) );
  XNOR2X1 U1379 ( .A(n2938), .B(n479), .Y(n2345) );
  XNOR2X1 U1380 ( .A(n2938), .B(n2980), .Y(n2346) );
  XNOR2X1 U1381 ( .A(n2939), .B(n475), .Y(n2347) );
  XNOR2X1 U1382 ( .A(n320), .B(n2983), .Y(n2348) );
  XNOR2X1 U1383 ( .A(n322), .B(n471), .Y(n2349) );
  XNOR2X1 U1384 ( .A(n322), .B(n2985), .Y(n2350) );
  XNOR2X1 U1385 ( .A(n320), .B(n467), .Y(n2351) );
  XNOR2X1 U1386 ( .A(n2939), .B(n2988), .Y(n2352) );
  XNOR2X1 U1387 ( .A(n320), .B(n463), .Y(n2353) );
  XNOR2X1 U1388 ( .A(n322), .B(n2991), .Y(n2354) );
  XNOR2X1 U1389 ( .A(n2939), .B(n459), .Y(n2355) );
  XNOR2X1 U1390 ( .A(n2938), .B(n2994), .Y(n2356) );
  XNOR2X1 U1391 ( .A(n320), .B(n455), .Y(n2357) );
  XNOR2X1 U1392 ( .A(n2939), .B(n2997), .Y(n2358) );
  XNOR2X1 U1393 ( .A(n2939), .B(n451), .Y(n2359) );
  XNOR2X1 U1394 ( .A(n320), .B(n3000), .Y(n2360) );
  XNOR2X1 U1395 ( .A(n320), .B(n447), .Y(n2361) );
  XNOR2X1 U1396 ( .A(n2938), .B(n3003), .Y(n2362) );
  XNOR2X1 U1397 ( .A(n322), .B(n443), .Y(n2363) );
  XNOR2X1 U1398 ( .A(n2938), .B(n3006), .Y(n2364) );
  XNOR2X1 U1399 ( .A(n320), .B(n439), .Y(n2365) );
  XNOR2X1 U1400 ( .A(n2939), .B(n3009), .Y(n2366) );
  XNOR2X1 U1401 ( .A(n2938), .B(n3012), .Y(n2367) );
  OAI22X1 U1402 ( .A(n367), .B(n2397), .C(n2801), .D(n417), .Y(n1748) );
  OAI22X1 U1403 ( .A(n2369), .B(n367), .C(n2370), .D(n417), .Y(n1878) );
  OAI22X1 U1404 ( .A(n2370), .B(n367), .C(n2371), .D(n417), .Y(n1879) );
  OAI22X1 U1405 ( .A(n2371), .B(n367), .C(n2372), .D(n417), .Y(n1880) );
  OAI22X1 U1406 ( .A(n2372), .B(n367), .C(n2373), .D(n417), .Y(n1881) );
  OAI22X1 U1407 ( .A(n2373), .B(n366), .C(n2374), .D(n417), .Y(n1882) );
  OAI22X1 U1408 ( .A(n2374), .B(n366), .C(n2375), .D(n416), .Y(n1883) );
  OAI22X1 U1409 ( .A(n2375), .B(n366), .C(n2376), .D(n416), .Y(n1884) );
  OAI22X1 U1410 ( .A(n2376), .B(n366), .C(n2377), .D(n416), .Y(n1885) );
  OAI22X1 U1411 ( .A(n2377), .B(n366), .C(n2378), .D(n416), .Y(n1886) );
  OAI22X1 U1412 ( .A(n2378), .B(n366), .C(n2379), .D(n416), .Y(n1887) );
  OAI22X1 U1413 ( .A(n2379), .B(n366), .C(n2380), .D(n416), .Y(n1888) );
  OAI22X1 U1414 ( .A(n2380), .B(n366), .C(n2381), .D(n416), .Y(n1889) );
  OAI22X1 U1415 ( .A(n2381), .B(n366), .C(n2382), .D(n416), .Y(n1890) );
  OAI22X1 U1416 ( .A(n2382), .B(n366), .C(n2383), .D(n416), .Y(n1891) );
  OAI22X1 U1417 ( .A(n2383), .B(n366), .C(n2384), .D(n416), .Y(n1892) );
  OAI22X1 U1418 ( .A(n2384), .B(n366), .C(n2385), .D(n416), .Y(n1893) );
  OAI22X1 U1419 ( .A(n2385), .B(n365), .C(n2386), .D(n416), .Y(n1894) );
  OAI22X1 U1420 ( .A(n2386), .B(n365), .C(n2387), .D(n415), .Y(n1895) );
  OAI22X1 U1421 ( .A(n2387), .B(n365), .C(n2388), .D(n415), .Y(n1896) );
  OAI22X1 U1422 ( .A(n2388), .B(n365), .C(n2389), .D(n415), .Y(n1897) );
  OAI22X1 U1423 ( .A(n2389), .B(n365), .C(n2390), .D(n415), .Y(n1898) );
  OAI22X1 U1424 ( .A(n2390), .B(n365), .C(n2391), .D(n415), .Y(n1899) );
  OAI22X1 U1425 ( .A(n2391), .B(n365), .C(n2392), .D(n415), .Y(n1900) );
  OAI22X1 U1426 ( .A(n2392), .B(n365), .C(n2393), .D(n415), .Y(n1901) );
  OAI22X1 U1427 ( .A(n2393), .B(n365), .C(n2394), .D(n415), .Y(n1902) );
  OAI22X1 U1428 ( .A(n2394), .B(n365), .C(n2395), .D(n415), .Y(n1903) );
  OAI22X1 U1429 ( .A(n2395), .B(n365), .C(n2396), .D(n415), .Y(n1904) );
  XNOR2X1 U1430 ( .A(n319), .B(n2973), .Y(n2369) );
  XNOR2X1 U1431 ( .A(n319), .B(b[26]), .Y(n2370) );
  XNOR2X1 U1432 ( .A(n319), .B(n2975), .Y(n2371) );
  XNOR2X1 U1433 ( .A(n319), .B(n483), .Y(n2372) );
  XNOR2X1 U1434 ( .A(n319), .B(n2977), .Y(n2373) );
  XNOR2X1 U1435 ( .A(n319), .B(n479), .Y(n2374) );
  XNOR2X1 U1436 ( .A(n319), .B(n2980), .Y(n2375) );
  XNOR2X1 U1437 ( .A(n2916), .B(n475), .Y(n2376) );
  XNOR2X1 U1438 ( .A(n2916), .B(n2983), .Y(n2377) );
  XNOR2X1 U1439 ( .A(n2917), .B(n471), .Y(n2378) );
  XNOR2X1 U1440 ( .A(n2917), .B(n2985), .Y(n2379) );
  XNOR2X1 U1441 ( .A(n2917), .B(n467), .Y(n2380) );
  XNOR2X1 U1442 ( .A(n2916), .B(n2988), .Y(n2381) );
  XNOR2X1 U1443 ( .A(n2917), .B(n463), .Y(n2382) );
  XNOR2X1 U1444 ( .A(n2915), .B(n2991), .Y(n2383) );
  XNOR2X1 U1445 ( .A(n2916), .B(n459), .Y(n2384) );
  XNOR2X1 U1446 ( .A(n2916), .B(n2994), .Y(n2385) );
  XNOR2X1 U1447 ( .A(n2915), .B(n455), .Y(n2386) );
  XNOR2X1 U1448 ( .A(n2915), .B(n2997), .Y(n2387) );
  XNOR2X1 U1449 ( .A(n317), .B(n451), .Y(n2388) );
  XNOR2X1 U1450 ( .A(n317), .B(n3000), .Y(n2389) );
  XNOR2X1 U1451 ( .A(n317), .B(n447), .Y(n2390) );
  XNOR2X1 U1452 ( .A(n317), .B(n3003), .Y(n2391) );
  XNOR2X1 U1453 ( .A(n317), .B(n443), .Y(n2392) );
  XNOR2X1 U1454 ( .A(n317), .B(n3006), .Y(n2393) );
  XNOR2X1 U1455 ( .A(n317), .B(n439), .Y(n2394) );
  XNOR2X1 U1456 ( .A(n317), .B(n3009), .Y(n2395) );
  XNOR2X1 U1457 ( .A(n317), .B(n3011), .Y(n2396) );
  OAI22X1 U1458 ( .A(n364), .B(n2428), .C(n2802), .D(n414), .Y(n1749) );
  OAI22X1 U1459 ( .A(n2398), .B(n364), .C(n2399), .D(n414), .Y(n1906) );
  OAI22X1 U1460 ( .A(n2399), .B(n364), .C(n2400), .D(n414), .Y(n1907) );
  OAI22X1 U1461 ( .A(n2400), .B(n364), .C(n2401), .D(n414), .Y(n1908) );
  OAI22X1 U1462 ( .A(n2401), .B(n364), .C(n2402), .D(n414), .Y(n1909) );
  OAI22X1 U1463 ( .A(n2402), .B(n364), .C(n2403), .D(n414), .Y(n1910) );
  OAI22X1 U1464 ( .A(n2403), .B(n364), .C(n2404), .D(n414), .Y(n1911) );
  OAI22X1 U1465 ( .A(n2404), .B(n363), .C(n2405), .D(n414), .Y(n1912) );
  OAI22X1 U1466 ( .A(n2405), .B(n363), .C(n2406), .D(n413), .Y(n1913) );
  OAI22X1 U1467 ( .A(n2406), .B(n363), .C(n2407), .D(n413), .Y(n1914) );
  OAI22X1 U1468 ( .A(n2407), .B(n363), .C(n2408), .D(n413), .Y(n1915) );
  OAI22X1 U1469 ( .A(n2408), .B(n363), .C(n2409), .D(n413), .Y(n1916) );
  OAI22X1 U1470 ( .A(n2409), .B(n363), .C(n2410), .D(n413), .Y(n1917) );
  OAI22X1 U1471 ( .A(n2410), .B(n363), .C(n2411), .D(n413), .Y(n1918) );
  OAI22X1 U1472 ( .A(n2411), .B(n363), .C(n2412), .D(n413), .Y(n1919) );
  OAI22X1 U1473 ( .A(n2412), .B(n363), .C(n2413), .D(n413), .Y(n1920) );
  OAI22X1 U1474 ( .A(n2413), .B(n363), .C(n2414), .D(n413), .Y(n1921) );
  OAI22X1 U1475 ( .A(n2414), .B(n363), .C(n2415), .D(n413), .Y(n1922) );
  OAI22X1 U1476 ( .A(n2415), .B(n363), .C(n2416), .D(n413), .Y(n1923) );
  OAI22X1 U1477 ( .A(n2416), .B(n362), .C(n2417), .D(n413), .Y(n1924) );
  OAI22X1 U1478 ( .A(n2417), .B(n362), .C(n2418), .D(n412), .Y(n1925) );
  OAI22X1 U1479 ( .A(n2418), .B(n362), .C(n2419), .D(n412), .Y(n1926) );
  OAI22X1 U1480 ( .A(n2419), .B(n362), .C(n2420), .D(n412), .Y(n1927) );
  OAI22X1 U1481 ( .A(n2420), .B(n362), .C(n2421), .D(n412), .Y(n1928) );
  OAI22X1 U1482 ( .A(n2421), .B(n362), .C(n2422), .D(n412), .Y(n1929) );
  OAI22X1 U1483 ( .A(n2422), .B(n362), .C(n2423), .D(n412), .Y(n1930) );
  OAI22X1 U1484 ( .A(n2423), .B(n362), .C(n2424), .D(n412), .Y(n1931) );
  OAI22X1 U1485 ( .A(n2424), .B(n362), .C(n2425), .D(n412), .Y(n1932) );
  OAI22X1 U1486 ( .A(n2425), .B(n362), .C(n2426), .D(n412), .Y(n1933) );
  OAI22X1 U1487 ( .A(n2426), .B(n362), .C(n2427), .D(n412), .Y(n1934) );
  XNOR2X1 U1488 ( .A(n316), .B(n2971), .Y(n2398) );
  XNOR2X1 U1489 ( .A(n316), .B(b[28]), .Y(n2399) );
  XNOR2X1 U1490 ( .A(n316), .B(n2973), .Y(n2400) );
  XNOR2X1 U1491 ( .A(n316), .B(b[26]), .Y(n2401) );
  XNOR2X1 U1492 ( .A(n316), .B(n2975), .Y(n2402) );
  XNOR2X1 U1493 ( .A(n316), .B(n483), .Y(n2403) );
  XNOR2X1 U1494 ( .A(n316), .B(n2977), .Y(n2404) );
  XNOR2X1 U1495 ( .A(n316), .B(n479), .Y(n2405) );
  XNOR2X1 U1496 ( .A(n316), .B(n2980), .Y(n2406) );
  XNOR2X1 U1497 ( .A(n315), .B(n475), .Y(n2407) );
  XNOR2X1 U1498 ( .A(n315), .B(n2983), .Y(n2408) );
  XNOR2X1 U1499 ( .A(n315), .B(n471), .Y(n2409) );
  XNOR2X1 U1500 ( .A(n315), .B(n2985), .Y(n2410) );
  XNOR2X1 U1501 ( .A(n315), .B(n467), .Y(n2411) );
  XNOR2X1 U1502 ( .A(n315), .B(n2988), .Y(n2412) );
  XNOR2X1 U1503 ( .A(n315), .B(n463), .Y(n2413) );
  XNOR2X1 U1504 ( .A(n315), .B(n2991), .Y(n2414) );
  XNOR2X1 U1505 ( .A(n315), .B(n459), .Y(n2415) );
  XNOR2X1 U1506 ( .A(n315), .B(n2994), .Y(n2416) );
  XNOR2X1 U1507 ( .A(n315), .B(n455), .Y(n2417) );
  XNOR2X1 U1508 ( .A(n315), .B(n2997), .Y(n2418) );
  XNOR2X1 U1509 ( .A(n314), .B(n451), .Y(n2419) );
  XNOR2X1 U1510 ( .A(n314), .B(n3000), .Y(n2420) );
  XNOR2X1 U1511 ( .A(n314), .B(n447), .Y(n2421) );
  XNOR2X1 U1512 ( .A(n314), .B(n3003), .Y(n2422) );
  XNOR2X1 U1513 ( .A(n314), .B(n443), .Y(n2423) );
  XNOR2X1 U1514 ( .A(n314), .B(n3006), .Y(n2424) );
  XNOR2X1 U1515 ( .A(n314), .B(n439), .Y(n2425) );
  XNOR2X1 U1516 ( .A(n314), .B(n3009), .Y(n2426) );
  XNOR2X1 U1517 ( .A(n314), .B(n3011), .Y(n2427) );
  OAI22X1 U1518 ( .A(n361), .B(n2461), .C(n2803), .D(n411), .Y(n1750) );
  OAI22X1 U1519 ( .A(n2429), .B(n361), .C(n2430), .D(n410), .Y(n1936) );
  OAI22X1 U1520 ( .A(n2430), .B(n361), .C(n2431), .D(n410), .Y(n1937) );
  OAI22X1 U1521 ( .A(n2431), .B(n361), .C(n2432), .D(n410), .Y(n1938) );
  OAI22X1 U1522 ( .A(n2432), .B(n361), .C(n2433), .D(n409), .Y(n1939) );
  OAI22X1 U1523 ( .A(n2433), .B(n361), .C(n2434), .D(n410), .Y(n1940) );
  OAI22X1 U1524 ( .A(n2434), .B(n361), .C(n2435), .D(n409), .Y(n1941) );
  OAI22X1 U1525 ( .A(n2435), .B(n361), .C(n2436), .D(n409), .Y(n1942) );
  OAI22X1 U1526 ( .A(n2436), .B(n361), .C(n2437), .D(n410), .Y(n1943) );
  OAI22X1 U1527 ( .A(n2437), .B(n360), .C(n2438), .D(n410), .Y(n1944) );
  OAI22X1 U1528 ( .A(n2438), .B(n360), .C(n2439), .D(n410), .Y(n1945) );
  OAI22X1 U1529 ( .A(n2439), .B(n360), .C(n2440), .D(n409), .Y(n1946) );
  OAI22X1 U1530 ( .A(n2440), .B(n360), .C(n2441), .D(n409), .Y(n1947) );
  OAI22X1 U1531 ( .A(n2441), .B(n360), .C(n2442), .D(n409), .Y(n1948) );
  OAI22X1 U1532 ( .A(n2442), .B(n360), .C(n2443), .D(n410), .Y(n1949) );
  OAI22X1 U1533 ( .A(n2443), .B(n360), .C(n2444), .D(n409), .Y(n1950) );
  OAI22X1 U1534 ( .A(n2444), .B(n360), .C(n2445), .D(n410), .Y(n1951) );
  OAI22X1 U1535 ( .A(n2445), .B(n360), .C(n2446), .D(n410), .Y(n1952) );
  OAI22X1 U1536 ( .A(n2446), .B(n360), .C(n2447), .D(n411), .Y(n1953) );
  OAI22X1 U1537 ( .A(n2447), .B(n360), .C(n2448), .D(n411), .Y(n1954) );
  OAI22X1 U1538 ( .A(n2448), .B(n360), .C(n2449), .D(n410), .Y(n1955) );
  OAI22X1 U1539 ( .A(n2449), .B(n359), .C(n2450), .D(n410), .Y(n1956) );
  OAI22X1 U1540 ( .A(n2450), .B(n359), .C(n2451), .D(n409), .Y(n1957) );
  OAI22X1 U1541 ( .A(n2451), .B(n359), .C(n2452), .D(n409), .Y(n1958) );
  OAI22X1 U1542 ( .A(n2452), .B(n359), .C(n2453), .D(n410), .Y(n1959) );
  OAI22X1 U1543 ( .A(n2453), .B(n359), .C(n2454), .D(n409), .Y(n1960) );
  OAI22X1 U1544 ( .A(n2454), .B(n359), .C(n2455), .D(n410), .Y(n1961) );
  OAI22X1 U1545 ( .A(n2455), .B(n359), .C(n2456), .D(n410), .Y(n1962) );
  OAI22X1 U1546 ( .A(n2456), .B(n359), .C(n2457), .D(n409), .Y(n1963) );
  OAI22X1 U1547 ( .A(n2457), .B(n359), .C(n2458), .D(n409), .Y(n1964) );
  OAI22X1 U1548 ( .A(n2458), .B(n359), .C(n2459), .D(n411), .Y(n1965) );
  OAI22X1 U1549 ( .A(n2459), .B(n359), .C(n2460), .D(n411), .Y(n1966) );
  XNOR2X1 U1550 ( .A(n313), .B(n2969), .Y(n2429) );
  XNOR2X1 U1551 ( .A(n313), .B(b[30]), .Y(n2430) );
  XNOR2X1 U1552 ( .A(n313), .B(n2971), .Y(n2431) );
  XNOR2X1 U1553 ( .A(n313), .B(b[28]), .Y(n2432) );
  XNOR2X1 U1554 ( .A(n313), .B(n2973), .Y(n2433) );
  XNOR2X1 U1555 ( .A(n313), .B(b[26]), .Y(n2434) );
  XNOR2X1 U1556 ( .A(n313), .B(n2975), .Y(n2435) );
  XNOR2X1 U1557 ( .A(n313), .B(n483), .Y(n2436) );
  XNOR2X1 U1558 ( .A(n313), .B(n2977), .Y(n2437) );
  XNOR2X1 U1559 ( .A(n313), .B(n479), .Y(n2438) );
  XNOR2X1 U1560 ( .A(n313), .B(n2980), .Y(n2439) );
  XNOR2X1 U1561 ( .A(n312), .B(n475), .Y(n2440) );
  XNOR2X1 U1562 ( .A(n312), .B(n2983), .Y(n2441) );
  XNOR2X1 U1563 ( .A(n312), .B(n471), .Y(n2442) );
  XNOR2X1 U1564 ( .A(n312), .B(n2985), .Y(n2443) );
  XNOR2X1 U1565 ( .A(n312), .B(n467), .Y(n2444) );
  XNOR2X1 U1566 ( .A(n312), .B(n2988), .Y(n2445) );
  XNOR2X1 U1567 ( .A(n312), .B(n463), .Y(n2446) );
  XNOR2X1 U1568 ( .A(n312), .B(n2991), .Y(n2447) );
  XNOR2X1 U1569 ( .A(n312), .B(n459), .Y(n2448) );
  XNOR2X1 U1570 ( .A(n312), .B(n2994), .Y(n2449) );
  XNOR2X1 U1571 ( .A(n312), .B(n455), .Y(n2450) );
  XNOR2X1 U1572 ( .A(n312), .B(n2997), .Y(n2451) );
  XNOR2X1 U1573 ( .A(n311), .B(n451), .Y(n2452) );
  XNOR2X1 U1574 ( .A(n311), .B(n3000), .Y(n2453) );
  XNOR2X1 U1575 ( .A(n311), .B(n447), .Y(n2454) );
  XNOR2X1 U1576 ( .A(n311), .B(n3003), .Y(n2455) );
  XNOR2X1 U1577 ( .A(n311), .B(n443), .Y(n2456) );
  XNOR2X1 U1578 ( .A(n311), .B(n3006), .Y(n2457) );
  XNOR2X1 U1579 ( .A(n311), .B(n439), .Y(n2458) );
  XNOR2X1 U1580 ( .A(n311), .B(n3009), .Y(n2459) );
  XNOR2X1 U1581 ( .A(n311), .B(n3011), .Y(n2460) );
  OAI22X1 U1582 ( .A(n358), .B(n2494), .C(n2804), .D(n408), .Y(n1751) );
  OAI22X1 U1583 ( .A(n2804), .B(n358), .C(n2462), .D(n408), .Y(n1969) );
  OAI22X1 U1584 ( .A(n2462), .B(n358), .C(n2463), .D(n408), .Y(n1970) );
  OAI22X1 U1585 ( .A(n2463), .B(n358), .C(n2464), .D(n408), .Y(n1971) );
  OAI22X1 U1586 ( .A(n2464), .B(n358), .C(n2465), .D(n408), .Y(n1972) );
  OAI22X1 U1587 ( .A(n2465), .B(n358), .C(n2466), .D(n408), .Y(n1973) );
  OAI22X1 U1588 ( .A(n2466), .B(n358), .C(n2467), .D(n408), .Y(n1974) );
  OAI22X1 U1589 ( .A(n2467), .B(n358), .C(n2468), .D(n408), .Y(n1975) );
  OAI22X1 U1590 ( .A(n2468), .B(n358), .C(n2469), .D(n408), .Y(n1976) );
  OAI22X1 U1591 ( .A(n2469), .B(n358), .C(n2470), .D(n408), .Y(n1977) );
  OAI22X1 U1592 ( .A(n2470), .B(n357), .C(n2471), .D(n408), .Y(n1978) );
  OAI22X1 U1593 ( .A(n2471), .B(n357), .C(n2472), .D(n407), .Y(n1979) );
  OAI22X1 U1594 ( .A(n2472), .B(n357), .C(n2473), .D(n407), .Y(n1980) );
  OAI22X1 U1595 ( .A(n2473), .B(n357), .C(n2474), .D(n407), .Y(n1981) );
  OAI22X1 U1596 ( .A(n2474), .B(n357), .C(n2475), .D(n407), .Y(n1982) );
  OAI22X1 U1597 ( .A(n2475), .B(n357), .C(n2476), .D(n407), .Y(n1983) );
  OAI22X1 U1598 ( .A(n2476), .B(n357), .C(n2477), .D(n407), .Y(n1984) );
  OAI22X1 U1599 ( .A(n2477), .B(n357), .C(n2478), .D(n407), .Y(n1985) );
  OAI22X1 U1600 ( .A(n2478), .B(n357), .C(n2479), .D(n407), .Y(n1986) );
  OAI22X1 U1601 ( .A(n2479), .B(n357), .C(n2480), .D(n407), .Y(n1987) );
  OAI22X1 U1602 ( .A(n2480), .B(n357), .C(n2481), .D(n407), .Y(n1988) );
  OAI22X1 U1603 ( .A(n2481), .B(n357), .C(n2482), .D(n407), .Y(n1989) );
  OAI22X1 U1604 ( .A(n2482), .B(n356), .C(n2483), .D(n407), .Y(n1990) );
  OAI22X1 U1605 ( .A(n2483), .B(n356), .C(n2484), .D(n406), .Y(n1991) );
  OAI22X1 U1606 ( .A(n2484), .B(n356), .C(n2485), .D(n406), .Y(n1992) );
  OAI22X1 U1607 ( .A(n2485), .B(n356), .C(n2486), .D(n406), .Y(n1993) );
  OAI22X1 U1608 ( .A(n2486), .B(n356), .C(n2487), .D(n406), .Y(n1994) );
  OAI22X1 U1609 ( .A(n2487), .B(n356), .C(n2488), .D(n406), .Y(n1995) );
  OAI22X1 U1610 ( .A(n2488), .B(n356), .C(n2489), .D(n406), .Y(n1996) );
  OAI22X1 U1611 ( .A(n2489), .B(n356), .C(n2490), .D(n406), .Y(n1997) );
  OAI22X1 U1612 ( .A(n2490), .B(n356), .C(n2491), .D(n406), .Y(n1998) );
  OAI22X1 U1613 ( .A(n2491), .B(n356), .C(n2492), .D(n406), .Y(n1999) );
  OAI22X1 U1614 ( .A(n2492), .B(n356), .C(n2493), .D(n406), .Y(n2000) );
  XNOR2X1 U1615 ( .A(n310), .B(n2969), .Y(n2462) );
  XNOR2X1 U1616 ( .A(n310), .B(n495), .Y(n2463) );
  XNOR2X1 U1617 ( .A(n310), .B(n2971), .Y(n2464) );
  XNOR2X1 U1618 ( .A(n310), .B(n491), .Y(n2465) );
  XNOR2X1 U1619 ( .A(n310), .B(n2973), .Y(n2466) );
  XNOR2X1 U1620 ( .A(n310), .B(n487), .Y(n2467) );
  XNOR2X1 U1621 ( .A(n310), .B(n2975), .Y(n2468) );
  XNOR2X1 U1622 ( .A(n310), .B(n483), .Y(n2469) );
  XNOR2X1 U1623 ( .A(n310), .B(n2977), .Y(n2470) );
  XNOR2X1 U1624 ( .A(n310), .B(n479), .Y(n2471) );
  XNOR2X1 U1625 ( .A(n310), .B(n2980), .Y(n2472) );
  XNOR2X1 U1626 ( .A(n309), .B(n475), .Y(n2473) );
  XNOR2X1 U1627 ( .A(n309), .B(n2983), .Y(n2474) );
  XNOR2X1 U1628 ( .A(n309), .B(n471), .Y(n2475) );
  XNOR2X1 U1629 ( .A(n309), .B(n2985), .Y(n2476) );
  XNOR2X1 U1630 ( .A(n309), .B(n467), .Y(n2477) );
  XNOR2X1 U1631 ( .A(n309), .B(n2989), .Y(n2478) );
  XNOR2X1 U1632 ( .A(n309), .B(n463), .Y(n2479) );
  XNOR2X1 U1633 ( .A(n309), .B(n2992), .Y(n2480) );
  XNOR2X1 U1634 ( .A(n309), .B(n459), .Y(n2481) );
  XNOR2X1 U1635 ( .A(n309), .B(n2995), .Y(n2482) );
  XNOR2X1 U1636 ( .A(n309), .B(n455), .Y(n2483) );
  XNOR2X1 U1637 ( .A(n309), .B(n2998), .Y(n2484) );
  XNOR2X1 U1638 ( .A(n308), .B(n451), .Y(n2485) );
  XNOR2X1 U1639 ( .A(n308), .B(n3001), .Y(n2486) );
  XNOR2X1 U1640 ( .A(n308), .B(n447), .Y(n2487) );
  XNOR2X1 U1641 ( .A(n308), .B(n3004), .Y(n2488) );
  XNOR2X1 U1642 ( .A(n308), .B(n443), .Y(n2489) );
  XNOR2X1 U1643 ( .A(n308), .B(n3007), .Y(n2490) );
  XNOR2X1 U1644 ( .A(n308), .B(n439), .Y(n2491) );
  XNOR2X1 U1645 ( .A(n308), .B(b[1]), .Y(n2492) );
  XNOR2X1 U1646 ( .A(n308), .B(n3011), .Y(n2493) );
  OAI22X1 U1647 ( .A(n355), .B(n2527), .C(n2805), .D(n405), .Y(n1752) );
  OAI22X1 U1648 ( .A(n2805), .B(n355), .C(n2495), .D(n404), .Y(n2003) );
  OAI22X1 U1649 ( .A(n2495), .B(n355), .C(n2496), .D(n404), .Y(n2004) );
  OAI22X1 U1650 ( .A(n2496), .B(n355), .C(n2497), .D(n404), .Y(n2005) );
  OAI22X1 U1651 ( .A(n2497), .B(n355), .C(n2498), .D(n405), .Y(n2006) );
  OAI22X1 U1652 ( .A(n2498), .B(n355), .C(n2499), .D(n405), .Y(n2007) );
  OAI22X1 U1653 ( .A(n2499), .B(n355), .C(n2500), .D(n404), .Y(n2008) );
  OAI22X1 U1654 ( .A(n2500), .B(n355), .C(n2501), .D(n405), .Y(n2009) );
  OAI22X1 U1655 ( .A(n2501), .B(n355), .C(n2502), .D(n405), .Y(n2010) );
  OAI22X1 U1656 ( .A(n2502), .B(n355), .C(n2503), .D(n404), .Y(n2011) );
  OAI22X1 U1657 ( .A(n2503), .B(n354), .C(n2504), .D(n405), .Y(n2012) );
  OAI22X1 U1658 ( .A(n2504), .B(n354), .C(n2505), .D(n404), .Y(n2013) );
  OAI22X1 U1659 ( .A(n2505), .B(n354), .C(n2506), .D(n405), .Y(n2014) );
  OAI22X1 U1660 ( .A(n2506), .B(n354), .C(n2507), .D(n404), .Y(n2015) );
  OAI22X1 U1661 ( .A(n2507), .B(n354), .C(n2508), .D(n403), .Y(n2016) );
  OAI22X1 U1662 ( .A(n2508), .B(n354), .C(n2509), .D(n403), .Y(n2017) );
  OAI22X1 U1663 ( .A(n2509), .B(n354), .C(n2510), .D(n405), .Y(n2018) );
  OAI22X1 U1664 ( .A(n2510), .B(n354), .C(n2511), .D(n404), .Y(n2019) );
  OAI22X1 U1665 ( .A(n2511), .B(n354), .C(n2512), .D(n405), .Y(n2020) );
  OAI22X1 U1666 ( .A(n2512), .B(n354), .C(n2513), .D(n403), .Y(n2021) );
  OAI22X1 U1667 ( .A(n2513), .B(n354), .C(n2514), .D(n403), .Y(n2022) );
  OAI22X1 U1668 ( .A(n2514), .B(n354), .C(n2515), .D(n403), .Y(n2023) );
  OAI22X1 U1669 ( .A(n2515), .B(n353), .C(n2516), .D(n403), .Y(n2024) );
  OAI22X1 U1670 ( .A(n2516), .B(n353), .C(n2517), .D(n404), .Y(n2025) );
  OAI22X1 U1671 ( .A(n2517), .B(n353), .C(n2518), .D(n403), .Y(n2026) );
  OAI22X1 U1672 ( .A(n2518), .B(n353), .C(n2519), .D(n404), .Y(n2027) );
  OAI22X1 U1673 ( .A(n2519), .B(n353), .C(n2520), .D(n405), .Y(n2028) );
  OAI22X1 U1674 ( .A(n2520), .B(n353), .C(n2521), .D(n405), .Y(n2029) );
  OAI22X1 U1675 ( .A(n2521), .B(n353), .C(n2522), .D(n405), .Y(n2030) );
  OAI22X1 U1676 ( .A(n2522), .B(n353), .C(n2523), .D(n404), .Y(n2031) );
  OAI22X1 U1677 ( .A(n2523), .B(n353), .C(n2524), .D(n404), .Y(n2032) );
  OAI22X1 U1678 ( .A(n2524), .B(n353), .C(n2525), .D(n403), .Y(n2033) );
  OAI22X1 U1679 ( .A(n2525), .B(n353), .C(n2526), .D(n404), .Y(n2034) );
  XNOR2X1 U1680 ( .A(n307), .B(n2969), .Y(n2495) );
  XNOR2X1 U1681 ( .A(n307), .B(n495), .Y(n2496) );
  XNOR2X1 U1682 ( .A(n307), .B(n2971), .Y(n2497) );
  XNOR2X1 U1683 ( .A(n307), .B(n491), .Y(n2498) );
  XNOR2X1 U1684 ( .A(n307), .B(n2973), .Y(n2499) );
  XNOR2X1 U1685 ( .A(n307), .B(n487), .Y(n2500) );
  XNOR2X1 U1686 ( .A(n307), .B(n2975), .Y(n2501) );
  XNOR2X1 U1687 ( .A(n307), .B(n483), .Y(n2502) );
  XNOR2X1 U1688 ( .A(n307), .B(n2977), .Y(n2503) );
  XNOR2X1 U1689 ( .A(n307), .B(n479), .Y(n2504) );
  XNOR2X1 U1690 ( .A(n307), .B(n2980), .Y(n2505) );
  XNOR2X1 U1691 ( .A(n306), .B(n475), .Y(n2506) );
  XNOR2X1 U1692 ( .A(n306), .B(n2983), .Y(n2507) );
  XNOR2X1 U1693 ( .A(n306), .B(n471), .Y(n2508) );
  XNOR2X1 U1694 ( .A(n306), .B(n2985), .Y(n2509) );
  XNOR2X1 U1695 ( .A(n306), .B(n467), .Y(n2510) );
  XNOR2X1 U1696 ( .A(n306), .B(n2989), .Y(n2511) );
  XNOR2X1 U1697 ( .A(n306), .B(n463), .Y(n2512) );
  XNOR2X1 U1698 ( .A(n306), .B(n2992), .Y(n2513) );
  XNOR2X1 U1699 ( .A(n306), .B(n459), .Y(n2514) );
  XNOR2X1 U1700 ( .A(n306), .B(n2995), .Y(n2515) );
  XNOR2X1 U1701 ( .A(n306), .B(n455), .Y(n2516) );
  XNOR2X1 U1702 ( .A(n306), .B(n2998), .Y(n2517) );
  XNOR2X1 U1703 ( .A(n305), .B(n451), .Y(n2518) );
  XNOR2X1 U1704 ( .A(n305), .B(n3001), .Y(n2519) );
  XNOR2X1 U1705 ( .A(n305), .B(n447), .Y(n2520) );
  XNOR2X1 U1706 ( .A(n305), .B(n3004), .Y(n2521) );
  XNOR2X1 U1707 ( .A(n305), .B(n443), .Y(n2522) );
  XNOR2X1 U1708 ( .A(n305), .B(n3007), .Y(n2523) );
  XNOR2X1 U1709 ( .A(n305), .B(n439), .Y(n2524) );
  XNOR2X1 U1710 ( .A(n305), .B(b[1]), .Y(n2525) );
  XNOR2X1 U1711 ( .A(n305), .B(n3011), .Y(n2526) );
  OAI22X1 U1712 ( .A(n352), .B(n2560), .C(n2806), .D(n402), .Y(n1753) );
  OAI22X1 U1713 ( .A(n2806), .B(n352), .C(n2528), .D(n402), .Y(n2037) );
  OAI22X1 U1714 ( .A(n2528), .B(n352), .C(n2529), .D(n402), .Y(n2038) );
  OAI22X1 U1715 ( .A(n2529), .B(n352), .C(n2530), .D(n402), .Y(n2039) );
  OAI22X1 U1716 ( .A(n2530), .B(n352), .C(n2531), .D(n402), .Y(n2040) );
  OAI22X1 U1717 ( .A(n2531), .B(n352), .C(n2532), .D(n402), .Y(n2041) );
  OAI22X1 U1718 ( .A(n2532), .B(n352), .C(n2533), .D(n402), .Y(n2042) );
  OAI22X1 U1719 ( .A(n2533), .B(n352), .C(n2534), .D(n402), .Y(n2043) );
  OAI22X1 U1720 ( .A(n2534), .B(n352), .C(n2535), .D(n402), .Y(n2044) );
  OAI22X1 U1721 ( .A(n2535), .B(n352), .C(n2536), .D(n402), .Y(n2045) );
  OAI22X1 U1722 ( .A(n2536), .B(n351), .C(n2537), .D(n402), .Y(n2046) );
  OAI22X1 U1723 ( .A(n2537), .B(n351), .C(n2538), .D(n401), .Y(n2047) );
  OAI22X1 U1724 ( .A(n2538), .B(n351), .C(n2539), .D(n401), .Y(n2048) );
  OAI22X1 U1725 ( .A(n2539), .B(n351), .C(n2540), .D(n401), .Y(n2049) );
  OAI22X1 U1726 ( .A(n2540), .B(n351), .C(n2541), .D(n401), .Y(n2050) );
  OAI22X1 U1727 ( .A(n2541), .B(n351), .C(n2542), .D(n401), .Y(n2051) );
  OAI22X1 U1728 ( .A(n2542), .B(n351), .C(n2543), .D(n401), .Y(n2052) );
  OAI22X1 U1729 ( .A(n2543), .B(n351), .C(n2544), .D(n401), .Y(n2053) );
  OAI22X1 U1730 ( .A(n2544), .B(n351), .C(n2545), .D(n401), .Y(n2054) );
  OAI22X1 U1731 ( .A(n2545), .B(n351), .C(n2546), .D(n401), .Y(n2055) );
  OAI22X1 U1732 ( .A(n2546), .B(n351), .C(n2547), .D(n401), .Y(n2056) );
  OAI22X1 U1733 ( .A(n2547), .B(n351), .C(n2548), .D(n401), .Y(n2057) );
  OAI22X1 U1734 ( .A(n2548), .B(n350), .C(n2549), .D(n401), .Y(n2058) );
  OAI22X1 U1735 ( .A(n2549), .B(n350), .C(n2550), .D(n400), .Y(n2059) );
  OAI22X1 U1736 ( .A(n2550), .B(n350), .C(n2551), .D(n400), .Y(n2060) );
  OAI22X1 U1737 ( .A(n2551), .B(n350), .C(n2552), .D(n400), .Y(n2061) );
  OAI22X1 U1738 ( .A(n2552), .B(n350), .C(n2553), .D(n400), .Y(n2062) );
  OAI22X1 U1739 ( .A(n2553), .B(n350), .C(n2554), .D(n400), .Y(n2063) );
  OAI22X1 U1740 ( .A(n2554), .B(n350), .C(n2555), .D(n400), .Y(n2064) );
  OAI22X1 U1741 ( .A(n2555), .B(n350), .C(n2556), .D(n400), .Y(n2065) );
  OAI22X1 U1742 ( .A(n2556), .B(n350), .C(n2557), .D(n400), .Y(n2066) );
  OAI22X1 U1743 ( .A(n2557), .B(n350), .C(n2558), .D(n400), .Y(n2067) );
  OAI22X1 U1744 ( .A(n2558), .B(n350), .C(n2559), .D(n400), .Y(n2068) );
  XNOR2X1 U1745 ( .A(n304), .B(n2969), .Y(n2528) );
  XNOR2X1 U1746 ( .A(n304), .B(n495), .Y(n2529) );
  XNOR2X1 U1747 ( .A(n304), .B(n2971), .Y(n2530) );
  XNOR2X1 U1748 ( .A(n304), .B(n491), .Y(n2531) );
  XNOR2X1 U1749 ( .A(n304), .B(n2973), .Y(n2532) );
  XNOR2X1 U1750 ( .A(n304), .B(n487), .Y(n2533) );
  XNOR2X1 U1751 ( .A(n304), .B(n2975), .Y(n2534) );
  XNOR2X1 U1752 ( .A(n304), .B(n483), .Y(n2535) );
  XNOR2X1 U1753 ( .A(n304), .B(n2977), .Y(n2536) );
  XNOR2X1 U1754 ( .A(n304), .B(n479), .Y(n2537) );
  XNOR2X1 U1755 ( .A(n304), .B(n2980), .Y(n2538) );
  XNOR2X1 U1756 ( .A(n303), .B(n475), .Y(n2539) );
  XNOR2X1 U1757 ( .A(n303), .B(n2983), .Y(n2540) );
  XNOR2X1 U1758 ( .A(n303), .B(n471), .Y(n2541) );
  XNOR2X1 U1759 ( .A(n303), .B(n2985), .Y(n2542) );
  XNOR2X1 U1760 ( .A(n303), .B(n467), .Y(n2543) );
  XNOR2X1 U1761 ( .A(n303), .B(n2989), .Y(n2544) );
  XNOR2X1 U1762 ( .A(n303), .B(n463), .Y(n2545) );
  XNOR2X1 U1763 ( .A(n303), .B(n2992), .Y(n2546) );
  XNOR2X1 U1764 ( .A(n303), .B(n459), .Y(n2547) );
  XNOR2X1 U1765 ( .A(n303), .B(n2995), .Y(n2548) );
  XNOR2X1 U1766 ( .A(n303), .B(n455), .Y(n2549) );
  XNOR2X1 U1767 ( .A(n303), .B(n2998), .Y(n2550) );
  XNOR2X1 U1768 ( .A(n302), .B(n451), .Y(n2551) );
  XNOR2X1 U1769 ( .A(n302), .B(n3001), .Y(n2552) );
  XNOR2X1 U1770 ( .A(n302), .B(n447), .Y(n2553) );
  XNOR2X1 U1771 ( .A(n302), .B(n3004), .Y(n2554) );
  XNOR2X1 U1772 ( .A(n302), .B(n443), .Y(n2555) );
  XNOR2X1 U1773 ( .A(n302), .B(n3007), .Y(n2556) );
  XNOR2X1 U1774 ( .A(n302), .B(n439), .Y(n2557) );
  XNOR2X1 U1775 ( .A(n302), .B(b[1]), .Y(n2558) );
  XNOR2X1 U1776 ( .A(n302), .B(n3011), .Y(n2559) );
  OAI22X1 U1777 ( .A(n349), .B(n2593), .C(n2807), .D(n399), .Y(n1754) );
  OAI22X1 U1778 ( .A(n2807), .B(n349), .C(n2561), .D(n399), .Y(n2071) );
  OAI22X1 U1779 ( .A(n2561), .B(n349), .C(n2562), .D(n399), .Y(n2072) );
  OAI22X1 U1780 ( .A(n2562), .B(n349), .C(n2563), .D(n399), .Y(n2073) );
  OAI22X1 U1781 ( .A(n2563), .B(n349), .C(n2564), .D(n399), .Y(n2074) );
  OAI22X1 U1782 ( .A(n2564), .B(n349), .C(n2565), .D(n399), .Y(n2075) );
  OAI22X1 U1783 ( .A(n2565), .B(n349), .C(n2566), .D(n399), .Y(n2076) );
  OAI22X1 U1784 ( .A(n2566), .B(n349), .C(n2567), .D(n399), .Y(n2077) );
  OAI22X1 U1785 ( .A(n2567), .B(n349), .C(n2568), .D(n399), .Y(n2078) );
  OAI22X1 U1786 ( .A(n2568), .B(n349), .C(n2569), .D(n399), .Y(n2079) );
  OAI22X1 U1787 ( .A(n2569), .B(n348), .C(n2570), .D(n399), .Y(n2080) );
  OAI22X1 U1788 ( .A(n2570), .B(n348), .C(n2571), .D(n398), .Y(n2081) );
  OAI22X1 U1789 ( .A(n2571), .B(n348), .C(n2572), .D(n398), .Y(n2082) );
  OAI22X1 U1790 ( .A(n2572), .B(n348), .C(n2573), .D(n398), .Y(n2083) );
  OAI22X1 U1791 ( .A(n2573), .B(n348), .C(n2574), .D(n398), .Y(n2084) );
  OAI22X1 U1792 ( .A(n2574), .B(n348), .C(n2575), .D(n398), .Y(n2085) );
  OAI22X1 U1793 ( .A(n2575), .B(n348), .C(n2576), .D(n398), .Y(n2086) );
  OAI22X1 U1794 ( .A(n2576), .B(n348), .C(n2577), .D(n398), .Y(n2087) );
  OAI22X1 U1795 ( .A(n2577), .B(n348), .C(n2578), .D(n398), .Y(n2088) );
  OAI22X1 U1796 ( .A(n2578), .B(n348), .C(n2579), .D(n398), .Y(n2089) );
  OAI22X1 U1797 ( .A(n2579), .B(n348), .C(n2580), .D(n398), .Y(n2090) );
  OAI22X1 U1798 ( .A(n2580), .B(n348), .C(n2581), .D(n398), .Y(n2091) );
  OAI22X1 U1799 ( .A(n2581), .B(n347), .C(n2582), .D(n398), .Y(n2092) );
  OAI22X1 U1800 ( .A(n2582), .B(n347), .C(n2583), .D(n397), .Y(n2093) );
  OAI22X1 U1801 ( .A(n2583), .B(n347), .C(n2584), .D(n397), .Y(n2094) );
  OAI22X1 U1802 ( .A(n2584), .B(n347), .C(n2585), .D(n397), .Y(n2095) );
  OAI22X1 U1803 ( .A(n2585), .B(n347), .C(n2586), .D(n397), .Y(n2096) );
  OAI22X1 U1804 ( .A(n2586), .B(n347), .C(n2587), .D(n397), .Y(n2097) );
  OAI22X1 U1805 ( .A(n2587), .B(n347), .C(n2588), .D(n397), .Y(n2098) );
  OAI22X1 U1806 ( .A(n2588), .B(n347), .C(n2589), .D(n397), .Y(n2099) );
  OAI22X1 U1807 ( .A(n2589), .B(n347), .C(n2590), .D(n397), .Y(n2100) );
  OAI22X1 U1808 ( .A(n2590), .B(n347), .C(n2591), .D(n397), .Y(n2101) );
  OAI22X1 U1809 ( .A(n2591), .B(n347), .C(n2592), .D(n397), .Y(n2102) );
  XNOR2X1 U1810 ( .A(n301), .B(n2969), .Y(n2561) );
  XNOR2X1 U1811 ( .A(n301), .B(n495), .Y(n2562) );
  XNOR2X1 U1812 ( .A(n301), .B(n2971), .Y(n2563) );
  XNOR2X1 U1813 ( .A(n301), .B(n491), .Y(n2564) );
  XNOR2X1 U1814 ( .A(n301), .B(n2973), .Y(n2565) );
  XNOR2X1 U1815 ( .A(n301), .B(n487), .Y(n2566) );
  XNOR2X1 U1816 ( .A(n301), .B(n2975), .Y(n2567) );
  XNOR2X1 U1817 ( .A(n301), .B(n483), .Y(n2568) );
  XNOR2X1 U1818 ( .A(n301), .B(n2977), .Y(n2569) );
  XNOR2X1 U1819 ( .A(n301), .B(n479), .Y(n2570) );
  XNOR2X1 U1820 ( .A(n301), .B(n2980), .Y(n2571) );
  XNOR2X1 U1821 ( .A(n300), .B(n475), .Y(n2572) );
  XNOR2X1 U1822 ( .A(n300), .B(n2983), .Y(n2573) );
  XNOR2X1 U1823 ( .A(n300), .B(n471), .Y(n2574) );
  XNOR2X1 U1824 ( .A(n300), .B(n2985), .Y(n2575) );
  XNOR2X1 U1825 ( .A(n300), .B(n467), .Y(n2576) );
  XNOR2X1 U1826 ( .A(n300), .B(n2989), .Y(n2577) );
  XNOR2X1 U1827 ( .A(n300), .B(n463), .Y(n2578) );
  XNOR2X1 U1828 ( .A(n300), .B(n2992), .Y(n2579) );
  XNOR2X1 U1829 ( .A(n300), .B(n459), .Y(n2580) );
  XNOR2X1 U1830 ( .A(n300), .B(n2995), .Y(n2581) );
  XNOR2X1 U1831 ( .A(n300), .B(n455), .Y(n2582) );
  XNOR2X1 U1832 ( .A(n300), .B(n2998), .Y(n2583) );
  XNOR2X1 U1833 ( .A(n299), .B(n451), .Y(n2584) );
  XNOR2X1 U1834 ( .A(n299), .B(n3001), .Y(n2585) );
  XNOR2X1 U1835 ( .A(n299), .B(n447), .Y(n2586) );
  XNOR2X1 U1836 ( .A(n299), .B(n3004), .Y(n2587) );
  XNOR2X1 U1837 ( .A(n299), .B(n443), .Y(n2588) );
  XNOR2X1 U1838 ( .A(n299), .B(n3007), .Y(n2589) );
  XNOR2X1 U1839 ( .A(n299), .B(n439), .Y(n2590) );
  XNOR2X1 U1840 ( .A(n299), .B(b[1]), .Y(n2591) );
  XNOR2X1 U1841 ( .A(n299), .B(n3011), .Y(n2592) );
  OAI22X1 U1842 ( .A(n346), .B(n2626), .C(n2808), .D(n396), .Y(n1755) );
  OAI22X1 U1843 ( .A(n2808), .B(n346), .C(n2594), .D(n396), .Y(n2105) );
  OAI22X1 U1844 ( .A(n2594), .B(n346), .C(n2595), .D(n396), .Y(n2106) );
  OAI22X1 U1845 ( .A(n2595), .B(n346), .C(n2596), .D(n396), .Y(n2107) );
  OAI22X1 U1846 ( .A(n2596), .B(n346), .C(n2597), .D(n396), .Y(n2108) );
  OAI22X1 U1847 ( .A(n2597), .B(n346), .C(n2598), .D(n396), .Y(n2109) );
  OAI22X1 U1848 ( .A(n2598), .B(n346), .C(n2599), .D(n396), .Y(n2110) );
  OAI22X1 U1849 ( .A(n2599), .B(n346), .C(n2600), .D(n396), .Y(n2111) );
  OAI22X1 U1850 ( .A(n2600), .B(n346), .C(n2601), .D(n396), .Y(n2112) );
  OAI22X1 U1851 ( .A(n2601), .B(n346), .C(n2602), .D(n396), .Y(n2113) );
  OAI22X1 U1852 ( .A(n2602), .B(n345), .C(n2603), .D(n396), .Y(n2114) );
  OAI22X1 U1853 ( .A(n2603), .B(n345), .C(n2604), .D(n395), .Y(n2115) );
  OAI22X1 U1854 ( .A(n2604), .B(n345), .C(n2605), .D(n395), .Y(n2116) );
  OAI22X1 U1855 ( .A(n2605), .B(n345), .C(n2606), .D(n395), .Y(n2117) );
  OAI22X1 U1856 ( .A(n2606), .B(n345), .C(n2607), .D(n395), .Y(n2118) );
  OAI22X1 U1857 ( .A(n2607), .B(n345), .C(n2608), .D(n395), .Y(n2119) );
  OAI22X1 U1858 ( .A(n2608), .B(n345), .C(n2609), .D(n395), .Y(n2120) );
  OAI22X1 U1859 ( .A(n2609), .B(n345), .C(n2610), .D(n395), .Y(n2121) );
  OAI22X1 U1860 ( .A(n2610), .B(n345), .C(n2611), .D(n395), .Y(n2122) );
  OAI22X1 U1861 ( .A(n2611), .B(n345), .C(n2612), .D(n395), .Y(n2123) );
  OAI22X1 U1862 ( .A(n2612), .B(n345), .C(n2613), .D(n395), .Y(n2124) );
  OAI22X1 U1863 ( .A(n2613), .B(n345), .C(n2614), .D(n395), .Y(n2125) );
  OAI22X1 U1864 ( .A(n2614), .B(n344), .C(n2615), .D(n395), .Y(n2126) );
  OAI22X1 U1865 ( .A(n2615), .B(n344), .C(n2616), .D(n394), .Y(n2127) );
  OAI22X1 U1866 ( .A(n2616), .B(n344), .C(n2617), .D(n394), .Y(n2128) );
  OAI22X1 U1867 ( .A(n2617), .B(n344), .C(n2618), .D(n394), .Y(n2129) );
  OAI22X1 U1868 ( .A(n2618), .B(n344), .C(n2619), .D(n394), .Y(n2130) );
  OAI22X1 U1869 ( .A(n2619), .B(n344), .C(n2620), .D(n394), .Y(n2131) );
  OAI22X1 U1870 ( .A(n2620), .B(n344), .C(n2621), .D(n394), .Y(n2132) );
  OAI22X1 U1871 ( .A(n2621), .B(n344), .C(n2622), .D(n394), .Y(n2133) );
  OAI22X1 U1872 ( .A(n2622), .B(n344), .C(n2623), .D(n394), .Y(n2134) );
  OAI22X1 U1873 ( .A(n2623), .B(n344), .C(n2624), .D(n394), .Y(n2135) );
  OAI22X1 U1874 ( .A(n2624), .B(n344), .C(n2625), .D(n394), .Y(n2136) );
  XNOR2X1 U1875 ( .A(n297), .B(n2969), .Y(n2594) );
  XNOR2X1 U1876 ( .A(n298), .B(n495), .Y(n2595) );
  XNOR2X1 U1877 ( .A(n297), .B(n2971), .Y(n2596) );
  XNOR2X1 U1878 ( .A(n297), .B(n491), .Y(n2597) );
  XNOR2X1 U1879 ( .A(n298), .B(n2973), .Y(n2598) );
  XNOR2X1 U1880 ( .A(n298), .B(n487), .Y(n2599) );
  XNOR2X1 U1881 ( .A(n297), .B(n2975), .Y(n2600) );
  XNOR2X1 U1882 ( .A(n297), .B(n483), .Y(n2601) );
  XNOR2X1 U1883 ( .A(n298), .B(n2977), .Y(n2602) );
  XNOR2X1 U1884 ( .A(n298), .B(n479), .Y(n2603) );
  XNOR2X1 U1885 ( .A(n297), .B(n2980), .Y(n2604) );
  XNOR2X1 U1886 ( .A(n297), .B(n475), .Y(n2605) );
  XNOR2X1 U1887 ( .A(n298), .B(n2983), .Y(n2606) );
  XNOR2X1 U1888 ( .A(n297), .B(n471), .Y(n2607) );
  XNOR2X1 U1889 ( .A(n298), .B(n2985), .Y(n2608) );
  XNOR2X1 U1890 ( .A(n297), .B(n467), .Y(n2609) );
  XNOR2X1 U1891 ( .A(n296), .B(n2988), .Y(n2610) );
  XNOR2X1 U1892 ( .A(n297), .B(n463), .Y(n2611) );
  XNOR2X1 U1893 ( .A(n297), .B(n2991), .Y(n2612) );
  XNOR2X1 U1894 ( .A(n296), .B(n459), .Y(n2613) );
  XNOR2X1 U1895 ( .A(n296), .B(n2994), .Y(n2614) );
  XNOR2X1 U1896 ( .A(n296), .B(n455), .Y(n2615) );
  XNOR2X1 U1897 ( .A(n298), .B(n2997), .Y(n2616) );
  XNOR2X1 U1898 ( .A(n297), .B(n451), .Y(n2617) );
  XNOR2X1 U1899 ( .A(n296), .B(n3000), .Y(n2618) );
  XNOR2X1 U1900 ( .A(n298), .B(n447), .Y(n2619) );
  XNOR2X1 U1901 ( .A(n296), .B(n3003), .Y(n2620) );
  XNOR2X1 U1902 ( .A(n296), .B(n443), .Y(n2621) );
  XNOR2X1 U1903 ( .A(n298), .B(n3006), .Y(n2622) );
  XNOR2X1 U1904 ( .A(n298), .B(n439), .Y(n2623) );
  XNOR2X1 U1905 ( .A(n296), .B(n3009), .Y(n2624) );
  XNOR2X1 U1906 ( .A(n296), .B(n3011), .Y(n2625) );
  OAI22X1 U1907 ( .A(n343), .B(n2659), .C(n2809), .D(n393), .Y(n1756) );
  OAI22X1 U1908 ( .A(n2809), .B(n343), .C(n2627), .D(n393), .Y(n2139) );
  OAI22X1 U1909 ( .A(n2627), .B(n343), .C(n2628), .D(n393), .Y(n2140) );
  OAI22X1 U1910 ( .A(n2628), .B(n343), .C(n2629), .D(n393), .Y(n2141) );
  OAI22X1 U1911 ( .A(n2629), .B(n343), .C(n2630), .D(n393), .Y(n2142) );
  OAI22X1 U1912 ( .A(n2630), .B(n343), .C(n2631), .D(n393), .Y(n2143) );
  OAI22X1 U1913 ( .A(n2631), .B(n343), .C(n2632), .D(n393), .Y(n2144) );
  OAI22X1 U1914 ( .A(n2632), .B(n343), .C(n2633), .D(n393), .Y(n2145) );
  OAI22X1 U1915 ( .A(n2633), .B(n343), .C(n2634), .D(n393), .Y(n2146) );
  OAI22X1 U1916 ( .A(n2634), .B(n343), .C(n2635), .D(n393), .Y(n2147) );
  OAI22X1 U1917 ( .A(n2635), .B(n342), .C(n2636), .D(n393), .Y(n2148) );
  OAI22X1 U1918 ( .A(n2636), .B(n342), .C(n2637), .D(n392), .Y(n2149) );
  OAI22X1 U1919 ( .A(n2637), .B(n342), .C(n2638), .D(n392), .Y(n2150) );
  OAI22X1 U1920 ( .A(n2638), .B(n342), .C(n2639), .D(n392), .Y(n2151) );
  OAI22X1 U1921 ( .A(n2639), .B(n342), .C(n2640), .D(n392), .Y(n2152) );
  OAI22X1 U1922 ( .A(n2640), .B(n342), .C(n2641), .D(n392), .Y(n2153) );
  OAI22X1 U1923 ( .A(n2641), .B(n342), .C(n2642), .D(n392), .Y(n2154) );
  OAI22X1 U1924 ( .A(n2642), .B(n342), .C(n2643), .D(n392), .Y(n2155) );
  OAI22X1 U1925 ( .A(n2643), .B(n342), .C(n2644), .D(n392), .Y(n2156) );
  OAI22X1 U1926 ( .A(n2644), .B(n342), .C(n2645), .D(n392), .Y(n2157) );
  OAI22X1 U1927 ( .A(n2645), .B(n342), .C(n2646), .D(n392), .Y(n2158) );
  OAI22X1 U1928 ( .A(n2646), .B(n342), .C(n2647), .D(n392), .Y(n2159) );
  OAI22X1 U1929 ( .A(n2647), .B(n341), .C(n2648), .D(n392), .Y(n2160) );
  OAI22X1 U1930 ( .A(n2648), .B(n341), .C(n2649), .D(n391), .Y(n2161) );
  OAI22X1 U1931 ( .A(n2649), .B(n341), .C(n2650), .D(n391), .Y(n2162) );
  OAI22X1 U1932 ( .A(n2650), .B(n341), .C(n2651), .D(n391), .Y(n2163) );
  OAI22X1 U1933 ( .A(n2651), .B(n341), .C(n2652), .D(n391), .Y(n2164) );
  OAI22X1 U1934 ( .A(n2652), .B(n341), .C(n2653), .D(n391), .Y(n2165) );
  OAI22X1 U1935 ( .A(n2653), .B(n341), .C(n2654), .D(n391), .Y(n2166) );
  OAI22X1 U1936 ( .A(n2654), .B(n341), .C(n2655), .D(n391), .Y(n2167) );
  OAI22X1 U1937 ( .A(n2655), .B(n341), .C(n2656), .D(n391), .Y(n2168) );
  OAI22X1 U1938 ( .A(n2656), .B(n341), .C(n2657), .D(n391), .Y(n2169) );
  OAI22X1 U1939 ( .A(n2657), .B(n341), .C(n2658), .D(n391), .Y(n2170) );
  XNOR2X1 U1940 ( .A(n295), .B(n2969), .Y(n2627) );
  XNOR2X1 U1941 ( .A(n295), .B(n495), .Y(n2628) );
  XNOR2X1 U1942 ( .A(n295), .B(n2971), .Y(n2629) );
  XNOR2X1 U1943 ( .A(n295), .B(n491), .Y(n2630) );
  XNOR2X1 U1944 ( .A(n295), .B(n2973), .Y(n2631) );
  XNOR2X1 U1945 ( .A(n295), .B(n487), .Y(n2632) );
  XNOR2X1 U1946 ( .A(n295), .B(n2975), .Y(n2633) );
  XNOR2X1 U1947 ( .A(n295), .B(n483), .Y(n2634) );
  XNOR2X1 U1948 ( .A(n295), .B(n2977), .Y(n2635) );
  XNOR2X1 U1949 ( .A(n295), .B(n479), .Y(n2636) );
  XNOR2X1 U1950 ( .A(n295), .B(n2980), .Y(n2637) );
  XNOR2X1 U1951 ( .A(n294), .B(n475), .Y(n2638) );
  XNOR2X1 U1952 ( .A(n294), .B(n2983), .Y(n2639) );
  XNOR2X1 U1953 ( .A(n294), .B(n471), .Y(n2640) );
  XNOR2X1 U1954 ( .A(n294), .B(n2985), .Y(n2641) );
  XNOR2X1 U1955 ( .A(n294), .B(n467), .Y(n2642) );
  XNOR2X1 U1956 ( .A(n294), .B(n2988), .Y(n2643) );
  XNOR2X1 U1957 ( .A(n294), .B(n463), .Y(n2644) );
  XNOR2X1 U1958 ( .A(n294), .B(n2991), .Y(n2645) );
  XNOR2X1 U1959 ( .A(n294), .B(n459), .Y(n2646) );
  XNOR2X1 U1960 ( .A(n294), .B(n2994), .Y(n2647) );
  XNOR2X1 U1961 ( .A(n294), .B(n455), .Y(n2648) );
  XNOR2X1 U1962 ( .A(n294), .B(n2997), .Y(n2649) );
  XNOR2X1 U1963 ( .A(n293), .B(n451), .Y(n2650) );
  XNOR2X1 U1964 ( .A(n293), .B(n3000), .Y(n2651) );
  XNOR2X1 U1965 ( .A(n293), .B(n447), .Y(n2652) );
  XNOR2X1 U1966 ( .A(n293), .B(n3003), .Y(n2653) );
  XNOR2X1 U1967 ( .A(n293), .B(n443), .Y(n2654) );
  XNOR2X1 U1968 ( .A(n293), .B(n3006), .Y(n2655) );
  XNOR2X1 U1969 ( .A(n293), .B(n439), .Y(n2656) );
  XNOR2X1 U1970 ( .A(n293), .B(n3009), .Y(n2657) );
  XNOR2X1 U1971 ( .A(n293), .B(n3011), .Y(n2658) );
  OAI22X1 U1972 ( .A(n340), .B(n2692), .C(n2810), .D(n390), .Y(n1757) );
  OAI22X1 U1973 ( .A(n2810), .B(n340), .C(n2660), .D(n390), .Y(n2173) );
  OAI22X1 U1974 ( .A(n2660), .B(n340), .C(n2661), .D(n390), .Y(n2174) );
  OAI22X1 U1975 ( .A(n2661), .B(n340), .C(n2662), .D(n390), .Y(n2175) );
  OAI22X1 U1976 ( .A(n2662), .B(n340), .C(n2663), .D(n390), .Y(n2176) );
  OAI22X1 U1977 ( .A(n2663), .B(n340), .C(n2664), .D(n390), .Y(n2177) );
  OAI22X1 U1978 ( .A(n2664), .B(n340), .C(n2665), .D(n390), .Y(n2178) );
  OAI22X1 U1979 ( .A(n2665), .B(n340), .C(n2666), .D(n390), .Y(n2179) );
  OAI22X1 U1980 ( .A(n2666), .B(n340), .C(n2667), .D(n390), .Y(n2180) );
  OAI22X1 U1981 ( .A(n2667), .B(n340), .C(n2668), .D(n390), .Y(n2181) );
  OAI22X1 U1982 ( .A(n2668), .B(n339), .C(n2669), .D(n390), .Y(n2182) );
  OAI22X1 U1983 ( .A(n2669), .B(n339), .C(n2670), .D(n389), .Y(n2183) );
  OAI22X1 U1984 ( .A(n2670), .B(n339), .C(n2671), .D(n389), .Y(n2184) );
  OAI22X1 U1985 ( .A(n2671), .B(n339), .C(n2672), .D(n389), .Y(n2185) );
  OAI22X1 U1986 ( .A(n2672), .B(n339), .C(n2673), .D(n389), .Y(n2186) );
  OAI22X1 U1987 ( .A(n2673), .B(n339), .C(n2674), .D(n389), .Y(n2187) );
  OAI22X1 U1988 ( .A(n2674), .B(n339), .C(n2675), .D(n389), .Y(n2188) );
  OAI22X1 U1989 ( .A(n2675), .B(n339), .C(n2676), .D(n389), .Y(n2189) );
  OAI22X1 U1990 ( .A(n2676), .B(n339), .C(n2677), .D(n389), .Y(n2190) );
  OAI22X1 U1991 ( .A(n2677), .B(n339), .C(n2678), .D(n389), .Y(n2191) );
  OAI22X1 U1992 ( .A(n2678), .B(n339), .C(n2679), .D(n389), .Y(n2192) );
  OAI22X1 U1993 ( .A(n2679), .B(n339), .C(n2680), .D(n389), .Y(n2193) );
  OAI22X1 U1994 ( .A(n2680), .B(n338), .C(n2681), .D(n389), .Y(n2194) );
  OAI22X1 U1995 ( .A(n2681), .B(n338), .C(n2682), .D(n388), .Y(n2195) );
  OAI22X1 U1996 ( .A(n2682), .B(n338), .C(n2683), .D(n388), .Y(n2196) );
  OAI22X1 U1997 ( .A(n2683), .B(n338), .C(n2684), .D(n388), .Y(n2197) );
  OAI22X1 U1998 ( .A(n2684), .B(n338), .C(n2685), .D(n388), .Y(n2198) );
  OAI22X1 U1999 ( .A(n2685), .B(n338), .C(n2686), .D(n388), .Y(n2199) );
  OAI22X1 U2000 ( .A(n2686), .B(n338), .C(n2687), .D(n388), .Y(n2200) );
  OAI22X1 U2001 ( .A(n2687), .B(n338), .C(n2688), .D(n388), .Y(n2201) );
  OAI22X1 U2002 ( .A(n2688), .B(n338), .C(n2689), .D(n388), .Y(n2202) );
  OAI22X1 U2003 ( .A(n2689), .B(n338), .C(n2690), .D(n388), .Y(n2203) );
  OAI22X1 U2004 ( .A(n2690), .B(n338), .C(n2691), .D(n388), .Y(n2204) );
  XNOR2X1 U2005 ( .A(n292), .B(n2969), .Y(n2660) );
  XNOR2X1 U2006 ( .A(n292), .B(n495), .Y(n2661) );
  XNOR2X1 U2007 ( .A(n292), .B(n2971), .Y(n2662) );
  XNOR2X1 U2008 ( .A(n292), .B(n491), .Y(n2663) );
  XNOR2X1 U2009 ( .A(n292), .B(n2973), .Y(n2664) );
  XNOR2X1 U2010 ( .A(n292), .B(n487), .Y(n2665) );
  XNOR2X1 U2011 ( .A(n292), .B(n2975), .Y(n2666) );
  XNOR2X1 U2012 ( .A(n292), .B(n483), .Y(n2667) );
  XNOR2X1 U2013 ( .A(n292), .B(n2977), .Y(n2668) );
  XNOR2X1 U2014 ( .A(n292), .B(n479), .Y(n2669) );
  XNOR2X1 U2015 ( .A(n292), .B(n2980), .Y(n2670) );
  XNOR2X1 U2016 ( .A(n2912), .B(n475), .Y(n2671) );
  XNOR2X1 U2017 ( .A(n2912), .B(n2983), .Y(n2672) );
  XNOR2X1 U2018 ( .A(n2912), .B(n471), .Y(n2673) );
  XNOR2X1 U2019 ( .A(n2912), .B(n2985), .Y(n2674) );
  XNOR2X1 U2020 ( .A(n2912), .B(n467), .Y(n2675) );
  XNOR2X1 U2021 ( .A(n2912), .B(n2988), .Y(n2676) );
  XNOR2X1 U2022 ( .A(n2912), .B(n463), .Y(n2677) );
  XNOR2X1 U2023 ( .A(n2912), .B(n2991), .Y(n2678) );
  XNOR2X1 U2024 ( .A(n2912), .B(n459), .Y(n2679) );
  XNOR2X1 U2025 ( .A(n2912), .B(n2994), .Y(n2680) );
  XNOR2X1 U2026 ( .A(n2912), .B(n455), .Y(n2681) );
  XNOR2X1 U2027 ( .A(n2912), .B(n2997), .Y(n2682) );
  XNOR2X1 U2028 ( .A(n2910), .B(n451), .Y(n2683) );
  XNOR2X1 U2029 ( .A(n2910), .B(n3000), .Y(n2684) );
  XNOR2X1 U2030 ( .A(n2910), .B(n447), .Y(n2685) );
  XNOR2X1 U2031 ( .A(n2909), .B(n3003), .Y(n2686) );
  XNOR2X1 U2032 ( .A(n2909), .B(n443), .Y(n2687) );
  XNOR2X1 U2033 ( .A(n2909), .B(n3006), .Y(n2688) );
  XNOR2X1 U2034 ( .A(n2910), .B(n439), .Y(n2689) );
  XNOR2X1 U2035 ( .A(n2910), .B(n3009), .Y(n2690) );
  XNOR2X1 U2036 ( .A(n2910), .B(n3011), .Y(n2691) );
  OAI22X1 U2037 ( .A(n3018), .B(n2725), .C(n3017), .D(n387), .Y(n1758) );
  OAI22X1 U2038 ( .A(n3018), .B(n3017), .C(n2693), .D(n387), .Y(n2207) );
  OAI22X1 U2039 ( .A(n3018), .B(n2693), .C(n2694), .D(n387), .Y(n2208) );
  OAI22X1 U2040 ( .A(n3018), .B(n2694), .C(n2695), .D(n387), .Y(n2209) );
  OAI22X1 U2041 ( .A(n3018), .B(n2695), .C(n2696), .D(n387), .Y(n2210) );
  OAI22X1 U2042 ( .A(n3018), .B(n2696), .C(n2697), .D(n387), .Y(n2211) );
  OAI22X1 U2043 ( .A(n3018), .B(n2697), .C(n2698), .D(n387), .Y(n2212) );
  OAI22X1 U2044 ( .A(n3018), .B(n2698), .C(n2699), .D(n387), .Y(n2213) );
  OAI22X1 U2045 ( .A(n3018), .B(n2699), .C(n2700), .D(n387), .Y(n2214) );
  OAI22X1 U2046 ( .A(n3018), .B(n2700), .C(n2701), .D(n387), .Y(n2215) );
  OAI22X1 U2047 ( .A(n3018), .B(n2701), .C(n2702), .D(n387), .Y(n2216) );
  OAI22X1 U2048 ( .A(n3018), .B(n2702), .C(n2703), .D(n386), .Y(n2217) );
  OAI22X1 U2049 ( .A(n3018), .B(n2703), .C(n2704), .D(n386), .Y(n2218) );
  OAI22X1 U2050 ( .A(n3019), .B(n2704), .C(n2705), .D(n386), .Y(n2219) );
  OAI22X1 U2051 ( .A(n3019), .B(n2705), .C(n2706), .D(n386), .Y(n2220) );
  OAI22X1 U2052 ( .A(n3019), .B(n2706), .C(n2707), .D(n386), .Y(n2221) );
  OAI22X1 U2053 ( .A(n3019), .B(n2707), .C(n2708), .D(n386), .Y(n2222) );
  OAI22X1 U2054 ( .A(n3019), .B(n2708), .C(n2709), .D(n386), .Y(n2223) );
  OAI22X1 U2055 ( .A(n3019), .B(n2709), .C(n2710), .D(n386), .Y(n2224) );
  OAI22X1 U2056 ( .A(n3019), .B(n2710), .C(n2711), .D(n386), .Y(n2225) );
  OAI22X1 U2057 ( .A(n3019), .B(n2711), .C(n2712), .D(n386), .Y(n2226) );
  OAI22X1 U2058 ( .A(n3019), .B(n2712), .C(n2713), .D(n386), .Y(n2227) );
  OAI22X1 U2059 ( .A(n3019), .B(n2713), .C(n2714), .D(n386), .Y(n2228) );
  OAI22X1 U2060 ( .A(n3019), .B(n2714), .C(n2715), .D(n385), .Y(n2229) );
  OAI22X1 U2061 ( .A(n3019), .B(n2715), .C(n2716), .D(n385), .Y(n2230) );
  OAI22X1 U2062 ( .A(n3019), .B(n2716), .C(n2717), .D(n385), .Y(n2231) );
  OAI22X1 U2063 ( .A(n3020), .B(n2717), .C(n2718), .D(n385), .Y(n2232) );
  OAI22X1 U2064 ( .A(n3020), .B(n2718), .C(n2719), .D(n385), .Y(n2233) );
  OAI22X1 U2065 ( .A(n3020), .B(n2719), .C(n2720), .D(n385), .Y(n2234) );
  OAI22X1 U2066 ( .A(n3020), .B(n2720), .C(n2721), .D(n385), .Y(n2235) );
  OAI22X1 U2067 ( .A(n3020), .B(n2721), .C(n2722), .D(n385), .Y(n2236) );
  OAI22X1 U2068 ( .A(n3020), .B(n2722), .C(n2723), .D(n385), .Y(n2237) );
  OAI22X1 U2069 ( .A(n3020), .B(n2723), .C(n2724), .D(n385), .Y(n2238) );
  XNOR2X1 U2070 ( .A(n3014), .B(n2969), .Y(n2693) );
  XNOR2X1 U2071 ( .A(n3014), .B(n495), .Y(n2694) );
  XNOR2X1 U2072 ( .A(n3014), .B(n2971), .Y(n2695) );
  XNOR2X1 U2073 ( .A(n3014), .B(n491), .Y(n2696) );
  XNOR2X1 U2074 ( .A(n3014), .B(n2973), .Y(n2697) );
  XNOR2X1 U2075 ( .A(n3014), .B(n487), .Y(n2698) );
  XNOR2X1 U2076 ( .A(n3015), .B(n2975), .Y(n2699) );
  XNOR2X1 U2077 ( .A(n3014), .B(n483), .Y(n2700) );
  XNOR2X1 U2078 ( .A(n3014), .B(n2977), .Y(n2701) );
  XNOR2X1 U2079 ( .A(n3014), .B(n479), .Y(n2702) );
  XNOR2X1 U2080 ( .A(n3014), .B(n2980), .Y(n2703) );
  XNOR2X1 U2081 ( .A(n3014), .B(n475), .Y(n2704) );
  XNOR2X1 U2082 ( .A(n3014), .B(n2983), .Y(n2705) );
  XNOR2X1 U2083 ( .A(n3015), .B(n471), .Y(n2706) );
  XNOR2X1 U2084 ( .A(n3015), .B(n2985), .Y(n2707) );
  XNOR2X1 U2085 ( .A(n3015), .B(n467), .Y(n2708) );
  XNOR2X1 U2086 ( .A(n3015), .B(n2988), .Y(n2709) );
  XNOR2X1 U2087 ( .A(n3015), .B(n463), .Y(n2710) );
  XNOR2X1 U2088 ( .A(n3015), .B(n2991), .Y(n2711) );
  XNOR2X1 U2089 ( .A(n3015), .B(n459), .Y(n2712) );
  XNOR2X1 U2090 ( .A(n3015), .B(n2994), .Y(n2713) );
  XNOR2X1 U2091 ( .A(n3015), .B(n455), .Y(n2714) );
  XNOR2X1 U2092 ( .A(n3015), .B(n2997), .Y(n2715) );
  XNOR2X1 U2093 ( .A(n3015), .B(n451), .Y(n2716) );
  XNOR2X1 U2094 ( .A(n3015), .B(n3000), .Y(n2717) );
  XNOR2X1 U2095 ( .A(n3015), .B(n447), .Y(n2718) );
  XNOR2X1 U2096 ( .A(n3015), .B(n3003), .Y(n2719) );
  XNOR2X1 U2097 ( .A(n3015), .B(n443), .Y(n2720) );
  XNOR2X1 U2098 ( .A(n3015), .B(n3006), .Y(n2721) );
  XNOR2X1 U2099 ( .A(n3015), .B(n439), .Y(n2722) );
  XNOR2X1 U2100 ( .A(n3015), .B(n3009), .Y(n2723) );
  XNOR2X1 U2101 ( .A(n3015), .B(n3011), .Y(n2724) );
  INVX2 U2102 ( .A(n334), .Y(n2796) );
  INVX2 U2104 ( .A(n2959), .Y(n2797) );
  INVX2 U2106 ( .A(n2965), .Y(n2798) );
  INVX2 U2108 ( .A(n325), .Y(n2799) );
  INVX2 U2110 ( .A(n2938), .Y(n2800) );
  INVX2 U2112 ( .A(n317), .Y(n2801) );
  INVX2 U2114 ( .A(n314), .Y(n2802) );
  INVX2 U2116 ( .A(n311), .Y(n2803) );
  INVX2 U2118 ( .A(n308), .Y(n2804) );
  INVX2 U2120 ( .A(n305), .Y(n2805) );
  INVX2 U2122 ( .A(n302), .Y(n2806) );
  INVX2 U2124 ( .A(n299), .Y(n2807) );
  INVX2 U2126 ( .A(n298), .Y(n2808) );
  INVX2 U2128 ( .A(n293), .Y(n2809) );
  INVX2 U2130 ( .A(n2910), .Y(n2810) );
  NAND2X1 U2135 ( .A(n2752), .B(n2780), .Y(n432) );
  XOR2X1 U2136 ( .A(a[30]), .B(a[31]), .Y(n2752) );
  XNOR2X1 U2137 ( .A(a[30]), .B(a[29]), .Y(n2780) );
  NAND2X1 U2138 ( .A(n2753), .B(n2781), .Y(n429) );
  XOR2X1 U2139 ( .A(a[28]), .B(a[29]), .Y(n2753) );
  XNOR2X1 U2140 ( .A(a[28]), .B(a[27]), .Y(n2781) );
  NAND2X1 U2141 ( .A(n2754), .B(n2782), .Y(n426) );
  XOR2X1 U2142 ( .A(a[26]), .B(a[27]), .Y(n2754) );
  XNOR2X1 U2143 ( .A(a[26]), .B(a[25]), .Y(n2782) );
  NAND2X1 U2144 ( .A(n2755), .B(n2783), .Y(n423) );
  XOR2X1 U2145 ( .A(a[24]), .B(a[25]), .Y(n2755) );
  XNOR2X1 U2146 ( .A(a[24]), .B(a[23]), .Y(n2783) );
  NAND2X1 U2147 ( .A(n2756), .B(n2784), .Y(n2768) );
  XOR2X1 U2148 ( .A(a[22]), .B(a[23]), .Y(n2756) );
  XNOR2X1 U2149 ( .A(a[22]), .B(a[21]), .Y(n2784) );
  NAND2X1 U2150 ( .A(n2757), .B(n2785), .Y(n2769) );
  XOR2X1 U2151 ( .A(a[20]), .B(a[21]), .Y(n2757) );
  XNOR2X1 U2152 ( .A(a[20]), .B(a[19]), .Y(n2785) );
  NAND2X1 U2153 ( .A(n2758), .B(n2786), .Y(n2770) );
  XOR2X1 U2154 ( .A(a[18]), .B(a[19]), .Y(n2758) );
  XNOR2X1 U2155 ( .A(a[18]), .B(a[17]), .Y(n2786) );
  NAND2X1 U2156 ( .A(n2759), .B(n2787), .Y(n2771) );
  XOR2X1 U2157 ( .A(a[16]), .B(a[17]), .Y(n2759) );
  XNOR2X1 U2158 ( .A(a[16]), .B(a[15]), .Y(n2787) );
  NAND2X1 U2159 ( .A(n2760), .B(n2788), .Y(n2772) );
  XOR2X1 U2160 ( .A(a[14]), .B(a[15]), .Y(n2760) );
  XNOR2X1 U2161 ( .A(a[14]), .B(a[13]), .Y(n2788) );
  NAND2X1 U2162 ( .A(n2761), .B(n2789), .Y(n2773) );
  XOR2X1 U2163 ( .A(a[12]), .B(a[13]), .Y(n2761) );
  XNOR2X1 U2164 ( .A(a[12]), .B(a[11]), .Y(n2789) );
  NAND2X1 U2165 ( .A(n2762), .B(n2790), .Y(n2774) );
  XOR2X1 U2166 ( .A(a[10]), .B(a[11]), .Y(n2762) );
  XNOR2X1 U2167 ( .A(a[10]), .B(a[9]), .Y(n2790) );
  NAND2X1 U2168 ( .A(n2763), .B(n2791), .Y(n2775) );
  XOR2X1 U2169 ( .A(a[8]), .B(a[9]), .Y(n2763) );
  XNOR2X1 U2170 ( .A(a[8]), .B(a[7]), .Y(n2791) );
  NAND2X1 U2171 ( .A(n2764), .B(n2792), .Y(n2776) );
  XOR2X1 U2172 ( .A(a[6]), .B(a[7]), .Y(n2764) );
  XNOR2X1 U2173 ( .A(a[6]), .B(a[5]), .Y(n2792) );
  NAND2X1 U2174 ( .A(n2765), .B(n2793), .Y(n2777) );
  XOR2X1 U2175 ( .A(a[4]), .B(a[5]), .Y(n2765) );
  XNOR2X1 U2176 ( .A(a[4]), .B(a[3]), .Y(n2793) );
  NAND2X1 U2177 ( .A(n2766), .B(n2794), .Y(n2778) );
  XOR2X1 U2178 ( .A(a[2]), .B(a[3]), .Y(n2766) );
  XNOR2X1 U2179 ( .A(a[2]), .B(n3014), .Y(n2794) );
  NAND2X1 U2180 ( .A(n3020), .B(n2767), .Y(n2779) );
  XOR2X1 U2181 ( .A(a[0]), .B(n3014), .Y(n2767) );
  INVX1 U2185 ( .A(n404), .Y(n179) );
  BUFX4 U2186 ( .A(n2779), .Y(n386) );
  BUFX4 U2187 ( .A(n2776), .Y(n395) );
  BUFX4 U2188 ( .A(n2813), .Y(n322) );
  BUFX4 U2189 ( .A(n2815), .Y(n315) );
  BUFX4 U2190 ( .A(n423), .Y(n422) );
  BUFX4 U2191 ( .A(n423), .Y(n421) );
  BUFX4 U2192 ( .A(n426), .Y(n424) );
  INVX1 U2193 ( .A(n650), .Y(n648) );
  BUFX2 U2194 ( .A(n290), .Y(n2909) );
  BUFX2 U2195 ( .A(n290), .Y(n2910) );
  INVX4 U2196 ( .A(n291), .Y(n2911) );
  INVX8 U2197 ( .A(n2911), .Y(n2912) );
  BUFX4 U2198 ( .A(n2813), .Y(n2938) );
  BUFX4 U2199 ( .A(n2813), .Y(n2939) );
  BUFX4 U2200 ( .A(n2813), .Y(n320) );
  BUFX4 U2201 ( .A(n330), .Y(n2913) );
  BUFX4 U2202 ( .A(n330), .Y(n2914) );
  BUFX4 U2203 ( .A(n2814), .Y(n317) );
  BUFX4 U2204 ( .A(n318), .Y(n2915) );
  BUFX4 U2205 ( .A(n318), .Y(n2916) );
  BUFX4 U2206 ( .A(n318), .Y(n2917) );
  BUFX2 U2207 ( .A(a[29]), .Y(n331) );
  BUFX2 U2208 ( .A(n329), .Y(n2958) );
  BUFX2 U2209 ( .A(n2815), .Y(n314) );
  BUFX2 U2210 ( .A(n2816), .Y(n311) );
  BUFX2 U2211 ( .A(n331), .Y(n329) );
  BUFX2 U2212 ( .A(n324), .Y(n2961) );
  BUFX2 U2213 ( .A(n2816), .Y(n312) );
  BUFX2 U2214 ( .A(n2823), .Y(n291) );
  BUFX2 U2215 ( .A(n329), .Y(n2960) );
  BUFX2 U2216 ( .A(n2818), .Y(n306) );
  BUFX2 U2217 ( .A(n2770), .Y(n412) );
  BUFX2 U2218 ( .A(a[7]), .Y(n2821) );
  BUFX2 U2219 ( .A(n327), .Y(n2940) );
  BUFX2 U2220 ( .A(n2774), .Y(n400) );
  BUFX2 U2221 ( .A(n2777), .Y(n392) );
  BUFX2 U2222 ( .A(n2772), .Y(n407) );
  BUFX2 U2223 ( .A(n2775), .Y(n398) );
  BUFX2 U2224 ( .A(n2768), .Y(n418) );
  BUFX2 U2225 ( .A(n2769), .Y(n415) );
  BUFX2 U2226 ( .A(n2774), .Y(n401) );
  BUFX2 U2227 ( .A(n2814), .Y(n318) );
  BUFX2 U2228 ( .A(n2772), .Y(n406) );
  BUFX2 U2229 ( .A(n2775), .Y(n397) );
  BUFX2 U2230 ( .A(a[3]), .Y(n2823) );
  BUFX2 U2231 ( .A(n2776), .Y(n396) );
  BUFX2 U2232 ( .A(n432), .Y(n430) );
  BUFX2 U2233 ( .A(n2777), .Y(n393) );
  BUFX2 U2234 ( .A(n2770), .Y(n413) );
  BUFX2 U2235 ( .A(n2780), .Y(n380) );
  BUFX2 U2236 ( .A(n2775), .Y(n399) );
  BUFX2 U2237 ( .A(n2773), .Y(n405) );
  BUFX2 U2238 ( .A(n2778), .Y(n390) );
  BUFX2 U2239 ( .A(n2823), .Y(n290) );
  BUFX2 U2240 ( .A(n2777), .Y(n391) );
  BUFX2 U2241 ( .A(n2769), .Y(n416) );
  BUFX2 U2242 ( .A(n325), .Y(n2962) );
  BUFX2 U2243 ( .A(a[17]), .Y(n2816) );
  BUFX2 U2244 ( .A(a[23]), .Y(n2813) );
  BUFX2 U2245 ( .A(a[19]), .Y(n2815) );
  BUFX2 U2246 ( .A(a[13]), .Y(n2818) );
  BUFX2 U2247 ( .A(n2771), .Y(n409) );
  BUFX2 U2248 ( .A(n2773), .Y(n404) );
  BUFX2 U2249 ( .A(n2774), .Y(n402) );
  INVX2 U2250 ( .A(a[0]), .Y(n3020) );
  BUFX2 U2251 ( .A(n2779), .Y(n387) );
  INVX4 U2252 ( .A(n3017), .Y(n3015) );
  BUFX2 U2253 ( .A(n2816), .Y(n313) );
  BUFX2 U2254 ( .A(n327), .Y(n2942) );
  BUFX2 U2255 ( .A(n327), .Y(n2941) );
  BUFX2 U2256 ( .A(a[21]), .Y(n2814) );
  BUFX2 U2257 ( .A(n2812), .Y(n323) );
  BUFX2 U2258 ( .A(n2812), .Y(n2937) );
  BUFX2 U2259 ( .A(n2772), .Y(n408) );
  BUFX2 U2260 ( .A(n2770), .Y(n414) );
  BUFX2 U2261 ( .A(n2771), .Y(n410) );
  BUFX2 U2262 ( .A(n331), .Y(n330) );
  INVX1 U2263 ( .A(n634), .Y(n632) );
  BUFX2 U2264 ( .A(n1230), .Y(n2918) );
  INVX1 U2265 ( .A(n615), .Y(n852) );
  OR2X2 U2266 ( .A(n1741), .B(n1740), .Y(n2919) );
  OR2X2 U2267 ( .A(n1719), .B(n1712), .Y(n2920) );
  OR2X2 U2268 ( .A(n1711), .B(n1704), .Y(n2921) );
  OR2X2 U2269 ( .A(n1645), .B(n1632), .Y(n2922) );
  OR2X2 U2270 ( .A(n1455), .B(n1432), .Y(n2923) );
  OR2X2 U2271 ( .A(n920), .B(n901), .Y(n2924) );
  OR2X2 U2272 ( .A(n1631), .B(n1616), .Y(n2925) );
  OR2X2 U2273 ( .A(n1501), .B(n1480), .Y(n2926) );
  OR2X2 U2274 ( .A(n2237), .B(n2953), .Y(n2927) );
  AND2X2 U2275 ( .A(n3012), .B(n2968), .Y(n2928) );
  AND2X2 U2276 ( .A(n3012), .B(n242), .Y(n2929) );
  AND2X2 U2277 ( .A(n3012), .B(n194), .Y(n2930) );
  AND2X2 U2278 ( .A(n3012), .B(n152), .Y(n2931) );
  AND2X2 U2279 ( .A(n3012), .B(n125), .Y(n2932) );
  AND2X2 U2280 ( .A(n3012), .B(n98), .Y(n2933) );
  BUFX2 U2281 ( .A(n2819), .Y(n303) );
  INVX2 U2282 ( .A(n582), .Y(n580) );
  BUFX2 U2283 ( .A(n2823), .Y(n292) );
  INVX2 U2284 ( .A(n667), .Y(n665) );
  AND2X2 U2285 ( .A(n843), .B(n2954), .Y(product[1]) );
  OR2X2 U2286 ( .A(n900), .B(n891), .Y(n2935) );
  INVX2 U2287 ( .A(n727), .Y(n726) );
  INVX2 U2288 ( .A(n698), .Y(n697) );
  BUFX4 U2289 ( .A(n84), .Y(n2967) );
  BUFX2 U2290 ( .A(n2817), .Y(n309) );
  BUFX2 U2291 ( .A(n2812), .Y(n2936) );
  BUFX4 U2292 ( .A(n84), .Y(n2968) );
  BUFX4 U2293 ( .A(n2821), .Y(n297) );
  BUFX4 U2294 ( .A(n2821), .Y(n298) );
  BUFX4 U2295 ( .A(n2821), .Y(n296) );
  BUFX2 U2296 ( .A(n2818), .Y(n307) );
  BUFX2 U2297 ( .A(n2817), .Y(n310) );
  BUFX2 U2298 ( .A(n2819), .Y(n304) );
  OR2X2 U2299 ( .A(n1758), .B(n2238), .Y(n2954) );
  INVX1 U2300 ( .A(n2926), .Y(n720) );
  INVX1 U2301 ( .A(n553), .Y(n551) );
  INVX1 U2302 ( .A(n623), .Y(n622) );
  INVX1 U2303 ( .A(n2925), .Y(n761) );
  BUFX2 U2304 ( .A(n2818), .Y(n305) );
  BUFX2 U2305 ( .A(n2817), .Y(n308) );
  INVX1 U2306 ( .A(n559), .Y(n557) );
  BUFX2 U2307 ( .A(n328), .Y(n327) );
  BUFX2 U2308 ( .A(a[9]), .Y(n2820) );
  BUFX2 U2309 ( .A(a[5]), .Y(n2822) );
  AND2X2 U2310 ( .A(n3012), .B(n143), .Y(n2946) );
  INVX1 U2311 ( .A(n364), .Y(n143) );
  AND2X2 U2312 ( .A(n3012), .B(n89), .Y(n2948) );
  INVX1 U2313 ( .A(n382), .Y(n89) );
  AND2X2 U2314 ( .A(n3012), .B(n168), .Y(n2947) );
  AND2X2 U2315 ( .A(n3012), .B(n184), .Y(n2949) );
  INVX1 U2316 ( .A(n355), .Y(n184) );
  AND2X2 U2317 ( .A(n3012), .B(n116), .Y(n2951) );
  INVX1 U2318 ( .A(n373), .Y(n116) );
  AND2X2 U2319 ( .A(n3012), .B(n210), .Y(n2950) );
  AND2X2 U2320 ( .A(n3012), .B(n232), .Y(n2952) );
  INVX1 U2321 ( .A(n346), .Y(n232) );
  AND2X2 U2322 ( .A(n3012), .B(n258), .Y(n2953) );
  AND2X2 U2323 ( .A(n3012), .B(a[0]), .Y(product[0]) );
  XNOR2X1 U2324 ( .A(n549), .B(n500), .Y(product[47]) );
  AND2X2 U2325 ( .A(n3012), .B(n134), .Y(n2956) );
  AND2X2 U2326 ( .A(n3012), .B(n107), .Y(n2957) );
  BUFX4 U2327 ( .A(a[27]), .Y(n328) );
  INVX2 U2328 ( .A(n581), .Y(n579) );
  INVX1 U2329 ( .A(n631), .Y(n629) );
  INVX1 U2330 ( .A(n648), .Y(n646) );
  INVX1 U2331 ( .A(n602), .Y(n596) );
  INVX2 U2332 ( .A(n668), .Y(n666) );
  INVX1 U2333 ( .A(n601), .Y(n599) );
  INVX1 U2334 ( .A(n669), .Y(n667) );
  XNOR2X1 U2335 ( .A(n707), .B(n2944), .Y(product[27]) );
  AND2X2 U2336 ( .A(n706), .B(n703), .Y(n2944) );
  OR2X2 U2337 ( .A(n554), .B(n581), .Y(n2945) );
  INVX1 U2338 ( .A(n718), .Y(n716) );
  BUFX2 U2339 ( .A(n323), .Y(n2963) );
  INVX1 U2340 ( .A(n592), .Y(n590) );
  INVX2 U2341 ( .A(n725), .Y(n723) );
  INVX1 U2342 ( .A(n696), .Y(n694) );
  INVX1 U2343 ( .A(n593), .Y(n591) );
  INVX1 U2344 ( .A(n706), .Y(n704) );
  INVX2 U2345 ( .A(n711), .Y(n709) );
  INVX1 U2346 ( .A(n624), .Y(n623) );
  BUFX2 U2347 ( .A(n2822), .Y(n294) );
  BUFX2 U2348 ( .A(n2820), .Y(n300) );
  BUFX2 U2349 ( .A(n2822), .Y(n295) );
  BUFX2 U2350 ( .A(n2820), .Y(n301) );
  BUFX2 U2351 ( .A(n2822), .Y(n293) );
  BUFX2 U2352 ( .A(n2820), .Y(n299) );
  BUFX2 U2353 ( .A(n2819), .Y(n302) );
  BUFX2 U2354 ( .A(n2815), .Y(n316) );
  BUFX2 U2355 ( .A(n2783), .Y(n372) );
  BUFX2 U2356 ( .A(n2794), .Y(n339) );
  BUFX2 U2357 ( .A(n2792), .Y(n345) );
  BUFX2 U2358 ( .A(n2791), .Y(n348) );
  BUFX2 U2359 ( .A(n2793), .Y(n342) );
  BUFX2 U2360 ( .A(n2788), .Y(n357) );
  BUFX2 U2361 ( .A(n2790), .Y(n351) );
  BUFX2 U2362 ( .A(n2784), .Y(n369) );
  BUFX2 U2363 ( .A(n2785), .Y(n366) );
  BUFX2 U2364 ( .A(n2786), .Y(n363) );
  BUFX2 U2365 ( .A(n2794), .Y(n340) );
  BUFX2 U2366 ( .A(n2792), .Y(n346) );
  BUFX2 U2367 ( .A(n2793), .Y(n343) );
  BUFX2 U2368 ( .A(n2791), .Y(n349) );
  BUFX2 U2369 ( .A(n2790), .Y(n352) );
  BUFX2 U2370 ( .A(n2788), .Y(n358) );
  BUFX2 U2371 ( .A(n2814), .Y(n319) );
  BUFX2 U2372 ( .A(n2789), .Y(n354) );
  BUFX2 U2373 ( .A(n2787), .Y(n360) );
  BUFX2 U2374 ( .A(n2789), .Y(n355) );
  BUFX2 U2375 ( .A(n426), .Y(n425) );
  BUFX2 U2376 ( .A(n2784), .Y(n368) );
  BUFX2 U2377 ( .A(n2785), .Y(n365) );
  BUFX2 U2378 ( .A(n2782), .Y(n374) );
  BUFX2 U2379 ( .A(n2783), .Y(n371) );
  BUFX2 U2380 ( .A(n2794), .Y(n338) );
  BUFX2 U2381 ( .A(n2792), .Y(n344) );
  BUFX2 U2382 ( .A(n2793), .Y(n341) );
  BUFX2 U2383 ( .A(n2781), .Y(n377) );
  BUFX2 U2384 ( .A(n2791), .Y(n347) );
  BUFX2 U2385 ( .A(n2788), .Y(n356) );
  BUFX2 U2386 ( .A(n2790), .Y(n350) );
  BUFX2 U2387 ( .A(n2786), .Y(n362) );
  BUFX2 U2388 ( .A(n2787), .Y(n359) );
  BUFX2 U2389 ( .A(n2789), .Y(n353) );
  BUFX2 U2390 ( .A(n2782), .Y(n375) );
  BUFX2 U2391 ( .A(n2779), .Y(n385) );
  BUFX2 U2392 ( .A(n2787), .Y(n361) );
  BUFX2 U2393 ( .A(n429), .Y(n428) );
  BUFX2 U2394 ( .A(n2781), .Y(n378) );
  BUFX2 U2395 ( .A(n2786), .Y(n364) );
  INVX1 U2396 ( .A(n759), .Y(n757) );
  BUFX2 U2397 ( .A(n2769), .Y(n417) );
  BUFX2 U2398 ( .A(n2780), .Y(n381) );
  BUFX2 U2399 ( .A(n2785), .Y(n367) );
  BUFX2 U2400 ( .A(n2812), .Y(n325) );
  INVX1 U2401 ( .A(n825), .Y(n824) );
  INVX1 U2402 ( .A(n574), .Y(n572) );
  BUFX2 U2403 ( .A(n2768), .Y(n420) );
  BUFX2 U2404 ( .A(n2784), .Y(n370) );
  INVX2 U2405 ( .A(n766), .Y(n764) );
  INVX1 U2406 ( .A(n783), .Y(n781) );
  INVX1 U2407 ( .A(n745), .Y(n743) );
  INVX1 U2408 ( .A(n784), .Y(n782) );
  INVX1 U2409 ( .A(n746), .Y(n744) );
  INVX1 U2410 ( .A(n575), .Y(n573) );
  INVX2 U2411 ( .A(n758), .Y(n756) );
  INVX1 U2412 ( .A(n774), .Y(n772) );
  BUFX2 U2413 ( .A(n2781), .Y(n379) );
  BUFX2 U2414 ( .A(n2782), .Y(n376) );
  INVX1 U2415 ( .A(n832), .Y(n830) );
  INVX1 U2416 ( .A(n840), .Y(n838) );
  INVX1 U2417 ( .A(n801), .Y(n799) );
  INVX1 U2418 ( .A(n812), .Y(n810) );
  INVX1 U2419 ( .A(a[0]), .Y(n3019) );
  INVX1 U2420 ( .A(a[0]), .Y(n3018) );
  BUFX2 U2421 ( .A(a[11]), .Y(n2819) );
  INVX2 U2422 ( .A(n800), .Y(n798) );
  INVX2 U2423 ( .A(n806), .Y(n804) );
  INVX2 U2424 ( .A(n843), .Y(n841) );
  INVX2 U2425 ( .A(n3013), .Y(n3011) );
  INVX2 U2426 ( .A(n3005), .Y(n3003) );
  INVX2 U2427 ( .A(n2970), .Y(n2969) );
  INVX1 U2428 ( .A(b[31]), .Y(n2970) );
  INVX2 U2429 ( .A(n3005), .Y(n3004) );
  INVX2 U2430 ( .A(n3013), .Y(n3012) );
  BUFX2 U2431 ( .A(b[2]), .Y(n439) );
  BUFX2 U2432 ( .A(b[14]), .Y(n463) );
  BUFX2 U2433 ( .A(b[26]), .Y(n487) );
  INVX2 U2434 ( .A(n3002), .Y(n3000) );
  INVX2 U2435 ( .A(n2996), .Y(n2994) );
  INVX2 U2436 ( .A(n2999), .Y(n2997) );
  INVX2 U2437 ( .A(n2990), .Y(n2988) );
  INVX2 U2438 ( .A(n2993), .Y(n2991) );
  INVX2 U2439 ( .A(n2984), .Y(n2983) );
  INVX2 U2440 ( .A(n2987), .Y(n2985) );
  INVX2 U2441 ( .A(n2982), .Y(n2980) );
  INVX2 U2442 ( .A(n3010), .Y(n3009) );
  INVX2 U2443 ( .A(n3008), .Y(n3006) );
  INVX2 U2444 ( .A(n2979), .Y(n2977) );
  INVX2 U2445 ( .A(n3002), .Y(n3001) );
  INVX2 U2446 ( .A(n2993), .Y(n2992) );
  INVX2 U2447 ( .A(n2999), .Y(n2998) );
  INVX2 U2448 ( .A(n2996), .Y(n2995) );
  INVX2 U2449 ( .A(n2990), .Y(n2989) );
  INVX2 U2450 ( .A(n2987), .Y(n2986) );
  INVX1 U2451 ( .A(b[5]), .Y(n3005) );
  INVX2 U2452 ( .A(n3008), .Y(n3007) );
  INVX1 U2453 ( .A(b[0]), .Y(n3013) );
  INVX2 U2454 ( .A(n2982), .Y(n2981) );
  INVX2 U2455 ( .A(n2979), .Y(n2978) );
  BUFX2 U2456 ( .A(b[28]), .Y(n491) );
  INVX2 U2457 ( .A(n2974), .Y(n2973) );
  INVX1 U2458 ( .A(b[27]), .Y(n2974) );
  INVX2 U2459 ( .A(n2972), .Y(n2971) );
  INVX1 U2460 ( .A(b[29]), .Y(n2972) );
  INVX1 U2461 ( .A(b[21]), .Y(n2982) );
  INVX1 U2462 ( .A(b[1]), .Y(n3010) );
  INVX1 U2463 ( .A(b[3]), .Y(n3008) );
  INVX1 U2464 ( .A(b[23]), .Y(n2979) );
  INVX2 U2465 ( .A(n2976), .Y(n2975) );
  INVX1 U2466 ( .A(b[25]), .Y(n2976) );
  INVX1 U2467 ( .A(b[17]), .Y(n2987) );
  BUFX2 U2468 ( .A(b[4]), .Y(n443) );
  INVX1 U2469 ( .A(b[7]), .Y(n3002) );
  INVX1 U2470 ( .A(b[11]), .Y(n2996) );
  INVX1 U2471 ( .A(b[13]), .Y(n2993) );
  INVX1 U2472 ( .A(b[9]), .Y(n2999) );
  INVX1 U2473 ( .A(b[15]), .Y(n2990) );
  INVX1 U2474 ( .A(b[19]), .Y(n2984) );
  BUFX4 U2475 ( .A(n329), .Y(n2959) );
  BUFX2 U2476 ( .A(n2812), .Y(n324) );
  BUFX2 U2477 ( .A(n326), .Y(n2964) );
  BUFX4 U2478 ( .A(n326), .Y(n2965) );
  BUFX4 U2479 ( .A(n326), .Y(n2966) );
  BUFX2 U2480 ( .A(n328), .Y(n326) );
  INVX1 U2481 ( .A(n384), .Y(n84) );
  BUFX4 U2482 ( .A(n334), .Y(n333) );
  BUFX2 U2483 ( .A(a[31]), .Y(n334) );
  BUFX2 U2484 ( .A(n2780), .Y(n382) );
  BUFX2 U2485 ( .A(b[24]), .Y(n483) );
  BUFX4 U2486 ( .A(n384), .Y(n383) );
  BUFX2 U2487 ( .A(b[8]), .Y(n451) );
  BUFX2 U2488 ( .A(b[6]), .Y(n447) );
  BUFX2 U2489 ( .A(b[18]), .Y(n471) );
  BUFX2 U2490 ( .A(n2783), .Y(n373) );
  BUFX2 U2491 ( .A(b[22]), .Y(n479) );
  BUFX2 U2492 ( .A(b[16]), .Y(n467) );
  BUFX2 U2493 ( .A(b[20]), .Y(n475) );
  BUFX2 U2494 ( .A(b[30]), .Y(n495) );
  BUFX2 U2495 ( .A(b[10]), .Y(n455) );
  BUFX2 U2496 ( .A(b[12]), .Y(n459) );
  BUFX2 U2497 ( .A(n2771), .Y(n411) );
  INVX1 U2498 ( .A(a[1]), .Y(n3017) );
  INVX1 U2499 ( .A(n633), .Y(n631) );
  INVX2 U2500 ( .A(n2918), .Y(n1231) );
  INVX2 U2501 ( .A(n705), .Y(n703) );
  BUFX2 U2502 ( .A(n2773), .Y(n403) );
  INVX1 U2503 ( .A(n682), .Y(n860) );
  INVX1 U2504 ( .A(n695), .Y(n693) );
  BUFX2 U2505 ( .A(a[15]), .Y(n2817) );
  INVX2 U2506 ( .A(n717), .Y(n715) );
  BUFX4 U2507 ( .A(a[25]), .Y(n2812) );
  BUFX2 U2508 ( .A(n432), .Y(n431) );
  INVX1 U2509 ( .A(n661), .Y(n659) );
  INVX2 U2510 ( .A(n643), .Y(n641) );
  INVX1 U2511 ( .A(n632), .Y(n630) );
  INVX1 U2512 ( .A(n653), .Y(n856) );
  INVX1 U2513 ( .A(n671), .Y(n858) );
  INVX1 U2514 ( .A(n390), .Y(n259) );
  INVX1 U2515 ( .A(n649), .Y(n647) );
  BUFX4 U2516 ( .A(n608), .Y(n499) );
  INVX1 U2517 ( .A(a[31]), .Y(n384) );
  INVX2 U2518 ( .A(n748), .Y(n747) );
  INVX1 U2519 ( .A(n660), .Y(n658) );
  BUFX4 U2520 ( .A(n429), .Y(n427) );
  INVX1 U2521 ( .A(n642), .Y(n640) );
  BUFX4 U2522 ( .A(n2768), .Y(n419) );
  INVX1 U2523 ( .A(n808), .Y(n807) );
  INVX1 U2524 ( .A(n786), .Y(n785) );
  BUFX4 U2525 ( .A(n2776), .Y(n394) );
  INVX1 U2526 ( .A(n670), .Y(n668) );
  BUFX4 U2527 ( .A(n2778), .Y(n389) );
  BUFX4 U2528 ( .A(n2778), .Y(n388) );
  INVX1 U2529 ( .A(n768), .Y(n767) );
  INVX1 U2530 ( .A(n795), .Y(n794) );
  INVX8 U2531 ( .A(n3016), .Y(n3014) );
  INVX4 U2532 ( .A(a[1]), .Y(n3016) );
endmodule


module poly5_DW01_sub_49 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   n1, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n42, n45, n46, n47, n48, n50,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n89, n90, n91, n92, n94, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282;

  XOR2X1 U3 ( .A(n3), .B(B[47]), .Y(DIFF[47]) );
  XOR2X1 U4 ( .A(n9), .B(B[46]), .Y(DIFF[46]) );
  NAND2X1 U7 ( .A(n6), .B(n32), .Y(n5) );
  NOR2X1 U8 ( .A(n7), .B(n19), .Y(n6) );
  NAND2X1 U9 ( .A(n8), .B(n12), .Y(n7) );
  XOR2X1 U11 ( .A(n13), .B(B[45]), .Y(DIFF[45]) );
  NAND2X1 U12 ( .A(n277), .B(n10), .Y(n9) );
  NOR2X1 U13 ( .A(n11), .B(n17), .Y(n10) );
  NOR2X1 U15 ( .A(B[45]), .B(B[44]), .Y(n12) );
  XOR2X1 U16 ( .A(B[44]), .B(n15), .Y(DIFF[44]) );
  NAND2X1 U17 ( .A(n276), .B(n14), .Y(n13) );
  NOR2X1 U18 ( .A(B[44]), .B(n17), .Y(n14) );
  XOR2X1 U19 ( .A(n21), .B(B[43]), .Y(DIFF[43]) );
  NAND2X1 U20 ( .A(n16), .B(n276), .Y(n15) );
  NAND2X1 U22 ( .A(n18), .B(n32), .Y(n17) );
  NAND2X1 U24 ( .A(n20), .B(n26), .Y(n19) );
  NOR2X1 U25 ( .A(B[43]), .B(B[42]), .Y(n20) );
  XOR2X1 U26 ( .A(n23), .B(B[42]), .Y(DIFF[42]) );
  NAND2X1 U27 ( .A(n277), .B(n22), .Y(n21) );
  NOR2X1 U28 ( .A(B[42]), .B(n25), .Y(n22) );
  XOR2X1 U29 ( .A(n27), .B(n273), .Y(DIFF[41]) );
  NAND2X1 U30 ( .A(n24), .B(n277), .Y(n23) );
  NAND2X1 U32 ( .A(n26), .B(n32), .Y(n25) );
  NOR2X1 U33 ( .A(B[41]), .B(B[40]), .Y(n26) );
  XOR2X1 U34 ( .A(n29), .B(B[40]), .Y(DIFF[40]) );
  NAND2X1 U35 ( .A(n28), .B(n276), .Y(n27) );
  NOR2X1 U36 ( .A(B[40]), .B(n31), .Y(n28) );
  XOR2X1 U37 ( .A(n35), .B(B[39]), .Y(DIFF[39]) );
  NAND2X1 U38 ( .A(n32), .B(n277), .Y(n29) );
  NOR2X1 U41 ( .A(n33), .B(n47), .Y(n32) );
  NAND2X1 U42 ( .A(n34), .B(n40), .Y(n33) );
  NOR2X1 U43 ( .A(B[39]), .B(B[38]), .Y(n34) );
  XOR2X1 U44 ( .A(n37), .B(B[38]), .Y(DIFF[38]) );
  NAND2X1 U45 ( .A(n36), .B(n276), .Y(n35) );
  NOR2X1 U46 ( .A(B[38]), .B(n39), .Y(n36) );
  NAND2X1 U48 ( .A(n38), .B(n277), .Y(n37) );
  NAND2X1 U50 ( .A(n40), .B(n46), .Y(n39) );
  NOR2X1 U51 ( .A(B[37]), .B(B[36]), .Y(n40) );
  NOR2X1 U54 ( .A(B[36]), .B(n45), .Y(n42) );
  NAND2X1 U60 ( .A(n48), .B(n54), .Y(n47) );
  NOR2X1 U61 ( .A(B[35]), .B(B[34]), .Y(n48) );
  NOR2X1 U64 ( .A(B[34]), .B(n53), .Y(n50) );
  XOR2X1 U65 ( .A(n55), .B(B[33]), .Y(DIFF[33]) );
  NOR2X1 U69 ( .A(B[33]), .B(B[32]), .Y(n54) );
  XNOR2X1 U70 ( .A(n1), .B(B[32]), .Y(DIFF[32]) );
  NAND2X1 U71 ( .A(n56), .B(n277), .Y(n55) );
  XOR2X1 U73 ( .A(n62), .B(B[31]), .Y(DIFF[31]) );
  NOR2X1 U74 ( .A(n123), .B(n58), .Y(n57) );
  NAND2X1 U75 ( .A(n59), .B(n97), .Y(n58) );
  NOR2X1 U76 ( .A(n60), .B(n80), .Y(n59) );
  NAND2X1 U77 ( .A(n61), .B(n71), .Y(n60) );
  NOR2X1 U78 ( .A(B[31]), .B(B[30]), .Y(n61) );
  XOR2X1 U79 ( .A(n66), .B(B[30]), .Y(DIFF[30]) );
  NAND2X1 U80 ( .A(n122), .B(n63), .Y(n62) );
  NOR2X1 U81 ( .A(n64), .B(n96), .Y(n63) );
  NAND2X1 U82 ( .A(n79), .B(n65), .Y(n64) );
  NOR2X1 U83 ( .A(B[30]), .B(n70), .Y(n65) );
  XOR2X1 U84 ( .A(n72), .B(B[29]), .Y(DIFF[29]) );
  NAND2X1 U85 ( .A(n122), .B(n67), .Y(n66) );
  NOR2X1 U86 ( .A(n68), .B(n96), .Y(n67) );
  NAND2X1 U87 ( .A(n71), .B(n79), .Y(n68) );
  NOR2X1 U90 ( .A(B[29]), .B(B[28]), .Y(n71) );
  XOR2X1 U91 ( .A(n76), .B(B[28]), .Y(DIFF[28]) );
  NAND2X1 U92 ( .A(n122), .B(n73), .Y(n72) );
  NOR2X1 U93 ( .A(n74), .B(n96), .Y(n73) );
  NAND2X1 U94 ( .A(n75), .B(n79), .Y(n74) );
  XOR2X1 U96 ( .A(n82), .B(B[27]), .Y(DIFF[27]) );
  NAND2X1 U97 ( .A(n122), .B(n77), .Y(n76) );
  NOR2X1 U98 ( .A(n80), .B(n96), .Y(n77) );
  NAND2X1 U101 ( .A(n81), .B(n91), .Y(n80) );
  NOR2X1 U102 ( .A(B[27]), .B(B[26]), .Y(n81) );
  XOR2X1 U103 ( .A(n86), .B(B[26]), .Y(DIFF[26]) );
  NAND2X1 U104 ( .A(n122), .B(n83), .Y(n82) );
  NOR2X1 U105 ( .A(n84), .B(n96), .Y(n83) );
  NAND2X1 U106 ( .A(n85), .B(n89), .Y(n84) );
  XOR2X1 U108 ( .A(n92), .B(B[25]), .Y(DIFF[25]) );
  NAND2X1 U109 ( .A(n122), .B(n87), .Y(n86) );
  NOR2X1 U110 ( .A(n90), .B(n96), .Y(n87) );
  NOR2X1 U114 ( .A(B[25]), .B(B[24]), .Y(n91) );
  XOR2X1 U115 ( .A(n94), .B(B[24]), .Y(DIFF[24]) );
  XOR2X1 U118 ( .A(n100), .B(B[23]), .Y(DIFF[23]) );
  NAND2X1 U119 ( .A(n97), .B(n122), .Y(n94) );
  NOR2X1 U122 ( .A(n98), .B(n112), .Y(n97) );
  NAND2X1 U123 ( .A(n99), .B(n105), .Y(n98) );
  NOR2X1 U124 ( .A(B[23]), .B(B[22]), .Y(n99) );
  XOR2X1 U125 ( .A(n102), .B(B[22]), .Y(DIFF[22]) );
  NAND2X1 U126 ( .A(n122), .B(n101), .Y(n100) );
  NOR2X1 U127 ( .A(B[22]), .B(n104), .Y(n101) );
  XOR2X1 U128 ( .A(n106), .B(B[21]), .Y(DIFF[21]) );
  NAND2X1 U129 ( .A(n103), .B(n122), .Y(n102) );
  NAND2X1 U131 ( .A(n105), .B(n111), .Y(n104) );
  NOR2X1 U132 ( .A(B[21]), .B(B[20]), .Y(n105) );
  XOR2X1 U133 ( .A(n108), .B(B[20]), .Y(DIFF[20]) );
  NAND2X1 U134 ( .A(n107), .B(n122), .Y(n106) );
  NOR2X1 U135 ( .A(B[20]), .B(n110), .Y(n107) );
  XOR2X1 U136 ( .A(n114), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U137 ( .A(n111), .B(n122), .Y(n108) );
  NAND2X1 U141 ( .A(n113), .B(n119), .Y(n112) );
  NOR2X1 U142 ( .A(B[19]), .B(B[18]), .Y(n113) );
  XOR2X1 U143 ( .A(n116), .B(B[18]), .Y(DIFF[18]) );
  NAND2X1 U144 ( .A(n115), .B(n122), .Y(n114) );
  NOR2X1 U145 ( .A(B[18]), .B(n118), .Y(n115) );
  XOR2X1 U146 ( .A(n120), .B(B[17]), .Y(DIFF[17]) );
  NAND2X1 U147 ( .A(n119), .B(n122), .Y(n116) );
  NOR2X1 U150 ( .A(B[17]), .B(B[16]), .Y(n119) );
  XNOR2X1 U151 ( .A(n122), .B(B[16]), .Y(DIFF[16]) );
  NAND2X1 U152 ( .A(n121), .B(n122), .Y(n120) );
  INVX4 U154 ( .A(n123), .Y(n122) );
  NAND2X1 U155 ( .A(n131), .B(n124), .Y(n123) );
  NOR2X1 U156 ( .A(n125), .B(n128), .Y(n124) );
  NAND2X1 U157 ( .A(n126), .B(n127), .Y(n125) );
  NOR2X1 U158 ( .A(B[15]), .B(B[14]), .Y(n126) );
  NOR2X1 U159 ( .A(B[13]), .B(B[12]), .Y(n127) );
  NAND2X1 U160 ( .A(n129), .B(n130), .Y(n128) );
  NOR2X1 U161 ( .A(B[11]), .B(B[10]), .Y(n129) );
  NOR2X1 U162 ( .A(B[9]), .B(B[8]), .Y(n130) );
  NOR2X1 U163 ( .A(n135), .B(n132), .Y(n131) );
  NAND2X1 U164 ( .A(n133), .B(n134), .Y(n132) );
  NOR2X1 U165 ( .A(B[7]), .B(B[6]), .Y(n133) );
  NOR2X1 U166 ( .A(B[5]), .B(B[4]), .Y(n134) );
  NAND2X1 U167 ( .A(n137), .B(n136), .Y(n135) );
  NOR2X1 U168 ( .A(B[3]), .B(B[2]), .Y(n136) );
  NOR2X1 U169 ( .A(B[0]), .B(B[1]), .Y(n137) );
  BUFX2 U173 ( .A(B[41]), .Y(n273) );
  INVX2 U174 ( .A(B[24]), .Y(n275) );
  BUFX2 U175 ( .A(n1), .Y(n276) );
  BUFX2 U176 ( .A(n1), .Y(n277) );
  INVX1 U177 ( .A(n32), .Y(n31) );
  INVX2 U178 ( .A(n97), .Y(n96) );
  NAND2X1 U179 ( .A(n275), .B(n122), .Y(n274) );
  INVX2 U180 ( .A(n90), .Y(n89) );
  OR2X2 U181 ( .A(n96), .B(n274), .Y(n92) );
  INVX2 U182 ( .A(n71), .Y(n70) );
  INVX2 U183 ( .A(n91), .Y(n90) );
  INVX2 U184 ( .A(n119), .Y(n118) );
  XOR2X1 U185 ( .A(n278), .B(B[36]), .Y(DIFF[36]) );
  NAND2X1 U186 ( .A(n46), .B(n276), .Y(n278) );
  XOR2X1 U187 ( .A(n279), .B(B[34]), .Y(DIFF[34]) );
  NAND2X1 U188 ( .A(n54), .B(n277), .Y(n279) );
  XOR2X1 U189 ( .A(n280), .B(B[35]), .Y(DIFF[35]) );
  NAND2X1 U190 ( .A(n50), .B(n276), .Y(n280) );
  XOR2X1 U191 ( .A(n281), .B(B[37]), .Y(DIFF[37]) );
  NAND2X1 U192 ( .A(n42), .B(n276), .Y(n281) );
  INVX1 U193 ( .A(n17), .Y(n16) );
  INVX2 U194 ( .A(n46), .Y(n45) );
  INVX1 U195 ( .A(n39), .Y(n38) );
  INVX1 U196 ( .A(n25), .Y(n24) );
  INVX2 U197 ( .A(n80), .Y(n79) );
  INVX1 U198 ( .A(n54), .Y(n53) );
  INVX2 U199 ( .A(n111), .Y(n110) );
  INVX1 U200 ( .A(B[32]), .Y(n56) );
  INVX1 U201 ( .A(B[28]), .Y(n75) );
  INVX1 U202 ( .A(B[26]), .Y(n85) );
  INVX2 U203 ( .A(n112), .Y(n111) );
  INVX1 U204 ( .A(B[16]), .Y(n121) );
  INVX1 U205 ( .A(B[46]), .Y(n8) );
  OR2X2 U206 ( .A(n282), .B(n5), .Y(n3) );
  INVX1 U207 ( .A(n57), .Y(n282) );
  BUFX2 U208 ( .A(n57), .Y(n1) );
  INVX1 U209 ( .A(n47), .Y(n46) );
  INVX1 U210 ( .A(n19), .Y(n18) );
  INVX1 U211 ( .A(n12), .Y(n11) );
  INVX1 U212 ( .A(n104), .Y(n103) );
endmodule


module poly5_DW01_sub_52 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, \B[0] ;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2X1 U1 ( .A(n1), .B(B[31]), .Y(DIFF[31]) );
  XOR2X1 U2 ( .A(n2), .B(B[30]), .Y(DIFF[30]) );
  NOR2X1 U3 ( .A(B[30]), .B(n2), .Y(n1) );
  XNOR2X1 U4 ( .A(n6), .B(B[29]), .Y(DIFF[29]) );
  NAND2X1 U5 ( .A(n24), .B(n3), .Y(n2) );
  NOR2X1 U6 ( .A(n10), .B(n4), .Y(n3) );
  NAND2X1 U7 ( .A(n8), .B(n5), .Y(n4) );
  XNOR2X1 U9 ( .A(n9), .B(B[28]), .Y(DIFF[28]) );
  NOR2X1 U10 ( .A(n23), .B(n7), .Y(n6) );
  NAND2X1 U11 ( .A(n8), .B(n11), .Y(n7) );
  XNOR2X1 U13 ( .A(n14), .B(B[27]), .Y(DIFF[27]) );
  NOR2X1 U14 ( .A(n10), .B(n23), .Y(n9) );
  NAND2X1 U17 ( .A(n19), .B(n13), .Y(n10) );
  NOR2X1 U18 ( .A(B[26]), .B(B[27]), .Y(n13) );
  XNOR2X1 U19 ( .A(n17), .B(B[26]), .Y(DIFF[26]) );
  NOR2X1 U20 ( .A(n15), .B(n23), .Y(n14) );
  NAND2X1 U21 ( .A(n16), .B(n19), .Y(n15) );
  XNOR2X1 U23 ( .A(n22), .B(B[25]), .Y(DIFF[25]) );
  NOR2X1 U24 ( .A(n18), .B(n23), .Y(n17) );
  NOR2X1 U28 ( .A(B[25]), .B(B[24]), .Y(n19) );
  XOR2X1 U29 ( .A(n23), .B(B[24]), .Y(DIFF[24]) );
  NOR2X1 U30 ( .A(B[24]), .B(n23), .Y(n22) );
  XOR2X1 U31 ( .A(n27), .B(B[23]), .Y(DIFF[23]) );
  NOR2X1 U33 ( .A(n36), .B(n25), .Y(n24) );
  NAND2X1 U34 ( .A(n26), .B(n30), .Y(n25) );
  NOR2X1 U35 ( .A(B[23]), .B(B[22]), .Y(n26) );
  XOR2X1 U36 ( .A(n29), .B(B[22]), .Y(DIFF[22]) );
  NAND2X1 U37 ( .A(n35), .B(n28), .Y(n27) );
  NOR2X1 U38 ( .A(B[22]), .B(n31), .Y(n28) );
  XOR2X1 U39 ( .A(n33), .B(B[21]), .Y(DIFF[21]) );
  NAND2X1 U40 ( .A(n30), .B(n35), .Y(n29) );
  NOR2X1 U43 ( .A(B[21]), .B(B[20]), .Y(n30) );
  XNOR2X1 U44 ( .A(n35), .B(B[20]), .Y(DIFF[20]) );
  NAND2X1 U45 ( .A(n34), .B(n35), .Y(n33) );
  XNOR2X1 U47 ( .A(n38), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U49 ( .A(n37), .B(n40), .Y(n36) );
  NOR2X1 U50 ( .A(B[19]), .B(B[18]), .Y(n37) );
  XOR2X1 U51 ( .A(n39), .B(B[18]), .Y(DIFF[18]) );
  NOR2X1 U52 ( .A(B[18]), .B(n39), .Y(n38) );
  XOR2X1 U53 ( .A(B[17]), .B(n41), .Y(DIFF[17]) );
  NOR2X1 U55 ( .A(B[17]), .B(n41), .Y(n40) );
  XNOR2X1 U56 ( .A(B[16]), .B(n43), .Y(DIFF[16]) );
  NAND2X1 U57 ( .A(n43), .B(n42), .Y(n41) );
  XOR2X1 U59 ( .A(n46), .B(B[15]), .Y(DIFF[15]) );
  NOR2X1 U60 ( .A(n51), .B(n44), .Y(n43) );
  NAND2X1 U61 ( .A(n45), .B(n47), .Y(n44) );
  XOR2X1 U63 ( .A(n48), .B(B[14]), .Y(DIFF[14]) );
  NAND2X1 U64 ( .A(n50), .B(n47), .Y(n46) );
  NOR2X1 U65 ( .A(B[13]), .B(B[14]), .Y(n47) );
  XNOR2X1 U66 ( .A(n50), .B(B[13]), .Y(DIFF[13]) );
  NAND2X1 U67 ( .A(n49), .B(n50), .Y(n48) );
  XNOR2X1 U69 ( .A(n53), .B(B[12]), .Y(DIFF[12]) );
  NAND2X1 U71 ( .A(n55), .B(n52), .Y(n51) );
  NOR2X1 U72 ( .A(B[11]), .B(B[12]), .Y(n52) );
  XOR2X1 U73 ( .A(n54), .B(B[11]), .Y(DIFF[11]) );
  NOR2X1 U74 ( .A(B[11]), .B(n54), .Y(n53) );
  XOR2X1 U75 ( .A(n58), .B(B[10]), .Y(DIFF[10]) );
  NOR2X1 U77 ( .A(n61), .B(n56), .Y(n55) );
  NAND2X1 U78 ( .A(n59), .B(n57), .Y(n56) );
  XNOR2X1 U80 ( .A(n60), .B(B[9]), .Y(DIFF[9]) );
  NAND2X1 U81 ( .A(n59), .B(n60), .Y(n58) );
  XNOR2X1 U83 ( .A(B[8]), .B(n63), .Y(DIFF[8]) );
  NAND2X1 U85 ( .A(n62), .B(n63), .Y(n61) );
  XOR2X1 U87 ( .A(n66), .B(B[7]), .Y(DIFF[7]) );
  NOR2X1 U88 ( .A(n64), .B(n69), .Y(n63) );
  NAND2X1 U89 ( .A(n67), .B(n65), .Y(n64) );
  XNOR2X1 U91 ( .A(n68), .B(B[6]), .Y(DIFF[6]) );
  NAND2X1 U92 ( .A(n67), .B(n68), .Y(n66) );
  XNOR2X1 U94 ( .A(n71), .B(B[5]), .Y(DIFF[5]) );
  NAND2X1 U96 ( .A(n73), .B(n70), .Y(n69) );
  NOR2X1 U97 ( .A(B[4]), .B(B[5]), .Y(n70) );
  XOR2X1 U98 ( .A(n72), .B(B[4]), .Y(DIFF[4]) );
  NOR2X1 U99 ( .A(B[4]), .B(n72), .Y(n71) );
  XOR2X1 U100 ( .A(n76), .B(B[3]), .Y(DIFF[3]) );
  NOR2X1 U102 ( .A(n79), .B(n74), .Y(n73) );
  NAND2X1 U103 ( .A(n75), .B(n77), .Y(n74) );
  XNOR2X1 U105 ( .A(n78), .B(B[2]), .Y(DIFF[2]) );
  NAND2X1 U106 ( .A(n77), .B(n78), .Y(n76) );
  XNOR2X1 U108 ( .A(B[1]), .B(n81), .Y(DIFF[1]) );
  NAND2X1 U110 ( .A(n81), .B(n80), .Y(n79) );
  INVX1 U116 ( .A(B[13]), .Y(n49) );
  INVX1 U117 ( .A(n55), .Y(n54) );
  INVX4 U118 ( .A(n24), .Y(n23) );
  INVX1 U119 ( .A(n40), .Y(n39) );
  INVX1 U120 ( .A(n51), .Y(n50) );
  INVX1 U121 ( .A(n69), .Y(n68) );
  INVX1 U122 ( .A(n61), .Y(n60) );
  INVX2 U123 ( .A(\B[0] ), .Y(n81) );
  INVX2 U124 ( .A(B[1]), .Y(n80) );
  INVX2 U125 ( .A(B[28]), .Y(n8) );
  INVX2 U126 ( .A(n79), .Y(n78) );
  INVX2 U127 ( .A(B[2]), .Y(n77) );
  INVX2 U128 ( .A(B[3]), .Y(n75) );
  INVX2 U129 ( .A(n73), .Y(n72) );
  INVX2 U130 ( .A(B[6]), .Y(n67) );
  INVX2 U131 ( .A(B[7]), .Y(n65) );
  INVX2 U132 ( .A(B[8]), .Y(n62) );
  INVX2 U133 ( .A(B[9]), .Y(n59) );
  INVX2 U134 ( .A(B[10]), .Y(n57) );
  INVX2 U135 ( .A(B[29]), .Y(n5) );
  INVX2 U136 ( .A(B[15]), .Y(n45) );
  INVX2 U137 ( .A(B[16]), .Y(n42) );
  INVX2 U138 ( .A(n36), .Y(n35) );
  INVX2 U139 ( .A(B[20]), .Y(n34) );
  INVX2 U140 ( .A(n30), .Y(n31) );
  INVX2 U141 ( .A(n19), .Y(n18) );
  INVX2 U142 ( .A(B[26]), .Y(n16) );
  INVX2 U143 ( .A(n10), .Y(n11) );
endmodule


module poly5_DW_mult_uns_41 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n8, n13, n18, n23, n28, n33, n38, n68, n80, n84, n89, n98, n107, n116,
         n125, n134, n143, n152, n162, n163, n178, n179, n194, n195, n210,
         n211, n227, n232, n242, n243, n258, n259, n274, n275, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n439, n443, n447, n451, n455, n459, n463, n467, n471, n475, n479,
         n483, n487, n491, n495, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n548, n549, n551, n553, n554,
         n555, n557, n559, n560, n561, n562, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n596, n599, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n664, n665, n667,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n709, n711, n712, n713, n714,
         n716, n718, n719, n720, n723, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n757, n759, n760, n761, n764, n766, n767, n768,
         n769, n770, n772, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n799, n801, n802, n804, n806, n807,
         n808, n810, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n830, n832, n833,
         n834, n835, n836, n838, n840, n841, n843, n846, n848, n850, n851,
         n852, n854, n856, n858, n859, n860, n861, n862, n864, n868, n869,
         n870, n872, n876, n878, n879, n883, n884, n885, n886, n888, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2240, n2242, n2244, n2246, n2248, n2250, n2252, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021;

  NAND2X1 OR_NOTi ( .A(n3021), .B(n289), .Y(n2725) );
  INVX2 U21 ( .A(n387), .Y(n275) );
  INVX2 U12 ( .A(n337), .Y(n274) );
  OAI21X1 AO21i ( .A(n274), .B(n275), .C(n288), .Y(n2206) );
  NAND2X1 OR_NOTi1 ( .A(n3021), .B(n292), .Y(n2692) );
  INVX2 U23 ( .A(n390), .Y(n259) );
  INVX2 U15 ( .A(n340), .Y(n258) );
  OAI21X1 AO21i1 ( .A(n258), .B(n259), .C(n290), .Y(n2172) );
  NAND2X1 OR_NOTi2 ( .A(n3021), .B(n295), .Y(n2659) );
  INVX2 U25 ( .A(n393), .Y(n243) );
  INVX2 U18 ( .A(n343), .Y(n242) );
  OAI21X1 AO21i2 ( .A(n242), .B(n243), .C(n294), .Y(n2138) );
  NAND2X1 OR_NOTi3 ( .A(n3021), .B(n298), .Y(n2626) );
  INVX2 U27 ( .A(n396), .Y(n227) );
  OAI21X1 AO21i3 ( .A(n232), .B(n227), .C(n298), .Y(n2104) );
  NAND2X1 OR_NOTi4 ( .A(n3021), .B(n301), .Y(n2593) );
  INVX2 U29 ( .A(n399), .Y(n211) );
  INVX2 U114 ( .A(n349), .Y(n210) );
  OAI21X1 AO21i4 ( .A(n210), .B(n211), .C(n301), .Y(n2070) );
  NAND2X1 OR_NOTi5 ( .A(n3021), .B(n304), .Y(n2560) );
  INVX2 U211 ( .A(n402), .Y(n195) );
  INVX2 U117 ( .A(n352), .Y(n194) );
  OAI21X1 AO21i5 ( .A(n194), .B(n195), .C(n303), .Y(n2036) );
  NAND2X1 OR_NOTi6 ( .A(n3021), .B(n307), .Y(n2527) );
  INVX2 U213 ( .A(n405), .Y(n179) );
  INVX2 U120 ( .A(n355), .Y(n178) );
  OAI21X1 AO21i6 ( .A(n178), .B(n179), .C(n306), .Y(n2002) );
  NAND2X1 OR_NOTi7 ( .A(n3021), .B(n310), .Y(n2494) );
  INVX2 U215 ( .A(n408), .Y(n163) );
  INVX2 U123 ( .A(n358), .Y(n162) );
  OAI21X1 AO21i7 ( .A(n162), .B(n163), .C(n309), .Y(n1968) );
  NAND2X1 OR_NOTi8 ( .A(n3021), .B(n311), .Y(n2461) );
  INVX2 U125 ( .A(n361), .Y(n152) );
  NAND2X1 OR_NOTi9 ( .A(n3021), .B(n316), .Y(n2428) );
  NAND2X1 OR_NOTi10 ( .A(n3021), .B(n319), .Y(n2397) );
  INVX2 U129 ( .A(n367), .Y(n134) );
  NAND2X1 OR_NOTi11 ( .A(n3021), .B(n322), .Y(n2368) );
  INVX2 U131 ( .A(n370), .Y(n125) );
  NAND2X1 OR_NOTi12 ( .A(n3021), .B(n324), .Y(n2341) );
  NAND2X1 OR_NOTi13 ( .A(n3021), .B(n328), .Y(n2316) );
  INVX2 U135 ( .A(n376), .Y(n107) );
  NAND2X1 OR_NOTi14 ( .A(n3021), .B(n331), .Y(n2293) );
  INVX2 U137 ( .A(n379), .Y(n98) );
  NAND2X1 OR_NOTi15 ( .A(n3021), .B(n334), .Y(n2272) );
  INVX2 U140 ( .A(n384), .Y(n84) );
  XOR2X1 U225 ( .A(n1759), .B(n918), .Y(n80) );
  XOR2X1 U141 ( .A(n1852), .B(n80), .Y(n899) );
  XOR2X1 U226 ( .A(n1768), .B(n1828), .Y(n68) );
  XOR2X1 U142 ( .A(n1786), .B(n68), .Y(n898) );
  XOR2X1 U227 ( .A(n1906), .B(n1806), .Y(n38) );
  XOR2X1 U143 ( .A(n1878), .B(n38), .Y(n897) );
  XOR2X1 U228 ( .A(n1968), .B(n1936), .Y(n33) );
  XOR2X1 U144 ( .A(n899), .B(n33), .Y(n896) );
  XOR2X1 U229 ( .A(n914), .B(n916), .Y(n28) );
  XOR2X1 U145 ( .A(n912), .B(n28), .Y(n895) );
  XOR2X1 U230 ( .A(n898), .B(n897), .Y(n23) );
  XOR2X1 U146 ( .A(n910), .B(n23), .Y(n894) );
  XOR2X1 U231 ( .A(n908), .B(n896), .Y(n18) );
  XOR2X1 U147 ( .A(n895), .B(n18), .Y(n893) );
  XOR2X1 U232 ( .A(n894), .B(n906), .Y(n13) );
  XOR2X1 U148 ( .A(n904), .B(n13), .Y(n892) );
  XOR2X1 U233 ( .A(n902), .B(n893), .Y(n8) );
  XOR2X1 U149 ( .A(n892), .B(n8), .Y(n891) );
  XNOR2X1 U292 ( .A(n549), .B(n500), .Y(product[47]) );
  NAND2X1 U293 ( .A(n548), .B(n2942), .Y(n500) );
  NAND2X1 U296 ( .A(n900), .B(n891), .Y(n548) );
  XNOR2X1 U297 ( .A(n560), .B(n501), .Y(product[46]) );
  OAI21X1 U298 ( .A(n2969), .B(n499), .C(n551), .Y(n549) );
  OAI21X1 U302 ( .A(n554), .B(n582), .C(n555), .Y(n553) );
  NAND2X1 U303 ( .A(n2931), .B(n565), .Y(n554) );
  AOI21X1 U304 ( .A(n2931), .B(n566), .C(n557), .Y(n555) );
  NAND2X1 U307 ( .A(n559), .B(n2931), .Y(n501) );
  NAND2X1 U310 ( .A(n920), .B(n901), .Y(n559) );
  XNOR2X1 U311 ( .A(n569), .B(n502), .Y(product[45]) );
  OAI21X1 U312 ( .A(n561), .B(n499), .C(n562), .Y(n560) );
  NAND2X1 U313 ( .A(n565), .B(n579), .Y(n561) );
  AOI21X1 U314 ( .A(n565), .B(n580), .C(n566), .Y(n562) );
  NOR2X1 U317 ( .A(n567), .B(n574), .Y(n565) );
  OAI21X1 U318 ( .A(n567), .B(n575), .C(n568), .Y(n566) );
  NAND2X1 U319 ( .A(n568), .B(n846), .Y(n502) );
  INVX2 U320 ( .A(n567), .Y(n846) );
  NOR2X1 U321 ( .A(n921), .B(n940), .Y(n567) );
  NAND2X1 U322 ( .A(n921), .B(n940), .Y(n568) );
  XNOR2X1 U323 ( .A(n576), .B(n503), .Y(product[44]) );
  OAI21X1 U324 ( .A(n570), .B(n499), .C(n571), .Y(n569) );
  NAND2X1 U325 ( .A(n572), .B(n579), .Y(n570) );
  AOI21X1 U326 ( .A(n572), .B(n580), .C(n573), .Y(n571) );
  NAND2X1 U329 ( .A(n575), .B(n572), .Y(n503) );
  NOR2X1 U331 ( .A(n962), .B(n941), .Y(n574) );
  NAND2X1 U332 ( .A(n962), .B(n941), .Y(n575) );
  XNOR2X1 U333 ( .A(n587), .B(n504), .Y(product[43]) );
  OAI21X1 U334 ( .A(n581), .B(n499), .C(n582), .Y(n576) );
  NAND2X1 U339 ( .A(n583), .B(n601), .Y(n581) );
  AOI21X1 U340 ( .A(n583), .B(n602), .C(n584), .Y(n582) );
  NOR2X1 U341 ( .A(n585), .B(n592), .Y(n583) );
  OAI21X1 U342 ( .A(n593), .B(n585), .C(n586), .Y(n584) );
  NAND2X1 U343 ( .A(n586), .B(n848), .Y(n504) );
  INVX2 U344 ( .A(n585), .Y(n848) );
  NOR2X1 U345 ( .A(n984), .B(n963), .Y(n585) );
  NAND2X1 U346 ( .A(n984), .B(n963), .Y(n586) );
  XNOR2X1 U347 ( .A(n594), .B(n505), .Y(product[42]) );
  OAI21X1 U348 ( .A(n588), .B(n499), .C(n589), .Y(n587) );
  NAND2X1 U349 ( .A(n590), .B(n601), .Y(n588) );
  AOI21X1 U350 ( .A(n590), .B(n602), .C(n591), .Y(n589) );
  NAND2X1 U353 ( .A(n593), .B(n590), .Y(n505) );
  NOR2X1 U355 ( .A(n1008), .B(n985), .Y(n592) );
  NAND2X1 U356 ( .A(n1008), .B(n985), .Y(n593) );
  XNOR2X1 U357 ( .A(n605), .B(n506), .Y(product[41]) );
  OAI21X1 U358 ( .A(n599), .B(n499), .C(n596), .Y(n594) );
  NOR2X1 U365 ( .A(n603), .B(n606), .Y(n601) );
  OAI21X1 U366 ( .A(n607), .B(n603), .C(n604), .Y(n602) );
  NAND2X1 U367 ( .A(n604), .B(n850), .Y(n506) );
  INVX2 U368 ( .A(n603), .Y(n850) );
  NOR2X1 U369 ( .A(n1032), .B(n1009), .Y(n603) );
  NAND2X1 U370 ( .A(n1032), .B(n1009), .Y(n604) );
  XOR2X1 U371 ( .A(n499), .B(n507), .Y(product[40]) );
  OAI21X1 U372 ( .A(n606), .B(n499), .C(n607), .Y(n605) );
  NAND2X1 U373 ( .A(n607), .B(n851), .Y(n507) );
  INVX2 U374 ( .A(n606), .Y(n851) );
  NOR2X1 U375 ( .A(n1058), .B(n1033), .Y(n606) );
  NAND2X1 U376 ( .A(n1058), .B(n1033), .Y(n607) );
  XNOR2X1 U377 ( .A(n617), .B(n508), .Y(product[39]) );
  AOI21X1 U378 ( .A(n677), .B(n609), .C(n610), .Y(n608) );
  NOR2X1 U379 ( .A(n649), .B(n611), .Y(n609) );
  OAI21X1 U380 ( .A(n611), .B(n650), .C(n612), .Y(n610) );
  NAND2X1 U381 ( .A(n613), .B(n633), .Y(n611) );
  AOI21X1 U382 ( .A(n634), .B(n613), .C(n614), .Y(n612) );
  NOR2X1 U383 ( .A(n615), .B(n624), .Y(n613) );
  OAI21X1 U384 ( .A(n625), .B(n615), .C(n616), .Y(n614) );
  NAND2X1 U385 ( .A(n616), .B(n852), .Y(n508) );
  INVX2 U386 ( .A(n615), .Y(n852) );
  NOR2X1 U387 ( .A(n1084), .B(n1059), .Y(n615) );
  NAND2X1 U388 ( .A(n1084), .B(n1059), .Y(n616) );
  XNOR2X1 U389 ( .A(n626), .B(n509), .Y(product[38]) );
  OAI21X1 U390 ( .A(n676), .B(n618), .C(n619), .Y(n617) );
  NAND2X1 U391 ( .A(n647), .B(n620), .Y(n618) );
  AOI21X1 U392 ( .A(n648), .B(n620), .C(n621), .Y(n619) );
  NOR2X1 U393 ( .A(n622), .B(n631), .Y(n620) );
  OAI21X1 U394 ( .A(n622), .B(n632), .C(n625), .Y(n621) );
  NAND2X1 U397 ( .A(n625), .B(n623), .Y(n509) );
  NOR2X1 U399 ( .A(n1112), .B(n1085), .Y(n624) );
  NAND2X1 U400 ( .A(n1112), .B(n1085), .Y(n625) );
  XNOR2X1 U401 ( .A(n637), .B(n510), .Y(product[37]) );
  OAI21X1 U402 ( .A(n676), .B(n627), .C(n628), .Y(n626) );
  NAND2X1 U403 ( .A(n629), .B(n647), .Y(n627) );
  AOI21X1 U404 ( .A(n629), .B(n648), .C(n634), .Y(n628) );
  NOR2X1 U409 ( .A(n635), .B(n642), .Y(n633) );
  OAI21X1 U410 ( .A(n643), .B(n635), .C(n636), .Y(n634) );
  NAND2X1 U411 ( .A(n636), .B(n854), .Y(n510) );
  INVX2 U412 ( .A(n635), .Y(n854) );
  NOR2X1 U413 ( .A(n1140), .B(n1113), .Y(n635) );
  NAND2X1 U414 ( .A(n1140), .B(n1113), .Y(n636) );
  XNOR2X1 U415 ( .A(n644), .B(n511), .Y(product[36]) );
  OAI21X1 U416 ( .A(n676), .B(n638), .C(n639), .Y(n637) );
  NAND2X1 U417 ( .A(n640), .B(n647), .Y(n638) );
  AOI21X1 U418 ( .A(n640), .B(n648), .C(n641), .Y(n639) );
  NAND2X1 U421 ( .A(n643), .B(n640), .Y(n511) );
  NOR2X1 U423 ( .A(n1170), .B(n1141), .Y(n642) );
  NAND2X1 U424 ( .A(n1170), .B(n1141), .Y(n643) );
  XNOR2X1 U425 ( .A(n655), .B(n512), .Y(product[35]) );
  OAI21X1 U426 ( .A(n649), .B(n676), .C(n646), .Y(n644) );
  NAND2X1 U431 ( .A(n669), .B(n651), .Y(n649) );
  AOI21X1 U432 ( .A(n670), .B(n651), .C(n652), .Y(n650) );
  NOR2X1 U433 ( .A(n653), .B(n660), .Y(n651) );
  OAI21X1 U434 ( .A(n661), .B(n653), .C(n654), .Y(n652) );
  NAND2X1 U435 ( .A(n654), .B(n856), .Y(n512) );
  INVX2 U436 ( .A(n653), .Y(n856) );
  NOR2X1 U437 ( .A(n1200), .B(n1171), .Y(n653) );
  NAND2X1 U438 ( .A(n1200), .B(n1171), .Y(n654) );
  XNOR2X1 U439 ( .A(n662), .B(n513), .Y(product[34]) );
  OAI21X1 U440 ( .A(n656), .B(n676), .C(n657), .Y(n655) );
  NAND2X1 U441 ( .A(n658), .B(n665), .Y(n656) );
  AOI21X1 U442 ( .A(n658), .B(n670), .C(n659), .Y(n657) );
  NAND2X1 U445 ( .A(n661), .B(n658), .Y(n513) );
  NOR2X1 U447 ( .A(n1232), .B(n1201), .Y(n660) );
  NAND2X1 U448 ( .A(n1232), .B(n1201), .Y(n661) );
  XNOR2X1 U449 ( .A(n673), .B(n514), .Y(product[33]) );
  OAI21X1 U450 ( .A(n667), .B(n676), .C(n664), .Y(n662) );
  NOR2X1 U457 ( .A(n674), .B(n671), .Y(n669) );
  OAI21X1 U458 ( .A(n675), .B(n671), .C(n672), .Y(n670) );
  NAND2X1 U459 ( .A(n672), .B(n858), .Y(n514) );
  INVX2 U460 ( .A(n671), .Y(n858) );
  NOR2X1 U461 ( .A(n1263), .B(n1233), .Y(n671) );
  NAND2X1 U462 ( .A(n1263), .B(n1233), .Y(n672) );
  XOR2X1 U463 ( .A(n676), .B(n515), .Y(product[32]) );
  OAI21X1 U464 ( .A(n674), .B(n676), .C(n675), .Y(n673) );
  NAND2X1 U465 ( .A(n675), .B(n859), .Y(n515) );
  INVX2 U466 ( .A(n674), .Y(n859) );
  NOR2X1 U467 ( .A(n1293), .B(n1264), .Y(n674) );
  NAND2X1 U468 ( .A(n1293), .B(n1264), .Y(n675) );
  XNOR2X1 U469 ( .A(n684), .B(n516), .Y(product[31]) );
  INVX4 U470 ( .A(n677), .Y(n676) );
  OAI21X1 U471 ( .A(n698), .B(n678), .C(n679), .Y(n677) );
  NAND2X1 U472 ( .A(n688), .B(n680), .Y(n678) );
  AOI21X1 U473 ( .A(n689), .B(n680), .C(n681), .Y(n679) );
  NOR2X1 U474 ( .A(n685), .B(n682), .Y(n680) );
  OAI21X1 U475 ( .A(n686), .B(n682), .C(n683), .Y(n681) );
  NAND2X1 U476 ( .A(n683), .B(n860), .Y(n516) );
  NOR2X1 U478 ( .A(n1323), .B(n1294), .Y(n682) );
  NAND2X1 U479 ( .A(n1323), .B(n1294), .Y(n683) );
  XOR2X1 U480 ( .A(n687), .B(n517), .Y(product[30]) );
  OAI21X1 U481 ( .A(n685), .B(n687), .C(n686), .Y(n684) );
  NAND2X1 U482 ( .A(n686), .B(n861), .Y(n517) );
  INVX2 U483 ( .A(n685), .Y(n861) );
  NOR2X1 U484 ( .A(n1351), .B(n1324), .Y(n685) );
  NAND2X1 U485 ( .A(n1351), .B(n1324), .Y(n686) );
  XOR2X1 U486 ( .A(n692), .B(n518), .Y(product[29]) );
  AOI21X1 U487 ( .A(n688), .B(n697), .C(n689), .Y(n687) );
  NOR2X1 U488 ( .A(n695), .B(n690), .Y(n688) );
  OAI21X1 U489 ( .A(n696), .B(n690), .C(n691), .Y(n689) );
  NAND2X1 U490 ( .A(n691), .B(n862), .Y(n518) );
  INVX2 U491 ( .A(n690), .Y(n862) );
  NOR2X1 U492 ( .A(n1379), .B(n1352), .Y(n690) );
  NAND2X1 U493 ( .A(n1379), .B(n1352), .Y(n691) );
  XNOR2X1 U494 ( .A(n697), .B(n519), .Y(product[28]) );
  AOI21X1 U495 ( .A(n693), .B(n697), .C(n694), .Y(n692) );
  NAND2X1 U498 ( .A(n696), .B(n693), .Y(n519) );
  NOR2X1 U500 ( .A(n1405), .B(n1380), .Y(n695) );
  NAND2X1 U501 ( .A(n1405), .B(n1380), .Y(n696) );
  AOI21X1 U504 ( .A(n699), .B(n727), .C(n700), .Y(n698) );
  NOR2X1 U505 ( .A(n713), .B(n701), .Y(n699) );
  OAI21X1 U506 ( .A(n714), .B(n701), .C(n702), .Y(n700) );
  NAND2X1 U507 ( .A(n2930), .B(n703), .Y(n701) );
  AOI21X1 U508 ( .A(n709), .B(n864), .C(n704), .Y(n702) );
  NOR2X1 U513 ( .A(n1431), .B(n1406), .Y(n705) );
  NAND2X1 U514 ( .A(n1431), .B(n1406), .Y(n706) );
  XNOR2X1 U515 ( .A(n712), .B(n521), .Y(product[26]) );
  AOI21X1 U516 ( .A(n2930), .B(n712), .C(n709), .Y(n707) );
  NAND2X1 U519 ( .A(n711), .B(n2930), .Y(n521) );
  NAND2X1 U522 ( .A(n1455), .B(n1432), .Y(n711) );
  XNOR2X1 U523 ( .A(n719), .B(n522), .Y(product[25]) );
  OAI21X1 U524 ( .A(n713), .B(n726), .C(n714), .Y(n712) );
  NAND2X1 U525 ( .A(n2932), .B(n2923), .Y(n713) );
  AOI21X1 U526 ( .A(n723), .B(n2923), .C(n716), .Y(n714) );
  NAND2X1 U529 ( .A(n718), .B(n2923), .Y(n522) );
  NAND2X1 U532 ( .A(n1479), .B(n1456), .Y(n718) );
  XOR2X1 U533 ( .A(n726), .B(n523), .Y(product[24]) );
  OAI21X1 U534 ( .A(n720), .B(n726), .C(n725), .Y(n719) );
  NAND2X1 U539 ( .A(n725), .B(n2932), .Y(n523) );
  NAND2X1 U542 ( .A(n1501), .B(n1480), .Y(n725) );
  XNOR2X1 U543 ( .A(n734), .B(n524), .Y(product[23]) );
  OAI21X1 U545 ( .A(n748), .B(n728), .C(n729), .Y(n727) );
  NAND2X1 U546 ( .A(n738), .B(n730), .Y(n728) );
  AOI21X1 U547 ( .A(n730), .B(n739), .C(n731), .Y(n729) );
  NOR2X1 U548 ( .A(n735), .B(n732), .Y(n730) );
  OAI21X1 U549 ( .A(n736), .B(n732), .C(n733), .Y(n731) );
  NAND2X1 U550 ( .A(n733), .B(n868), .Y(n524) );
  NOR2X1 U552 ( .A(n1523), .B(n1502), .Y(n732) );
  NAND2X1 U553 ( .A(n1523), .B(n1502), .Y(n733) );
  XOR2X1 U554 ( .A(n737), .B(n525), .Y(product[22]) );
  OAI21X1 U555 ( .A(n735), .B(n737), .C(n736), .Y(n734) );
  NAND2X1 U556 ( .A(n736), .B(n869), .Y(n525) );
  INVX2 U557 ( .A(n735), .Y(n869) );
  NOR2X1 U558 ( .A(n1543), .B(n1524), .Y(n735) );
  NAND2X1 U559 ( .A(n1543), .B(n1524), .Y(n736) );
  XOR2X1 U560 ( .A(n742), .B(n526), .Y(product[21]) );
  AOI21X1 U561 ( .A(n738), .B(n747), .C(n739), .Y(n737) );
  NOR2X1 U562 ( .A(n745), .B(n740), .Y(n738) );
  OAI21X1 U563 ( .A(n746), .B(n740), .C(n741), .Y(n739) );
  NAND2X1 U564 ( .A(n741), .B(n870), .Y(n526) );
  INVX2 U565 ( .A(n740), .Y(n870) );
  NOR2X1 U566 ( .A(n1563), .B(n1544), .Y(n740) );
  NAND2X1 U567 ( .A(n1563), .B(n1544), .Y(n741) );
  XNOR2X1 U568 ( .A(n747), .B(n527), .Y(product[20]) );
  AOI21X1 U569 ( .A(n743), .B(n747), .C(n744), .Y(n742) );
  NAND2X1 U572 ( .A(n746), .B(n743), .Y(n527) );
  NOR2X1 U574 ( .A(n1581), .B(n1564), .Y(n745) );
  NAND2X1 U575 ( .A(n1581), .B(n1564), .Y(n746) );
  XNOR2X1 U576 ( .A(n753), .B(n528), .Y(product[19]) );
  AOI21X1 U578 ( .A(n749), .B(n768), .C(n750), .Y(n748) );
  NOR2X1 U579 ( .A(n751), .B(n754), .Y(n749) );
  OAI21X1 U580 ( .A(n751), .B(n755), .C(n752), .Y(n750) );
  NAND2X1 U581 ( .A(n752), .B(n872), .Y(n528) );
  INVX2 U582 ( .A(n751), .Y(n872) );
  NOR2X1 U583 ( .A(n1599), .B(n1582), .Y(n751) );
  NAND2X1 U584 ( .A(n1599), .B(n1582), .Y(n752) );
  XNOR2X1 U585 ( .A(n760), .B(n529), .Y(product[18]) );
  OAI21X1 U586 ( .A(n754), .B(n767), .C(n755), .Y(n753) );
  NAND2X1 U587 ( .A(n2933), .B(n2925), .Y(n754) );
  AOI21X1 U588 ( .A(n764), .B(n2925), .C(n757), .Y(n755) );
  NAND2X1 U591 ( .A(n759), .B(n2925), .Y(n529) );
  NAND2X1 U594 ( .A(n1615), .B(n1600), .Y(n759) );
  XOR2X1 U595 ( .A(n767), .B(n530), .Y(product[17]) );
  OAI21X1 U596 ( .A(n761), .B(n767), .C(n766), .Y(n760) );
  NAND2X1 U601 ( .A(n766), .B(n2933), .Y(n530) );
  NAND2X1 U604 ( .A(n1631), .B(n1616), .Y(n766) );
  XOR2X1 U605 ( .A(n775), .B(n531), .Y(product[16]) );
  OAI21X1 U607 ( .A(n786), .B(n769), .C(n770), .Y(n768) );
  NAND2X1 U608 ( .A(n2929), .B(n776), .Y(n769) );
  AOI21X1 U609 ( .A(n2929), .B(n777), .C(n772), .Y(n770) );
  NAND2X1 U612 ( .A(n774), .B(n2929), .Y(n531) );
  NAND2X1 U615 ( .A(n1645), .B(n1632), .Y(n774) );
  XOR2X1 U616 ( .A(n780), .B(n532), .Y(product[15]) );
  AOI21X1 U617 ( .A(n776), .B(n785), .C(n777), .Y(n775) );
  NOR2X1 U618 ( .A(n783), .B(n778), .Y(n776) );
  OAI21X1 U619 ( .A(n784), .B(n778), .C(n779), .Y(n777) );
  NAND2X1 U620 ( .A(n779), .B(n876), .Y(n532) );
  NOR2X1 U622 ( .A(n1659), .B(n1646), .Y(n778) );
  NAND2X1 U623 ( .A(n1659), .B(n1646), .Y(n779) );
  XNOR2X1 U624 ( .A(n785), .B(n533), .Y(product[14]) );
  AOI21X1 U625 ( .A(n781), .B(n785), .C(n782), .Y(n780) );
  NAND2X1 U628 ( .A(n784), .B(n781), .Y(n533) );
  NOR2X1 U630 ( .A(n1671), .B(n1660), .Y(n783) );
  NAND2X1 U631 ( .A(n1671), .B(n1660), .Y(n784) );
  XNOR2X1 U632 ( .A(n791), .B(n534), .Y(product[13]) );
  AOI21X1 U634 ( .A(n787), .B(n795), .C(n788), .Y(n786) );
  NOR2X1 U635 ( .A(n792), .B(n789), .Y(n787) );
  OAI21X1 U636 ( .A(n793), .B(n789), .C(n790), .Y(n788) );
  NAND2X1 U637 ( .A(n790), .B(n878), .Y(n534) );
  INVX2 U638 ( .A(n789), .Y(n878) );
  NOR2X1 U639 ( .A(n1683), .B(n1672), .Y(n789) );
  NAND2X1 U640 ( .A(n1683), .B(n1672), .Y(n790) );
  XOR2X1 U641 ( .A(n794), .B(n535), .Y(product[12]) );
  OAI21X1 U642 ( .A(n792), .B(n794), .C(n793), .Y(n791) );
  NAND2X1 U643 ( .A(n793), .B(n879), .Y(n535) );
  INVX2 U644 ( .A(n792), .Y(n879) );
  NOR2X1 U645 ( .A(n1693), .B(n1684), .Y(n792) );
  NAND2X1 U646 ( .A(n1693), .B(n1684), .Y(n793) );
  XOR2X1 U647 ( .A(n802), .B(n536), .Y(product[11]) );
  OAI21X1 U649 ( .A(n796), .B(n808), .C(n797), .Y(n795) );
  NAND2X1 U650 ( .A(n2928), .B(n2924), .Y(n796) );
  AOI21X1 U651 ( .A(n804), .B(n2924), .C(n799), .Y(n797) );
  NAND2X1 U654 ( .A(n801), .B(n2924), .Y(n536) );
  NAND2X1 U657 ( .A(n1703), .B(n1694), .Y(n801) );
  XNOR2X1 U658 ( .A(n807), .B(n537), .Y(product[10]) );
  AOI21X1 U659 ( .A(n2928), .B(n807), .C(n804), .Y(n802) );
  NAND2X1 U662 ( .A(n806), .B(n2928), .Y(n537) );
  NAND2X1 U665 ( .A(n1711), .B(n1704), .Y(n806) );
  XNOR2X1 U666 ( .A(n813), .B(n538), .Y(product[9]) );
  AOI21X1 U668 ( .A(n2927), .B(n813), .C(n810), .Y(n808) );
  NAND2X1 U671 ( .A(n812), .B(n2927), .Y(n538) );
  NAND2X1 U674 ( .A(n1719), .B(n1712), .Y(n812) );
  XOR2X1 U675 ( .A(n816), .B(n539), .Y(product[8]) );
  OAI21X1 U676 ( .A(n814), .B(n816), .C(n815), .Y(n813) );
  NAND2X1 U677 ( .A(n815), .B(n883), .Y(n539) );
  INVX2 U678 ( .A(n814), .Y(n883) );
  NOR2X1 U679 ( .A(n1725), .B(n1720), .Y(n814) );
  NAND2X1 U680 ( .A(n1725), .B(n1720), .Y(n815) );
  XNOR2X1 U681 ( .A(n821), .B(n540), .Y(product[7]) );
  AOI21X1 U682 ( .A(n825), .B(n817), .C(n818), .Y(n816) );
  NOR2X1 U683 ( .A(n822), .B(n819), .Y(n817) );
  OAI21X1 U684 ( .A(n823), .B(n819), .C(n820), .Y(n818) );
  NAND2X1 U685 ( .A(n820), .B(n884), .Y(n540) );
  INVX2 U686 ( .A(n819), .Y(n884) );
  NOR2X1 U687 ( .A(n1731), .B(n1726), .Y(n819) );
  NAND2X1 U688 ( .A(n1731), .B(n1726), .Y(n820) );
  XOR2X1 U689 ( .A(n541), .B(n824), .Y(product[6]) );
  OAI21X1 U690 ( .A(n822), .B(n824), .C(n823), .Y(n821) );
  NAND2X1 U691 ( .A(n823), .B(n885), .Y(n541) );
  INVX2 U692 ( .A(n822), .Y(n885) );
  NOR2X1 U693 ( .A(n1735), .B(n1732), .Y(n822) );
  NAND2X1 U694 ( .A(n1735), .B(n1732), .Y(n823) );
  XOR2X1 U695 ( .A(n542), .B(n828), .Y(product[5]) );
  OAI21X1 U697 ( .A(n826), .B(n828), .C(n827), .Y(n825) );
  NAND2X1 U698 ( .A(n827), .B(n886), .Y(n542) );
  INVX2 U699 ( .A(n826), .Y(n886) );
  NOR2X1 U700 ( .A(n1739), .B(n1736), .Y(n826) );
  NAND2X1 U701 ( .A(n1739), .B(n1736), .Y(n827) );
  XNOR2X1 U702 ( .A(n543), .B(n833), .Y(product[4]) );
  AOI21X1 U703 ( .A(n833), .B(n2926), .C(n830), .Y(n828) );
  NAND2X1 U706 ( .A(n832), .B(n2926), .Y(n543) );
  NAND2X1 U709 ( .A(n1741), .B(n1740), .Y(n832) );
  XOR2X1 U710 ( .A(n544), .B(n836), .Y(product[3]) );
  OAI21X1 U711 ( .A(n834), .B(n836), .C(n835), .Y(n833) );
  NAND2X1 U712 ( .A(n835), .B(n888), .Y(n544) );
  INVX2 U713 ( .A(n834), .Y(n888) );
  NOR2X1 U714 ( .A(n1757), .B(n1742), .Y(n834) );
  NAND2X1 U715 ( .A(n1757), .B(n1742), .Y(n835) );
  XNOR2X1 U716 ( .A(n545), .B(n841), .Y(product[2]) );
  AOI21X1 U717 ( .A(n841), .B(n2934), .C(n838), .Y(n836) );
  NAND2X1 U720 ( .A(n840), .B(n2934), .Y(n545) );
  NAND2X1 U723 ( .A(n2237), .B(n2977), .Y(n840) );
  NAND2X1 U729 ( .A(n1758), .B(n2238), .Y(n843) );
  FAX1 U730 ( .A(n905), .B(n922), .C(n903), .YC(n900), .YS(n901) );
  FAX1 U731 ( .A(n926), .B(n907), .C(n924), .YC(n902), .YS(n903) );
  FAX1 U732 ( .A(n911), .B(n928), .C(n909), .YC(n904), .YS(n905) );
  FAX1 U733 ( .A(n915), .B(n932), .C(n930), .YC(n906), .YS(n907) );
  FAX1 U734 ( .A(n934), .B(n917), .C(n913), .YC(n908), .YS(n909) );
  FAX1 U735 ( .A(n1829), .B(n938), .C(n936), .YC(n910), .YS(n911) );
  FAX1 U736 ( .A(n1853), .B(n1787), .C(n1807), .YC(n912), .YS(n913) );
  FAX1 U737 ( .A(n1907), .B(n1769), .C(n1879), .YC(n914), .YS(n915) );
  FAX1 U738 ( .A(n919), .B(n1969), .C(n1937), .YC(n916), .YS(n917) );
  INVX2 U739 ( .A(n918), .Y(n919) );
  FAX1 U740 ( .A(n925), .B(n942), .C(n923), .YC(n920), .YS(n921) );
  FAX1 U741 ( .A(n946), .B(n927), .C(n944), .YC(n922), .YS(n923) );
  FAX1 U742 ( .A(n948), .B(n931), .C(n929), .YC(n924), .YS(n925) );
  FAX1 U743 ( .A(n933), .B(n952), .C(n950), .YC(n926), .YS(n927) );
  FAX1 U744 ( .A(n954), .B(n935), .C(n937), .YC(n928), .YS(n929) );
  FAX1 U745 ( .A(n958), .B(n956), .C(n939), .YC(n930), .YS(n931) );
  FAX1 U746 ( .A(n1970), .B(n1938), .C(n2002), .YC(n932), .YS(n933) );
  FAX1 U747 ( .A(n1788), .B(n1908), .C(n1830), .YC(n934), .YS(n935) );
  FAX1 U748 ( .A(n1854), .B(n1770), .C(n1808), .YC(n936), .YS(n937) );
  FAX1 U749 ( .A(n960), .B(n1760), .C(n1880), .YC(n938), .YS(n939) );
  FAX1 U750 ( .A(n945), .B(n964), .C(n943), .YC(n940), .YS(n941) );
  FAX1 U751 ( .A(n968), .B(n947), .C(n966), .YC(n942), .YS(n943) );
  FAX1 U752 ( .A(n970), .B(n951), .C(n949), .YC(n944), .YS(n945) );
  FAX1 U753 ( .A(n953), .B(n974), .C(n972), .YC(n946), .YS(n947) );
  FAX1 U754 ( .A(n959), .B(n955), .C(n957), .YC(n948), .YS(n949) );
  FAX1 U755 ( .A(n980), .B(n976), .C(n978), .YC(n950), .YS(n951) );
  FAX1 U756 ( .A(n1909), .B(n1881), .C(n982), .YC(n952), .YS(n953) );
  FAX1 U757 ( .A(n1855), .B(n1809), .C(n1831), .YC(n954), .YS(n955) );
  FAX1 U758 ( .A(n1939), .B(n1771), .C(n1789), .YC(n956), .YS(n957) );
  FAX1 U759 ( .A(n961), .B(n2003), .C(n1971), .YC(n958), .YS(n959) );
  INVX2 U760 ( .A(n960), .Y(n961) );
  FAX1 U761 ( .A(n988), .B(n986), .C(n965), .YC(n962), .YS(n963) );
  FAX1 U762 ( .A(n990), .B(n969), .C(n967), .YC(n964), .YS(n965) );
  FAX1 U763 ( .A(n973), .B(n971), .C(n992), .YC(n966), .YS(n967) );
  FAX1 U764 ( .A(n996), .B(n994), .C(n975), .YC(n968), .YS(n969) );
  FAX1 U765 ( .A(n977), .B(n981), .C(n979), .YC(n970), .YS(n971) );
  FAX1 U766 ( .A(n1000), .B(n998), .C(n983), .YC(n972), .YS(n973) );
  FAX1 U767 ( .A(n2036), .B(n1004), .C(n1002), .YC(n974), .YS(n975) );
  FAX1 U768 ( .A(n2004), .B(n1832), .C(n1972), .YC(n976), .YS(n977) );
  FAX1 U769 ( .A(n1910), .B(n1810), .C(n1940), .YC(n978), .YS(n979) );
  FAX1 U770 ( .A(n1856), .B(n1772), .C(n1790), .YC(n980), .YS(n981) );
  FAX1 U771 ( .A(n1006), .B(n1761), .C(n1882), .YC(n982), .YS(n983) );
  FAX1 U772 ( .A(n989), .B(n1010), .C(n987), .YC(n984), .YS(n985) );
  FAX1 U773 ( .A(n1014), .B(n991), .C(n1012), .YC(n986), .YS(n987) );
  FAX1 U774 ( .A(n995), .B(n1016), .C(n993), .YC(n988), .YS(n989) );
  FAX1 U775 ( .A(n1020), .B(n1018), .C(n997), .YC(n990), .YS(n991) );
  FAX1 U776 ( .A(n1003), .B(n1001), .C(n1022), .YC(n992), .YS(n993) );
  FAX1 U777 ( .A(n1024), .B(n1005), .C(n999), .YC(n994), .YS(n995) );
  FAX1 U778 ( .A(n1030), .B(n1028), .C(n1026), .YC(n996), .YS(n997) );
  FAX1 U779 ( .A(n1911), .B(n1857), .C(n1883), .YC(n998), .YS(n999) );
  FAX1 U780 ( .A(n1811), .B(n1941), .C(n1833), .YC(n1000), .YS(n1001) );
  FAX1 U781 ( .A(n1973), .B(n1773), .C(n1791), .YC(n1002), .YS(n1003) );
  FAX1 U782 ( .A(n1007), .B(n2037), .C(n2005), .YC(n1004), .YS(n1005) );
  INVX2 U783 ( .A(n1006), .Y(n1007) );
  FAX1 U784 ( .A(n1013), .B(n1034), .C(n1011), .YC(n1008), .YS(n1009) );
  FAX1 U785 ( .A(n1038), .B(n1015), .C(n1036), .YC(n1010), .YS(n1011) );
  FAX1 U786 ( .A(n1019), .B(n1040), .C(n1017), .YC(n1012), .YS(n1013) );
  FAX1 U787 ( .A(n1023), .B(n1042), .C(n1021), .YC(n1014), .YS(n1015) );
  FAX1 U788 ( .A(n1029), .B(n1046), .C(n1044), .YC(n1016), .YS(n1017) );
  FAX1 U789 ( .A(n1050), .B(n1025), .C(n1027), .YC(n1018), .YS(n1019) );
  FAX1 U790 ( .A(n1052), .B(n1048), .C(n1031), .YC(n1020), .YS(n1021) );
  FAX1 U791 ( .A(n2038), .B(n2070), .C(n1054), .YC(n1022), .YS(n1023) );
  FAX1 U792 ( .A(n2006), .B(n1834), .C(n1974), .YC(n1024), .YS(n1025) );
  FAX1 U793 ( .A(n1942), .B(n1774), .C(n1858), .YC(n1026), .YS(n1027) );
  FAX1 U794 ( .A(n1884), .B(n1792), .C(n1812), .YC(n1028), .YS(n1029) );
  FAX1 U795 ( .A(n1056), .B(n1762), .C(n1912), .YC(n1030), .YS(n1031) );
  FAX1 U796 ( .A(n1037), .B(n1060), .C(n1035), .YC(n1032), .YS(n1033) );
  FAX1 U797 ( .A(n1064), .B(n1039), .C(n1062), .YC(n1034), .YS(n1035) );
  FAX1 U798 ( .A(n1043), .B(n1066), .C(n1041), .YC(n1036), .YS(n1037) );
  FAX1 U799 ( .A(n1047), .B(n1045), .C(n1068), .YC(n1038), .YS(n1039) );
  FAX1 U800 ( .A(n1053), .B(n1072), .C(n1070), .YC(n1040), .YS(n1041) );
  FAX1 U801 ( .A(n1051), .B(n1049), .C(n1074), .YC(n1042), .YS(n1043) );
  FAX1 U802 ( .A(n1078), .B(n1076), .C(n1055), .YC(n1044), .YS(n1045) );
  FAX1 U803 ( .A(n1943), .B(n1082), .C(n1080), .YC(n1046), .YS(n1047) );
  FAX1 U804 ( .A(n1975), .B(n1859), .C(n1913), .YC(n1048), .YS(n1049) );
  FAX1 U805 ( .A(n1835), .B(n2007), .C(n1813), .YC(n1050), .YS(n1051) );
  FAX1 U806 ( .A(n2039), .B(n1775), .C(n1793), .YC(n1052), .YS(n1053) );
  FAX1 U807 ( .A(n1057), .B(n2071), .C(n1885), .YC(n1054), .YS(n1055) );
  INVX2 U808 ( .A(n1056), .Y(n1057) );
  FAX1 U809 ( .A(n1063), .B(n1086), .C(n1061), .YC(n1058), .YS(n1059) );
  FAX1 U810 ( .A(n1090), .B(n1065), .C(n1088), .YC(n1060), .YS(n1061) );
  FAX1 U811 ( .A(n1094), .B(n1092), .C(n1067), .YC(n1062), .YS(n1063) );
  FAX1 U812 ( .A(n1073), .B(n1071), .C(n1069), .YC(n1064), .YS(n1065) );
  FAX1 U813 ( .A(n1100), .B(n1098), .C(n1096), .YC(n1066), .YS(n1067) );
  FAX1 U814 ( .A(n1079), .B(n1081), .C(n1075), .YC(n1068), .YS(n1069) );
  FAX1 U815 ( .A(n1104), .B(n1102), .C(n1077), .YC(n1070), .YS(n1071) );
  FAX1 U816 ( .A(n1108), .B(n1106), .C(n1083), .YC(n1072), .YS(n1073) );
  FAX1 U817 ( .A(n2072), .B(n2040), .C(n2104), .YC(n1074), .YS(n1075) );
  FAX1 U818 ( .A(n1860), .B(n2008), .C(n1976), .YC(n1076), .YS(n1077) );
  FAX1 U819 ( .A(n1914), .B(n1776), .C(n1836), .YC(n1078), .YS(n1079) );
  FAX1 U820 ( .A(n1886), .B(n1794), .C(n1814), .YC(n1080), .YS(n1081) );
  FAX1 U821 ( .A(n1110), .B(n1763), .C(n1944), .YC(n1082), .YS(n1083) );
  FAX1 U822 ( .A(n1089), .B(n1114), .C(n1087), .YC(n1084), .YS(n1085) );
  FAX1 U823 ( .A(n1118), .B(n1091), .C(n1116), .YC(n1086), .YS(n1087) );
  FAX1 U824 ( .A(n1095), .B(n1120), .C(n1093), .YC(n1088), .YS(n1089) );
  FAX1 U825 ( .A(n1099), .B(n1097), .C(n1122), .YC(n1090), .YS(n1091) );
  FAX1 U826 ( .A(n1128), .B(n1126), .C(n1124), .YC(n1092), .YS(n1093) );
  FAX1 U827 ( .A(n1105), .B(n1107), .C(n1101), .YC(n1094), .YS(n1095) );
  FAX1 U828 ( .A(n1132), .B(n1109), .C(n1103), .YC(n1096), .YS(n1097) );
  FAX1 U829 ( .A(n1136), .B(n1130), .C(n1134), .YC(n1098), .YS(n1099) );
  FAX1 U830 ( .A(n1915), .B(n1861), .C(n1138), .YC(n1100), .YS(n1101) );
  FAX1 U831 ( .A(n1945), .B(n1815), .C(n1837), .YC(n1102), .YS(n1103) );
  FAX1 U832 ( .A(n2009), .B(n1795), .C(n1977), .YC(n1104), .YS(n1105) );
  FAX1 U833 ( .A(n1887), .B(n2041), .C(n1777), .YC(n1106), .YS(n1107) );
  FAX1 U834 ( .A(n1111), .B(n2105), .C(n2073), .YC(n1108), .YS(n1109) );
  INVX2 U835 ( .A(n1110), .Y(n1111) );
  FAX1 U836 ( .A(n1117), .B(n1142), .C(n1115), .YC(n1112), .YS(n1113) );
  FAX1 U837 ( .A(n1146), .B(n1119), .C(n1144), .YC(n1114), .YS(n1115) );
  FAX1 U838 ( .A(n1123), .B(n1148), .C(n1121), .YC(n1116), .YS(n1117) );
  FAX1 U839 ( .A(n1127), .B(n1125), .C(n1150), .YC(n1118), .YS(n1119) );
  FAX1 U840 ( .A(n1154), .B(n1129), .C(n1152), .YC(n1120), .YS(n1121) );
  FAX1 U841 ( .A(n1137), .B(n1135), .C(n1156), .YC(n1122), .YS(n1123) );
  FAX1 U842 ( .A(n1162), .B(n1131), .C(n1133), .YC(n1124), .YS(n1125) );
  FAX1 U843 ( .A(n1160), .B(n1164), .C(n1139), .YC(n1126), .YS(n1127) );
  FAX1 U844 ( .A(n2138), .B(n1166), .C(n1158), .YC(n1128), .YS(n1129) );
  FAX1 U845 ( .A(n2074), .B(n2106), .C(n1888), .YC(n1130), .YS(n1131) );
  FAX1 U846 ( .A(n1862), .B(n2010), .C(n2042), .YC(n1132), .YS(n1133) );
  FAX1 U847 ( .A(n1978), .B(n1796), .C(n1838), .YC(n1134), .YS(n1135) );
  FAX1 U848 ( .A(n1916), .B(n1778), .C(n1816), .YC(n1136), .YS(n1137) );
  FAX1 U849 ( .A(n1168), .B(n1764), .C(n1946), .YC(n1138), .YS(n1139) );
  FAX1 U850 ( .A(n1145), .B(n1172), .C(n1143), .YC(n1140), .YS(n1141) );
  FAX1 U851 ( .A(n1176), .B(n1147), .C(n1174), .YC(n1142), .YS(n1143) );
  FAX1 U852 ( .A(n1151), .B(n1178), .C(n1149), .YC(n1144), .YS(n1145) );
  FAX1 U853 ( .A(n1155), .B(n1153), .C(n1180), .YC(n1146), .YS(n1147) );
  FAX1 U854 ( .A(n1184), .B(n1157), .C(n1182), .YC(n1148), .YS(n1149) );
  FAX1 U855 ( .A(n1163), .B(n1188), .C(n1186), .YC(n1150), .YS(n1151) );
  FAX1 U856 ( .A(n1159), .B(n1165), .C(n1161), .YC(n1152), .YS(n1153) );
  FAX1 U857 ( .A(n1194), .B(n1196), .C(n1167), .YC(n1154), .YS(n1155) );
  FAX1 U858 ( .A(n1198), .B(n1190), .C(n1192), .YC(n1156), .YS(n1157) );
  FAX1 U859 ( .A(n1947), .B(n1863), .C(n1917), .YC(n1158), .YS(n1159) );
  FAX1 U860 ( .A(n1979), .B(n1817), .C(n1839), .YC(n1160), .YS(n1161) );
  FAX1 U861 ( .A(n2043), .B(n1797), .C(n2011), .YC(n1162), .YS(n1163) );
  FAX1 U862 ( .A(n1889), .B(n2075), .C(n1779), .YC(n1164), .YS(n1165) );
  FAX1 U863 ( .A(n1169), .B(n2139), .C(n2107), .YC(n1166), .YS(n1167) );
  INVX2 U864 ( .A(n1168), .Y(n1169) );
  FAX1 U865 ( .A(n1175), .B(n1202), .C(n1173), .YC(n1170), .YS(n1171) );
  FAX1 U866 ( .A(n1206), .B(n1177), .C(n1204), .YC(n1172), .YS(n1173) );
  FAX1 U867 ( .A(n1181), .B(n1208), .C(n1179), .YC(n1174), .YS(n1175) );
  FAX1 U868 ( .A(n1185), .B(n1183), .C(n1210), .YC(n1176), .YS(n1177) );
  FAX1 U869 ( .A(n1214), .B(n1212), .C(n1187), .YC(n1178), .YS(n1179) );
  FAX1 U870 ( .A(n1218), .B(n1189), .C(n1216), .YC(n1180), .YS(n1181) );
  FAX1 U871 ( .A(n1195), .B(n1197), .C(n1193), .YC(n1182), .YS(n1183) );
  FAX1 U872 ( .A(n1224), .B(n1222), .C(n1191), .YC(n1184), .YS(n1185) );
  FAX1 U873 ( .A(n1220), .B(n1226), .C(n1199), .YC(n1186), .YS(n1187) );
  FAX1 U874 ( .A(n2076), .B(n2172), .C(n1228), .YC(n1188), .YS(n1189) );
  FAX1 U875 ( .A(n2108), .B(n2044), .C(n2140), .YC(n1190), .YS(n1191) );
  FAX1 U876 ( .A(n1864), .B(n1948), .C(n1890), .YC(n1192), .YS(n1193) );
  FAX1 U877 ( .A(n2012), .B(n1840), .C(n1818), .YC(n1194), .YS(n1195) );
  FAX1 U878 ( .A(n1918), .B(n1798), .C(n1780), .YC(n1196), .YS(n1197) );
  FAX1 U879 ( .A(n1230), .B(n1765), .C(n1980), .YC(n1198), .YS(n1199) );
  FAX1 U880 ( .A(n1205), .B(n1234), .C(n1203), .YC(n1200), .YS(n1201) );
  FAX1 U881 ( .A(n1238), .B(n1207), .C(n1236), .YC(n1202), .YS(n1203) );
  FAX1 U882 ( .A(n1240), .B(n1211), .C(n1209), .YC(n1204), .YS(n1205) );
  FAX1 U883 ( .A(n1217), .B(n1213), .C(n1242), .YC(n1206), .YS(n1207) );
  FAX1 U884 ( .A(n1246), .B(n1244), .C(n1215), .YC(n1208), .YS(n1209) );
  FAX1 U885 ( .A(n1250), .B(n1248), .C(n1219), .YC(n1210), .YS(n1211) );
  FAX1 U886 ( .A(n1225), .B(n1227), .C(n1223), .YC(n1212), .YS(n1213) );
  FAX1 U887 ( .A(n1256), .B(n1254), .C(n1221), .YC(n1214), .YS(n1215) );
  FAX1 U888 ( .A(n1252), .B(n1258), .C(n1229), .YC(n1216), .YS(n1217) );
  FAX1 U889 ( .A(n1981), .B(n2013), .C(n1260), .YC(n1218), .YS(n1219) );
  FAX1 U890 ( .A(n2045), .B(n1919), .C(n1949), .YC(n1220), .YS(n1221) );
  FAX1 U891 ( .A(n1865), .B(n2077), .C(n1891), .YC(n1222), .YS(n1223) );
  FAX1 U892 ( .A(n2109), .B(n1819), .C(n1841), .YC(n1224), .YS(n1225) );
  FAX1 U893 ( .A(n2141), .B(n1781), .C(n1799), .YC(n1226), .YS(n1227) );
  FAX1 U894 ( .A(n1766), .B(n1262), .C(n2173), .YC(n1228), .YS(n1229) );
  FAX1 U896 ( .A(n1237), .B(n1265), .C(n1235), .YC(n1232), .YS(n1233) );
  FAX1 U897 ( .A(n1269), .B(n1239), .C(n1267), .YC(n1234), .YS(n1235) );
  FAX1 U898 ( .A(n1271), .B(n1243), .C(n1241), .YC(n1236), .YS(n1237) );
  FAX1 U899 ( .A(n1247), .B(n1245), .C(n1273), .YC(n1238), .YS(n1239) );
  FAX1 U900 ( .A(n1251), .B(n1275), .C(n1249), .YC(n1240), .YS(n1241) );
  FAX1 U901 ( .A(n1255), .B(n1279), .C(n1277), .YC(n1242), .YS(n1243) );
  FAX1 U902 ( .A(n1257), .B(n1259), .C(n1281), .YC(n1244), .YS(n1245) );
  FAX1 U903 ( .A(n1285), .B(n1261), .C(n1253), .YC(n1246), .YS(n1247) );
  FAX1 U904 ( .A(n1283), .B(n1289), .C(n1287), .YC(n1248), .YS(n1249) );
  FAX1 U905 ( .A(n2110), .B(n2206), .C(n1291), .YC(n1250), .YS(n1251) );
  FAX1 U906 ( .A(n2142), .B(n2078), .C(n2174), .YC(n1252), .YS(n1253) );
  FAX1 U907 ( .A(n1892), .B(n1982), .C(n1920), .YC(n1254), .YS(n1255) );
  FAX1 U908 ( .A(n2046), .B(n1866), .C(n1842), .YC(n1256), .YS(n1257) );
  FAX1 U909 ( .A(n1950), .B(n1820), .C(n1782), .YC(n1258), .YS(n1259) );
  FAX1 U910 ( .A(n1262), .B(n1800), .C(n2014), .YC(n1260), .YS(n1261) );
  INVX2 U911 ( .A(n1230), .Y(n1262) );
  FAX1 U912 ( .A(n1268), .B(n1295), .C(n1266), .YC(n1263), .YS(n1264) );
  FAX1 U913 ( .A(n1272), .B(n1270), .C(n1297), .YC(n1265), .YS(n1266) );
  FAX1 U914 ( .A(n1274), .B(n1301), .C(n1299), .YC(n1267), .YS(n1268) );
  FAX1 U915 ( .A(n1278), .B(n1276), .C(n1303), .YC(n1269), .YS(n1270) );
  FAX1 U916 ( .A(n1307), .B(n1305), .C(n1280), .YC(n1271), .YS(n1272) );
  FAX1 U917 ( .A(n1288), .B(n1282), .C(n1309), .YC(n1273), .YS(n1274) );
  FAX1 U918 ( .A(n1284), .B(n1290), .C(n1286), .YC(n1275), .YS(n1276) );
  FAX1 U919 ( .A(n1311), .B(n1315), .C(n1292), .YC(n1277), .YS(n1278) );
  FAX1 U920 ( .A(n1313), .B(n1319), .C(n1317), .YC(n1279), .YS(n1280) );
  FAX1 U921 ( .A(n2015), .B(n2047), .C(n1321), .YC(n1281), .YS(n1282) );
  FAX1 U922 ( .A(n2079), .B(n1921), .C(n1951), .YC(n1283), .YS(n1284) );
  FAX1 U923 ( .A(n2111), .B(n1867), .C(n1893), .YC(n1285), .YS(n1286) );
  FAX1 U924 ( .A(n1983), .B(n2143), .C(n1843), .YC(n1287), .YS(n1288) );
  FAX1 U925 ( .A(n2175), .B(n1801), .C(n1821), .YC(n1289), .YS(n1290) );
  FAX1 U926 ( .A(n2936), .B(n2207), .C(n1783), .YC(n1291), .YS(n1292) );
  FAX1 U927 ( .A(n1298), .B(n1325), .C(n1296), .YC(n1293), .YS(n1294) );
  FAX1 U928 ( .A(n1302), .B(n1300), .C(n1327), .YC(n1295), .YS(n1296) );
  FAX1 U929 ( .A(n1304), .B(n1331), .C(n1329), .YC(n1297), .YS(n1298) );
  FAX1 U930 ( .A(n1308), .B(n1333), .C(n1306), .YC(n1299), .YS(n1300) );
  FAX1 U931 ( .A(n1337), .B(n1310), .C(n1335), .YC(n1301), .YS(n1302) );
  FAX1 U932 ( .A(n1314), .B(n1316), .C(n1339), .YC(n1303), .YS(n1304) );
  FAX1 U933 ( .A(n1312), .B(n1320), .C(n1318), .YC(n1305), .YS(n1306) );
  FAX1 U934 ( .A(n1341), .B(n1345), .C(n1343), .YC(n1307), .YS(n1308) );
  FAX1 U935 ( .A(n1322), .B(n1349), .C(n1347), .YC(n1309), .YS(n1310) );
  FAX1 U936 ( .A(n1868), .B(n2016), .C(n1922), .YC(n1311), .YS(n1312) );
  FAX1 U937 ( .A(n2048), .B(n1822), .C(n1844), .YC(n1313), .YS(n1314) );
  FAX1 U938 ( .A(n1894), .B(n2112), .C(n2080), .YC(n1315), .YS(n1316) );
  FAX1 U939 ( .A(n1984), .B(n2176), .C(n2144), .YC(n1317), .YS(n1318) );
  FAX1 U940 ( .A(n1952), .B(n1784), .C(n1802), .YC(n1319), .YS(n1320) );
  HAX1 U941 ( .A(n2208), .B(n1743), .YC(n1321), .YS(n1322) );
  FAX1 U942 ( .A(n1328), .B(n1353), .C(n1326), .YC(n1323), .YS(n1324) );
  FAX1 U943 ( .A(n1332), .B(n1330), .C(n1355), .YC(n1325), .YS(n1326) );
  FAX1 U944 ( .A(n1334), .B(n1359), .C(n1357), .YC(n1327), .YS(n1328) );
  FAX1 U945 ( .A(n1361), .B(n1338), .C(n1336), .YC(n1329), .YS(n1330) );
  FAX1 U946 ( .A(n1365), .B(n1340), .C(n1363), .YC(n1331), .YS(n1332) );
  FAX1 U947 ( .A(n1344), .B(n1346), .C(n1367), .YC(n1333), .YS(n1334) );
  FAX1 U948 ( .A(n1350), .B(n1342), .C(n1348), .YC(n1335), .YS(n1336) );
  FAX1 U949 ( .A(n1371), .B(n1375), .C(n1373), .YC(n1337), .YS(n1338) );
  FAX1 U950 ( .A(n2972), .B(n1377), .C(n1369), .YC(n1339), .YS(n1340) );
  FAX1 U951 ( .A(n2017), .B(n1953), .C(n1985), .YC(n1341), .YS(n1342) );
  FAX1 U952 ( .A(n2049), .B(n1895), .C(n1923), .YC(n1343), .YS(n1344) );
  FAX1 U953 ( .A(n2081), .B(n1845), .C(n1869), .YC(n1345), .YS(n1346) );
  FAX1 U954 ( .A(n2145), .B(n1823), .C(n2113), .YC(n1347), .YS(n1348) );
  FAX1 U955 ( .A(n2209), .B(n2177), .C(n1803), .YC(n1349), .YS(n1350) );
  FAX1 U956 ( .A(n1356), .B(n1381), .C(n1354), .YC(n1351), .YS(n1352) );
  FAX1 U957 ( .A(n1385), .B(n1358), .C(n1383), .YC(n1353), .YS(n1354) );
  FAX1 U958 ( .A(n1362), .B(n1387), .C(n1360), .YC(n1355), .YS(n1356) );
  FAX1 U959 ( .A(n1366), .B(n1389), .C(n1364), .YC(n1357), .YS(n1358) );
  FAX1 U960 ( .A(n1368), .B(n1393), .C(n1391), .YC(n1359), .YS(n1360) );
  FAX1 U961 ( .A(n1374), .B(n1376), .C(n1395), .YC(n1361), .YS(n1362) );
  FAX1 U962 ( .A(n1401), .B(n1370), .C(n1372), .YC(n1363), .YS(n1364) );
  FAX1 U963 ( .A(n1403), .B(n1397), .C(n1399), .YC(n1365), .YS(n1366) );
  FAX1 U964 ( .A(n2018), .B(n2050), .C(n1378), .YC(n1367), .YS(n1368) );
  FAX1 U965 ( .A(n2082), .B(n1924), .C(n1954), .YC(n1369), .YS(n1370) );
  FAX1 U966 ( .A(n1846), .B(n1824), .C(n1870), .YC(n1371), .YS(n1372) );
  FAX1 U967 ( .A(n1896), .B(n2114), .C(n1804), .YC(n1373), .YS(n1374) );
  FAX1 U968 ( .A(n1986), .B(n2178), .C(n2146), .YC(n1375), .YS(n1376) );
  HAX1 U969 ( .A(n2210), .B(n1744), .YC(n1377), .YS(n1378) );
  FAX1 U970 ( .A(n1384), .B(n1407), .C(n1382), .YC(n1379), .YS(n1380) );
  FAX1 U971 ( .A(n1411), .B(n1386), .C(n1409), .YC(n1381), .YS(n1382) );
  FAX1 U972 ( .A(n1390), .B(n1413), .C(n1388), .YC(n1383), .YS(n1384) );
  FAX1 U973 ( .A(n1394), .B(n1415), .C(n1392), .YC(n1385), .YS(n1386) );
  FAX1 U974 ( .A(n1396), .B(n1419), .C(n1417), .YC(n1387), .YS(n1388) );
  FAX1 U975 ( .A(n1400), .B(n1398), .C(n1402), .YC(n1389), .YS(n1390) );
  FAX1 U976 ( .A(n1421), .B(n1423), .C(n1404), .YC(n1391), .YS(n1392) );
  FAX1 U977 ( .A(n1429), .B(n1427), .C(n1425), .YC(n1393), .YS(n1394) );
  FAX1 U978 ( .A(n2019), .B(n1987), .C(n2941), .YC(n1395), .YS(n1396) );
  FAX1 U979 ( .A(n2051), .B(n1925), .C(n1955), .YC(n1397), .YS(n1398) );
  FAX1 U980 ( .A(n2083), .B(n1871), .C(n1897), .YC(n1399), .YS(n1400) );
  FAX1 U981 ( .A(n2147), .B(n1847), .C(n2115), .YC(n1401), .YS(n1402) );
  FAX1 U982 ( .A(n2211), .B(n2179), .C(n1825), .YC(n1403), .YS(n1404) );
  FAX1 U983 ( .A(n1410), .B(n1433), .C(n1408), .YC(n1405), .YS(n1406) );
  FAX1 U984 ( .A(n1414), .B(n1412), .C(n1435), .YC(n1407), .YS(n1408) );
  FAX1 U985 ( .A(n1416), .B(n1439), .C(n1437), .YC(n1409), .YS(n1410) );
  FAX1 U986 ( .A(n1420), .B(n1418), .C(n1441), .YC(n1411), .YS(n1412) );
  FAX1 U987 ( .A(n1424), .B(n1445), .C(n1443), .YC(n1413), .YS(n1414) );
  FAX1 U988 ( .A(n1422), .B(n1428), .C(n1426), .YC(n1415), .YS(n1416) );
  FAX1 U989 ( .A(n1447), .B(n1449), .C(n1451), .YC(n1417), .YS(n1418) );
  FAX1 U990 ( .A(n2084), .B(n1430), .C(n1453), .YC(n1419), .YS(n1420) );
  FAX1 U991 ( .A(n2116), .B(n1956), .C(n2052), .YC(n1421), .YS(n1422) );
  FAX1 U992 ( .A(n2148), .B(n1898), .C(n1926), .YC(n1423), .YS(n1424) );
  FAX1 U993 ( .A(n2020), .B(n1872), .C(n2180), .YC(n1425), .YS(n1426) );
  FAX1 U994 ( .A(n1988), .B(n1826), .C(n1848), .YC(n1427), .YS(n1428) );
  HAX1 U995 ( .A(n2212), .B(n1745), .YC(n1429), .YS(n1430) );
  FAX1 U998 ( .A(n1444), .B(n1442), .C(n1440), .YC(n1435), .YS(n1436) );
  FAX1 U999 ( .A(n1467), .B(n1465), .C(n1463), .YC(n1437), .YS(n1438) );
  FAX1 U1000 ( .A(n1452), .B(n1450), .C(n1446), .YC(n1439), .YS(n1440) );
  FAX1 U1001 ( .A(n1473), .B(n1454), .C(n1448), .YC(n1441), .YS(n1442) );
  FAX1 U1002 ( .A(n1475), .B(n1469), .C(n1471), .YC(n1443), .YS(n1444) );
  FAX1 U1003 ( .A(n2053), .B(n2980), .C(n1477), .YC(n1445), .YS(n1446) );
  FAX1 U1004 ( .A(n2085), .B(n1989), .C(n2021), .YC(n1447), .YS(n1448) );
  FAX1 U1005 ( .A(n2117), .B(n1927), .C(n1957), .YC(n1449), .YS(n1450) );
  FAX1 U1006 ( .A(n2149), .B(n1873), .C(n1899), .YC(n1451), .YS(n1452) );
  FAX1 U1007 ( .A(n2213), .B(n2181), .C(n1849), .YC(n1453), .YS(n1454) );
  FAX1 U1008 ( .A(n1460), .B(n1481), .C(n1458), .YC(n1455), .YS(n1456) );
  FAX1 U1009 ( .A(n1485), .B(n1483), .C(n1462), .YC(n1457), .YS(n1458) );
  FAX1 U1010 ( .A(n1487), .B(n1466), .C(n1464), .YC(n1459), .YS(n1460) );
  FAX1 U1011 ( .A(n1491), .B(n1489), .C(n1468), .YC(n1461), .YS(n1462) );
  FAX1 U1012 ( .A(n1472), .B(n1476), .C(n1474), .YC(n1463), .YS(n1464) );
  FAX1 U1013 ( .A(n1495), .B(n1493), .C(n1470), .YC(n1465), .YS(n1466) );
  FAX1 U1014 ( .A(n1478), .B(n1499), .C(n1497), .YC(n1467), .YS(n1468) );
  FAX1 U1015 ( .A(n2086), .B(n1990), .C(n2054), .YC(n1469), .YS(n1470) );
  FAX1 U1016 ( .A(n2118), .B(n1900), .C(n1958), .YC(n1471), .YS(n1472) );
  FAX1 U1018 ( .A(n2022), .B(n2182), .C(n2150), .YC(n1475), .YS(n1476) );
  HAX1 U1019 ( .A(n2214), .B(n1746), .YC(n1477), .YS(n1478) );
  FAX1 U1020 ( .A(n1484), .B(n1503), .C(n1482), .YC(n1479), .YS(n1480) );
  FAX1 U1021 ( .A(n1507), .B(n1486), .C(n1505), .YC(n1481), .YS(n1482) );
  FAX1 U1022 ( .A(n1509), .B(n1490), .C(n1488), .YC(n1483), .YS(n1484) );
  FAX1 U1023 ( .A(n1513), .B(n1511), .C(n1492), .YC(n1485), .YS(n1486) );
  FAX1 U1024 ( .A(n1494), .B(n1498), .C(n1496), .YC(n1487), .YS(n1488) );
  FAX1 U1025 ( .A(n1517), .B(n1515), .C(n1500), .YC(n1489), .YS(n1490) );
  FAX1 U1026 ( .A(n2975), .B(n1521), .C(n1519), .YC(n1491), .YS(n1492) );
  FAX1 U1027 ( .A(n2087), .B(n2023), .C(n2055), .YC(n1493), .YS(n1494) );
  FAX1 U1028 ( .A(n2119), .B(n1959), .C(n1991), .YC(n1495), .YS(n1496) );
  FAX1 U1029 ( .A(n2151), .B(n1901), .C(n1929), .YC(n1497), .YS(n1498) );
  FAX1 U1030 ( .A(n2215), .B(n2183), .C(n1875), .YC(n1499), .YS(n1500) );
  FAX1 U1033 ( .A(n1531), .B(n1512), .C(n1510), .YC(n1505), .YS(n1506) );
  FAX1 U1034 ( .A(n1518), .B(n1514), .C(n1533), .YC(n1507), .YS(n1508) );
  FAX1 U1035 ( .A(n1516), .B(n1520), .C(n1535), .YC(n1509), .YS(n1510) );
  FAX1 U1036 ( .A(n1541), .B(n1539), .C(n1537), .YC(n1511), .YS(n1512) );
  FAX1 U1037 ( .A(n2088), .B(n1992), .C(n1522), .YC(n1513), .YS(n1514) );
  FAX1 U1038 ( .A(n2120), .B(n1930), .C(n1960), .YC(n1515), .YS(n1516) );
  FAX1 U1039 ( .A(n2056), .B(n2184), .C(n2152), .YC(n1517), .YS(n1518) );
  FAX1 U1040 ( .A(n2024), .B(n1876), .C(n1902), .YC(n1519), .YS(n1520) );
  HAX1 U1041 ( .A(n2216), .B(n1747), .YC(n1521), .YS(n1522) );
  FAX1 U1042 ( .A(n1528), .B(n1545), .C(n1526), .YC(n1523), .YS(n1524) );
  FAX1 U1043 ( .A(n1532), .B(n1530), .C(n1547), .YC(n1525), .YS(n1526) );
  FAX1 U1044 ( .A(n1551), .B(n1534), .C(n1549), .YC(n1527), .YS(n1528) );
  FAX1 U1045 ( .A(n1540), .B(n1536), .C(n1553), .YC(n1529), .YS(n1530) );
  FAX1 U1046 ( .A(n1555), .B(n1542), .C(n1538), .YC(n1531), .YS(n1532) );
  FAX1 U1047 ( .A(n1561), .B(n1559), .C(n1557), .YC(n1533), .YS(n1534) );
  FAX1 U1048 ( .A(n2089), .B(n2057), .C(n2940), .YC(n1535), .YS(n1536) );
  FAX1 U1049 ( .A(n2121), .B(n1993), .C(n2025), .YC(n1537), .YS(n1538) );
  FAX1 U1050 ( .A(n2153), .B(n1931), .C(n1961), .YC(n1539), .YS(n1540) );
  FAX1 U1051 ( .A(n2217), .B(n2185), .C(n1903), .YC(n1541), .YS(n1542) );
  FAX1 U1052 ( .A(n1548), .B(n1565), .C(n1546), .YC(n1543), .YS(n1544) );
  FAX1 U1053 ( .A(n1552), .B(n1550), .C(n1567), .YC(n1545), .YS(n1546) );
  FAX1 U1054 ( .A(n1571), .B(n1554), .C(n1569), .YC(n1547), .YS(n1548) );
  FAX1 U1055 ( .A(n1558), .B(n1560), .C(n1573), .YC(n1549), .YS(n1550) );
  FAX1 U1056 ( .A(n1577), .B(n1575), .C(n1556), .YC(n1551), .YS(n1552) );
  FAX1 U1057 ( .A(n1994), .B(n1562), .C(n1579), .YC(n1553), .YS(n1554) );
  FAX1 U1058 ( .A(n2058), .B(n1904), .C(n1932), .YC(n1555), .YS(n1556) );
  FAX1 U1059 ( .A(n1962), .B(n2122), .C(n2090), .YC(n1557), .YS(n1558) );
  FAX1 U1060 ( .A(n2026), .B(n2186), .C(n2154), .YC(n1559), .YS(n1560) );
  HAX1 U1061 ( .A(n2218), .B(n1748), .YC(n1561), .YS(n1562) );
  FAX1 U1062 ( .A(n1568), .B(n1583), .C(n1566), .YC(n1563), .YS(n1564) );
  FAX1 U1063 ( .A(n1572), .B(n1570), .C(n1585), .YC(n1565), .YS(n1566) );
  FAX1 U1064 ( .A(n1574), .B(n1589), .C(n1587), .YC(n1567), .YS(n1568) );
  FAX1 U1065 ( .A(n1580), .B(n1576), .C(n1578), .YC(n1569), .YS(n1570) );
  FAX1 U1066 ( .A(n1595), .B(n1591), .C(n1593), .YC(n1571), .YS(n1572) );
  FAX1 U1067 ( .A(n2091), .B(n2979), .C(n1597), .YC(n1573), .YS(n1574) );
  FAX1 U1068 ( .A(n2123), .B(n2027), .C(n2059), .YC(n1575), .YS(n1576) );
  FAX1 U1069 ( .A(n2155), .B(n1963), .C(n1995), .YC(n1577), .YS(n1578) );
  FAX1 U1070 ( .A(n2219), .B(n2187), .C(n1933), .YC(n1579), .YS(n1580) );
  FAX1 U1071 ( .A(n1586), .B(n1601), .C(n1584), .YC(n1581), .YS(n1582) );
  FAX1 U1072 ( .A(n1590), .B(n1588), .C(n1603), .YC(n1583), .YS(n1584) );
  FAX1 U1073 ( .A(n1596), .B(n1607), .C(n1605), .YC(n1585), .YS(n1586) );
  FAX1 U1074 ( .A(n1609), .B(n1592), .C(n1594), .YC(n1587), .YS(n1588) );
  FAX1 U1075 ( .A(n1598), .B(n1613), .C(n1611), .YC(n1589), .YS(n1590) );
  FAX1 U1076 ( .A(n2156), .B(n2028), .C(n2124), .YC(n1591), .YS(n1592) );
  FAX1 U1077 ( .A(n2092), .B(n2188), .C(n1996), .YC(n1593), .YS(n1594) );
  FAX1 U1078 ( .A(n2060), .B(n1934), .C(n1964), .YC(n1595), .YS(n1596) );
  HAX1 U1079 ( .A(n2220), .B(n1749), .YC(n1597), .YS(n1598) );
  FAX1 U1080 ( .A(n1604), .B(n1617), .C(n1602), .YC(n1599), .YS(n1600) );
  FAX1 U1081 ( .A(n1608), .B(n1606), .C(n1619), .YC(n1601), .YS(n1602) );
  FAX1 U1082 ( .A(n1612), .B(n1623), .C(n1621), .YC(n1603), .YS(n1604) );
  FAX1 U1083 ( .A(n1625), .B(n1614), .C(n1610), .YC(n1605), .YS(n1606) );
  FAX1 U1084 ( .A(n2970), .B(n1629), .C(n1627), .YC(n1607), .YS(n1608) );
  FAX1 U1085 ( .A(n2125), .B(n2061), .C(n2093), .YC(n1609), .YS(n1610) );
  FAX1 U1086 ( .A(n2157), .B(n1997), .C(n2029), .YC(n1611), .YS(n1612) );
  FAX1 U1087 ( .A(n2221), .B(n2189), .C(n1965), .YC(n1613), .YS(n1614) );
  FAX1 U1088 ( .A(n1620), .B(n1633), .C(n1618), .YC(n1615), .YS(n1616) );
  FAX1 U1089 ( .A(n1637), .B(n1622), .C(n1635), .YC(n1617), .YS(n1618) );
  FAX1 U1090 ( .A(n1628), .B(n1639), .C(n1624), .YC(n1619), .YS(n1620) );
  FAX1 U1091 ( .A(n1643), .B(n1641), .C(n1626), .YC(n1621), .YS(n1622) );
  FAX1 U1092 ( .A(n2094), .B(n2030), .C(n1630), .YC(n1623), .YS(n1624) );
  FAX1 U1093 ( .A(n2126), .B(n1966), .C(n1998), .YC(n1625), .YS(n1626) );
  FAX1 U1094 ( .A(n2062), .B(n2190), .C(n2158), .YC(n1627), .YS(n1628) );
  HAX1 U1095 ( .A(n2222), .B(n1750), .YC(n1629), .YS(n1630) );
  FAX1 U1096 ( .A(n1636), .B(n1647), .C(n1634), .YC(n1631), .YS(n1632) );
  FAX1 U1097 ( .A(n1651), .B(n1649), .C(n1638), .YC(n1633), .YS(n1634) );
  FAX1 U1098 ( .A(n1644), .B(n1642), .C(n1640), .YC(n1635), .YS(n1636) );
  FAX1 U1099 ( .A(n1657), .B(n1655), .C(n1653), .YC(n1637), .YS(n1638) );
  FAX1 U1100 ( .A(n2127), .B(n2095), .C(n2939), .YC(n1639), .YS(n1640) );
  FAX1 U1101 ( .A(n2159), .B(n2031), .C(n2063), .YC(n1641), .YS(n1642) );
  FAX1 U1102 ( .A(n2223), .B(n2191), .C(n1999), .YC(n1643), .YS(n1644) );
  FAX1 U1103 ( .A(n1650), .B(n1661), .C(n1648), .YC(n1645), .YS(n1646) );
  FAX1 U1104 ( .A(n1665), .B(n1663), .C(n1652), .YC(n1647), .YS(n1648) );
  FAX1 U1105 ( .A(n1667), .B(n1654), .C(n1656), .YC(n1649), .YS(n1650) );
  FAX1 U1106 ( .A(n2160), .B(n1658), .C(n1669), .YC(n1651), .YS(n1652) );
  FAX1 U1107 ( .A(n2192), .B(n2064), .C(n2128), .YC(n1653), .YS(n1654) );
  FAX1 U1108 ( .A(n2096), .B(n2000), .C(n2032), .YC(n1655), .YS(n1656) );
  HAX1 U1109 ( .A(n2224), .B(n1751), .YC(n1657), .YS(n1658) );
  FAX1 U1110 ( .A(n1664), .B(n1673), .C(n1662), .YC(n1659), .YS(n1660) );
  FAX1 U1111 ( .A(n1668), .B(n1666), .C(n1675), .YC(n1661), .YS(n1662) );
  FAX1 U1112 ( .A(n1679), .B(n1677), .C(n1670), .YC(n1663), .YS(n1664) );
  FAX1 U1113 ( .A(n2129), .B(n2971), .C(n1681), .YC(n1665), .YS(n1666) );
  FAX1 U1114 ( .A(n2161), .B(n2065), .C(n2097), .YC(n1667), .YS(n1668) );
  FAX1 U1115 ( .A(n2225), .B(n2193), .C(n2033), .YC(n1669), .YS(n1670) );
  FAX1 U1116 ( .A(n1676), .B(n1685), .C(n1674), .YC(n1671), .YS(n1672) );
  FAX1 U1117 ( .A(n1678), .B(n1680), .C(n1687), .YC(n1673), .YS(n1674) );
  FAX1 U1118 ( .A(n1682), .B(n1691), .C(n1689), .YC(n1675), .YS(n1676) );
  FAX1 U1119 ( .A(n2130), .B(n2034), .C(n2066), .YC(n1677), .YS(n1678) );
  FAX1 U1120 ( .A(n2098), .B(n2194), .C(n2162), .YC(n1679), .YS(n1680) );
  HAX1 U1121 ( .A(n2226), .B(n1752), .YC(n1681), .YS(n1682) );
  FAX1 U1122 ( .A(n1688), .B(n1695), .C(n1686), .YC(n1683), .YS(n1684) );
  FAX1 U1123 ( .A(n1692), .B(n1690), .C(n1697), .YC(n1685), .YS(n1686) );
  FAX1 U1124 ( .A(n2973), .B(n1701), .C(n1699), .YC(n1687), .YS(n1688) );
  FAX1 U1125 ( .A(n2163), .B(n2099), .C(n2131), .YC(n1689), .YS(n1690) );
  FAX1 U1126 ( .A(n2227), .B(n2195), .C(n2067), .YC(n1691), .YS(n1692) );
  FAX1 U1127 ( .A(n1698), .B(n1705), .C(n1696), .YC(n1693), .YS(n1694) );
  FAX1 U1128 ( .A(n1709), .B(n1700), .C(n1707), .YC(n1695), .YS(n1696) );
  FAX1 U1129 ( .A(n2164), .B(n2100), .C(n1702), .YC(n1697), .YS(n1698) );
  FAX1 U1130 ( .A(n2132), .B(n2068), .C(n2196), .YC(n1699), .YS(n1700) );
  HAX1 U1131 ( .A(n2228), .B(n1753), .YC(n1701), .YS(n1702) );
  FAX1 U1132 ( .A(n1708), .B(n1713), .C(n1706), .YC(n1703), .YS(n1704) );
  FAX1 U1133 ( .A(n1717), .B(n1715), .C(n1710), .YC(n1705), .YS(n1706) );
  FAX1 U1134 ( .A(n2165), .B(n2133), .C(n2938), .YC(n1707), .YS(n1708) );
  FAX1 U1135 ( .A(n2229), .B(n2197), .C(n2101), .YC(n1709), .YS(n1710) );
  FAX1 U1136 ( .A(n1716), .B(n1721), .C(n1714), .YC(n1711), .YS(n1712) );
  FAX1 U1137 ( .A(n2198), .B(n1718), .C(n1723), .YC(n1713), .YS(n1714) );
  FAX1 U1138 ( .A(n2134), .B(n2102), .C(n2166), .YC(n1715), .YS(n1716) );
  HAX1 U1139 ( .A(n2230), .B(n1754), .YC(n1717), .YS(n1718) );
  FAX1 U1140 ( .A(n1727), .B(n1724), .C(n1722), .YC(n1719), .YS(n1720) );
  FAX1 U1141 ( .A(n2167), .B(n2974), .C(n1729), .YC(n1721), .YS(n1722) );
  FAX1 U1142 ( .A(n2231), .B(n2199), .C(n2135), .YC(n1723), .YS(n1724) );
  FAX1 U1143 ( .A(n1730), .B(n1733), .C(n1728), .YC(n1725), .YS(n1726) );
  FAX1 U1144 ( .A(n2200), .B(n2136), .C(n2168), .YC(n1727), .YS(n1728) );
  HAX1 U1145 ( .A(n2232), .B(n1755), .YC(n1729), .YS(n1730) );
  FAX1 U1146 ( .A(n2976), .B(n1737), .C(n1734), .YC(n1731), .YS(n1732) );
  FAX1 U1147 ( .A(n2233), .B(n2201), .C(n2169), .YC(n1733), .YS(n1734) );
  FAX1 U1148 ( .A(n2202), .B(n2170), .C(n1738), .YC(n1735), .YS(n1736) );
  HAX1 U1149 ( .A(n2234), .B(n1756), .YC(n1737), .YS(n1738) );
  FAX1 U1150 ( .A(n2235), .B(n2203), .C(n2937), .YC(n1739), .YS(n1740) );
  HAX1 U1151 ( .A(n2236), .B(n2204), .YC(n1741), .YS(n1742) );
  NOR2X1 U1152 ( .A(n3001), .B(n2922), .Y(n1759) );
  NOR2X1 U1153 ( .A(n2240), .B(n2922), .Y(n918) );
  NOR2X1 U1154 ( .A(n3003), .B(n2922), .Y(n1760) );
  NOR2X1 U1155 ( .A(n2242), .B(n2922), .Y(n960) );
  NOR2X1 U1156 ( .A(n3006), .B(n2922), .Y(n1761) );
  NOR2X1 U1157 ( .A(n2244), .B(n2922), .Y(n1006) );
  NOR2X1 U1158 ( .A(n3009), .B(n2922), .Y(n1762) );
  NOR2X1 U1159 ( .A(n2246), .B(n2922), .Y(n1056) );
  NOR2X1 U1160 ( .A(n3012), .B(n2922), .Y(n1763) );
  NOR2X1 U1161 ( .A(n2248), .B(n2922), .Y(n1110) );
  NOR2X1 U1162 ( .A(n3014), .B(n2922), .Y(n1764) );
  NOR2X1 U1163 ( .A(n2250), .B(n2922), .Y(n1168) );
  NOR2X1 U1164 ( .A(n3016), .B(n2922), .Y(n1765) );
  NOR2X1 U1165 ( .A(n2252), .B(n2922), .Y(n1766) );
  NOR2X1 U1166 ( .A(n3018), .B(n2921), .Y(n1230) );
  INVX2 U1168 ( .A(n463), .Y(n2240) );
  INVX2 U1170 ( .A(n459), .Y(n2242) );
  INVX2 U1172 ( .A(n455), .Y(n2244) );
  INVX2 U1174 ( .A(n451), .Y(n2246) );
  INVX2 U1176 ( .A(n447), .Y(n2248) );
  INVX2 U1178 ( .A(n443), .Y(n2250) );
  INVX2 U1180 ( .A(n439), .Y(n2252) );
  OAI22X1 U1182 ( .A(n382), .B(n2272), .C(n2922), .D(n432), .Y(n1743) );
  OAI22X1 U1183 ( .A(n2254), .B(n381), .C(n2255), .D(n431), .Y(n1768) );
  OAI22X1 U1184 ( .A(n2255), .B(n381), .C(n2256), .D(n431), .Y(n1769) );
  OAI22X1 U1185 ( .A(n2256), .B(n381), .C(n2257), .D(n431), .Y(n1770) );
  OAI22X1 U1186 ( .A(n2257), .B(n381), .C(n2258), .D(n431), .Y(n1771) );
  OAI22X1 U1187 ( .A(n2258), .B(n381), .C(n2259), .D(n431), .Y(n1772) );
  OAI22X1 U1188 ( .A(n2259), .B(n381), .C(n2260), .D(n431), .Y(n1773) );
  OAI22X1 U1189 ( .A(n2260), .B(n380), .C(n2261), .D(n431), .Y(n1774) );
  OAI22X1 U1190 ( .A(n2261), .B(n380), .C(n2262), .D(n431), .Y(n1775) );
  OAI22X1 U1191 ( .A(n2262), .B(n380), .C(n2263), .D(n431), .Y(n1776) );
  OAI22X1 U1192 ( .A(n2263), .B(n380), .C(n2264), .D(n431), .Y(n1777) );
  OAI22X1 U1193 ( .A(n2264), .B(n380), .C(n2265), .D(n431), .Y(n1778) );
  OAI22X1 U1194 ( .A(n2265), .B(n380), .C(n2266), .D(n430), .Y(n1779) );
  OAI22X1 U1195 ( .A(n2266), .B(n380), .C(n2267), .D(n430), .Y(n1780) );
  OAI22X1 U1196 ( .A(n2267), .B(n380), .C(n2268), .D(n430), .Y(n1781) );
  OAI22X1 U1197 ( .A(n2268), .B(n380), .C(n2269), .D(n430), .Y(n1782) );
  OAI22X1 U1198 ( .A(n2269), .B(n380), .C(n2270), .D(n430), .Y(n1783) );
  OAI22X1 U1199 ( .A(n2270), .B(n380), .C(n2271), .D(n430), .Y(n1784) );
  XNOR2X1 U1200 ( .A(n333), .B(b[17]), .Y(n2254) );
  XNOR2X1 U1201 ( .A(n333), .B(n467), .Y(n2255) );
  XNOR2X1 U1202 ( .A(n333), .B(n3000), .Y(n2256) );
  XNOR2X1 U1203 ( .A(n333), .B(n463), .Y(n2257) );
  XNOR2X1 U1204 ( .A(n333), .B(n3002), .Y(n2258) );
  XNOR2X1 U1205 ( .A(n333), .B(n459), .Y(n2259) );
  XNOR2X1 U1206 ( .A(n333), .B(n3004), .Y(n2260) );
  XNOR2X1 U1207 ( .A(n333), .B(n455), .Y(n2261) );
  XNOR2X1 U1208 ( .A(n333), .B(n3007), .Y(n2262) );
  XNOR2X1 U1209 ( .A(n334), .B(n451), .Y(n2263) );
  XNOR2X1 U1210 ( .A(n334), .B(n3010), .Y(n2264) );
  XNOR2X1 U1211 ( .A(n84), .B(n447), .Y(n2265) );
  XNOR2X1 U1212 ( .A(n84), .B(n3013), .Y(n2266) );
  XNOR2X1 U1213 ( .A(n84), .B(n443), .Y(n2267) );
  XNOR2X1 U1214 ( .A(n84), .B(n3015), .Y(n2268) );
  XNOR2X1 U1215 ( .A(n84), .B(n439), .Y(n2269) );
  XNOR2X1 U1216 ( .A(n84), .B(n3017), .Y(n2270) );
  XNOR2X1 U1217 ( .A(n84), .B(n3020), .Y(n2271) );
  OAI22X1 U1218 ( .A(n379), .B(n2293), .C(n2797), .D(n429), .Y(n1744) );
  OAI22X1 U1219 ( .A(n2273), .B(n378), .C(n2274), .D(n428), .Y(n1786) );
  OAI22X1 U1220 ( .A(n2274), .B(n378), .C(n2275), .D(n428), .Y(n1787) );
  OAI22X1 U1221 ( .A(n2275), .B(n378), .C(n2276), .D(n428), .Y(n1788) );
  OAI22X1 U1222 ( .A(n2276), .B(n378), .C(n2277), .D(n428), .Y(n1789) );
  OAI22X1 U1223 ( .A(n2277), .B(n378), .C(n2278), .D(n428), .Y(n1790) );
  OAI22X1 U1224 ( .A(n2278), .B(n378), .C(n2279), .D(n428), .Y(n1791) );
  OAI22X1 U1225 ( .A(n2279), .B(n378), .C(n2280), .D(n428), .Y(n1792) );
  OAI22X1 U1226 ( .A(n2280), .B(n378), .C(n2281), .D(n428), .Y(n1793) );
  OAI22X1 U1227 ( .A(n2281), .B(n377), .C(n2282), .D(n428), .Y(n1794) );
  OAI22X1 U1228 ( .A(n2282), .B(n377), .C(n2283), .D(n427), .Y(n1795) );
  OAI22X1 U1229 ( .A(n2283), .B(n377), .C(n2284), .D(n427), .Y(n1796) );
  OAI22X1 U1230 ( .A(n2284), .B(n377), .C(n2285), .D(n427), .Y(n1797) );
  OAI22X1 U1231 ( .A(n2285), .B(n377), .C(n2286), .D(n427), .Y(n1798) );
  OAI22X1 U1232 ( .A(n2286), .B(n377), .C(n2287), .D(n427), .Y(n1799) );
  OAI22X1 U1233 ( .A(n2287), .B(n377), .C(n2288), .D(n427), .Y(n1800) );
  OAI22X1 U1234 ( .A(n2288), .B(n377), .C(n2289), .D(n427), .Y(n1801) );
  OAI22X1 U1235 ( .A(n2289), .B(n377), .C(n2290), .D(n427), .Y(n1802) );
  OAI22X1 U1236 ( .A(n2290), .B(n377), .C(n2291), .D(n427), .Y(n1803) );
  OAI22X1 U1237 ( .A(n2291), .B(n377), .C(n2292), .D(n427), .Y(n1804) );
  XNOR2X1 U1238 ( .A(n330), .B(b[19]), .Y(n2273) );
  XNOR2X1 U1239 ( .A(n330), .B(n471), .Y(n2274) );
  XNOR2X1 U1240 ( .A(n330), .B(b[17]), .Y(n2275) );
  XNOR2X1 U1241 ( .A(n330), .B(n467), .Y(n2276) );
  XNOR2X1 U1242 ( .A(n330), .B(n3000), .Y(n2277) );
  XNOR2X1 U1243 ( .A(n330), .B(n463), .Y(n2278) );
  XNOR2X1 U1244 ( .A(n330), .B(n3002), .Y(n2279) );
  XNOR2X1 U1245 ( .A(n330), .B(n459), .Y(n2280) );
  XNOR2X1 U1246 ( .A(n330), .B(n3004), .Y(n2281) );
  XNOR2X1 U1247 ( .A(n330), .B(n455), .Y(n2282) );
  XNOR2X1 U1248 ( .A(n330), .B(n3007), .Y(n2283) );
  XNOR2X1 U1249 ( .A(n329), .B(n451), .Y(n2284) );
  XNOR2X1 U1250 ( .A(n329), .B(n3010), .Y(n2285) );
  XNOR2X1 U1251 ( .A(n329), .B(n447), .Y(n2286) );
  XNOR2X1 U1252 ( .A(n329), .B(n3013), .Y(n2287) );
  XNOR2X1 U1253 ( .A(n329), .B(n443), .Y(n2288) );
  XNOR2X1 U1254 ( .A(n329), .B(n3015), .Y(n2289) );
  XNOR2X1 U1255 ( .A(n329), .B(n439), .Y(n2290) );
  XNOR2X1 U1256 ( .A(n329), .B(n3017), .Y(n2291) );
  XNOR2X1 U1257 ( .A(n329), .B(n3019), .Y(n2292) );
  OAI22X1 U1258 ( .A(n376), .B(n2316), .C(n2798), .D(n426), .Y(n1745) );
  OAI22X1 U1259 ( .A(n2294), .B(n375), .C(n2295), .D(n425), .Y(n1806) );
  OAI22X1 U1260 ( .A(n2295), .B(n375), .C(n2296), .D(n425), .Y(n1807) );
  OAI22X1 U1261 ( .A(n2296), .B(n375), .C(n2297), .D(n425), .Y(n1808) );
  OAI22X1 U1262 ( .A(n2297), .B(n375), .C(n2298), .D(n425), .Y(n1809) );
  OAI22X1 U1263 ( .A(n2298), .B(n375), .C(n2299), .D(n425), .Y(n1810) );
  OAI22X1 U1264 ( .A(n2299), .B(n375), .C(n2300), .D(n425), .Y(n1811) );
  OAI22X1 U1265 ( .A(n2300), .B(n375), .C(n2301), .D(n425), .Y(n1812) );
  OAI22X1 U1266 ( .A(n2301), .B(n375), .C(n2302), .D(n425), .Y(n1813) );
  OAI22X1 U1267 ( .A(n2302), .B(n375), .C(n2303), .D(n425), .Y(n1814) );
  OAI22X1 U1268 ( .A(n2303), .B(n375), .C(n2304), .D(n425), .Y(n1815) );
  OAI22X1 U1269 ( .A(n2304), .B(n2909), .C(n2305), .D(n425), .Y(n1816) );
  OAI22X1 U1270 ( .A(n2305), .B(n2909), .C(n2306), .D(n425), .Y(n1817) );
  OAI22X1 U1271 ( .A(n2306), .B(n2909), .C(n2307), .D(n425), .Y(n1818) );
  OAI22X1 U1272 ( .A(n2307), .B(n2909), .C(n2308), .D(n424), .Y(n1819) );
  OAI22X1 U1273 ( .A(n2308), .B(n2909), .C(n2309), .D(n424), .Y(n1820) );
  OAI22X1 U1274 ( .A(n2309), .B(n2909), .C(n2310), .D(n425), .Y(n1821) );
  OAI22X1 U1275 ( .A(n2310), .B(n2909), .C(n2311), .D(n425), .Y(n1822) );
  OAI22X1 U1276 ( .A(n2311), .B(n2909), .C(n2312), .D(n424), .Y(n1823) );
  OAI22X1 U1277 ( .A(n2312), .B(n2909), .C(n2313), .D(n424), .Y(n1824) );
  OAI22X1 U1278 ( .A(n2313), .B(n2909), .C(n2314), .D(n424), .Y(n1825) );
  OAI22X1 U1279 ( .A(n2314), .B(n2909), .C(n2315), .D(n424), .Y(n1826) );
  XNOR2X1 U1280 ( .A(n328), .B(n2994), .Y(n2294) );
  XNOR2X1 U1281 ( .A(n2982), .B(n475), .Y(n2295) );
  XNOR2X1 U1282 ( .A(n2983), .B(b[19]), .Y(n2296) );
  XNOR2X1 U1283 ( .A(n2982), .B(n471), .Y(n2297) );
  XNOR2X1 U1284 ( .A(n2983), .B(b[17]), .Y(n2298) );
  XNOR2X1 U1285 ( .A(n2982), .B(n467), .Y(n2299) );
  XNOR2X1 U1286 ( .A(n2983), .B(n3000), .Y(n2300) );
  XNOR2X1 U1287 ( .A(n2982), .B(n463), .Y(n2301) );
  XNOR2X1 U1288 ( .A(n2983), .B(n3002), .Y(n2302) );
  XNOR2X1 U1289 ( .A(n2983), .B(n459), .Y(n2303) );
  XNOR2X1 U1290 ( .A(n2982), .B(n3004), .Y(n2304) );
  XNOR2X1 U1291 ( .A(n2982), .B(n455), .Y(n2305) );
  XNOR2X1 U1292 ( .A(n2983), .B(n3007), .Y(n2306) );
  XNOR2X1 U1293 ( .A(n2981), .B(n451), .Y(n2307) );
  XNOR2X1 U1294 ( .A(n326), .B(n3010), .Y(n2308) );
  XNOR2X1 U1295 ( .A(n326), .B(n447), .Y(n2309) );
  XNOR2X1 U1296 ( .A(n2981), .B(n3013), .Y(n2310) );
  XNOR2X1 U1297 ( .A(n326), .B(n443), .Y(n2311) );
  XNOR2X1 U1298 ( .A(n326), .B(n3015), .Y(n2312) );
  XNOR2X1 U1299 ( .A(n326), .B(n439), .Y(n2313) );
  XNOR2X1 U1300 ( .A(n326), .B(n3017), .Y(n2314) );
  XNOR2X1 U1301 ( .A(n326), .B(n3020), .Y(n2315) );
  OAI22X1 U1302 ( .A(n373), .B(n2341), .C(n2799), .D(n423), .Y(n1746) );
  OAI22X1 U1303 ( .A(n2317), .B(n372), .C(n2318), .D(n423), .Y(n1828) );
  OAI22X1 U1304 ( .A(n2318), .B(n372), .C(n2319), .D(n422), .Y(n1829) );
  OAI22X1 U1305 ( .A(n2319), .B(n372), .C(n2320), .D(n422), .Y(n1830) );
  OAI22X1 U1306 ( .A(n2320), .B(n372), .C(n2321), .D(n422), .Y(n1831) );
  OAI22X1 U1307 ( .A(n2321), .B(n372), .C(n2322), .D(n422), .Y(n1832) );
  OAI22X1 U1308 ( .A(n2322), .B(n372), .C(n2323), .D(n422), .Y(n1833) );
  OAI22X1 U1309 ( .A(n2323), .B(n372), .C(n2324), .D(n422), .Y(n1834) );
  OAI22X1 U1310 ( .A(n2324), .B(n372), .C(n2325), .D(n422), .Y(n1835) );
  OAI22X1 U1311 ( .A(n2325), .B(n372), .C(n2326), .D(n422), .Y(n1836) );
  OAI22X1 U1312 ( .A(n2326), .B(n372), .C(n2327), .D(n422), .Y(n1837) );
  OAI22X1 U1313 ( .A(n2327), .B(n372), .C(n2328), .D(n422), .Y(n1838) );
  OAI22X1 U1314 ( .A(n2328), .B(n372), .C(n2329), .D(n422), .Y(n1839) );
  OAI22X1 U1315 ( .A(n2329), .B(n371), .C(n2330), .D(n422), .Y(n1840) );
  OAI22X1 U1316 ( .A(n2330), .B(n371), .C(n2331), .D(n421), .Y(n1841) );
  OAI22X1 U1317 ( .A(n2331), .B(n371), .C(n2332), .D(n421), .Y(n1842) );
  OAI22X1 U1318 ( .A(n2332), .B(n371), .C(n2333), .D(n421), .Y(n1843) );
  OAI22X1 U1319 ( .A(n2333), .B(n371), .C(n2334), .D(n421), .Y(n1844) );
  OAI22X1 U1320 ( .A(n2334), .B(n371), .C(n2335), .D(n421), .Y(n1845) );
  OAI22X1 U1321 ( .A(n2335), .B(n371), .C(n2336), .D(n421), .Y(n1846) );
  OAI22X1 U1322 ( .A(n2336), .B(n371), .C(n2337), .D(n421), .Y(n1847) );
  OAI22X1 U1323 ( .A(n2337), .B(n371), .C(n2338), .D(n421), .Y(n1848) );
  OAI22X1 U1324 ( .A(n2338), .B(n371), .C(n2339), .D(n421), .Y(n1849) );
  OAI22X1 U1325 ( .A(n2339), .B(n371), .C(n2340), .D(n421), .Y(n1850) );
  XNOR2X1 U1326 ( .A(n325), .B(n2991), .Y(n2317) );
  XNOR2X1 U1327 ( .A(n324), .B(n479), .Y(n2318) );
  XNOR2X1 U1328 ( .A(n2966), .B(n2994), .Y(n2319) );
  XNOR2X1 U1329 ( .A(n2967), .B(n475), .Y(n2320) );
  XNOR2X1 U1330 ( .A(n2967), .B(b[19]), .Y(n2321) );
  XNOR2X1 U1331 ( .A(n2966), .B(n471), .Y(n2322) );
  XNOR2X1 U1332 ( .A(n325), .B(b[17]), .Y(n2323) );
  XNOR2X1 U1333 ( .A(n324), .B(n467), .Y(n2324) );
  XNOR2X1 U1334 ( .A(n2966), .B(n3000), .Y(n2325) );
  XNOR2X1 U1335 ( .A(n324), .B(n463), .Y(n2326) );
  XNOR2X1 U1336 ( .A(n325), .B(n3002), .Y(n2327) );
  XNOR2X1 U1337 ( .A(n2967), .B(n459), .Y(n2328) );
  XNOR2X1 U1338 ( .A(n2966), .B(n3004), .Y(n2329) );
  XNOR2X1 U1339 ( .A(n324), .B(n455), .Y(n2330) );
  XNOR2X1 U1340 ( .A(n2966), .B(n3007), .Y(n2331) );
  XNOR2X1 U1341 ( .A(n2967), .B(n451), .Y(n2332) );
  XNOR2X1 U1342 ( .A(n325), .B(n3010), .Y(n2333) );
  XNOR2X1 U1343 ( .A(n325), .B(n447), .Y(n2334) );
  XNOR2X1 U1344 ( .A(n325), .B(n3013), .Y(n2335) );
  XNOR2X1 U1345 ( .A(n324), .B(n443), .Y(n2336) );
  XNOR2X1 U1346 ( .A(n2967), .B(n3015), .Y(n2337) );
  XNOR2X1 U1347 ( .A(n323), .B(n439), .Y(n2338) );
  XNOR2X1 U1348 ( .A(n323), .B(n3017), .Y(n2339) );
  XNOR2X1 U1349 ( .A(n323), .B(n3020), .Y(n2340) );
  OAI22X1 U1350 ( .A(n370), .B(n2368), .C(n2800), .D(n420), .Y(n1747) );
  OAI22X1 U1351 ( .A(n2342), .B(n370), .C(n2343), .D(n420), .Y(n1852) );
  OAI22X1 U1352 ( .A(n2343), .B(n370), .C(n2344), .D(n420), .Y(n1853) );
  OAI22X1 U1353 ( .A(n2344), .B(n369), .C(n2345), .D(n420), .Y(n1854) );
  OAI22X1 U1354 ( .A(n2345), .B(n369), .C(n2346), .D(n419), .Y(n1855) );
  OAI22X1 U1355 ( .A(n2346), .B(n369), .C(n2347), .D(n419), .Y(n1856) );
  OAI22X1 U1356 ( .A(n2347), .B(n369), .C(n2348), .D(n419), .Y(n1857) );
  OAI22X1 U1357 ( .A(n2348), .B(n369), .C(n2349), .D(n419), .Y(n1858) );
  OAI22X1 U1358 ( .A(n2349), .B(n369), .C(n2350), .D(n419), .Y(n1859) );
  OAI22X1 U1359 ( .A(n2350), .B(n369), .C(n2351), .D(n419), .Y(n1860) );
  OAI22X1 U1360 ( .A(n2351), .B(n369), .C(n2352), .D(n419), .Y(n1861) );
  OAI22X1 U1361 ( .A(n2352), .B(n369), .C(n2353), .D(n419), .Y(n1862) );
  OAI22X1 U1362 ( .A(n2353), .B(n369), .C(n2354), .D(n419), .Y(n1863) );
  OAI22X1 U1363 ( .A(n2354), .B(n369), .C(n2355), .D(n419), .Y(n1864) );
  OAI22X1 U1364 ( .A(n2355), .B(n369), .C(n2356), .D(n419), .Y(n1865) );
  OAI22X1 U1365 ( .A(n2356), .B(n368), .C(n2357), .D(n419), .Y(n1866) );
  OAI22X1 U1366 ( .A(n2357), .B(n368), .C(n2358), .D(n418), .Y(n1867) );
  OAI22X1 U1367 ( .A(n2358), .B(n368), .C(n2359), .D(n418), .Y(n1868) );
  OAI22X1 U1368 ( .A(n2359), .B(n368), .C(n2360), .D(n418), .Y(n1869) );
  OAI22X1 U1369 ( .A(n2360), .B(n368), .C(n2361), .D(n418), .Y(n1870) );
  OAI22X1 U1370 ( .A(n2361), .B(n368), .C(n2362), .D(n418), .Y(n1871) );
  OAI22X1 U1371 ( .A(n2362), .B(n368), .C(n2363), .D(n418), .Y(n1872) );
  OAI22X1 U1372 ( .A(n2363), .B(n368), .C(n2364), .D(n418), .Y(n1873) );
  OAI22X1 U1373 ( .A(n2364), .B(n368), .C(n2365), .D(n418), .Y(n1874) );
  OAI22X1 U1374 ( .A(n2365), .B(n368), .C(n2366), .D(n418), .Y(n1875) );
  OAI22X1 U1375 ( .A(n2366), .B(n368), .C(n2367), .D(n418), .Y(n1876) );
  XNOR2X1 U1376 ( .A(n322), .B(n2988), .Y(n2342) );
  XNOR2X1 U1377 ( .A(n322), .B(n483), .Y(n2343) );
  XNOR2X1 U1378 ( .A(n322), .B(n2990), .Y(n2344) );
  XNOR2X1 U1379 ( .A(n322), .B(n479), .Y(n2345) );
  XNOR2X1 U1380 ( .A(n322), .B(n2993), .Y(n2346) );
  XNOR2X1 U1381 ( .A(n2920), .B(n475), .Y(n2347) );
  XNOR2X1 U1382 ( .A(n2920), .B(n2996), .Y(n2348) );
  XNOR2X1 U1383 ( .A(n2920), .B(n471), .Y(n2349) );
  XNOR2X1 U1384 ( .A(n2920), .B(n2998), .Y(n2350) );
  XNOR2X1 U1385 ( .A(n2920), .B(n467), .Y(n2351) );
  XNOR2X1 U1386 ( .A(n2920), .B(n3000), .Y(n2352) );
  XNOR2X1 U1387 ( .A(n2920), .B(n463), .Y(n2353) );
  XNOR2X1 U1388 ( .A(n2920), .B(n3002), .Y(n2354) );
  XNOR2X1 U1389 ( .A(n2920), .B(n459), .Y(n2355) );
  XNOR2X1 U1390 ( .A(n2919), .B(n3004), .Y(n2356) );
  XNOR2X1 U1391 ( .A(n2919), .B(n455), .Y(n2357) );
  XNOR2X1 U1392 ( .A(n2919), .B(n3007), .Y(n2358) );
  XNOR2X1 U1393 ( .A(n320), .B(n451), .Y(n2359) );
  XNOR2X1 U1394 ( .A(n320), .B(n3010), .Y(n2360) );
  XNOR2X1 U1395 ( .A(n320), .B(n447), .Y(n2361) );
  XNOR2X1 U1396 ( .A(n320), .B(n3013), .Y(n2362) );
  XNOR2X1 U1397 ( .A(n320), .B(n443), .Y(n2363) );
  XNOR2X1 U1398 ( .A(n320), .B(n3015), .Y(n2364) );
  XNOR2X1 U1399 ( .A(n320), .B(n439), .Y(n2365) );
  XNOR2X1 U1400 ( .A(n320), .B(n3017), .Y(n2366) );
  XNOR2X1 U1401 ( .A(n320), .B(n3020), .Y(n2367) );
  OAI22X1 U1402 ( .A(n367), .B(n2397), .C(n2801), .D(n417), .Y(n1748) );
  OAI22X1 U1403 ( .A(n2369), .B(n367), .C(n2370), .D(n417), .Y(n1878) );
  OAI22X1 U1404 ( .A(n2370), .B(n367), .C(n2371), .D(n417), .Y(n1879) );
  OAI22X1 U1405 ( .A(n2371), .B(n367), .C(n2372), .D(n417), .Y(n1880) );
  OAI22X1 U1406 ( .A(n2372), .B(n367), .C(n2373), .D(n417), .Y(n1881) );
  OAI22X1 U1407 ( .A(n2373), .B(n366), .C(n2374), .D(n417), .Y(n1882) );
  OAI22X1 U1408 ( .A(n2374), .B(n366), .C(n2375), .D(n416), .Y(n1883) );
  OAI22X1 U1409 ( .A(n2375), .B(n366), .C(n2376), .D(n416), .Y(n1884) );
  OAI22X1 U1410 ( .A(n2376), .B(n366), .C(n2377), .D(n416), .Y(n1885) );
  OAI22X1 U1411 ( .A(n2377), .B(n366), .C(n2378), .D(n416), .Y(n1886) );
  OAI22X1 U1412 ( .A(n2378), .B(n366), .C(n2379), .D(n416), .Y(n1887) );
  OAI22X1 U1413 ( .A(n2379), .B(n366), .C(n2380), .D(n416), .Y(n1888) );
  OAI22X1 U1414 ( .A(n2380), .B(n366), .C(n2381), .D(n416), .Y(n1889) );
  OAI22X1 U1415 ( .A(n2381), .B(n366), .C(n2382), .D(n416), .Y(n1890) );
  OAI22X1 U1416 ( .A(n2382), .B(n366), .C(n2383), .D(n416), .Y(n1891) );
  OAI22X1 U1417 ( .A(n2383), .B(n366), .C(n2384), .D(n416), .Y(n1892) );
  OAI22X1 U1418 ( .A(n2384), .B(n366), .C(n2385), .D(n416), .Y(n1893) );
  OAI22X1 U1419 ( .A(n2385), .B(n365), .C(n2386), .D(n416), .Y(n1894) );
  OAI22X1 U1420 ( .A(n2386), .B(n365), .C(n2387), .D(n415), .Y(n1895) );
  OAI22X1 U1421 ( .A(n2387), .B(n365), .C(n2388), .D(n415), .Y(n1896) );
  OAI22X1 U1422 ( .A(n2388), .B(n365), .C(n2389), .D(n415), .Y(n1897) );
  OAI22X1 U1423 ( .A(n2389), .B(n365), .C(n2390), .D(n415), .Y(n1898) );
  OAI22X1 U1424 ( .A(n2390), .B(n365), .C(n2391), .D(n415), .Y(n1899) );
  OAI22X1 U1425 ( .A(n2391), .B(n365), .C(n2392), .D(n415), .Y(n1900) );
  OAI22X1 U1426 ( .A(n2392), .B(n365), .C(n2393), .D(n415), .Y(n1901) );
  OAI22X1 U1427 ( .A(n2393), .B(n365), .C(n2394), .D(n415), .Y(n1902) );
  OAI22X1 U1428 ( .A(n2394), .B(n365), .C(n2395), .D(n415), .Y(n1903) );
  OAI22X1 U1429 ( .A(n2395), .B(n365), .C(n2396), .D(n415), .Y(n1904) );
  XNOR2X1 U1430 ( .A(n319), .B(n2986), .Y(n2369) );
  XNOR2X1 U1431 ( .A(n319), .B(b[26]), .Y(n2370) );
  XNOR2X1 U1432 ( .A(n319), .B(n2988), .Y(n2371) );
  XNOR2X1 U1433 ( .A(n319), .B(n483), .Y(n2372) );
  XNOR2X1 U1434 ( .A(n319), .B(n2990), .Y(n2373) );
  XNOR2X1 U1435 ( .A(n319), .B(n479), .Y(n2374) );
  XNOR2X1 U1436 ( .A(n319), .B(n2993), .Y(n2375) );
  XNOR2X1 U1437 ( .A(n2918), .B(n475), .Y(n2376) );
  XNOR2X1 U1438 ( .A(n2918), .B(n2996), .Y(n2377) );
  XNOR2X1 U1439 ( .A(n2918), .B(n471), .Y(n2378) );
  XNOR2X1 U1440 ( .A(n2918), .B(n2998), .Y(n2379) );
  XNOR2X1 U1441 ( .A(n2918), .B(n467), .Y(n2380) );
  XNOR2X1 U1442 ( .A(n2918), .B(n3000), .Y(n2381) );
  XNOR2X1 U1443 ( .A(n2918), .B(n463), .Y(n2382) );
  XNOR2X1 U1444 ( .A(n2918), .B(n3002), .Y(n2383) );
  XNOR2X1 U1445 ( .A(n2918), .B(n459), .Y(n2384) );
  XNOR2X1 U1446 ( .A(n2918), .B(n3004), .Y(n2385) );
  XNOR2X1 U1447 ( .A(n2918), .B(n455), .Y(n2386) );
  XNOR2X1 U1448 ( .A(n2918), .B(n3007), .Y(n2387) );
  XNOR2X1 U1449 ( .A(n317), .B(n451), .Y(n2388) );
  XNOR2X1 U1450 ( .A(n317), .B(n3010), .Y(n2389) );
  XNOR2X1 U1451 ( .A(n317), .B(n447), .Y(n2390) );
  XNOR2X1 U1452 ( .A(n317), .B(n3013), .Y(n2391) );
  XNOR2X1 U1453 ( .A(n317), .B(n443), .Y(n2392) );
  XNOR2X1 U1454 ( .A(n317), .B(n3015), .Y(n2393) );
  XNOR2X1 U1455 ( .A(n317), .B(n439), .Y(n2394) );
  XNOR2X1 U1456 ( .A(n317), .B(n3017), .Y(n2395) );
  XNOR2X1 U1457 ( .A(n317), .B(n3019), .Y(n2396) );
  OAI22X1 U1458 ( .A(n364), .B(n2428), .C(n2802), .D(n414), .Y(n1749) );
  OAI22X1 U1459 ( .A(n2398), .B(n364), .C(n2399), .D(n414), .Y(n1906) );
  OAI22X1 U1460 ( .A(n2399), .B(n364), .C(n2400), .D(n414), .Y(n1907) );
  OAI22X1 U1461 ( .A(n2400), .B(n364), .C(n2401), .D(n414), .Y(n1908) );
  OAI22X1 U1462 ( .A(n2401), .B(n364), .C(n2402), .D(n414), .Y(n1909) );
  OAI22X1 U1463 ( .A(n2402), .B(n364), .C(n2403), .D(n414), .Y(n1910) );
  OAI22X1 U1464 ( .A(n2403), .B(n364), .C(n2404), .D(n414), .Y(n1911) );
  OAI22X1 U1465 ( .A(n2404), .B(n363), .C(n2405), .D(n414), .Y(n1912) );
  OAI22X1 U1466 ( .A(n2405), .B(n363), .C(n2406), .D(n413), .Y(n1913) );
  OAI22X1 U1467 ( .A(n2406), .B(n363), .C(n2407), .D(n413), .Y(n1914) );
  OAI22X1 U1468 ( .A(n2407), .B(n363), .C(n2408), .D(n413), .Y(n1915) );
  OAI22X1 U1469 ( .A(n2408), .B(n363), .C(n2409), .D(n413), .Y(n1916) );
  OAI22X1 U1470 ( .A(n2409), .B(n363), .C(n2410), .D(n413), .Y(n1917) );
  OAI22X1 U1471 ( .A(n2410), .B(n363), .C(n2411), .D(n413), .Y(n1918) );
  OAI22X1 U1472 ( .A(n2411), .B(n363), .C(n2412), .D(n413), .Y(n1919) );
  OAI22X1 U1473 ( .A(n2412), .B(n363), .C(n2413), .D(n413), .Y(n1920) );
  OAI22X1 U1474 ( .A(n2413), .B(n363), .C(n2414), .D(n413), .Y(n1921) );
  OAI22X1 U1475 ( .A(n2414), .B(n363), .C(n2415), .D(n413), .Y(n1922) );
  OAI22X1 U1476 ( .A(n2415), .B(n363), .C(n2416), .D(n413), .Y(n1923) );
  OAI22X1 U1477 ( .A(n2416), .B(n362), .C(n2417), .D(n413), .Y(n1924) );
  OAI22X1 U1478 ( .A(n2417), .B(n362), .C(n2418), .D(n412), .Y(n1925) );
  OAI22X1 U1479 ( .A(n2418), .B(n362), .C(n2419), .D(n412), .Y(n1926) );
  OAI22X1 U1480 ( .A(n2419), .B(n362), .C(n2420), .D(n412), .Y(n1927) );
  OAI22X1 U1481 ( .A(n2420), .B(n362), .C(n2421), .D(n412), .Y(n1928) );
  OAI22X1 U1482 ( .A(n2421), .B(n362), .C(n2422), .D(n412), .Y(n1929) );
  OAI22X1 U1483 ( .A(n2422), .B(n362), .C(n2423), .D(n412), .Y(n1930) );
  OAI22X1 U1484 ( .A(n2423), .B(n362), .C(n2424), .D(n412), .Y(n1931) );
  OAI22X1 U1485 ( .A(n2424), .B(n362), .C(n2425), .D(n412), .Y(n1932) );
  OAI22X1 U1486 ( .A(n2425), .B(n362), .C(n2426), .D(n412), .Y(n1933) );
  OAI22X1 U1487 ( .A(n2426), .B(n362), .C(n2427), .D(n412), .Y(n1934) );
  XNOR2X1 U1488 ( .A(n316), .B(b[29]), .Y(n2398) );
  XNOR2X1 U1489 ( .A(n316), .B(b[28]), .Y(n2399) );
  XNOR2X1 U1490 ( .A(n316), .B(n2986), .Y(n2400) );
  XNOR2X1 U1491 ( .A(n316), .B(b[26]), .Y(n2401) );
  XNOR2X1 U1492 ( .A(n316), .B(n2988), .Y(n2402) );
  XNOR2X1 U1493 ( .A(n316), .B(n483), .Y(n2403) );
  XNOR2X1 U1494 ( .A(n316), .B(n2990), .Y(n2404) );
  XNOR2X1 U1495 ( .A(n316), .B(n479), .Y(n2405) );
  XNOR2X1 U1496 ( .A(n316), .B(n2993), .Y(n2406) );
  XNOR2X1 U1497 ( .A(n315), .B(n475), .Y(n2407) );
  XNOR2X1 U1498 ( .A(n315), .B(n2996), .Y(n2408) );
  XNOR2X1 U1499 ( .A(n315), .B(n471), .Y(n2409) );
  XNOR2X1 U1500 ( .A(n315), .B(n2998), .Y(n2410) );
  XNOR2X1 U1501 ( .A(n315), .B(n467), .Y(n2411) );
  XNOR2X1 U1502 ( .A(n315), .B(n3000), .Y(n2412) );
  XNOR2X1 U1503 ( .A(n315), .B(n463), .Y(n2413) );
  XNOR2X1 U1504 ( .A(n315), .B(n3002), .Y(n2414) );
  XNOR2X1 U1505 ( .A(n315), .B(n459), .Y(n2415) );
  XNOR2X1 U1506 ( .A(n315), .B(n3004), .Y(n2416) );
  XNOR2X1 U1507 ( .A(n315), .B(n455), .Y(n2417) );
  XNOR2X1 U1508 ( .A(n315), .B(n3007), .Y(n2418) );
  XNOR2X1 U1509 ( .A(n314), .B(n451), .Y(n2419) );
  XNOR2X1 U1510 ( .A(n314), .B(n3010), .Y(n2420) );
  XNOR2X1 U1511 ( .A(n314), .B(n447), .Y(n2421) );
  XNOR2X1 U1512 ( .A(n314), .B(n3013), .Y(n2422) );
  XNOR2X1 U1513 ( .A(n314), .B(n443), .Y(n2423) );
  XNOR2X1 U1514 ( .A(n314), .B(n3015), .Y(n2424) );
  XNOR2X1 U1515 ( .A(n314), .B(n439), .Y(n2425) );
  XNOR2X1 U1516 ( .A(n314), .B(n3017), .Y(n2426) );
  XNOR2X1 U1517 ( .A(n314), .B(n3019), .Y(n2427) );
  OAI22X1 U1518 ( .A(n361), .B(n2461), .C(n2803), .D(n411), .Y(n1750) );
  OAI22X1 U1519 ( .A(n2429), .B(n361), .C(n2430), .D(n411), .Y(n1936) );
  OAI22X1 U1520 ( .A(n2430), .B(n361), .C(n2431), .D(n411), .Y(n1937) );
  OAI22X1 U1521 ( .A(n2431), .B(n361), .C(n2432), .D(n411), .Y(n1938) );
  OAI22X1 U1522 ( .A(n2432), .B(n361), .C(n2433), .D(n411), .Y(n1939) );
  OAI22X1 U1523 ( .A(n2433), .B(n361), .C(n2434), .D(n411), .Y(n1940) );
  OAI22X1 U1524 ( .A(n2434), .B(n361), .C(n2435), .D(n411), .Y(n1941) );
  OAI22X1 U1525 ( .A(n2435), .B(n361), .C(n2436), .D(n411), .Y(n1942) );
  OAI22X1 U1526 ( .A(n2436), .B(n361), .C(n2437), .D(n411), .Y(n1943) );
  OAI22X1 U1527 ( .A(n2437), .B(n360), .C(n2438), .D(n411), .Y(n1944) );
  OAI22X1 U1528 ( .A(n2438), .B(n360), .C(n2439), .D(n410), .Y(n1945) );
  OAI22X1 U1529 ( .A(n2439), .B(n360), .C(n2440), .D(n410), .Y(n1946) );
  OAI22X1 U1530 ( .A(n2440), .B(n360), .C(n2441), .D(n410), .Y(n1947) );
  OAI22X1 U1531 ( .A(n2441), .B(n360), .C(n2442), .D(n410), .Y(n1948) );
  OAI22X1 U1532 ( .A(n2442), .B(n360), .C(n2443), .D(n410), .Y(n1949) );
  OAI22X1 U1533 ( .A(n2443), .B(n360), .C(n2444), .D(n410), .Y(n1950) );
  OAI22X1 U1534 ( .A(n2444), .B(n360), .C(n2445), .D(n410), .Y(n1951) );
  OAI22X1 U1535 ( .A(n2445), .B(n360), .C(n2446), .D(n410), .Y(n1952) );
  OAI22X1 U1536 ( .A(n2446), .B(n360), .C(n2447), .D(n410), .Y(n1953) );
  OAI22X1 U1537 ( .A(n2447), .B(n360), .C(n2448), .D(n410), .Y(n1954) );
  OAI22X1 U1538 ( .A(n2448), .B(n360), .C(n2449), .D(n410), .Y(n1955) );
  OAI22X1 U1539 ( .A(n2449), .B(n359), .C(n2450), .D(n410), .Y(n1956) );
  OAI22X1 U1540 ( .A(n2450), .B(n359), .C(n2451), .D(n409), .Y(n1957) );
  OAI22X1 U1541 ( .A(n2451), .B(n359), .C(n2452), .D(n409), .Y(n1958) );
  OAI22X1 U1542 ( .A(n2452), .B(n359), .C(n2453), .D(n409), .Y(n1959) );
  OAI22X1 U1543 ( .A(n2453), .B(n359), .C(n2454), .D(n409), .Y(n1960) );
  OAI22X1 U1544 ( .A(n2454), .B(n359), .C(n2455), .D(n409), .Y(n1961) );
  OAI22X1 U1545 ( .A(n2455), .B(n359), .C(n2456), .D(n409), .Y(n1962) );
  OAI22X1 U1546 ( .A(n2456), .B(n359), .C(n2457), .D(n409), .Y(n1963) );
  OAI22X1 U1547 ( .A(n2457), .B(n359), .C(n2458), .D(n409), .Y(n1964) );
  OAI22X1 U1548 ( .A(n2458), .B(n359), .C(n2459), .D(n409), .Y(n1965) );
  OAI22X1 U1549 ( .A(n2459), .B(n359), .C(n2460), .D(n409), .Y(n1966) );
  XNOR2X1 U1550 ( .A(n2964), .B(n2984), .Y(n2429) );
  XNOR2X1 U1551 ( .A(n2965), .B(b[30]), .Y(n2430) );
  XNOR2X1 U1552 ( .A(n313), .B(b[29]), .Y(n2431) );
  XNOR2X1 U1553 ( .A(n312), .B(b[28]), .Y(n2432) );
  XNOR2X1 U1554 ( .A(n312), .B(n2986), .Y(n2433) );
  XNOR2X1 U1555 ( .A(n313), .B(b[26]), .Y(n2434) );
  XNOR2X1 U1556 ( .A(n2965), .B(n2988), .Y(n2435) );
  XNOR2X1 U1557 ( .A(n2964), .B(n483), .Y(n2436) );
  XNOR2X1 U1558 ( .A(n2964), .B(n2990), .Y(n2437) );
  XNOR2X1 U1559 ( .A(n2965), .B(n479), .Y(n2438) );
  XNOR2X1 U1560 ( .A(n313), .B(n2993), .Y(n2439) );
  XNOR2X1 U1561 ( .A(n2964), .B(n475), .Y(n2440) );
  XNOR2X1 U1562 ( .A(n312), .B(n2996), .Y(n2441) );
  XNOR2X1 U1563 ( .A(n2965), .B(n471), .Y(n2442) );
  XNOR2X1 U1564 ( .A(n2965), .B(n2998), .Y(n2443) );
  XNOR2X1 U1565 ( .A(n313), .B(n467), .Y(n2444) );
  XNOR2X1 U1566 ( .A(n312), .B(n3000), .Y(n2445) );
  XNOR2X1 U1567 ( .A(n2964), .B(n463), .Y(n2446) );
  XNOR2X1 U1568 ( .A(n312), .B(n3002), .Y(n2447) );
  XNOR2X1 U1569 ( .A(n313), .B(n459), .Y(n2448) );
  XNOR2X1 U1570 ( .A(n2964), .B(n3004), .Y(n2449) );
  XNOR2X1 U1571 ( .A(n2965), .B(n455), .Y(n2450) );
  XNOR2X1 U1572 ( .A(n2965), .B(n3007), .Y(n2451) );
  XNOR2X1 U1573 ( .A(n2964), .B(n451), .Y(n2452) );
  XNOR2X1 U1574 ( .A(n312), .B(n3010), .Y(n2453) );
  XNOR2X1 U1575 ( .A(n313), .B(n447), .Y(n2454) );
  XNOR2X1 U1576 ( .A(n2964), .B(n3013), .Y(n2455) );
  XNOR2X1 U1577 ( .A(n312), .B(n443), .Y(n2456) );
  XNOR2X1 U1578 ( .A(n313), .B(n3015), .Y(n2457) );
  XNOR2X1 U1579 ( .A(n311), .B(n439), .Y(n2458) );
  XNOR2X1 U1580 ( .A(n311), .B(n3017), .Y(n2459) );
  XNOR2X1 U1581 ( .A(n311), .B(n3019), .Y(n2460) );
  OAI22X1 U1582 ( .A(n358), .B(n2494), .C(n2804), .D(n408), .Y(n1751) );
  OAI22X1 U1583 ( .A(n2804), .B(n358), .C(n2462), .D(n408), .Y(n1969) );
  OAI22X1 U1584 ( .A(n2462), .B(n358), .C(n2463), .D(n408), .Y(n1970) );
  OAI22X1 U1585 ( .A(n2463), .B(n358), .C(n2464), .D(n408), .Y(n1971) );
  OAI22X1 U1586 ( .A(n2464), .B(n358), .C(n2465), .D(n408), .Y(n1972) );
  OAI22X1 U1587 ( .A(n2465), .B(n358), .C(n2466), .D(n408), .Y(n1973) );
  OAI22X1 U1588 ( .A(n2466), .B(n358), .C(n2467), .D(n408), .Y(n1974) );
  OAI22X1 U1589 ( .A(n2467), .B(n358), .C(n2468), .D(n408), .Y(n1975) );
  OAI22X1 U1590 ( .A(n2468), .B(n358), .C(n2469), .D(n408), .Y(n1976) );
  OAI22X1 U1591 ( .A(n2469), .B(n358), .C(n2470), .D(n408), .Y(n1977) );
  OAI22X1 U1592 ( .A(n2470), .B(n357), .C(n2471), .D(n408), .Y(n1978) );
  OAI22X1 U1593 ( .A(n2471), .B(n357), .C(n2472), .D(n407), .Y(n1979) );
  OAI22X1 U1594 ( .A(n2472), .B(n357), .C(n2473), .D(n407), .Y(n1980) );
  OAI22X1 U1595 ( .A(n2473), .B(n357), .C(n2474), .D(n407), .Y(n1981) );
  OAI22X1 U1596 ( .A(n2474), .B(n357), .C(n2475), .D(n407), .Y(n1982) );
  OAI22X1 U1597 ( .A(n2475), .B(n357), .C(n2476), .D(n407), .Y(n1983) );
  OAI22X1 U1598 ( .A(n2476), .B(n357), .C(n2477), .D(n407), .Y(n1984) );
  OAI22X1 U1599 ( .A(n2477), .B(n357), .C(n2478), .D(n407), .Y(n1985) );
  OAI22X1 U1600 ( .A(n2478), .B(n357), .C(n2479), .D(n407), .Y(n1986) );
  OAI22X1 U1601 ( .A(n2479), .B(n357), .C(n2480), .D(n407), .Y(n1987) );
  OAI22X1 U1602 ( .A(n2480), .B(n357), .C(n2481), .D(n407), .Y(n1988) );
  OAI22X1 U1603 ( .A(n2481), .B(n357), .C(n2482), .D(n407), .Y(n1989) );
  OAI22X1 U1604 ( .A(n2482), .B(n356), .C(n2483), .D(n407), .Y(n1990) );
  OAI22X1 U1605 ( .A(n2483), .B(n356), .C(n2484), .D(n406), .Y(n1991) );
  OAI22X1 U1606 ( .A(n2484), .B(n356), .C(n2485), .D(n406), .Y(n1992) );
  OAI22X1 U1607 ( .A(n2485), .B(n356), .C(n2486), .D(n406), .Y(n1993) );
  OAI22X1 U1608 ( .A(n2486), .B(n356), .C(n2487), .D(n406), .Y(n1994) );
  OAI22X1 U1609 ( .A(n2487), .B(n356), .C(n2488), .D(n406), .Y(n1995) );
  OAI22X1 U1610 ( .A(n2488), .B(n356), .C(n2489), .D(n406), .Y(n1996) );
  OAI22X1 U1611 ( .A(n2489), .B(n356), .C(n2490), .D(n406), .Y(n1997) );
  OAI22X1 U1612 ( .A(n2490), .B(n356), .C(n2491), .D(n406), .Y(n1998) );
  OAI22X1 U1613 ( .A(n2491), .B(n356), .C(n2492), .D(n406), .Y(n1999) );
  OAI22X1 U1614 ( .A(n2492), .B(n356), .C(n2493), .D(n406), .Y(n2000) );
  XNOR2X1 U1615 ( .A(n310), .B(n2984), .Y(n2462) );
  XNOR2X1 U1616 ( .A(n310), .B(n495), .Y(n2463) );
  XNOR2X1 U1617 ( .A(n310), .B(b[29]), .Y(n2464) );
  XNOR2X1 U1618 ( .A(n310), .B(n491), .Y(n2465) );
  XNOR2X1 U1619 ( .A(n310), .B(n2986), .Y(n2466) );
  XNOR2X1 U1620 ( .A(n310), .B(n487), .Y(n2467) );
  XNOR2X1 U1621 ( .A(n310), .B(n2988), .Y(n2468) );
  XNOR2X1 U1622 ( .A(n310), .B(n483), .Y(n2469) );
  XNOR2X1 U1623 ( .A(n310), .B(n2990), .Y(n2470) );
  XNOR2X1 U1624 ( .A(n310), .B(n479), .Y(n2471) );
  XNOR2X1 U1625 ( .A(n310), .B(n2993), .Y(n2472) );
  XNOR2X1 U1626 ( .A(n309), .B(n475), .Y(n2473) );
  XNOR2X1 U1627 ( .A(n309), .B(n2996), .Y(n2474) );
  XNOR2X1 U1628 ( .A(n309), .B(n471), .Y(n2475) );
  XNOR2X1 U1629 ( .A(n309), .B(n2998), .Y(n2476) );
  XNOR2X1 U1630 ( .A(n309), .B(n467), .Y(n2477) );
  XNOR2X1 U1631 ( .A(n309), .B(b[15]), .Y(n2478) );
  XNOR2X1 U1632 ( .A(n309), .B(n463), .Y(n2479) );
  XNOR2X1 U1633 ( .A(n309), .B(b[13]), .Y(n2480) );
  XNOR2X1 U1634 ( .A(n309), .B(n459), .Y(n2481) );
  XNOR2X1 U1635 ( .A(n309), .B(n3005), .Y(n2482) );
  XNOR2X1 U1636 ( .A(n309), .B(n455), .Y(n2483) );
  XNOR2X1 U1637 ( .A(n309), .B(n3008), .Y(n2484) );
  XNOR2X1 U1638 ( .A(n2911), .B(n451), .Y(n2485) );
  XNOR2X1 U1639 ( .A(n2911), .B(n3011), .Y(n2486) );
  XNOR2X1 U1640 ( .A(n2911), .B(n447), .Y(n2487) );
  XNOR2X1 U1641 ( .A(n2911), .B(b[5]), .Y(n2488) );
  XNOR2X1 U1642 ( .A(n2911), .B(n443), .Y(n2489) );
  XNOR2X1 U1643 ( .A(n2910), .B(b[3]), .Y(n2490) );
  XNOR2X1 U1644 ( .A(n2910), .B(n439), .Y(n2491) );
  XNOR2X1 U1645 ( .A(n2910), .B(b[1]), .Y(n2492) );
  XNOR2X1 U1646 ( .A(n2911), .B(n3019), .Y(n2493) );
  OAI22X1 U1647 ( .A(n355), .B(n2527), .C(n2805), .D(n405), .Y(n1752) );
  OAI22X1 U1648 ( .A(n2805), .B(n355), .C(n2495), .D(n405), .Y(n2003) );
  OAI22X1 U1649 ( .A(n2495), .B(n355), .C(n2496), .D(n405), .Y(n2004) );
  OAI22X1 U1650 ( .A(n2496), .B(n355), .C(n2497), .D(n405), .Y(n2005) );
  OAI22X1 U1651 ( .A(n2497), .B(n355), .C(n2498), .D(n405), .Y(n2006) );
  OAI22X1 U1652 ( .A(n2498), .B(n355), .C(n2499), .D(n405), .Y(n2007) );
  OAI22X1 U1653 ( .A(n2499), .B(n355), .C(n2500), .D(n405), .Y(n2008) );
  OAI22X1 U1654 ( .A(n2500), .B(n355), .C(n2501), .D(n405), .Y(n2009) );
  OAI22X1 U1655 ( .A(n2501), .B(n355), .C(n2502), .D(n405), .Y(n2010) );
  OAI22X1 U1656 ( .A(n2502), .B(n355), .C(n2503), .D(n405), .Y(n2011) );
  OAI22X1 U1657 ( .A(n2503), .B(n354), .C(n2504), .D(n405), .Y(n2012) );
  OAI22X1 U1658 ( .A(n2504), .B(n354), .C(n2505), .D(n404), .Y(n2013) );
  OAI22X1 U1659 ( .A(n2505), .B(n354), .C(n2506), .D(n404), .Y(n2014) );
  OAI22X1 U1660 ( .A(n2506), .B(n354), .C(n2507), .D(n404), .Y(n2015) );
  OAI22X1 U1661 ( .A(n2507), .B(n354), .C(n2508), .D(n404), .Y(n2016) );
  OAI22X1 U1662 ( .A(n2508), .B(n354), .C(n2509), .D(n404), .Y(n2017) );
  OAI22X1 U1663 ( .A(n2509), .B(n354), .C(n2510), .D(n404), .Y(n2018) );
  OAI22X1 U1664 ( .A(n2510), .B(n354), .C(n2511), .D(n404), .Y(n2019) );
  OAI22X1 U1665 ( .A(n2511), .B(n354), .C(n2512), .D(n404), .Y(n2020) );
  OAI22X1 U1666 ( .A(n2512), .B(n354), .C(n2513), .D(n404), .Y(n2021) );
  OAI22X1 U1667 ( .A(n2513), .B(n354), .C(n2514), .D(n404), .Y(n2022) );
  OAI22X1 U1668 ( .A(n2514), .B(n354), .C(n2515), .D(n404), .Y(n2023) );
  OAI22X1 U1669 ( .A(n2515), .B(n353), .C(n2516), .D(n404), .Y(n2024) );
  OAI22X1 U1670 ( .A(n2516), .B(n353), .C(n2517), .D(n403), .Y(n2025) );
  OAI22X1 U1671 ( .A(n2517), .B(n353), .C(n2518), .D(n403), .Y(n2026) );
  OAI22X1 U1672 ( .A(n2518), .B(n353), .C(n2519), .D(n403), .Y(n2027) );
  OAI22X1 U1673 ( .A(n2519), .B(n353), .C(n2520), .D(n403), .Y(n2028) );
  OAI22X1 U1674 ( .A(n2520), .B(n353), .C(n2521), .D(n403), .Y(n2029) );
  OAI22X1 U1675 ( .A(n2521), .B(n353), .C(n2522), .D(n403), .Y(n2030) );
  OAI22X1 U1676 ( .A(n2522), .B(n353), .C(n2523), .D(n403), .Y(n2031) );
  OAI22X1 U1677 ( .A(n2523), .B(n353), .C(n2524), .D(n403), .Y(n2032) );
  OAI22X1 U1678 ( .A(n2524), .B(n353), .C(n2525), .D(n403), .Y(n2033) );
  OAI22X1 U1679 ( .A(n2525), .B(n353), .C(n2526), .D(n403), .Y(n2034) );
  XNOR2X1 U1680 ( .A(n307), .B(n2984), .Y(n2495) );
  XNOR2X1 U1681 ( .A(n307), .B(n495), .Y(n2496) );
  XNOR2X1 U1682 ( .A(n307), .B(b[29]), .Y(n2497) );
  XNOR2X1 U1683 ( .A(n307), .B(n491), .Y(n2498) );
  XNOR2X1 U1684 ( .A(n307), .B(n2986), .Y(n2499) );
  XNOR2X1 U1685 ( .A(n307), .B(n487), .Y(n2500) );
  XNOR2X1 U1686 ( .A(n307), .B(n2988), .Y(n2501) );
  XNOR2X1 U1687 ( .A(n307), .B(n483), .Y(n2502) );
  XNOR2X1 U1688 ( .A(n307), .B(n2990), .Y(n2503) );
  XNOR2X1 U1689 ( .A(n307), .B(n479), .Y(n2504) );
  XNOR2X1 U1690 ( .A(n307), .B(n2993), .Y(n2505) );
  XNOR2X1 U1691 ( .A(n306), .B(n475), .Y(n2506) );
  XNOR2X1 U1692 ( .A(n306), .B(n2996), .Y(n2507) );
  XNOR2X1 U1693 ( .A(n306), .B(n471), .Y(n2508) );
  XNOR2X1 U1694 ( .A(n306), .B(n2998), .Y(n2509) );
  XNOR2X1 U1695 ( .A(n306), .B(n467), .Y(n2510) );
  XNOR2X1 U1696 ( .A(n306), .B(b[15]), .Y(n2511) );
  XNOR2X1 U1697 ( .A(n306), .B(n463), .Y(n2512) );
  XNOR2X1 U1698 ( .A(n306), .B(b[13]), .Y(n2513) );
  XNOR2X1 U1699 ( .A(n306), .B(n459), .Y(n2514) );
  XNOR2X1 U1700 ( .A(n306), .B(n3005), .Y(n2515) );
  XNOR2X1 U1701 ( .A(n306), .B(n455), .Y(n2516) );
  XNOR2X1 U1702 ( .A(n306), .B(n3008), .Y(n2517) );
  XNOR2X1 U1703 ( .A(n305), .B(n451), .Y(n2518) );
  XNOR2X1 U1704 ( .A(n305), .B(n3011), .Y(n2519) );
  XNOR2X1 U1705 ( .A(n305), .B(n447), .Y(n2520) );
  XNOR2X1 U1706 ( .A(n305), .B(b[5]), .Y(n2521) );
  XNOR2X1 U1707 ( .A(n305), .B(n443), .Y(n2522) );
  XNOR2X1 U1708 ( .A(n305), .B(b[3]), .Y(n2523) );
  XNOR2X1 U1709 ( .A(n305), .B(n439), .Y(n2524) );
  XNOR2X1 U1710 ( .A(n305), .B(b[1]), .Y(n2525) );
  XNOR2X1 U1711 ( .A(n305), .B(n3019), .Y(n2526) );
  OAI22X1 U1712 ( .A(n352), .B(n2560), .C(n2806), .D(n402), .Y(n1753) );
  OAI22X1 U1713 ( .A(n2806), .B(n352), .C(n2528), .D(n402), .Y(n2037) );
  OAI22X1 U1714 ( .A(n2528), .B(n352), .C(n2529), .D(n402), .Y(n2038) );
  OAI22X1 U1715 ( .A(n2529), .B(n352), .C(n2530), .D(n402), .Y(n2039) );
  OAI22X1 U1716 ( .A(n2530), .B(n352), .C(n2531), .D(n402), .Y(n2040) );
  OAI22X1 U1717 ( .A(n2531), .B(n352), .C(n2532), .D(n402), .Y(n2041) );
  OAI22X1 U1718 ( .A(n2532), .B(n352), .C(n2533), .D(n402), .Y(n2042) );
  OAI22X1 U1719 ( .A(n2533), .B(n352), .C(n2534), .D(n402), .Y(n2043) );
  OAI22X1 U1720 ( .A(n2534), .B(n352), .C(n2535), .D(n402), .Y(n2044) );
  OAI22X1 U1721 ( .A(n2535), .B(n352), .C(n2536), .D(n402), .Y(n2045) );
  OAI22X1 U1722 ( .A(n2536), .B(n351), .C(n2537), .D(n402), .Y(n2046) );
  OAI22X1 U1723 ( .A(n2537), .B(n351), .C(n2538), .D(n401), .Y(n2047) );
  OAI22X1 U1724 ( .A(n2538), .B(n351), .C(n2539), .D(n401), .Y(n2048) );
  OAI22X1 U1725 ( .A(n2539), .B(n351), .C(n2540), .D(n401), .Y(n2049) );
  OAI22X1 U1726 ( .A(n2540), .B(n351), .C(n2541), .D(n401), .Y(n2050) );
  OAI22X1 U1727 ( .A(n2541), .B(n351), .C(n2542), .D(n401), .Y(n2051) );
  OAI22X1 U1728 ( .A(n2542), .B(n351), .C(n2543), .D(n401), .Y(n2052) );
  OAI22X1 U1729 ( .A(n2543), .B(n351), .C(n2544), .D(n401), .Y(n2053) );
  OAI22X1 U1730 ( .A(n2544), .B(n351), .C(n2545), .D(n401), .Y(n2054) );
  OAI22X1 U1731 ( .A(n2545), .B(n351), .C(n2546), .D(n401), .Y(n2055) );
  OAI22X1 U1732 ( .A(n2546), .B(n351), .C(n2547), .D(n401), .Y(n2056) );
  OAI22X1 U1733 ( .A(n2547), .B(n351), .C(n2548), .D(n401), .Y(n2057) );
  OAI22X1 U1734 ( .A(n2548), .B(n350), .C(n2549), .D(n401), .Y(n2058) );
  OAI22X1 U1735 ( .A(n2549), .B(n350), .C(n2550), .D(n400), .Y(n2059) );
  OAI22X1 U1736 ( .A(n2550), .B(n350), .C(n2551), .D(n400), .Y(n2060) );
  OAI22X1 U1737 ( .A(n2551), .B(n350), .C(n2552), .D(n400), .Y(n2061) );
  OAI22X1 U1738 ( .A(n2552), .B(n350), .C(n2553), .D(n400), .Y(n2062) );
  OAI22X1 U1739 ( .A(n2553), .B(n350), .C(n2554), .D(n400), .Y(n2063) );
  OAI22X1 U1740 ( .A(n2554), .B(n350), .C(n2555), .D(n400), .Y(n2064) );
  OAI22X1 U1741 ( .A(n2555), .B(n350), .C(n2556), .D(n400), .Y(n2065) );
  OAI22X1 U1742 ( .A(n2556), .B(n350), .C(n2557), .D(n400), .Y(n2066) );
  OAI22X1 U1743 ( .A(n2557), .B(n350), .C(n2558), .D(n400), .Y(n2067) );
  OAI22X1 U1744 ( .A(n2558), .B(n350), .C(n2559), .D(n400), .Y(n2068) );
  XNOR2X1 U1745 ( .A(n304), .B(n2984), .Y(n2528) );
  XNOR2X1 U1746 ( .A(n304), .B(n495), .Y(n2529) );
  XNOR2X1 U1747 ( .A(n304), .B(b[29]), .Y(n2530) );
  XNOR2X1 U1748 ( .A(n304), .B(n491), .Y(n2531) );
  XNOR2X1 U1749 ( .A(n304), .B(n2986), .Y(n2532) );
  XNOR2X1 U1750 ( .A(n304), .B(n487), .Y(n2533) );
  XNOR2X1 U1751 ( .A(n304), .B(n2988), .Y(n2534) );
  XNOR2X1 U1752 ( .A(n304), .B(n483), .Y(n2535) );
  XNOR2X1 U1753 ( .A(n304), .B(n2990), .Y(n2536) );
  XNOR2X1 U1754 ( .A(n304), .B(n479), .Y(n2537) );
  XNOR2X1 U1755 ( .A(n304), .B(n2993), .Y(n2538) );
  XNOR2X1 U1756 ( .A(n303), .B(n475), .Y(n2539) );
  XNOR2X1 U1757 ( .A(n303), .B(n2996), .Y(n2540) );
  XNOR2X1 U1758 ( .A(n303), .B(n471), .Y(n2541) );
  XNOR2X1 U1759 ( .A(n303), .B(n2998), .Y(n2542) );
  XNOR2X1 U1760 ( .A(n303), .B(n467), .Y(n2543) );
  XNOR2X1 U1761 ( .A(n303), .B(b[15]), .Y(n2544) );
  XNOR2X1 U1762 ( .A(n303), .B(n463), .Y(n2545) );
  XNOR2X1 U1763 ( .A(n303), .B(b[13]), .Y(n2546) );
  XNOR2X1 U1764 ( .A(n303), .B(n459), .Y(n2547) );
  XNOR2X1 U1765 ( .A(n303), .B(n3005), .Y(n2548) );
  XNOR2X1 U1766 ( .A(n303), .B(n455), .Y(n2549) );
  XNOR2X1 U1767 ( .A(n303), .B(n3008), .Y(n2550) );
  XNOR2X1 U1768 ( .A(n302), .B(n451), .Y(n2551) );
  XNOR2X1 U1769 ( .A(n302), .B(n3011), .Y(n2552) );
  XNOR2X1 U1770 ( .A(n302), .B(n447), .Y(n2553) );
  XNOR2X1 U1771 ( .A(n302), .B(b[5]), .Y(n2554) );
  XNOR2X1 U1772 ( .A(n302), .B(n443), .Y(n2555) );
  XNOR2X1 U1773 ( .A(n302), .B(b[3]), .Y(n2556) );
  XNOR2X1 U1774 ( .A(n302), .B(n439), .Y(n2557) );
  XNOR2X1 U1775 ( .A(n302), .B(b[1]), .Y(n2558) );
  XNOR2X1 U1776 ( .A(n302), .B(n3019), .Y(n2559) );
  OAI22X1 U1777 ( .A(n349), .B(n2593), .C(n2807), .D(n399), .Y(n1754) );
  OAI22X1 U1778 ( .A(n2807), .B(n349), .C(n2561), .D(n399), .Y(n2071) );
  OAI22X1 U1779 ( .A(n2561), .B(n349), .C(n2562), .D(n399), .Y(n2072) );
  OAI22X1 U1780 ( .A(n2562), .B(n349), .C(n2563), .D(n399), .Y(n2073) );
  OAI22X1 U1781 ( .A(n2563), .B(n349), .C(n2564), .D(n399), .Y(n2074) );
  OAI22X1 U1782 ( .A(n2564), .B(n349), .C(n2565), .D(n399), .Y(n2075) );
  OAI22X1 U1783 ( .A(n2565), .B(n349), .C(n2566), .D(n399), .Y(n2076) );
  OAI22X1 U1784 ( .A(n2566), .B(n349), .C(n2567), .D(n399), .Y(n2077) );
  OAI22X1 U1785 ( .A(n2567), .B(n349), .C(n2568), .D(n399), .Y(n2078) );
  OAI22X1 U1786 ( .A(n2568), .B(n349), .C(n2569), .D(n399), .Y(n2079) );
  OAI22X1 U1787 ( .A(n2569), .B(n348), .C(n2570), .D(n399), .Y(n2080) );
  OAI22X1 U1788 ( .A(n2570), .B(n348), .C(n2571), .D(n398), .Y(n2081) );
  OAI22X1 U1789 ( .A(n2571), .B(n348), .C(n2572), .D(n398), .Y(n2082) );
  OAI22X1 U1790 ( .A(n2572), .B(n348), .C(n2573), .D(n398), .Y(n2083) );
  OAI22X1 U1791 ( .A(n2573), .B(n348), .C(n2574), .D(n398), .Y(n2084) );
  OAI22X1 U1792 ( .A(n2574), .B(n348), .C(n2575), .D(n398), .Y(n2085) );
  OAI22X1 U1793 ( .A(n2575), .B(n348), .C(n2576), .D(n398), .Y(n2086) );
  OAI22X1 U1794 ( .A(n2576), .B(n348), .C(n2577), .D(n398), .Y(n2087) );
  OAI22X1 U1795 ( .A(n2577), .B(n348), .C(n2578), .D(n398), .Y(n2088) );
  OAI22X1 U1796 ( .A(n2578), .B(n348), .C(n2579), .D(n398), .Y(n2089) );
  OAI22X1 U1797 ( .A(n2579), .B(n348), .C(n2580), .D(n398), .Y(n2090) );
  OAI22X1 U1798 ( .A(n2580), .B(n348), .C(n2581), .D(n398), .Y(n2091) );
  OAI22X1 U1799 ( .A(n2581), .B(n347), .C(n2582), .D(n398), .Y(n2092) );
  OAI22X1 U1800 ( .A(n2582), .B(n347), .C(n2583), .D(n397), .Y(n2093) );
  OAI22X1 U1801 ( .A(n2583), .B(n347), .C(n2584), .D(n397), .Y(n2094) );
  OAI22X1 U1802 ( .A(n2584), .B(n347), .C(n2585), .D(n397), .Y(n2095) );
  OAI22X1 U1803 ( .A(n2585), .B(n347), .C(n2586), .D(n397), .Y(n2096) );
  OAI22X1 U1804 ( .A(n2586), .B(n347), .C(n2587), .D(n397), .Y(n2097) );
  OAI22X1 U1805 ( .A(n2587), .B(n347), .C(n2588), .D(n397), .Y(n2098) );
  OAI22X1 U1806 ( .A(n2588), .B(n347), .C(n2589), .D(n397), .Y(n2099) );
  OAI22X1 U1807 ( .A(n2589), .B(n347), .C(n2590), .D(n397), .Y(n2100) );
  OAI22X1 U1808 ( .A(n2590), .B(n347), .C(n2591), .D(n397), .Y(n2101) );
  OAI22X1 U1809 ( .A(n2591), .B(n347), .C(n2592), .D(n397), .Y(n2102) );
  XNOR2X1 U1810 ( .A(n301), .B(n2984), .Y(n2561) );
  XNOR2X1 U1811 ( .A(n301), .B(n495), .Y(n2562) );
  XNOR2X1 U1812 ( .A(n301), .B(b[29]), .Y(n2563) );
  XNOR2X1 U1813 ( .A(n301), .B(n491), .Y(n2564) );
  XNOR2X1 U1814 ( .A(n301), .B(n2986), .Y(n2565) );
  XNOR2X1 U1815 ( .A(n301), .B(n487), .Y(n2566) );
  XNOR2X1 U1816 ( .A(n301), .B(n2988), .Y(n2567) );
  XNOR2X1 U1817 ( .A(n301), .B(n483), .Y(n2568) );
  XNOR2X1 U1818 ( .A(n301), .B(n2990), .Y(n2569) );
  XNOR2X1 U1819 ( .A(n301), .B(n479), .Y(n2570) );
  XNOR2X1 U1820 ( .A(n301), .B(n2993), .Y(n2571) );
  XNOR2X1 U1821 ( .A(n300), .B(n475), .Y(n2572) );
  XNOR2X1 U1822 ( .A(n300), .B(n2996), .Y(n2573) );
  XNOR2X1 U1823 ( .A(n300), .B(n471), .Y(n2574) );
  XNOR2X1 U1824 ( .A(n300), .B(n2998), .Y(n2575) );
  XNOR2X1 U1825 ( .A(n300), .B(n467), .Y(n2576) );
  XNOR2X1 U1826 ( .A(n300), .B(b[15]), .Y(n2577) );
  XNOR2X1 U1827 ( .A(n300), .B(n463), .Y(n2578) );
  XNOR2X1 U1828 ( .A(n300), .B(b[13]), .Y(n2579) );
  XNOR2X1 U1829 ( .A(n300), .B(n459), .Y(n2580) );
  XNOR2X1 U1830 ( .A(n300), .B(n3005), .Y(n2581) );
  XNOR2X1 U1831 ( .A(n300), .B(n455), .Y(n2582) );
  XNOR2X1 U1832 ( .A(n300), .B(n3008), .Y(n2583) );
  XNOR2X1 U1833 ( .A(n299), .B(n451), .Y(n2584) );
  XNOR2X1 U1834 ( .A(n299), .B(n3011), .Y(n2585) );
  XNOR2X1 U1835 ( .A(n299), .B(n447), .Y(n2586) );
  XNOR2X1 U1836 ( .A(n299), .B(b[5]), .Y(n2587) );
  XNOR2X1 U1837 ( .A(n299), .B(n443), .Y(n2588) );
  XNOR2X1 U1838 ( .A(n299), .B(b[3]), .Y(n2589) );
  XNOR2X1 U1839 ( .A(n299), .B(n439), .Y(n2590) );
  XNOR2X1 U1840 ( .A(n299), .B(b[1]), .Y(n2591) );
  XNOR2X1 U1841 ( .A(n299), .B(n3019), .Y(n2592) );
  OAI22X1 U1842 ( .A(n346), .B(n2626), .C(n2808), .D(n396), .Y(n1755) );
  OAI22X1 U1843 ( .A(n2808), .B(n346), .C(n2594), .D(n396), .Y(n2105) );
  OAI22X1 U1844 ( .A(n2594), .B(n346), .C(n2595), .D(n396), .Y(n2106) );
  OAI22X1 U1845 ( .A(n2595), .B(n346), .C(n2596), .D(n396), .Y(n2107) );
  OAI22X1 U1846 ( .A(n2596), .B(n346), .C(n2597), .D(n396), .Y(n2108) );
  OAI22X1 U1847 ( .A(n2597), .B(n346), .C(n2598), .D(n396), .Y(n2109) );
  OAI22X1 U1848 ( .A(n2598), .B(n346), .C(n2599), .D(n396), .Y(n2110) );
  OAI22X1 U1849 ( .A(n2599), .B(n346), .C(n2600), .D(n396), .Y(n2111) );
  OAI22X1 U1850 ( .A(n2600), .B(n346), .C(n2601), .D(n396), .Y(n2112) );
  OAI22X1 U1851 ( .A(n2601), .B(n346), .C(n2602), .D(n396), .Y(n2113) );
  OAI22X1 U1852 ( .A(n2602), .B(n345), .C(n2603), .D(n396), .Y(n2114) );
  OAI22X1 U1853 ( .A(n2603), .B(n345), .C(n2604), .D(n395), .Y(n2115) );
  OAI22X1 U1854 ( .A(n2604), .B(n345), .C(n2605), .D(n395), .Y(n2116) );
  OAI22X1 U1855 ( .A(n2605), .B(n345), .C(n2606), .D(n395), .Y(n2117) );
  OAI22X1 U1856 ( .A(n2606), .B(n345), .C(n2607), .D(n395), .Y(n2118) );
  OAI22X1 U1857 ( .A(n2607), .B(n345), .C(n2608), .D(n395), .Y(n2119) );
  OAI22X1 U1858 ( .A(n2608), .B(n345), .C(n2609), .D(n395), .Y(n2120) );
  OAI22X1 U1859 ( .A(n2609), .B(n345), .C(n2610), .D(n395), .Y(n2121) );
  OAI22X1 U1860 ( .A(n2610), .B(n345), .C(n2611), .D(n395), .Y(n2122) );
  OAI22X1 U1861 ( .A(n2611), .B(n345), .C(n2612), .D(n395), .Y(n2123) );
  OAI22X1 U1862 ( .A(n2612), .B(n345), .C(n2613), .D(n395), .Y(n2124) );
  OAI22X1 U1863 ( .A(n2613), .B(n345), .C(n2614), .D(n395), .Y(n2125) );
  OAI22X1 U1864 ( .A(n2614), .B(n344), .C(n2615), .D(n395), .Y(n2126) );
  OAI22X1 U1865 ( .A(n2615), .B(n344), .C(n2616), .D(n394), .Y(n2127) );
  OAI22X1 U1866 ( .A(n2616), .B(n344), .C(n2617), .D(n394), .Y(n2128) );
  OAI22X1 U1867 ( .A(n2617), .B(n344), .C(n2618), .D(n394), .Y(n2129) );
  OAI22X1 U1868 ( .A(n2618), .B(n344), .C(n2619), .D(n394), .Y(n2130) );
  OAI22X1 U1869 ( .A(n2619), .B(n344), .C(n2620), .D(n394), .Y(n2131) );
  OAI22X1 U1870 ( .A(n2620), .B(n344), .C(n2621), .D(n394), .Y(n2132) );
  OAI22X1 U1871 ( .A(n2621), .B(n344), .C(n2622), .D(n394), .Y(n2133) );
  OAI22X1 U1872 ( .A(n2622), .B(n344), .C(n2623), .D(n394), .Y(n2134) );
  OAI22X1 U1873 ( .A(n2623), .B(n344), .C(n2624), .D(n394), .Y(n2135) );
  OAI22X1 U1874 ( .A(n2624), .B(n344), .C(n2625), .D(n394), .Y(n2136) );
  XNOR2X1 U1875 ( .A(n298), .B(n2984), .Y(n2594) );
  XNOR2X1 U1876 ( .A(n298), .B(n495), .Y(n2595) );
  XNOR2X1 U1877 ( .A(n298), .B(b[29]), .Y(n2596) );
  XNOR2X1 U1878 ( .A(n298), .B(n491), .Y(n2597) );
  XNOR2X1 U1879 ( .A(n298), .B(n2986), .Y(n2598) );
  XNOR2X1 U1880 ( .A(n298), .B(n487), .Y(n2599) );
  XNOR2X1 U1881 ( .A(n298), .B(n2988), .Y(n2600) );
  XNOR2X1 U1882 ( .A(n298), .B(n483), .Y(n2601) );
  XNOR2X1 U1883 ( .A(n298), .B(n2990), .Y(n2602) );
  XNOR2X1 U1884 ( .A(n298), .B(n479), .Y(n2603) );
  XNOR2X1 U1885 ( .A(n298), .B(n2993), .Y(n2604) );
  XNOR2X1 U1886 ( .A(n297), .B(n475), .Y(n2605) );
  XNOR2X1 U1887 ( .A(n297), .B(n2996), .Y(n2606) );
  XNOR2X1 U1888 ( .A(n297), .B(n471), .Y(n2607) );
  XNOR2X1 U1889 ( .A(n297), .B(n2998), .Y(n2608) );
  XNOR2X1 U1890 ( .A(n297), .B(n467), .Y(n2609) );
  XNOR2X1 U1891 ( .A(n297), .B(n3000), .Y(n2610) );
  XNOR2X1 U1892 ( .A(n297), .B(n463), .Y(n2611) );
  XNOR2X1 U1893 ( .A(n297), .B(n3002), .Y(n2612) );
  XNOR2X1 U1894 ( .A(n297), .B(n459), .Y(n2613) );
  XNOR2X1 U1895 ( .A(n297), .B(n3004), .Y(n2614) );
  XNOR2X1 U1896 ( .A(n297), .B(n455), .Y(n2615) );
  XNOR2X1 U1897 ( .A(n297), .B(n3007), .Y(n2616) );
  XNOR2X1 U1898 ( .A(n2913), .B(n451), .Y(n2617) );
  XNOR2X1 U1899 ( .A(n2913), .B(n3010), .Y(n2618) );
  XNOR2X1 U1900 ( .A(n2914), .B(n447), .Y(n2619) );
  XNOR2X1 U1901 ( .A(n2913), .B(n3013), .Y(n2620) );
  XNOR2X1 U1902 ( .A(n2914), .B(n443), .Y(n2621) );
  XNOR2X1 U1903 ( .A(n2914), .B(n3015), .Y(n2622) );
  XNOR2X1 U1904 ( .A(n2913), .B(n439), .Y(n2623) );
  XNOR2X1 U1905 ( .A(n2912), .B(n3017), .Y(n2624) );
  XNOR2X1 U1906 ( .A(n2914), .B(n3019), .Y(n2625) );
  OAI22X1 U1907 ( .A(n343), .B(n2659), .C(n2809), .D(n393), .Y(n1756) );
  OAI22X1 U1908 ( .A(n2809), .B(n343), .C(n2627), .D(n393), .Y(n2139) );
  OAI22X1 U1909 ( .A(n2627), .B(n343), .C(n2628), .D(n393), .Y(n2140) );
  OAI22X1 U1910 ( .A(n2628), .B(n343), .C(n2629), .D(n393), .Y(n2141) );
  OAI22X1 U1911 ( .A(n2629), .B(n343), .C(n2630), .D(n393), .Y(n2142) );
  OAI22X1 U1912 ( .A(n2630), .B(n343), .C(n2631), .D(n393), .Y(n2143) );
  OAI22X1 U1913 ( .A(n2631), .B(n343), .C(n2632), .D(n393), .Y(n2144) );
  OAI22X1 U1914 ( .A(n2632), .B(n343), .C(n2633), .D(n393), .Y(n2145) );
  OAI22X1 U1915 ( .A(n2633), .B(n343), .C(n2634), .D(n393), .Y(n2146) );
  OAI22X1 U1916 ( .A(n2634), .B(n343), .C(n2635), .D(n393), .Y(n2147) );
  OAI22X1 U1917 ( .A(n2635), .B(n342), .C(n2636), .D(n393), .Y(n2148) );
  OAI22X1 U1918 ( .A(n2636), .B(n342), .C(n2637), .D(n392), .Y(n2149) );
  OAI22X1 U1919 ( .A(n2637), .B(n342), .C(n2638), .D(n392), .Y(n2150) );
  OAI22X1 U1920 ( .A(n2638), .B(n342), .C(n2639), .D(n392), .Y(n2151) );
  OAI22X1 U1921 ( .A(n2639), .B(n342), .C(n2640), .D(n392), .Y(n2152) );
  OAI22X1 U1922 ( .A(n2640), .B(n342), .C(n2641), .D(n392), .Y(n2153) );
  OAI22X1 U1923 ( .A(n2641), .B(n342), .C(n2642), .D(n392), .Y(n2154) );
  OAI22X1 U1924 ( .A(n2642), .B(n342), .C(n2643), .D(n392), .Y(n2155) );
  OAI22X1 U1925 ( .A(n2643), .B(n342), .C(n2644), .D(n392), .Y(n2156) );
  OAI22X1 U1926 ( .A(n2644), .B(n342), .C(n2645), .D(n392), .Y(n2157) );
  OAI22X1 U1927 ( .A(n2645), .B(n342), .C(n2646), .D(n392), .Y(n2158) );
  OAI22X1 U1928 ( .A(n2646), .B(n342), .C(n2647), .D(n392), .Y(n2159) );
  OAI22X1 U1929 ( .A(n2647), .B(n341), .C(n2648), .D(n392), .Y(n2160) );
  OAI22X1 U1930 ( .A(n2648), .B(n341), .C(n2649), .D(n391), .Y(n2161) );
  OAI22X1 U1931 ( .A(n2649), .B(n341), .C(n2650), .D(n391), .Y(n2162) );
  OAI22X1 U1932 ( .A(n2650), .B(n341), .C(n2651), .D(n391), .Y(n2163) );
  OAI22X1 U1933 ( .A(n2651), .B(n341), .C(n2652), .D(n391), .Y(n2164) );
  OAI22X1 U1934 ( .A(n2652), .B(n341), .C(n2653), .D(n391), .Y(n2165) );
  OAI22X1 U1935 ( .A(n2653), .B(n341), .C(n2654), .D(n391), .Y(n2166) );
  OAI22X1 U1936 ( .A(n2654), .B(n341), .C(n2655), .D(n391), .Y(n2167) );
  OAI22X1 U1937 ( .A(n2655), .B(n341), .C(n2656), .D(n391), .Y(n2168) );
  OAI22X1 U1938 ( .A(n2656), .B(n341), .C(n2657), .D(n391), .Y(n2169) );
  OAI22X1 U1939 ( .A(n2657), .B(n341), .C(n2658), .D(n391), .Y(n2170) );
  XNOR2X1 U1940 ( .A(n295), .B(n2984), .Y(n2627) );
  XNOR2X1 U1941 ( .A(n295), .B(n495), .Y(n2628) );
  XNOR2X1 U1942 ( .A(n295), .B(b[29]), .Y(n2629) );
  XNOR2X1 U1943 ( .A(n295), .B(n491), .Y(n2630) );
  XNOR2X1 U1944 ( .A(n295), .B(n2986), .Y(n2631) );
  XNOR2X1 U1945 ( .A(n295), .B(n487), .Y(n2632) );
  XNOR2X1 U1946 ( .A(n295), .B(n2988), .Y(n2633) );
  XNOR2X1 U1947 ( .A(n295), .B(n483), .Y(n2634) );
  XNOR2X1 U1948 ( .A(n295), .B(n2990), .Y(n2635) );
  XNOR2X1 U1949 ( .A(n295), .B(n479), .Y(n2636) );
  XNOR2X1 U1950 ( .A(n295), .B(n2993), .Y(n2637) );
  XNOR2X1 U1951 ( .A(n294), .B(n475), .Y(n2638) );
  XNOR2X1 U1952 ( .A(n294), .B(n2996), .Y(n2639) );
  XNOR2X1 U1953 ( .A(n294), .B(n471), .Y(n2640) );
  XNOR2X1 U1954 ( .A(n294), .B(n2998), .Y(n2641) );
  XNOR2X1 U1955 ( .A(n294), .B(n467), .Y(n2642) );
  XNOR2X1 U1956 ( .A(n294), .B(n3000), .Y(n2643) );
  XNOR2X1 U1957 ( .A(n294), .B(n463), .Y(n2644) );
  XNOR2X1 U1958 ( .A(n294), .B(n3002), .Y(n2645) );
  XNOR2X1 U1959 ( .A(n294), .B(n459), .Y(n2646) );
  XNOR2X1 U1960 ( .A(n294), .B(n3004), .Y(n2647) );
  XNOR2X1 U1961 ( .A(n294), .B(n455), .Y(n2648) );
  XNOR2X1 U1962 ( .A(n294), .B(n3007), .Y(n2649) );
  XNOR2X1 U1963 ( .A(n293), .B(n451), .Y(n2650) );
  XNOR2X1 U1964 ( .A(n293), .B(n3010), .Y(n2651) );
  XNOR2X1 U1965 ( .A(n293), .B(n447), .Y(n2652) );
  XNOR2X1 U1966 ( .A(n293), .B(n3013), .Y(n2653) );
  XNOR2X1 U1967 ( .A(n293), .B(n443), .Y(n2654) );
  XNOR2X1 U1968 ( .A(n293), .B(n3015), .Y(n2655) );
  XNOR2X1 U1969 ( .A(n293), .B(n439), .Y(n2656) );
  XNOR2X1 U1970 ( .A(n293), .B(n3017), .Y(n2657) );
  XNOR2X1 U1971 ( .A(n293), .B(n3019), .Y(n2658) );
  OAI22X1 U1972 ( .A(n340), .B(n2692), .C(n2810), .D(n390), .Y(n1757) );
  OAI22X1 U1973 ( .A(n2810), .B(n340), .C(n2660), .D(n390), .Y(n2173) );
  OAI22X1 U1974 ( .A(n2660), .B(n340), .C(n2661), .D(n390), .Y(n2174) );
  OAI22X1 U1975 ( .A(n2661), .B(n340), .C(n2662), .D(n390), .Y(n2175) );
  OAI22X1 U1976 ( .A(n2662), .B(n340), .C(n2663), .D(n390), .Y(n2176) );
  OAI22X1 U1977 ( .A(n2663), .B(n340), .C(n2664), .D(n390), .Y(n2177) );
  OAI22X1 U1978 ( .A(n2664), .B(n340), .C(n2665), .D(n390), .Y(n2178) );
  OAI22X1 U1979 ( .A(n2665), .B(n340), .C(n2666), .D(n390), .Y(n2179) );
  OAI22X1 U1980 ( .A(n2666), .B(n340), .C(n2667), .D(n390), .Y(n2180) );
  OAI22X1 U1981 ( .A(n2667), .B(n340), .C(n2668), .D(n390), .Y(n2181) );
  OAI22X1 U1982 ( .A(n2668), .B(n339), .C(n2669), .D(n390), .Y(n2182) );
  OAI22X1 U1983 ( .A(n2669), .B(n339), .C(n2670), .D(n389), .Y(n2183) );
  OAI22X1 U1984 ( .A(n2670), .B(n339), .C(n2671), .D(n389), .Y(n2184) );
  OAI22X1 U1985 ( .A(n2671), .B(n339), .C(n2672), .D(n389), .Y(n2185) );
  OAI22X1 U1986 ( .A(n2672), .B(n339), .C(n2673), .D(n389), .Y(n2186) );
  OAI22X1 U1987 ( .A(n2673), .B(n339), .C(n2674), .D(n389), .Y(n2187) );
  OAI22X1 U1988 ( .A(n2674), .B(n339), .C(n2675), .D(n389), .Y(n2188) );
  OAI22X1 U1989 ( .A(n2675), .B(n339), .C(n2676), .D(n389), .Y(n2189) );
  OAI22X1 U1990 ( .A(n2676), .B(n339), .C(n2677), .D(n389), .Y(n2190) );
  OAI22X1 U1991 ( .A(n2677), .B(n339), .C(n2678), .D(n389), .Y(n2191) );
  OAI22X1 U1992 ( .A(n2678), .B(n339), .C(n2679), .D(n389), .Y(n2192) );
  OAI22X1 U1993 ( .A(n2679), .B(n339), .C(n2680), .D(n389), .Y(n2193) );
  OAI22X1 U1994 ( .A(n2680), .B(n338), .C(n2681), .D(n389), .Y(n2194) );
  OAI22X1 U1995 ( .A(n2681), .B(n338), .C(n2682), .D(n388), .Y(n2195) );
  OAI22X1 U1996 ( .A(n2682), .B(n338), .C(n2683), .D(n388), .Y(n2196) );
  OAI22X1 U1997 ( .A(n2683), .B(n338), .C(n2684), .D(n388), .Y(n2197) );
  OAI22X1 U1998 ( .A(n2684), .B(n338), .C(n2685), .D(n388), .Y(n2198) );
  OAI22X1 U1999 ( .A(n2685), .B(n338), .C(n2686), .D(n388), .Y(n2199) );
  OAI22X1 U2000 ( .A(n2686), .B(n338), .C(n2687), .D(n388), .Y(n2200) );
  OAI22X1 U2001 ( .A(n2687), .B(n338), .C(n2688), .D(n388), .Y(n2201) );
  OAI22X1 U2002 ( .A(n2688), .B(n338), .C(n2689), .D(n388), .Y(n2202) );
  OAI22X1 U2003 ( .A(n2689), .B(n338), .C(n2690), .D(n388), .Y(n2203) );
  OAI22X1 U2004 ( .A(n2690), .B(n338), .C(n2691), .D(n388), .Y(n2204) );
  XNOR2X1 U2005 ( .A(n292), .B(n2984), .Y(n2660) );
  XNOR2X1 U2006 ( .A(n292), .B(n495), .Y(n2661) );
  XNOR2X1 U2007 ( .A(n292), .B(b[29]), .Y(n2662) );
  XNOR2X1 U2008 ( .A(n292), .B(n491), .Y(n2663) );
  XNOR2X1 U2009 ( .A(n292), .B(n2986), .Y(n2664) );
  XNOR2X1 U2010 ( .A(n292), .B(n487), .Y(n2665) );
  XNOR2X1 U2011 ( .A(n292), .B(n2988), .Y(n2666) );
  XNOR2X1 U2012 ( .A(n292), .B(n483), .Y(n2667) );
  XNOR2X1 U2013 ( .A(n292), .B(n2990), .Y(n2668) );
  XNOR2X1 U2014 ( .A(n292), .B(n479), .Y(n2669) );
  XNOR2X1 U2015 ( .A(n292), .B(n2993), .Y(n2670) );
  XNOR2X1 U2016 ( .A(n2916), .B(n475), .Y(n2671) );
  XNOR2X1 U2017 ( .A(n2917), .B(n2996), .Y(n2672) );
  XNOR2X1 U2018 ( .A(n2917), .B(n471), .Y(n2673) );
  XNOR2X1 U2019 ( .A(n2916), .B(n2998), .Y(n2674) );
  XNOR2X1 U2020 ( .A(n2915), .B(n467), .Y(n2675) );
  XNOR2X1 U2021 ( .A(n2915), .B(n3000), .Y(n2676) );
  XNOR2X1 U2022 ( .A(n2917), .B(n463), .Y(n2677) );
  XNOR2X1 U2023 ( .A(n2916), .B(n3002), .Y(n2678) );
  XNOR2X1 U2024 ( .A(n2915), .B(n459), .Y(n2679) );
  XNOR2X1 U2025 ( .A(n2916), .B(n3004), .Y(n2680) );
  XNOR2X1 U2026 ( .A(n2917), .B(n455), .Y(n2681) );
  XNOR2X1 U2027 ( .A(n2916), .B(n3007), .Y(n2682) );
  XNOR2X1 U2028 ( .A(n290), .B(n451), .Y(n2683) );
  XNOR2X1 U2029 ( .A(n290), .B(n3010), .Y(n2684) );
  XNOR2X1 U2030 ( .A(n290), .B(n447), .Y(n2685) );
  XNOR2X1 U2031 ( .A(n290), .B(n3013), .Y(n2686) );
  XNOR2X1 U2032 ( .A(n290), .B(n443), .Y(n2687) );
  XNOR2X1 U2033 ( .A(n290), .B(n3015), .Y(n2688) );
  XNOR2X1 U2034 ( .A(n290), .B(n439), .Y(n2689) );
  XNOR2X1 U2035 ( .A(n290), .B(n3017), .Y(n2690) );
  XNOR2X1 U2036 ( .A(n290), .B(n3019), .Y(n2691) );
  OAI22X1 U2037 ( .A(n337), .B(n2725), .C(n2811), .D(n387), .Y(n1758) );
  OAI22X1 U2038 ( .A(n337), .B(n2811), .C(n2693), .D(n387), .Y(n2207) );
  OAI22X1 U2039 ( .A(n337), .B(n2693), .C(n2694), .D(n387), .Y(n2208) );
  OAI22X1 U2040 ( .A(n337), .B(n2694), .C(n2695), .D(n387), .Y(n2209) );
  OAI22X1 U2041 ( .A(n337), .B(n2695), .C(n2696), .D(n387), .Y(n2210) );
  OAI22X1 U2042 ( .A(n337), .B(n2696), .C(n2697), .D(n387), .Y(n2211) );
  OAI22X1 U2043 ( .A(n337), .B(n2697), .C(n2698), .D(n387), .Y(n2212) );
  OAI22X1 U2044 ( .A(n337), .B(n2698), .C(n2699), .D(n387), .Y(n2213) );
  OAI22X1 U2045 ( .A(n337), .B(n2699), .C(n2700), .D(n387), .Y(n2214) );
  OAI22X1 U2046 ( .A(n337), .B(n2700), .C(n2701), .D(n387), .Y(n2215) );
  OAI22X1 U2047 ( .A(n336), .B(n2701), .C(n2702), .D(n387), .Y(n2216) );
  OAI22X1 U2048 ( .A(n336), .B(n2702), .C(n2703), .D(n386), .Y(n2217) );
  OAI22X1 U2049 ( .A(n336), .B(n2703), .C(n2704), .D(n386), .Y(n2218) );
  OAI22X1 U2050 ( .A(n336), .B(n2704), .C(n2705), .D(n386), .Y(n2219) );
  OAI22X1 U2051 ( .A(n336), .B(n2705), .C(n2706), .D(n386), .Y(n2220) );
  OAI22X1 U2052 ( .A(n336), .B(n2706), .C(n2707), .D(n386), .Y(n2221) );
  OAI22X1 U2053 ( .A(n336), .B(n2707), .C(n2708), .D(n386), .Y(n2222) );
  OAI22X1 U2054 ( .A(n336), .B(n2708), .C(n2709), .D(n386), .Y(n2223) );
  OAI22X1 U2055 ( .A(n336), .B(n2709), .C(n2710), .D(n386), .Y(n2224) );
  OAI22X1 U2056 ( .A(n336), .B(n2710), .C(n2711), .D(n386), .Y(n2225) );
  OAI22X1 U2057 ( .A(n336), .B(n2711), .C(n2712), .D(n386), .Y(n2226) );
  OAI22X1 U2058 ( .A(n336), .B(n2712), .C(n2713), .D(n386), .Y(n2227) );
  OAI22X1 U2059 ( .A(n335), .B(n2713), .C(n2714), .D(n386), .Y(n2228) );
  OAI22X1 U2060 ( .A(n335), .B(n2714), .C(n2715), .D(n385), .Y(n2229) );
  OAI22X1 U2061 ( .A(n335), .B(n2715), .C(n2716), .D(n385), .Y(n2230) );
  OAI22X1 U2062 ( .A(n335), .B(n2716), .C(n2717), .D(n385), .Y(n2231) );
  OAI22X1 U2063 ( .A(n335), .B(n2717), .C(n2718), .D(n385), .Y(n2232) );
  OAI22X1 U2064 ( .A(n335), .B(n2718), .C(n2719), .D(n385), .Y(n2233) );
  OAI22X1 U2065 ( .A(n335), .B(n2719), .C(n2720), .D(n385), .Y(n2234) );
  OAI22X1 U2066 ( .A(n335), .B(n2720), .C(n2721), .D(n385), .Y(n2235) );
  OAI22X1 U2067 ( .A(n335), .B(n2721), .C(n2722), .D(n385), .Y(n2236) );
  OAI22X1 U2068 ( .A(n335), .B(n2722), .C(n2723), .D(n385), .Y(n2237) );
  OAI22X1 U2069 ( .A(n335), .B(n2723), .C(n2724), .D(n385), .Y(n2238) );
  XNOR2X1 U2070 ( .A(n289), .B(n2984), .Y(n2693) );
  XNOR2X1 U2071 ( .A(n289), .B(n495), .Y(n2694) );
  XNOR2X1 U2072 ( .A(n289), .B(b[29]), .Y(n2695) );
  XNOR2X1 U2073 ( .A(n289), .B(n491), .Y(n2696) );
  XNOR2X1 U2074 ( .A(n289), .B(n2986), .Y(n2697) );
  XNOR2X1 U2075 ( .A(n289), .B(n487), .Y(n2698) );
  XNOR2X1 U2076 ( .A(n289), .B(n2988), .Y(n2699) );
  XNOR2X1 U2077 ( .A(n289), .B(n483), .Y(n2700) );
  XNOR2X1 U2078 ( .A(n289), .B(n2990), .Y(n2701) );
  XNOR2X1 U2079 ( .A(n289), .B(n479), .Y(n2702) );
  XNOR2X1 U2080 ( .A(n289), .B(n2993), .Y(n2703) );
  XNOR2X1 U2081 ( .A(n288), .B(n475), .Y(n2704) );
  XNOR2X1 U2082 ( .A(n288), .B(n2996), .Y(n2705) );
  XNOR2X1 U2083 ( .A(n288), .B(n471), .Y(n2706) );
  XNOR2X1 U2084 ( .A(n288), .B(n2998), .Y(n2707) );
  XNOR2X1 U2085 ( .A(n288), .B(n467), .Y(n2708) );
  XNOR2X1 U2086 ( .A(n288), .B(n3000), .Y(n2709) );
  XNOR2X1 U2087 ( .A(n288), .B(n463), .Y(n2710) );
  XNOR2X1 U2088 ( .A(n288), .B(n3002), .Y(n2711) );
  XNOR2X1 U2089 ( .A(n288), .B(n459), .Y(n2712) );
  XNOR2X1 U2090 ( .A(n288), .B(n3004), .Y(n2713) );
  XNOR2X1 U2091 ( .A(n288), .B(n455), .Y(n2714) );
  XNOR2X1 U2092 ( .A(n288), .B(n3007), .Y(n2715) );
  XNOR2X1 U2093 ( .A(n287), .B(n451), .Y(n2716) );
  XNOR2X1 U2094 ( .A(n287), .B(n3010), .Y(n2717) );
  XNOR2X1 U2095 ( .A(n287), .B(n447), .Y(n2718) );
  XNOR2X1 U2096 ( .A(n287), .B(n3013), .Y(n2719) );
  XNOR2X1 U2097 ( .A(n287), .B(n443), .Y(n2720) );
  XNOR2X1 U2098 ( .A(n287), .B(n3015), .Y(n2721) );
  XNOR2X1 U2099 ( .A(n287), .B(n439), .Y(n2722) );
  XNOR2X1 U2100 ( .A(n287), .B(n3017), .Y(n2723) );
  XNOR2X1 U2101 ( .A(n287), .B(n3019), .Y(n2724) );
  INVX2 U2104 ( .A(n329), .Y(n2797) );
  INVX2 U2108 ( .A(n2966), .Y(n2799) );
  INVX2 U2110 ( .A(n320), .Y(n2800) );
  INVX2 U2112 ( .A(n317), .Y(n2801) );
  INVX2 U2114 ( .A(n314), .Y(n2802) );
  INVX2 U2116 ( .A(n2965), .Y(n2803) );
  INVX2 U2118 ( .A(n2911), .Y(n2804) );
  INVX2 U2120 ( .A(n305), .Y(n2805) );
  INVX2 U2122 ( .A(n302), .Y(n2806) );
  INVX2 U2124 ( .A(n299), .Y(n2807) );
  INVX2 U2126 ( .A(n2914), .Y(n2808) );
  INVX2 U2128 ( .A(n293), .Y(n2809) );
  INVX2 U2130 ( .A(n290), .Y(n2810) );
  INVX2 U2132 ( .A(n287), .Y(n2811) );
  INVX2 U2134 ( .A(a[31]), .Y(n384) );
  NAND2X1 U2135 ( .A(n2752), .B(n2780), .Y(n432) );
  XOR2X1 U2136 ( .A(a[30]), .B(a[31]), .Y(n2752) );
  XNOR2X1 U2137 ( .A(a[30]), .B(a[29]), .Y(n2780) );
  NAND2X1 U2138 ( .A(n2753), .B(n2781), .Y(n429) );
  XOR2X1 U2139 ( .A(a[28]), .B(a[29]), .Y(n2753) );
  XNOR2X1 U2140 ( .A(a[28]), .B(a[27]), .Y(n2781) );
  NAND2X1 U2141 ( .A(n2754), .B(n2782), .Y(n426) );
  XOR2X1 U2142 ( .A(a[26]), .B(a[27]), .Y(n2754) );
  XNOR2X1 U2143 ( .A(a[26]), .B(a[25]), .Y(n2782) );
  NAND2X1 U2144 ( .A(n2755), .B(n2783), .Y(n423) );
  XOR2X1 U2145 ( .A(a[25]), .B(a[24]), .Y(n2755) );
  XNOR2X1 U2146 ( .A(a[24]), .B(a[23]), .Y(n2783) );
  NAND2X1 U2147 ( .A(n2756), .B(n2784), .Y(n2768) );
  XOR2X1 U2148 ( .A(a[22]), .B(a[23]), .Y(n2756) );
  XNOR2X1 U2149 ( .A(a[22]), .B(a[21]), .Y(n2784) );
  NAND2X1 U2150 ( .A(n2757), .B(n2785), .Y(n2769) );
  XOR2X1 U2151 ( .A(a[20]), .B(a[21]), .Y(n2757) );
  XNOR2X1 U2152 ( .A(a[20]), .B(a[19]), .Y(n2785) );
  NAND2X1 U2153 ( .A(n2758), .B(n2786), .Y(n2770) );
  XOR2X1 U2154 ( .A(a[18]), .B(a[19]), .Y(n2758) );
  XNOR2X1 U2155 ( .A(a[18]), .B(a[17]), .Y(n2786) );
  NAND2X1 U2156 ( .A(n2759), .B(n2787), .Y(n2771) );
  XOR2X1 U2157 ( .A(a[16]), .B(a[17]), .Y(n2759) );
  XNOR2X1 U2158 ( .A(a[16]), .B(a[15]), .Y(n2787) );
  NAND2X1 U2159 ( .A(n2760), .B(n2788), .Y(n2772) );
  XOR2X1 U2160 ( .A(a[14]), .B(a[15]), .Y(n2760) );
  XNOR2X1 U2161 ( .A(a[14]), .B(a[13]), .Y(n2788) );
  NAND2X1 U2162 ( .A(n2761), .B(n2789), .Y(n2773) );
  XOR2X1 U2163 ( .A(a[12]), .B(a[13]), .Y(n2761) );
  XNOR2X1 U2164 ( .A(a[12]), .B(a[11]), .Y(n2789) );
  NAND2X1 U2165 ( .A(n2762), .B(n2790), .Y(n2774) );
  XOR2X1 U2166 ( .A(a[10]), .B(a[11]), .Y(n2762) );
  XNOR2X1 U2167 ( .A(a[10]), .B(a[9]), .Y(n2790) );
  NAND2X1 U2168 ( .A(n2763), .B(n2791), .Y(n2775) );
  XOR2X1 U2169 ( .A(a[8]), .B(a[9]), .Y(n2763) );
  XNOR2X1 U2170 ( .A(a[8]), .B(a[7]), .Y(n2791) );
  NAND2X1 U2171 ( .A(n2764), .B(n2792), .Y(n2776) );
  XOR2X1 U2172 ( .A(a[6]), .B(a[7]), .Y(n2764) );
  XNOR2X1 U2173 ( .A(a[6]), .B(a[5]), .Y(n2792) );
  NAND2X1 U2174 ( .A(n2765), .B(n2793), .Y(n2777) );
  XOR2X1 U2175 ( .A(a[4]), .B(a[5]), .Y(n2765) );
  XNOR2X1 U2176 ( .A(a[4]), .B(a[3]), .Y(n2793) );
  NAND2X1 U2177 ( .A(n2766), .B(n2794), .Y(n2778) );
  XOR2X1 U2178 ( .A(a[2]), .B(a[3]), .Y(n2766) );
  XNOR2X1 U2179 ( .A(a[2]), .B(a[1]), .Y(n2794) );
  NAND2X1 U2180 ( .A(n2795), .B(n2767), .Y(n2779) );
  XOR2X1 U2181 ( .A(a[0]), .B(a[1]), .Y(n2767) );
  BUFX4 U2185 ( .A(n374), .Y(n2909) );
  BUFX4 U2186 ( .A(n308), .Y(n2910) );
  BUFX4 U2187 ( .A(n308), .Y(n2911) );
  BUFX2 U2188 ( .A(n296), .Y(n2912) );
  BUFX4 U2189 ( .A(n296), .Y(n2913) );
  BUFX4 U2190 ( .A(n296), .Y(n2914) );
  BUFX4 U2191 ( .A(n291), .Y(n2915) );
  BUFX4 U2192 ( .A(n291), .Y(n2916) );
  BUFX4 U2193 ( .A(n291), .Y(n2917) );
  BUFX2 U2194 ( .A(a[23]), .Y(n2813) );
  BUFX2 U2195 ( .A(a[19]), .Y(n2815) );
  BUFX2 U2196 ( .A(n2823), .Y(n291) );
  BUFX2 U2197 ( .A(n327), .Y(n2981) );
  BUFX2 U2198 ( .A(n2820), .Y(n300) );
  BUFX2 U2199 ( .A(n432), .Y(n430) );
  BUFX2 U2200 ( .A(n2812), .Y(n323) );
  BUFX2 U2201 ( .A(n2770), .Y(n412) );
  BUFX2 U2202 ( .A(n2786), .Y(n362) );
  BUFX2 U2203 ( .A(n2771), .Y(n409) );
  BUFX2 U2204 ( .A(n2776), .Y(n395) );
  BUFX2 U2205 ( .A(n2777), .Y(n392) );
  BUFX2 U2206 ( .A(n2778), .Y(n389) );
  BUFX2 U2207 ( .A(n2773), .Y(n403) );
  BUFX2 U2208 ( .A(n2779), .Y(n386) );
  BUFX2 U2209 ( .A(n2774), .Y(n400) );
  BUFX2 U2210 ( .A(n2820), .Y(n299) );
  BUFX2 U2211 ( .A(n2821), .Y(n296) );
  BUFX2 U2212 ( .A(n2769), .Y(n415) );
  BUFX2 U2213 ( .A(n2785), .Y(n365) );
  BUFX2 U2214 ( .A(n2775), .Y(n398) );
  BUFX2 U2215 ( .A(n2781), .Y(n377) );
  BUFX2 U2216 ( .A(n2772), .Y(n406) );
  BUFX2 U2217 ( .A(n2775), .Y(n397) );
  BUFX2 U2218 ( .A(a[3]), .Y(n2823) );
  BUFX2 U2219 ( .A(n2776), .Y(n396) );
  BUFX2 U2220 ( .A(n2776), .Y(n394) );
  BUFX2 U2221 ( .A(n2819), .Y(n302) );
  BUFX2 U2222 ( .A(n2822), .Y(n293) );
  BUFX2 U2223 ( .A(n2778), .Y(n388) );
  BUFX2 U2224 ( .A(n2777), .Y(n391) );
  BUFX2 U2225 ( .A(n2818), .Y(n305) );
  BUFX2 U2226 ( .A(a[17]), .Y(n2816) );
  BUFX2 U2227 ( .A(n2816), .Y(n2964) );
  BUFX2 U2228 ( .A(n2816), .Y(n2965) );
  BUFX2 U2229 ( .A(n2813), .Y(n322) );
  BUFX2 U2230 ( .A(n383), .Y(n2922) );
  BUFX2 U2231 ( .A(n2772), .Y(n408) );
  BUFX2 U2232 ( .A(n2770), .Y(n414) );
  BUFX2 U2233 ( .A(n2771), .Y(n411) );
  BUFX2 U2234 ( .A(a[15]), .Y(n2817) );
  BUFX4 U2235 ( .A(n318), .Y(n2918) );
  BUFX2 U2236 ( .A(n321), .Y(n2919) );
  BUFX2 U2237 ( .A(n321), .Y(n2920) );
  BUFX2 U2238 ( .A(n383), .Y(n2921) );
  BUFX2 U2239 ( .A(a[31]), .Y(n334) );
  OR2X2 U2240 ( .A(n1479), .B(n1456), .Y(n2923) );
  OR2X2 U2241 ( .A(n1703), .B(n1694), .Y(n2924) );
  OR2X2 U2242 ( .A(n1615), .B(n1600), .Y(n2925) );
  OR2X2 U2243 ( .A(n1741), .B(n1740), .Y(n2926) );
  OR2X2 U2244 ( .A(n1719), .B(n1712), .Y(n2927) );
  OR2X2 U2245 ( .A(n1711), .B(n1704), .Y(n2928) );
  OR2X2 U2246 ( .A(n1645), .B(n1632), .Y(n2929) );
  OR2X2 U2247 ( .A(n1455), .B(n1432), .Y(n2930) );
  OR2X2 U2248 ( .A(n920), .B(n901), .Y(n2931) );
  OR2X2 U2249 ( .A(n1501), .B(n1480), .Y(n2932) );
  OR2X2 U2250 ( .A(n1631), .B(n1616), .Y(n2933) );
  OR2X2 U2251 ( .A(n2237), .B(n2977), .Y(n2934) );
  BUFX2 U2252 ( .A(n2824), .Y(n288) );
  BUFX2 U2253 ( .A(n2821), .Y(n298) );
  BUFX2 U2254 ( .A(n2822), .Y(n294) );
  AND2X2 U2255 ( .A(n843), .B(n2978), .Y(product[1]) );
  AND2X2 U2256 ( .A(n3020), .B(n84), .Y(n2936) );
  AND2X2 U2257 ( .A(n3020), .B(n242), .Y(n2937) );
  AND2X2 U2258 ( .A(n3020), .B(n194), .Y(n2938) );
  AND2X2 U2259 ( .A(n3020), .B(n152), .Y(n2939) );
  AND2X2 U2260 ( .A(n3020), .B(n125), .Y(n2940) );
  AND2X2 U2261 ( .A(n3020), .B(n98), .Y(n2941) );
  BUFX2 U2262 ( .A(n384), .Y(n383) );
  INVX2 U2263 ( .A(n582), .Y(n580) );
  BUFX2 U2264 ( .A(n2823), .Y(n290) );
  INVX2 U2265 ( .A(n667), .Y(n665) );
  BUFX2 U2266 ( .A(n2818), .Y(n306) );
  BUFX2 U2267 ( .A(n2819), .Y(n303) );
  OR2X2 U2268 ( .A(n900), .B(n891), .Y(n2942) );
  AND2X2 U2269 ( .A(n3020), .B(n274), .Y(product[0]) );
  INVX1 U2270 ( .A(n778), .Y(n876) );
  BUFX4 U2271 ( .A(n2812), .Y(n324) );
  BUFX4 U2272 ( .A(n2814), .Y(n319) );
  XOR2X1 U2273 ( .A(n1461), .B(n1459), .Y(n2944) );
  XOR2X1 U2274 ( .A(n2944), .B(n1438), .Y(n1434) );
  XOR2X1 U2275 ( .A(n1436), .B(n1457), .Y(n2945) );
  XOR2X1 U2276 ( .A(n2945), .B(n1434), .Y(n1432) );
  NAND2X1 U2277 ( .A(n1461), .B(n1459), .Y(n2946) );
  NAND2X1 U2278 ( .A(n1461), .B(n1438), .Y(n2947) );
  NAND2X1 U2279 ( .A(n1459), .B(n1438), .Y(n2948) );
  NAND3X1 U2280 ( .A(n2946), .B(n2947), .C(n2948), .Y(n1433) );
  NAND2X1 U2281 ( .A(n1436), .B(n1457), .Y(n2949) );
  NAND2X1 U2282 ( .A(n1436), .B(n1434), .Y(n2950) );
  NAND2X1 U2283 ( .A(n1457), .B(n1434), .Y(n2951) );
  NAND3X1 U2284 ( .A(n2949), .B(n2950), .C(n2951), .Y(n1431) );
  XOR2X1 U2285 ( .A(n1874), .B(n1928), .Y(n2952) );
  XOR2X1 U2286 ( .A(n1850), .B(n2952), .Y(n1474) );
  NAND2X1 U2287 ( .A(n1850), .B(n1874), .Y(n2953) );
  NAND2X1 U2288 ( .A(n1850), .B(n1928), .Y(n2954) );
  NAND2X1 U2289 ( .A(n1874), .B(n1928), .Y(n2955) );
  NAND3X1 U2290 ( .A(n2953), .B(n2954), .C(n2955), .Y(n1473) );
  XOR2X1 U2291 ( .A(n1529), .B(n1508), .Y(n2956) );
  XOR2X1 U2292 ( .A(n2956), .B(n1527), .Y(n1504) );
  XOR2X1 U2293 ( .A(n1506), .B(n1525), .Y(n2957) );
  XOR2X1 U2294 ( .A(n2957), .B(n1504), .Y(n1502) );
  NAND2X1 U2295 ( .A(n1529), .B(n1508), .Y(n2958) );
  NAND2X1 U2296 ( .A(n1529), .B(n1527), .Y(n2959) );
  NAND2X1 U2297 ( .A(n1508), .B(n1527), .Y(n2960) );
  NAND3X1 U2298 ( .A(n2958), .B(n2959), .C(n2960), .Y(n1503) );
  NAND2X1 U2299 ( .A(n1506), .B(n1525), .Y(n2961) );
  NAND2X1 U2300 ( .A(n1506), .B(n1504), .Y(n2962) );
  NAND2X1 U2301 ( .A(n1525), .B(n1504), .Y(n2963) );
  NAND3X1 U2302 ( .A(n2961), .B(n2962), .C(n2963), .Y(n1501) );
  BUFX4 U2303 ( .A(n2815), .Y(n314) );
  BUFX2 U2304 ( .A(n2774), .Y(n402) );
  BUFX2 U2305 ( .A(n2779), .Y(n385) );
  BUFX2 U2306 ( .A(n2816), .Y(n311) );
  INVX1 U2307 ( .A(n670), .Y(n664) );
  INVX1 U2308 ( .A(n2932), .Y(n720) );
  INVX1 U2309 ( .A(n553), .Y(n551) );
  INVX1 U2310 ( .A(n623), .Y(n622) );
  INVX1 U2311 ( .A(n2933), .Y(n761) );
  INVX1 U2312 ( .A(n575), .Y(n573) );
  BUFX2 U2313 ( .A(n2814), .Y(n318) );
  BUFX2 U2314 ( .A(n2813), .Y(n321) );
  BUFX2 U2315 ( .A(n331), .Y(n330) );
  BUFX2 U2316 ( .A(n2775), .Y(n399) );
  BUFX2 U2317 ( .A(n2773), .Y(n405) );
  BUFX2 U2318 ( .A(n2779), .Y(n387) );
  BUFX2 U2319 ( .A(n2777), .Y(n393) );
  BUFX2 U2320 ( .A(n2812), .Y(n2966) );
  BUFX2 U2321 ( .A(n2812), .Y(n2967) );
  AND2X2 U2322 ( .A(n3020), .B(n143), .Y(n2970) );
  INVX1 U2323 ( .A(n364), .Y(n143) );
  AND2X2 U2324 ( .A(n3020), .B(n89), .Y(n2972) );
  INVX1 U2325 ( .A(n382), .Y(n89) );
  AND2X2 U2326 ( .A(n3020), .B(n162), .Y(n2971) );
  AND2X2 U2327 ( .A(n3020), .B(n178), .Y(n2973) );
  AND2X2 U2328 ( .A(n3020), .B(n116), .Y(n2975) );
  INVX1 U2329 ( .A(n373), .Y(n116) );
  AND2X2 U2330 ( .A(n3020), .B(n210), .Y(n2974) );
  AND2X2 U2331 ( .A(n3020), .B(n232), .Y(n2976) );
  INVX1 U2332 ( .A(n346), .Y(n232) );
  AND2X2 U2333 ( .A(n3020), .B(n258), .Y(n2977) );
  AND2X2 U2334 ( .A(n3020), .B(n134), .Y(n2979) );
  AND2X2 U2335 ( .A(n3020), .B(n107), .Y(n2980) );
  BUFX4 U2336 ( .A(a[25]), .Y(n2812) );
  INVX1 U2337 ( .A(n649), .Y(n647) );
  INVX2 U2338 ( .A(n581), .Y(n579) );
  INVX1 U2339 ( .A(n648), .Y(n646) );
  INVX1 U2340 ( .A(n631), .Y(n629) );
  INVX1 U2341 ( .A(n602), .Y(n596) );
  INVX1 U2342 ( .A(n634), .Y(n632) );
  INVX1 U2343 ( .A(n601), .Y(n599) );
  INVX1 U2344 ( .A(n669), .Y(n667) );
  XNOR2X1 U2345 ( .A(n707), .B(n2968), .Y(product[27]) );
  AND2X2 U2346 ( .A(n706), .B(n864), .Y(n2968) );
  OR2X2 U2347 ( .A(n554), .B(n581), .Y(n2969) );
  INVX1 U2348 ( .A(n718), .Y(n716) );
  INVX1 U2349 ( .A(n643), .Y(n641) );
  INVX1 U2350 ( .A(n642), .Y(n640) );
  INVX1 U2351 ( .A(n592), .Y(n590) );
  INVX2 U2352 ( .A(n725), .Y(n723) );
  INVX1 U2353 ( .A(n695), .Y(n693) );
  INVX1 U2354 ( .A(n661), .Y(n659) );
  INVX1 U2355 ( .A(n696), .Y(n694) );
  INVX1 U2356 ( .A(n593), .Y(n591) );
  INVX2 U2357 ( .A(n711), .Y(n709) );
  INVX1 U2358 ( .A(n706), .Y(n704) );
  INVX1 U2359 ( .A(n624), .Y(n623) );
  BUFX2 U2360 ( .A(n2819), .Y(n304) );
  BUFX2 U2361 ( .A(n334), .Y(n333) );
  INVX2 U2362 ( .A(n559), .Y(n557) );
  INVX1 U2363 ( .A(n759), .Y(n757) );
  INVX1 U2364 ( .A(n825), .Y(n824) );
  INVX1 U2365 ( .A(n574), .Y(n572) );
  INVX2 U2366 ( .A(n766), .Y(n764) );
  INVX1 U2367 ( .A(n783), .Y(n781) );
  INVX1 U2368 ( .A(n745), .Y(n743) );
  INVX1 U2369 ( .A(n784), .Y(n782) );
  INVX1 U2370 ( .A(n746), .Y(n744) );
  INVX1 U2371 ( .A(n774), .Y(n772) );
  BUFX2 U2372 ( .A(n2816), .Y(n312) );
  BUFX2 U2373 ( .A(n2815), .Y(n315) );
  BUFX2 U2374 ( .A(n2817), .Y(n309) );
  BUFX4 U2375 ( .A(n2821), .Y(n297) );
  BUFX2 U2376 ( .A(n2820), .Y(n301) );
  BUFX2 U2377 ( .A(n2816), .Y(n313) );
  BUFX2 U2378 ( .A(n2817), .Y(n310) );
  BUFX2 U2379 ( .A(n2823), .Y(n292) );
  BUFX2 U2380 ( .A(n2824), .Y(n289) );
  BUFX2 U2381 ( .A(n2818), .Y(n307) );
  BUFX2 U2382 ( .A(n2822), .Y(n295) );
  BUFX4 U2383 ( .A(n2813), .Y(n320) );
  BUFX4 U2384 ( .A(n2814), .Y(n317) );
  BUFX2 U2385 ( .A(n2817), .Y(n308) );
  BUFX2 U2386 ( .A(n2824), .Y(n287) );
  BUFX4 U2387 ( .A(n331), .Y(n329) );
  BUFX2 U2388 ( .A(n2815), .Y(n316) );
  INVX1 U2389 ( .A(n832), .Y(n830) );
  INVX1 U2390 ( .A(n840), .Y(n838) );
  BUFX2 U2391 ( .A(n2778), .Y(n390) );
  BUFX2 U2392 ( .A(n2771), .Y(n410) );
  BUFX2 U2393 ( .A(n2768), .Y(n419) );
  BUFX2 U2394 ( .A(n2770), .Y(n413) );
  BUFX2 U2395 ( .A(n2769), .Y(n416) );
  BUFX2 U2396 ( .A(n423), .Y(n422) );
  BUFX2 U2397 ( .A(n2787), .Y(n360) );
  BUFX2 U2398 ( .A(n2794), .Y(n339) );
  BUFX2 U2399 ( .A(n2793), .Y(n342) );
  BUFX2 U2400 ( .A(n2784), .Y(n369) );
  BUFX2 U2401 ( .A(n2785), .Y(n366) );
  BUFX2 U2402 ( .A(n2783), .Y(n372) );
  BUFX2 U2403 ( .A(n2786), .Y(n363) );
  BUFX2 U2404 ( .A(n2794), .Y(n340) );
  BUFX2 U2405 ( .A(n2793), .Y(n343) );
  BUFX2 U2406 ( .A(n2774), .Y(n401) );
  BUFX2 U2407 ( .A(n2773), .Y(n404) );
  BUFX2 U2408 ( .A(n2772), .Y(n407) );
  BUFX2 U2409 ( .A(n2790), .Y(n351) );
  BUFX2 U2410 ( .A(n2792), .Y(n345) );
  BUFX2 U2411 ( .A(n2789), .Y(n354) );
  BUFX2 U2412 ( .A(n2791), .Y(n348) );
  BUFX2 U2413 ( .A(n2788), .Y(n357) );
  BUFX2 U2414 ( .A(n2789), .Y(n355) );
  BUFX2 U2415 ( .A(n2788), .Y(n358) );
  BUFX2 U2416 ( .A(n2791), .Y(n349) );
  BUFX2 U2417 ( .A(n2790), .Y(n352) );
  BUFX2 U2418 ( .A(n2792), .Y(n346) );
  BUFX2 U2419 ( .A(n2795), .Y(n337) );
  BUFX2 U2420 ( .A(n2784), .Y(n368) );
  BUFX2 U2421 ( .A(n2783), .Y(n371) );
  BUFX2 U2422 ( .A(n2787), .Y(n359) );
  BUFX2 U2423 ( .A(n2794), .Y(n338) );
  BUFX2 U2424 ( .A(n2793), .Y(n341) );
  BUFX2 U2425 ( .A(n2795), .Y(n336) );
  BUFX2 U2426 ( .A(n2780), .Y(n380) );
  BUFX2 U2427 ( .A(n2790), .Y(n350) );
  BUFX2 U2428 ( .A(n2788), .Y(n356) );
  BUFX2 U2429 ( .A(n2789), .Y(n353) );
  BUFX2 U2430 ( .A(n2791), .Y(n347) );
  BUFX2 U2431 ( .A(n2792), .Y(n344) );
  BUFX2 U2432 ( .A(n2782), .Y(n374) );
  BUFX2 U2433 ( .A(n2787), .Y(n361) );
  BUFX2 U2434 ( .A(n2795), .Y(n335) );
  BUFX2 U2435 ( .A(n2782), .Y(n375) );
  BUFX2 U2436 ( .A(n429), .Y(n428) );
  BUFX2 U2437 ( .A(n2781), .Y(n378) );
  BUFX2 U2438 ( .A(n2786), .Y(n364) );
  INVX1 U2439 ( .A(n801), .Y(n799) );
  INVX1 U2440 ( .A(n812), .Y(n810) );
  BUFX2 U2441 ( .A(n426), .Y(n424) );
  BUFX2 U2442 ( .A(a[11]), .Y(n2819) );
  BUFX2 U2443 ( .A(n2769), .Y(n417) );
  BUFX2 U2444 ( .A(n2785), .Y(n367) );
  BUFX2 U2445 ( .A(n2812), .Y(n325) );
  BUFX2 U2446 ( .A(n2780), .Y(n381) );
  BUFX2 U2447 ( .A(n2768), .Y(n420) );
  BUFX2 U2448 ( .A(n2784), .Y(n370) );
  INVX2 U2449 ( .A(n806), .Y(n804) );
  BUFX2 U2450 ( .A(n2783), .Y(n373) );
  BUFX2 U2451 ( .A(n2781), .Y(n379) );
  BUFX2 U2452 ( .A(n2780), .Y(n382) );
  BUFX2 U2453 ( .A(a[1]), .Y(n2824) );
  BUFX2 U2454 ( .A(a[13]), .Y(n2818) );
  INVX2 U2455 ( .A(n843), .Y(n841) );
  OR2X2 U2456 ( .A(n1758), .B(n2238), .Y(n2978) );
  INVX2 U2457 ( .A(n3021), .Y(n3019) );
  INVX2 U2458 ( .A(n3014), .Y(n3013) );
  INVX2 U2459 ( .A(n3021), .Y(n3020) );
  INVX2 U2460 ( .A(n2985), .Y(n2984) );
  INVX1 U2461 ( .A(b[31]), .Y(n2985) );
  BUFX2 U2462 ( .A(b[8]), .Y(n451) );
  BUFX2 U2463 ( .A(b[4]), .Y(n443) );
  BUFX2 U2464 ( .A(b[2]), .Y(n439) );
  BUFX2 U2465 ( .A(b[14]), .Y(n463) );
  BUFX2 U2466 ( .A(b[26]), .Y(n487) );
  INVX2 U2467 ( .A(n3006), .Y(n3004) );
  INVX2 U2468 ( .A(n3003), .Y(n3002) );
  INVX2 U2469 ( .A(n3001), .Y(n3000) );
  INVX2 U2470 ( .A(n3012), .Y(n3010) );
  INVX2 U2471 ( .A(n3009), .Y(n3007) );
  INVX2 U2472 ( .A(n2997), .Y(n2996) );
  INVX2 U2473 ( .A(n2999), .Y(n2998) );
  INVX2 U2474 ( .A(n2995), .Y(n2993) );
  INVX2 U2475 ( .A(n3018), .Y(n3017) );
  INVX2 U2476 ( .A(n3016), .Y(n3015) );
  INVX2 U2477 ( .A(n2992), .Y(n2990) );
  INVX2 U2478 ( .A(n3012), .Y(n3011) );
  INVX2 U2479 ( .A(n3006), .Y(n3005) );
  INVX2 U2480 ( .A(n3009), .Y(n3008) );
  INVX1 U2481 ( .A(b[0]), .Y(n3021) );
  INVX1 U2482 ( .A(b[5]), .Y(n3014) );
  INVX2 U2483 ( .A(n2995), .Y(n2994) );
  INVX2 U2484 ( .A(n2992), .Y(n2991) );
  BUFX2 U2485 ( .A(b[6]), .Y(n447) );
  BUFX2 U2486 ( .A(b[12]), .Y(n459) );
  BUFX2 U2487 ( .A(b[28]), .Y(n491) );
  INVX2 U2488 ( .A(n2989), .Y(n2988) );
  INVX1 U2489 ( .A(b[25]), .Y(n2989) );
  INVX2 U2490 ( .A(n2987), .Y(n2986) );
  INVX1 U2491 ( .A(b[27]), .Y(n2987) );
  INVX1 U2492 ( .A(b[21]), .Y(n2995) );
  INVX1 U2493 ( .A(b[1]), .Y(n3018) );
  INVX1 U2494 ( .A(b[3]), .Y(n3016) );
  INVX1 U2495 ( .A(b[23]), .Y(n2992) );
  BUFX2 U2496 ( .A(b[10]), .Y(n455) );
  BUFX2 U2497 ( .A(b[16]), .Y(n467) );
  BUFX2 U2498 ( .A(a[7]), .Y(n2821) );
  INVX1 U2499 ( .A(b[17]), .Y(n2999) );
  INVX1 U2500 ( .A(b[7]), .Y(n3012) );
  INVX1 U2501 ( .A(b[11]), .Y(n3006) );
  INVX1 U2502 ( .A(b[13]), .Y(n3003) );
  INVX1 U2503 ( .A(b[9]), .Y(n3009) );
  INVX1 U2504 ( .A(b[15]), .Y(n3001) );
  INVX1 U2505 ( .A(b[19]), .Y(n2997) );
  BUFX4 U2506 ( .A(n327), .Y(n2982) );
  BUFX4 U2507 ( .A(n327), .Y(n2983) );
  BUFX2 U2508 ( .A(n328), .Y(n327) );
  BUFX2 U2509 ( .A(b[24]), .Y(n483) );
  BUFX2 U2510 ( .A(b[18]), .Y(n471) );
  BUFX2 U2511 ( .A(b[22]), .Y(n479) );
  BUFX2 U2512 ( .A(b[20]), .Y(n475) );
  BUFX2 U2513 ( .A(b[30]), .Y(n495) );
  INVX1 U2514 ( .A(n705), .Y(n703) );
  INVX1 U2515 ( .A(n705), .Y(n864) );
  BUFX2 U2516 ( .A(a[9]), .Y(n2820) );
  BUFX4 U2517 ( .A(n426), .Y(n425) );
  INVX2 U2518 ( .A(n727), .Y(n726) );
  BUFX4 U2519 ( .A(n328), .Y(n326) );
  INVX1 U2520 ( .A(n326), .Y(n2798) );
  BUFX2 U2521 ( .A(n432), .Y(n431) );
  BUFX2 U2522 ( .A(n2782), .Y(n376) );
  BUFX4 U2523 ( .A(a[21]), .Y(n2814) );
  BUFX2 U2524 ( .A(a[5]), .Y(n2822) );
  INVX1 U2525 ( .A(n682), .Y(n860) );
  INVX1 U2526 ( .A(n732), .Y(n868) );
  INVX1 U2527 ( .A(a[0]), .Y(n2795) );
  BUFX4 U2528 ( .A(n423), .Y(n421) );
  BUFX4 U2529 ( .A(n608), .Y(n499) );
  INVX1 U2530 ( .A(n633), .Y(n631) );
  INVX2 U2531 ( .A(n748), .Y(n747) );
  INVX1 U2532 ( .A(n650), .Y(n648) );
  INVX1 U2533 ( .A(n660), .Y(n658) );
  BUFX2 U2534 ( .A(a[29]), .Y(n331) );
  INVX1 U2535 ( .A(n808), .Y(n807) );
  INVX2 U2536 ( .A(n786), .Y(n785) );
  BUFX4 U2537 ( .A(n429), .Y(n427) );
  BUFX4 U2538 ( .A(a[27]), .Y(n328) );
  INVX2 U2539 ( .A(n768), .Y(n767) );
  INVX1 U2540 ( .A(n795), .Y(n794) );
  BUFX4 U2541 ( .A(n2768), .Y(n418) );
  INVX2 U2542 ( .A(n698), .Y(n697) );
endmodule


module poly5_DW01_sub_56 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n46, n47, n48,
         n49, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n111, n112, n113, n114, n115, n116, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n273;

  XOR2X1 U3 ( .A(n3), .B(B[47]), .Y(DIFF[47]) );
  XOR2X1 U4 ( .A(n9), .B(B[46]), .Y(DIFF[46]) );
  NAND2X1 U5 ( .A(n273), .B(n2), .Y(n3) );
  NOR2X1 U8 ( .A(n7), .B(n19), .Y(n6) );
  NAND2X1 U9 ( .A(n8), .B(n12), .Y(n7) );
  XOR2X1 U11 ( .A(n13), .B(B[45]), .Y(DIFF[45]) );
  NAND2X1 U12 ( .A(n2), .B(n10), .Y(n9) );
  NOR2X1 U13 ( .A(n11), .B(n17), .Y(n10) );
  NOR2X1 U15 ( .A(B[45]), .B(B[44]), .Y(n12) );
  XOR2X1 U16 ( .A(n15), .B(B[44]), .Y(DIFF[44]) );
  NAND2X1 U17 ( .A(n2), .B(n14), .Y(n13) );
  NOR2X1 U18 ( .A(B[44]), .B(n17), .Y(n14) );
  XOR2X1 U19 ( .A(n21), .B(B[43]), .Y(DIFF[43]) );
  NAND2X1 U20 ( .A(n16), .B(n2), .Y(n15) );
  NAND2X1 U22 ( .A(n18), .B(n32), .Y(n17) );
  NAND2X1 U24 ( .A(n20), .B(n26), .Y(n19) );
  NOR2X1 U25 ( .A(B[43]), .B(B[42]), .Y(n20) );
  XOR2X1 U26 ( .A(n23), .B(B[42]), .Y(DIFF[42]) );
  NAND2X1 U27 ( .A(n2), .B(n22), .Y(n21) );
  NOR2X1 U28 ( .A(B[42]), .B(n25), .Y(n22) );
  XOR2X1 U29 ( .A(n27), .B(B[41]), .Y(DIFF[41]) );
  NAND2X1 U30 ( .A(n24), .B(n2), .Y(n23) );
  NAND2X1 U32 ( .A(n26), .B(n32), .Y(n25) );
  NOR2X1 U33 ( .A(B[41]), .B(B[40]), .Y(n26) );
  XOR2X1 U34 ( .A(n29), .B(B[40]), .Y(DIFF[40]) );
  NAND2X1 U35 ( .A(n28), .B(n2), .Y(n27) );
  NOR2X1 U36 ( .A(B[40]), .B(n31), .Y(n28) );
  XOR2X1 U37 ( .A(n35), .B(B[39]), .Y(DIFF[39]) );
  NAND2X1 U38 ( .A(n32), .B(n2), .Y(n29) );
  NOR2X1 U41 ( .A(n33), .B(n47), .Y(n32) );
  NAND2X1 U42 ( .A(n34), .B(n40), .Y(n33) );
  NOR2X1 U43 ( .A(B[39]), .B(B[38]), .Y(n34) );
  XOR2X1 U44 ( .A(n37), .B(B[38]), .Y(DIFF[38]) );
  NAND2X1 U45 ( .A(n36), .B(n1), .Y(n35) );
  NOR2X1 U46 ( .A(B[38]), .B(n39), .Y(n36) );
  XOR2X1 U47 ( .A(n41), .B(B[37]), .Y(DIFF[37]) );
  NAND2X1 U48 ( .A(n38), .B(n1), .Y(n37) );
  NAND2X1 U50 ( .A(n40), .B(n46), .Y(n39) );
  NOR2X1 U51 ( .A(B[37]), .B(B[36]), .Y(n40) );
  XOR2X1 U52 ( .A(n43), .B(B[36]), .Y(DIFF[36]) );
  NAND2X1 U53 ( .A(n42), .B(n1), .Y(n41) );
  NOR2X1 U54 ( .A(B[36]), .B(n47), .Y(n42) );
  XOR2X1 U55 ( .A(n49), .B(B[35]), .Y(DIFF[35]) );
  NAND2X1 U56 ( .A(n46), .B(n1), .Y(n43) );
  NAND2X1 U60 ( .A(n48), .B(n54), .Y(n47) );
  NOR2X1 U61 ( .A(B[35]), .B(B[34]), .Y(n48) );
  XOR2X1 U62 ( .A(n51), .B(B[34]), .Y(DIFF[34]) );
  NAND2X1 U63 ( .A(n50), .B(n1), .Y(n49) );
  NOR2X1 U64 ( .A(B[34]), .B(n53), .Y(n50) );
  XOR2X1 U65 ( .A(n55), .B(B[33]), .Y(DIFF[33]) );
  NAND2X1 U66 ( .A(n54), .B(n1), .Y(n51) );
  NOR2X1 U69 ( .A(B[33]), .B(B[32]), .Y(n54) );
  XNOR2X1 U70 ( .A(n1), .B(B[32]), .Y(DIFF[32]) );
  NAND2X1 U71 ( .A(n56), .B(n1), .Y(n55) );
  XOR2X1 U73 ( .A(n62), .B(B[31]), .Y(DIFF[31]) );
  NOR2X1 U74 ( .A(n123), .B(n58), .Y(n57) );
  NAND2X1 U75 ( .A(n59), .B(n97), .Y(n58) );
  NOR2X1 U76 ( .A(n60), .B(n80), .Y(n59) );
  NAND2X1 U77 ( .A(n61), .B(n71), .Y(n60) );
  NOR2X1 U78 ( .A(B[31]), .B(B[30]), .Y(n61) );
  XOR2X1 U79 ( .A(n66), .B(B[30]), .Y(DIFF[30]) );
  NAND2X1 U80 ( .A(n122), .B(n63), .Y(n62) );
  NOR2X1 U81 ( .A(n64), .B(n96), .Y(n63) );
  NAND2X1 U82 ( .A(n79), .B(n65), .Y(n64) );
  NOR2X1 U83 ( .A(B[30]), .B(n70), .Y(n65) );
  XOR2X1 U84 ( .A(n72), .B(B[29]), .Y(DIFF[29]) );
  NAND2X1 U85 ( .A(n122), .B(n67), .Y(n66) );
  NOR2X1 U86 ( .A(n68), .B(n96), .Y(n67) );
  NAND2X1 U87 ( .A(n69), .B(n79), .Y(n68) );
  NOR2X1 U90 ( .A(B[29]), .B(B[28]), .Y(n71) );
  XOR2X1 U91 ( .A(n76), .B(B[28]), .Y(DIFF[28]) );
  NAND2X1 U92 ( .A(n122), .B(n73), .Y(n72) );
  NOR2X1 U93 ( .A(n74), .B(n96), .Y(n73) );
  NAND2X1 U94 ( .A(n75), .B(n79), .Y(n74) );
  XOR2X1 U96 ( .A(n82), .B(B[27]), .Y(DIFF[27]) );
  NAND2X1 U97 ( .A(n122), .B(n77), .Y(n76) );
  NOR2X1 U98 ( .A(n78), .B(n96), .Y(n77) );
  NAND2X1 U101 ( .A(n81), .B(n91), .Y(n80) );
  NOR2X1 U102 ( .A(B[27]), .B(B[26]), .Y(n81) );
  XOR2X1 U103 ( .A(n86), .B(B[26]), .Y(DIFF[26]) );
  NAND2X1 U104 ( .A(n122), .B(n83), .Y(n82) );
  NOR2X1 U105 ( .A(n84), .B(n96), .Y(n83) );
  NAND2X1 U106 ( .A(n85), .B(n91), .Y(n84) );
  XOR2X1 U108 ( .A(n92), .B(B[25]), .Y(DIFF[25]) );
  NAND2X1 U109 ( .A(n122), .B(n87), .Y(n86) );
  NOR2X1 U110 ( .A(n90), .B(n96), .Y(n87) );
  NOR2X1 U114 ( .A(B[25]), .B(B[24]), .Y(n91) );
  XOR2X1 U115 ( .A(n94), .B(B[24]), .Y(DIFF[24]) );
  NAND2X1 U116 ( .A(n122), .B(n93), .Y(n92) );
  NOR2X1 U117 ( .A(B[24]), .B(n96), .Y(n93) );
  XOR2X1 U118 ( .A(n100), .B(B[23]), .Y(DIFF[23]) );
  NAND2X1 U119 ( .A(n95), .B(n122), .Y(n94) );
  NOR2X1 U122 ( .A(n98), .B(n112), .Y(n97) );
  NAND2X1 U123 ( .A(n99), .B(n105), .Y(n98) );
  NOR2X1 U124 ( .A(B[23]), .B(B[22]), .Y(n99) );
  XOR2X1 U125 ( .A(n102), .B(B[22]), .Y(DIFF[22]) );
  NAND2X1 U126 ( .A(n122), .B(n101), .Y(n100) );
  NOR2X1 U127 ( .A(B[22]), .B(n104), .Y(n101) );
  XOR2X1 U128 ( .A(n106), .B(B[21]), .Y(DIFF[21]) );
  NAND2X1 U129 ( .A(n103), .B(n122), .Y(n102) );
  NAND2X1 U131 ( .A(n105), .B(n111), .Y(n104) );
  NOR2X1 U132 ( .A(B[21]), .B(B[20]), .Y(n105) );
  XOR2X1 U133 ( .A(n108), .B(B[20]), .Y(DIFF[20]) );
  NAND2X1 U134 ( .A(n107), .B(n122), .Y(n106) );
  NOR2X1 U135 ( .A(B[20]), .B(n112), .Y(n107) );
  XOR2X1 U136 ( .A(n114), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U137 ( .A(n111), .B(n122), .Y(n108) );
  NAND2X1 U141 ( .A(n113), .B(n119), .Y(n112) );
  NOR2X1 U142 ( .A(B[19]), .B(B[18]), .Y(n113) );
  XOR2X1 U143 ( .A(n116), .B(B[18]), .Y(DIFF[18]) );
  NAND2X1 U144 ( .A(n115), .B(n122), .Y(n114) );
  NOR2X1 U145 ( .A(B[18]), .B(n118), .Y(n115) );
  XOR2X1 U146 ( .A(n120), .B(B[17]), .Y(DIFF[17]) );
  NAND2X1 U147 ( .A(n119), .B(n122), .Y(n116) );
  NOR2X1 U150 ( .A(B[17]), .B(B[16]), .Y(n119) );
  XNOR2X1 U151 ( .A(n122), .B(B[16]), .Y(DIFF[16]) );
  NAND2X1 U152 ( .A(n121), .B(n122), .Y(n120) );
  INVX4 U154 ( .A(n123), .Y(n122) );
  NAND2X1 U155 ( .A(n131), .B(n124), .Y(n123) );
  NOR2X1 U156 ( .A(n125), .B(n128), .Y(n124) );
  NAND2X1 U157 ( .A(n126), .B(n127), .Y(n125) );
  NOR2X1 U158 ( .A(B[15]), .B(B[14]), .Y(n126) );
  NOR2X1 U159 ( .A(B[13]), .B(B[12]), .Y(n127) );
  NAND2X1 U160 ( .A(n129), .B(n130), .Y(n128) );
  NOR2X1 U161 ( .A(B[11]), .B(B[10]), .Y(n129) );
  NOR2X1 U162 ( .A(B[9]), .B(B[8]), .Y(n130) );
  NOR2X1 U163 ( .A(n135), .B(n132), .Y(n131) );
  NAND2X1 U164 ( .A(n133), .B(n134), .Y(n132) );
  NOR2X1 U165 ( .A(B[7]), .B(B[6]), .Y(n133) );
  NOR2X1 U166 ( .A(B[5]), .B(B[4]), .Y(n134) );
  NAND2X1 U167 ( .A(n137), .B(n136), .Y(n135) );
  NOR2X1 U168 ( .A(B[3]), .B(B[2]), .Y(n136) );
  NOR2X1 U169 ( .A(B[0]), .B(B[1]), .Y(n137) );
  INVX2 U173 ( .A(n97), .Y(n96) );
  INVX1 U174 ( .A(n47), .Y(n46) );
  AND2X2 U175 ( .A(n6), .B(n32), .Y(n273) );
  INVX2 U176 ( .A(n119), .Y(n118) );
  INVX2 U177 ( .A(n32), .Y(n31) );
  INVX1 U178 ( .A(n54), .Y(n53) );
  INVX2 U179 ( .A(n91), .Y(n90) );
  INVX2 U180 ( .A(n112), .Y(n111) );
  INVX1 U181 ( .A(B[28]), .Y(n75) );
  INVX1 U182 ( .A(B[26]), .Y(n85) );
  INVX1 U183 ( .A(n12), .Y(n11) );
  INVX1 U184 ( .A(B[46]), .Y(n8) );
  BUFX2 U185 ( .A(n57), .Y(n2) );
  INVX2 U186 ( .A(n96), .Y(n95) );
  INVX1 U187 ( .A(n25), .Y(n24) );
  INVX1 U188 ( .A(B[16]), .Y(n121) );
  INVX1 U189 ( .A(B[32]), .Y(n56) );
  INVX1 U190 ( .A(n70), .Y(n69) );
  INVX1 U191 ( .A(n39), .Y(n38) );
  INVX1 U192 ( .A(n79), .Y(n78) );
  INVX2 U193 ( .A(n80), .Y(n79) );
  INVX2 U194 ( .A(n71), .Y(n70) );
  INVX1 U195 ( .A(n17), .Y(n16) );
  INVX1 U196 ( .A(n19), .Y(n18) );
  INVX1 U197 ( .A(n104), .Y(n103) );
  BUFX4 U198 ( .A(n57), .Y(n1) );
endmodule


module poly5_DW_mult_uns_43 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n8, n13, n18, n23, n28, n33, n38, n68, n80, n85, n89, n98, n107, n116,
         n125, n134, n143, n152, n162, n163, n178, n179, n194, n195, n201,
         n210, n211, n226, n227, n242, n243, n249, n258, n259, n275, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n437, n439, n441, n443, n445, n447, n449, n451, n453,
         n455, n457, n459, n461, n463, n465, n467, n469, n471, n473, n475,
         n477, n479, n481, n483, n485, n489, n491, n493, n495, n497, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n548, n549, n551, n553, n554, n555, n557, n559, n560,
         n561, n562, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n596, n599, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n709, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n723, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n764, n766, n767,
         n768, n769, n770, n772, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n799, n801, n802, n804, n806,
         n807, n808, n810, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n830, n832,
         n833, n834, n835, n836, n838, n840, n841, n843, n846, n848, n850,
         n851, n852, n854, n856, n858, n859, n860, n861, n862, n868, n869,
         n870, n872, n876, n878, n879, n883, n884, n885, n886, n888, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953;

  NAND2X1 OR_NOTi ( .A(n2953), .B(n289), .Y(n2725) );
  INVX2 U21 ( .A(n387), .Y(n275) );
  OAI21X1 AO21i ( .A(a[0]), .B(n275), .C(n287), .Y(n2206) );
  NAND2X1 OR_NOTi1 ( .A(n2953), .B(n292), .Y(n2692) );
  INVX2 U23 ( .A(n390), .Y(n259) );
  INVX2 U15 ( .A(n340), .Y(n258) );
  OAI21X1 AO21i1 ( .A(n258), .B(n259), .C(n290), .Y(n2172) );
  NAND2X1 OR_NOTi2 ( .A(n2953), .B(n295), .Y(n2659) );
  INVX2 U24 ( .A(n249), .Y(n2171) );
  NAND2X1 AND_NOTi2 ( .A(n2951), .B(n242), .Y(n249) );
  INVX2 U25 ( .A(n393), .Y(n243) );
  INVX2 U18 ( .A(n343), .Y(n242) );
  OAI21X1 AO21i2 ( .A(n242), .B(n243), .C(n293), .Y(n2138) );
  NAND2X1 OR_NOTi3 ( .A(n2953), .B(n298), .Y(n2626) );
  INVX2 U27 ( .A(n396), .Y(n227) );
  INVX2 U111 ( .A(n346), .Y(n226) );
  OAI21X1 AO21i3 ( .A(n226), .B(n227), .C(n298), .Y(n2104) );
  NAND2X1 OR_NOTi4 ( .A(n2953), .B(n301), .Y(n2593) );
  INVX2 U29 ( .A(n399), .Y(n211) );
  INVX2 U114 ( .A(n349), .Y(n210) );
  OAI21X1 AO21i4 ( .A(n210), .B(n211), .C(n299), .Y(n2070) );
  NAND2X1 OR_NOTi5 ( .A(n2953), .B(n304), .Y(n2560) );
  INVX2 U210 ( .A(n201), .Y(n2069) );
  NAND2X1 AND_NOTi5 ( .A(n2951), .B(n194), .Y(n201) );
  INVX2 U211 ( .A(n402), .Y(n195) );
  INVX2 U117 ( .A(n352), .Y(n194) );
  OAI21X1 AO21i5 ( .A(n194), .B(n195), .C(n304), .Y(n2036) );
  NAND2X1 OR_NOTi6 ( .A(n2953), .B(n307), .Y(n2527) );
  INVX2 U213 ( .A(n405), .Y(n179) );
  INVX2 U120 ( .A(n355), .Y(n178) );
  OAI21X1 AO21i6 ( .A(n178), .B(n179), .C(n307), .Y(n2002) );
  NAND2X1 OR_NOTi7 ( .A(n2953), .B(n310), .Y(n2494) );
  INVX2 U215 ( .A(n408), .Y(n163) );
  INVX2 U123 ( .A(n358), .Y(n162) );
  OAI21X1 AO21i7 ( .A(n162), .B(n163), .C(n310), .Y(n1968) );
  NAND2X1 OR_NOTi8 ( .A(n2953), .B(n313), .Y(n2461) );
  INVX2 U125 ( .A(n361), .Y(n152) );
  NAND2X1 OR_NOTi9 ( .A(n2953), .B(n316), .Y(n2428) );
  INVX2 U127 ( .A(n364), .Y(n143) );
  NAND2X1 OR_NOTi10 ( .A(n2952), .B(n319), .Y(n2397) );
  INVX2 U129 ( .A(n367), .Y(n134) );
  NAND2X1 OR_NOTi11 ( .A(n2952), .B(n322), .Y(n2368) );
  INVX2 U131 ( .A(n370), .Y(n125) );
  NAND2X1 OR_NOTi12 ( .A(n2952), .B(n325), .Y(n2341) );
  INVX2 U133 ( .A(n373), .Y(n116) );
  NAND2X1 OR_NOTi13 ( .A(n2952), .B(n328), .Y(n2316) );
  INVX2 U135 ( .A(n376), .Y(n107) );
  NAND2X1 OR_NOTi14 ( .A(n2952), .B(n331), .Y(n2293) );
  INVX2 U137 ( .A(n379), .Y(n98) );
  NAND2X1 OR_NOTi15 ( .A(n2952), .B(n334), .Y(n2272) );
  INVX2 U139 ( .A(n382), .Y(n89) );
  INVX2 U224 ( .A(n85), .Y(n1767) );
  NAND2X1 AND_NOTi16 ( .A(n2951), .B(n333), .Y(n85) );
  XOR2X1 U225 ( .A(n1759), .B(n918), .Y(n80) );
  XOR2X1 U141 ( .A(n1852), .B(n80), .Y(n899) );
  XOR2X1 U226 ( .A(n1768), .B(n1828), .Y(n68) );
  XOR2X1 U142 ( .A(n1786), .B(n68), .Y(n898) );
  XOR2X1 U227 ( .A(n1906), .B(n1806), .Y(n38) );
  XOR2X1 U143 ( .A(n1878), .B(n38), .Y(n897) );
  XOR2X1 U228 ( .A(n1968), .B(n1936), .Y(n33) );
  XOR2X1 U144 ( .A(n899), .B(n33), .Y(n896) );
  XOR2X1 U229 ( .A(n914), .B(n916), .Y(n28) );
  XOR2X1 U145 ( .A(n912), .B(n28), .Y(n895) );
  XOR2X1 U230 ( .A(n898), .B(n897), .Y(n23) );
  XOR2X1 U146 ( .A(n910), .B(n23), .Y(n894) );
  XOR2X1 U231 ( .A(n908), .B(n896), .Y(n18) );
  XOR2X1 U147 ( .A(n895), .B(n18), .Y(n893) );
  XOR2X1 U232 ( .A(n894), .B(n906), .Y(n13) );
  XOR2X1 U148 ( .A(n904), .B(n13), .Y(n892) );
  XOR2X1 U233 ( .A(n902), .B(n893), .Y(n8) );
  XOR2X1 U149 ( .A(n892), .B(n8), .Y(n891) );
  XNOR2X1 U292 ( .A(n549), .B(n500), .Y(product[47]) );
  NAND2X1 U293 ( .A(n548), .B(n2932), .Y(n500) );
  NAND2X1 U296 ( .A(n900), .B(n891), .Y(n548) );
  XNOR2X1 U297 ( .A(n560), .B(n501), .Y(product[46]) );
  OAI21X1 U298 ( .A(n2934), .B(n499), .C(n551), .Y(n549) );
  OAI21X1 U302 ( .A(n554), .B(n582), .C(n555), .Y(n553) );
  NAND2X1 U303 ( .A(n2928), .B(n565), .Y(n554) );
  AOI21X1 U304 ( .A(n2928), .B(n566), .C(n557), .Y(n555) );
  NAND2X1 U307 ( .A(n559), .B(n2928), .Y(n501) );
  NAND2X1 U310 ( .A(n920), .B(n901), .Y(n559) );
  XNOR2X1 U311 ( .A(n569), .B(n502), .Y(product[45]) );
  OAI21X1 U312 ( .A(n561), .B(n499), .C(n562), .Y(n560) );
  NAND2X1 U313 ( .A(n565), .B(n579), .Y(n561) );
  AOI21X1 U314 ( .A(n565), .B(n580), .C(n566), .Y(n562) );
  NOR2X1 U317 ( .A(n567), .B(n574), .Y(n565) );
  OAI21X1 U318 ( .A(n567), .B(n575), .C(n568), .Y(n566) );
  NAND2X1 U319 ( .A(n568), .B(n846), .Y(n502) );
  INVX2 U320 ( .A(n567), .Y(n846) );
  NOR2X1 U321 ( .A(n921), .B(n940), .Y(n567) );
  NAND2X1 U322 ( .A(n921), .B(n940), .Y(n568) );
  XNOR2X1 U323 ( .A(n576), .B(n503), .Y(product[44]) );
  OAI21X1 U324 ( .A(n570), .B(n499), .C(n571), .Y(n569) );
  NAND2X1 U325 ( .A(n572), .B(n579), .Y(n570) );
  AOI21X1 U326 ( .A(n572), .B(n580), .C(n573), .Y(n571) );
  NAND2X1 U329 ( .A(n575), .B(n572), .Y(n503) );
  NOR2X1 U331 ( .A(n962), .B(n941), .Y(n574) );
  NAND2X1 U332 ( .A(n962), .B(n941), .Y(n575) );
  XNOR2X1 U333 ( .A(n587), .B(n504), .Y(product[43]) );
  OAI21X1 U334 ( .A(n581), .B(n499), .C(n582), .Y(n576) );
  NAND2X1 U339 ( .A(n583), .B(n601), .Y(n581) );
  AOI21X1 U340 ( .A(n583), .B(n602), .C(n584), .Y(n582) );
  NOR2X1 U341 ( .A(n585), .B(n592), .Y(n583) );
  OAI21X1 U342 ( .A(n593), .B(n585), .C(n586), .Y(n584) );
  NAND2X1 U343 ( .A(n586), .B(n848), .Y(n504) );
  INVX2 U344 ( .A(n585), .Y(n848) );
  NOR2X1 U345 ( .A(n984), .B(n963), .Y(n585) );
  NAND2X1 U346 ( .A(n984), .B(n963), .Y(n586) );
  XNOR2X1 U347 ( .A(n594), .B(n505), .Y(product[42]) );
  OAI21X1 U348 ( .A(n588), .B(n499), .C(n589), .Y(n587) );
  NAND2X1 U349 ( .A(n590), .B(n601), .Y(n588) );
  AOI21X1 U350 ( .A(n590), .B(n602), .C(n591), .Y(n589) );
  NAND2X1 U353 ( .A(n593), .B(n590), .Y(n505) );
  NOR2X1 U355 ( .A(n1008), .B(n985), .Y(n592) );
  NAND2X1 U356 ( .A(n1008), .B(n985), .Y(n593) );
  XNOR2X1 U357 ( .A(n605), .B(n506), .Y(product[41]) );
  OAI21X1 U358 ( .A(n599), .B(n499), .C(n596), .Y(n594) );
  NOR2X1 U365 ( .A(n603), .B(n606), .Y(n601) );
  OAI21X1 U366 ( .A(n607), .B(n603), .C(n604), .Y(n602) );
  NAND2X1 U367 ( .A(n604), .B(n850), .Y(n506) );
  INVX2 U368 ( .A(n603), .Y(n850) );
  NOR2X1 U369 ( .A(n1032), .B(n1009), .Y(n603) );
  NAND2X1 U370 ( .A(n1032), .B(n1009), .Y(n604) );
  XOR2X1 U371 ( .A(n499), .B(n507), .Y(product[40]) );
  OAI21X1 U372 ( .A(n606), .B(n499), .C(n607), .Y(n605) );
  NAND2X1 U373 ( .A(n607), .B(n851), .Y(n507) );
  INVX2 U374 ( .A(n606), .Y(n851) );
  NOR2X1 U375 ( .A(n1058), .B(n1033), .Y(n606) );
  NAND2X1 U376 ( .A(n1058), .B(n1033), .Y(n607) );
  XNOR2X1 U377 ( .A(n617), .B(n508), .Y(product[39]) );
  AOI21X1 U378 ( .A(n677), .B(n609), .C(n610), .Y(n608) );
  NOR2X1 U379 ( .A(n649), .B(n611), .Y(n609) );
  OAI21X1 U380 ( .A(n611), .B(n650), .C(n612), .Y(n610) );
  NAND2X1 U381 ( .A(n613), .B(n633), .Y(n611) );
  AOI21X1 U382 ( .A(n634), .B(n613), .C(n614), .Y(n612) );
  NOR2X1 U383 ( .A(n615), .B(n624), .Y(n613) );
  OAI21X1 U384 ( .A(n625), .B(n615), .C(n616), .Y(n614) );
  NAND2X1 U385 ( .A(n616), .B(n852), .Y(n508) );
  INVX2 U386 ( .A(n615), .Y(n852) );
  NOR2X1 U387 ( .A(n1084), .B(n1059), .Y(n615) );
  NAND2X1 U388 ( .A(n1084), .B(n1059), .Y(n616) );
  XNOR2X1 U389 ( .A(n626), .B(n509), .Y(product[38]) );
  OAI21X1 U390 ( .A(n676), .B(n618), .C(n619), .Y(n617) );
  NAND2X1 U391 ( .A(n647), .B(n620), .Y(n618) );
  AOI21X1 U392 ( .A(n648), .B(n620), .C(n621), .Y(n619) );
  NOR2X1 U393 ( .A(n622), .B(n631), .Y(n620) );
  OAI21X1 U394 ( .A(n622), .B(n632), .C(n625), .Y(n621) );
  NAND2X1 U397 ( .A(n625), .B(n623), .Y(n509) );
  NOR2X1 U399 ( .A(n1112), .B(n1085), .Y(n624) );
  NAND2X1 U400 ( .A(n1112), .B(n1085), .Y(n625) );
  XNOR2X1 U401 ( .A(n637), .B(n510), .Y(product[37]) );
  OAI21X1 U402 ( .A(n676), .B(n627), .C(n628), .Y(n626) );
  NAND2X1 U403 ( .A(n629), .B(n647), .Y(n627) );
  AOI21X1 U404 ( .A(n629), .B(n648), .C(n634), .Y(n628) );
  NOR2X1 U409 ( .A(n635), .B(n642), .Y(n633) );
  OAI21X1 U410 ( .A(n643), .B(n635), .C(n636), .Y(n634) );
  NAND2X1 U411 ( .A(n636), .B(n854), .Y(n510) );
  INVX2 U412 ( .A(n635), .Y(n854) );
  NOR2X1 U413 ( .A(n1140), .B(n1113), .Y(n635) );
  NAND2X1 U414 ( .A(n1140), .B(n1113), .Y(n636) );
  XNOR2X1 U415 ( .A(n644), .B(n511), .Y(product[36]) );
  OAI21X1 U416 ( .A(n676), .B(n638), .C(n639), .Y(n637) );
  NAND2X1 U417 ( .A(n640), .B(n647), .Y(n638) );
  AOI21X1 U418 ( .A(n640), .B(n648), .C(n641), .Y(n639) );
  NAND2X1 U421 ( .A(n643), .B(n640), .Y(n511) );
  NOR2X1 U423 ( .A(n1170), .B(n1141), .Y(n642) );
  NAND2X1 U424 ( .A(n1170), .B(n1141), .Y(n643) );
  XNOR2X1 U425 ( .A(n655), .B(n512), .Y(product[35]) );
  OAI21X1 U426 ( .A(n649), .B(n676), .C(n650), .Y(n644) );
  NAND2X1 U431 ( .A(n669), .B(n651), .Y(n649) );
  AOI21X1 U432 ( .A(n670), .B(n651), .C(n652), .Y(n650) );
  NOR2X1 U433 ( .A(n653), .B(n660), .Y(n651) );
  OAI21X1 U434 ( .A(n661), .B(n653), .C(n654), .Y(n652) );
  NAND2X1 U435 ( .A(n654), .B(n856), .Y(n512) );
  INVX2 U436 ( .A(n653), .Y(n856) );
  NOR2X1 U437 ( .A(n1200), .B(n1171), .Y(n653) );
  NAND2X1 U438 ( .A(n1200), .B(n1171), .Y(n654) );
  XNOR2X1 U439 ( .A(n662), .B(n513), .Y(product[34]) );
  OAI21X1 U440 ( .A(n656), .B(n676), .C(n657), .Y(n655) );
  NAND2X1 U441 ( .A(n658), .B(n665), .Y(n656) );
  AOI21X1 U442 ( .A(n658), .B(n666), .C(n659), .Y(n657) );
  NAND2X1 U445 ( .A(n661), .B(n658), .Y(n513) );
  NOR2X1 U447 ( .A(n1232), .B(n1201), .Y(n660) );
  NAND2X1 U448 ( .A(n1232), .B(n1201), .Y(n661) );
  XNOR2X1 U449 ( .A(n673), .B(n514), .Y(product[33]) );
  OAI21X1 U450 ( .A(n667), .B(n676), .C(n664), .Y(n662) );
  NOR2X1 U457 ( .A(n674), .B(n671), .Y(n669) );
  OAI21X1 U458 ( .A(n675), .B(n671), .C(n672), .Y(n670) );
  NAND2X1 U459 ( .A(n672), .B(n858), .Y(n514) );
  NOR2X1 U461 ( .A(n1263), .B(n1233), .Y(n671) );
  NAND2X1 U462 ( .A(n1263), .B(n1233), .Y(n672) );
  XOR2X1 U463 ( .A(n676), .B(n515), .Y(product[32]) );
  OAI21X1 U464 ( .A(n674), .B(n676), .C(n675), .Y(n673) );
  NAND2X1 U465 ( .A(n675), .B(n859), .Y(n515) );
  INVX2 U466 ( .A(n674), .Y(n859) );
  NOR2X1 U467 ( .A(n1293), .B(n1264), .Y(n674) );
  NAND2X1 U468 ( .A(n1293), .B(n1264), .Y(n675) );
  XNOR2X1 U469 ( .A(n684), .B(n516), .Y(product[31]) );
  INVX4 U470 ( .A(n677), .Y(n676) );
  OAI21X1 U471 ( .A(n698), .B(n678), .C(n679), .Y(n677) );
  NAND2X1 U472 ( .A(n688), .B(n680), .Y(n678) );
  AOI21X1 U473 ( .A(n689), .B(n680), .C(n681), .Y(n679) );
  NOR2X1 U474 ( .A(n685), .B(n682), .Y(n680) );
  OAI21X1 U475 ( .A(n686), .B(n682), .C(n683), .Y(n681) );
  NAND2X1 U476 ( .A(n683), .B(n860), .Y(n516) );
  NOR2X1 U478 ( .A(n1323), .B(n1294), .Y(n682) );
  NAND2X1 U479 ( .A(n1323), .B(n1294), .Y(n683) );
  XOR2X1 U480 ( .A(n687), .B(n517), .Y(product[30]) );
  OAI21X1 U481 ( .A(n685), .B(n687), .C(n686), .Y(n684) );
  NAND2X1 U482 ( .A(n686), .B(n861), .Y(n517) );
  INVX2 U483 ( .A(n685), .Y(n861) );
  NOR2X1 U484 ( .A(n1351), .B(n1324), .Y(n685) );
  NAND2X1 U485 ( .A(n1351), .B(n1324), .Y(n686) );
  XOR2X1 U486 ( .A(n692), .B(n518), .Y(product[29]) );
  AOI21X1 U487 ( .A(n688), .B(n697), .C(n689), .Y(n687) );
  NOR2X1 U488 ( .A(n695), .B(n690), .Y(n688) );
  OAI21X1 U489 ( .A(n696), .B(n690), .C(n691), .Y(n689) );
  NAND2X1 U490 ( .A(n691), .B(n862), .Y(n518) );
  INVX2 U491 ( .A(n690), .Y(n862) );
  NOR2X1 U492 ( .A(n1379), .B(n1352), .Y(n690) );
  NAND2X1 U493 ( .A(n1379), .B(n1352), .Y(n691) );
  XNOR2X1 U494 ( .A(n697), .B(n519), .Y(product[28]) );
  AOI21X1 U495 ( .A(n693), .B(n697), .C(n694), .Y(n692) );
  NAND2X1 U498 ( .A(n696), .B(n693), .Y(n519) );
  NOR2X1 U500 ( .A(n1405), .B(n1380), .Y(n695) );
  NAND2X1 U501 ( .A(n1405), .B(n1380), .Y(n696) );
  XOR2X1 U502 ( .A(n707), .B(n520), .Y(product[27]) );
  AOI21X1 U504 ( .A(n699), .B(n727), .C(n700), .Y(n698) );
  NOR2X1 U505 ( .A(n713), .B(n701), .Y(n699) );
  OAI21X1 U506 ( .A(n714), .B(n701), .C(n702), .Y(n700) );
  NAND2X1 U507 ( .A(n2924), .B(n703), .Y(n701) );
  AOI21X1 U508 ( .A(n709), .B(n703), .C(n704), .Y(n702) );
  NAND2X1 U511 ( .A(n706), .B(n703), .Y(n520) );
  NOR2X1 U513 ( .A(n1431), .B(n1406), .Y(n705) );
  NAND2X1 U514 ( .A(n1431), .B(n1406), .Y(n706) );
  XNOR2X1 U515 ( .A(n712), .B(n521), .Y(product[26]) );
  AOI21X1 U516 ( .A(n2924), .B(n712), .C(n709), .Y(n707) );
  NAND2X1 U519 ( .A(n711), .B(n2924), .Y(n521) );
  NAND2X1 U522 ( .A(n1455), .B(n1432), .Y(n711) );
  XNOR2X1 U523 ( .A(n719), .B(n522), .Y(product[25]) );
  OAI21X1 U524 ( .A(n713), .B(n726), .C(n714), .Y(n712) );
  NAND2X1 U525 ( .A(n2926), .B(n715), .Y(n713) );
  AOI21X1 U526 ( .A(n723), .B(n715), .C(n716), .Y(n714) );
  NAND2X1 U529 ( .A(n718), .B(n715), .Y(n522) );
  NOR2X1 U531 ( .A(n1479), .B(n1456), .Y(n717) );
  NAND2X1 U532 ( .A(n1479), .B(n1456), .Y(n718) );
  XOR2X1 U533 ( .A(n726), .B(n523), .Y(product[24]) );
  OAI21X1 U534 ( .A(n720), .B(n726), .C(n725), .Y(n719) );
  NAND2X1 U539 ( .A(n725), .B(n2926), .Y(n523) );
  NAND2X1 U542 ( .A(n1501), .B(n1480), .Y(n725) );
  XNOR2X1 U543 ( .A(n734), .B(n524), .Y(product[23]) );
  OAI21X1 U545 ( .A(n748), .B(n728), .C(n729), .Y(n727) );
  NAND2X1 U546 ( .A(n738), .B(n730), .Y(n728) );
  AOI21X1 U547 ( .A(n739), .B(n730), .C(n731), .Y(n729) );
  NOR2X1 U548 ( .A(n735), .B(n732), .Y(n730) );
  OAI21X1 U549 ( .A(n736), .B(n732), .C(n733), .Y(n731) );
  NAND2X1 U550 ( .A(n733), .B(n868), .Y(n524) );
  INVX2 U551 ( .A(n732), .Y(n868) );
  NOR2X1 U552 ( .A(n1523), .B(n1502), .Y(n732) );
  NAND2X1 U553 ( .A(n1523), .B(n1502), .Y(n733) );
  XOR2X1 U554 ( .A(n737), .B(n525), .Y(product[22]) );
  OAI21X1 U555 ( .A(n735), .B(n737), .C(n736), .Y(n734) );
  NAND2X1 U556 ( .A(n736), .B(n869), .Y(n525) );
  INVX2 U557 ( .A(n735), .Y(n869) );
  NOR2X1 U558 ( .A(n1543), .B(n1524), .Y(n735) );
  NAND2X1 U559 ( .A(n1543), .B(n1524), .Y(n736) );
  XOR2X1 U560 ( .A(n742), .B(n526), .Y(product[21]) );
  AOI21X1 U561 ( .A(n738), .B(n747), .C(n739), .Y(n737) );
  NOR2X1 U562 ( .A(n745), .B(n740), .Y(n738) );
  OAI21X1 U563 ( .A(n746), .B(n740), .C(n741), .Y(n739) );
  NAND2X1 U564 ( .A(n741), .B(n870), .Y(n526) );
  INVX2 U565 ( .A(n740), .Y(n870) );
  NOR2X1 U566 ( .A(n1563), .B(n1544), .Y(n740) );
  NAND2X1 U567 ( .A(n1563), .B(n1544), .Y(n741) );
  XNOR2X1 U568 ( .A(n747), .B(n527), .Y(product[20]) );
  AOI21X1 U569 ( .A(n743), .B(n747), .C(n744), .Y(n742) );
  NAND2X1 U572 ( .A(n746), .B(n743), .Y(n527) );
  NOR2X1 U574 ( .A(n1581), .B(n1564), .Y(n745) );
  NAND2X1 U575 ( .A(n1581), .B(n1564), .Y(n746) );
  XNOR2X1 U576 ( .A(n753), .B(n528), .Y(product[19]) );
  AOI21X1 U578 ( .A(n749), .B(n768), .C(n750), .Y(n748) );
  NOR2X1 U579 ( .A(n751), .B(n754), .Y(n749) );
  OAI21X1 U580 ( .A(n751), .B(n755), .C(n752), .Y(n750) );
  NAND2X1 U581 ( .A(n752), .B(n872), .Y(n528) );
  INVX2 U582 ( .A(n751), .Y(n872) );
  NOR2X1 U583 ( .A(n1599), .B(n1582), .Y(n751) );
  NAND2X1 U584 ( .A(n1599), .B(n1582), .Y(n752) );
  XNOR2X1 U585 ( .A(n760), .B(n529), .Y(product[18]) );
  OAI21X1 U586 ( .A(n754), .B(n767), .C(n755), .Y(n753) );
  NAND2X1 U587 ( .A(n2925), .B(n756), .Y(n754) );
  AOI21X1 U588 ( .A(n764), .B(n756), .C(n757), .Y(n755) );
  NAND2X1 U591 ( .A(n759), .B(n756), .Y(n529) );
  NOR2X1 U593 ( .A(n1615), .B(n1600), .Y(n758) );
  NAND2X1 U594 ( .A(n1615), .B(n1600), .Y(n759) );
  XOR2X1 U595 ( .A(n767), .B(n530), .Y(product[17]) );
  OAI21X1 U596 ( .A(n761), .B(n767), .C(n766), .Y(n760) );
  NAND2X1 U601 ( .A(n766), .B(n2925), .Y(n530) );
  NAND2X1 U604 ( .A(n1631), .B(n1616), .Y(n766) );
  XOR2X1 U605 ( .A(n775), .B(n531), .Y(product[16]) );
  OAI21X1 U607 ( .A(n786), .B(n769), .C(n770), .Y(n768) );
  NAND2X1 U608 ( .A(n2923), .B(n776), .Y(n769) );
  AOI21X1 U609 ( .A(n2923), .B(n777), .C(n772), .Y(n770) );
  NAND2X1 U612 ( .A(n774), .B(n2923), .Y(n531) );
  NAND2X1 U615 ( .A(n1645), .B(n1632), .Y(n774) );
  XOR2X1 U616 ( .A(n780), .B(n532), .Y(product[15]) );
  AOI21X1 U617 ( .A(n776), .B(n785), .C(n777), .Y(n775) );
  NOR2X1 U618 ( .A(n783), .B(n778), .Y(n776) );
  OAI21X1 U619 ( .A(n784), .B(n778), .C(n779), .Y(n777) );
  NAND2X1 U620 ( .A(n779), .B(n876), .Y(n532) );
  INVX2 U621 ( .A(n778), .Y(n876) );
  NOR2X1 U622 ( .A(n1659), .B(n1646), .Y(n778) );
  NAND2X1 U623 ( .A(n1659), .B(n1646), .Y(n779) );
  XNOR2X1 U624 ( .A(n785), .B(n533), .Y(product[14]) );
  AOI21X1 U625 ( .A(n781), .B(n785), .C(n782), .Y(n780) );
  NAND2X1 U628 ( .A(n784), .B(n781), .Y(n533) );
  NOR2X1 U630 ( .A(n1671), .B(n1660), .Y(n783) );
  NAND2X1 U631 ( .A(n1671), .B(n1660), .Y(n784) );
  XNOR2X1 U632 ( .A(n791), .B(n534), .Y(product[13]) );
  AOI21X1 U634 ( .A(n787), .B(n795), .C(n788), .Y(n786) );
  NOR2X1 U635 ( .A(n792), .B(n789), .Y(n787) );
  OAI21X1 U636 ( .A(n793), .B(n789), .C(n790), .Y(n788) );
  NAND2X1 U637 ( .A(n790), .B(n878), .Y(n534) );
  INVX2 U638 ( .A(n789), .Y(n878) );
  NOR2X1 U639 ( .A(n1683), .B(n1672), .Y(n789) );
  NAND2X1 U640 ( .A(n1683), .B(n1672), .Y(n790) );
  XOR2X1 U641 ( .A(n794), .B(n535), .Y(product[12]) );
  OAI21X1 U642 ( .A(n792), .B(n794), .C(n793), .Y(n791) );
  NAND2X1 U643 ( .A(n793), .B(n879), .Y(n535) );
  INVX2 U644 ( .A(n792), .Y(n879) );
  NOR2X1 U645 ( .A(n1693), .B(n1684), .Y(n792) );
  NAND2X1 U646 ( .A(n1693), .B(n1684), .Y(n793) );
  XOR2X1 U647 ( .A(n802), .B(n536), .Y(product[11]) );
  OAI21X1 U649 ( .A(n796), .B(n808), .C(n797), .Y(n795) );
  NAND2X1 U650 ( .A(n2922), .B(n2919), .Y(n796) );
  AOI21X1 U651 ( .A(n804), .B(n2919), .C(n799), .Y(n797) );
  NAND2X1 U654 ( .A(n801), .B(n2919), .Y(n536) );
  NAND2X1 U657 ( .A(n1703), .B(n1694), .Y(n801) );
  XNOR2X1 U658 ( .A(n807), .B(n537), .Y(product[10]) );
  AOI21X1 U659 ( .A(n2922), .B(n807), .C(n804), .Y(n802) );
  NAND2X1 U662 ( .A(n806), .B(n2922), .Y(n537) );
  NAND2X1 U665 ( .A(n1711), .B(n1704), .Y(n806) );
  XNOR2X1 U666 ( .A(n813), .B(n538), .Y(product[9]) );
  AOI21X1 U668 ( .A(n2921), .B(n813), .C(n810), .Y(n808) );
  NAND2X1 U671 ( .A(n812), .B(n2921), .Y(n538) );
  NAND2X1 U674 ( .A(n1719), .B(n1712), .Y(n812) );
  XOR2X1 U675 ( .A(n816), .B(n539), .Y(product[8]) );
  OAI21X1 U676 ( .A(n814), .B(n816), .C(n815), .Y(n813) );
  NAND2X1 U677 ( .A(n815), .B(n883), .Y(n539) );
  INVX2 U678 ( .A(n814), .Y(n883) );
  NOR2X1 U679 ( .A(n1725), .B(n1720), .Y(n814) );
  NAND2X1 U680 ( .A(n1725), .B(n1720), .Y(n815) );
  XNOR2X1 U681 ( .A(n821), .B(n540), .Y(product[7]) );
  AOI21X1 U682 ( .A(n825), .B(n817), .C(n818), .Y(n816) );
  NOR2X1 U683 ( .A(n822), .B(n819), .Y(n817) );
  OAI21X1 U684 ( .A(n823), .B(n819), .C(n820), .Y(n818) );
  NAND2X1 U685 ( .A(n820), .B(n884), .Y(n540) );
  NOR2X1 U687 ( .A(n1731), .B(n1726), .Y(n819) );
  NAND2X1 U688 ( .A(n1731), .B(n1726), .Y(n820) );
  XOR2X1 U689 ( .A(n541), .B(n824), .Y(product[6]) );
  OAI21X1 U690 ( .A(n822), .B(n824), .C(n823), .Y(n821) );
  NAND2X1 U691 ( .A(n823), .B(n885), .Y(n541) );
  INVX2 U692 ( .A(n822), .Y(n885) );
  NOR2X1 U693 ( .A(n1735), .B(n1732), .Y(n822) );
  NAND2X1 U694 ( .A(n1735), .B(n1732), .Y(n823) );
  XOR2X1 U695 ( .A(n542), .B(n828), .Y(product[5]) );
  OAI21X1 U697 ( .A(n826), .B(n828), .C(n827), .Y(n825) );
  NAND2X1 U698 ( .A(n827), .B(n886), .Y(n542) );
  INVX2 U699 ( .A(n826), .Y(n886) );
  NOR2X1 U700 ( .A(n1739), .B(n1736), .Y(n826) );
  NAND2X1 U701 ( .A(n1739), .B(n1736), .Y(n827) );
  XNOR2X1 U702 ( .A(n543), .B(n833), .Y(product[4]) );
  AOI21X1 U703 ( .A(n833), .B(n2920), .C(n830), .Y(n828) );
  NAND2X1 U706 ( .A(n832), .B(n2920), .Y(n543) );
  NAND2X1 U709 ( .A(n1741), .B(n1740), .Y(n832) );
  XOR2X1 U710 ( .A(n544), .B(n836), .Y(product[3]) );
  OAI21X1 U711 ( .A(n834), .B(n836), .C(n835), .Y(n833) );
  NAND2X1 U712 ( .A(n835), .B(n888), .Y(n544) );
  INVX2 U713 ( .A(n834), .Y(n888) );
  NOR2X1 U714 ( .A(n1757), .B(n1742), .Y(n834) );
  NAND2X1 U715 ( .A(n1757), .B(n1742), .Y(n835) );
  XNOR2X1 U716 ( .A(n545), .B(n841), .Y(product[2]) );
  AOI21X1 U717 ( .A(n841), .B(n2927), .C(n838), .Y(n836) );
  NAND2X1 U720 ( .A(n840), .B(n2927), .Y(n545) );
  NAND2X1 U723 ( .A(n2237), .B(n2944), .Y(n840) );
  NAND2X1 U729 ( .A(n1758), .B(n2238), .Y(n843) );
  FAX1 U730 ( .A(n905), .B(n922), .C(n903), .YC(n900), .YS(n901) );
  FAX1 U731 ( .A(n926), .B(n907), .C(n924), .YC(n902), .YS(n903) );
  FAX1 U732 ( .A(n911), .B(n928), .C(n909), .YC(n904), .YS(n905) );
  FAX1 U733 ( .A(n915), .B(n932), .C(n930), .YC(n906), .YS(n907) );
  FAX1 U734 ( .A(n934), .B(n917), .C(n913), .YC(n908), .YS(n909) );
  FAX1 U735 ( .A(n1829), .B(n938), .C(n936), .YC(n910), .YS(n911) );
  FAX1 U736 ( .A(n1853), .B(n1787), .C(n1807), .YC(n912), .YS(n913) );
  FAX1 U737 ( .A(n1907), .B(n1769), .C(n1879), .YC(n914), .YS(n915) );
  FAX1 U738 ( .A(n919), .B(n1969), .C(n1937), .YC(n916), .YS(n917) );
  INVX2 U739 ( .A(n918), .Y(n919) );
  FAX1 U740 ( .A(n925), .B(n942), .C(n923), .YC(n920), .YS(n921) );
  FAX1 U741 ( .A(n946), .B(n927), .C(n944), .YC(n922), .YS(n923) );
  FAX1 U742 ( .A(n948), .B(n931), .C(n929), .YC(n924), .YS(n925) );
  FAX1 U743 ( .A(n933), .B(n952), .C(n950), .YC(n926), .YS(n927) );
  FAX1 U744 ( .A(n954), .B(n935), .C(n937), .YC(n928), .YS(n929) );
  FAX1 U745 ( .A(n958), .B(n956), .C(n939), .YC(n930), .YS(n931) );
  FAX1 U746 ( .A(n1970), .B(n1938), .C(n2002), .YC(n932), .YS(n933) );
  FAX1 U747 ( .A(n1788), .B(n1908), .C(n1830), .YC(n934), .YS(n935) );
  FAX1 U748 ( .A(n1854), .B(n1770), .C(n1808), .YC(n936), .YS(n937) );
  FAX1 U749 ( .A(n960), .B(n1760), .C(n1880), .YC(n938), .YS(n939) );
  FAX1 U750 ( .A(n945), .B(n964), .C(n943), .YC(n940), .YS(n941) );
  FAX1 U751 ( .A(n968), .B(n947), .C(n966), .YC(n942), .YS(n943) );
  FAX1 U752 ( .A(n970), .B(n951), .C(n949), .YC(n944), .YS(n945) );
  FAX1 U753 ( .A(n953), .B(n974), .C(n972), .YC(n946), .YS(n947) );
  FAX1 U754 ( .A(n959), .B(n955), .C(n957), .YC(n948), .YS(n949) );
  FAX1 U755 ( .A(n980), .B(n976), .C(n978), .YC(n950), .YS(n951) );
  FAX1 U756 ( .A(n1909), .B(n1881), .C(n982), .YC(n952), .YS(n953) );
  FAX1 U757 ( .A(n1855), .B(n1809), .C(n1831), .YC(n954), .YS(n955) );
  FAX1 U758 ( .A(n1939), .B(n1771), .C(n1789), .YC(n956), .YS(n957) );
  FAX1 U759 ( .A(n961), .B(n2003), .C(n1971), .YC(n958), .YS(n959) );
  INVX2 U760 ( .A(n960), .Y(n961) );
  FAX1 U761 ( .A(n988), .B(n986), .C(n965), .YC(n962), .YS(n963) );
  FAX1 U762 ( .A(n990), .B(n969), .C(n967), .YC(n964), .YS(n965) );
  FAX1 U763 ( .A(n973), .B(n971), .C(n992), .YC(n966), .YS(n967) );
  FAX1 U764 ( .A(n996), .B(n994), .C(n975), .YC(n968), .YS(n969) );
  FAX1 U765 ( .A(n977), .B(n981), .C(n979), .YC(n970), .YS(n971) );
  FAX1 U766 ( .A(n1000), .B(n998), .C(n983), .YC(n972), .YS(n973) );
  FAX1 U767 ( .A(n2036), .B(n1004), .C(n1002), .YC(n974), .YS(n975) );
  FAX1 U768 ( .A(n2004), .B(n1832), .C(n1972), .YC(n976), .YS(n977) );
  FAX1 U769 ( .A(n1910), .B(n1810), .C(n1940), .YC(n978), .YS(n979) );
  FAX1 U770 ( .A(n1856), .B(n1772), .C(n1790), .YC(n980), .YS(n981) );
  FAX1 U771 ( .A(n1006), .B(n1761), .C(n1882), .YC(n982), .YS(n983) );
  FAX1 U772 ( .A(n989), .B(n1010), .C(n987), .YC(n984), .YS(n985) );
  FAX1 U773 ( .A(n1014), .B(n991), .C(n1012), .YC(n986), .YS(n987) );
  FAX1 U774 ( .A(n995), .B(n1016), .C(n993), .YC(n988), .YS(n989) );
  FAX1 U775 ( .A(n1020), .B(n1018), .C(n997), .YC(n990), .YS(n991) );
  FAX1 U776 ( .A(n1003), .B(n1001), .C(n1022), .YC(n992), .YS(n993) );
  FAX1 U777 ( .A(n1024), .B(n1005), .C(n999), .YC(n994), .YS(n995) );
  FAX1 U778 ( .A(n1030), .B(n1028), .C(n1026), .YC(n996), .YS(n997) );
  FAX1 U779 ( .A(n1911), .B(n1857), .C(n1883), .YC(n998), .YS(n999) );
  FAX1 U780 ( .A(n1811), .B(n1941), .C(n1833), .YC(n1000), .YS(n1001) );
  FAX1 U781 ( .A(n1973), .B(n1773), .C(n1791), .YC(n1002), .YS(n1003) );
  FAX1 U782 ( .A(n1007), .B(n2037), .C(n2005), .YC(n1004), .YS(n1005) );
  INVX2 U783 ( .A(n1006), .Y(n1007) );
  FAX1 U784 ( .A(n1013), .B(n1034), .C(n1011), .YC(n1008), .YS(n1009) );
  FAX1 U785 ( .A(n1038), .B(n1015), .C(n1036), .YC(n1010), .YS(n1011) );
  FAX1 U786 ( .A(n1019), .B(n1040), .C(n1017), .YC(n1012), .YS(n1013) );
  FAX1 U787 ( .A(n1023), .B(n1042), .C(n1021), .YC(n1014), .YS(n1015) );
  FAX1 U788 ( .A(n1029), .B(n1046), .C(n1044), .YC(n1016), .YS(n1017) );
  FAX1 U789 ( .A(n1050), .B(n1025), .C(n1027), .YC(n1018), .YS(n1019) );
  FAX1 U790 ( .A(n1052), .B(n1048), .C(n1031), .YC(n1020), .YS(n1021) );
  FAX1 U791 ( .A(n2038), .B(n2070), .C(n1054), .YC(n1022), .YS(n1023) );
  FAX1 U792 ( .A(n2006), .B(n1834), .C(n1974), .YC(n1024), .YS(n1025) );
  FAX1 U793 ( .A(n1942), .B(n1774), .C(n1858), .YC(n1026), .YS(n1027) );
  FAX1 U794 ( .A(n1884), .B(n1792), .C(n1812), .YC(n1028), .YS(n1029) );
  FAX1 U795 ( .A(n1056), .B(n1762), .C(n1912), .YC(n1030), .YS(n1031) );
  FAX1 U796 ( .A(n1037), .B(n1060), .C(n1035), .YC(n1032), .YS(n1033) );
  FAX1 U797 ( .A(n1064), .B(n1039), .C(n1062), .YC(n1034), .YS(n1035) );
  FAX1 U798 ( .A(n1043), .B(n1066), .C(n1041), .YC(n1036), .YS(n1037) );
  FAX1 U799 ( .A(n1047), .B(n1045), .C(n1068), .YC(n1038), .YS(n1039) );
  FAX1 U800 ( .A(n1053), .B(n1072), .C(n1070), .YC(n1040), .YS(n1041) );
  FAX1 U801 ( .A(n1051), .B(n1049), .C(n1074), .YC(n1042), .YS(n1043) );
  FAX1 U802 ( .A(n1078), .B(n1076), .C(n1055), .YC(n1044), .YS(n1045) );
  FAX1 U803 ( .A(n1943), .B(n1082), .C(n1080), .YC(n1046), .YS(n1047) );
  FAX1 U804 ( .A(n1975), .B(n1859), .C(n1913), .YC(n1048), .YS(n1049) );
  FAX1 U805 ( .A(n1835), .B(n2007), .C(n1813), .YC(n1050), .YS(n1051) );
  FAX1 U806 ( .A(n2039), .B(n1775), .C(n1793), .YC(n1052), .YS(n1053) );
  FAX1 U807 ( .A(n1057), .B(n2071), .C(n1885), .YC(n1054), .YS(n1055) );
  INVX2 U808 ( .A(n1056), .Y(n1057) );
  FAX1 U809 ( .A(n1063), .B(n1086), .C(n1061), .YC(n1058), .YS(n1059) );
  FAX1 U810 ( .A(n1090), .B(n1065), .C(n1088), .YC(n1060), .YS(n1061) );
  FAX1 U811 ( .A(n1094), .B(n1092), .C(n1067), .YC(n1062), .YS(n1063) );
  FAX1 U812 ( .A(n1073), .B(n1071), .C(n1069), .YC(n1064), .YS(n1065) );
  FAX1 U813 ( .A(n1100), .B(n1098), .C(n1096), .YC(n1066), .YS(n1067) );
  FAX1 U814 ( .A(n1079), .B(n1081), .C(n1075), .YC(n1068), .YS(n1069) );
  FAX1 U815 ( .A(n1104), .B(n1102), .C(n1077), .YC(n1070), .YS(n1071) );
  FAX1 U816 ( .A(n1108), .B(n1106), .C(n1083), .YC(n1072), .YS(n1073) );
  FAX1 U817 ( .A(n2072), .B(n2040), .C(n2104), .YC(n1074), .YS(n1075) );
  FAX1 U818 ( .A(n1860), .B(n2008), .C(n1976), .YC(n1076), .YS(n1077) );
  FAX1 U819 ( .A(n1914), .B(n1776), .C(n1836), .YC(n1078), .YS(n1079) );
  FAX1 U820 ( .A(n1886), .B(n1794), .C(n1814), .YC(n1080), .YS(n1081) );
  FAX1 U821 ( .A(n1110), .B(n1763), .C(n1944), .YC(n1082), .YS(n1083) );
  FAX1 U822 ( .A(n1089), .B(n1114), .C(n1087), .YC(n1084), .YS(n1085) );
  FAX1 U823 ( .A(n1118), .B(n1091), .C(n1116), .YC(n1086), .YS(n1087) );
  FAX1 U824 ( .A(n1095), .B(n1120), .C(n1093), .YC(n1088), .YS(n1089) );
  FAX1 U825 ( .A(n1099), .B(n1097), .C(n1122), .YC(n1090), .YS(n1091) );
  FAX1 U826 ( .A(n1128), .B(n1126), .C(n1124), .YC(n1092), .YS(n1093) );
  FAX1 U827 ( .A(n1105), .B(n1107), .C(n1101), .YC(n1094), .YS(n1095) );
  FAX1 U828 ( .A(n1132), .B(n1109), .C(n1103), .YC(n1096), .YS(n1097) );
  FAX1 U829 ( .A(n1136), .B(n1130), .C(n1134), .YC(n1098), .YS(n1099) );
  FAX1 U830 ( .A(n1915), .B(n1861), .C(n1138), .YC(n1100), .YS(n1101) );
  FAX1 U831 ( .A(n1945), .B(n1815), .C(n1837), .YC(n1102), .YS(n1103) );
  FAX1 U832 ( .A(n2009), .B(n1795), .C(n1977), .YC(n1104), .YS(n1105) );
  FAX1 U833 ( .A(n1887), .B(n2041), .C(n1777), .YC(n1106), .YS(n1107) );
  FAX1 U834 ( .A(n1111), .B(n2105), .C(n2073), .YC(n1108), .YS(n1109) );
  INVX2 U835 ( .A(n1110), .Y(n1111) );
  FAX1 U836 ( .A(n1117), .B(n1142), .C(n1115), .YC(n1112), .YS(n1113) );
  FAX1 U837 ( .A(n1146), .B(n1119), .C(n1144), .YC(n1114), .YS(n1115) );
  FAX1 U838 ( .A(n1123), .B(n1148), .C(n1121), .YC(n1116), .YS(n1117) );
  FAX1 U839 ( .A(n1127), .B(n1125), .C(n1150), .YC(n1118), .YS(n1119) );
  FAX1 U840 ( .A(n1154), .B(n1129), .C(n1152), .YC(n1120), .YS(n1121) );
  FAX1 U841 ( .A(n1137), .B(n1135), .C(n1156), .YC(n1122), .YS(n1123) );
  FAX1 U842 ( .A(n1162), .B(n1131), .C(n1133), .YC(n1124), .YS(n1125) );
  FAX1 U843 ( .A(n1160), .B(n1164), .C(n1139), .YC(n1126), .YS(n1127) );
  FAX1 U844 ( .A(n2138), .B(n1166), .C(n1158), .YC(n1128), .YS(n1129) );
  FAX1 U845 ( .A(n2074), .B(n2106), .C(n1888), .YC(n1130), .YS(n1131) );
  FAX1 U846 ( .A(n1862), .B(n2010), .C(n2042), .YC(n1132), .YS(n1133) );
  FAX1 U847 ( .A(n1978), .B(n1796), .C(n1838), .YC(n1134), .YS(n1135) );
  FAX1 U848 ( .A(n1916), .B(n1778), .C(n1816), .YC(n1136), .YS(n1137) );
  FAX1 U849 ( .A(n1168), .B(n1764), .C(n1946), .YC(n1138), .YS(n1139) );
  FAX1 U850 ( .A(n1145), .B(n1172), .C(n1143), .YC(n1140), .YS(n1141) );
  FAX1 U851 ( .A(n1176), .B(n1147), .C(n1174), .YC(n1142), .YS(n1143) );
  FAX1 U852 ( .A(n1151), .B(n1178), .C(n1149), .YC(n1144), .YS(n1145) );
  FAX1 U853 ( .A(n1155), .B(n1153), .C(n1180), .YC(n1146), .YS(n1147) );
  FAX1 U854 ( .A(n1184), .B(n1157), .C(n1182), .YC(n1148), .YS(n1149) );
  FAX1 U855 ( .A(n1163), .B(n1188), .C(n1186), .YC(n1150), .YS(n1151) );
  FAX1 U856 ( .A(n1159), .B(n1165), .C(n1161), .YC(n1152), .YS(n1153) );
  FAX1 U857 ( .A(n1194), .B(n1196), .C(n1167), .YC(n1154), .YS(n1155) );
  FAX1 U858 ( .A(n1198), .B(n1190), .C(n1192), .YC(n1156), .YS(n1157) );
  FAX1 U859 ( .A(n1947), .B(n1863), .C(n1917), .YC(n1158), .YS(n1159) );
  FAX1 U860 ( .A(n1979), .B(n1817), .C(n1839), .YC(n1160), .YS(n1161) );
  FAX1 U861 ( .A(n2043), .B(n1797), .C(n2011), .YC(n1162), .YS(n1163) );
  FAX1 U862 ( .A(n1889), .B(n2075), .C(n1779), .YC(n1164), .YS(n1165) );
  FAX1 U863 ( .A(n1169), .B(n2139), .C(n2107), .YC(n1166), .YS(n1167) );
  INVX2 U864 ( .A(n1168), .Y(n1169) );
  FAX1 U865 ( .A(n1175), .B(n1202), .C(n1173), .YC(n1170), .YS(n1171) );
  FAX1 U866 ( .A(n1206), .B(n1177), .C(n1204), .YC(n1172), .YS(n1173) );
  FAX1 U867 ( .A(n1181), .B(n1208), .C(n1179), .YC(n1174), .YS(n1175) );
  FAX1 U868 ( .A(n1185), .B(n1183), .C(n1210), .YC(n1176), .YS(n1177) );
  FAX1 U869 ( .A(n1214), .B(n1212), .C(n1187), .YC(n1178), .YS(n1179) );
  FAX1 U870 ( .A(n1218), .B(n1189), .C(n1216), .YC(n1180), .YS(n1181) );
  FAX1 U871 ( .A(n1195), .B(n1197), .C(n1193), .YC(n1182), .YS(n1183) );
  FAX1 U872 ( .A(n1224), .B(n1222), .C(n1191), .YC(n1184), .YS(n1185) );
  FAX1 U873 ( .A(n1220), .B(n1226), .C(n1199), .YC(n1186), .YS(n1187) );
  FAX1 U874 ( .A(n2076), .B(n2172), .C(n1228), .YC(n1188), .YS(n1189) );
  FAX1 U875 ( .A(n2108), .B(n2044), .C(n2140), .YC(n1190), .YS(n1191) );
  FAX1 U876 ( .A(n1864), .B(n1948), .C(n1890), .YC(n1192), .YS(n1193) );
  FAX1 U877 ( .A(n2012), .B(n1840), .C(n1818), .YC(n1194), .YS(n1195) );
  FAX1 U878 ( .A(n1918), .B(n1798), .C(n1780), .YC(n1196), .YS(n1197) );
  FAX1 U879 ( .A(n1230), .B(n1765), .C(n1980), .YC(n1198), .YS(n1199) );
  FAX1 U880 ( .A(n1205), .B(n1234), .C(n1203), .YC(n1200), .YS(n1201) );
  FAX1 U881 ( .A(n1238), .B(n1207), .C(n1236), .YC(n1202), .YS(n1203) );
  FAX1 U882 ( .A(n1240), .B(n1211), .C(n1209), .YC(n1204), .YS(n1205) );
  FAX1 U883 ( .A(n1217), .B(n1213), .C(n1242), .YC(n1206), .YS(n1207) );
  FAX1 U884 ( .A(n1246), .B(n1244), .C(n1215), .YC(n1208), .YS(n1209) );
  FAX1 U885 ( .A(n1250), .B(n1248), .C(n1219), .YC(n1210), .YS(n1211) );
  FAX1 U886 ( .A(n1225), .B(n1227), .C(n1223), .YC(n1212), .YS(n1213) );
  FAX1 U887 ( .A(n1256), .B(n1254), .C(n1221), .YC(n1214), .YS(n1215) );
  FAX1 U888 ( .A(n1252), .B(n1258), .C(n1229), .YC(n1216), .YS(n1217) );
  FAX1 U889 ( .A(n1981), .B(n2013), .C(n1260), .YC(n1218), .YS(n1219) );
  FAX1 U890 ( .A(n2045), .B(n1919), .C(n1949), .YC(n1220), .YS(n1221) );
  FAX1 U891 ( .A(n1865), .B(n2077), .C(n1891), .YC(n1222), .YS(n1223) );
  FAX1 U892 ( .A(n2109), .B(n1819), .C(n1841), .YC(n1224), .YS(n1225) );
  FAX1 U893 ( .A(n2141), .B(n1781), .C(n1799), .YC(n1226), .YS(n1227) );
  FAX1 U894 ( .A(n1766), .B(n1262), .C(n2173), .YC(n1228), .YS(n1229) );
  FAX1 U896 ( .A(n1237), .B(n1265), .C(n1235), .YC(n1232), .YS(n1233) );
  FAX1 U897 ( .A(n1269), .B(n1239), .C(n1267), .YC(n1234), .YS(n1235) );
  FAX1 U898 ( .A(n1271), .B(n1243), .C(n1241), .YC(n1236), .YS(n1237) );
  FAX1 U899 ( .A(n1247), .B(n1245), .C(n1273), .YC(n1238), .YS(n1239) );
  FAX1 U900 ( .A(n1251), .B(n1275), .C(n1249), .YC(n1240), .YS(n1241) );
  FAX1 U901 ( .A(n1255), .B(n1279), .C(n1277), .YC(n1242), .YS(n1243) );
  FAX1 U902 ( .A(n1257), .B(n1259), .C(n1281), .YC(n1244), .YS(n1245) );
  FAX1 U903 ( .A(n1285), .B(n1261), .C(n1253), .YC(n1246), .YS(n1247) );
  FAX1 U904 ( .A(n1283), .B(n1289), .C(n1287), .YC(n1248), .YS(n1249) );
  FAX1 U905 ( .A(n2110), .B(n2206), .C(n1291), .YC(n1250), .YS(n1251) );
  FAX1 U906 ( .A(n2142), .B(n2078), .C(n2174), .YC(n1252), .YS(n1253) );
  FAX1 U907 ( .A(n1892), .B(n1982), .C(n1920), .YC(n1254), .YS(n1255) );
  FAX1 U908 ( .A(n2046), .B(n1866), .C(n1842), .YC(n1256), .YS(n1257) );
  FAX1 U909 ( .A(n1950), .B(n1820), .C(n1782), .YC(n1258), .YS(n1259) );
  FAX1 U910 ( .A(n1262), .B(n1800), .C(n2014), .YC(n1260), .YS(n1261) );
  INVX2 U911 ( .A(n1230), .Y(n1262) );
  FAX1 U912 ( .A(n1268), .B(n1295), .C(n1266), .YC(n1263), .YS(n1264) );
  FAX1 U913 ( .A(n1272), .B(n1270), .C(n1297), .YC(n1265), .YS(n1266) );
  FAX1 U914 ( .A(n1274), .B(n1301), .C(n1299), .YC(n1267), .YS(n1268) );
  FAX1 U915 ( .A(n1278), .B(n1276), .C(n1303), .YC(n1269), .YS(n1270) );
  FAX1 U916 ( .A(n1307), .B(n1305), .C(n1280), .YC(n1271), .YS(n1272) );
  FAX1 U917 ( .A(n1288), .B(n1282), .C(n1309), .YC(n1273), .YS(n1274) );
  FAX1 U918 ( .A(n1284), .B(n1290), .C(n1286), .YC(n1275), .YS(n1276) );
  FAX1 U919 ( .A(n1311), .B(n1315), .C(n1292), .YC(n1277), .YS(n1278) );
  FAX1 U920 ( .A(n1313), .B(n1319), .C(n1317), .YC(n1279), .YS(n1280) );
  FAX1 U921 ( .A(n2015), .B(n2047), .C(n1321), .YC(n1281), .YS(n1282) );
  FAX1 U922 ( .A(n2079), .B(n1921), .C(n1951), .YC(n1283), .YS(n1284) );
  FAX1 U923 ( .A(n2111), .B(n1867), .C(n1893), .YC(n1285), .YS(n1286) );
  FAX1 U924 ( .A(n1983), .B(n2143), .C(n1843), .YC(n1287), .YS(n1288) );
  FAX1 U925 ( .A(n2175), .B(n1801), .C(n1821), .YC(n1289), .YS(n1290) );
  FAX1 U926 ( .A(n1767), .B(n2207), .C(n1783), .YC(n1291), .YS(n1292) );
  FAX1 U927 ( .A(n1298), .B(n1325), .C(n1296), .YC(n1293), .YS(n1294) );
  FAX1 U928 ( .A(n1302), .B(n1300), .C(n1327), .YC(n1295), .YS(n1296) );
  FAX1 U929 ( .A(n1304), .B(n1331), .C(n1329), .YC(n1297), .YS(n1298) );
  FAX1 U930 ( .A(n1308), .B(n1333), .C(n1306), .YC(n1299), .YS(n1300) );
  FAX1 U931 ( .A(n1337), .B(n1310), .C(n1335), .YC(n1301), .YS(n1302) );
  FAX1 U932 ( .A(n1314), .B(n1316), .C(n1339), .YC(n1303), .YS(n1304) );
  FAX1 U933 ( .A(n1312), .B(n1320), .C(n1318), .YC(n1305), .YS(n1306) );
  FAX1 U934 ( .A(n1341), .B(n1345), .C(n1343), .YC(n1307), .YS(n1308) );
  FAX1 U935 ( .A(n1322), .B(n1349), .C(n1347), .YC(n1309), .YS(n1310) );
  FAX1 U936 ( .A(n1868), .B(n2016), .C(n1922), .YC(n1311), .YS(n1312) );
  FAX1 U937 ( .A(n2048), .B(n1822), .C(n1844), .YC(n1313), .YS(n1314) );
  FAX1 U938 ( .A(n1894), .B(n2112), .C(n2080), .YC(n1315), .YS(n1316) );
  FAX1 U939 ( .A(n1984), .B(n2176), .C(n2144), .YC(n1317), .YS(n1318) );
  FAX1 U940 ( .A(n1952), .B(n1784), .C(n1802), .YC(n1319), .YS(n1320) );
  HAX1 U941 ( .A(n2208), .B(n1743), .YC(n1321), .YS(n1322) );
  FAX1 U942 ( .A(n1328), .B(n1353), .C(n1326), .YC(n1323), .YS(n1324) );
  FAX1 U943 ( .A(n1332), .B(n1330), .C(n1355), .YC(n1325), .YS(n1326) );
  FAX1 U944 ( .A(n1334), .B(n1359), .C(n1357), .YC(n1327), .YS(n1328) );
  FAX1 U945 ( .A(n1361), .B(n1338), .C(n1336), .YC(n1329), .YS(n1330) );
  FAX1 U946 ( .A(n1365), .B(n1340), .C(n1363), .YC(n1331), .YS(n1332) );
  FAX1 U947 ( .A(n1344), .B(n1346), .C(n1367), .YC(n1333), .YS(n1334) );
  FAX1 U948 ( .A(n1350), .B(n1342), .C(n1348), .YC(n1335), .YS(n1336) );
  FAX1 U949 ( .A(n1371), .B(n1375), .C(n1373), .YC(n1337), .YS(n1338) );
  FAX1 U950 ( .A(n2937), .B(n1377), .C(n1369), .YC(n1339), .YS(n1340) );
  FAX1 U951 ( .A(n2017), .B(n1953), .C(n1985), .YC(n1341), .YS(n1342) );
  FAX1 U952 ( .A(n2049), .B(n1895), .C(n1923), .YC(n1343), .YS(n1344) );
  FAX1 U953 ( .A(n2081), .B(n1845), .C(n1869), .YC(n1345), .YS(n1346) );
  FAX1 U954 ( .A(n2145), .B(n1823), .C(n2113), .YC(n1347), .YS(n1348) );
  FAX1 U955 ( .A(n2209), .B(n2177), .C(n1803), .YC(n1349), .YS(n1350) );
  FAX1 U956 ( .A(n1356), .B(n1381), .C(n1354), .YC(n1351), .YS(n1352) );
  FAX1 U957 ( .A(n1385), .B(n1358), .C(n1383), .YC(n1353), .YS(n1354) );
  FAX1 U958 ( .A(n1362), .B(n1387), .C(n1360), .YC(n1355), .YS(n1356) );
  FAX1 U959 ( .A(n1366), .B(n1389), .C(n1364), .YC(n1357), .YS(n1358) );
  FAX1 U960 ( .A(n1368), .B(n1393), .C(n1391), .YC(n1359), .YS(n1360) );
  FAX1 U961 ( .A(n1374), .B(n1376), .C(n1395), .YC(n1361), .YS(n1362) );
  FAX1 U962 ( .A(n1401), .B(n1370), .C(n1372), .YC(n1363), .YS(n1364) );
  FAX1 U963 ( .A(n1403), .B(n1397), .C(n1399), .YC(n1365), .YS(n1366) );
  FAX1 U964 ( .A(n2018), .B(n2050), .C(n1378), .YC(n1367), .YS(n1368) );
  FAX1 U965 ( .A(n2082), .B(n1924), .C(n1954), .YC(n1369), .YS(n1370) );
  FAX1 U966 ( .A(n1846), .B(n1824), .C(n1870), .YC(n1371), .YS(n1372) );
  FAX1 U967 ( .A(n1896), .B(n2114), .C(n1804), .YC(n1373), .YS(n1374) );
  FAX1 U968 ( .A(n1986), .B(n2178), .C(n2146), .YC(n1375), .YS(n1376) );
  HAX1 U969 ( .A(n2210), .B(n1744), .YC(n1377), .YS(n1378) );
  FAX1 U970 ( .A(n1384), .B(n1407), .C(n1382), .YC(n1379), .YS(n1380) );
  FAX1 U971 ( .A(n1411), .B(n1386), .C(n1409), .YC(n1381), .YS(n1382) );
  FAX1 U972 ( .A(n1390), .B(n1413), .C(n1388), .YC(n1383), .YS(n1384) );
  FAX1 U973 ( .A(n1394), .B(n1415), .C(n1392), .YC(n1385), .YS(n1386) );
  FAX1 U974 ( .A(n1396), .B(n1419), .C(n1417), .YC(n1387), .YS(n1388) );
  FAX1 U975 ( .A(n1400), .B(n1398), .C(n1402), .YC(n1389), .YS(n1390) );
  FAX1 U976 ( .A(n1421), .B(n1423), .C(n1404), .YC(n1391), .YS(n1392) );
  FAX1 U977 ( .A(n1429), .B(n1427), .C(n1425), .YC(n1393), .YS(n1394) );
  FAX1 U978 ( .A(n2019), .B(n1987), .C(n2931), .YC(n1395), .YS(n1396) );
  FAX1 U979 ( .A(n2051), .B(n1925), .C(n1955), .YC(n1397), .YS(n1398) );
  FAX1 U980 ( .A(n2083), .B(n1871), .C(n1897), .YC(n1399), .YS(n1400) );
  FAX1 U981 ( .A(n2147), .B(n1847), .C(n2115), .YC(n1401), .YS(n1402) );
  FAX1 U982 ( .A(n2211), .B(n2179), .C(n1825), .YC(n1403), .YS(n1404) );
  FAX1 U983 ( .A(n1410), .B(n1433), .C(n1408), .YC(n1405), .YS(n1406) );
  FAX1 U984 ( .A(n1414), .B(n1412), .C(n1435), .YC(n1407), .YS(n1408) );
  FAX1 U985 ( .A(n1416), .B(n1439), .C(n1437), .YC(n1409), .YS(n1410) );
  FAX1 U986 ( .A(n1420), .B(n1441), .C(n1418), .YC(n1411), .YS(n1412) );
  FAX1 U987 ( .A(n1424), .B(n1445), .C(n1443), .YC(n1413), .YS(n1414) );
  FAX1 U988 ( .A(n1422), .B(n1428), .C(n1426), .YC(n1415), .YS(n1416) );
  FAX1 U989 ( .A(n1447), .B(n1449), .C(n1451), .YC(n1417), .YS(n1418) );
  FAX1 U990 ( .A(n2084), .B(n1430), .C(n1453), .YC(n1419), .YS(n1420) );
  FAX1 U991 ( .A(n2116), .B(n1956), .C(n2052), .YC(n1421), .YS(n1422) );
  FAX1 U992 ( .A(n2148), .B(n1898), .C(n1926), .YC(n1423), .YS(n1424) );
  FAX1 U993 ( .A(n2020), .B(n1872), .C(n2180), .YC(n1425), .YS(n1426) );
  FAX1 U994 ( .A(n1988), .B(n1826), .C(n1848), .YC(n1427), .YS(n1428) );
  HAX1 U995 ( .A(n2212), .B(n1745), .YC(n1429), .YS(n1430) );
  FAX1 U996 ( .A(n1436), .B(n1457), .C(n1434), .YC(n1431), .YS(n1432) );
  FAX1 U997 ( .A(n1461), .B(n1459), .C(n1438), .YC(n1433), .YS(n1434) );
  FAX1 U998 ( .A(n1444), .B(n1442), .C(n1440), .YC(n1435), .YS(n1436) );
  FAX1 U999 ( .A(n1467), .B(n1465), .C(n1463), .YC(n1437), .YS(n1438) );
  FAX1 U1000 ( .A(n1452), .B(n1450), .C(n1446), .YC(n1439), .YS(n1440) );
  FAX1 U1001 ( .A(n1473), .B(n1454), .C(n1448), .YC(n1441), .YS(n1442) );
  FAX1 U1002 ( .A(n1475), .B(n1469), .C(n1471), .YC(n1443), .YS(n1444) );
  FAX1 U1003 ( .A(n2053), .B(n2940), .C(n1477), .YC(n1445), .YS(n1446) );
  FAX1 U1004 ( .A(n2085), .B(n1989), .C(n2021), .YC(n1447), .YS(n1448) );
  FAX1 U1005 ( .A(n2117), .B(n1927), .C(n1957), .YC(n1449), .YS(n1450) );
  FAX1 U1006 ( .A(n2149), .B(n1873), .C(n1899), .YC(n1451), .YS(n1452) );
  FAX1 U1007 ( .A(n1849), .B(n2181), .C(n2213), .YC(n1453), .YS(n1454) );
  FAX1 U1008 ( .A(n1460), .B(n1481), .C(n1458), .YC(n1455), .YS(n1456) );
  FAX1 U1009 ( .A(n1485), .B(n1483), .C(n1462), .YC(n1457), .YS(n1458) );
  FAX1 U1010 ( .A(n1487), .B(n1466), .C(n1464), .YC(n1459), .YS(n1460) );
  FAX1 U1011 ( .A(n1491), .B(n1489), .C(n1468), .YC(n1461), .YS(n1462) );
  FAX1 U1012 ( .A(n1472), .B(n1476), .C(n1474), .YC(n1463), .YS(n1464) );
  FAX1 U1013 ( .A(n1495), .B(n1493), .C(n1470), .YC(n1465), .YS(n1466) );
  FAX1 U1014 ( .A(n1478), .B(n1499), .C(n1497), .YC(n1467), .YS(n1468) );
  FAX1 U1015 ( .A(n2086), .B(n1990), .C(n2054), .YC(n1469), .YS(n1470) );
  FAX1 U1016 ( .A(n2118), .B(n1900), .C(n1958), .YC(n1471), .YS(n1472) );
  FAX1 U1017 ( .A(n1928), .B(n1850), .C(n1874), .YC(n1473), .YS(n1474) );
  FAX1 U1018 ( .A(n2022), .B(n2182), .C(n2150), .YC(n1475), .YS(n1476) );
  HAX1 U1019 ( .A(n2214), .B(n1746), .YC(n1477), .YS(n1478) );
  FAX1 U1020 ( .A(n1484), .B(n1503), .C(n1482), .YC(n1479), .YS(n1480) );
  FAX1 U1021 ( .A(n1507), .B(n1486), .C(n1505), .YC(n1481), .YS(n1482) );
  FAX1 U1022 ( .A(n1509), .B(n1490), .C(n1488), .YC(n1483), .YS(n1484) );
  FAX1 U1023 ( .A(n1513), .B(n1511), .C(n1492), .YC(n1485), .YS(n1486) );
  FAX1 U1024 ( .A(n1494), .B(n1498), .C(n1496), .YC(n1487), .YS(n1488) );
  FAX1 U1025 ( .A(n1517), .B(n1515), .C(n1500), .YC(n1489), .YS(n1490) );
  FAX1 U1026 ( .A(n2942), .B(n1521), .C(n1519), .YC(n1491), .YS(n1492) );
  FAX1 U1027 ( .A(n2087), .B(n2023), .C(n2055), .YC(n1493), .YS(n1494) );
  FAX1 U1028 ( .A(n2119), .B(n1959), .C(n1991), .YC(n1495), .YS(n1496) );
  FAX1 U1029 ( .A(n2151), .B(n1901), .C(n1929), .YC(n1497), .YS(n1498) );
  FAX1 U1030 ( .A(n2215), .B(n2183), .C(n1875), .YC(n1499), .YS(n1500) );
  FAX1 U1031 ( .A(n1506), .B(n1525), .C(n1504), .YC(n1501), .YS(n1502) );
  FAX1 U1032 ( .A(n1529), .B(n1508), .C(n1527), .YC(n1503), .YS(n1504) );
  FAX1 U1033 ( .A(n1531), .B(n1512), .C(n1510), .YC(n1505), .YS(n1506) );
  FAX1 U1034 ( .A(n1518), .B(n1514), .C(n1533), .YC(n1507), .YS(n1508) );
  FAX1 U1035 ( .A(n1516), .B(n1520), .C(n1535), .YC(n1509), .YS(n1510) );
  FAX1 U1036 ( .A(n1541), .B(n1539), .C(n1537), .YC(n1511), .YS(n1512) );
  FAX1 U1037 ( .A(n2088), .B(n1992), .C(n1522), .YC(n1513), .YS(n1514) );
  FAX1 U1038 ( .A(n2120), .B(n1930), .C(n1960), .YC(n1515), .YS(n1516) );
  FAX1 U1039 ( .A(n2056), .B(n2184), .C(n2152), .YC(n1517), .YS(n1518) );
  FAX1 U1040 ( .A(n2024), .B(n1876), .C(n1902), .YC(n1519), .YS(n1520) );
  HAX1 U1041 ( .A(n2216), .B(n1747), .YC(n1521), .YS(n1522) );
  FAX1 U1042 ( .A(n1528), .B(n1545), .C(n1526), .YC(n1523), .YS(n1524) );
  FAX1 U1043 ( .A(n1532), .B(n1530), .C(n1547), .YC(n1525), .YS(n1526) );
  FAX1 U1044 ( .A(n1551), .B(n1534), .C(n1549), .YC(n1527), .YS(n1528) );
  FAX1 U1045 ( .A(n1540), .B(n1536), .C(n1553), .YC(n1529), .YS(n1530) );
  FAX1 U1046 ( .A(n1555), .B(n1542), .C(n1538), .YC(n1531), .YS(n1532) );
  FAX1 U1047 ( .A(n1561), .B(n1559), .C(n1557), .YC(n1533), .YS(n1534) );
  FAX1 U1048 ( .A(n2089), .B(n2057), .C(n2930), .YC(n1535), .YS(n1536) );
  FAX1 U1049 ( .A(n2121), .B(n1993), .C(n2025), .YC(n1537), .YS(n1538) );
  FAX1 U1050 ( .A(n2153), .B(n1931), .C(n1961), .YC(n1539), .YS(n1540) );
  FAX1 U1051 ( .A(n2217), .B(n2185), .C(n1903), .YC(n1541), .YS(n1542) );
  FAX1 U1052 ( .A(n1548), .B(n1565), .C(n1546), .YC(n1543), .YS(n1544) );
  FAX1 U1053 ( .A(n1552), .B(n1550), .C(n1567), .YC(n1545), .YS(n1546) );
  FAX1 U1054 ( .A(n1571), .B(n1554), .C(n1569), .YC(n1547), .YS(n1548) );
  FAX1 U1055 ( .A(n1558), .B(n1560), .C(n1573), .YC(n1549), .YS(n1550) );
  FAX1 U1056 ( .A(n1577), .B(n1575), .C(n1556), .YC(n1551), .YS(n1552) );
  FAX1 U1057 ( .A(n1994), .B(n1562), .C(n1579), .YC(n1553), .YS(n1554) );
  FAX1 U1058 ( .A(n2058), .B(n1904), .C(n1932), .YC(n1555), .YS(n1556) );
  FAX1 U1059 ( .A(n1962), .B(n2122), .C(n2090), .YC(n1557), .YS(n1558) );
  FAX1 U1060 ( .A(n2026), .B(n2186), .C(n2154), .YC(n1559), .YS(n1560) );
  HAX1 U1061 ( .A(n2218), .B(n1748), .YC(n1561), .YS(n1562) );
  FAX1 U1062 ( .A(n1568), .B(n1583), .C(n1566), .YC(n1563), .YS(n1564) );
  FAX1 U1063 ( .A(n1572), .B(n1570), .C(n1585), .YC(n1565), .YS(n1566) );
  FAX1 U1064 ( .A(n1574), .B(n1589), .C(n1587), .YC(n1567), .YS(n1568) );
  FAX1 U1065 ( .A(n1580), .B(n1576), .C(n1578), .YC(n1569), .YS(n1570) );
  FAX1 U1066 ( .A(n1595), .B(n1591), .C(n1593), .YC(n1571), .YS(n1572) );
  FAX1 U1067 ( .A(n2091), .B(n2938), .C(n1597), .YC(n1573), .YS(n1574) );
  FAX1 U1068 ( .A(n2123), .B(n2027), .C(n2059), .YC(n1575), .YS(n1576) );
  FAX1 U1069 ( .A(n2155), .B(n1963), .C(n1995), .YC(n1577), .YS(n1578) );
  FAX1 U1070 ( .A(n2219), .B(n2187), .C(n1933), .YC(n1579), .YS(n1580) );
  FAX1 U1071 ( .A(n1586), .B(n1601), .C(n1584), .YC(n1581), .YS(n1582) );
  FAX1 U1072 ( .A(n1590), .B(n1588), .C(n1603), .YC(n1583), .YS(n1584) );
  FAX1 U1073 ( .A(n1596), .B(n1607), .C(n1605), .YC(n1585), .YS(n1586) );
  FAX1 U1074 ( .A(n1609), .B(n1592), .C(n1594), .YC(n1587), .YS(n1588) );
  FAX1 U1075 ( .A(n1598), .B(n1613), .C(n1611), .YC(n1589), .YS(n1590) );
  FAX1 U1076 ( .A(n2156), .B(n2028), .C(n2124), .YC(n1591), .YS(n1592) );
  FAX1 U1077 ( .A(n2092), .B(n2188), .C(n1996), .YC(n1593), .YS(n1594) );
  FAX1 U1078 ( .A(n2060), .B(n1934), .C(n1964), .YC(n1595), .YS(n1596) );
  HAX1 U1079 ( .A(n2220), .B(n1749), .YC(n1597), .YS(n1598) );
  FAX1 U1080 ( .A(n1604), .B(n1617), .C(n1602), .YC(n1599), .YS(n1600) );
  FAX1 U1081 ( .A(n1608), .B(n1606), .C(n1619), .YC(n1601), .YS(n1602) );
  FAX1 U1082 ( .A(n1612), .B(n1623), .C(n1621), .YC(n1603), .YS(n1604) );
  FAX1 U1083 ( .A(n1625), .B(n1614), .C(n1610), .YC(n1605), .YS(n1606) );
  FAX1 U1084 ( .A(n2935), .B(n1629), .C(n1627), .YC(n1607), .YS(n1608) );
  FAX1 U1085 ( .A(n2125), .B(n2061), .C(n2093), .YC(n1609), .YS(n1610) );
  FAX1 U1086 ( .A(n2157), .B(n1997), .C(n2029), .YC(n1611), .YS(n1612) );
  FAX1 U1087 ( .A(n2221), .B(n2189), .C(n1965), .YC(n1613), .YS(n1614) );
  FAX1 U1088 ( .A(n1620), .B(n1633), .C(n1618), .YC(n1615), .YS(n1616) );
  FAX1 U1089 ( .A(n1637), .B(n1622), .C(n1635), .YC(n1617), .YS(n1618) );
  FAX1 U1090 ( .A(n1628), .B(n1639), .C(n1624), .YC(n1619), .YS(n1620) );
  FAX1 U1091 ( .A(n1643), .B(n1641), .C(n1626), .YC(n1621), .YS(n1622) );
  FAX1 U1092 ( .A(n2094), .B(n2030), .C(n1630), .YC(n1623), .YS(n1624) );
  FAX1 U1093 ( .A(n2126), .B(n1966), .C(n1998), .YC(n1625), .YS(n1626) );
  FAX1 U1094 ( .A(n2062), .B(n2190), .C(n2158), .YC(n1627), .YS(n1628) );
  HAX1 U1095 ( .A(n2222), .B(n1750), .YC(n1629), .YS(n1630) );
  FAX1 U1096 ( .A(n1636), .B(n1647), .C(n1634), .YC(n1631), .YS(n1632) );
  FAX1 U1097 ( .A(n1651), .B(n1649), .C(n1638), .YC(n1633), .YS(n1634) );
  FAX1 U1098 ( .A(n1644), .B(n1642), .C(n1640), .YC(n1635), .YS(n1636) );
  FAX1 U1099 ( .A(n1657), .B(n1655), .C(n1653), .YC(n1637), .YS(n1638) );
  FAX1 U1100 ( .A(n2127), .B(n2095), .C(n2929), .YC(n1639), .YS(n1640) );
  FAX1 U1101 ( .A(n2159), .B(n2031), .C(n2063), .YC(n1641), .YS(n1642) );
  FAX1 U1102 ( .A(n2223), .B(n2191), .C(n1999), .YC(n1643), .YS(n1644) );
  FAX1 U1103 ( .A(n1650), .B(n1661), .C(n1648), .YC(n1645), .YS(n1646) );
  FAX1 U1104 ( .A(n1665), .B(n1663), .C(n1652), .YC(n1647), .YS(n1648) );
  FAX1 U1105 ( .A(n1667), .B(n1654), .C(n1656), .YC(n1649), .YS(n1650) );
  FAX1 U1106 ( .A(n2160), .B(n1658), .C(n1669), .YC(n1651), .YS(n1652) );
  FAX1 U1107 ( .A(n2192), .B(n2064), .C(n2128), .YC(n1653), .YS(n1654) );
  FAX1 U1108 ( .A(n2096), .B(n2000), .C(n2032), .YC(n1655), .YS(n1656) );
  HAX1 U1109 ( .A(n2224), .B(n1751), .YC(n1657), .YS(n1658) );
  FAX1 U1110 ( .A(n1664), .B(n1673), .C(n1662), .YC(n1659), .YS(n1660) );
  FAX1 U1111 ( .A(n1668), .B(n1666), .C(n1675), .YC(n1661), .YS(n1662) );
  FAX1 U1112 ( .A(n1679), .B(n1677), .C(n1670), .YC(n1663), .YS(n1664) );
  FAX1 U1113 ( .A(n2129), .B(n2936), .C(n1681), .YC(n1665), .YS(n1666) );
  FAX1 U1114 ( .A(n2161), .B(n2065), .C(n2097), .YC(n1667), .YS(n1668) );
  FAX1 U1115 ( .A(n2225), .B(n2193), .C(n2033), .YC(n1669), .YS(n1670) );
  FAX1 U1116 ( .A(n1676), .B(n1685), .C(n1674), .YC(n1671), .YS(n1672) );
  FAX1 U1117 ( .A(n1678), .B(n1680), .C(n1687), .YC(n1673), .YS(n1674) );
  FAX1 U1118 ( .A(n1682), .B(n1691), .C(n1689), .YC(n1675), .YS(n1676) );
  FAX1 U1119 ( .A(n2130), .B(n2034), .C(n2066), .YC(n1677), .YS(n1678) );
  FAX1 U1120 ( .A(n2098), .B(n2194), .C(n2162), .YC(n1679), .YS(n1680) );
  HAX1 U1121 ( .A(n2226), .B(n1752), .YC(n1681), .YS(n1682) );
  FAX1 U1122 ( .A(n1688), .B(n1695), .C(n1686), .YC(n1683), .YS(n1684) );
  FAX1 U1123 ( .A(n1692), .B(n1690), .C(n1697), .YC(n1685), .YS(n1686) );
  FAX1 U1124 ( .A(n2939), .B(n1701), .C(n1699), .YC(n1687), .YS(n1688) );
  FAX1 U1125 ( .A(n2163), .B(n2099), .C(n2131), .YC(n1689), .YS(n1690) );
  FAX1 U1126 ( .A(n2227), .B(n2195), .C(n2067), .YC(n1691), .YS(n1692) );
  FAX1 U1127 ( .A(n1698), .B(n1705), .C(n1696), .YC(n1693), .YS(n1694) );
  FAX1 U1128 ( .A(n1709), .B(n1700), .C(n1707), .YC(n1695), .YS(n1696) );
  FAX1 U1129 ( .A(n2164), .B(n2100), .C(n1702), .YC(n1697), .YS(n1698) );
  FAX1 U1130 ( .A(n2132), .B(n2068), .C(n2196), .YC(n1699), .YS(n1700) );
  HAX1 U1131 ( .A(n2228), .B(n1753), .YC(n1701), .YS(n1702) );
  FAX1 U1132 ( .A(n1708), .B(n1713), .C(n1706), .YC(n1703), .YS(n1704) );
  FAX1 U1133 ( .A(n1717), .B(n1715), .C(n1710), .YC(n1705), .YS(n1706) );
  FAX1 U1134 ( .A(n2165), .B(n2133), .C(n2069), .YC(n1707), .YS(n1708) );
  FAX1 U1135 ( .A(n2229), .B(n2197), .C(n2101), .YC(n1709), .YS(n1710) );
  FAX1 U1136 ( .A(n1716), .B(n1721), .C(n1714), .YC(n1711), .YS(n1712) );
  FAX1 U1137 ( .A(n2198), .B(n1718), .C(n1723), .YC(n1713), .YS(n1714) );
  FAX1 U1138 ( .A(n2134), .B(n2102), .C(n2166), .YC(n1715), .YS(n1716) );
  HAX1 U1139 ( .A(n2230), .B(n1754), .YC(n1717), .YS(n1718) );
  FAX1 U1140 ( .A(n1727), .B(n1724), .C(n1722), .YC(n1719), .YS(n1720) );
  FAX1 U1141 ( .A(n2167), .B(n2941), .C(n1729), .YC(n1721), .YS(n1722) );
  FAX1 U1142 ( .A(n2231), .B(n2199), .C(n2135), .YC(n1723), .YS(n1724) );
  FAX1 U1143 ( .A(n1730), .B(n1733), .C(n1728), .YC(n1725), .YS(n1726) );
  FAX1 U1144 ( .A(n2200), .B(n2136), .C(n2168), .YC(n1727), .YS(n1728) );
  HAX1 U1145 ( .A(n2232), .B(n1755), .YC(n1729), .YS(n1730) );
  FAX1 U1146 ( .A(n2943), .B(n1737), .C(n1734), .YC(n1731), .YS(n1732) );
  FAX1 U1147 ( .A(n2233), .B(n2201), .C(n2169), .YC(n1733), .YS(n1734) );
  FAX1 U1148 ( .A(n2202), .B(n2170), .C(n1738), .YC(n1735), .YS(n1736) );
  HAX1 U1149 ( .A(n2234), .B(n1756), .YC(n1737), .YS(n1738) );
  FAX1 U1150 ( .A(n2235), .B(n2203), .C(n2171), .YC(n1739), .YS(n1740) );
  HAX1 U1151 ( .A(n2236), .B(n2204), .YC(n1741), .YS(n1742) );
  NOR2X1 U1152 ( .A(n2239), .B(n383), .Y(n1759) );
  NOR2X1 U1153 ( .A(n2240), .B(n383), .Y(n918) );
  NOR2X1 U1154 ( .A(n2241), .B(n383), .Y(n1760) );
  NOR2X1 U1155 ( .A(n2242), .B(n383), .Y(n960) );
  NOR2X1 U1156 ( .A(n2243), .B(n383), .Y(n1761) );
  NOR2X1 U1157 ( .A(n2244), .B(n383), .Y(n1006) );
  NOR2X1 U1158 ( .A(n2245), .B(n383), .Y(n1762) );
  NOR2X1 U1159 ( .A(n2246), .B(n383), .Y(n1056) );
  NOR2X1 U1160 ( .A(n2247), .B(n383), .Y(n1763) );
  NOR2X1 U1161 ( .A(n2248), .B(n383), .Y(n1110) );
  NOR2X1 U1162 ( .A(n2249), .B(n383), .Y(n1764) );
  NOR2X1 U1163 ( .A(n2250), .B(n383), .Y(n1168) );
  NOR2X1 U1164 ( .A(n2251), .B(n383), .Y(n1765) );
  NOR2X1 U1165 ( .A(n2252), .B(n383), .Y(n1766) );
  NOR2X1 U1166 ( .A(n2253), .B(n383), .Y(n1230) );
  INVX2 U1167 ( .A(n465), .Y(n2239) );
  INVX2 U1168 ( .A(n463), .Y(n2240) );
  INVX2 U1169 ( .A(n461), .Y(n2241) );
  INVX2 U1170 ( .A(n459), .Y(n2242) );
  INVX2 U1171 ( .A(n457), .Y(n2243) );
  INVX2 U1172 ( .A(n455), .Y(n2244) );
  INVX2 U1173 ( .A(n453), .Y(n2245) );
  INVX2 U1174 ( .A(n451), .Y(n2246) );
  INVX2 U1175 ( .A(n449), .Y(n2247) );
  INVX2 U1176 ( .A(n447), .Y(n2248) );
  INVX2 U1177 ( .A(n445), .Y(n2249) );
  INVX2 U1178 ( .A(n443), .Y(n2250) );
  INVX2 U1179 ( .A(n441), .Y(n2251) );
  INVX2 U1180 ( .A(n439), .Y(n2252) );
  INVX2 U1181 ( .A(n437), .Y(n2253) );
  OAI22X1 U1182 ( .A(n382), .B(n2272), .C(n2796), .D(n432), .Y(n1743) );
  OAI22X1 U1183 ( .A(n2254), .B(n381), .C(n2255), .D(n431), .Y(n1768) );
  OAI22X1 U1184 ( .A(n2255), .B(n381), .C(n2256), .D(n431), .Y(n1769) );
  OAI22X1 U1185 ( .A(n2256), .B(n381), .C(n2257), .D(n431), .Y(n1770) );
  OAI22X1 U1186 ( .A(n2257), .B(n381), .C(n2258), .D(n431), .Y(n1771) );
  OAI22X1 U1187 ( .A(n2258), .B(n381), .C(n2259), .D(n431), .Y(n1772) );
  OAI22X1 U1188 ( .A(n2259), .B(n381), .C(n2260), .D(n431), .Y(n1773) );
  OAI22X1 U1189 ( .A(n2260), .B(n380), .C(n2261), .D(n431), .Y(n1774) );
  OAI22X1 U1190 ( .A(n2261), .B(n380), .C(n2262), .D(n430), .Y(n1775) );
  OAI22X1 U1191 ( .A(n2262), .B(n380), .C(n2263), .D(n430), .Y(n1776) );
  OAI22X1 U1192 ( .A(n2263), .B(n380), .C(n2264), .D(n430), .Y(n1777) );
  OAI22X1 U1193 ( .A(n2264), .B(n380), .C(n2265), .D(n430), .Y(n1778) );
  OAI22X1 U1194 ( .A(n2265), .B(n380), .C(n2266), .D(n430), .Y(n1779) );
  OAI22X1 U1195 ( .A(n2266), .B(n380), .C(n2267), .D(n430), .Y(n1780) );
  OAI22X1 U1196 ( .A(n2267), .B(n380), .C(n2268), .D(n430), .Y(n1781) );
  OAI22X1 U1197 ( .A(n2268), .B(n380), .C(n2269), .D(n430), .Y(n1782) );
  OAI22X1 U1198 ( .A(n2269), .B(n380), .C(n2270), .D(n430), .Y(n1783) );
  OAI22X1 U1199 ( .A(n2270), .B(n380), .C(n2271), .D(n430), .Y(n1784) );
  XNOR2X1 U1200 ( .A(n333), .B(n469), .Y(n2254) );
  XNOR2X1 U1201 ( .A(n333), .B(n467), .Y(n2255) );
  XNOR2X1 U1202 ( .A(n333), .B(n465), .Y(n2256) );
  XNOR2X1 U1203 ( .A(n333), .B(n463), .Y(n2257) );
  XNOR2X1 U1204 ( .A(n333), .B(n461), .Y(n2258) );
  XNOR2X1 U1205 ( .A(n333), .B(n459), .Y(n2259) );
  XNOR2X1 U1206 ( .A(n333), .B(n457), .Y(n2260) );
  XNOR2X1 U1207 ( .A(n333), .B(n455), .Y(n2261) );
  XNOR2X1 U1208 ( .A(n333), .B(n453), .Y(n2262) );
  XNOR2X1 U1209 ( .A(n332), .B(n451), .Y(n2263) );
  XNOR2X1 U1210 ( .A(n332), .B(n449), .Y(n2264) );
  XNOR2X1 U1211 ( .A(n332), .B(n447), .Y(n2265) );
  XNOR2X1 U1212 ( .A(n332), .B(n445), .Y(n2266) );
  XNOR2X1 U1213 ( .A(n332), .B(n443), .Y(n2267) );
  XNOR2X1 U1214 ( .A(n332), .B(n441), .Y(n2268) );
  XNOR2X1 U1215 ( .A(n332), .B(n439), .Y(n2269) );
  XNOR2X1 U1216 ( .A(n332), .B(n437), .Y(n2270) );
  XNOR2X1 U1217 ( .A(n332), .B(n2951), .Y(n2271) );
  OAI22X1 U1218 ( .A(n379), .B(n2293), .C(n2797), .D(n429), .Y(n1744) );
  OAI22X1 U1219 ( .A(n2273), .B(n378), .C(n2274), .D(n428), .Y(n1786) );
  OAI22X1 U1220 ( .A(n2274), .B(n378), .C(n2275), .D(n428), .Y(n1787) );
  OAI22X1 U1221 ( .A(n2275), .B(n378), .C(n2276), .D(n428), .Y(n1788) );
  OAI22X1 U1222 ( .A(n2276), .B(n378), .C(n2277), .D(n428), .Y(n1789) );
  OAI22X1 U1223 ( .A(n2277), .B(n378), .C(n2278), .D(n428), .Y(n1790) );
  OAI22X1 U1224 ( .A(n2278), .B(n378), .C(n2279), .D(n428), .Y(n1791) );
  OAI22X1 U1225 ( .A(n2279), .B(n378), .C(n2280), .D(n428), .Y(n1792) );
  OAI22X1 U1226 ( .A(n2280), .B(n378), .C(n2281), .D(n428), .Y(n1793) );
  OAI22X1 U1227 ( .A(n2281), .B(n377), .C(n2282), .D(n428), .Y(n1794) );
  OAI22X1 U1228 ( .A(n2282), .B(n377), .C(n2283), .D(n427), .Y(n1795) );
  OAI22X1 U1229 ( .A(n2283), .B(n377), .C(n2284), .D(n427), .Y(n1796) );
  OAI22X1 U1230 ( .A(n2284), .B(n377), .C(n2285), .D(n427), .Y(n1797) );
  OAI22X1 U1231 ( .A(n2285), .B(n377), .C(n2286), .D(n427), .Y(n1798) );
  OAI22X1 U1232 ( .A(n2286), .B(n377), .C(n2287), .D(n427), .Y(n1799) );
  OAI22X1 U1233 ( .A(n2287), .B(n377), .C(n2288), .D(n427), .Y(n1800) );
  OAI22X1 U1234 ( .A(n2288), .B(n377), .C(n2289), .D(n427), .Y(n1801) );
  OAI22X1 U1235 ( .A(n2289), .B(n377), .C(n2290), .D(n427), .Y(n1802) );
  OAI22X1 U1236 ( .A(n2290), .B(n377), .C(n2291), .D(n427), .Y(n1803) );
  OAI22X1 U1237 ( .A(n2291), .B(n377), .C(n2292), .D(n427), .Y(n1804) );
  XNOR2X1 U1238 ( .A(n330), .B(n473), .Y(n2273) );
  XNOR2X1 U1239 ( .A(n330), .B(n471), .Y(n2274) );
  XNOR2X1 U1240 ( .A(n330), .B(n469), .Y(n2275) );
  XNOR2X1 U1241 ( .A(n330), .B(n467), .Y(n2276) );
  XNOR2X1 U1242 ( .A(n330), .B(n465), .Y(n2277) );
  XNOR2X1 U1243 ( .A(n330), .B(n463), .Y(n2278) );
  XNOR2X1 U1244 ( .A(n330), .B(n461), .Y(n2279) );
  XNOR2X1 U1245 ( .A(n330), .B(n459), .Y(n2280) );
  XNOR2X1 U1246 ( .A(n330), .B(n457), .Y(n2281) );
  XNOR2X1 U1247 ( .A(n330), .B(n455), .Y(n2282) );
  XNOR2X1 U1248 ( .A(n330), .B(n453), .Y(n2283) );
  XNOR2X1 U1249 ( .A(n329), .B(n451), .Y(n2284) );
  XNOR2X1 U1250 ( .A(n329), .B(n449), .Y(n2285) );
  XNOR2X1 U1251 ( .A(n329), .B(n447), .Y(n2286) );
  XNOR2X1 U1252 ( .A(n329), .B(n445), .Y(n2287) );
  XNOR2X1 U1253 ( .A(n329), .B(n443), .Y(n2288) );
  XNOR2X1 U1254 ( .A(n329), .B(n441), .Y(n2289) );
  XNOR2X1 U1255 ( .A(n329), .B(n439), .Y(n2290) );
  XNOR2X1 U1256 ( .A(n329), .B(n437), .Y(n2291) );
  XNOR2X1 U1257 ( .A(n329), .B(n2950), .Y(n2292) );
  OAI22X1 U1258 ( .A(n376), .B(n2316), .C(n2798), .D(n426), .Y(n1745) );
  OAI22X1 U1259 ( .A(n2294), .B(n375), .C(n2295), .D(n425), .Y(n1806) );
  OAI22X1 U1260 ( .A(n2295), .B(n375), .C(n2296), .D(n425), .Y(n1807) );
  OAI22X1 U1261 ( .A(n2296), .B(n375), .C(n2297), .D(n425), .Y(n1808) );
  OAI22X1 U1262 ( .A(n2297), .B(n375), .C(n2298), .D(n425), .Y(n1809) );
  OAI22X1 U1263 ( .A(n2298), .B(n375), .C(n2299), .D(n425), .Y(n1810) );
  OAI22X1 U1264 ( .A(n2299), .B(n375), .C(n2300), .D(n425), .Y(n1811) );
  OAI22X1 U1265 ( .A(n2300), .B(n375), .C(n2301), .D(n425), .Y(n1812) );
  OAI22X1 U1266 ( .A(n2301), .B(n375), .C(n2302), .D(n425), .Y(n1813) );
  OAI22X1 U1267 ( .A(n2302), .B(n375), .C(n2303), .D(n425), .Y(n1814) );
  OAI22X1 U1268 ( .A(n2303), .B(n375), .C(n2304), .D(n425), .Y(n1815) );
  OAI22X1 U1269 ( .A(n2304), .B(n374), .C(n2305), .D(n425), .Y(n1816) );
  OAI22X1 U1270 ( .A(n2305), .B(n374), .C(n2306), .D(n424), .Y(n1817) );
  OAI22X1 U1271 ( .A(n2306), .B(n374), .C(n2307), .D(n424), .Y(n1818) );
  OAI22X1 U1272 ( .A(n2307), .B(n374), .C(n2308), .D(n424), .Y(n1819) );
  OAI22X1 U1273 ( .A(n2308), .B(n374), .C(n2309), .D(n424), .Y(n1820) );
  OAI22X1 U1274 ( .A(n2309), .B(n374), .C(n2310), .D(n424), .Y(n1821) );
  OAI22X1 U1275 ( .A(n2310), .B(n374), .C(n2311), .D(n424), .Y(n1822) );
  OAI22X1 U1276 ( .A(n2311), .B(n374), .C(n2312), .D(n424), .Y(n1823) );
  OAI22X1 U1277 ( .A(n2312), .B(n374), .C(n2313), .D(n424), .Y(n1824) );
  OAI22X1 U1278 ( .A(n2313), .B(n374), .C(n2314), .D(n424), .Y(n1825) );
  OAI22X1 U1279 ( .A(n2314), .B(n374), .C(n2315), .D(n424), .Y(n1826) );
  XNOR2X1 U1280 ( .A(n328), .B(n477), .Y(n2294) );
  XNOR2X1 U1281 ( .A(n327), .B(n475), .Y(n2295) );
  XNOR2X1 U1282 ( .A(n327), .B(n473), .Y(n2296) );
  XNOR2X1 U1283 ( .A(n327), .B(n471), .Y(n2297) );
  XNOR2X1 U1284 ( .A(n327), .B(n469), .Y(n2298) );
  XNOR2X1 U1285 ( .A(n327), .B(n467), .Y(n2299) );
  XNOR2X1 U1286 ( .A(n327), .B(n465), .Y(n2300) );
  XNOR2X1 U1287 ( .A(n327), .B(n463), .Y(n2301) );
  XNOR2X1 U1288 ( .A(n327), .B(n461), .Y(n2302) );
  XNOR2X1 U1289 ( .A(n327), .B(n459), .Y(n2303) );
  XNOR2X1 U1290 ( .A(n327), .B(n457), .Y(n2304) );
  XNOR2X1 U1291 ( .A(n327), .B(n455), .Y(n2305) );
  XNOR2X1 U1292 ( .A(n327), .B(n453), .Y(n2306) );
  XNOR2X1 U1293 ( .A(n326), .B(n451), .Y(n2307) );
  XNOR2X1 U1294 ( .A(n326), .B(n449), .Y(n2308) );
  XNOR2X1 U1295 ( .A(n326), .B(n447), .Y(n2309) );
  XNOR2X1 U1296 ( .A(n326), .B(n445), .Y(n2310) );
  XNOR2X1 U1297 ( .A(n326), .B(n443), .Y(n2311) );
  XNOR2X1 U1298 ( .A(n326), .B(n441), .Y(n2312) );
  XNOR2X1 U1299 ( .A(n326), .B(n439), .Y(n2313) );
  XNOR2X1 U1300 ( .A(n326), .B(n437), .Y(n2314) );
  XNOR2X1 U1301 ( .A(n326), .B(n2951), .Y(n2315) );
  OAI22X1 U1302 ( .A(n373), .B(n2341), .C(n2799), .D(n423), .Y(n1746) );
  OAI22X1 U1303 ( .A(n2317), .B(n372), .C(n2318), .D(n423), .Y(n1828) );
  OAI22X1 U1304 ( .A(n2318), .B(n372), .C(n2319), .D(n422), .Y(n1829) );
  OAI22X1 U1305 ( .A(n2319), .B(n372), .C(n2320), .D(n422), .Y(n1830) );
  OAI22X1 U1306 ( .A(n2320), .B(n372), .C(n2321), .D(n422), .Y(n1831) );
  OAI22X1 U1307 ( .A(n2321), .B(n372), .C(n2322), .D(n422), .Y(n1832) );
  OAI22X1 U1308 ( .A(n2322), .B(n372), .C(n2323), .D(n422), .Y(n1833) );
  OAI22X1 U1309 ( .A(n2323), .B(n372), .C(n2324), .D(n422), .Y(n1834) );
  OAI22X1 U1310 ( .A(n2324), .B(n372), .C(n2325), .D(n422), .Y(n1835) );
  OAI22X1 U1311 ( .A(n2325), .B(n372), .C(n2326), .D(n422), .Y(n1836) );
  OAI22X1 U1312 ( .A(n2326), .B(n372), .C(n2327), .D(n422), .Y(n1837) );
  OAI22X1 U1313 ( .A(n2327), .B(n372), .C(n2328), .D(n422), .Y(n1838) );
  OAI22X1 U1314 ( .A(n2328), .B(n372), .C(n2329), .D(n422), .Y(n1839) );
  OAI22X1 U1315 ( .A(n2329), .B(n371), .C(n2330), .D(n422), .Y(n1840) );
  OAI22X1 U1316 ( .A(n2330), .B(n371), .C(n2331), .D(n421), .Y(n1841) );
  OAI22X1 U1317 ( .A(n2331), .B(n371), .C(n2332), .D(n421), .Y(n1842) );
  OAI22X1 U1318 ( .A(n2332), .B(n371), .C(n2333), .D(n421), .Y(n1843) );
  OAI22X1 U1319 ( .A(n2333), .B(n371), .C(n2334), .D(n421), .Y(n1844) );
  OAI22X1 U1320 ( .A(n2334), .B(n371), .C(n2335), .D(n421), .Y(n1845) );
  OAI22X1 U1321 ( .A(n2335), .B(n371), .C(n2336), .D(n421), .Y(n1846) );
  OAI22X1 U1322 ( .A(n2336), .B(n371), .C(n2337), .D(n421), .Y(n1847) );
  OAI22X1 U1323 ( .A(n2337), .B(n371), .C(n2338), .D(n421), .Y(n1848) );
  OAI22X1 U1324 ( .A(n2338), .B(n371), .C(n2339), .D(n421), .Y(n1849) );
  OAI22X1 U1325 ( .A(n2339), .B(n371), .C(n2340), .D(n421), .Y(n1850) );
  XNOR2X1 U1326 ( .A(n325), .B(n2913), .Y(n2317) );
  XNOR2X1 U1327 ( .A(n325), .B(n2909), .Y(n2318) );
  XNOR2X1 U1328 ( .A(n325), .B(n477), .Y(n2319) );
  XNOR2X1 U1329 ( .A(n324), .B(n475), .Y(n2320) );
  XNOR2X1 U1330 ( .A(n324), .B(n473), .Y(n2321) );
  XNOR2X1 U1331 ( .A(n324), .B(n471), .Y(n2322) );
  XNOR2X1 U1332 ( .A(n324), .B(n469), .Y(n2323) );
  XNOR2X1 U1333 ( .A(n324), .B(n467), .Y(n2324) );
  XNOR2X1 U1334 ( .A(n324), .B(n465), .Y(n2325) );
  XNOR2X1 U1335 ( .A(n324), .B(n463), .Y(n2326) );
  XNOR2X1 U1336 ( .A(n324), .B(n461), .Y(n2327) );
  XNOR2X1 U1337 ( .A(n324), .B(n459), .Y(n2328) );
  XNOR2X1 U1338 ( .A(n324), .B(n457), .Y(n2329) );
  XNOR2X1 U1339 ( .A(n324), .B(n455), .Y(n2330) );
  XNOR2X1 U1340 ( .A(n324), .B(n453), .Y(n2331) );
  XNOR2X1 U1341 ( .A(n323), .B(n451), .Y(n2332) );
  XNOR2X1 U1342 ( .A(n323), .B(n449), .Y(n2333) );
  XNOR2X1 U1343 ( .A(n323), .B(n447), .Y(n2334) );
  XNOR2X1 U1344 ( .A(n323), .B(n445), .Y(n2335) );
  XNOR2X1 U1345 ( .A(n323), .B(n443), .Y(n2336) );
  XNOR2X1 U1346 ( .A(n323), .B(n441), .Y(n2337) );
  XNOR2X1 U1347 ( .A(n323), .B(n439), .Y(n2338) );
  XNOR2X1 U1348 ( .A(n323), .B(n437), .Y(n2339) );
  XNOR2X1 U1349 ( .A(n323), .B(n2951), .Y(n2340) );
  OAI22X1 U1350 ( .A(n370), .B(n2368), .C(n2800), .D(n420), .Y(n1747) );
  OAI22X1 U1351 ( .A(n2342), .B(n370), .C(n2343), .D(n420), .Y(n1852) );
  OAI22X1 U1352 ( .A(n2343), .B(n370), .C(n2344), .D(n420), .Y(n1853) );
  OAI22X1 U1353 ( .A(n2344), .B(n369), .C(n2345), .D(n420), .Y(n1854) );
  OAI22X1 U1354 ( .A(n2345), .B(n369), .C(n2346), .D(n419), .Y(n1855) );
  OAI22X1 U1355 ( .A(n2346), .B(n369), .C(n2347), .D(n419), .Y(n1856) );
  OAI22X1 U1356 ( .A(n2347), .B(n369), .C(n2348), .D(n419), .Y(n1857) );
  OAI22X1 U1357 ( .A(n2348), .B(n369), .C(n2349), .D(n419), .Y(n1858) );
  OAI22X1 U1358 ( .A(n2349), .B(n369), .C(n2350), .D(n419), .Y(n1859) );
  OAI22X1 U1359 ( .A(n2350), .B(n369), .C(n2351), .D(n419), .Y(n1860) );
  OAI22X1 U1360 ( .A(n2351), .B(n369), .C(n2352), .D(n419), .Y(n1861) );
  OAI22X1 U1361 ( .A(n2352), .B(n369), .C(n2353), .D(n419), .Y(n1862) );
  OAI22X1 U1362 ( .A(n2353), .B(n369), .C(n2354), .D(n419), .Y(n1863) );
  OAI22X1 U1363 ( .A(n2354), .B(n369), .C(n2355), .D(n419), .Y(n1864) );
  OAI22X1 U1364 ( .A(n2355), .B(n369), .C(n2356), .D(n419), .Y(n1865) );
  OAI22X1 U1365 ( .A(n2356), .B(n368), .C(n2357), .D(n419), .Y(n1866) );
  OAI22X1 U1366 ( .A(n2357), .B(n368), .C(n2358), .D(n418), .Y(n1867) );
  OAI22X1 U1367 ( .A(n2358), .B(n368), .C(n2359), .D(n418), .Y(n1868) );
  OAI22X1 U1368 ( .A(n2359), .B(n368), .C(n2360), .D(n418), .Y(n1869) );
  OAI22X1 U1369 ( .A(n2360), .B(n368), .C(n2361), .D(n418), .Y(n1870) );
  OAI22X1 U1370 ( .A(n2361), .B(n368), .C(n2362), .D(n418), .Y(n1871) );
  OAI22X1 U1371 ( .A(n2362), .B(n368), .C(n2363), .D(n418), .Y(n1872) );
  OAI22X1 U1372 ( .A(n2363), .B(n368), .C(n2364), .D(n418), .Y(n1873) );
  OAI22X1 U1373 ( .A(n2364), .B(n368), .C(n2365), .D(n418), .Y(n1874) );
  OAI22X1 U1374 ( .A(n2365), .B(n368), .C(n2366), .D(n418), .Y(n1875) );
  OAI22X1 U1375 ( .A(n2366), .B(n368), .C(n2367), .D(n418), .Y(n1876) );
  XNOR2X1 U1376 ( .A(n322), .B(n485), .Y(n2342) );
  XNOR2X1 U1377 ( .A(n322), .B(n483), .Y(n2343) );
  XNOR2X1 U1378 ( .A(n322), .B(n2913), .Y(n2344) );
  XNOR2X1 U1379 ( .A(n322), .B(n2909), .Y(n2345) );
  XNOR2X1 U1380 ( .A(n322), .B(n477), .Y(n2346) );
  XNOR2X1 U1381 ( .A(n321), .B(n475), .Y(n2347) );
  XNOR2X1 U1382 ( .A(n321), .B(n473), .Y(n2348) );
  XNOR2X1 U1383 ( .A(n321), .B(n471), .Y(n2349) );
  XNOR2X1 U1384 ( .A(n321), .B(n469), .Y(n2350) );
  XNOR2X1 U1385 ( .A(n321), .B(n467), .Y(n2351) );
  XNOR2X1 U1386 ( .A(n321), .B(n465), .Y(n2352) );
  XNOR2X1 U1387 ( .A(n321), .B(n463), .Y(n2353) );
  XNOR2X1 U1388 ( .A(n321), .B(n461), .Y(n2354) );
  XNOR2X1 U1389 ( .A(n321), .B(n459), .Y(n2355) );
  XNOR2X1 U1390 ( .A(n321), .B(n457), .Y(n2356) );
  XNOR2X1 U1391 ( .A(n321), .B(n455), .Y(n2357) );
  XNOR2X1 U1392 ( .A(n321), .B(n453), .Y(n2358) );
  XNOR2X1 U1393 ( .A(n320), .B(n451), .Y(n2359) );
  XNOR2X1 U1394 ( .A(n320), .B(n449), .Y(n2360) );
  XNOR2X1 U1395 ( .A(n320), .B(n447), .Y(n2361) );
  XNOR2X1 U1396 ( .A(n320), .B(n445), .Y(n2362) );
  XNOR2X1 U1397 ( .A(n320), .B(n443), .Y(n2363) );
  XNOR2X1 U1398 ( .A(n320), .B(n441), .Y(n2364) );
  XNOR2X1 U1399 ( .A(n320), .B(n439), .Y(n2365) );
  XNOR2X1 U1400 ( .A(n320), .B(n437), .Y(n2366) );
  XNOR2X1 U1401 ( .A(n320), .B(n2951), .Y(n2367) );
  OAI22X1 U1402 ( .A(n367), .B(n2397), .C(n2801), .D(n417), .Y(n1748) );
  OAI22X1 U1403 ( .A(n2369), .B(n367), .C(n2370), .D(n417), .Y(n1878) );
  OAI22X1 U1404 ( .A(n2370), .B(n367), .C(n2371), .D(n417), .Y(n1879) );
  OAI22X1 U1405 ( .A(n2371), .B(n367), .C(n2372), .D(n417), .Y(n1880) );
  OAI22X1 U1406 ( .A(n2372), .B(n367), .C(n2373), .D(n417), .Y(n1881) );
  OAI22X1 U1407 ( .A(n2373), .B(n366), .C(n2374), .D(n417), .Y(n1882) );
  OAI22X1 U1408 ( .A(n2374), .B(n366), .C(n2375), .D(n416), .Y(n1883) );
  OAI22X1 U1409 ( .A(n2375), .B(n366), .C(n2376), .D(n416), .Y(n1884) );
  OAI22X1 U1410 ( .A(n2376), .B(n366), .C(n2377), .D(n416), .Y(n1885) );
  OAI22X1 U1411 ( .A(n2377), .B(n366), .C(n2378), .D(n416), .Y(n1886) );
  OAI22X1 U1412 ( .A(n2378), .B(n366), .C(n2379), .D(n416), .Y(n1887) );
  OAI22X1 U1413 ( .A(n2379), .B(n366), .C(n2380), .D(n416), .Y(n1888) );
  OAI22X1 U1414 ( .A(n2380), .B(n366), .C(n2381), .D(n416), .Y(n1889) );
  OAI22X1 U1415 ( .A(n2381), .B(n366), .C(n2382), .D(n416), .Y(n1890) );
  OAI22X1 U1416 ( .A(n2382), .B(n366), .C(n2383), .D(n416), .Y(n1891) );
  OAI22X1 U1417 ( .A(n2383), .B(n366), .C(n2384), .D(n416), .Y(n1892) );
  OAI22X1 U1418 ( .A(n2384), .B(n366), .C(n2385), .D(n416), .Y(n1893) );
  OAI22X1 U1419 ( .A(n2385), .B(n365), .C(n2386), .D(n416), .Y(n1894) );
  OAI22X1 U1420 ( .A(n2386), .B(n365), .C(n2387), .D(n415), .Y(n1895) );
  OAI22X1 U1421 ( .A(n2387), .B(n365), .C(n2388), .D(n415), .Y(n1896) );
  OAI22X1 U1422 ( .A(n2388), .B(n365), .C(n2389), .D(n415), .Y(n1897) );
  OAI22X1 U1423 ( .A(n2389), .B(n365), .C(n2390), .D(n415), .Y(n1898) );
  OAI22X1 U1424 ( .A(n2390), .B(n365), .C(n2391), .D(n415), .Y(n1899) );
  OAI22X1 U1425 ( .A(n2391), .B(n365), .C(n2392), .D(n415), .Y(n1900) );
  OAI22X1 U1426 ( .A(n2392), .B(n365), .C(n2393), .D(n415), .Y(n1901) );
  OAI22X1 U1427 ( .A(n2393), .B(n365), .C(n2394), .D(n415), .Y(n1902) );
  OAI22X1 U1428 ( .A(n2394), .B(n365), .C(n2395), .D(n415), .Y(n1903) );
  OAI22X1 U1429 ( .A(n2395), .B(n365), .C(n2396), .D(n415), .Y(n1904) );
  XNOR2X1 U1430 ( .A(n319), .B(n2947), .Y(n2369) );
  XNOR2X1 U1431 ( .A(n319), .B(n2949), .Y(n2370) );
  XNOR2X1 U1432 ( .A(n319), .B(n485), .Y(n2371) );
  XNOR2X1 U1433 ( .A(n319), .B(n483), .Y(n2372) );
  XNOR2X1 U1434 ( .A(n319), .B(n2913), .Y(n2373) );
  XNOR2X1 U1435 ( .A(n319), .B(n479), .Y(n2374) );
  XNOR2X1 U1436 ( .A(n319), .B(n477), .Y(n2375) );
  XNOR2X1 U1437 ( .A(n318), .B(n475), .Y(n2376) );
  XNOR2X1 U1438 ( .A(n318), .B(n473), .Y(n2377) );
  XNOR2X1 U1439 ( .A(n318), .B(n471), .Y(n2378) );
  XNOR2X1 U1440 ( .A(n318), .B(n469), .Y(n2379) );
  XNOR2X1 U1441 ( .A(n318), .B(n467), .Y(n2380) );
  XNOR2X1 U1442 ( .A(n318), .B(n465), .Y(n2381) );
  XNOR2X1 U1443 ( .A(n318), .B(n463), .Y(n2382) );
  XNOR2X1 U1444 ( .A(n318), .B(n461), .Y(n2383) );
  XNOR2X1 U1445 ( .A(n318), .B(n459), .Y(n2384) );
  XNOR2X1 U1446 ( .A(n318), .B(n457), .Y(n2385) );
  XNOR2X1 U1447 ( .A(n318), .B(n455), .Y(n2386) );
  XNOR2X1 U1448 ( .A(n318), .B(n453), .Y(n2387) );
  XNOR2X1 U1449 ( .A(n317), .B(n451), .Y(n2388) );
  XNOR2X1 U1450 ( .A(n317), .B(n449), .Y(n2389) );
  XNOR2X1 U1451 ( .A(n317), .B(n447), .Y(n2390) );
  XNOR2X1 U1452 ( .A(n317), .B(n445), .Y(n2391) );
  XNOR2X1 U1453 ( .A(n317), .B(n443), .Y(n2392) );
  XNOR2X1 U1454 ( .A(n317), .B(n441), .Y(n2393) );
  XNOR2X1 U1455 ( .A(n317), .B(n439), .Y(n2394) );
  XNOR2X1 U1456 ( .A(n317), .B(n437), .Y(n2395) );
  XNOR2X1 U1457 ( .A(n317), .B(n2950), .Y(n2396) );
  OAI22X1 U1458 ( .A(n364), .B(n2428), .C(n2802), .D(n414), .Y(n1749) );
  OAI22X1 U1459 ( .A(n2398), .B(n364), .C(n2399), .D(n414), .Y(n1906) );
  OAI22X1 U1460 ( .A(n2399), .B(n364), .C(n2400), .D(n414), .Y(n1907) );
  OAI22X1 U1461 ( .A(n2400), .B(n364), .C(n2401), .D(n414), .Y(n1908) );
  OAI22X1 U1462 ( .A(n2401), .B(n364), .C(n2402), .D(n414), .Y(n1909) );
  OAI22X1 U1463 ( .A(n2402), .B(n364), .C(n2403), .D(n414), .Y(n1910) );
  OAI22X1 U1464 ( .A(n2403), .B(n364), .C(n2404), .D(n414), .Y(n1911) );
  OAI22X1 U1465 ( .A(n2404), .B(n363), .C(n2405), .D(n414), .Y(n1912) );
  OAI22X1 U1466 ( .A(n2405), .B(n363), .C(n2406), .D(n413), .Y(n1913) );
  OAI22X1 U1467 ( .A(n2406), .B(n363), .C(n2407), .D(n413), .Y(n1914) );
  OAI22X1 U1468 ( .A(n2407), .B(n363), .C(n2408), .D(n413), .Y(n1915) );
  OAI22X1 U1469 ( .A(n2408), .B(n363), .C(n2409), .D(n413), .Y(n1916) );
  OAI22X1 U1470 ( .A(n2409), .B(n363), .C(n2410), .D(n413), .Y(n1917) );
  OAI22X1 U1471 ( .A(n2410), .B(n363), .C(n2411), .D(n413), .Y(n1918) );
  OAI22X1 U1472 ( .A(n2411), .B(n363), .C(n2412), .D(n413), .Y(n1919) );
  OAI22X1 U1473 ( .A(n2412), .B(n363), .C(n2413), .D(n413), .Y(n1920) );
  OAI22X1 U1474 ( .A(n2413), .B(n363), .C(n2414), .D(n413), .Y(n1921) );
  OAI22X1 U1475 ( .A(n2414), .B(n363), .C(n2415), .D(n413), .Y(n1922) );
  OAI22X1 U1476 ( .A(n2415), .B(n363), .C(n2416), .D(n413), .Y(n1923) );
  OAI22X1 U1477 ( .A(n2416), .B(n362), .C(n2417), .D(n413), .Y(n1924) );
  OAI22X1 U1478 ( .A(n2417), .B(n362), .C(n2418), .D(n412), .Y(n1925) );
  OAI22X1 U1479 ( .A(n2418), .B(n362), .C(n2419), .D(n412), .Y(n1926) );
  OAI22X1 U1480 ( .A(n2419), .B(n362), .C(n2420), .D(n412), .Y(n1927) );
  OAI22X1 U1481 ( .A(n2420), .B(n362), .C(n2421), .D(n412), .Y(n1928) );
  OAI22X1 U1482 ( .A(n2421), .B(n362), .C(n2422), .D(n412), .Y(n1929) );
  OAI22X1 U1483 ( .A(n2422), .B(n362), .C(n2423), .D(n412), .Y(n1930) );
  OAI22X1 U1484 ( .A(n2423), .B(n362), .C(n2424), .D(n412), .Y(n1931) );
  OAI22X1 U1485 ( .A(n2424), .B(n362), .C(n2425), .D(n412), .Y(n1932) );
  OAI22X1 U1486 ( .A(n2425), .B(n362), .C(n2426), .D(n412), .Y(n1933) );
  OAI22X1 U1487 ( .A(n2426), .B(n362), .C(n2427), .D(n412), .Y(n1934) );
  XNOR2X1 U1488 ( .A(n316), .B(n2948), .Y(n2398) );
  XNOR2X1 U1489 ( .A(n316), .B(n2910), .Y(n2399) );
  XNOR2X1 U1490 ( .A(n316), .B(n2947), .Y(n2400) );
  XNOR2X1 U1491 ( .A(n316), .B(n2949), .Y(n2401) );
  XNOR2X1 U1492 ( .A(n316), .B(n485), .Y(n2402) );
  XNOR2X1 U1493 ( .A(n316), .B(n483), .Y(n2403) );
  XNOR2X1 U1494 ( .A(n316), .B(n2913), .Y(n2404) );
  XNOR2X1 U1495 ( .A(n316), .B(n479), .Y(n2405) );
  XNOR2X1 U1496 ( .A(n316), .B(n477), .Y(n2406) );
  XNOR2X1 U1497 ( .A(n315), .B(n475), .Y(n2407) );
  XNOR2X1 U1498 ( .A(n315), .B(n473), .Y(n2408) );
  XNOR2X1 U1499 ( .A(n315), .B(n471), .Y(n2409) );
  XNOR2X1 U1500 ( .A(n315), .B(n469), .Y(n2410) );
  XNOR2X1 U1501 ( .A(n315), .B(n467), .Y(n2411) );
  XNOR2X1 U1502 ( .A(n315), .B(n465), .Y(n2412) );
  XNOR2X1 U1503 ( .A(n315), .B(n463), .Y(n2413) );
  XNOR2X1 U1504 ( .A(n315), .B(n461), .Y(n2414) );
  XNOR2X1 U1505 ( .A(n315), .B(n459), .Y(n2415) );
  XNOR2X1 U1506 ( .A(n315), .B(n457), .Y(n2416) );
  XNOR2X1 U1507 ( .A(n315), .B(n455), .Y(n2417) );
  XNOR2X1 U1508 ( .A(n315), .B(n453), .Y(n2418) );
  XNOR2X1 U1509 ( .A(n314), .B(n451), .Y(n2419) );
  XNOR2X1 U1510 ( .A(n314), .B(n449), .Y(n2420) );
  XNOR2X1 U1511 ( .A(n314), .B(n447), .Y(n2421) );
  XNOR2X1 U1512 ( .A(n314), .B(n445), .Y(n2422) );
  XNOR2X1 U1513 ( .A(n314), .B(n443), .Y(n2423) );
  XNOR2X1 U1514 ( .A(n314), .B(n441), .Y(n2424) );
  XNOR2X1 U1515 ( .A(n314), .B(n439), .Y(n2425) );
  XNOR2X1 U1516 ( .A(n314), .B(n437), .Y(n2426) );
  XNOR2X1 U1517 ( .A(n314), .B(n2950), .Y(n2427) );
  OAI22X1 U1518 ( .A(n361), .B(n2461), .C(n2803), .D(n411), .Y(n1750) );
  OAI22X1 U1519 ( .A(n2429), .B(n361), .C(n2430), .D(n411), .Y(n1936) );
  OAI22X1 U1520 ( .A(n2430), .B(n361), .C(n2431), .D(n411), .Y(n1937) );
  OAI22X1 U1521 ( .A(n2431), .B(n361), .C(n2432), .D(n411), .Y(n1938) );
  OAI22X1 U1522 ( .A(n2432), .B(n361), .C(n2433), .D(n411), .Y(n1939) );
  OAI22X1 U1523 ( .A(n2433), .B(n361), .C(n2434), .D(n411), .Y(n1940) );
  OAI22X1 U1524 ( .A(n2434), .B(n361), .C(n2435), .D(n411), .Y(n1941) );
  OAI22X1 U1525 ( .A(n2435), .B(n361), .C(n2436), .D(n411), .Y(n1942) );
  OAI22X1 U1526 ( .A(n2436), .B(n361), .C(n2437), .D(n411), .Y(n1943) );
  OAI22X1 U1527 ( .A(n2437), .B(n360), .C(n2438), .D(n411), .Y(n1944) );
  OAI22X1 U1528 ( .A(n2438), .B(n360), .C(n2439), .D(n410), .Y(n1945) );
  OAI22X1 U1529 ( .A(n2439), .B(n360), .C(n2440), .D(n410), .Y(n1946) );
  OAI22X1 U1530 ( .A(n2440), .B(n360), .C(n2441), .D(n410), .Y(n1947) );
  OAI22X1 U1531 ( .A(n2441), .B(n360), .C(n2442), .D(n410), .Y(n1948) );
  OAI22X1 U1532 ( .A(n2442), .B(n360), .C(n2443), .D(n410), .Y(n1949) );
  OAI22X1 U1533 ( .A(n2443), .B(n360), .C(n2444), .D(n410), .Y(n1950) );
  OAI22X1 U1534 ( .A(n2444), .B(n360), .C(n2445), .D(n410), .Y(n1951) );
  OAI22X1 U1535 ( .A(n2445), .B(n360), .C(n2446), .D(n410), .Y(n1952) );
  OAI22X1 U1536 ( .A(n2446), .B(n360), .C(n2447), .D(n410), .Y(n1953) );
  OAI22X1 U1537 ( .A(n2447), .B(n360), .C(n2448), .D(n410), .Y(n1954) );
  OAI22X1 U1538 ( .A(n2448), .B(n360), .C(n2449), .D(n410), .Y(n1955) );
  OAI22X1 U1539 ( .A(n2449), .B(n359), .C(n2450), .D(n410), .Y(n1956) );
  OAI22X1 U1540 ( .A(n2450), .B(n359), .C(n2451), .D(n409), .Y(n1957) );
  OAI22X1 U1541 ( .A(n2451), .B(n359), .C(n2452), .D(n409), .Y(n1958) );
  OAI22X1 U1542 ( .A(n2452), .B(n359), .C(n2453), .D(n409), .Y(n1959) );
  OAI22X1 U1543 ( .A(n2453), .B(n359), .C(n2454), .D(n409), .Y(n1960) );
  OAI22X1 U1544 ( .A(n2454), .B(n359), .C(n2455), .D(n409), .Y(n1961) );
  OAI22X1 U1545 ( .A(n2455), .B(n359), .C(n2456), .D(n409), .Y(n1962) );
  OAI22X1 U1546 ( .A(n2456), .B(n359), .C(n2457), .D(n409), .Y(n1963) );
  OAI22X1 U1547 ( .A(n2457), .B(n359), .C(n2458), .D(n409), .Y(n1964) );
  OAI22X1 U1548 ( .A(n2458), .B(n359), .C(n2459), .D(n409), .Y(n1965) );
  OAI22X1 U1549 ( .A(n2459), .B(n359), .C(n2460), .D(n409), .Y(n1966) );
  XNOR2X1 U1550 ( .A(n313), .B(b[31]), .Y(n2429) );
  XNOR2X1 U1551 ( .A(n313), .B(b[30]), .Y(n2430) );
  XNOR2X1 U1552 ( .A(n313), .B(n2948), .Y(n2431) );
  XNOR2X1 U1553 ( .A(n313), .B(n2910), .Y(n2432) );
  XNOR2X1 U1554 ( .A(n313), .B(n2947), .Y(n2433) );
  XNOR2X1 U1555 ( .A(n313), .B(n2949), .Y(n2434) );
  XNOR2X1 U1556 ( .A(n313), .B(n485), .Y(n2435) );
  XNOR2X1 U1557 ( .A(n313), .B(n483), .Y(n2436) );
  XNOR2X1 U1558 ( .A(n313), .B(n2913), .Y(n2437) );
  XNOR2X1 U1559 ( .A(n313), .B(n479), .Y(n2438) );
  XNOR2X1 U1560 ( .A(n313), .B(n477), .Y(n2439) );
  XNOR2X1 U1561 ( .A(n312), .B(n475), .Y(n2440) );
  XNOR2X1 U1562 ( .A(n312), .B(n473), .Y(n2441) );
  XNOR2X1 U1563 ( .A(n312), .B(n471), .Y(n2442) );
  XNOR2X1 U1564 ( .A(n312), .B(n469), .Y(n2443) );
  XNOR2X1 U1565 ( .A(n312), .B(n467), .Y(n2444) );
  XNOR2X1 U1566 ( .A(n312), .B(n465), .Y(n2445) );
  XNOR2X1 U1567 ( .A(n312), .B(n463), .Y(n2446) );
  XNOR2X1 U1568 ( .A(n312), .B(n461), .Y(n2447) );
  XNOR2X1 U1569 ( .A(n312), .B(n459), .Y(n2448) );
  XNOR2X1 U1570 ( .A(n312), .B(n457), .Y(n2449) );
  XNOR2X1 U1571 ( .A(n312), .B(n455), .Y(n2450) );
  XNOR2X1 U1572 ( .A(n312), .B(n453), .Y(n2451) );
  XNOR2X1 U1573 ( .A(n311), .B(n451), .Y(n2452) );
  XNOR2X1 U1574 ( .A(n311), .B(n449), .Y(n2453) );
  XNOR2X1 U1575 ( .A(n311), .B(n447), .Y(n2454) );
  XNOR2X1 U1576 ( .A(n311), .B(n445), .Y(n2455) );
  XNOR2X1 U1577 ( .A(n311), .B(n443), .Y(n2456) );
  XNOR2X1 U1578 ( .A(n311), .B(n441), .Y(n2457) );
  XNOR2X1 U1579 ( .A(n311), .B(n439), .Y(n2458) );
  XNOR2X1 U1580 ( .A(n311), .B(n437), .Y(n2459) );
  XNOR2X1 U1581 ( .A(n311), .B(n2950), .Y(n2460) );
  OAI22X1 U1582 ( .A(n358), .B(n2494), .C(n2804), .D(n408), .Y(n1751) );
  OAI22X1 U1583 ( .A(n2804), .B(n358), .C(n2462), .D(n408), .Y(n1969) );
  OAI22X1 U1584 ( .A(n2462), .B(n358), .C(n2463), .D(n408), .Y(n1970) );
  OAI22X1 U1585 ( .A(n2463), .B(n358), .C(n2464), .D(n408), .Y(n1971) );
  OAI22X1 U1586 ( .A(n2464), .B(n358), .C(n2465), .D(n408), .Y(n1972) );
  OAI22X1 U1587 ( .A(n2465), .B(n358), .C(n2466), .D(n408), .Y(n1973) );
  OAI22X1 U1588 ( .A(n2466), .B(n358), .C(n2467), .D(n408), .Y(n1974) );
  OAI22X1 U1589 ( .A(n2467), .B(n358), .C(n2468), .D(n408), .Y(n1975) );
  OAI22X1 U1590 ( .A(n2468), .B(n358), .C(n2469), .D(n408), .Y(n1976) );
  OAI22X1 U1591 ( .A(n2469), .B(n358), .C(n2470), .D(n408), .Y(n1977) );
  OAI22X1 U1592 ( .A(n2470), .B(n357), .C(n2471), .D(n408), .Y(n1978) );
  OAI22X1 U1593 ( .A(n2471), .B(n357), .C(n2472), .D(n407), .Y(n1979) );
  OAI22X1 U1594 ( .A(n2472), .B(n357), .C(n2473), .D(n407), .Y(n1980) );
  OAI22X1 U1595 ( .A(n2473), .B(n357), .C(n2474), .D(n407), .Y(n1981) );
  OAI22X1 U1596 ( .A(n2474), .B(n357), .C(n2475), .D(n407), .Y(n1982) );
  OAI22X1 U1597 ( .A(n2475), .B(n357), .C(n2476), .D(n407), .Y(n1983) );
  OAI22X1 U1598 ( .A(n2476), .B(n357), .C(n2477), .D(n407), .Y(n1984) );
  OAI22X1 U1599 ( .A(n2477), .B(n357), .C(n2478), .D(n407), .Y(n1985) );
  OAI22X1 U1600 ( .A(n2478), .B(n357), .C(n2479), .D(n407), .Y(n1986) );
  OAI22X1 U1601 ( .A(n2479), .B(n357), .C(n2480), .D(n407), .Y(n1987) );
  OAI22X1 U1602 ( .A(n2480), .B(n357), .C(n2481), .D(n407), .Y(n1988) );
  OAI22X1 U1603 ( .A(n2481), .B(n357), .C(n2482), .D(n407), .Y(n1989) );
  OAI22X1 U1604 ( .A(n2482), .B(n356), .C(n2483), .D(n407), .Y(n1990) );
  OAI22X1 U1605 ( .A(n2483), .B(n356), .C(n2484), .D(n406), .Y(n1991) );
  OAI22X1 U1606 ( .A(n2484), .B(n356), .C(n2485), .D(n406), .Y(n1992) );
  OAI22X1 U1607 ( .A(n2485), .B(n356), .C(n2486), .D(n406), .Y(n1993) );
  OAI22X1 U1608 ( .A(n2486), .B(n356), .C(n2487), .D(n406), .Y(n1994) );
  OAI22X1 U1609 ( .A(n2487), .B(n356), .C(n2488), .D(n406), .Y(n1995) );
  OAI22X1 U1610 ( .A(n2488), .B(n356), .C(n2489), .D(n406), .Y(n1996) );
  OAI22X1 U1611 ( .A(n2489), .B(n356), .C(n2490), .D(n406), .Y(n1997) );
  OAI22X1 U1612 ( .A(n2490), .B(n356), .C(n2491), .D(n406), .Y(n1998) );
  OAI22X1 U1613 ( .A(n2491), .B(n356), .C(n2492), .D(n406), .Y(n1999) );
  OAI22X1 U1614 ( .A(n2492), .B(n356), .C(n2493), .D(n406), .Y(n2000) );
  XNOR2X1 U1615 ( .A(n310), .B(n497), .Y(n2462) );
  XNOR2X1 U1616 ( .A(n310), .B(n495), .Y(n2463) );
  XNOR2X1 U1617 ( .A(n310), .B(n2918), .Y(n2464) );
  XNOR2X1 U1618 ( .A(n310), .B(n491), .Y(n2465) );
  XNOR2X1 U1619 ( .A(n310), .B(n489), .Y(n2466) );
  XNOR2X1 U1620 ( .A(n310), .B(n2949), .Y(n2467) );
  XNOR2X1 U1621 ( .A(n310), .B(n485), .Y(n2468) );
  XNOR2X1 U1622 ( .A(n310), .B(n483), .Y(n2469) );
  XNOR2X1 U1623 ( .A(n310), .B(n2913), .Y(n2470) );
  XNOR2X1 U1624 ( .A(n310), .B(n479), .Y(n2471) );
  XNOR2X1 U1625 ( .A(n310), .B(n477), .Y(n2472) );
  XNOR2X1 U1626 ( .A(n309), .B(n475), .Y(n2473) );
  XNOR2X1 U1627 ( .A(n309), .B(n473), .Y(n2474) );
  XNOR2X1 U1628 ( .A(n309), .B(n471), .Y(n2475) );
  XNOR2X1 U1629 ( .A(n309), .B(n469), .Y(n2476) );
  XNOR2X1 U1630 ( .A(n309), .B(n467), .Y(n2477) );
  XNOR2X1 U1631 ( .A(n309), .B(n465), .Y(n2478) );
  XNOR2X1 U1632 ( .A(n309), .B(n463), .Y(n2479) );
  XNOR2X1 U1633 ( .A(n309), .B(n461), .Y(n2480) );
  XNOR2X1 U1634 ( .A(n309), .B(n459), .Y(n2481) );
  XNOR2X1 U1635 ( .A(n309), .B(n457), .Y(n2482) );
  XNOR2X1 U1636 ( .A(n309), .B(n455), .Y(n2483) );
  XNOR2X1 U1637 ( .A(n309), .B(n453), .Y(n2484) );
  XNOR2X1 U1638 ( .A(n308), .B(n451), .Y(n2485) );
  XNOR2X1 U1639 ( .A(n308), .B(n449), .Y(n2486) );
  XNOR2X1 U1640 ( .A(n308), .B(n447), .Y(n2487) );
  XNOR2X1 U1641 ( .A(n308), .B(n445), .Y(n2488) );
  XNOR2X1 U1642 ( .A(n308), .B(n443), .Y(n2489) );
  XNOR2X1 U1643 ( .A(n308), .B(n441), .Y(n2490) );
  XNOR2X1 U1644 ( .A(n308), .B(n439), .Y(n2491) );
  XNOR2X1 U1645 ( .A(n308), .B(n437), .Y(n2492) );
  XNOR2X1 U1646 ( .A(n308), .B(n2950), .Y(n2493) );
  OAI22X1 U1647 ( .A(n355), .B(n2527), .C(n2805), .D(n405), .Y(n1752) );
  OAI22X1 U1648 ( .A(n2805), .B(n355), .C(n2495), .D(n405), .Y(n2003) );
  OAI22X1 U1649 ( .A(n2495), .B(n355), .C(n2496), .D(n405), .Y(n2004) );
  OAI22X1 U1650 ( .A(n2496), .B(n355), .C(n2497), .D(n405), .Y(n2005) );
  OAI22X1 U1651 ( .A(n2497), .B(n355), .C(n2498), .D(n405), .Y(n2006) );
  OAI22X1 U1652 ( .A(n2498), .B(n355), .C(n2499), .D(n405), .Y(n2007) );
  OAI22X1 U1653 ( .A(n2499), .B(n355), .C(n2500), .D(n405), .Y(n2008) );
  OAI22X1 U1654 ( .A(n2500), .B(n355), .C(n2501), .D(n405), .Y(n2009) );
  OAI22X1 U1655 ( .A(n2501), .B(n355), .C(n2502), .D(n405), .Y(n2010) );
  OAI22X1 U1656 ( .A(n2502), .B(n355), .C(n2503), .D(n405), .Y(n2011) );
  OAI22X1 U1657 ( .A(n2503), .B(n354), .C(n2504), .D(n405), .Y(n2012) );
  OAI22X1 U1658 ( .A(n2504), .B(n354), .C(n2505), .D(n404), .Y(n2013) );
  OAI22X1 U1659 ( .A(n2505), .B(n354), .C(n2506), .D(n404), .Y(n2014) );
  OAI22X1 U1660 ( .A(n2506), .B(n354), .C(n2507), .D(n404), .Y(n2015) );
  OAI22X1 U1661 ( .A(n2507), .B(n354), .C(n2508), .D(n404), .Y(n2016) );
  OAI22X1 U1662 ( .A(n2508), .B(n354), .C(n2509), .D(n404), .Y(n2017) );
  OAI22X1 U1663 ( .A(n2509), .B(n354), .C(n2510), .D(n404), .Y(n2018) );
  OAI22X1 U1664 ( .A(n2510), .B(n354), .C(n2511), .D(n404), .Y(n2019) );
  OAI22X1 U1665 ( .A(n2511), .B(n354), .C(n2512), .D(n404), .Y(n2020) );
  OAI22X1 U1666 ( .A(n2512), .B(n354), .C(n2513), .D(n404), .Y(n2021) );
  OAI22X1 U1667 ( .A(n2513), .B(n354), .C(n2514), .D(n404), .Y(n2022) );
  OAI22X1 U1668 ( .A(n2514), .B(n354), .C(n2515), .D(n404), .Y(n2023) );
  OAI22X1 U1669 ( .A(n2515), .B(n353), .C(n2516), .D(n404), .Y(n2024) );
  OAI22X1 U1670 ( .A(n2516), .B(n353), .C(n2517), .D(n403), .Y(n2025) );
  OAI22X1 U1671 ( .A(n2517), .B(n353), .C(n2518), .D(n403), .Y(n2026) );
  OAI22X1 U1672 ( .A(n2518), .B(n353), .C(n2519), .D(n403), .Y(n2027) );
  OAI22X1 U1673 ( .A(n2519), .B(n353), .C(n2520), .D(n403), .Y(n2028) );
  OAI22X1 U1674 ( .A(n2520), .B(n353), .C(n2521), .D(n403), .Y(n2029) );
  OAI22X1 U1675 ( .A(n2521), .B(n353), .C(n2522), .D(n403), .Y(n2030) );
  OAI22X1 U1676 ( .A(n2522), .B(n353), .C(n2523), .D(n403), .Y(n2031) );
  OAI22X1 U1677 ( .A(n2523), .B(n353), .C(n2524), .D(n403), .Y(n2032) );
  OAI22X1 U1678 ( .A(n2524), .B(n353), .C(n2525), .D(n403), .Y(n2033) );
  OAI22X1 U1679 ( .A(n2525), .B(n353), .C(n2526), .D(n403), .Y(n2034) );
  XNOR2X1 U1680 ( .A(n307), .B(n497), .Y(n2495) );
  XNOR2X1 U1681 ( .A(n307), .B(n495), .Y(n2496) );
  XNOR2X1 U1682 ( .A(n307), .B(n2917), .Y(n2497) );
  XNOR2X1 U1683 ( .A(n307), .B(n491), .Y(n2498) );
  XNOR2X1 U1684 ( .A(n307), .B(n489), .Y(n2499) );
  XNOR2X1 U1685 ( .A(n307), .B(n2949), .Y(n2500) );
  XNOR2X1 U1686 ( .A(n307), .B(n485), .Y(n2501) );
  XNOR2X1 U1687 ( .A(n307), .B(n483), .Y(n2502) );
  XNOR2X1 U1688 ( .A(n307), .B(n2913), .Y(n2503) );
  XNOR2X1 U1689 ( .A(n307), .B(n479), .Y(n2504) );
  XNOR2X1 U1690 ( .A(n307), .B(n477), .Y(n2505) );
  XNOR2X1 U1691 ( .A(n306), .B(n475), .Y(n2506) );
  XNOR2X1 U1692 ( .A(n306), .B(n473), .Y(n2507) );
  XNOR2X1 U1693 ( .A(n306), .B(n471), .Y(n2508) );
  XNOR2X1 U1694 ( .A(n306), .B(n469), .Y(n2509) );
  XNOR2X1 U1695 ( .A(n306), .B(n467), .Y(n2510) );
  XNOR2X1 U1696 ( .A(n306), .B(n465), .Y(n2511) );
  XNOR2X1 U1697 ( .A(n306), .B(n463), .Y(n2512) );
  XNOR2X1 U1698 ( .A(n306), .B(n461), .Y(n2513) );
  XNOR2X1 U1699 ( .A(n306), .B(n459), .Y(n2514) );
  XNOR2X1 U1700 ( .A(n306), .B(n457), .Y(n2515) );
  XNOR2X1 U1701 ( .A(n306), .B(n455), .Y(n2516) );
  XNOR2X1 U1702 ( .A(n306), .B(n453), .Y(n2517) );
  XNOR2X1 U1703 ( .A(n305), .B(n451), .Y(n2518) );
  XNOR2X1 U1704 ( .A(n305), .B(n449), .Y(n2519) );
  XNOR2X1 U1705 ( .A(n305), .B(n447), .Y(n2520) );
  XNOR2X1 U1706 ( .A(n305), .B(n445), .Y(n2521) );
  XNOR2X1 U1707 ( .A(n305), .B(n443), .Y(n2522) );
  XNOR2X1 U1708 ( .A(n305), .B(n441), .Y(n2523) );
  XNOR2X1 U1709 ( .A(n305), .B(n439), .Y(n2524) );
  XNOR2X1 U1710 ( .A(n305), .B(n437), .Y(n2525) );
  XNOR2X1 U1711 ( .A(n305), .B(n2950), .Y(n2526) );
  OAI22X1 U1712 ( .A(n352), .B(n2560), .C(n2806), .D(n402), .Y(n1753) );
  OAI22X1 U1713 ( .A(n2806), .B(n352), .C(n2528), .D(n402), .Y(n2037) );
  OAI22X1 U1714 ( .A(n2528), .B(n352), .C(n2529), .D(n402), .Y(n2038) );
  OAI22X1 U1715 ( .A(n2529), .B(n352), .C(n2530), .D(n402), .Y(n2039) );
  OAI22X1 U1716 ( .A(n2530), .B(n352), .C(n2531), .D(n402), .Y(n2040) );
  OAI22X1 U1717 ( .A(n2531), .B(n352), .C(n2532), .D(n402), .Y(n2041) );
  OAI22X1 U1718 ( .A(n2532), .B(n352), .C(n2533), .D(n402), .Y(n2042) );
  OAI22X1 U1719 ( .A(n2533), .B(n352), .C(n2534), .D(n402), .Y(n2043) );
  OAI22X1 U1720 ( .A(n2534), .B(n352), .C(n2535), .D(n402), .Y(n2044) );
  OAI22X1 U1721 ( .A(n2535), .B(n352), .C(n2536), .D(n402), .Y(n2045) );
  OAI22X1 U1722 ( .A(n2536), .B(n351), .C(n2537), .D(n402), .Y(n2046) );
  OAI22X1 U1723 ( .A(n2537), .B(n351), .C(n2538), .D(n401), .Y(n2047) );
  OAI22X1 U1724 ( .A(n2538), .B(n351), .C(n2539), .D(n401), .Y(n2048) );
  OAI22X1 U1725 ( .A(n2539), .B(n351), .C(n2540), .D(n401), .Y(n2049) );
  OAI22X1 U1726 ( .A(n2540), .B(n351), .C(n2541), .D(n401), .Y(n2050) );
  OAI22X1 U1727 ( .A(n2541), .B(n351), .C(n2542), .D(n401), .Y(n2051) );
  OAI22X1 U1728 ( .A(n2542), .B(n351), .C(n2543), .D(n401), .Y(n2052) );
  OAI22X1 U1729 ( .A(n2543), .B(n351), .C(n2544), .D(n401), .Y(n2053) );
  OAI22X1 U1730 ( .A(n2544), .B(n351), .C(n2545), .D(n401), .Y(n2054) );
  OAI22X1 U1731 ( .A(n2545), .B(n351), .C(n2546), .D(n401), .Y(n2055) );
  OAI22X1 U1732 ( .A(n2546), .B(n351), .C(n2547), .D(n401), .Y(n2056) );
  OAI22X1 U1733 ( .A(n2547), .B(n351), .C(n2548), .D(n401), .Y(n2057) );
  OAI22X1 U1734 ( .A(n2548), .B(n350), .C(n2549), .D(n401), .Y(n2058) );
  OAI22X1 U1735 ( .A(n2549), .B(n350), .C(n2550), .D(n400), .Y(n2059) );
  OAI22X1 U1736 ( .A(n2550), .B(n350), .C(n2551), .D(n400), .Y(n2060) );
  OAI22X1 U1737 ( .A(n2551), .B(n350), .C(n2552), .D(n400), .Y(n2061) );
  OAI22X1 U1738 ( .A(n2552), .B(n350), .C(n2553), .D(n400), .Y(n2062) );
  OAI22X1 U1739 ( .A(n2553), .B(n350), .C(n2554), .D(n400), .Y(n2063) );
  OAI22X1 U1740 ( .A(n2554), .B(n350), .C(n2555), .D(n400), .Y(n2064) );
  OAI22X1 U1741 ( .A(n2555), .B(n350), .C(n2556), .D(n400), .Y(n2065) );
  OAI22X1 U1742 ( .A(n2556), .B(n350), .C(n2557), .D(n400), .Y(n2066) );
  OAI22X1 U1743 ( .A(n2557), .B(n350), .C(n2558), .D(n400), .Y(n2067) );
  OAI22X1 U1744 ( .A(n2558), .B(n350), .C(n2559), .D(n400), .Y(n2068) );
  XNOR2X1 U1745 ( .A(n304), .B(n497), .Y(n2528) );
  XNOR2X1 U1746 ( .A(n304), .B(n495), .Y(n2529) );
  XNOR2X1 U1747 ( .A(n304), .B(n2917), .Y(n2530) );
  XNOR2X1 U1748 ( .A(n304), .B(n491), .Y(n2531) );
  XNOR2X1 U1749 ( .A(n304), .B(n2947), .Y(n2532) );
  XNOR2X1 U1750 ( .A(n304), .B(n2949), .Y(n2533) );
  XNOR2X1 U1751 ( .A(n304), .B(n485), .Y(n2534) );
  XNOR2X1 U1752 ( .A(n304), .B(n483), .Y(n2535) );
  XNOR2X1 U1753 ( .A(n304), .B(n2913), .Y(n2536) );
  XNOR2X1 U1754 ( .A(n304), .B(n479), .Y(n2537) );
  XNOR2X1 U1755 ( .A(n304), .B(n477), .Y(n2538) );
  XNOR2X1 U1756 ( .A(n303), .B(n475), .Y(n2539) );
  XNOR2X1 U1757 ( .A(n303), .B(n473), .Y(n2540) );
  XNOR2X1 U1758 ( .A(n303), .B(n471), .Y(n2541) );
  XNOR2X1 U1759 ( .A(n303), .B(n469), .Y(n2542) );
  XNOR2X1 U1760 ( .A(n303), .B(n467), .Y(n2543) );
  XNOR2X1 U1761 ( .A(n303), .B(n465), .Y(n2544) );
  XNOR2X1 U1762 ( .A(n303), .B(n463), .Y(n2545) );
  XNOR2X1 U1763 ( .A(n303), .B(n461), .Y(n2546) );
  XNOR2X1 U1764 ( .A(n303), .B(n459), .Y(n2547) );
  XNOR2X1 U1765 ( .A(n303), .B(n457), .Y(n2548) );
  XNOR2X1 U1766 ( .A(n303), .B(n455), .Y(n2549) );
  XNOR2X1 U1767 ( .A(n303), .B(n453), .Y(n2550) );
  XNOR2X1 U1768 ( .A(n302), .B(n451), .Y(n2551) );
  XNOR2X1 U1769 ( .A(n302), .B(n449), .Y(n2552) );
  XNOR2X1 U1770 ( .A(n302), .B(n447), .Y(n2553) );
  XNOR2X1 U1771 ( .A(n302), .B(n445), .Y(n2554) );
  XNOR2X1 U1772 ( .A(n302), .B(n443), .Y(n2555) );
  XNOR2X1 U1773 ( .A(n302), .B(n441), .Y(n2556) );
  XNOR2X1 U1774 ( .A(n302), .B(n439), .Y(n2557) );
  XNOR2X1 U1775 ( .A(n302), .B(n437), .Y(n2558) );
  XNOR2X1 U1776 ( .A(n302), .B(n2950), .Y(n2559) );
  OAI22X1 U1777 ( .A(n349), .B(n2593), .C(n2807), .D(n399), .Y(n1754) );
  OAI22X1 U1778 ( .A(n2807), .B(n349), .C(n2561), .D(n399), .Y(n2071) );
  OAI22X1 U1779 ( .A(n2561), .B(n349), .C(n2562), .D(n399), .Y(n2072) );
  OAI22X1 U1780 ( .A(n2562), .B(n349), .C(n2563), .D(n399), .Y(n2073) );
  OAI22X1 U1781 ( .A(n2563), .B(n349), .C(n2564), .D(n399), .Y(n2074) );
  OAI22X1 U1782 ( .A(n2564), .B(n349), .C(n2565), .D(n399), .Y(n2075) );
  OAI22X1 U1783 ( .A(n2565), .B(n349), .C(n2566), .D(n399), .Y(n2076) );
  OAI22X1 U1784 ( .A(n2566), .B(n349), .C(n2567), .D(n399), .Y(n2077) );
  OAI22X1 U1785 ( .A(n2567), .B(n349), .C(n2568), .D(n399), .Y(n2078) );
  OAI22X1 U1786 ( .A(n2568), .B(n349), .C(n2569), .D(n399), .Y(n2079) );
  OAI22X1 U1787 ( .A(n2569), .B(n348), .C(n2570), .D(n399), .Y(n2080) );
  OAI22X1 U1788 ( .A(n2570), .B(n348), .C(n2571), .D(n398), .Y(n2081) );
  OAI22X1 U1789 ( .A(n2571), .B(n348), .C(n2572), .D(n398), .Y(n2082) );
  OAI22X1 U1790 ( .A(n2572), .B(n348), .C(n2573), .D(n398), .Y(n2083) );
  OAI22X1 U1791 ( .A(n2573), .B(n348), .C(n2574), .D(n398), .Y(n2084) );
  OAI22X1 U1792 ( .A(n2574), .B(n348), .C(n2575), .D(n398), .Y(n2085) );
  OAI22X1 U1793 ( .A(n2575), .B(n348), .C(n2576), .D(n398), .Y(n2086) );
  OAI22X1 U1794 ( .A(n2576), .B(n348), .C(n2577), .D(n398), .Y(n2087) );
  OAI22X1 U1795 ( .A(n2577), .B(n348), .C(n2578), .D(n398), .Y(n2088) );
  OAI22X1 U1796 ( .A(n2578), .B(n348), .C(n2579), .D(n398), .Y(n2089) );
  OAI22X1 U1797 ( .A(n2579), .B(n348), .C(n2580), .D(n398), .Y(n2090) );
  OAI22X1 U1798 ( .A(n2580), .B(n348), .C(n2581), .D(n398), .Y(n2091) );
  OAI22X1 U1799 ( .A(n2581), .B(n347), .C(n2582), .D(n398), .Y(n2092) );
  OAI22X1 U1800 ( .A(n2582), .B(n347), .C(n2583), .D(n397), .Y(n2093) );
  OAI22X1 U1801 ( .A(n2583), .B(n347), .C(n2584), .D(n397), .Y(n2094) );
  OAI22X1 U1802 ( .A(n2584), .B(n347), .C(n2585), .D(n397), .Y(n2095) );
  OAI22X1 U1803 ( .A(n2585), .B(n347), .C(n2586), .D(n397), .Y(n2096) );
  OAI22X1 U1804 ( .A(n2586), .B(n347), .C(n2587), .D(n397), .Y(n2097) );
  OAI22X1 U1805 ( .A(n2587), .B(n347), .C(n2588), .D(n397), .Y(n2098) );
  OAI22X1 U1806 ( .A(n2588), .B(n347), .C(n2589), .D(n397), .Y(n2099) );
  OAI22X1 U1807 ( .A(n2589), .B(n347), .C(n2590), .D(n397), .Y(n2100) );
  OAI22X1 U1808 ( .A(n2590), .B(n347), .C(n2591), .D(n397), .Y(n2101) );
  OAI22X1 U1809 ( .A(n2591), .B(n347), .C(n2592), .D(n397), .Y(n2102) );
  XNOR2X1 U1810 ( .A(n301), .B(n497), .Y(n2561) );
  XNOR2X1 U1811 ( .A(n301), .B(n495), .Y(n2562) );
  XNOR2X1 U1812 ( .A(n301), .B(n2918), .Y(n2563) );
  XNOR2X1 U1813 ( .A(n301), .B(n491), .Y(n2564) );
  XNOR2X1 U1814 ( .A(n301), .B(n2947), .Y(n2565) );
  XNOR2X1 U1815 ( .A(n301), .B(n2914), .Y(n2566) );
  XNOR2X1 U1816 ( .A(n301), .B(n485), .Y(n2567) );
  XNOR2X1 U1817 ( .A(n301), .B(n483), .Y(n2568) );
  XNOR2X1 U1818 ( .A(n301), .B(n2913), .Y(n2569) );
  XNOR2X1 U1819 ( .A(n301), .B(n479), .Y(n2570) );
  XNOR2X1 U1820 ( .A(n301), .B(n477), .Y(n2571) );
  XNOR2X1 U1821 ( .A(n300), .B(n475), .Y(n2572) );
  XNOR2X1 U1822 ( .A(n300), .B(n473), .Y(n2573) );
  XNOR2X1 U1823 ( .A(n300), .B(n471), .Y(n2574) );
  XNOR2X1 U1824 ( .A(n300), .B(n469), .Y(n2575) );
  XNOR2X1 U1825 ( .A(n300), .B(n467), .Y(n2576) );
  XNOR2X1 U1826 ( .A(n300), .B(n465), .Y(n2577) );
  XNOR2X1 U1827 ( .A(n300), .B(n463), .Y(n2578) );
  XNOR2X1 U1828 ( .A(n300), .B(n461), .Y(n2579) );
  XNOR2X1 U1829 ( .A(n300), .B(n459), .Y(n2580) );
  XNOR2X1 U1830 ( .A(n300), .B(n457), .Y(n2581) );
  XNOR2X1 U1831 ( .A(n300), .B(n455), .Y(n2582) );
  XNOR2X1 U1832 ( .A(n300), .B(n453), .Y(n2583) );
  XNOR2X1 U1833 ( .A(n299), .B(n451), .Y(n2584) );
  XNOR2X1 U1834 ( .A(n299), .B(n449), .Y(n2585) );
  XNOR2X1 U1835 ( .A(n299), .B(n447), .Y(n2586) );
  XNOR2X1 U1836 ( .A(n299), .B(n445), .Y(n2587) );
  XNOR2X1 U1837 ( .A(n299), .B(n443), .Y(n2588) );
  XNOR2X1 U1838 ( .A(n299), .B(n441), .Y(n2589) );
  XNOR2X1 U1839 ( .A(n299), .B(n439), .Y(n2590) );
  XNOR2X1 U1840 ( .A(n299), .B(n437), .Y(n2591) );
  XNOR2X1 U1841 ( .A(n299), .B(n2950), .Y(n2592) );
  OAI22X1 U1842 ( .A(n346), .B(n2626), .C(n2808), .D(n396), .Y(n1755) );
  OAI22X1 U1843 ( .A(n2808), .B(n346), .C(n2594), .D(n396), .Y(n2105) );
  OAI22X1 U1844 ( .A(n2594), .B(n346), .C(n2595), .D(n396), .Y(n2106) );
  OAI22X1 U1845 ( .A(n2595), .B(n346), .C(n2596), .D(n396), .Y(n2107) );
  OAI22X1 U1846 ( .A(n2596), .B(n346), .C(n2597), .D(n396), .Y(n2108) );
  OAI22X1 U1847 ( .A(n2597), .B(n346), .C(n2598), .D(n396), .Y(n2109) );
  OAI22X1 U1848 ( .A(n2598), .B(n346), .C(n2599), .D(n396), .Y(n2110) );
  OAI22X1 U1849 ( .A(n2599), .B(n346), .C(n2600), .D(n396), .Y(n2111) );
  OAI22X1 U1850 ( .A(n2600), .B(n346), .C(n2601), .D(n396), .Y(n2112) );
  OAI22X1 U1851 ( .A(n2601), .B(n346), .C(n2602), .D(n396), .Y(n2113) );
  OAI22X1 U1852 ( .A(n2602), .B(n345), .C(n2603), .D(n396), .Y(n2114) );
  OAI22X1 U1853 ( .A(n2603), .B(n345), .C(n2604), .D(n395), .Y(n2115) );
  OAI22X1 U1854 ( .A(n2604), .B(n345), .C(n2605), .D(n395), .Y(n2116) );
  OAI22X1 U1855 ( .A(n2605), .B(n345), .C(n2606), .D(n395), .Y(n2117) );
  OAI22X1 U1856 ( .A(n2606), .B(n345), .C(n2607), .D(n395), .Y(n2118) );
  OAI22X1 U1857 ( .A(n2607), .B(n345), .C(n2608), .D(n395), .Y(n2119) );
  OAI22X1 U1858 ( .A(n2608), .B(n345), .C(n2609), .D(n395), .Y(n2120) );
  OAI22X1 U1859 ( .A(n2609), .B(n345), .C(n2610), .D(n395), .Y(n2121) );
  OAI22X1 U1860 ( .A(n2610), .B(n345), .C(n2611), .D(n395), .Y(n2122) );
  OAI22X1 U1861 ( .A(n2611), .B(n345), .C(n2612), .D(n395), .Y(n2123) );
  OAI22X1 U1862 ( .A(n2612), .B(n345), .C(n2613), .D(n395), .Y(n2124) );
  OAI22X1 U1863 ( .A(n2613), .B(n345), .C(n2614), .D(n395), .Y(n2125) );
  OAI22X1 U1864 ( .A(n2614), .B(n344), .C(n2615), .D(n395), .Y(n2126) );
  OAI22X1 U1865 ( .A(n2615), .B(n344), .C(n2616), .D(n394), .Y(n2127) );
  OAI22X1 U1866 ( .A(n2616), .B(n344), .C(n2617), .D(n394), .Y(n2128) );
  OAI22X1 U1867 ( .A(n2617), .B(n344), .C(n2618), .D(n394), .Y(n2129) );
  OAI22X1 U1868 ( .A(n2618), .B(n344), .C(n2619), .D(n394), .Y(n2130) );
  OAI22X1 U1869 ( .A(n2619), .B(n344), .C(n2620), .D(n394), .Y(n2131) );
  OAI22X1 U1870 ( .A(n2620), .B(n344), .C(n2621), .D(n394), .Y(n2132) );
  OAI22X1 U1871 ( .A(n2621), .B(n344), .C(n2622), .D(n394), .Y(n2133) );
  OAI22X1 U1872 ( .A(n2622), .B(n344), .C(n2623), .D(n394), .Y(n2134) );
  OAI22X1 U1873 ( .A(n2623), .B(n344), .C(n2624), .D(n394), .Y(n2135) );
  OAI22X1 U1874 ( .A(n2624), .B(n344), .C(n2625), .D(n394), .Y(n2136) );
  XNOR2X1 U1875 ( .A(n298), .B(n497), .Y(n2594) );
  XNOR2X1 U1876 ( .A(n298), .B(n495), .Y(n2595) );
  XNOR2X1 U1877 ( .A(n298), .B(n2917), .Y(n2596) );
  XNOR2X1 U1878 ( .A(n298), .B(n491), .Y(n2597) );
  XNOR2X1 U1879 ( .A(n298), .B(n2947), .Y(n2598) );
  XNOR2X1 U1880 ( .A(n298), .B(n2914), .Y(n2599) );
  XNOR2X1 U1881 ( .A(n298), .B(n485), .Y(n2600) );
  XNOR2X1 U1882 ( .A(n298), .B(n483), .Y(n2601) );
  XNOR2X1 U1883 ( .A(n298), .B(n2913), .Y(n2602) );
  XNOR2X1 U1884 ( .A(n298), .B(n479), .Y(n2603) );
  XNOR2X1 U1885 ( .A(n298), .B(n477), .Y(n2604) );
  XNOR2X1 U1886 ( .A(n297), .B(n475), .Y(n2605) );
  XNOR2X1 U1887 ( .A(n297), .B(n473), .Y(n2606) );
  XNOR2X1 U1888 ( .A(n297), .B(n471), .Y(n2607) );
  XNOR2X1 U1889 ( .A(n297), .B(n469), .Y(n2608) );
  XNOR2X1 U1890 ( .A(n297), .B(n467), .Y(n2609) );
  XNOR2X1 U1891 ( .A(n297), .B(n465), .Y(n2610) );
  XNOR2X1 U1892 ( .A(n297), .B(n463), .Y(n2611) );
  XNOR2X1 U1893 ( .A(n297), .B(n461), .Y(n2612) );
  XNOR2X1 U1894 ( .A(n297), .B(n459), .Y(n2613) );
  XNOR2X1 U1895 ( .A(n297), .B(n457), .Y(n2614) );
  XNOR2X1 U1896 ( .A(n297), .B(n455), .Y(n2615) );
  XNOR2X1 U1897 ( .A(n297), .B(n453), .Y(n2616) );
  XNOR2X1 U1898 ( .A(n296), .B(n451), .Y(n2617) );
  XNOR2X1 U1899 ( .A(n296), .B(n449), .Y(n2618) );
  XNOR2X1 U1900 ( .A(n296), .B(n447), .Y(n2619) );
  XNOR2X1 U1901 ( .A(n296), .B(n445), .Y(n2620) );
  XNOR2X1 U1902 ( .A(n296), .B(n443), .Y(n2621) );
  XNOR2X1 U1903 ( .A(n296), .B(n441), .Y(n2622) );
  XNOR2X1 U1904 ( .A(n296), .B(n439), .Y(n2623) );
  XNOR2X1 U1905 ( .A(n296), .B(n437), .Y(n2624) );
  XNOR2X1 U1906 ( .A(n296), .B(n2950), .Y(n2625) );
  OAI22X1 U1907 ( .A(n343), .B(n2659), .C(n2809), .D(n393), .Y(n1756) );
  OAI22X1 U1908 ( .A(n2809), .B(n343), .C(n2627), .D(n393), .Y(n2139) );
  OAI22X1 U1909 ( .A(n2627), .B(n343), .C(n2628), .D(n393), .Y(n2140) );
  OAI22X1 U1910 ( .A(n2628), .B(n343), .C(n2629), .D(n393), .Y(n2141) );
  OAI22X1 U1911 ( .A(n2629), .B(n343), .C(n2630), .D(n393), .Y(n2142) );
  OAI22X1 U1912 ( .A(n2630), .B(n343), .C(n2631), .D(n393), .Y(n2143) );
  OAI22X1 U1913 ( .A(n2631), .B(n343), .C(n2632), .D(n393), .Y(n2144) );
  OAI22X1 U1914 ( .A(n2632), .B(n343), .C(n2633), .D(n393), .Y(n2145) );
  OAI22X1 U1915 ( .A(n2633), .B(n343), .C(n2634), .D(n393), .Y(n2146) );
  OAI22X1 U1916 ( .A(n2634), .B(n343), .C(n2635), .D(n393), .Y(n2147) );
  OAI22X1 U1917 ( .A(n2635), .B(n342), .C(n2636), .D(n393), .Y(n2148) );
  OAI22X1 U1918 ( .A(n2636), .B(n342), .C(n2637), .D(n392), .Y(n2149) );
  OAI22X1 U1919 ( .A(n2637), .B(n342), .C(n2638), .D(n392), .Y(n2150) );
  OAI22X1 U1920 ( .A(n2638), .B(n342), .C(n2639), .D(n392), .Y(n2151) );
  OAI22X1 U1921 ( .A(n2639), .B(n342), .C(n2640), .D(n392), .Y(n2152) );
  OAI22X1 U1922 ( .A(n2640), .B(n342), .C(n2641), .D(n392), .Y(n2153) );
  OAI22X1 U1923 ( .A(n2641), .B(n342), .C(n2642), .D(n392), .Y(n2154) );
  OAI22X1 U1924 ( .A(n2642), .B(n342), .C(n2643), .D(n392), .Y(n2155) );
  OAI22X1 U1925 ( .A(n2643), .B(n342), .C(n2644), .D(n392), .Y(n2156) );
  OAI22X1 U1926 ( .A(n2644), .B(n342), .C(n2645), .D(n392), .Y(n2157) );
  OAI22X1 U1927 ( .A(n2645), .B(n342), .C(n2646), .D(n392), .Y(n2158) );
  OAI22X1 U1928 ( .A(n2646), .B(n342), .C(n2647), .D(n392), .Y(n2159) );
  OAI22X1 U1929 ( .A(n2647), .B(n341), .C(n2648), .D(n392), .Y(n2160) );
  OAI22X1 U1930 ( .A(n2648), .B(n341), .C(n2649), .D(n391), .Y(n2161) );
  OAI22X1 U1931 ( .A(n2649), .B(n341), .C(n2650), .D(n391), .Y(n2162) );
  OAI22X1 U1932 ( .A(n2650), .B(n341), .C(n2651), .D(n391), .Y(n2163) );
  OAI22X1 U1933 ( .A(n2651), .B(n341), .C(n2652), .D(n391), .Y(n2164) );
  OAI22X1 U1934 ( .A(n2652), .B(n341), .C(n2653), .D(n391), .Y(n2165) );
  OAI22X1 U1935 ( .A(n2653), .B(n341), .C(n2654), .D(n391), .Y(n2166) );
  OAI22X1 U1936 ( .A(n2654), .B(n341), .C(n2655), .D(n391), .Y(n2167) );
  OAI22X1 U1937 ( .A(n2655), .B(n341), .C(n2656), .D(n391), .Y(n2168) );
  OAI22X1 U1938 ( .A(n2656), .B(n341), .C(n2657), .D(n391), .Y(n2169) );
  OAI22X1 U1939 ( .A(n2657), .B(n341), .C(n2658), .D(n391), .Y(n2170) );
  XNOR2X1 U1940 ( .A(n295), .B(n497), .Y(n2627) );
  XNOR2X1 U1941 ( .A(n295), .B(n495), .Y(n2628) );
  XNOR2X1 U1942 ( .A(n295), .B(n2918), .Y(n2629) );
  XNOR2X1 U1943 ( .A(n295), .B(n491), .Y(n2630) );
  XNOR2X1 U1944 ( .A(n295), .B(n2947), .Y(n2631) );
  XNOR2X1 U1945 ( .A(n295), .B(n2914), .Y(n2632) );
  XNOR2X1 U1946 ( .A(n295), .B(n485), .Y(n2633) );
  XNOR2X1 U1947 ( .A(n295), .B(n483), .Y(n2634) );
  XNOR2X1 U1948 ( .A(n295), .B(n2913), .Y(n2635) );
  XNOR2X1 U1949 ( .A(n295), .B(n479), .Y(n2636) );
  XNOR2X1 U1950 ( .A(n295), .B(n477), .Y(n2637) );
  XNOR2X1 U1951 ( .A(n294), .B(n475), .Y(n2638) );
  XNOR2X1 U1952 ( .A(n294), .B(n473), .Y(n2639) );
  XNOR2X1 U1953 ( .A(n294), .B(n471), .Y(n2640) );
  XNOR2X1 U1954 ( .A(n294), .B(n469), .Y(n2641) );
  XNOR2X1 U1955 ( .A(n294), .B(n467), .Y(n2642) );
  XNOR2X1 U1956 ( .A(n294), .B(n465), .Y(n2643) );
  XNOR2X1 U1957 ( .A(n294), .B(n463), .Y(n2644) );
  XNOR2X1 U1958 ( .A(n294), .B(n461), .Y(n2645) );
  XNOR2X1 U1959 ( .A(n294), .B(n459), .Y(n2646) );
  XNOR2X1 U1960 ( .A(n294), .B(n457), .Y(n2647) );
  XNOR2X1 U1961 ( .A(n294), .B(n455), .Y(n2648) );
  XNOR2X1 U1962 ( .A(n294), .B(n453), .Y(n2649) );
  XNOR2X1 U1963 ( .A(n293), .B(n451), .Y(n2650) );
  XNOR2X1 U1964 ( .A(n293), .B(n449), .Y(n2651) );
  XNOR2X1 U1965 ( .A(n293), .B(n447), .Y(n2652) );
  XNOR2X1 U1966 ( .A(n293), .B(n445), .Y(n2653) );
  XNOR2X1 U1967 ( .A(n293), .B(n443), .Y(n2654) );
  XNOR2X1 U1968 ( .A(n293), .B(n441), .Y(n2655) );
  XNOR2X1 U1969 ( .A(n293), .B(n439), .Y(n2656) );
  XNOR2X1 U1970 ( .A(n293), .B(n437), .Y(n2657) );
  XNOR2X1 U1971 ( .A(n293), .B(n2950), .Y(n2658) );
  OAI22X1 U1972 ( .A(n340), .B(n2692), .C(n2810), .D(n390), .Y(n1757) );
  OAI22X1 U1973 ( .A(n2810), .B(n340), .C(n2660), .D(n390), .Y(n2173) );
  OAI22X1 U1974 ( .A(n2660), .B(n340), .C(n2661), .D(n390), .Y(n2174) );
  OAI22X1 U1975 ( .A(n2661), .B(n340), .C(n2662), .D(n390), .Y(n2175) );
  OAI22X1 U1976 ( .A(n2662), .B(n340), .C(n2663), .D(n390), .Y(n2176) );
  OAI22X1 U1977 ( .A(n2663), .B(n340), .C(n2664), .D(n390), .Y(n2177) );
  OAI22X1 U1978 ( .A(n2664), .B(n340), .C(n2665), .D(n390), .Y(n2178) );
  OAI22X1 U1979 ( .A(n2665), .B(n340), .C(n2666), .D(n390), .Y(n2179) );
  OAI22X1 U1980 ( .A(n2666), .B(n340), .C(n2667), .D(n390), .Y(n2180) );
  OAI22X1 U1981 ( .A(n2667), .B(n340), .C(n2668), .D(n390), .Y(n2181) );
  OAI22X1 U1982 ( .A(n2668), .B(n339), .C(n2669), .D(n390), .Y(n2182) );
  OAI22X1 U1983 ( .A(n2669), .B(n339), .C(n2670), .D(n389), .Y(n2183) );
  OAI22X1 U1984 ( .A(n2670), .B(n339), .C(n2671), .D(n389), .Y(n2184) );
  OAI22X1 U1985 ( .A(n2671), .B(n339), .C(n2672), .D(n389), .Y(n2185) );
  OAI22X1 U1986 ( .A(n2672), .B(n339), .C(n2673), .D(n389), .Y(n2186) );
  OAI22X1 U1987 ( .A(n2673), .B(n339), .C(n2674), .D(n389), .Y(n2187) );
  OAI22X1 U1988 ( .A(n2674), .B(n339), .C(n2675), .D(n389), .Y(n2188) );
  OAI22X1 U1989 ( .A(n2675), .B(n339), .C(n2676), .D(n389), .Y(n2189) );
  OAI22X1 U1990 ( .A(n2676), .B(n339), .C(n2677), .D(n389), .Y(n2190) );
  OAI22X1 U1991 ( .A(n2677), .B(n339), .C(n2678), .D(n389), .Y(n2191) );
  OAI22X1 U1992 ( .A(n2678), .B(n339), .C(n2679), .D(n389), .Y(n2192) );
  OAI22X1 U1993 ( .A(n2679), .B(n339), .C(n2680), .D(n389), .Y(n2193) );
  OAI22X1 U1994 ( .A(n2680), .B(n338), .C(n2681), .D(n389), .Y(n2194) );
  OAI22X1 U1995 ( .A(n2681), .B(n338), .C(n2682), .D(n388), .Y(n2195) );
  OAI22X1 U1996 ( .A(n2682), .B(n338), .C(n2683), .D(n388), .Y(n2196) );
  OAI22X1 U1997 ( .A(n2683), .B(n338), .C(n2684), .D(n388), .Y(n2197) );
  OAI22X1 U1998 ( .A(n2684), .B(n338), .C(n2685), .D(n388), .Y(n2198) );
  OAI22X1 U1999 ( .A(n2685), .B(n338), .C(n2686), .D(n388), .Y(n2199) );
  OAI22X1 U2000 ( .A(n2686), .B(n338), .C(n2687), .D(n388), .Y(n2200) );
  OAI22X1 U2001 ( .A(n2687), .B(n338), .C(n2688), .D(n388), .Y(n2201) );
  OAI22X1 U2002 ( .A(n2688), .B(n338), .C(n2689), .D(n388), .Y(n2202) );
  OAI22X1 U2003 ( .A(n2689), .B(n338), .C(n2690), .D(n388), .Y(n2203) );
  OAI22X1 U2004 ( .A(n2690), .B(n338), .C(n2691), .D(n388), .Y(n2204) );
  XNOR2X1 U2005 ( .A(n292), .B(n497), .Y(n2660) );
  XNOR2X1 U2006 ( .A(n292), .B(n495), .Y(n2661) );
  XNOR2X1 U2007 ( .A(n292), .B(n2917), .Y(n2662) );
  XNOR2X1 U2008 ( .A(n292), .B(n491), .Y(n2663) );
  XNOR2X1 U2009 ( .A(n292), .B(n2947), .Y(n2664) );
  XNOR2X1 U2010 ( .A(n292), .B(n2914), .Y(n2665) );
  XNOR2X1 U2011 ( .A(n292), .B(n485), .Y(n2666) );
  XNOR2X1 U2012 ( .A(n292), .B(n483), .Y(n2667) );
  XNOR2X1 U2013 ( .A(n292), .B(n2912), .Y(n2668) );
  XNOR2X1 U2014 ( .A(n292), .B(n479), .Y(n2669) );
  XNOR2X1 U2015 ( .A(n292), .B(n477), .Y(n2670) );
  XNOR2X1 U2016 ( .A(n291), .B(n475), .Y(n2671) );
  XNOR2X1 U2017 ( .A(n291), .B(n473), .Y(n2672) );
  XNOR2X1 U2018 ( .A(n291), .B(n471), .Y(n2673) );
  XNOR2X1 U2019 ( .A(n291), .B(n469), .Y(n2674) );
  XNOR2X1 U2020 ( .A(n291), .B(n467), .Y(n2675) );
  XNOR2X1 U2021 ( .A(n291), .B(n465), .Y(n2676) );
  XNOR2X1 U2022 ( .A(n291), .B(n463), .Y(n2677) );
  XNOR2X1 U2023 ( .A(n291), .B(n461), .Y(n2678) );
  XNOR2X1 U2024 ( .A(n291), .B(n459), .Y(n2679) );
  XNOR2X1 U2025 ( .A(n291), .B(n457), .Y(n2680) );
  XNOR2X1 U2026 ( .A(n291), .B(n455), .Y(n2681) );
  XNOR2X1 U2027 ( .A(n291), .B(n453), .Y(n2682) );
  XNOR2X1 U2028 ( .A(n290), .B(n451), .Y(n2683) );
  XNOR2X1 U2029 ( .A(n290), .B(n449), .Y(n2684) );
  XNOR2X1 U2030 ( .A(n290), .B(n447), .Y(n2685) );
  XNOR2X1 U2031 ( .A(n290), .B(n445), .Y(n2686) );
  XNOR2X1 U2032 ( .A(n290), .B(n443), .Y(n2687) );
  XNOR2X1 U2033 ( .A(n290), .B(n441), .Y(n2688) );
  XNOR2X1 U2034 ( .A(n290), .B(n439), .Y(n2689) );
  XNOR2X1 U2035 ( .A(n290), .B(n437), .Y(n2690) );
  XNOR2X1 U2036 ( .A(n290), .B(n2950), .Y(n2691) );
  OAI22X1 U2037 ( .A(n337), .B(n2725), .C(n2811), .D(n387), .Y(n1758) );
  OAI22X1 U2038 ( .A(n337), .B(n2811), .C(n2693), .D(n387), .Y(n2207) );
  OAI22X1 U2039 ( .A(n337), .B(n2693), .C(n2694), .D(n387), .Y(n2208) );
  OAI22X1 U2040 ( .A(n337), .B(n2694), .C(n2695), .D(n387), .Y(n2209) );
  OAI22X1 U2041 ( .A(n337), .B(n2695), .C(n2696), .D(n387), .Y(n2210) );
  OAI22X1 U2042 ( .A(n337), .B(n2696), .C(n2697), .D(n387), .Y(n2211) );
  OAI22X1 U2043 ( .A(n337), .B(n2697), .C(n2698), .D(n387), .Y(n2212) );
  OAI22X1 U2044 ( .A(n337), .B(n2698), .C(n2699), .D(n387), .Y(n2213) );
  OAI22X1 U2045 ( .A(n337), .B(n2699), .C(n2700), .D(n387), .Y(n2214) );
  OAI22X1 U2046 ( .A(n337), .B(n2700), .C(n2701), .D(n387), .Y(n2215) );
  OAI22X1 U2047 ( .A(n336), .B(n2701), .C(n2702), .D(n387), .Y(n2216) );
  OAI22X1 U2048 ( .A(n336), .B(n2702), .C(n2703), .D(n386), .Y(n2217) );
  OAI22X1 U2049 ( .A(n336), .B(n2703), .C(n2704), .D(n386), .Y(n2218) );
  OAI22X1 U2050 ( .A(n336), .B(n2704), .C(n2705), .D(n386), .Y(n2219) );
  OAI22X1 U2051 ( .A(n336), .B(n2705), .C(n2706), .D(n386), .Y(n2220) );
  OAI22X1 U2052 ( .A(n336), .B(n2706), .C(n2707), .D(n386), .Y(n2221) );
  OAI22X1 U2053 ( .A(n336), .B(n2707), .C(n2708), .D(n386), .Y(n2222) );
  OAI22X1 U2054 ( .A(n336), .B(n2708), .C(n2709), .D(n386), .Y(n2223) );
  OAI22X1 U2055 ( .A(n336), .B(n2709), .C(n2710), .D(n386), .Y(n2224) );
  OAI22X1 U2056 ( .A(n336), .B(n2710), .C(n2711), .D(n386), .Y(n2225) );
  OAI22X1 U2057 ( .A(n336), .B(n2711), .C(n2712), .D(n386), .Y(n2226) );
  OAI22X1 U2058 ( .A(n336), .B(n2712), .C(n2713), .D(n386), .Y(n2227) );
  OAI22X1 U2059 ( .A(n335), .B(n2713), .C(n2714), .D(n386), .Y(n2228) );
  OAI22X1 U2060 ( .A(n335), .B(n2714), .C(n2715), .D(n385), .Y(n2229) );
  OAI22X1 U2061 ( .A(n335), .B(n2715), .C(n2716), .D(n385), .Y(n2230) );
  OAI22X1 U2062 ( .A(n335), .B(n2716), .C(n2717), .D(n385), .Y(n2231) );
  OAI22X1 U2063 ( .A(n335), .B(n2717), .C(n2718), .D(n385), .Y(n2232) );
  OAI22X1 U2064 ( .A(n335), .B(n2718), .C(n2719), .D(n385), .Y(n2233) );
  OAI22X1 U2065 ( .A(n335), .B(n2719), .C(n2720), .D(n385), .Y(n2234) );
  OAI22X1 U2066 ( .A(n335), .B(n2720), .C(n2721), .D(n385), .Y(n2235) );
  OAI22X1 U2067 ( .A(n335), .B(n2721), .C(n2722), .D(n385), .Y(n2236) );
  OAI22X1 U2068 ( .A(n335), .B(n2722), .C(n2723), .D(n385), .Y(n2237) );
  OAI22X1 U2069 ( .A(n335), .B(n2723), .C(n2724), .D(n385), .Y(n2238) );
  XNOR2X1 U2070 ( .A(n289), .B(n497), .Y(n2693) );
  XNOR2X1 U2071 ( .A(n289), .B(n495), .Y(n2694) );
  XNOR2X1 U2072 ( .A(n289), .B(n2916), .Y(n2695) );
  XNOR2X1 U2073 ( .A(n289), .B(n491), .Y(n2696) );
  XNOR2X1 U2074 ( .A(n289), .B(n2947), .Y(n2697) );
  XNOR2X1 U2075 ( .A(n289), .B(n2914), .Y(n2698) );
  XNOR2X1 U2076 ( .A(n289), .B(n485), .Y(n2699) );
  XNOR2X1 U2077 ( .A(n289), .B(n483), .Y(n2700) );
  XNOR2X1 U2078 ( .A(n289), .B(n2912), .Y(n2701) );
  XNOR2X1 U2079 ( .A(n289), .B(n479), .Y(n2702) );
  XNOR2X1 U2080 ( .A(n289), .B(n477), .Y(n2703) );
  XNOR2X1 U2081 ( .A(n288), .B(n475), .Y(n2704) );
  XNOR2X1 U2082 ( .A(n288), .B(n473), .Y(n2705) );
  XNOR2X1 U2083 ( .A(n288), .B(n471), .Y(n2706) );
  XNOR2X1 U2084 ( .A(n288), .B(n469), .Y(n2707) );
  XNOR2X1 U2085 ( .A(n288), .B(n467), .Y(n2708) );
  XNOR2X1 U2086 ( .A(n288), .B(n465), .Y(n2709) );
  XNOR2X1 U2087 ( .A(n288), .B(n463), .Y(n2710) );
  XNOR2X1 U2088 ( .A(n288), .B(n461), .Y(n2711) );
  XNOR2X1 U2089 ( .A(n288), .B(n459), .Y(n2712) );
  XNOR2X1 U2090 ( .A(n288), .B(n457), .Y(n2713) );
  XNOR2X1 U2091 ( .A(n288), .B(n455), .Y(n2714) );
  XNOR2X1 U2092 ( .A(n288), .B(n453), .Y(n2715) );
  XNOR2X1 U2093 ( .A(n287), .B(n451), .Y(n2716) );
  XNOR2X1 U2094 ( .A(n287), .B(n449), .Y(n2717) );
  XNOR2X1 U2095 ( .A(n287), .B(n447), .Y(n2718) );
  XNOR2X1 U2096 ( .A(n287), .B(n445), .Y(n2719) );
  XNOR2X1 U2097 ( .A(n287), .B(n443), .Y(n2720) );
  XNOR2X1 U2098 ( .A(n287), .B(n441), .Y(n2721) );
  XNOR2X1 U2099 ( .A(n287), .B(n439), .Y(n2722) );
  XNOR2X1 U2100 ( .A(n287), .B(n437), .Y(n2723) );
  XNOR2X1 U2101 ( .A(n287), .B(n2950), .Y(n2724) );
  INVX2 U2102 ( .A(n332), .Y(n2796) );
  INVX2 U2104 ( .A(n329), .Y(n2797) );
  INVX2 U2106 ( .A(n326), .Y(n2798) );
  INVX2 U2108 ( .A(n323), .Y(n2799) );
  INVX2 U2110 ( .A(n320), .Y(n2800) );
  INVX2 U2112 ( .A(n317), .Y(n2801) );
  INVX2 U2114 ( .A(n314), .Y(n2802) );
  INVX2 U2116 ( .A(n311), .Y(n2803) );
  INVX2 U2118 ( .A(n308), .Y(n2804) );
  INVX2 U2120 ( .A(n305), .Y(n2805) );
  INVX2 U2122 ( .A(n302), .Y(n2806) );
  INVX2 U2124 ( .A(n299), .Y(n2807) );
  INVX2 U2126 ( .A(n296), .Y(n2808) );
  INVX2 U2128 ( .A(n293), .Y(n2809) );
  INVX2 U2130 ( .A(n290), .Y(n2810) );
  INVX2 U2132 ( .A(n287), .Y(n2811) );
  NAND2X1 U2135 ( .A(n2752), .B(n2780), .Y(n432) );
  XOR2X1 U2136 ( .A(a[30]), .B(a[31]), .Y(n2752) );
  XNOR2X1 U2137 ( .A(a[30]), .B(a[29]), .Y(n2780) );
  NAND2X1 U2138 ( .A(n2753), .B(n2781), .Y(n429) );
  XOR2X1 U2139 ( .A(a[28]), .B(a[29]), .Y(n2753) );
  XNOR2X1 U2140 ( .A(a[28]), .B(a[27]), .Y(n2781) );
  NAND2X1 U2141 ( .A(n2754), .B(n2782), .Y(n426) );
  XOR2X1 U2142 ( .A(a[26]), .B(a[27]), .Y(n2754) );
  XNOR2X1 U2143 ( .A(a[26]), .B(a[25]), .Y(n2782) );
  NAND2X1 U2144 ( .A(n2755), .B(n2783), .Y(n423) );
  XOR2X1 U2145 ( .A(a[24]), .B(a[25]), .Y(n2755) );
  XNOR2X1 U2146 ( .A(a[24]), .B(a[23]), .Y(n2783) );
  NAND2X1 U2147 ( .A(n2756), .B(n2784), .Y(n2768) );
  XOR2X1 U2148 ( .A(a[22]), .B(a[23]), .Y(n2756) );
  XNOR2X1 U2149 ( .A(a[22]), .B(a[21]), .Y(n2784) );
  NAND2X1 U2150 ( .A(n2757), .B(n2785), .Y(n2769) );
  XOR2X1 U2151 ( .A(a[20]), .B(a[21]), .Y(n2757) );
  XNOR2X1 U2152 ( .A(a[20]), .B(a[19]), .Y(n2785) );
  NAND2X1 U2153 ( .A(n2758), .B(n2786), .Y(n2770) );
  XOR2X1 U2154 ( .A(a[18]), .B(a[19]), .Y(n2758) );
  XNOR2X1 U2155 ( .A(a[18]), .B(a[17]), .Y(n2786) );
  NAND2X1 U2156 ( .A(n2759), .B(n2787), .Y(n2771) );
  XOR2X1 U2157 ( .A(a[16]), .B(a[17]), .Y(n2759) );
  XNOR2X1 U2158 ( .A(a[16]), .B(a[15]), .Y(n2787) );
  NAND2X1 U2159 ( .A(n2760), .B(n2788), .Y(n2772) );
  XOR2X1 U2160 ( .A(a[14]), .B(a[15]), .Y(n2760) );
  XNOR2X1 U2161 ( .A(a[14]), .B(a[13]), .Y(n2788) );
  NAND2X1 U2162 ( .A(n2761), .B(n2789), .Y(n2773) );
  XOR2X1 U2163 ( .A(a[12]), .B(a[13]), .Y(n2761) );
  XNOR2X1 U2164 ( .A(a[12]), .B(a[11]), .Y(n2789) );
  NAND2X1 U2165 ( .A(n2762), .B(n2790), .Y(n2774) );
  XOR2X1 U2166 ( .A(a[10]), .B(a[11]), .Y(n2762) );
  XNOR2X1 U2167 ( .A(a[10]), .B(a[9]), .Y(n2790) );
  NAND2X1 U2168 ( .A(n2763), .B(n2791), .Y(n2775) );
  XOR2X1 U2169 ( .A(a[8]), .B(a[9]), .Y(n2763) );
  XNOR2X1 U2170 ( .A(a[8]), .B(a[7]), .Y(n2791) );
  NAND2X1 U2171 ( .A(n2764), .B(n2792), .Y(n2776) );
  XOR2X1 U2172 ( .A(a[6]), .B(a[7]), .Y(n2764) );
  XNOR2X1 U2173 ( .A(a[6]), .B(a[5]), .Y(n2792) );
  NAND2X1 U2174 ( .A(n2765), .B(n2793), .Y(n2777) );
  XOR2X1 U2175 ( .A(a[4]), .B(a[5]), .Y(n2765) );
  XNOR2X1 U2176 ( .A(a[4]), .B(a[3]), .Y(n2793) );
  NAND2X1 U2177 ( .A(n2766), .B(n2794), .Y(n2778) );
  XOR2X1 U2178 ( .A(a[2]), .B(a[3]), .Y(n2766) );
  XNOR2X1 U2179 ( .A(a[2]), .B(a[1]), .Y(n2794) );
  NAND2X1 U2180 ( .A(n2795), .B(n2767), .Y(n2779) );
  XOR2X1 U2181 ( .A(a[0]), .B(a[1]), .Y(n2767) );
  INVX2 U2182 ( .A(a[0]), .Y(n2795) );
  BUFX2 U2185 ( .A(n479), .Y(n2909) );
  BUFX4 U2186 ( .A(b[28]), .Y(n2910) );
  INVX8 U2187 ( .A(n481), .Y(n2911) );
  INVX8 U2188 ( .A(n2911), .Y(n2912) );
  INVX8 U2189 ( .A(n2911), .Y(n2913) );
  INVX4 U2190 ( .A(n2952), .Y(n2951) );
  INVX4 U2191 ( .A(n433), .Y(n2952) );
  BUFX2 U2192 ( .A(n2914), .Y(n2949) );
  INVX2 U2193 ( .A(n698), .Y(n697) );
  BUFX2 U2194 ( .A(b[26]), .Y(n2914) );
  INVX8 U2195 ( .A(n493), .Y(n2915) );
  INVX4 U2196 ( .A(n2915), .Y(n2916) );
  INVX8 U2197 ( .A(n2915), .Y(n2917) );
  INVX4 U2198 ( .A(n2915), .Y(n2918) );
  OR2X2 U2199 ( .A(n1703), .B(n1694), .Y(n2919) );
  OR2X2 U2200 ( .A(n1741), .B(n1740), .Y(n2920) );
  OR2X2 U2201 ( .A(n1719), .B(n1712), .Y(n2921) );
  OR2X2 U2202 ( .A(n1711), .B(n1704), .Y(n2922) );
  OR2X2 U2203 ( .A(n1645), .B(n1632), .Y(n2923) );
  OR2X2 U2204 ( .A(n1455), .B(n1432), .Y(n2924) );
  INVX2 U2205 ( .A(n650), .Y(n648) );
  OR2X2 U2206 ( .A(n1631), .B(n1616), .Y(n2925) );
  OR2X2 U2207 ( .A(n1501), .B(n1480), .Y(n2926) );
  OR2X2 U2208 ( .A(n2237), .B(n2944), .Y(n2927) );
  OR2X2 U2209 ( .A(n920), .B(n901), .Y(n2928) );
  AND2X2 U2210 ( .A(n2951), .B(n152), .Y(n2929) );
  AND2X2 U2211 ( .A(n2951), .B(n125), .Y(n2930) );
  AND2X2 U2212 ( .A(n2951), .B(n98), .Y(n2931) );
  INVX2 U2213 ( .A(n667), .Y(n665) );
  OR2X2 U2214 ( .A(n900), .B(n891), .Y(n2932) );
  AND2X2 U2215 ( .A(n843), .B(n2945), .Y(product[1]) );
  BUFX2 U2216 ( .A(n2947), .Y(n489) );
  INVX4 U2217 ( .A(n2952), .Y(n2950) );
  INVX2 U2218 ( .A(n593), .Y(n591) );
  INVX1 U2219 ( .A(n602), .Y(n596) );
  INVX1 U2220 ( .A(n666), .Y(n664) );
  INVX1 U2221 ( .A(n623), .Y(n622) );
  INVX1 U2222 ( .A(n2926), .Y(n720) );
  INVX1 U2223 ( .A(n2925), .Y(n761) );
  AND2X2 U2224 ( .A(n2951), .B(n143), .Y(n2935) );
  AND2X2 U2225 ( .A(n2951), .B(n89), .Y(n2937) );
  AND2X2 U2226 ( .A(n2951), .B(n162), .Y(n2936) );
  AND2X2 U2227 ( .A(n2951), .B(n134), .Y(n2938) );
  AND2X2 U2228 ( .A(n2951), .B(n178), .Y(n2939) );
  AND2X2 U2229 ( .A(n2951), .B(n116), .Y(n2942) );
  AND2X2 U2230 ( .A(n2951), .B(n107), .Y(n2940) );
  AND2X2 U2231 ( .A(n2951), .B(n210), .Y(n2941) );
  AND2X2 U2232 ( .A(n2951), .B(n226), .Y(n2943) );
  BUFX2 U2233 ( .A(b[0]), .Y(n433) );
  AND2X2 U2234 ( .A(n2951), .B(a[0]), .Y(product[0]) );
  INVX2 U2235 ( .A(n581), .Y(n579) );
  INVX1 U2236 ( .A(n631), .Y(n629) );
  INVX2 U2237 ( .A(n582), .Y(n580) );
  INVX1 U2238 ( .A(n634), .Y(n632) );
  INVX1 U2239 ( .A(n601), .Y(n599) );
  OR2X2 U2240 ( .A(n554), .B(n581), .Y(n2934) );
  INVX1 U2241 ( .A(n643), .Y(n641) );
  INVX2 U2242 ( .A(n592), .Y(n590) );
  INVX2 U2243 ( .A(n574), .Y(n572) );
  INVX1 U2244 ( .A(n695), .Y(n693) );
  INVX1 U2245 ( .A(n696), .Y(n694) );
  INVX2 U2246 ( .A(n575), .Y(n573) );
  INVX2 U2247 ( .A(n668), .Y(n666) );
  INVX1 U2248 ( .A(n669), .Y(n667) );
  INVX1 U2249 ( .A(n624), .Y(n623) );
  INVX1 U2250 ( .A(n759), .Y(n757) );
  INVX1 U2251 ( .A(n718), .Y(n716) );
  INVX1 U2252 ( .A(n786), .Y(n785) );
  INVX2 U2253 ( .A(n725), .Y(n723) );
  INVX1 U2254 ( .A(n745), .Y(n743) );
  INVX1 U2255 ( .A(n661), .Y(n659) );
  INVX1 U2256 ( .A(n746), .Y(n744) );
  INVX2 U2257 ( .A(n717), .Y(n715) );
  INVX2 U2258 ( .A(n758), .Y(n756) );
  INVX1 U2259 ( .A(n706), .Y(n704) );
  INVX2 U2260 ( .A(n711), .Y(n709) );
  INVX2 U2261 ( .A(n553), .Y(n551) );
  INVX2 U2262 ( .A(n559), .Y(n557) );
  INVX1 U2263 ( .A(n801), .Y(n799) );
  INVX2 U2264 ( .A(n766), .Y(n764) );
  INVX1 U2265 ( .A(n783), .Y(n781) );
  INVX1 U2266 ( .A(n784), .Y(n782) );
  INVX2 U2267 ( .A(n806), .Y(n804) );
  INVX1 U2268 ( .A(n774), .Y(n772) );
  INVX1 U2269 ( .A(n812), .Y(n810) );
  INVX1 U2270 ( .A(n825), .Y(n824) );
  INVX1 U2271 ( .A(n832), .Y(n830) );
  INVX1 U2272 ( .A(n840), .Y(n838) );
  INVX2 U2273 ( .A(n843), .Y(n841) );
  INVX2 U2274 ( .A(n433), .Y(n2953) );
  BUFX4 U2275 ( .A(b[15]), .Y(n465) );
  BUFX4 U2276 ( .A(b[13]), .Y(n461) );
  BUFX4 U2277 ( .A(b[14]), .Y(n463) );
  BUFX4 U2278 ( .A(b[1]), .Y(n437) );
  BUFX4 U2279 ( .A(b[2]), .Y(n439) );
  BUFX4 U2280 ( .A(b[10]), .Y(n455) );
  BUFX4 U2281 ( .A(b[8]), .Y(n451) );
  BUFX4 U2282 ( .A(b[11]), .Y(n457) );
  BUFX4 U2283 ( .A(b[5]), .Y(n445) );
  BUFX4 U2284 ( .A(b[3]), .Y(n441) );
  BUFX4 U2285 ( .A(b[4]), .Y(n443) );
  BUFX4 U2286 ( .A(b[6]), .Y(n447) );
  BUFX4 U2287 ( .A(b[9]), .Y(n453) );
  BUFX4 U2288 ( .A(b[12]), .Y(n459) );
  BUFX4 U2289 ( .A(b[7]), .Y(n449) );
  BUFX4 U2290 ( .A(b[17]), .Y(n469) );
  BUFX4 U2291 ( .A(b[16]), .Y(n467) );
  BUFX4 U2292 ( .A(b[18]), .Y(n471) );
  BUFX4 U2293 ( .A(b[19]), .Y(n473) );
  BUFX4 U2294 ( .A(b[21]), .Y(n477) );
  BUFX4 U2295 ( .A(b[20]), .Y(n475) );
  BUFX4 U2296 ( .A(b[23]), .Y(n481) );
  BUFX4 U2297 ( .A(b[22]), .Y(n479) );
  BUFX4 U2298 ( .A(b[25]), .Y(n485) );
  BUFX4 U2299 ( .A(b[24]), .Y(n483) );
  AND2X1 U2300 ( .A(n2951), .B(n258), .Y(n2944) );
  OR2X2 U2301 ( .A(n1758), .B(n2238), .Y(n2945) );
  BUFX2 U2302 ( .A(n334), .Y(n332) );
  BUFX2 U2303 ( .A(n334), .Y(n333) );
  BUFX2 U2304 ( .A(n2796), .Y(n383) );
  BUFX2 U2305 ( .A(n331), .Y(n329) );
  BUFX2 U2306 ( .A(n2780), .Y(n380) );
  BUFX2 U2307 ( .A(n429), .Y(n427) );
  BUFX2 U2308 ( .A(n432), .Y(n430) );
  BUFX2 U2309 ( .A(a[31]), .Y(n334) );
  BUFX2 U2310 ( .A(n2780), .Y(n382) );
  BUFX2 U2311 ( .A(n2813), .Y(n321) );
  BUFX2 U2312 ( .A(n2812), .Y(n324) );
  BUFX2 U2313 ( .A(n328), .Y(n327) );
  BUFX2 U2314 ( .A(n331), .Y(n330) );
  BUFX2 U2315 ( .A(n2813), .Y(n320) );
  BUFX2 U2316 ( .A(n2814), .Y(n317) );
  BUFX2 U2317 ( .A(n2812), .Y(n323) );
  BUFX2 U2318 ( .A(n328), .Y(n326) );
  BUFX2 U2319 ( .A(n2814), .Y(n319) );
  BUFX2 U2320 ( .A(n2768), .Y(n419) );
  BUFX2 U2321 ( .A(n423), .Y(n422) );
  BUFX2 U2322 ( .A(n2783), .Y(n372) );
  BUFX2 U2323 ( .A(n426), .Y(n425) );
  BUFX2 U2324 ( .A(n2784), .Y(n368) );
  BUFX2 U2325 ( .A(n2783), .Y(n371) );
  BUFX2 U2326 ( .A(n2782), .Y(n374) );
  BUFX2 U2327 ( .A(n2781), .Y(n377) );
  BUFX2 U2328 ( .A(n2769), .Y(n415) );
  BUFX2 U2329 ( .A(n2768), .Y(n418) );
  BUFX2 U2330 ( .A(n423), .Y(n421) );
  BUFX2 U2331 ( .A(n426), .Y(n424) );
  BUFX2 U2332 ( .A(n2782), .Y(n375) );
  BUFX2 U2333 ( .A(n429), .Y(n428) );
  BUFX2 U2334 ( .A(n2813), .Y(n322) );
  BUFX2 U2335 ( .A(n2781), .Y(n378) );
  BUFX2 U2336 ( .A(n432), .Y(n431) );
  BUFX2 U2337 ( .A(n2769), .Y(n417) );
  BUFX2 U2338 ( .A(n2780), .Y(n381) );
  BUFX2 U2339 ( .A(n2812), .Y(n325) );
  BUFX2 U2340 ( .A(n2768), .Y(n420) );
  BUFX2 U2341 ( .A(n2784), .Y(n370) );
  BUFX2 U2342 ( .A(n2781), .Y(n379) );
  BUFX2 U2343 ( .A(n2782), .Y(n376) );
  BUFX2 U2344 ( .A(n2783), .Y(n373) );
  BUFX2 U2345 ( .A(n2817), .Y(n309) );
  BUFX2 U2346 ( .A(n2815), .Y(n315) );
  BUFX2 U2347 ( .A(n2816), .Y(n312) );
  BUFX2 U2348 ( .A(n2814), .Y(n318) );
  BUFX2 U2349 ( .A(n2817), .Y(n310) );
  BUFX2 U2350 ( .A(n2816), .Y(n313) );
  BUFX2 U2351 ( .A(n2815), .Y(n314) );
  BUFX2 U2352 ( .A(n2816), .Y(n311) );
  BUFX2 U2353 ( .A(n2817), .Y(n308) );
  BUFX2 U2354 ( .A(n2815), .Y(n316) );
  BUFX2 U2355 ( .A(n2772), .Y(n408) );
  BUFX2 U2356 ( .A(n2772), .Y(n407) );
  BUFX2 U2357 ( .A(n2771), .Y(n410) );
  BUFX2 U2358 ( .A(n2770), .Y(n413) );
  BUFX2 U2359 ( .A(n2769), .Y(n416) );
  BUFX2 U2360 ( .A(n2787), .Y(n360) );
  BUFX2 U2361 ( .A(n2786), .Y(n363) );
  BUFX2 U2362 ( .A(n2785), .Y(n366) );
  BUFX2 U2363 ( .A(n2784), .Y(n369) );
  BUFX2 U2364 ( .A(n2787), .Y(n359) );
  BUFX2 U2365 ( .A(n2786), .Y(n362) );
  BUFX2 U2366 ( .A(n2785), .Y(n365) );
  BUFX2 U2367 ( .A(n2772), .Y(n406) );
  BUFX2 U2368 ( .A(n2771), .Y(n409) );
  BUFX2 U2369 ( .A(n2770), .Y(n412) );
  BUFX2 U2370 ( .A(n2771), .Y(n411) );
  BUFX2 U2371 ( .A(n2787), .Y(n361) );
  BUFX2 U2372 ( .A(n2770), .Y(n414) );
  BUFX2 U2373 ( .A(n2786), .Y(n364) );
  BUFX2 U2374 ( .A(n2785), .Y(n367) );
  BUFX2 U2375 ( .A(n2819), .Y(n303) );
  BUFX2 U2376 ( .A(n2818), .Y(n306) );
  BUFX2 U2377 ( .A(n2821), .Y(n297) );
  BUFX2 U2378 ( .A(n2820), .Y(n300) );
  BUFX2 U2379 ( .A(n2821), .Y(n298) );
  BUFX2 U2380 ( .A(n2819), .Y(n304) );
  BUFX2 U2381 ( .A(n2820), .Y(n301) );
  BUFX2 U2382 ( .A(n2818), .Y(n307) );
  BUFX2 U2383 ( .A(n2821), .Y(n296) );
  BUFX2 U2384 ( .A(n2818), .Y(n305) );
  BUFX2 U2385 ( .A(n2820), .Y(n299) );
  BUFX2 U2386 ( .A(n2819), .Y(n302) );
  BUFX2 U2387 ( .A(n2775), .Y(n399) );
  BUFX2 U2388 ( .A(n2773), .Y(n405) );
  BUFX2 U2389 ( .A(n2774), .Y(n402) );
  BUFX2 U2390 ( .A(n2776), .Y(n395) );
  BUFX2 U2391 ( .A(n2775), .Y(n398) );
  BUFX2 U2392 ( .A(n2773), .Y(n404) );
  BUFX2 U2393 ( .A(n2774), .Y(n401) );
  BUFX2 U2394 ( .A(n2791), .Y(n348) );
  BUFX2 U2395 ( .A(n2789), .Y(n354) );
  BUFX2 U2396 ( .A(n2788), .Y(n357) );
  BUFX2 U2397 ( .A(n2790), .Y(n351) );
  BUFX2 U2398 ( .A(n2789), .Y(n355) );
  BUFX2 U2399 ( .A(n2790), .Y(n352) );
  BUFX2 U2400 ( .A(n2788), .Y(n358) );
  BUFX2 U2401 ( .A(n2789), .Y(n353) );
  BUFX2 U2402 ( .A(n2791), .Y(n347) );
  BUFX2 U2403 ( .A(n2790), .Y(n350) );
  BUFX2 U2404 ( .A(n2788), .Y(n356) );
  BUFX2 U2405 ( .A(n2776), .Y(n394) );
  BUFX2 U2406 ( .A(n2773), .Y(n403) );
  BUFX2 U2407 ( .A(n2775), .Y(n397) );
  BUFX2 U2408 ( .A(n2774), .Y(n400) );
  BUFX2 U2409 ( .A(n2823), .Y(n291) );
  BUFX2 U2410 ( .A(n2824), .Y(n288) );
  BUFX2 U2411 ( .A(n2822), .Y(n294) );
  BUFX2 U2412 ( .A(n2822), .Y(n295) );
  BUFX2 U2413 ( .A(n2824), .Y(n289) );
  BUFX2 U2414 ( .A(n2823), .Y(n292) );
  BUFX2 U2415 ( .A(n2823), .Y(n290) );
  BUFX2 U2416 ( .A(n2822), .Y(n293) );
  BUFX2 U2417 ( .A(n2824), .Y(n287) );
  BUFX2 U2418 ( .A(n2777), .Y(n393) );
  BUFX2 U2419 ( .A(n2778), .Y(n390) );
  BUFX2 U2420 ( .A(n2776), .Y(n396) );
  BUFX2 U2421 ( .A(n2778), .Y(n389) );
  BUFX2 U2422 ( .A(n2777), .Y(n392) );
  BUFX2 U2423 ( .A(n2794), .Y(n339) );
  BUFX2 U2424 ( .A(n2793), .Y(n342) );
  BUFX2 U2425 ( .A(n2792), .Y(n345) );
  BUFX2 U2426 ( .A(n2793), .Y(n343) );
  BUFX2 U2427 ( .A(n2794), .Y(n340) );
  BUFX2 U2428 ( .A(n2792), .Y(n346) );
  BUFX2 U2429 ( .A(n2791), .Y(n349) );
  BUFX2 U2430 ( .A(n2794), .Y(n338) );
  BUFX2 U2431 ( .A(n2793), .Y(n341) );
  BUFX2 U2432 ( .A(n2792), .Y(n344) );
  BUFX2 U2433 ( .A(n2777), .Y(n391) );
  BUFX2 U2434 ( .A(n2778), .Y(n388) );
  BUFX2 U2435 ( .A(a[29]), .Y(n331) );
  BUFX2 U2436 ( .A(a[27]), .Y(n328) );
  BUFX2 U2437 ( .A(a[23]), .Y(n2813) );
  BUFX2 U2438 ( .A(a[21]), .Y(n2814) );
  BUFX2 U2439 ( .A(a[25]), .Y(n2812) );
  BUFX2 U2440 ( .A(a[15]), .Y(n2817) );
  BUFX2 U2441 ( .A(a[17]), .Y(n2816) );
  BUFX2 U2442 ( .A(a[19]), .Y(n2815) );
  BUFX2 U2443 ( .A(a[7]), .Y(n2821) );
  BUFX2 U2444 ( .A(a[11]), .Y(n2819) );
  BUFX2 U2445 ( .A(a[9]), .Y(n2820) );
  BUFX2 U2446 ( .A(a[13]), .Y(n2818) );
  BUFX2 U2447 ( .A(n2779), .Y(n387) );
  BUFX2 U2448 ( .A(n2779), .Y(n386) );
  BUFX2 U2449 ( .A(n2795), .Y(n337) );
  BUFX2 U2450 ( .A(n2795), .Y(n336) );
  BUFX2 U2451 ( .A(n2795), .Y(n335) );
  BUFX2 U2452 ( .A(n2779), .Y(n385) );
  BUFX2 U2453 ( .A(a[3]), .Y(n2823) );
  BUFX2 U2454 ( .A(a[5]), .Y(n2822) );
  BUFX2 U2455 ( .A(a[1]), .Y(n2824) );
  BUFX4 U2456 ( .A(b[27]), .Y(n2947) );
  BUFX4 U2457 ( .A(b[29]), .Y(n2948) );
  BUFX4 U2458 ( .A(b[31]), .Y(n497) );
  INVX2 U2459 ( .A(n649), .Y(n647) );
  INVX1 U2460 ( .A(n808), .Y(n807) );
  INVX2 U2461 ( .A(n748), .Y(n747) );
  INVX1 U2462 ( .A(n682), .Y(n860) );
  BUFX4 U2463 ( .A(n2910), .Y(n491) );
  INVX1 U2464 ( .A(n671), .Y(n858) );
  BUFX4 U2465 ( .A(n2948), .Y(n493) );
  INVX1 U2466 ( .A(n819), .Y(n884) );
  INVX2 U2467 ( .A(n727), .Y(n726) );
  INVX2 U2468 ( .A(n705), .Y(n703) );
  BUFX4 U2469 ( .A(n608), .Y(n499) );
  INVX1 U2470 ( .A(n660), .Y(n658) );
  BUFX4 U2471 ( .A(b[30]), .Y(n495) );
  INVX1 U2472 ( .A(n642), .Y(n640) );
  INVX1 U2473 ( .A(n633), .Y(n631) );
  INVX1 U2474 ( .A(n795), .Y(n794) );
  INVX1 U2475 ( .A(n768), .Y(n767) );
  INVX1 U2476 ( .A(n670), .Y(n668) );
endmodule


module poly5_DW01_sub_59 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, \B[0] , n184;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2X1 U1 ( .A(n1), .B(B[31]), .Y(DIFF[31]) );
  XOR2X1 U2 ( .A(n2), .B(B[30]), .Y(DIFF[30]) );
  NOR2X1 U3 ( .A(B[30]), .B(n2), .Y(n1) );
  XNOR2X1 U4 ( .A(n6), .B(B[29]), .Y(DIFF[29]) );
  NAND2X1 U5 ( .A(n24), .B(n3), .Y(n2) );
  NOR2X1 U6 ( .A(n10), .B(n4), .Y(n3) );
  NAND2X1 U7 ( .A(n8), .B(n5), .Y(n4) );
  XNOR2X1 U9 ( .A(n9), .B(B[28]), .Y(DIFF[28]) );
  NOR2X1 U10 ( .A(n23), .B(n7), .Y(n6) );
  NAND2X1 U11 ( .A(n8), .B(n11), .Y(n7) );
  XNOR2X1 U13 ( .A(n14), .B(B[27]), .Y(DIFF[27]) );
  NOR2X1 U14 ( .A(n10), .B(n23), .Y(n9) );
  NAND2X1 U17 ( .A(n19), .B(n13), .Y(n10) );
  NOR2X1 U18 ( .A(B[26]), .B(B[27]), .Y(n13) );
  XNOR2X1 U19 ( .A(n17), .B(B[26]), .Y(DIFF[26]) );
  NOR2X1 U20 ( .A(n15), .B(n23), .Y(n14) );
  NAND2X1 U21 ( .A(n16), .B(n19), .Y(n15) );
  XNOR2X1 U23 ( .A(n22), .B(B[25]), .Y(DIFF[25]) );
  NOR2X1 U24 ( .A(n18), .B(n23), .Y(n17) );
  NOR2X1 U28 ( .A(B[25]), .B(B[24]), .Y(n19) );
  XOR2X1 U29 ( .A(n23), .B(B[24]), .Y(DIFF[24]) );
  NOR2X1 U30 ( .A(B[24]), .B(n23), .Y(n22) );
  XOR2X1 U31 ( .A(n27), .B(B[23]), .Y(DIFF[23]) );
  NOR2X1 U33 ( .A(n36), .B(n25), .Y(n24) );
  NAND2X1 U34 ( .A(n26), .B(n30), .Y(n25) );
  NOR2X1 U35 ( .A(B[23]), .B(B[22]), .Y(n26) );
  XOR2X1 U36 ( .A(n29), .B(B[22]), .Y(DIFF[22]) );
  NAND2X1 U37 ( .A(n35), .B(n28), .Y(n27) );
  NOR2X1 U38 ( .A(B[22]), .B(n31), .Y(n28) );
  XOR2X1 U39 ( .A(n33), .B(B[21]), .Y(DIFF[21]) );
  NAND2X1 U40 ( .A(n30), .B(n35), .Y(n29) );
  NOR2X1 U43 ( .A(B[21]), .B(B[20]), .Y(n30) );
  XNOR2X1 U44 ( .A(n35), .B(B[20]), .Y(DIFF[20]) );
  NAND2X1 U45 ( .A(n34), .B(n35), .Y(n33) );
  XNOR2X1 U47 ( .A(n38), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U49 ( .A(n40), .B(n37), .Y(n36) );
  NOR2X1 U50 ( .A(B[19]), .B(B[18]), .Y(n37) );
  XOR2X1 U51 ( .A(n39), .B(B[18]), .Y(DIFF[18]) );
  NOR2X1 U52 ( .A(B[18]), .B(n39), .Y(n38) );
  XOR2X1 U53 ( .A(B[17]), .B(n41), .Y(DIFF[17]) );
  NOR2X1 U55 ( .A(B[17]), .B(n41), .Y(n40) );
  XNOR2X1 U56 ( .A(B[16]), .B(n43), .Y(DIFF[16]) );
  NAND2X1 U57 ( .A(n43), .B(n42), .Y(n41) );
  XOR2X1 U59 ( .A(n46), .B(B[15]), .Y(DIFF[15]) );
  NOR2X1 U60 ( .A(n51), .B(n44), .Y(n43) );
  NAND2X1 U61 ( .A(n45), .B(n47), .Y(n44) );
  XOR2X1 U63 ( .A(n48), .B(n184), .Y(DIFF[14]) );
  NAND2X1 U64 ( .A(n50), .B(n47), .Y(n46) );
  NOR2X1 U65 ( .A(B[13]), .B(B[14]), .Y(n47) );
  XNOR2X1 U66 ( .A(n50), .B(B[13]), .Y(DIFF[13]) );
  NAND2X1 U67 ( .A(n49), .B(n50), .Y(n48) );
  XNOR2X1 U69 ( .A(n53), .B(B[12]), .Y(DIFF[12]) );
  NAND2X1 U71 ( .A(n55), .B(n52), .Y(n51) );
  NOR2X1 U72 ( .A(B[11]), .B(B[12]), .Y(n52) );
  XOR2X1 U73 ( .A(n54), .B(B[11]), .Y(DIFF[11]) );
  NOR2X1 U74 ( .A(B[11]), .B(n54), .Y(n53) );
  XOR2X1 U75 ( .A(n58), .B(B[10]), .Y(DIFF[10]) );
  NOR2X1 U77 ( .A(n61), .B(n56), .Y(n55) );
  NAND2X1 U78 ( .A(n59), .B(n57), .Y(n56) );
  XNOR2X1 U80 ( .A(n60), .B(B[9]), .Y(DIFF[9]) );
  NAND2X1 U81 ( .A(n59), .B(n60), .Y(n58) );
  XNOR2X1 U83 ( .A(B[8]), .B(n63), .Y(DIFF[8]) );
  NAND2X1 U85 ( .A(n62), .B(n63), .Y(n61) );
  XOR2X1 U87 ( .A(n66), .B(B[7]), .Y(DIFF[7]) );
  NOR2X1 U88 ( .A(n64), .B(n69), .Y(n63) );
  NAND2X1 U89 ( .A(n67), .B(n65), .Y(n64) );
  XNOR2X1 U91 ( .A(n68), .B(B[6]), .Y(DIFF[6]) );
  NAND2X1 U92 ( .A(n67), .B(n68), .Y(n66) );
  XNOR2X1 U94 ( .A(n71), .B(B[5]), .Y(DIFF[5]) );
  NAND2X1 U96 ( .A(n73), .B(n70), .Y(n69) );
  NOR2X1 U97 ( .A(B[4]), .B(B[5]), .Y(n70) );
  XOR2X1 U98 ( .A(n72), .B(B[4]), .Y(DIFF[4]) );
  NOR2X1 U99 ( .A(B[4]), .B(n72), .Y(n71) );
  XOR2X1 U100 ( .A(n76), .B(B[3]), .Y(DIFF[3]) );
  NOR2X1 U102 ( .A(n79), .B(n74), .Y(n73) );
  NAND2X1 U103 ( .A(n75), .B(n77), .Y(n74) );
  XNOR2X1 U105 ( .A(n78), .B(B[2]), .Y(DIFF[2]) );
  NAND2X1 U106 ( .A(n77), .B(n78), .Y(n76) );
  XNOR2X1 U108 ( .A(B[1]), .B(n81), .Y(DIFF[1]) );
  NAND2X1 U110 ( .A(n81), .B(n80), .Y(n79) );
  INVX1 U116 ( .A(n61), .Y(n60) );
  INVX1 U117 ( .A(n55), .Y(n54) );
  INVX1 U118 ( .A(n19), .Y(n18) );
  BUFX2 U119 ( .A(B[14]), .Y(n184) );
  INVX1 U120 ( .A(B[13]), .Y(n49) );
  INVX1 U121 ( .A(n30), .Y(n31) );
  INVX1 U122 ( .A(n51), .Y(n50) );
  INVX1 U123 ( .A(n40), .Y(n39) );
  INVX4 U124 ( .A(n24), .Y(n23) );
  INVX1 U125 ( .A(n36), .Y(n35) );
  INVX1 U126 ( .A(n10), .Y(n11) );
  INVX2 U127 ( .A(\B[0] ), .Y(n81) );
  INVX2 U128 ( .A(B[1]), .Y(n80) );
  INVX2 U129 ( .A(B[28]), .Y(n8) );
  INVX2 U130 ( .A(n79), .Y(n78) );
  INVX2 U131 ( .A(B[2]), .Y(n77) );
  INVX2 U132 ( .A(B[3]), .Y(n75) );
  INVX2 U133 ( .A(n73), .Y(n72) );
  INVX2 U134 ( .A(n69), .Y(n68) );
  INVX2 U135 ( .A(B[6]), .Y(n67) );
  INVX2 U136 ( .A(B[7]), .Y(n65) );
  INVX2 U137 ( .A(B[8]), .Y(n62) );
  INVX2 U138 ( .A(B[9]), .Y(n59) );
  INVX2 U139 ( .A(B[10]), .Y(n57) );
  INVX2 U140 ( .A(B[29]), .Y(n5) );
  INVX2 U141 ( .A(B[15]), .Y(n45) );
  INVX2 U142 ( .A(B[16]), .Y(n42) );
  INVX2 U143 ( .A(B[20]), .Y(n34) );
  INVX2 U144 ( .A(B[26]), .Y(n16) );
endmodule


module poly5_DW01_sub_60 ( A, B, CI, DIFF, CO );
  input [47:0] A;
  input [47:0] B;
  output [47:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n45, n46, n47,
         n48, n49, n50, n51, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n70, n71, n72, n73, n74, n75, n76, n77,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n111, n112, n113, n114, n115, n116, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n273, n274;

  XOR2X1 U3 ( .A(n3), .B(B[47]), .Y(DIFF[47]) );
  XOR2X1 U4 ( .A(n9), .B(B[46]), .Y(DIFF[46]) );
  NAND2X1 U5 ( .A(n274), .B(n2), .Y(n3) );
  NOR2X1 U8 ( .A(n7), .B(n19), .Y(n6) );
  NAND2X1 U9 ( .A(n8), .B(n12), .Y(n7) );
  XOR2X1 U11 ( .A(n13), .B(B[45]), .Y(DIFF[45]) );
  NAND2X1 U12 ( .A(n2), .B(n10), .Y(n9) );
  NOR2X1 U13 ( .A(n11), .B(n17), .Y(n10) );
  NOR2X1 U15 ( .A(B[45]), .B(B[44]), .Y(n12) );
  XOR2X1 U16 ( .A(n15), .B(B[44]), .Y(DIFF[44]) );
  NAND2X1 U17 ( .A(n2), .B(n14), .Y(n13) );
  NOR2X1 U18 ( .A(B[44]), .B(n17), .Y(n14) );
  XOR2X1 U19 ( .A(n21), .B(B[43]), .Y(DIFF[43]) );
  NAND2X1 U20 ( .A(n16), .B(n2), .Y(n15) );
  NAND2X1 U22 ( .A(n18), .B(n32), .Y(n17) );
  NAND2X1 U24 ( .A(n20), .B(n26), .Y(n19) );
  NOR2X1 U25 ( .A(B[43]), .B(B[42]), .Y(n20) );
  XOR2X1 U26 ( .A(n23), .B(B[42]), .Y(DIFF[42]) );
  NAND2X1 U27 ( .A(n2), .B(n22), .Y(n21) );
  NOR2X1 U28 ( .A(B[42]), .B(n25), .Y(n22) );
  XOR2X1 U29 ( .A(n27), .B(B[41]), .Y(DIFF[41]) );
  NAND2X1 U30 ( .A(n24), .B(n2), .Y(n23) );
  NAND2X1 U32 ( .A(n26), .B(n32), .Y(n25) );
  NOR2X1 U33 ( .A(B[41]), .B(B[40]), .Y(n26) );
  XOR2X1 U34 ( .A(n29), .B(B[40]), .Y(DIFF[40]) );
  NAND2X1 U35 ( .A(n28), .B(n2), .Y(n27) );
  NOR2X1 U36 ( .A(B[40]), .B(n31), .Y(n28) );
  XOR2X1 U37 ( .A(n35), .B(B[39]), .Y(DIFF[39]) );
  NAND2X1 U38 ( .A(n32), .B(n2), .Y(n29) );
  NOR2X1 U41 ( .A(n33), .B(n47), .Y(n32) );
  NAND2X1 U42 ( .A(n34), .B(n40), .Y(n33) );
  NOR2X1 U43 ( .A(B[39]), .B(B[38]), .Y(n34) );
  XOR2X1 U44 ( .A(n37), .B(B[38]), .Y(DIFF[38]) );
  NAND2X1 U45 ( .A(n36), .B(n1), .Y(n35) );
  NOR2X1 U46 ( .A(B[38]), .B(n39), .Y(n36) );
  XOR2X1 U47 ( .A(n41), .B(B[37]), .Y(DIFF[37]) );
  NAND2X1 U48 ( .A(n38), .B(n1), .Y(n37) );
  NAND2X1 U50 ( .A(n40), .B(n46), .Y(n39) );
  NOR2X1 U51 ( .A(B[37]), .B(B[36]), .Y(n40) );
  XOR2X1 U52 ( .A(n43), .B(B[36]), .Y(DIFF[36]) );
  NAND2X1 U53 ( .A(n42), .B(n1), .Y(n41) );
  NOR2X1 U54 ( .A(B[36]), .B(n45), .Y(n42) );
  XOR2X1 U55 ( .A(n49), .B(B[35]), .Y(DIFF[35]) );
  NAND2X1 U56 ( .A(n46), .B(n1), .Y(n43) );
  NAND2X1 U60 ( .A(n48), .B(n54), .Y(n47) );
  NOR2X1 U61 ( .A(B[35]), .B(B[34]), .Y(n48) );
  XOR2X1 U62 ( .A(n51), .B(B[34]), .Y(DIFF[34]) );
  NAND2X1 U63 ( .A(n50), .B(n1), .Y(n49) );
  NOR2X1 U64 ( .A(B[34]), .B(n53), .Y(n50) );
  XOR2X1 U65 ( .A(n55), .B(B[33]), .Y(DIFF[33]) );
  NAND2X1 U66 ( .A(n54), .B(n1), .Y(n51) );
  NOR2X1 U69 ( .A(B[33]), .B(B[32]), .Y(n54) );
  XNOR2X1 U70 ( .A(n1), .B(B[32]), .Y(DIFF[32]) );
  NAND2X1 U71 ( .A(n56), .B(n1), .Y(n55) );
  XOR2X1 U73 ( .A(n62), .B(n273), .Y(DIFF[31]) );
  NOR2X1 U74 ( .A(n123), .B(n58), .Y(n57) );
  NAND2X1 U75 ( .A(n59), .B(n97), .Y(n58) );
  NOR2X1 U76 ( .A(n60), .B(n80), .Y(n59) );
  NAND2X1 U77 ( .A(n61), .B(n71), .Y(n60) );
  NOR2X1 U78 ( .A(B[31]), .B(B[30]), .Y(n61) );
  XOR2X1 U79 ( .A(n66), .B(B[30]), .Y(DIFF[30]) );
  NAND2X1 U80 ( .A(n122), .B(n63), .Y(n62) );
  NOR2X1 U81 ( .A(n64), .B(n96), .Y(n63) );
  NAND2X1 U82 ( .A(n79), .B(n65), .Y(n64) );
  NOR2X1 U83 ( .A(B[30]), .B(n70), .Y(n65) );
  XOR2X1 U84 ( .A(n72), .B(B[29]), .Y(DIFF[29]) );
  NAND2X1 U85 ( .A(n122), .B(n67), .Y(n66) );
  NOR2X1 U86 ( .A(n68), .B(n96), .Y(n67) );
  NAND2X1 U87 ( .A(n71), .B(n79), .Y(n68) );
  NOR2X1 U90 ( .A(B[29]), .B(B[28]), .Y(n71) );
  XOR2X1 U91 ( .A(n76), .B(B[28]), .Y(DIFF[28]) );
  NAND2X1 U92 ( .A(n122), .B(n73), .Y(n72) );
  NOR2X1 U93 ( .A(n74), .B(n96), .Y(n73) );
  NAND2X1 U94 ( .A(n75), .B(n79), .Y(n74) );
  XOR2X1 U96 ( .A(n82), .B(B[27]), .Y(DIFF[27]) );
  NAND2X1 U97 ( .A(n122), .B(n77), .Y(n76) );
  NOR2X1 U98 ( .A(n80), .B(n96), .Y(n77) );
  NAND2X1 U101 ( .A(n81), .B(n91), .Y(n80) );
  NOR2X1 U102 ( .A(B[27]), .B(B[26]), .Y(n81) );
  XOR2X1 U103 ( .A(n86), .B(B[26]), .Y(DIFF[26]) );
  NAND2X1 U104 ( .A(n122), .B(n83), .Y(n82) );
  NOR2X1 U105 ( .A(n84), .B(n96), .Y(n83) );
  NAND2X1 U106 ( .A(n85), .B(n91), .Y(n84) );
  XOR2X1 U108 ( .A(n92), .B(B[25]), .Y(DIFF[25]) );
  NAND2X1 U109 ( .A(n122), .B(n87), .Y(n86) );
  NOR2X1 U110 ( .A(n90), .B(n96), .Y(n87) );
  NOR2X1 U114 ( .A(B[25]), .B(B[24]), .Y(n91) );
  XOR2X1 U115 ( .A(n94), .B(B[24]), .Y(DIFF[24]) );
  NAND2X1 U116 ( .A(n122), .B(n93), .Y(n92) );
  NOR2X1 U117 ( .A(B[24]), .B(n96), .Y(n93) );
  XOR2X1 U118 ( .A(n100), .B(B[23]), .Y(DIFF[23]) );
  NAND2X1 U119 ( .A(n97), .B(n122), .Y(n94) );
  NOR2X1 U122 ( .A(n98), .B(n112), .Y(n97) );
  NAND2X1 U123 ( .A(n99), .B(n105), .Y(n98) );
  NOR2X1 U124 ( .A(B[23]), .B(B[22]), .Y(n99) );
  XOR2X1 U125 ( .A(n102), .B(B[22]), .Y(DIFF[22]) );
  NAND2X1 U126 ( .A(n122), .B(n101), .Y(n100) );
  NOR2X1 U127 ( .A(B[22]), .B(n104), .Y(n101) );
  XOR2X1 U128 ( .A(n106), .B(B[21]), .Y(DIFF[21]) );
  NAND2X1 U129 ( .A(n103), .B(n122), .Y(n102) );
  NAND2X1 U131 ( .A(n105), .B(n111), .Y(n104) );
  NOR2X1 U132 ( .A(B[21]), .B(B[20]), .Y(n105) );
  XOR2X1 U133 ( .A(n108), .B(B[20]), .Y(DIFF[20]) );
  NAND2X1 U134 ( .A(n107), .B(n122), .Y(n106) );
  NOR2X1 U135 ( .A(B[20]), .B(n112), .Y(n107) );
  XOR2X1 U136 ( .A(n114), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U137 ( .A(n111), .B(n122), .Y(n108) );
  NAND2X1 U141 ( .A(n113), .B(n119), .Y(n112) );
  NOR2X1 U142 ( .A(B[19]), .B(B[18]), .Y(n113) );
  XOR2X1 U143 ( .A(n116), .B(B[18]), .Y(DIFF[18]) );
  NAND2X1 U144 ( .A(n115), .B(n122), .Y(n114) );
  NOR2X1 U145 ( .A(B[18]), .B(n118), .Y(n115) );
  XOR2X1 U146 ( .A(n120), .B(B[17]), .Y(DIFF[17]) );
  NAND2X1 U147 ( .A(n119), .B(n122), .Y(n116) );
  NOR2X1 U150 ( .A(B[17]), .B(B[16]), .Y(n119) );
  XNOR2X1 U151 ( .A(n122), .B(B[16]), .Y(DIFF[16]) );
  NAND2X1 U152 ( .A(n121), .B(n122), .Y(n120) );
  NAND2X1 U155 ( .A(n131), .B(n124), .Y(n123) );
  NOR2X1 U156 ( .A(n125), .B(n128), .Y(n124) );
  NAND2X1 U157 ( .A(n126), .B(n127), .Y(n125) );
  NOR2X1 U158 ( .A(B[15]), .B(B[14]), .Y(n126) );
  NOR2X1 U159 ( .A(B[13]), .B(B[12]), .Y(n127) );
  NAND2X1 U160 ( .A(n129), .B(n130), .Y(n128) );
  NOR2X1 U161 ( .A(B[11]), .B(B[10]), .Y(n129) );
  NOR2X1 U162 ( .A(B[9]), .B(B[8]), .Y(n130) );
  NOR2X1 U163 ( .A(n135), .B(n132), .Y(n131) );
  NAND2X1 U164 ( .A(n133), .B(n134), .Y(n132) );
  NOR2X1 U165 ( .A(B[7]), .B(B[6]), .Y(n133) );
  NOR2X1 U166 ( .A(B[5]), .B(B[4]), .Y(n134) );
  NAND2X1 U167 ( .A(n137), .B(n136), .Y(n135) );
  NOR2X1 U168 ( .A(B[3]), .B(B[2]), .Y(n136) );
  NOR2X1 U169 ( .A(B[0]), .B(B[1]), .Y(n137) );
  BUFX2 U173 ( .A(B[31]), .Y(n273) );
  INVX2 U174 ( .A(n47), .Y(n46) );
  AND2X2 U175 ( .A(n6), .B(n32), .Y(n274) );
  INVX1 U176 ( .A(n71), .Y(n70) );
  INVX2 U177 ( .A(n97), .Y(n96) );
  INVX1 U178 ( .A(n80), .Y(n79) );
  INVX1 U179 ( .A(n112), .Y(n111) );
  INVX1 U180 ( .A(n91), .Y(n90) );
  INVX1 U181 ( .A(B[46]), .Y(n8) );
  INVX1 U182 ( .A(n119), .Y(n118) );
  INVX1 U183 ( .A(n12), .Y(n11) );
  INVX1 U184 ( .A(B[32]), .Y(n56) );
  INVX1 U185 ( .A(B[28]), .Y(n75) );
  INVX1 U186 ( .A(B[26]), .Y(n85) );
  INVX1 U187 ( .A(n104), .Y(n103) );
  INVX1 U188 ( .A(B[16]), .Y(n121) );
  INVX2 U189 ( .A(n123), .Y(n122) );
  INVX2 U190 ( .A(n46), .Y(n45) );
  BUFX2 U191 ( .A(n57), .Y(n2) );
  INVX1 U192 ( .A(n25), .Y(n24) );
  INVX2 U193 ( .A(n32), .Y(n31) );
  INVX1 U194 ( .A(n19), .Y(n18) );
  INVX1 U195 ( .A(n17), .Y(n16) );
  INVX1 U196 ( .A(n39), .Y(n38) );
  INVX1 U197 ( .A(n54), .Y(n53) );
  BUFX4 U198 ( .A(n57), .Y(n1) );
endmodule


module poly5_DW01_add_19 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n168, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n193, n194, n195, n196, n197, n198,
         n199, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n281, n284, n286,
         n288, n290, n292, n294, n296, n297, n298, n300, n302, n304, n305,
         n306, n307, n308, n310, n311, n312, n417, n418, n420;

  XNOR2X1 U5 ( .A(n41), .B(n7), .Y(SUM[31]) );
  NAND2X1 U6 ( .A(n40), .B(n420), .Y(n7) );
  NAND2X1 U9 ( .A(B[31]), .B(A[31]), .Y(n40) );
  XNOR2X1 U10 ( .A(n52), .B(n8), .Y(SUM[30]) );
  OAI21X1 U11 ( .A(n42), .B(n2), .C(n43), .Y(n41) );
  NAND2X1 U12 ( .A(n44), .B(n4), .Y(n42) );
  AOI21X1 U13 ( .A(n3), .B(n44), .C(n45), .Y(n43) );
  NOR2X1 U14 ( .A(n46), .B(n6), .Y(n44) );
  OAI21X1 U15 ( .A(n46), .B(n5), .C(n47), .Y(n45) );
  NAND2X1 U16 ( .A(n417), .B(n59), .Y(n46) );
  AOI21X1 U17 ( .A(n417), .B(n60), .C(n49), .Y(n47) );
  NAND2X1 U20 ( .A(n51), .B(n417), .Y(n8) );
  NAND2X1 U23 ( .A(B[30]), .B(A[30]), .Y(n51) );
  XNOR2X1 U24 ( .A(n63), .B(n9), .Y(SUM[29]) );
  OAI21X1 U25 ( .A(n53), .B(n2), .C(n54), .Y(n52) );
  NAND2X1 U26 ( .A(n55), .B(n4), .Y(n53) );
  AOI21X1 U27 ( .A(n3), .B(n55), .C(n56), .Y(n54) );
  NOR2X1 U28 ( .A(n57), .B(n6), .Y(n55) );
  OAI21X1 U29 ( .A(n57), .B(n5), .C(n58), .Y(n56) );
  NOR2X1 U32 ( .A(n61), .B(n70), .Y(n59) );
  OAI21X1 U33 ( .A(n71), .B(n61), .C(n62), .Y(n60) );
  NAND2X1 U34 ( .A(n62), .B(n284), .Y(n9) );
  NOR2X1 U36 ( .A(B[29]), .B(A[29]), .Y(n61) );
  NAND2X1 U37 ( .A(B[29]), .B(A[29]), .Y(n62) );
  XNOR2X1 U38 ( .A(n72), .B(n10), .Y(SUM[28]) );
  OAI21X1 U39 ( .A(n64), .B(n2), .C(n65), .Y(n63) );
  NAND2X1 U40 ( .A(n66), .B(n4), .Y(n64) );
  AOI21X1 U41 ( .A(n3), .B(n66), .C(n67), .Y(n65) );
  NOR2X1 U42 ( .A(n68), .B(n6), .Y(n66) );
  OAI21X1 U43 ( .A(n68), .B(n5), .C(n71), .Y(n67) );
  NAND2X1 U46 ( .A(n71), .B(n69), .Y(n10) );
  NOR2X1 U48 ( .A(B[28]), .B(A[28]), .Y(n70) );
  NAND2X1 U49 ( .A(B[28]), .B(A[28]), .Y(n71) );
  XNOR2X1 U50 ( .A(n81), .B(n11), .Y(SUM[27]) );
  OAI21X1 U51 ( .A(n73), .B(n2), .C(n74), .Y(n72) );
  NAND2X1 U52 ( .A(n75), .B(n4), .Y(n73) );
  AOI21X1 U53 ( .A(n75), .B(n3), .C(n76), .Y(n74) );
  NAND2X1 U56 ( .A(n77), .B(n97), .Y(n6) );
  AOI21X1 U57 ( .A(n98), .B(n77), .C(n78), .Y(n5) );
  NOR2X1 U58 ( .A(n79), .B(n88), .Y(n77) );
  OAI21X1 U59 ( .A(n89), .B(n79), .C(n80), .Y(n78) );
  NAND2X1 U60 ( .A(n80), .B(n286), .Y(n11) );
  NOR2X1 U62 ( .A(B[27]), .B(A[27]), .Y(n79) );
  NAND2X1 U63 ( .A(B[27]), .B(A[27]), .Y(n80) );
  XNOR2X1 U64 ( .A(n90), .B(n12), .Y(SUM[26]) );
  OAI21X1 U65 ( .A(n82), .B(n2), .C(n83), .Y(n81) );
  NAND2X1 U66 ( .A(n84), .B(n4), .Y(n82) );
  AOI21X1 U67 ( .A(n84), .B(n3), .C(n85), .Y(n83) );
  NOR2X1 U68 ( .A(n86), .B(n95), .Y(n84) );
  OAI21X1 U69 ( .A(n86), .B(n96), .C(n89), .Y(n85) );
  NAND2X1 U72 ( .A(n89), .B(n87), .Y(n12) );
  NOR2X1 U74 ( .A(B[26]), .B(A[26]), .Y(n88) );
  NAND2X1 U75 ( .A(B[26]), .B(A[26]), .Y(n89) );
  XNOR2X1 U76 ( .A(n101), .B(n13), .Y(SUM[25]) );
  OAI21X1 U77 ( .A(n91), .B(n2), .C(n92), .Y(n90) );
  NAND2X1 U78 ( .A(n93), .B(n4), .Y(n91) );
  AOI21X1 U79 ( .A(n93), .B(n3), .C(n98), .Y(n92) );
  NOR2X1 U84 ( .A(n99), .B(n106), .Y(n97) );
  OAI21X1 U85 ( .A(n107), .B(n99), .C(n100), .Y(n98) );
  NAND2X1 U86 ( .A(n100), .B(n288), .Y(n13) );
  NOR2X1 U88 ( .A(B[25]), .B(A[25]), .Y(n99) );
  NAND2X1 U89 ( .A(B[25]), .B(A[25]), .Y(n100) );
  XNOR2X1 U90 ( .A(n108), .B(n14), .Y(SUM[24]) );
  OAI21X1 U91 ( .A(n102), .B(n2), .C(n103), .Y(n101) );
  NAND2X1 U92 ( .A(n104), .B(n4), .Y(n102) );
  AOI21X1 U93 ( .A(n104), .B(n3), .C(n105), .Y(n103) );
  NAND2X1 U96 ( .A(n107), .B(n104), .Y(n14) );
  NOR2X1 U98 ( .A(B[24]), .B(A[24]), .Y(n106) );
  NAND2X1 U99 ( .A(B[24]), .B(A[24]), .Y(n107) );
  XNOR2X1 U100 ( .A(n119), .B(n15), .Y(SUM[23]) );
  OAI21X1 U101 ( .A(n109), .B(n2), .C(n110), .Y(n108) );
  NOR2X1 U104 ( .A(n113), .B(n151), .Y(n111) );
  OAI21X1 U105 ( .A(n113), .B(n152), .C(n114), .Y(n112) );
  NAND2X1 U106 ( .A(n115), .B(n135), .Y(n113) );
  AOI21X1 U107 ( .A(n136), .B(n115), .C(n116), .Y(n114) );
  NOR2X1 U108 ( .A(n117), .B(n126), .Y(n115) );
  OAI21X1 U109 ( .A(n127), .B(n117), .C(n118), .Y(n116) );
  NAND2X1 U110 ( .A(n118), .B(n290), .Y(n15) );
  NOR2X1 U112 ( .A(B[23]), .B(A[23]), .Y(n117) );
  NAND2X1 U113 ( .A(B[23]), .B(A[23]), .Y(n118) );
  XNOR2X1 U114 ( .A(n128), .B(n16), .Y(SUM[22]) );
  OAI21X1 U115 ( .A(n120), .B(n1), .C(n121), .Y(n119) );
  NAND2X1 U116 ( .A(n149), .B(n122), .Y(n120) );
  AOI21X1 U117 ( .A(n150), .B(n122), .C(n123), .Y(n121) );
  NOR2X1 U118 ( .A(n124), .B(n133), .Y(n122) );
  OAI21X1 U119 ( .A(n124), .B(n134), .C(n127), .Y(n123) );
  NAND2X1 U122 ( .A(n127), .B(n125), .Y(n16) );
  NOR2X1 U124 ( .A(B[22]), .B(A[22]), .Y(n126) );
  NAND2X1 U125 ( .A(B[22]), .B(A[22]), .Y(n127) );
  XNOR2X1 U126 ( .A(n139), .B(n17), .Y(SUM[21]) );
  OAI21X1 U127 ( .A(n129), .B(n1), .C(n130), .Y(n128) );
  NAND2X1 U128 ( .A(n131), .B(n149), .Y(n129) );
  AOI21X1 U129 ( .A(n131), .B(n150), .C(n136), .Y(n130) );
  NOR2X1 U134 ( .A(n137), .B(n144), .Y(n135) );
  OAI21X1 U135 ( .A(n145), .B(n137), .C(n138), .Y(n136) );
  NAND2X1 U136 ( .A(n138), .B(n292), .Y(n17) );
  INVX2 U137 ( .A(n137), .Y(n292) );
  NOR2X1 U138 ( .A(B[21]), .B(A[21]), .Y(n137) );
  NAND2X1 U139 ( .A(B[21]), .B(A[21]), .Y(n138) );
  XNOR2X1 U140 ( .A(n146), .B(n18), .Y(SUM[20]) );
  OAI21X1 U141 ( .A(n140), .B(n1), .C(n141), .Y(n139) );
  NAND2X1 U142 ( .A(n142), .B(n149), .Y(n140) );
  AOI21X1 U143 ( .A(n142), .B(n150), .C(n143), .Y(n141) );
  NAND2X1 U146 ( .A(n145), .B(n142), .Y(n18) );
  NOR2X1 U148 ( .A(B[20]), .B(A[20]), .Y(n144) );
  NAND2X1 U149 ( .A(B[20]), .B(A[20]), .Y(n145) );
  XNOR2X1 U150 ( .A(n157), .B(n19), .Y(SUM[19]) );
  OAI21X1 U151 ( .A(n151), .B(n1), .C(n148), .Y(n146) );
  NAND2X1 U156 ( .A(n153), .B(n171), .Y(n151) );
  AOI21X1 U157 ( .A(n172), .B(n153), .C(n154), .Y(n152) );
  NOR2X1 U158 ( .A(n155), .B(n162), .Y(n153) );
  OAI21X1 U159 ( .A(n163), .B(n155), .C(n156), .Y(n154) );
  NAND2X1 U160 ( .A(n156), .B(n294), .Y(n19) );
  INVX2 U161 ( .A(n155), .Y(n294) );
  NOR2X1 U162 ( .A(B[19]), .B(A[19]), .Y(n155) );
  NAND2X1 U163 ( .A(B[19]), .B(A[19]), .Y(n156) );
  XNOR2X1 U164 ( .A(n164), .B(n20), .Y(SUM[18]) );
  OAI21X1 U165 ( .A(n158), .B(n1), .C(n159), .Y(n157) );
  NAND2X1 U166 ( .A(n160), .B(n171), .Y(n158) );
  AOI21X1 U167 ( .A(n160), .B(n168), .C(n161), .Y(n159) );
  NAND2X1 U170 ( .A(n163), .B(n160), .Y(n20) );
  NOR2X1 U172 ( .A(B[18]), .B(A[18]), .Y(n162) );
  NAND2X1 U173 ( .A(B[18]), .B(A[18]), .Y(n163) );
  XNOR2X1 U174 ( .A(n175), .B(n21), .Y(SUM[17]) );
  OAI21X1 U175 ( .A(n165), .B(n1), .C(n170), .Y(n164) );
  NOR2X1 U182 ( .A(n173), .B(n176), .Y(n171) );
  OAI21X1 U183 ( .A(n177), .B(n173), .C(n174), .Y(n172) );
  NAND2X1 U184 ( .A(n174), .B(n296), .Y(n21) );
  INVX2 U185 ( .A(n173), .Y(n296) );
  NOR2X1 U186 ( .A(B[17]), .B(A[17]), .Y(n173) );
  NAND2X1 U187 ( .A(B[17]), .B(A[17]), .Y(n174) );
  XOR2X1 U188 ( .A(n1), .B(n22), .Y(SUM[16]) );
  OAI21X1 U189 ( .A(n176), .B(n1), .C(n177), .Y(n175) );
  NAND2X1 U190 ( .A(n177), .B(n297), .Y(n22) );
  INVX2 U191 ( .A(n176), .Y(n297) );
  NOR2X1 U192 ( .A(B[16]), .B(A[16]), .Y(n176) );
  NAND2X1 U193 ( .A(B[16]), .B(A[16]), .Y(n177) );
  XNOR2X1 U194 ( .A(n187), .B(n23), .Y(SUM[15]) );
  AOI21X1 U195 ( .A(n247), .B(n179), .C(n180), .Y(n178) );
  NOR2X1 U196 ( .A(n181), .B(n219), .Y(n179) );
  OAI21X1 U197 ( .A(n181), .B(n220), .C(n182), .Y(n180) );
  NAND2X1 U198 ( .A(n183), .B(n203), .Y(n181) );
  AOI21X1 U199 ( .A(n204), .B(n183), .C(n184), .Y(n182) );
  NOR2X1 U200 ( .A(n185), .B(n194), .Y(n183) );
  OAI21X1 U201 ( .A(n195), .B(n185), .C(n186), .Y(n184) );
  NAND2X1 U202 ( .A(n186), .B(n298), .Y(n23) );
  INVX2 U203 ( .A(n185), .Y(n298) );
  NOR2X1 U204 ( .A(B[15]), .B(A[15]), .Y(n185) );
  NAND2X1 U205 ( .A(B[15]), .B(A[15]), .Y(n186) );
  XNOR2X1 U206 ( .A(n196), .B(n24), .Y(SUM[14]) );
  OAI21X1 U207 ( .A(n188), .B(n246), .C(n189), .Y(n187) );
  NAND2X1 U208 ( .A(n217), .B(n190), .Y(n188) );
  AOI21X1 U209 ( .A(n218), .B(n190), .C(n191), .Y(n189) );
  NOR2X1 U210 ( .A(n194), .B(n201), .Y(n190) );
  OAI21X1 U211 ( .A(n194), .B(n202), .C(n195), .Y(n191) );
  NAND2X1 U214 ( .A(n195), .B(n193), .Y(n24) );
  NOR2X1 U216 ( .A(B[14]), .B(A[14]), .Y(n194) );
  NAND2X1 U217 ( .A(B[14]), .B(A[14]), .Y(n195) );
  XNOR2X1 U218 ( .A(n207), .B(n25), .Y(SUM[13]) );
  OAI21X1 U219 ( .A(n197), .B(n246), .C(n198), .Y(n196) );
  NAND2X1 U220 ( .A(n199), .B(n217), .Y(n197) );
  AOI21X1 U221 ( .A(n199), .B(n218), .C(n204), .Y(n198) );
  NOR2X1 U226 ( .A(n205), .B(n212), .Y(n203) );
  OAI21X1 U227 ( .A(n213), .B(n205), .C(n206), .Y(n204) );
  NAND2X1 U228 ( .A(n206), .B(n300), .Y(n25) );
  INVX2 U229 ( .A(n205), .Y(n300) );
  NOR2X1 U230 ( .A(B[13]), .B(A[13]), .Y(n205) );
  NAND2X1 U231 ( .A(B[13]), .B(A[13]), .Y(n206) );
  XNOR2X1 U232 ( .A(n214), .B(n26), .Y(SUM[12]) );
  OAI21X1 U233 ( .A(n208), .B(n246), .C(n209), .Y(n207) );
  NAND2X1 U234 ( .A(n210), .B(n217), .Y(n208) );
  AOI21X1 U235 ( .A(n210), .B(n218), .C(n211), .Y(n209) );
  NAND2X1 U238 ( .A(n213), .B(n210), .Y(n26) );
  NOR2X1 U240 ( .A(B[12]), .B(A[12]), .Y(n212) );
  NAND2X1 U241 ( .A(B[12]), .B(A[12]), .Y(n213) );
  XNOR2X1 U242 ( .A(n225), .B(n27), .Y(SUM[11]) );
  OAI21X1 U243 ( .A(n219), .B(n246), .C(n220), .Y(n214) );
  NAND2X1 U248 ( .A(n221), .B(n239), .Y(n219) );
  AOI21X1 U249 ( .A(n240), .B(n221), .C(n222), .Y(n220) );
  NOR2X1 U250 ( .A(n223), .B(n230), .Y(n221) );
  OAI21X1 U251 ( .A(n231), .B(n223), .C(n224), .Y(n222) );
  NAND2X1 U252 ( .A(n224), .B(n302), .Y(n27) );
  INVX2 U253 ( .A(n223), .Y(n302) );
  NOR2X1 U254 ( .A(B[11]), .B(A[11]), .Y(n223) );
  NAND2X1 U255 ( .A(B[11]), .B(A[11]), .Y(n224) );
  XNOR2X1 U256 ( .A(n232), .B(n28), .Y(SUM[10]) );
  OAI21X1 U257 ( .A(n226), .B(n246), .C(n227), .Y(n225) );
  NAND2X1 U258 ( .A(n228), .B(n239), .Y(n226) );
  AOI21X1 U259 ( .A(n228), .B(n240), .C(n229), .Y(n227) );
  NAND2X1 U262 ( .A(n231), .B(n228), .Y(n28) );
  NOR2X1 U264 ( .A(B[10]), .B(A[10]), .Y(n230) );
  NAND2X1 U265 ( .A(B[10]), .B(A[10]), .Y(n231) );
  XNOR2X1 U266 ( .A(n243), .B(n29), .Y(SUM[9]) );
  OAI21X1 U267 ( .A(n233), .B(n246), .C(n238), .Y(n232) );
  NOR2X1 U274 ( .A(n241), .B(n244), .Y(n239) );
  OAI21X1 U275 ( .A(n245), .B(n241), .C(n242), .Y(n240) );
  NAND2X1 U276 ( .A(n242), .B(n304), .Y(n29) );
  INVX2 U277 ( .A(n241), .Y(n304) );
  NOR2X1 U278 ( .A(B[9]), .B(A[9]), .Y(n241) );
  NAND2X1 U279 ( .A(B[9]), .B(A[9]), .Y(n242) );
  XOR2X1 U280 ( .A(n246), .B(n30), .Y(SUM[8]) );
  OAI21X1 U281 ( .A(n244), .B(n246), .C(n245), .Y(n243) );
  NAND2X1 U282 ( .A(n245), .B(n305), .Y(n30) );
  INVX2 U283 ( .A(n244), .Y(n305) );
  NOR2X1 U284 ( .A(B[8]), .B(A[8]), .Y(n244) );
  NAND2X1 U285 ( .A(B[8]), .B(A[8]), .Y(n245) );
  XNOR2X1 U286 ( .A(n254), .B(n31), .Y(SUM[7]) );
  OAI21X1 U288 ( .A(n248), .B(n268), .C(n249), .Y(n247) );
  NAND2X1 U289 ( .A(n250), .B(n258), .Y(n248) );
  AOI21X1 U290 ( .A(n259), .B(n250), .C(n251), .Y(n249) );
  NOR2X1 U291 ( .A(n252), .B(n255), .Y(n250) );
  OAI21X1 U292 ( .A(n256), .B(n252), .C(n253), .Y(n251) );
  NAND2X1 U293 ( .A(n253), .B(n306), .Y(n31) );
  INVX2 U294 ( .A(n252), .Y(n306) );
  NOR2X1 U295 ( .A(B[7]), .B(A[7]), .Y(n252) );
  NAND2X1 U296 ( .A(B[7]), .B(A[7]), .Y(n253) );
  XOR2X1 U297 ( .A(n257), .B(n32), .Y(SUM[6]) );
  OAI21X1 U298 ( .A(n255), .B(n257), .C(n256), .Y(n254) );
  NAND2X1 U299 ( .A(n256), .B(n307), .Y(n32) );
  INVX2 U300 ( .A(n255), .Y(n307) );
  NOR2X1 U301 ( .A(B[6]), .B(A[6]), .Y(n255) );
  NAND2X1 U302 ( .A(B[6]), .B(A[6]), .Y(n256) );
  XOR2X1 U303 ( .A(n262), .B(n33), .Y(SUM[5]) );
  AOI21X1 U304 ( .A(n258), .B(n267), .C(n259), .Y(n257) );
  NOR2X1 U305 ( .A(n260), .B(n265), .Y(n258) );
  OAI21X1 U306 ( .A(n266), .B(n260), .C(n261), .Y(n259) );
  NAND2X1 U307 ( .A(n261), .B(n308), .Y(n33) );
  INVX2 U308 ( .A(n260), .Y(n308) );
  NOR2X1 U309 ( .A(B[5]), .B(A[5]), .Y(n260) );
  NAND2X1 U310 ( .A(B[5]), .B(A[5]), .Y(n261) );
  XNOR2X1 U311 ( .A(n267), .B(n34), .Y(SUM[4]) );
  AOI21X1 U312 ( .A(n263), .B(n267), .C(n264), .Y(n262) );
  NAND2X1 U315 ( .A(n266), .B(n263), .Y(n34) );
  NOR2X1 U317 ( .A(B[4]), .B(A[4]), .Y(n265) );
  NAND2X1 U318 ( .A(B[4]), .B(A[4]), .Y(n266) );
  XNOR2X1 U319 ( .A(n273), .B(n35), .Y(SUM[3]) );
  AOI21X1 U321 ( .A(n277), .B(n269), .C(n270), .Y(n268) );
  NOR2X1 U322 ( .A(n271), .B(n274), .Y(n269) );
  OAI21X1 U323 ( .A(n275), .B(n271), .C(n272), .Y(n270) );
  NAND2X1 U324 ( .A(n272), .B(n310), .Y(n35) );
  INVX2 U325 ( .A(n271), .Y(n310) );
  NOR2X1 U326 ( .A(B[3]), .B(A[3]), .Y(n271) );
  NAND2X1 U327 ( .A(B[3]), .B(A[3]), .Y(n272) );
  XOR2X1 U328 ( .A(n276), .B(n36), .Y(SUM[2]) );
  OAI21X1 U329 ( .A(n274), .B(n276), .C(n275), .Y(n273) );
  NAND2X1 U330 ( .A(n275), .B(n311), .Y(n36) );
  INVX2 U331 ( .A(n274), .Y(n311) );
  NOR2X1 U332 ( .A(B[2]), .B(A[2]), .Y(n274) );
  NAND2X1 U333 ( .A(B[2]), .B(A[2]), .Y(n275) );
  XOR2X1 U334 ( .A(n37), .B(n281), .Y(SUM[1]) );
  OAI21X1 U336 ( .A(n281), .B(n278), .C(n279), .Y(n277) );
  NAND2X1 U337 ( .A(n279), .B(n312), .Y(n37) );
  INVX2 U338 ( .A(n278), .Y(n312) );
  NOR2X1 U339 ( .A(B[1]), .B(A[1]), .Y(n278) );
  NAND2X1 U340 ( .A(B[1]), .B(A[1]), .Y(n279) );
  NAND2X1 U345 ( .A(B[0]), .B(A[0]), .Y(n281) );
  OR2X2 U349 ( .A(B[30]), .B(A[30]), .Y(n417) );
  OR2X2 U350 ( .A(B[0]), .B(A[0]), .Y(n418) );
  INVX1 U351 ( .A(n79), .Y(n286) );
  INVX1 U352 ( .A(n247), .Y(n246) );
  INVX1 U353 ( .A(n4), .Y(n109) );
  INVX1 U354 ( .A(n171), .Y(n165) );
  INVX1 U355 ( .A(n239), .Y(n233) );
  INVX1 U356 ( .A(n268), .Y(n267) );
  INVX1 U357 ( .A(n277), .Y(n276) );
  INVX1 U358 ( .A(n69), .Y(n68) );
  INVX1 U359 ( .A(n87), .Y(n86) );
  OR2X1 U360 ( .A(B[31]), .B(A[31]), .Y(n420) );
  BUFX2 U361 ( .A(n178), .Y(n1) );
  BUFX2 U362 ( .A(n178), .Y(n2) );
  INVX1 U363 ( .A(n219), .Y(n217) );
  BUFX2 U364 ( .A(n111), .Y(n4) );
  INVX1 U365 ( .A(n150), .Y(n148) );
  INVX1 U366 ( .A(n95), .Y(n93) );
  INVX1 U367 ( .A(n133), .Y(n131) );
  INVX1 U368 ( .A(n201), .Y(n199) );
  INVX1 U369 ( .A(n220), .Y(n218) );
  INVX1 U370 ( .A(n136), .Y(n134) );
  INVX1 U371 ( .A(n204), .Y(n202) );
  INVX1 U372 ( .A(n240), .Y(n238) );
  INVX2 U373 ( .A(n170), .Y(n168) );
  INVX1 U374 ( .A(n145), .Y(n143) );
  INVX1 U375 ( .A(n230), .Y(n228) );
  INVX1 U376 ( .A(n106), .Y(n104) );
  INVX1 U377 ( .A(n162), .Y(n160) );
  INVX1 U378 ( .A(n51), .Y(n49) );
  INVX1 U379 ( .A(n265), .Y(n263) );
  INVX1 U380 ( .A(n107), .Y(n105) );
  INVX1 U381 ( .A(n213), .Y(n211) );
  INVX1 U382 ( .A(n266), .Y(n264) );
  INVX1 U383 ( .A(n163), .Y(n161) );
  INVX1 U384 ( .A(n231), .Y(n229) );
  INVX1 U385 ( .A(n125), .Y(n124) );
  INVX1 U386 ( .A(n70), .Y(n69) );
  INVX1 U387 ( .A(n88), .Y(n87) );
  INVX1 U388 ( .A(n194), .Y(n193) );
  AND2X1 U389 ( .A(n281), .B(n418), .Y(SUM[0]) );
  INVX1 U390 ( .A(n212), .Y(n210) );
  INVX1 U391 ( .A(n203), .Y(n201) );
  INVX1 U392 ( .A(n3), .Y(n110) );
  INVX1 U393 ( .A(n126), .Y(n125) );
  INVX1 U394 ( .A(n99), .Y(n288) );
  INVX1 U395 ( .A(n97), .Y(n95) );
  INVX1 U396 ( .A(n144), .Y(n142) );
  INVX1 U397 ( .A(n135), .Y(n133) );
  INVX1 U398 ( .A(n5), .Y(n76) );
  INVX1 U399 ( .A(n98), .Y(n96) );
  INVX1 U400 ( .A(n6), .Y(n75) );
  INVX1 U401 ( .A(n60), .Y(n58) );
  INVX1 U402 ( .A(n151), .Y(n149) );
  INVX1 U403 ( .A(n61), .Y(n284) );
  INVX1 U404 ( .A(n59), .Y(n57) );
  INVX1 U405 ( .A(n117), .Y(n290) );
  BUFX4 U406 ( .A(n112), .Y(n3) );
  INVX1 U407 ( .A(n152), .Y(n150) );
  INVX1 U408 ( .A(n172), .Y(n170) );
endmodule


module poly5_DW_mult_uns_44 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n8, n13, n18, n23, n28, n33, n38, n68, n80, n85, n89, n98, n107, n116,
         n125, n134, n143, n152, n163, n168, n178, n179, n194, n195, n201,
         n211, n216, n226, n227, n242, n243, n249, n258, n259, n275, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n439, n441, n453, n459, n461, n463, n465, n467, n469,
         n471, n473, n475, n477, n479, n481, n483, n485, n487, n489, n491,
         n493, n495, n497, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n548, n549, n551, n553, n554, n555,
         n557, n559, n560, n561, n562, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n624, n625, n626, n627, n628, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n704, n706, n707, n709, n711,
         n712, n713, n714, n716, n718, n719, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n757, n759, n760, n761, n764,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n799,
         n801, n802, n803, n804, n805, n806, n807, n808, n810, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n830, n832, n833, n834, n835, n836, n838,
         n840, n841, n843, n846, n848, n850, n851, n852, n853, n854, n856,
         n858, n859, n860, n861, n862, n867, n868, n869, n870, n872, n876,
         n878, n879, n883, n884, n885, n886, n888, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2248, n2250, n2251,
         n2252, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000;

  NAND2X1 OR_NOTi ( .A(n2999), .B(n289), .Y(n2725) );
  INVX2 U21 ( .A(n387), .Y(n275) );
  OAI21X1 AO21i ( .A(a[0]), .B(n275), .C(n289), .Y(n2206) );
  NAND2X1 OR_NOTi1 ( .A(n3000), .B(n292), .Y(n2692) );
  INVX2 U23 ( .A(n390), .Y(n259) );
  INVX2 U15 ( .A(n340), .Y(n258) );
  OAI21X1 AO21i1 ( .A(n258), .B(n259), .C(n292), .Y(n2172) );
  NAND2X1 OR_NOTi2 ( .A(n2999), .B(n295), .Y(n2659) );
  INVX2 U24 ( .A(n249), .Y(n2171) );
  NAND2X1 AND_NOTi2 ( .A(n2913), .B(n242), .Y(n249) );
  INVX2 U25 ( .A(n393), .Y(n243) );
  INVX2 U18 ( .A(n343), .Y(n242) );
  OAI21X1 AO21i2 ( .A(n242), .B(n243), .C(n295), .Y(n2138) );
  NAND2X1 OR_NOTi3 ( .A(n2999), .B(n298), .Y(n2626) );
  INVX2 U27 ( .A(n396), .Y(n227) );
  INVX2 U111 ( .A(n346), .Y(n226) );
  OAI21X1 AO21i3 ( .A(n226), .B(n227), .C(n297), .Y(n2104) );
  NAND2X1 OR_NOTi4 ( .A(n3000), .B(n301), .Y(n2593) );
  INVX2 U113 ( .A(n349), .Y(n216) );
  INVX2 U29 ( .A(n399), .Y(n211) );
  OAI21X1 AO21i4 ( .A(n216), .B(n211), .C(n300), .Y(n2070) );
  NAND2X1 OR_NOTi5 ( .A(n2999), .B(n304), .Y(n2560) );
  INVX2 U210 ( .A(n201), .Y(n2069) );
  NAND2X1 AND_NOTi5 ( .A(n2913), .B(n194), .Y(n201) );
  INVX2 U211 ( .A(n402), .Y(n195) );
  INVX2 U117 ( .A(n352), .Y(n194) );
  OAI21X1 AO21i5 ( .A(n194), .B(n195), .C(n303), .Y(n2036) );
  NAND2X1 OR_NOTi6 ( .A(n3000), .B(n307), .Y(n2527) );
  INVX2 U213 ( .A(n405), .Y(n179) );
  INVX2 U120 ( .A(n355), .Y(n178) );
  OAI21X1 AO21i6 ( .A(n178), .B(n179), .C(n306), .Y(n2002) );
  NAND2X1 OR_NOTi7 ( .A(n3000), .B(n310), .Y(n2494) );
  INVX2 U122 ( .A(n358), .Y(n168) );
  INVX2 U215 ( .A(n408), .Y(n163) );
  OAI21X1 AO21i7 ( .A(n168), .B(n163), .C(n309), .Y(n1968) );
  NAND2X1 OR_NOTi8 ( .A(n3000), .B(n313), .Y(n2461) );
  INVX2 U125 ( .A(n361), .Y(n152) );
  NAND2X1 OR_NOTi9 ( .A(n3000), .B(n316), .Y(n2428) );
  INVX2 U127 ( .A(n364), .Y(n143) );
  NAND2X1 OR_NOTi10 ( .A(n3000), .B(n319), .Y(n2397) );
  INVX2 U129 ( .A(n367), .Y(n134) );
  NAND2X1 OR_NOTi11 ( .A(n3000), .B(n322), .Y(n2368) );
  INVX2 U131 ( .A(n370), .Y(n125) );
  NAND2X1 OR_NOTi12 ( .A(n3000), .B(n325), .Y(n2341) );
  INVX2 U133 ( .A(n373), .Y(n116) );
  NAND2X1 OR_NOTi13 ( .A(n3000), .B(n328), .Y(n2316) );
  INVX2 U135 ( .A(n376), .Y(n107) );
  NAND2X1 OR_NOTi14 ( .A(n3000), .B(n331), .Y(n2293) );
  INVX2 U137 ( .A(n379), .Y(n98) );
  NAND2X1 OR_NOTi15 ( .A(n3000), .B(n334), .Y(n2272) );
  INVX2 U139 ( .A(n382), .Y(n89) );
  INVX2 U224 ( .A(n85), .Y(n1767) );
  NAND2X1 AND_NOTi16 ( .A(n2944), .B(n333), .Y(n85) );
  XOR2X1 U225 ( .A(n1759), .B(n918), .Y(n80) );
  XOR2X1 U141 ( .A(n1852), .B(n80), .Y(n899) );
  XOR2X1 U226 ( .A(n1768), .B(n1828), .Y(n68) );
  XOR2X1 U142 ( .A(n1786), .B(n68), .Y(n898) );
  XOR2X1 U227 ( .A(n1906), .B(n1806), .Y(n38) );
  XOR2X1 U143 ( .A(n1878), .B(n38), .Y(n897) );
  XOR2X1 U228 ( .A(n1968), .B(n1936), .Y(n33) );
  XOR2X1 U144 ( .A(n899), .B(n33), .Y(n896) );
  XOR2X1 U229 ( .A(n914), .B(n916), .Y(n28) );
  XOR2X1 U145 ( .A(n912), .B(n28), .Y(n895) );
  XOR2X1 U230 ( .A(n898), .B(n897), .Y(n23) );
  XOR2X1 U146 ( .A(n910), .B(n23), .Y(n894) );
  XOR2X1 U231 ( .A(n908), .B(n896), .Y(n18) );
  XOR2X1 U147 ( .A(n895), .B(n18), .Y(n893) );
  XOR2X1 U232 ( .A(n894), .B(n906), .Y(n13) );
  XOR2X1 U148 ( .A(n904), .B(n13), .Y(n892) );
  XOR2X1 U233 ( .A(n902), .B(n893), .Y(n8) );
  XOR2X1 U149 ( .A(n892), .B(n8), .Y(n891) );
  XNOR2X1 U292 ( .A(n549), .B(n500), .Y(product[47]) );
  NAND2X1 U293 ( .A(n548), .B(n2931), .Y(n500) );
  NAND2X1 U296 ( .A(n900), .B(n891), .Y(n548) );
  XNOR2X1 U297 ( .A(n560), .B(n501), .Y(product[46]) );
  OAI21X1 U298 ( .A(n2946), .B(n499), .C(n551), .Y(n549) );
  OAI21X1 U302 ( .A(n554), .B(n582), .C(n555), .Y(n553) );
  NAND2X1 U303 ( .A(n2925), .B(n565), .Y(n554) );
  AOI21X1 U304 ( .A(n2925), .B(n566), .C(n557), .Y(n555) );
  NAND2X1 U307 ( .A(n559), .B(n2925), .Y(n501) );
  NAND2X1 U310 ( .A(n920), .B(n901), .Y(n559) );
  XNOR2X1 U311 ( .A(n569), .B(n502), .Y(product[45]) );
  OAI21X1 U312 ( .A(n561), .B(n499), .C(n562), .Y(n560) );
  NAND2X1 U313 ( .A(n565), .B(n579), .Y(n561) );
  AOI21X1 U314 ( .A(n565), .B(n580), .C(n566), .Y(n562) );
  NOR2X1 U317 ( .A(n567), .B(n574), .Y(n565) );
  OAI21X1 U318 ( .A(n567), .B(n575), .C(n568), .Y(n566) );
  NAND2X1 U319 ( .A(n568), .B(n846), .Y(n502) );
  INVX2 U320 ( .A(n567), .Y(n846) );
  NOR2X1 U321 ( .A(n921), .B(n940), .Y(n567) );
  NAND2X1 U322 ( .A(n921), .B(n940), .Y(n568) );
  XNOR2X1 U323 ( .A(n576), .B(n503), .Y(product[44]) );
  OAI21X1 U324 ( .A(n570), .B(n499), .C(n571), .Y(n569) );
  NAND2X1 U325 ( .A(n572), .B(n579), .Y(n570) );
  AOI21X1 U326 ( .A(n572), .B(n580), .C(n573), .Y(n571) );
  NAND2X1 U329 ( .A(n575), .B(n572), .Y(n503) );
  NOR2X1 U331 ( .A(n962), .B(n941), .Y(n574) );
  NAND2X1 U332 ( .A(n962), .B(n941), .Y(n575) );
  XNOR2X1 U333 ( .A(n587), .B(n504), .Y(product[43]) );
  OAI21X1 U334 ( .A(n581), .B(n499), .C(n582), .Y(n576) );
  NAND2X1 U339 ( .A(n583), .B(n601), .Y(n581) );
  AOI21X1 U340 ( .A(n583), .B(n602), .C(n584), .Y(n582) );
  NOR2X1 U341 ( .A(n585), .B(n592), .Y(n583) );
  OAI21X1 U342 ( .A(n593), .B(n585), .C(n586), .Y(n584) );
  NAND2X1 U343 ( .A(n586), .B(n848), .Y(n504) );
  INVX2 U344 ( .A(n585), .Y(n848) );
  NOR2X1 U345 ( .A(n984), .B(n963), .Y(n585) );
  NAND2X1 U346 ( .A(n984), .B(n963), .Y(n586) );
  XNOR2X1 U347 ( .A(n594), .B(n505), .Y(product[42]) );
  OAI21X1 U348 ( .A(n588), .B(n499), .C(n589), .Y(n587) );
  NAND2X1 U349 ( .A(n590), .B(n601), .Y(n588) );
  AOI21X1 U350 ( .A(n590), .B(n602), .C(n591), .Y(n589) );
  NAND2X1 U353 ( .A(n593), .B(n590), .Y(n505) );
  NOR2X1 U355 ( .A(n1008), .B(n985), .Y(n592) );
  NAND2X1 U356 ( .A(n1008), .B(n985), .Y(n593) );
  XNOR2X1 U357 ( .A(n605), .B(n506), .Y(product[41]) );
  OAI21X1 U358 ( .A(n595), .B(n499), .C(n600), .Y(n594) );
  NOR2X1 U365 ( .A(n603), .B(n606), .Y(n601) );
  OAI21X1 U366 ( .A(n607), .B(n603), .C(n604), .Y(n602) );
  NAND2X1 U367 ( .A(n604), .B(n850), .Y(n506) );
  INVX2 U368 ( .A(n603), .Y(n850) );
  NOR2X1 U369 ( .A(n1032), .B(n1009), .Y(n603) );
  NAND2X1 U370 ( .A(n1032), .B(n1009), .Y(n604) );
  XOR2X1 U371 ( .A(n499), .B(n507), .Y(product[40]) );
  OAI21X1 U372 ( .A(n606), .B(n499), .C(n607), .Y(n605) );
  NAND2X1 U373 ( .A(n607), .B(n851), .Y(n507) );
  INVX2 U374 ( .A(n606), .Y(n851) );
  NOR2X1 U375 ( .A(n1058), .B(n1033), .Y(n606) );
  NAND2X1 U376 ( .A(n1058), .B(n1033), .Y(n607) );
  XNOR2X1 U377 ( .A(n617), .B(n508), .Y(product[39]) );
  AOI21X1 U378 ( .A(n677), .B(n609), .C(n610), .Y(n608) );
  NOR2X1 U379 ( .A(n649), .B(n611), .Y(n609) );
  OAI21X1 U380 ( .A(n611), .B(n650), .C(n612), .Y(n610) );
  NAND2X1 U381 ( .A(n613), .B(n633), .Y(n611) );
  AOI21X1 U382 ( .A(n634), .B(n613), .C(n614), .Y(n612) );
  NOR2X1 U383 ( .A(n615), .B(n624), .Y(n613) );
  OAI21X1 U384 ( .A(n625), .B(n615), .C(n616), .Y(n614) );
  NAND2X1 U385 ( .A(n616), .B(n852), .Y(n508) );
  INVX2 U386 ( .A(n615), .Y(n852) );
  NOR2X1 U387 ( .A(n1084), .B(n1059), .Y(n615) );
  NAND2X1 U388 ( .A(n1084), .B(n1059), .Y(n616) );
  XNOR2X1 U389 ( .A(n626), .B(n509), .Y(product[38]) );
  OAI21X1 U390 ( .A(n676), .B(n618), .C(n619), .Y(n617) );
  NAND2X1 U391 ( .A(n647), .B(n620), .Y(n618) );
  AOI21X1 U392 ( .A(n648), .B(n620), .C(n621), .Y(n619) );
  NOR2X1 U393 ( .A(n624), .B(n631), .Y(n620) );
  OAI21X1 U394 ( .A(n624), .B(n632), .C(n625), .Y(n621) );
  NAND2X1 U397 ( .A(n625), .B(n853), .Y(n509) );
  INVX2 U398 ( .A(n624), .Y(n853) );
  NOR2X1 U399 ( .A(n1112), .B(n1085), .Y(n624) );
  NAND2X1 U400 ( .A(n1112), .B(n1085), .Y(n625) );
  XNOR2X1 U401 ( .A(n637), .B(n510), .Y(product[37]) );
  OAI21X1 U402 ( .A(n676), .B(n627), .C(n628), .Y(n626) );
  NAND2X1 U403 ( .A(n633), .B(n647), .Y(n627) );
  AOI21X1 U404 ( .A(n633), .B(n648), .C(n634), .Y(n628) );
  NOR2X1 U409 ( .A(n635), .B(n642), .Y(n633) );
  OAI21X1 U410 ( .A(n643), .B(n635), .C(n636), .Y(n634) );
  NAND2X1 U411 ( .A(n636), .B(n854), .Y(n510) );
  INVX2 U412 ( .A(n635), .Y(n854) );
  NOR2X1 U413 ( .A(n1140), .B(n1113), .Y(n635) );
  NAND2X1 U414 ( .A(n1140), .B(n1113), .Y(n636) );
  XNOR2X1 U415 ( .A(n644), .B(n511), .Y(product[36]) );
  OAI21X1 U416 ( .A(n676), .B(n638), .C(n639), .Y(n637) );
  NAND2X1 U417 ( .A(n640), .B(n647), .Y(n638) );
  AOI21X1 U418 ( .A(n640), .B(n648), .C(n641), .Y(n639) );
  NAND2X1 U421 ( .A(n643), .B(n640), .Y(n511) );
  NOR2X1 U423 ( .A(n1170), .B(n1141), .Y(n642) );
  NAND2X1 U424 ( .A(n1170), .B(n1141), .Y(n643) );
  XNOR2X1 U425 ( .A(n655), .B(n512), .Y(product[35]) );
  OAI21X1 U426 ( .A(n649), .B(n676), .C(n650), .Y(n644) );
  NAND2X1 U431 ( .A(n669), .B(n651), .Y(n649) );
  AOI21X1 U432 ( .A(n670), .B(n651), .C(n652), .Y(n650) );
  NOR2X1 U433 ( .A(n653), .B(n660), .Y(n651) );
  OAI21X1 U434 ( .A(n661), .B(n653), .C(n654), .Y(n652) );
  NAND2X1 U435 ( .A(n654), .B(n856), .Y(n512) );
  INVX2 U436 ( .A(n653), .Y(n856) );
  NOR2X1 U437 ( .A(n1200), .B(n1171), .Y(n653) );
  NAND2X1 U438 ( .A(n1200), .B(n1171), .Y(n654) );
  XNOR2X1 U439 ( .A(n662), .B(n513), .Y(product[34]) );
  OAI21X1 U440 ( .A(n656), .B(n676), .C(n657), .Y(n655) );
  NAND2X1 U441 ( .A(n658), .B(n669), .Y(n656) );
  AOI21X1 U442 ( .A(n658), .B(n670), .C(n659), .Y(n657) );
  NAND2X1 U445 ( .A(n661), .B(n658), .Y(n513) );
  NOR2X1 U447 ( .A(n1232), .B(n1201), .Y(n660) );
  NAND2X1 U448 ( .A(n1232), .B(n1201), .Y(n661) );
  XNOR2X1 U449 ( .A(n673), .B(n514), .Y(product[33]) );
  OAI21X1 U450 ( .A(n663), .B(n676), .C(n668), .Y(n662) );
  NOR2X1 U457 ( .A(n674), .B(n671), .Y(n669) );
  OAI21X1 U458 ( .A(n675), .B(n671), .C(n672), .Y(n670) );
  NAND2X1 U459 ( .A(n672), .B(n858), .Y(n514) );
  INVX2 U460 ( .A(n671), .Y(n858) );
  NOR2X1 U461 ( .A(n1263), .B(n1233), .Y(n671) );
  NAND2X1 U462 ( .A(n1263), .B(n1233), .Y(n672) );
  XOR2X1 U463 ( .A(n676), .B(n515), .Y(product[32]) );
  OAI21X1 U464 ( .A(n674), .B(n676), .C(n675), .Y(n673) );
  NAND2X1 U465 ( .A(n675), .B(n859), .Y(n515) );
  INVX2 U466 ( .A(n674), .Y(n859) );
  NOR2X1 U467 ( .A(n1293), .B(n1264), .Y(n674) );
  NAND2X1 U468 ( .A(n1293), .B(n1264), .Y(n675) );
  XNOR2X1 U469 ( .A(n684), .B(n516), .Y(product[31]) );
  OAI21X1 U471 ( .A(n698), .B(n678), .C(n679), .Y(n677) );
  NAND2X1 U472 ( .A(n688), .B(n680), .Y(n678) );
  AOI21X1 U473 ( .A(n689), .B(n680), .C(n681), .Y(n679) );
  NOR2X1 U474 ( .A(n685), .B(n682), .Y(n680) );
  OAI21X1 U475 ( .A(n686), .B(n682), .C(n683), .Y(n681) );
  NAND2X1 U476 ( .A(n683), .B(n860), .Y(n516) );
  INVX2 U477 ( .A(n682), .Y(n860) );
  NOR2X1 U478 ( .A(n1323), .B(n1294), .Y(n682) );
  NAND2X1 U479 ( .A(n1323), .B(n1294), .Y(n683) );
  XOR2X1 U480 ( .A(n687), .B(n517), .Y(product[30]) );
  OAI21X1 U481 ( .A(n685), .B(n687), .C(n686), .Y(n684) );
  NAND2X1 U482 ( .A(n686), .B(n861), .Y(n517) );
  INVX2 U483 ( .A(n685), .Y(n861) );
  NOR2X1 U484 ( .A(n1351), .B(n1324), .Y(n685) );
  NAND2X1 U485 ( .A(n1351), .B(n1324), .Y(n686) );
  XOR2X1 U486 ( .A(n692), .B(n518), .Y(product[29]) );
  AOI21X1 U487 ( .A(n688), .B(n697), .C(n689), .Y(n687) );
  NOR2X1 U488 ( .A(n695), .B(n690), .Y(n688) );
  OAI21X1 U489 ( .A(n696), .B(n690), .C(n691), .Y(n689) );
  NAND2X1 U490 ( .A(n691), .B(n862), .Y(n518) );
  INVX2 U491 ( .A(n690), .Y(n862) );
  NOR2X1 U492 ( .A(n1379), .B(n1352), .Y(n690) );
  NAND2X1 U493 ( .A(n1379), .B(n1352), .Y(n691) );
  XNOR2X1 U494 ( .A(n697), .B(n519), .Y(product[28]) );
  AOI21X1 U495 ( .A(n693), .B(n697), .C(n694), .Y(n692) );
  NAND2X1 U498 ( .A(n696), .B(n693), .Y(n519) );
  NOR2X1 U500 ( .A(n1405), .B(n1380), .Y(n695) );
  NAND2X1 U501 ( .A(n1405), .B(n1380), .Y(n696) );
  XOR2X1 U502 ( .A(n707), .B(n520), .Y(product[27]) );
  AOI21X1 U504 ( .A(n699), .B(n727), .C(n700), .Y(n698) );
  NOR2X1 U505 ( .A(n713), .B(n701), .Y(n699) );
  OAI21X1 U506 ( .A(n714), .B(n701), .C(n702), .Y(n700) );
  NAND2X1 U507 ( .A(n2924), .B(n2917), .Y(n701) );
  AOI21X1 U508 ( .A(n709), .B(n2917), .C(n704), .Y(n702) );
  NAND2X1 U511 ( .A(n706), .B(n2917), .Y(n520) );
  NAND2X1 U514 ( .A(n1431), .B(n1406), .Y(n706) );
  XNOR2X1 U515 ( .A(n712), .B(n521), .Y(product[26]) );
  AOI21X1 U516 ( .A(n2924), .B(n712), .C(n709), .Y(n707) );
  NAND2X1 U519 ( .A(n711), .B(n2924), .Y(n521) );
  NAND2X1 U522 ( .A(n1455), .B(n1432), .Y(n711) );
  XNOR2X1 U523 ( .A(n719), .B(n522), .Y(product[25]) );
  OAI21X1 U524 ( .A(n713), .B(n726), .C(n714), .Y(n712) );
  NAND2X1 U525 ( .A(n867), .B(n2923), .Y(n713) );
  AOI21X1 U526 ( .A(n723), .B(n2923), .C(n716), .Y(n714) );
  NAND2X1 U529 ( .A(n718), .B(n2923), .Y(n522) );
  NAND2X1 U532 ( .A(n1479), .B(n1456), .Y(n718) );
  XOR2X1 U533 ( .A(n726), .B(n523), .Y(product[24]) );
  OAI21X1 U534 ( .A(n724), .B(n726), .C(n725), .Y(n719) );
  NAND2X1 U539 ( .A(n725), .B(n867), .Y(n523) );
  INVX2 U540 ( .A(n724), .Y(n867) );
  NOR2X1 U541 ( .A(n1501), .B(n1480), .Y(n724) );
  NAND2X1 U542 ( .A(n1501), .B(n1480), .Y(n725) );
  XNOR2X1 U543 ( .A(n734), .B(n524), .Y(product[23]) );
  OAI21X1 U545 ( .A(n748), .B(n728), .C(n729), .Y(n727) );
  NAND2X1 U546 ( .A(n738), .B(n730), .Y(n728) );
  AOI21X1 U547 ( .A(n739), .B(n730), .C(n731), .Y(n729) );
  NOR2X1 U548 ( .A(n735), .B(n732), .Y(n730) );
  OAI21X1 U549 ( .A(n736), .B(n732), .C(n733), .Y(n731) );
  NAND2X1 U550 ( .A(n733), .B(n868), .Y(n524) );
  INVX2 U551 ( .A(n732), .Y(n868) );
  NOR2X1 U552 ( .A(n1523), .B(n1502), .Y(n732) );
  NAND2X1 U553 ( .A(n1523), .B(n1502), .Y(n733) );
  XOR2X1 U554 ( .A(n737), .B(n525), .Y(product[22]) );
  OAI21X1 U555 ( .A(n735), .B(n737), .C(n736), .Y(n734) );
  NAND2X1 U556 ( .A(n736), .B(n869), .Y(n525) );
  INVX2 U557 ( .A(n735), .Y(n869) );
  NOR2X1 U558 ( .A(n1543), .B(n1524), .Y(n735) );
  NAND2X1 U559 ( .A(n1543), .B(n1524), .Y(n736) );
  XOR2X1 U560 ( .A(n742), .B(n526), .Y(product[21]) );
  AOI21X1 U561 ( .A(n738), .B(n747), .C(n739), .Y(n737) );
  NOR2X1 U562 ( .A(n745), .B(n740), .Y(n738) );
  OAI21X1 U563 ( .A(n746), .B(n740), .C(n741), .Y(n739) );
  NAND2X1 U564 ( .A(n741), .B(n870), .Y(n526) );
  INVX2 U565 ( .A(n740), .Y(n870) );
  NOR2X1 U566 ( .A(n1563), .B(n1544), .Y(n740) );
  NAND2X1 U567 ( .A(n1563), .B(n1544), .Y(n741) );
  XNOR2X1 U568 ( .A(n747), .B(n527), .Y(product[20]) );
  AOI21X1 U569 ( .A(n743), .B(n747), .C(n744), .Y(n742) );
  NAND2X1 U572 ( .A(n746), .B(n743), .Y(n527) );
  NOR2X1 U574 ( .A(n1581), .B(n1564), .Y(n745) );
  NAND2X1 U575 ( .A(n1581), .B(n1564), .Y(n746) );
  XNOR2X1 U576 ( .A(n753), .B(n528), .Y(product[19]) );
  AOI21X1 U578 ( .A(n749), .B(n768), .C(n750), .Y(n748) );
  NOR2X1 U579 ( .A(n751), .B(n754), .Y(n749) );
  OAI21X1 U580 ( .A(n751), .B(n755), .C(n752), .Y(n750) );
  NAND2X1 U581 ( .A(n752), .B(n872), .Y(n528) );
  INVX2 U582 ( .A(n751), .Y(n872) );
  NOR2X1 U583 ( .A(n1599), .B(n1582), .Y(n751) );
  NAND2X1 U584 ( .A(n1599), .B(n1582), .Y(n752) );
  XNOR2X1 U585 ( .A(n760), .B(n529), .Y(product[18]) );
  OAI21X1 U586 ( .A(n754), .B(n767), .C(n755), .Y(n753) );
  NAND2X1 U587 ( .A(n2918), .B(n2916), .Y(n754) );
  AOI21X1 U588 ( .A(n764), .B(n2916), .C(n757), .Y(n755) );
  NAND2X1 U591 ( .A(n759), .B(n2916), .Y(n529) );
  NAND2X1 U594 ( .A(n1615), .B(n1600), .Y(n759) );
  XOR2X1 U595 ( .A(n767), .B(n530), .Y(product[17]) );
  OAI21X1 U596 ( .A(n761), .B(n767), .C(n766), .Y(n760) );
  NAND2X1 U601 ( .A(n766), .B(n2918), .Y(n530) );
  NAND2X1 U604 ( .A(n1631), .B(n1616), .Y(n766) );
  XOR2X1 U605 ( .A(n775), .B(n531), .Y(product[16]) );
  OAI21X1 U607 ( .A(n786), .B(n769), .C(n770), .Y(n768) );
  NAND2X1 U608 ( .A(n771), .B(n776), .Y(n769) );
  AOI21X1 U609 ( .A(n771), .B(n777), .C(n772), .Y(n770) );
  NAND2X1 U612 ( .A(n774), .B(n771), .Y(n531) );
  NOR2X1 U614 ( .A(n1645), .B(n1632), .Y(n773) );
  NAND2X1 U615 ( .A(n1645), .B(n1632), .Y(n774) );
  AOI21X1 U617 ( .A(n776), .B(n785), .C(n777), .Y(n775) );
  NOR2X1 U618 ( .A(n783), .B(n778), .Y(n776) );
  OAI21X1 U619 ( .A(n784), .B(n778), .C(n779), .Y(n777) );
  NOR2X1 U622 ( .A(n1659), .B(n1646), .Y(n778) );
  NAND2X1 U623 ( .A(n1659), .B(n1646), .Y(n779) );
  XNOR2X1 U624 ( .A(n785), .B(n533), .Y(product[14]) );
  AOI21X1 U625 ( .A(n781), .B(n785), .C(n782), .Y(n780) );
  NAND2X1 U628 ( .A(n784), .B(n781), .Y(n533) );
  NOR2X1 U630 ( .A(n1671), .B(n1660), .Y(n783) );
  NAND2X1 U631 ( .A(n1671), .B(n1660), .Y(n784) );
  XNOR2X1 U632 ( .A(n791), .B(n534), .Y(product[13]) );
  AOI21X1 U634 ( .A(n787), .B(n795), .C(n788), .Y(n786) );
  NOR2X1 U635 ( .A(n792), .B(n789), .Y(n787) );
  OAI21X1 U636 ( .A(n793), .B(n789), .C(n790), .Y(n788) );
  NAND2X1 U637 ( .A(n790), .B(n878), .Y(n534) );
  NOR2X1 U639 ( .A(n1683), .B(n1672), .Y(n789) );
  NAND2X1 U640 ( .A(n1683), .B(n1672), .Y(n790) );
  XOR2X1 U641 ( .A(n794), .B(n535), .Y(product[12]) );
  OAI21X1 U642 ( .A(n792), .B(n794), .C(n793), .Y(n791) );
  NAND2X1 U643 ( .A(n793), .B(n879), .Y(n535) );
  NOR2X1 U645 ( .A(n1693), .B(n1684), .Y(n792) );
  NAND2X1 U646 ( .A(n1684), .B(n1693), .Y(n793) );
  XOR2X1 U647 ( .A(n802), .B(n536), .Y(product[11]) );
  OAI21X1 U649 ( .A(n808), .B(n796), .C(n797), .Y(n795) );
  NAND2X1 U650 ( .A(n803), .B(n2921), .Y(n796) );
  AOI21X1 U651 ( .A(n804), .B(n2921), .C(n799), .Y(n797) );
  NAND2X1 U654 ( .A(n801), .B(n2921), .Y(n536) );
  NAND2X1 U657 ( .A(n1703), .B(n1694), .Y(n801) );
  XNOR2X1 U658 ( .A(n807), .B(n537), .Y(product[10]) );
  AOI21X1 U659 ( .A(n803), .B(n807), .C(n804), .Y(n802) );
  NAND2X1 U662 ( .A(n806), .B(n803), .Y(n537) );
  NOR2X1 U664 ( .A(n1704), .B(n1711), .Y(n805) );
  NAND2X1 U665 ( .A(n1711), .B(n1704), .Y(n806) );
  XNOR2X1 U666 ( .A(n813), .B(n538), .Y(product[9]) );
  AOI21X1 U668 ( .A(n2920), .B(n813), .C(n810), .Y(n808) );
  NAND2X1 U671 ( .A(n812), .B(n2920), .Y(n538) );
  NAND2X1 U674 ( .A(n1719), .B(n1712), .Y(n812) );
  XOR2X1 U675 ( .A(n816), .B(n539), .Y(product[8]) );
  OAI21X1 U676 ( .A(n814), .B(n816), .C(n815), .Y(n813) );
  NAND2X1 U677 ( .A(n815), .B(n883), .Y(n539) );
  INVX2 U678 ( .A(n814), .Y(n883) );
  NOR2X1 U679 ( .A(n1725), .B(n1720), .Y(n814) );
  NAND2X1 U680 ( .A(n1725), .B(n1720), .Y(n815) );
  XNOR2X1 U681 ( .A(n821), .B(n540), .Y(product[7]) );
  AOI21X1 U682 ( .A(n825), .B(n817), .C(n818), .Y(n816) );
  NOR2X1 U683 ( .A(n822), .B(n819), .Y(n817) );
  OAI21X1 U684 ( .A(n823), .B(n819), .C(n820), .Y(n818) );
  NAND2X1 U685 ( .A(n820), .B(n884), .Y(n540) );
  NOR2X1 U687 ( .A(n1731), .B(n1726), .Y(n819) );
  NAND2X1 U688 ( .A(n1731), .B(n1726), .Y(n820) );
  XOR2X1 U689 ( .A(n541), .B(n824), .Y(product[6]) );
  OAI21X1 U690 ( .A(n2990), .B(n824), .C(n2989), .Y(n821) );
  NAND2X1 U691 ( .A(n2989), .B(n885), .Y(n541) );
  NOR2X1 U693 ( .A(n1735), .B(n1732), .Y(n822) );
  NAND2X1 U694 ( .A(n1735), .B(n1732), .Y(n823) );
  XOR2X1 U695 ( .A(n542), .B(n828), .Y(product[5]) );
  OAI21X1 U697 ( .A(n826), .B(n828), .C(n827), .Y(n825) );
  NAND2X1 U698 ( .A(n827), .B(n886), .Y(n542) );
  INVX2 U699 ( .A(n826), .Y(n886) );
  NOR2X1 U700 ( .A(n1739), .B(n1736), .Y(n826) );
  NAND2X1 U701 ( .A(n1739), .B(n1736), .Y(n827) );
  XNOR2X1 U702 ( .A(n543), .B(n833), .Y(product[4]) );
  AOI21X1 U703 ( .A(n833), .B(n2919), .C(n830), .Y(n828) );
  NAND2X1 U706 ( .A(n832), .B(n2919), .Y(n543) );
  NAND2X1 U709 ( .A(n1741), .B(n1740), .Y(n832) );
  XOR2X1 U710 ( .A(n544), .B(n836), .Y(product[3]) );
  OAI21X1 U711 ( .A(n834), .B(n836), .C(n835), .Y(n833) );
  NAND2X1 U712 ( .A(n835), .B(n888), .Y(n544) );
  INVX2 U713 ( .A(n834), .Y(n888) );
  NOR2X1 U714 ( .A(n1757), .B(n1742), .Y(n834) );
  NAND2X1 U715 ( .A(n1757), .B(n1742), .Y(n835) );
  XNOR2X1 U716 ( .A(n545), .B(n841), .Y(product[2]) );
  AOI21X1 U717 ( .A(n841), .B(n2922), .C(n838), .Y(n836) );
  NAND2X1 U720 ( .A(n840), .B(n2922), .Y(n545) );
  NAND2X1 U723 ( .A(n2237), .B(n2954), .Y(n840) );
  NAND2X1 U729 ( .A(n1758), .B(n2238), .Y(n843) );
  FAX1 U730 ( .A(n905), .B(n922), .C(n903), .YC(n900), .YS(n901) );
  FAX1 U731 ( .A(n926), .B(n907), .C(n924), .YC(n902), .YS(n903) );
  FAX1 U732 ( .A(n911), .B(n928), .C(n909), .YC(n904), .YS(n905) );
  FAX1 U733 ( .A(n915), .B(n932), .C(n930), .YC(n906), .YS(n907) );
  FAX1 U734 ( .A(n934), .B(n917), .C(n913), .YC(n908), .YS(n909) );
  FAX1 U735 ( .A(n1829), .B(n938), .C(n936), .YC(n910), .YS(n911) );
  FAX1 U736 ( .A(n1853), .B(n1787), .C(n1807), .YC(n912), .YS(n913) );
  FAX1 U737 ( .A(n1907), .B(n1769), .C(n1879), .YC(n914), .YS(n915) );
  FAX1 U738 ( .A(n919), .B(n1969), .C(n1937), .YC(n916), .YS(n917) );
  INVX2 U739 ( .A(n918), .Y(n919) );
  FAX1 U740 ( .A(n925), .B(n942), .C(n923), .YC(n920), .YS(n921) );
  FAX1 U741 ( .A(n946), .B(n927), .C(n944), .YC(n922), .YS(n923) );
  FAX1 U742 ( .A(n948), .B(n931), .C(n929), .YC(n924), .YS(n925) );
  FAX1 U743 ( .A(n933), .B(n952), .C(n950), .YC(n926), .YS(n927) );
  FAX1 U744 ( .A(n954), .B(n935), .C(n937), .YC(n928), .YS(n929) );
  FAX1 U745 ( .A(n958), .B(n956), .C(n939), .YC(n930), .YS(n931) );
  FAX1 U746 ( .A(n1970), .B(n1938), .C(n2002), .YC(n932), .YS(n933) );
  FAX1 U747 ( .A(n1788), .B(n1908), .C(n1830), .YC(n934), .YS(n935) );
  FAX1 U748 ( .A(n1854), .B(n1770), .C(n1808), .YC(n936), .YS(n937) );
  FAX1 U749 ( .A(n960), .B(n1760), .C(n1880), .YC(n938), .YS(n939) );
  FAX1 U750 ( .A(n945), .B(n964), .C(n943), .YC(n940), .YS(n941) );
  FAX1 U751 ( .A(n968), .B(n947), .C(n966), .YC(n942), .YS(n943) );
  FAX1 U752 ( .A(n970), .B(n951), .C(n949), .YC(n944), .YS(n945) );
  FAX1 U753 ( .A(n953), .B(n974), .C(n972), .YC(n946), .YS(n947) );
  FAX1 U754 ( .A(n959), .B(n955), .C(n957), .YC(n948), .YS(n949) );
  FAX1 U755 ( .A(n980), .B(n976), .C(n978), .YC(n950), .YS(n951) );
  FAX1 U756 ( .A(n1909), .B(n1881), .C(n982), .YC(n952), .YS(n953) );
  FAX1 U757 ( .A(n1855), .B(n1809), .C(n1831), .YC(n954), .YS(n955) );
  FAX1 U758 ( .A(n1939), .B(n1771), .C(n1789), .YC(n956), .YS(n957) );
  FAX1 U759 ( .A(n961), .B(n2003), .C(n1971), .YC(n958), .YS(n959) );
  INVX2 U760 ( .A(n960), .Y(n961) );
  FAX1 U761 ( .A(n988), .B(n986), .C(n965), .YC(n962), .YS(n963) );
  FAX1 U762 ( .A(n990), .B(n969), .C(n967), .YC(n964), .YS(n965) );
  FAX1 U763 ( .A(n973), .B(n971), .C(n992), .YC(n966), .YS(n967) );
  FAX1 U764 ( .A(n996), .B(n994), .C(n975), .YC(n968), .YS(n969) );
  FAX1 U765 ( .A(n977), .B(n981), .C(n979), .YC(n970), .YS(n971) );
  FAX1 U766 ( .A(n1000), .B(n998), .C(n983), .YC(n972), .YS(n973) );
  FAX1 U767 ( .A(n2036), .B(n1004), .C(n1002), .YC(n974), .YS(n975) );
  FAX1 U768 ( .A(n2004), .B(n1832), .C(n1972), .YC(n976), .YS(n977) );
  FAX1 U769 ( .A(n1910), .B(n1810), .C(n1940), .YC(n978), .YS(n979) );
  FAX1 U770 ( .A(n1856), .B(n1772), .C(n1790), .YC(n980), .YS(n981) );
  FAX1 U771 ( .A(n1006), .B(n1761), .C(n1882), .YC(n982), .YS(n983) );
  FAX1 U772 ( .A(n989), .B(n1010), .C(n987), .YC(n984), .YS(n985) );
  FAX1 U773 ( .A(n1014), .B(n991), .C(n1012), .YC(n986), .YS(n987) );
  FAX1 U774 ( .A(n995), .B(n1016), .C(n993), .YC(n988), .YS(n989) );
  FAX1 U775 ( .A(n1020), .B(n1018), .C(n997), .YC(n990), .YS(n991) );
  FAX1 U776 ( .A(n1003), .B(n1001), .C(n1022), .YC(n992), .YS(n993) );
  FAX1 U777 ( .A(n1024), .B(n1005), .C(n999), .YC(n994), .YS(n995) );
  FAX1 U778 ( .A(n1030), .B(n1028), .C(n1026), .YC(n996), .YS(n997) );
  FAX1 U779 ( .A(n1911), .B(n1857), .C(n1883), .YC(n998), .YS(n999) );
  FAX1 U780 ( .A(n1811), .B(n1941), .C(n1833), .YC(n1000), .YS(n1001) );
  FAX1 U781 ( .A(n1973), .B(n1773), .C(n1791), .YC(n1002), .YS(n1003) );
  FAX1 U782 ( .A(n1007), .B(n2037), .C(n2005), .YC(n1004), .YS(n1005) );
  INVX2 U783 ( .A(n1006), .Y(n1007) );
  FAX1 U784 ( .A(n1013), .B(n1034), .C(n1011), .YC(n1008), .YS(n1009) );
  FAX1 U785 ( .A(n1038), .B(n1015), .C(n1036), .YC(n1010), .YS(n1011) );
  FAX1 U786 ( .A(n1019), .B(n1040), .C(n1017), .YC(n1012), .YS(n1013) );
  FAX1 U787 ( .A(n1023), .B(n1042), .C(n1021), .YC(n1014), .YS(n1015) );
  FAX1 U788 ( .A(n1029), .B(n1046), .C(n1044), .YC(n1016), .YS(n1017) );
  FAX1 U789 ( .A(n1050), .B(n1025), .C(n1027), .YC(n1018), .YS(n1019) );
  FAX1 U790 ( .A(n1052), .B(n1048), .C(n1031), .YC(n1020), .YS(n1021) );
  FAX1 U791 ( .A(n2038), .B(n2070), .C(n1054), .YC(n1022), .YS(n1023) );
  FAX1 U792 ( .A(n2006), .B(n1834), .C(n1974), .YC(n1024), .YS(n1025) );
  FAX1 U793 ( .A(n1942), .B(n1774), .C(n1858), .YC(n1026), .YS(n1027) );
  FAX1 U794 ( .A(n1884), .B(n1792), .C(n1812), .YC(n1028), .YS(n1029) );
  FAX1 U795 ( .A(n1056), .B(n1762), .C(n1912), .YC(n1030), .YS(n1031) );
  FAX1 U796 ( .A(n1037), .B(n1060), .C(n1035), .YC(n1032), .YS(n1033) );
  FAX1 U797 ( .A(n1064), .B(n1039), .C(n1062), .YC(n1034), .YS(n1035) );
  FAX1 U798 ( .A(n1043), .B(n1066), .C(n1041), .YC(n1036), .YS(n1037) );
  FAX1 U799 ( .A(n1047), .B(n1045), .C(n1068), .YC(n1038), .YS(n1039) );
  FAX1 U800 ( .A(n1053), .B(n1072), .C(n1070), .YC(n1040), .YS(n1041) );
  FAX1 U801 ( .A(n1051), .B(n1049), .C(n1074), .YC(n1042), .YS(n1043) );
  FAX1 U802 ( .A(n1078), .B(n1076), .C(n1055), .YC(n1044), .YS(n1045) );
  FAX1 U803 ( .A(n1943), .B(n1082), .C(n1080), .YC(n1046), .YS(n1047) );
  FAX1 U804 ( .A(n1975), .B(n1859), .C(n1913), .YC(n1048), .YS(n1049) );
  FAX1 U805 ( .A(n1835), .B(n2007), .C(n1813), .YC(n1050), .YS(n1051) );
  FAX1 U806 ( .A(n2039), .B(n1775), .C(n1793), .YC(n1052), .YS(n1053) );
  FAX1 U807 ( .A(n1057), .B(n2071), .C(n1885), .YC(n1054), .YS(n1055) );
  INVX2 U808 ( .A(n1056), .Y(n1057) );
  FAX1 U809 ( .A(n1063), .B(n1086), .C(n1061), .YC(n1058), .YS(n1059) );
  FAX1 U810 ( .A(n1090), .B(n1065), .C(n1088), .YC(n1060), .YS(n1061) );
  FAX1 U811 ( .A(n1094), .B(n1092), .C(n1067), .YC(n1062), .YS(n1063) );
  FAX1 U812 ( .A(n1073), .B(n1071), .C(n1069), .YC(n1064), .YS(n1065) );
  FAX1 U813 ( .A(n1100), .B(n1098), .C(n1096), .YC(n1066), .YS(n1067) );
  FAX1 U814 ( .A(n1079), .B(n1081), .C(n1075), .YC(n1068), .YS(n1069) );
  FAX1 U815 ( .A(n1104), .B(n1102), .C(n1077), .YC(n1070), .YS(n1071) );
  FAX1 U816 ( .A(n1108), .B(n1106), .C(n1083), .YC(n1072), .YS(n1073) );
  FAX1 U817 ( .A(n2072), .B(n2040), .C(n2104), .YC(n1074), .YS(n1075) );
  FAX1 U818 ( .A(n1860), .B(n2008), .C(n1976), .YC(n1076), .YS(n1077) );
  FAX1 U819 ( .A(n1914), .B(n1776), .C(n1836), .YC(n1078), .YS(n1079) );
  FAX1 U820 ( .A(n1886), .B(n1794), .C(n1814), .YC(n1080), .YS(n1081) );
  FAX1 U821 ( .A(n1110), .B(n1763), .C(n1944), .YC(n1082), .YS(n1083) );
  FAX1 U822 ( .A(n1089), .B(n1114), .C(n1087), .YC(n1084), .YS(n1085) );
  FAX1 U823 ( .A(n1118), .B(n1091), .C(n1116), .YC(n1086), .YS(n1087) );
  FAX1 U824 ( .A(n1095), .B(n1120), .C(n1093), .YC(n1088), .YS(n1089) );
  FAX1 U825 ( .A(n1099), .B(n1097), .C(n1122), .YC(n1090), .YS(n1091) );
  FAX1 U826 ( .A(n1128), .B(n1126), .C(n1124), .YC(n1092), .YS(n1093) );
  FAX1 U827 ( .A(n1105), .B(n1107), .C(n1101), .YC(n1094), .YS(n1095) );
  FAX1 U828 ( .A(n1132), .B(n1109), .C(n1103), .YC(n1096), .YS(n1097) );
  FAX1 U829 ( .A(n1136), .B(n1130), .C(n1134), .YC(n1098), .YS(n1099) );
  FAX1 U830 ( .A(n1915), .B(n1861), .C(n1138), .YC(n1100), .YS(n1101) );
  FAX1 U831 ( .A(n1945), .B(n1815), .C(n1837), .YC(n1102), .YS(n1103) );
  FAX1 U832 ( .A(n2009), .B(n1795), .C(n1977), .YC(n1104), .YS(n1105) );
  FAX1 U833 ( .A(n1887), .B(n2041), .C(n1777), .YC(n1106), .YS(n1107) );
  FAX1 U834 ( .A(n1111), .B(n2105), .C(n2073), .YC(n1108), .YS(n1109) );
  INVX2 U835 ( .A(n1110), .Y(n1111) );
  FAX1 U836 ( .A(n1117), .B(n1142), .C(n1115), .YC(n1112), .YS(n1113) );
  FAX1 U837 ( .A(n1146), .B(n1119), .C(n1144), .YC(n1114), .YS(n1115) );
  FAX1 U838 ( .A(n1123), .B(n1148), .C(n1121), .YC(n1116), .YS(n1117) );
  FAX1 U839 ( .A(n1127), .B(n1125), .C(n1150), .YC(n1118), .YS(n1119) );
  FAX1 U840 ( .A(n1154), .B(n1129), .C(n1152), .YC(n1120), .YS(n1121) );
  FAX1 U841 ( .A(n1137), .B(n1135), .C(n1156), .YC(n1122), .YS(n1123) );
  FAX1 U842 ( .A(n1162), .B(n1131), .C(n1133), .YC(n1124), .YS(n1125) );
  FAX1 U843 ( .A(n1160), .B(n1164), .C(n1139), .YC(n1126), .YS(n1127) );
  FAX1 U844 ( .A(n2138), .B(n1166), .C(n1158), .YC(n1128), .YS(n1129) );
  FAX1 U845 ( .A(n2074), .B(n2106), .C(n1888), .YC(n1130), .YS(n1131) );
  FAX1 U846 ( .A(n1862), .B(n2010), .C(n2042), .YC(n1132), .YS(n1133) );
  FAX1 U847 ( .A(n1978), .B(n1796), .C(n1838), .YC(n1134), .YS(n1135) );
  FAX1 U848 ( .A(n1916), .B(n1778), .C(n1816), .YC(n1136), .YS(n1137) );
  FAX1 U849 ( .A(n1168), .B(n1764), .C(n1946), .YC(n1138), .YS(n1139) );
  FAX1 U850 ( .A(n1145), .B(n1172), .C(n1143), .YC(n1140), .YS(n1141) );
  FAX1 U851 ( .A(n1176), .B(n1147), .C(n1174), .YC(n1142), .YS(n1143) );
  FAX1 U852 ( .A(n1151), .B(n1178), .C(n1149), .YC(n1144), .YS(n1145) );
  FAX1 U853 ( .A(n1155), .B(n1153), .C(n1180), .YC(n1146), .YS(n1147) );
  FAX1 U854 ( .A(n1184), .B(n1157), .C(n1182), .YC(n1148), .YS(n1149) );
  FAX1 U855 ( .A(n1163), .B(n1188), .C(n1186), .YC(n1150), .YS(n1151) );
  FAX1 U856 ( .A(n1159), .B(n1165), .C(n1161), .YC(n1152), .YS(n1153) );
  FAX1 U857 ( .A(n1194), .B(n1196), .C(n1167), .YC(n1154), .YS(n1155) );
  FAX1 U858 ( .A(n1198), .B(n1190), .C(n1192), .YC(n1156), .YS(n1157) );
  FAX1 U859 ( .A(n1947), .B(n1863), .C(n1917), .YC(n1158), .YS(n1159) );
  FAX1 U860 ( .A(n1979), .B(n1817), .C(n1839), .YC(n1160), .YS(n1161) );
  FAX1 U861 ( .A(n2043), .B(n1797), .C(n2011), .YC(n1162), .YS(n1163) );
  FAX1 U862 ( .A(n1889), .B(n2075), .C(n1779), .YC(n1164), .YS(n1165) );
  FAX1 U863 ( .A(n1169), .B(n2139), .C(n2107), .YC(n1166), .YS(n1167) );
  INVX2 U864 ( .A(n1168), .Y(n1169) );
  FAX1 U865 ( .A(n1175), .B(n1202), .C(n1173), .YC(n1170), .YS(n1171) );
  FAX1 U866 ( .A(n1206), .B(n1177), .C(n1204), .YC(n1172), .YS(n1173) );
  FAX1 U867 ( .A(n1181), .B(n1208), .C(n1179), .YC(n1174), .YS(n1175) );
  FAX1 U868 ( .A(n1185), .B(n1183), .C(n1210), .YC(n1176), .YS(n1177) );
  FAX1 U869 ( .A(n1214), .B(n1212), .C(n1187), .YC(n1178), .YS(n1179) );
  FAX1 U870 ( .A(n1218), .B(n1189), .C(n1216), .YC(n1180), .YS(n1181) );
  FAX1 U871 ( .A(n1195), .B(n1197), .C(n1193), .YC(n1182), .YS(n1183) );
  FAX1 U872 ( .A(n1224), .B(n1222), .C(n1191), .YC(n1184), .YS(n1185) );
  FAX1 U873 ( .A(n1220), .B(n1226), .C(n1199), .YC(n1186), .YS(n1187) );
  FAX1 U874 ( .A(n2076), .B(n2172), .C(n1228), .YC(n1188), .YS(n1189) );
  FAX1 U875 ( .A(n2108), .B(n2044), .C(n2140), .YC(n1190), .YS(n1191) );
  FAX1 U876 ( .A(n1864), .B(n1948), .C(n1890), .YC(n1192), .YS(n1193) );
  FAX1 U877 ( .A(n2012), .B(n1840), .C(n1818), .YC(n1194), .YS(n1195) );
  FAX1 U878 ( .A(n1918), .B(n1798), .C(n1780), .YC(n1196), .YS(n1197) );
  FAX1 U879 ( .A(n1230), .B(n1765), .C(n1980), .YC(n1198), .YS(n1199) );
  FAX1 U880 ( .A(n1205), .B(n1234), .C(n1203), .YC(n1200), .YS(n1201) );
  FAX1 U881 ( .A(n1238), .B(n1207), .C(n1236), .YC(n1202), .YS(n1203) );
  FAX1 U882 ( .A(n1240), .B(n1211), .C(n1209), .YC(n1204), .YS(n1205) );
  FAX1 U883 ( .A(n1217), .B(n1213), .C(n1242), .YC(n1206), .YS(n1207) );
  FAX1 U884 ( .A(n1246), .B(n1244), .C(n1215), .YC(n1208), .YS(n1209) );
  FAX1 U885 ( .A(n1250), .B(n1248), .C(n1219), .YC(n1210), .YS(n1211) );
  FAX1 U886 ( .A(n1225), .B(n1227), .C(n1223), .YC(n1212), .YS(n1213) );
  FAX1 U887 ( .A(n1256), .B(n1254), .C(n1221), .YC(n1214), .YS(n1215) );
  FAX1 U888 ( .A(n1252), .B(n1258), .C(n1229), .YC(n1216), .YS(n1217) );
  FAX1 U889 ( .A(n1981), .B(n2013), .C(n1260), .YC(n1218), .YS(n1219) );
  FAX1 U890 ( .A(n2045), .B(n1919), .C(n1949), .YC(n1220), .YS(n1221) );
  FAX1 U891 ( .A(n1865), .B(n2077), .C(n1891), .YC(n1222), .YS(n1223) );
  FAX1 U892 ( .A(n2109), .B(n1819), .C(n1841), .YC(n1224), .YS(n1225) );
  FAX1 U893 ( .A(n2141), .B(n1781), .C(n1799), .YC(n1226), .YS(n1227) );
  FAX1 U894 ( .A(n1766), .B(n1262), .C(n2173), .YC(n1228), .YS(n1229) );
  FAX1 U896 ( .A(n1237), .B(n1265), .C(n1235), .YC(n1232), .YS(n1233) );
  FAX1 U897 ( .A(n1269), .B(n1239), .C(n1267), .YC(n1234), .YS(n1235) );
  FAX1 U898 ( .A(n1271), .B(n1243), .C(n1241), .YC(n1236), .YS(n1237) );
  FAX1 U899 ( .A(n1247), .B(n1245), .C(n1273), .YC(n1238), .YS(n1239) );
  FAX1 U900 ( .A(n1251), .B(n1275), .C(n1249), .YC(n1240), .YS(n1241) );
  FAX1 U901 ( .A(n1255), .B(n1279), .C(n1277), .YC(n1242), .YS(n1243) );
  FAX1 U902 ( .A(n1257), .B(n1259), .C(n1281), .YC(n1244), .YS(n1245) );
  FAX1 U903 ( .A(n1285), .B(n1261), .C(n1253), .YC(n1246), .YS(n1247) );
  FAX1 U904 ( .A(n1283), .B(n1289), .C(n1287), .YC(n1248), .YS(n1249) );
  FAX1 U905 ( .A(n2110), .B(n2206), .C(n1291), .YC(n1250), .YS(n1251) );
  FAX1 U906 ( .A(n2142), .B(n2078), .C(n2174), .YC(n1252), .YS(n1253) );
  FAX1 U907 ( .A(n1892), .B(n1982), .C(n1920), .YC(n1254), .YS(n1255) );
  FAX1 U908 ( .A(n2046), .B(n1866), .C(n1842), .YC(n1256), .YS(n1257) );
  FAX1 U909 ( .A(n1950), .B(n1820), .C(n1782), .YC(n1258), .YS(n1259) );
  FAX1 U910 ( .A(n1262), .B(n1800), .C(n2014), .YC(n1260), .YS(n1261) );
  INVX2 U911 ( .A(n1230), .Y(n1262) );
  FAX1 U912 ( .A(n1268), .B(n1295), .C(n1266), .YC(n1263), .YS(n1264) );
  FAX1 U913 ( .A(n1272), .B(n1270), .C(n1297), .YC(n1265), .YS(n1266) );
  FAX1 U914 ( .A(n1274), .B(n1301), .C(n1299), .YC(n1267), .YS(n1268) );
  FAX1 U915 ( .A(n1278), .B(n1276), .C(n1303), .YC(n1269), .YS(n1270) );
  FAX1 U916 ( .A(n1307), .B(n1305), .C(n1280), .YC(n1271), .YS(n1272) );
  FAX1 U917 ( .A(n1288), .B(n1282), .C(n1309), .YC(n1273), .YS(n1274) );
  FAX1 U918 ( .A(n1284), .B(n1290), .C(n1286), .YC(n1275), .YS(n1276) );
  FAX1 U919 ( .A(n1311), .B(n1315), .C(n1292), .YC(n1277), .YS(n1278) );
  FAX1 U920 ( .A(n1313), .B(n1319), .C(n1317), .YC(n1279), .YS(n1280) );
  FAX1 U921 ( .A(n2015), .B(n2047), .C(n1321), .YC(n1281), .YS(n1282) );
  FAX1 U922 ( .A(n2079), .B(n1921), .C(n1951), .YC(n1283), .YS(n1284) );
  FAX1 U923 ( .A(n2111), .B(n1867), .C(n1893), .YC(n1285), .YS(n1286) );
  FAX1 U924 ( .A(n1983), .B(n2143), .C(n1843), .YC(n1287), .YS(n1288) );
  FAX1 U925 ( .A(n2175), .B(n1801), .C(n1821), .YC(n1289), .YS(n1290) );
  FAX1 U926 ( .A(n1767), .B(n2207), .C(n1783), .YC(n1291), .YS(n1292) );
  FAX1 U927 ( .A(n1298), .B(n1325), .C(n1296), .YC(n1293), .YS(n1294) );
  FAX1 U928 ( .A(n1302), .B(n1300), .C(n1327), .YC(n1295), .YS(n1296) );
  FAX1 U929 ( .A(n1304), .B(n1331), .C(n1329), .YC(n1297), .YS(n1298) );
  FAX1 U930 ( .A(n1308), .B(n1333), .C(n1306), .YC(n1299), .YS(n1300) );
  FAX1 U931 ( .A(n1337), .B(n1310), .C(n1335), .YC(n1301), .YS(n1302) );
  FAX1 U932 ( .A(n1314), .B(n1316), .C(n1339), .YC(n1303), .YS(n1304) );
  FAX1 U933 ( .A(n1312), .B(n1320), .C(n1318), .YC(n1305), .YS(n1306) );
  FAX1 U934 ( .A(n1341), .B(n1345), .C(n1343), .YC(n1307), .YS(n1308) );
  FAX1 U935 ( .A(n1322), .B(n1349), .C(n1347), .YC(n1309), .YS(n1310) );
  FAX1 U936 ( .A(n1868), .B(n2016), .C(n1922), .YC(n1311), .YS(n1312) );
  FAX1 U937 ( .A(n2048), .B(n1822), .C(n1844), .YC(n1313), .YS(n1314) );
  FAX1 U938 ( .A(n1894), .B(n2112), .C(n2080), .YC(n1315), .YS(n1316) );
  FAX1 U939 ( .A(n1984), .B(n2176), .C(n2144), .YC(n1317), .YS(n1318) );
  FAX1 U940 ( .A(n1952), .B(n1784), .C(n1802), .YC(n1319), .YS(n1320) );
  HAX1 U941 ( .A(n2208), .B(n1743), .YC(n1321), .YS(n1322) );
  FAX1 U942 ( .A(n1328), .B(n1353), .C(n1326), .YC(n1323), .YS(n1324) );
  FAX1 U943 ( .A(n1332), .B(n1330), .C(n1355), .YC(n1325), .YS(n1326) );
  FAX1 U944 ( .A(n1334), .B(n1359), .C(n1357), .YC(n1327), .YS(n1328) );
  FAX1 U945 ( .A(n1361), .B(n1338), .C(n1336), .YC(n1329), .YS(n1330) );
  FAX1 U946 ( .A(n1365), .B(n1340), .C(n1363), .YC(n1331), .YS(n1332) );
  FAX1 U947 ( .A(n1344), .B(n1346), .C(n1367), .YC(n1333), .YS(n1334) );
  FAX1 U948 ( .A(n1350), .B(n1342), .C(n1348), .YC(n1335), .YS(n1336) );
  FAX1 U949 ( .A(n1371), .B(n1375), .C(n1373), .YC(n1337), .YS(n1338) );
  FAX1 U950 ( .A(n2955), .B(n1377), .C(n1369), .YC(n1339), .YS(n1340) );
  FAX1 U951 ( .A(n2017), .B(n1953), .C(n1985), .YC(n1341), .YS(n1342) );
  FAX1 U952 ( .A(n2049), .B(n1895), .C(n1923), .YC(n1343), .YS(n1344) );
  FAX1 U953 ( .A(n2081), .B(n1845), .C(n1869), .YC(n1345), .YS(n1346) );
  FAX1 U954 ( .A(n2145), .B(n1823), .C(n2113), .YC(n1347), .YS(n1348) );
  FAX1 U955 ( .A(n2209), .B(n2177), .C(n1803), .YC(n1349), .YS(n1350) );
  FAX1 U956 ( .A(n1356), .B(n1381), .C(n1354), .YC(n1351), .YS(n1352) );
  FAX1 U957 ( .A(n1385), .B(n1358), .C(n1383), .YC(n1353), .YS(n1354) );
  FAX1 U958 ( .A(n1362), .B(n1387), .C(n1360), .YC(n1355), .YS(n1356) );
  FAX1 U959 ( .A(n1366), .B(n1389), .C(n1364), .YC(n1357), .YS(n1358) );
  FAX1 U960 ( .A(n1368), .B(n1393), .C(n1391), .YC(n1359), .YS(n1360) );
  FAX1 U961 ( .A(n1374), .B(n1376), .C(n1395), .YC(n1361), .YS(n1362) );
  FAX1 U962 ( .A(n1401), .B(n1370), .C(n1372), .YC(n1363), .YS(n1364) );
  FAX1 U963 ( .A(n1403), .B(n1397), .C(n1399), .YC(n1365), .YS(n1366) );
  FAX1 U964 ( .A(n2018), .B(n2050), .C(n1378), .YC(n1367), .YS(n1368) );
  FAX1 U965 ( .A(n2082), .B(n1924), .C(n1954), .YC(n1369), .YS(n1370) );
  FAX1 U966 ( .A(n1846), .B(n1824), .C(n1870), .YC(n1371), .YS(n1372) );
  FAX1 U967 ( .A(n1896), .B(n2114), .C(n1804), .YC(n1373), .YS(n1374) );
  FAX1 U968 ( .A(n1986), .B(n2178), .C(n2146), .YC(n1375), .YS(n1376) );
  HAX1 U969 ( .A(n2210), .B(n1744), .YC(n1377), .YS(n1378) );
  FAX1 U970 ( .A(n1384), .B(n1407), .C(n1382), .YC(n1379), .YS(n1380) );
  FAX1 U971 ( .A(n1411), .B(n1386), .C(n1409), .YC(n1381), .YS(n1382) );
  FAX1 U972 ( .A(n1390), .B(n1413), .C(n1388), .YC(n1383), .YS(n1384) );
  FAX1 U973 ( .A(n1394), .B(n1415), .C(n1392), .YC(n1385), .YS(n1386) );
  FAX1 U974 ( .A(n1396), .B(n1419), .C(n1417), .YC(n1387), .YS(n1388) );
  FAX1 U975 ( .A(n1400), .B(n1398), .C(n1402), .YC(n1389), .YS(n1390) );
  FAX1 U976 ( .A(n1421), .B(n1423), .C(n1404), .YC(n1391), .YS(n1392) );
  FAX1 U977 ( .A(n1429), .B(n1427), .C(n1425), .YC(n1393), .YS(n1394) );
  FAX1 U978 ( .A(n2019), .B(n1987), .C(n2930), .YC(n1395), .YS(n1396) );
  FAX1 U979 ( .A(n2051), .B(n1925), .C(n1955), .YC(n1397), .YS(n1398) );
  FAX1 U980 ( .A(n2083), .B(n1871), .C(n1897), .YC(n1399), .YS(n1400) );
  FAX1 U981 ( .A(n2147), .B(n1847), .C(n2115), .YC(n1401), .YS(n1402) );
  FAX1 U982 ( .A(n2211), .B(n2179), .C(n1825), .YC(n1403), .YS(n1404) );
  FAX1 U983 ( .A(n1410), .B(n1433), .C(n1408), .YC(n1405), .YS(n1406) );
  FAX1 U984 ( .A(n1414), .B(n1412), .C(n1435), .YC(n1407), .YS(n1408) );
  FAX1 U985 ( .A(n1416), .B(n1439), .C(n1437), .YC(n1409), .YS(n1410) );
  FAX1 U986 ( .A(n1420), .B(n1441), .C(n1418), .YC(n1411), .YS(n1412) );
  FAX1 U987 ( .A(n1424), .B(n1445), .C(n1443), .YC(n1413), .YS(n1414) );
  FAX1 U988 ( .A(n1422), .B(n1428), .C(n1426), .YC(n1415), .YS(n1416) );
  FAX1 U989 ( .A(n1447), .B(n1449), .C(n1451), .YC(n1417), .YS(n1418) );
  FAX1 U990 ( .A(n2084), .B(n1430), .C(n1453), .YC(n1419), .YS(n1420) );
  FAX1 U991 ( .A(n2116), .B(n1956), .C(n2052), .YC(n1421), .YS(n1422) );
  FAX1 U992 ( .A(n2148), .B(n1898), .C(n1926), .YC(n1423), .YS(n1424) );
  FAX1 U993 ( .A(n2020), .B(n1872), .C(n2180), .YC(n1425), .YS(n1426) );
  FAX1 U994 ( .A(n1988), .B(n1826), .C(n1848), .YC(n1427), .YS(n1428) );
  HAX1 U995 ( .A(n2212), .B(n1745), .YC(n1429), .YS(n1430) );
  FAX1 U996 ( .A(n1436), .B(n1457), .C(n1434), .YC(n1431), .YS(n1432) );
  FAX1 U997 ( .A(n1461), .B(n1459), .C(n1438), .YC(n1433), .YS(n1434) );
  FAX1 U998 ( .A(n1444), .B(n1442), .C(n1440), .YC(n1435), .YS(n1436) );
  FAX1 U999 ( .A(n1467), .B(n1465), .C(n1463), .YC(n1437), .YS(n1438) );
  FAX1 U1000 ( .A(n1452), .B(n1450), .C(n1446), .YC(n1439), .YS(n1440) );
  FAX1 U1001 ( .A(n1473), .B(n1454), .C(n1448), .YC(n1441), .YS(n1442) );
  FAX1 U1002 ( .A(n1475), .B(n1469), .C(n1471), .YC(n1443), .YS(n1444) );
  FAX1 U1003 ( .A(n2053), .B(n2956), .C(n1477), .YC(n1445), .YS(n1446) );
  FAX1 U1004 ( .A(n2085), .B(n1989), .C(n2021), .YC(n1447), .YS(n1448) );
  FAX1 U1005 ( .A(n2117), .B(n1927), .C(n1957), .YC(n1449), .YS(n1450) );
  FAX1 U1006 ( .A(n2149), .B(n1873), .C(n1899), .YC(n1451), .YS(n1452) );
  FAX1 U1007 ( .A(n2213), .B(n2181), .C(n1849), .YC(n1453), .YS(n1454) );
  FAX1 U1008 ( .A(n1460), .B(n1481), .C(n1458), .YC(n1455), .YS(n1456) );
  FAX1 U1009 ( .A(n1485), .B(n1483), .C(n1462), .YC(n1457), .YS(n1458) );
  FAX1 U1010 ( .A(n1487), .B(n1466), .C(n1464), .YC(n1459), .YS(n1460) );
  FAX1 U1011 ( .A(n1491), .B(n1489), .C(n1468), .YC(n1461), .YS(n1462) );
  FAX1 U1012 ( .A(n1472), .B(n1476), .C(n1474), .YC(n1463), .YS(n1464) );
  FAX1 U1013 ( .A(n1495), .B(n1493), .C(n1470), .YC(n1465), .YS(n1466) );
  FAX1 U1014 ( .A(n1478), .B(n1499), .C(n1497), .YC(n1467), .YS(n1468) );
  FAX1 U1015 ( .A(n2086), .B(n1990), .C(n2054), .YC(n1469), .YS(n1470) );
  FAX1 U1016 ( .A(n2118), .B(n1900), .C(n1958), .YC(n1471), .YS(n1472) );
  FAX1 U1017 ( .A(n1928), .B(n1850), .C(n1874), .YC(n1473), .YS(n1474) );
  FAX1 U1018 ( .A(n2022), .B(n2182), .C(n2150), .YC(n1475), .YS(n1476) );
  HAX1 U1019 ( .A(n2214), .B(n1746), .YC(n1477), .YS(n1478) );
  FAX1 U1020 ( .A(n1484), .B(n1503), .C(n1482), .YC(n1479), .YS(n1480) );
  FAX1 U1021 ( .A(n1507), .B(n1486), .C(n1505), .YC(n1481), .YS(n1482) );
  FAX1 U1022 ( .A(n1509), .B(n1490), .C(n1488), .YC(n1483), .YS(n1484) );
  FAX1 U1023 ( .A(n1513), .B(n1511), .C(n1492), .YC(n1485), .YS(n1486) );
  FAX1 U1024 ( .A(n1494), .B(n1498), .C(n1496), .YC(n1487), .YS(n1488) );
  FAX1 U1025 ( .A(n1517), .B(n1515), .C(n1500), .YC(n1489), .YS(n1490) );
  FAX1 U1026 ( .A(n2952), .B(n1521), .C(n1519), .YC(n1491), .YS(n1492) );
  FAX1 U1027 ( .A(n2087), .B(n2023), .C(n2055), .YC(n1493), .YS(n1494) );
  FAX1 U1028 ( .A(n2119), .B(n1959), .C(n1991), .YC(n1495), .YS(n1496) );
  FAX1 U1029 ( .A(n2151), .B(n1901), .C(n1929), .YC(n1497), .YS(n1498) );
  FAX1 U1030 ( .A(n2215), .B(n2183), .C(n1875), .YC(n1499), .YS(n1500) );
  FAX1 U1031 ( .A(n1506), .B(n1525), .C(n1504), .YC(n1501), .YS(n1502) );
  FAX1 U1032 ( .A(n1529), .B(n1508), .C(n1527), .YC(n1503), .YS(n1504) );
  FAX1 U1033 ( .A(n1531), .B(n1512), .C(n1510), .YC(n1505), .YS(n1506) );
  FAX1 U1034 ( .A(n1518), .B(n1514), .C(n1533), .YC(n1507), .YS(n1508) );
  FAX1 U1035 ( .A(n1516), .B(n1520), .C(n1535), .YC(n1509), .YS(n1510) );
  FAX1 U1036 ( .A(n1541), .B(n1539), .C(n1537), .YC(n1511), .YS(n1512) );
  FAX1 U1037 ( .A(n2088), .B(n1992), .C(n1522), .YC(n1513), .YS(n1514) );
  FAX1 U1038 ( .A(n2120), .B(n1930), .C(n1960), .YC(n1515), .YS(n1516) );
  FAX1 U1039 ( .A(n2056), .B(n2184), .C(n2152), .YC(n1517), .YS(n1518) );
  FAX1 U1040 ( .A(n2024), .B(n1876), .C(n1902), .YC(n1519), .YS(n1520) );
  HAX1 U1041 ( .A(n2216), .B(n1747), .YC(n1521), .YS(n1522) );
  FAX1 U1042 ( .A(n1528), .B(n1545), .C(n1526), .YC(n1523), .YS(n1524) );
  FAX1 U1043 ( .A(n1532), .B(n1530), .C(n1547), .YC(n1525), .YS(n1526) );
  FAX1 U1044 ( .A(n1551), .B(n1534), .C(n1549), .YC(n1527), .YS(n1528) );
  FAX1 U1045 ( .A(n1540), .B(n1536), .C(n1553), .YC(n1529), .YS(n1530) );
  FAX1 U1046 ( .A(n1555), .B(n1542), .C(n1538), .YC(n1531), .YS(n1532) );
  FAX1 U1047 ( .A(n1561), .B(n1559), .C(n1557), .YC(n1533), .YS(n1534) );
  FAX1 U1048 ( .A(n2089), .B(n2057), .C(n2927), .YC(n1535), .YS(n1536) );
  FAX1 U1049 ( .A(n2121), .B(n1993), .C(n2025), .YC(n1537), .YS(n1538) );
  FAX1 U1050 ( .A(n2153), .B(n1931), .C(n1961), .YC(n1539), .YS(n1540) );
  FAX1 U1051 ( .A(n2217), .B(n2185), .C(n1903), .YC(n1541), .YS(n1542) );
  FAX1 U1052 ( .A(n1548), .B(n1565), .C(n1546), .YC(n1543), .YS(n1544) );
  FAX1 U1053 ( .A(n1552), .B(n1550), .C(n1567), .YC(n1545), .YS(n1546) );
  FAX1 U1054 ( .A(n1571), .B(n1554), .C(n1569), .YC(n1547), .YS(n1548) );
  FAX1 U1055 ( .A(n1558), .B(n1560), .C(n1573), .YC(n1549), .YS(n1550) );
  FAX1 U1056 ( .A(n1577), .B(n1575), .C(n1556), .YC(n1551), .YS(n1552) );
  FAX1 U1057 ( .A(n1994), .B(n1562), .C(n1579), .YC(n1553), .YS(n1554) );
  FAX1 U1058 ( .A(n2058), .B(n1904), .C(n1932), .YC(n1555), .YS(n1556) );
  FAX1 U1059 ( .A(n1962), .B(n2122), .C(n2090), .YC(n1557), .YS(n1558) );
  FAX1 U1060 ( .A(n2026), .B(n2186), .C(n2154), .YC(n1559), .YS(n1560) );
  HAX1 U1061 ( .A(n2218), .B(n1748), .YC(n1561), .YS(n1562) );
  FAX1 U1062 ( .A(n1568), .B(n1583), .C(n1566), .YC(n1563), .YS(n1564) );
  FAX1 U1063 ( .A(n1572), .B(n1570), .C(n1585), .YC(n1565), .YS(n1566) );
  FAX1 U1064 ( .A(n1574), .B(n1589), .C(n1587), .YC(n1567), .YS(n1568) );
  FAX1 U1065 ( .A(n1580), .B(n1576), .C(n1578), .YC(n1569), .YS(n1570) );
  FAX1 U1066 ( .A(n1595), .B(n1591), .C(n1593), .YC(n1571), .YS(n1572) );
  FAX1 U1067 ( .A(n2091), .B(n2947), .C(n1597), .YC(n1573), .YS(n1574) );
  FAX1 U1068 ( .A(n2123), .B(n2027), .C(n2059), .YC(n1575), .YS(n1576) );
  FAX1 U1069 ( .A(n2155), .B(n1963), .C(n1995), .YC(n1577), .YS(n1578) );
  FAX1 U1070 ( .A(n2219), .B(n2187), .C(n1933), .YC(n1579), .YS(n1580) );
  FAX1 U1071 ( .A(n1586), .B(n1601), .C(n1584), .YC(n1581), .YS(n1582) );
  FAX1 U1072 ( .A(n1590), .B(n1588), .C(n1603), .YC(n1583), .YS(n1584) );
  FAX1 U1073 ( .A(n1596), .B(n1607), .C(n1605), .YC(n1585), .YS(n1586) );
  FAX1 U1074 ( .A(n1609), .B(n1592), .C(n1594), .YC(n1587), .YS(n1588) );
  FAX1 U1075 ( .A(n1598), .B(n1613), .C(n1611), .YC(n1589), .YS(n1590) );
  FAX1 U1076 ( .A(n2156), .B(n2028), .C(n2124), .YC(n1591), .YS(n1592) );
  FAX1 U1077 ( .A(n2092), .B(n2188), .C(n1996), .YC(n1593), .YS(n1594) );
  FAX1 U1078 ( .A(n2060), .B(n1934), .C(n1964), .YC(n1595), .YS(n1596) );
  HAX1 U1079 ( .A(n2220), .B(n1749), .YC(n1597), .YS(n1598) );
  FAX1 U1080 ( .A(n1604), .B(n1617), .C(n1602), .YC(n1599), .YS(n1600) );
  FAX1 U1081 ( .A(n1608), .B(n1606), .C(n1619), .YC(n1601), .YS(n1602) );
  FAX1 U1082 ( .A(n1612), .B(n1623), .C(n1621), .YC(n1603), .YS(n1604) );
  FAX1 U1083 ( .A(n1625), .B(n1614), .C(n1610), .YC(n1605), .YS(n1606) );
  FAX1 U1084 ( .A(n2948), .B(n1629), .C(n1627), .YC(n1607), .YS(n1608) );
  FAX1 U1085 ( .A(n2125), .B(n2061), .C(n2093), .YC(n1609), .YS(n1610) );
  FAX1 U1086 ( .A(n2157), .B(n1997), .C(n2029), .YC(n1611), .YS(n1612) );
  FAX1 U1087 ( .A(n2221), .B(n2189), .C(n1965), .YC(n1613), .YS(n1614) );
  FAX1 U1088 ( .A(n1620), .B(n1633), .C(n1618), .YC(n1615), .YS(n1616) );
  FAX1 U1089 ( .A(n1637), .B(n1622), .C(n1635), .YC(n1617), .YS(n1618) );
  FAX1 U1090 ( .A(n1628), .B(n1639), .C(n1624), .YC(n1619), .YS(n1620) );
  FAX1 U1091 ( .A(n1643), .B(n1641), .C(n1626), .YC(n1621), .YS(n1622) );
  FAX1 U1092 ( .A(n2094), .B(n2030), .C(n1630), .YC(n1623), .YS(n1624) );
  FAX1 U1093 ( .A(n2126), .B(n1966), .C(n1998), .YC(n1625), .YS(n1626) );
  FAX1 U1094 ( .A(n2062), .B(n2190), .C(n2158), .YC(n1627), .YS(n1628) );
  HAX1 U1095 ( .A(n2222), .B(n1750), .YC(n1629), .YS(n1630) );
  FAX1 U1096 ( .A(n1636), .B(n1647), .C(n1634), .YC(n1631), .YS(n1632) );
  FAX1 U1097 ( .A(n1651), .B(n1649), .C(n1638), .YC(n1633), .YS(n1634) );
  FAX1 U1098 ( .A(n1644), .B(n1642), .C(n1640), .YC(n1635), .YS(n1636) );
  FAX1 U1099 ( .A(n1657), .B(n1655), .C(n1653), .YC(n1637), .YS(n1638) );
  FAX1 U1100 ( .A(n2127), .B(n2095), .C(n2926), .YC(n1639), .YS(n1640) );
  FAX1 U1101 ( .A(n2159), .B(n2031), .C(n2063), .YC(n1641), .YS(n1642) );
  FAX1 U1102 ( .A(n2223), .B(n2191), .C(n1999), .YC(n1643), .YS(n1644) );
  FAX1 U1103 ( .A(n1650), .B(n1661), .C(n1648), .YC(n1645), .YS(n1646) );
  FAX1 U1104 ( .A(n1665), .B(n1652), .C(n1663), .YC(n1647), .YS(n1648) );
  FAX1 U1106 ( .A(n2160), .B(n1658), .C(n1669), .YC(n1651), .YS(n1652) );
  FAX1 U1107 ( .A(n2192), .B(n2064), .C(n2128), .YC(n1653), .YS(n1654) );
  FAX1 U1108 ( .A(n2096), .B(n2000), .C(n2032), .YC(n1655), .YS(n1656) );
  HAX1 U1109 ( .A(n2224), .B(n1751), .YC(n1657), .YS(n1658) );
  FAX1 U1110 ( .A(n1664), .B(n1673), .C(n1662), .YC(n1659), .YS(n1660) );
  FAX1 U1111 ( .A(n1668), .B(n1666), .C(n1675), .YC(n1661), .YS(n1662) );
  FAX1 U1112 ( .A(n1679), .B(n1677), .C(n1670), .YC(n1663), .YS(n1664) );
  FAX1 U1113 ( .A(n2129), .B(n2949), .C(n1681), .YC(n1665), .YS(n1666) );
  FAX1 U1114 ( .A(n2161), .B(n2065), .C(n2097), .YC(n1667), .YS(n1668) );
  FAX1 U1115 ( .A(n2033), .B(n2193), .C(n2225), .YC(n1669), .YS(n1670) );
  FAX1 U1116 ( .A(n1685), .B(n1676), .C(n1674), .YC(n1671), .YS(n1672) );
  FAX1 U1117 ( .A(n1678), .B(n1680), .C(n1687), .YC(n1673), .YS(n1674) );
  FAX1 U1119 ( .A(n2130), .B(n2034), .C(n2066), .YC(n1677), .YS(n1678) );
  FAX1 U1120 ( .A(n2098), .B(n2194), .C(n2162), .YC(n1679), .YS(n1680) );
  HAX1 U1121 ( .A(n2226), .B(n1752), .YC(n1681), .YS(n1682) );
  FAX1 U1122 ( .A(n1688), .B(n1695), .C(n1686), .YC(n1683), .YS(n1684) );
  FAX1 U1123 ( .A(n1692), .B(n1690), .C(n1697), .YC(n1685), .YS(n1686) );
  FAX1 U1124 ( .A(n2950), .B(n1701), .C(n1699), .YC(n1687), .YS(n1688) );
  FAX1 U1125 ( .A(n2163), .B(n2131), .C(n2099), .YC(n1689), .YS(n1690) );
  FAX1 U1126 ( .A(n2227), .B(n2195), .C(n2067), .YC(n1691), .YS(n1692) );
  FAX1 U1127 ( .A(n1698), .B(n1705), .C(n1696), .YC(n1693), .YS(n1694) );
  FAX1 U1128 ( .A(n1709), .B(n1700), .C(n1707), .YC(n1695), .YS(n1696) );
  FAX1 U1129 ( .A(n2164), .B(n2100), .C(n1702), .YC(n1697), .YS(n1698) );
  FAX1 U1130 ( .A(n2132), .B(n2068), .C(n2196), .YC(n1699), .YS(n1700) );
  HAX1 U1131 ( .A(n1753), .B(n2228), .YC(n1701), .YS(n1702) );
  FAX1 U1132 ( .A(n1708), .B(n1713), .C(n1706), .YC(n1703), .YS(n1704) );
  FAX1 U1133 ( .A(n1717), .B(n1715), .C(n1710), .YC(n1705), .YS(n1706) );
  FAX1 U1134 ( .A(n2165), .B(n2133), .C(n2069), .YC(n1707), .YS(n1708) );
  FAX1 U1135 ( .A(n2229), .B(n2197), .C(n2101), .YC(n1709), .YS(n1710) );
  FAX1 U1136 ( .A(n1716), .B(n1721), .C(n1714), .YC(n1711), .YS(n1712) );
  FAX1 U1137 ( .A(n2198), .B(n1718), .C(n1723), .YC(n1713), .YS(n1714) );
  FAX1 U1138 ( .A(n2134), .B(n2102), .C(n2166), .YC(n1715), .YS(n1716) );
  HAX1 U1139 ( .A(n2230), .B(n1754), .YC(n1717), .YS(n1718) );
  FAX1 U1140 ( .A(n1727), .B(n1724), .C(n1722), .YC(n1719), .YS(n1720) );
  FAX1 U1141 ( .A(n2167), .B(n2951), .C(n1729), .YC(n1721), .YS(n1722) );
  FAX1 U1142 ( .A(n2231), .B(n2199), .C(n2135), .YC(n1723), .YS(n1724) );
  FAX1 U1143 ( .A(n1730), .B(n1733), .C(n1728), .YC(n1725), .YS(n1726) );
  FAX1 U1144 ( .A(n2200), .B(n2136), .C(n2168), .YC(n1727), .YS(n1728) );
  HAX1 U1145 ( .A(n2232), .B(n1755), .YC(n1729), .YS(n1730) );
  FAX1 U1146 ( .A(n2953), .B(n1737), .C(n1734), .YC(n1731), .YS(n1732) );
  FAX1 U1147 ( .A(n2233), .B(n2201), .C(n2169), .YC(n1733), .YS(n1734) );
  FAX1 U1148 ( .A(n2202), .B(n2170), .C(n1738), .YC(n1735), .YS(n1736) );
  HAX1 U1149 ( .A(n2234), .B(n1756), .YC(n1737), .YS(n1738) );
  FAX1 U1150 ( .A(n2235), .B(n2203), .C(n2171), .YC(n1739), .YS(n1740) );
  HAX1 U1151 ( .A(n2236), .B(n2204), .YC(n1741), .YS(n1742) );
  NOR2X1 U1152 ( .A(n2239), .B(n383), .Y(n1759) );
  NOR2X1 U1153 ( .A(n2240), .B(n383), .Y(n918) );
  NOR2X1 U1154 ( .A(n2241), .B(n383), .Y(n1760) );
  NOR2X1 U1155 ( .A(n2242), .B(n383), .Y(n960) );
  NOR2X1 U1156 ( .A(n2243), .B(n383), .Y(n1761) );
  NOR2X1 U1157 ( .A(n2244), .B(n383), .Y(n1006) );
  NOR2X1 U1158 ( .A(n2245), .B(n383), .Y(n1762) );
  NOR2X1 U1159 ( .A(n2972), .B(n383), .Y(n1056) );
  NOR2X1 U1160 ( .A(n2992), .B(n383), .Y(n1763) );
  NOR2X1 U1161 ( .A(n2248), .B(n383), .Y(n1110) );
  NOR2X1 U1162 ( .A(n2966), .B(n383), .Y(n1764) );
  NOR2X1 U1163 ( .A(n2250), .B(n383), .Y(n1168) );
  NOR2X1 U1164 ( .A(n2251), .B(n383), .Y(n1765) );
  NOR2X1 U1165 ( .A(n2252), .B(n383), .Y(n1766) );
  NOR2X1 U1166 ( .A(n2984), .B(n383), .Y(n1230) );
  INVX2 U1178 ( .A(b[4]), .Y(n2250) );
  INVX2 U1180 ( .A(n439), .Y(n2252) );
  OAI22X1 U1182 ( .A(n382), .B(n2272), .C(n2796), .D(n432), .Y(n1743) );
  OAI22X1 U1183 ( .A(n2254), .B(n381), .C(n2255), .D(n431), .Y(n1768) );
  OAI22X1 U1184 ( .A(n2255), .B(n381), .C(n2256), .D(n431), .Y(n1769) );
  OAI22X1 U1185 ( .A(n2256), .B(n381), .C(n2257), .D(n431), .Y(n1770) );
  OAI22X1 U1186 ( .A(n2257), .B(n381), .C(n2258), .D(n431), .Y(n1771) );
  OAI22X1 U1187 ( .A(n2258), .B(n381), .C(n2259), .D(n431), .Y(n1772) );
  OAI22X1 U1188 ( .A(n2259), .B(n381), .C(n2260), .D(n431), .Y(n1773) );
  OAI22X1 U1189 ( .A(n2260), .B(n380), .C(n2261), .D(n431), .Y(n1774) );
  OAI22X1 U1190 ( .A(n2261), .B(n380), .C(n2262), .D(n430), .Y(n1775) );
  OAI22X1 U1191 ( .A(n2262), .B(n380), .C(n2263), .D(n430), .Y(n1776) );
  OAI22X1 U1192 ( .A(n2263), .B(n380), .C(n2264), .D(n430), .Y(n1777) );
  OAI22X1 U1193 ( .A(n2264), .B(n380), .C(n2265), .D(n430), .Y(n1778) );
  OAI22X1 U1194 ( .A(n2265), .B(n380), .C(n2266), .D(n430), .Y(n1779) );
  OAI22X1 U1195 ( .A(n2266), .B(n380), .C(n2267), .D(n430), .Y(n1780) );
  OAI22X1 U1196 ( .A(n2267), .B(n380), .C(n2268), .D(n430), .Y(n1781) );
  OAI22X1 U1197 ( .A(n2268), .B(n380), .C(n2269), .D(n430), .Y(n1782) );
  OAI22X1 U1198 ( .A(n2269), .B(n380), .C(n2270), .D(n430), .Y(n1783) );
  OAI22X1 U1199 ( .A(n2270), .B(n380), .C(n2271), .D(n430), .Y(n1784) );
  XNOR2X1 U1200 ( .A(n333), .B(n469), .Y(n2254) );
  XNOR2X1 U1201 ( .A(n333), .B(n467), .Y(n2255) );
  XNOR2X1 U1202 ( .A(n333), .B(n2983), .Y(n2256) );
  XNOR2X1 U1203 ( .A(n333), .B(n2962), .Y(n2257) );
  XNOR2X1 U1204 ( .A(n333), .B(n2976), .Y(n2258) );
  XNOR2X1 U1205 ( .A(n333), .B(n2991), .Y(n2259) );
  XNOR2X1 U1206 ( .A(n333), .B(n2965), .Y(n2260) );
  XNOR2X1 U1207 ( .A(n333), .B(n2978), .Y(n2261) );
  XNOR2X1 U1208 ( .A(n333), .B(n2970), .Y(n2262) );
  XNOR2X1 U1209 ( .A(n332), .B(n2973), .Y(n2263) );
  XNOR2X1 U1210 ( .A(n332), .B(n2994), .Y(n2264) );
  XNOR2X1 U1211 ( .A(n332), .B(n2960), .Y(n2265) );
  XNOR2X1 U1212 ( .A(n332), .B(n2968), .Y(n2266) );
  XNOR2X1 U1213 ( .A(n332), .B(n2996), .Y(n2267) );
  XNOR2X1 U1214 ( .A(n332), .B(n2981), .Y(n2268) );
  XNOR2X1 U1215 ( .A(n332), .B(n439), .Y(n2269) );
  XNOR2X1 U1216 ( .A(n332), .B(n2911), .Y(n2270) );
  XNOR2X1 U1217 ( .A(n332), .B(n2998), .Y(n2271) );
  OAI22X1 U1218 ( .A(n379), .B(n2293), .C(n2797), .D(n429), .Y(n1744) );
  OAI22X1 U1219 ( .A(n2273), .B(n378), .C(n2274), .D(n428), .Y(n1786) );
  OAI22X1 U1220 ( .A(n2274), .B(n378), .C(n2275), .D(n428), .Y(n1787) );
  OAI22X1 U1221 ( .A(n2275), .B(n378), .C(n2276), .D(n428), .Y(n1788) );
  OAI22X1 U1222 ( .A(n2276), .B(n378), .C(n2277), .D(n428), .Y(n1789) );
  OAI22X1 U1223 ( .A(n2277), .B(n378), .C(n2278), .D(n428), .Y(n1790) );
  OAI22X1 U1224 ( .A(n2278), .B(n378), .C(n2279), .D(n428), .Y(n1791) );
  OAI22X1 U1225 ( .A(n2279), .B(n378), .C(n2280), .D(n428), .Y(n1792) );
  OAI22X1 U1226 ( .A(n2280), .B(n378), .C(n2281), .D(n428), .Y(n1793) );
  OAI22X1 U1227 ( .A(n2281), .B(n377), .C(n2282), .D(n428), .Y(n1794) );
  OAI22X1 U1228 ( .A(n2282), .B(n377), .C(n2283), .D(n427), .Y(n1795) );
  OAI22X1 U1229 ( .A(n2283), .B(n377), .C(n2284), .D(n427), .Y(n1796) );
  OAI22X1 U1230 ( .A(n2284), .B(n377), .C(n2285), .D(n427), .Y(n1797) );
  OAI22X1 U1231 ( .A(n2285), .B(n377), .C(n2286), .D(n427), .Y(n1798) );
  OAI22X1 U1232 ( .A(n2286), .B(n377), .C(n2287), .D(n427), .Y(n1799) );
  OAI22X1 U1233 ( .A(n2287), .B(n377), .C(n2288), .D(n427), .Y(n1800) );
  OAI22X1 U1234 ( .A(n2288), .B(n377), .C(n2289), .D(n427), .Y(n1801) );
  OAI22X1 U1235 ( .A(n2289), .B(n377), .C(n2290), .D(n427), .Y(n1802) );
  OAI22X1 U1236 ( .A(n2290), .B(n377), .C(n2291), .D(n427), .Y(n1803) );
  OAI22X1 U1237 ( .A(n2291), .B(n377), .C(n2292), .D(n427), .Y(n1804) );
  XNOR2X1 U1238 ( .A(n330), .B(n473), .Y(n2273) );
  XNOR2X1 U1239 ( .A(n330), .B(n471), .Y(n2274) );
  XNOR2X1 U1240 ( .A(n330), .B(n469), .Y(n2275) );
  XNOR2X1 U1241 ( .A(n330), .B(n467), .Y(n2276) );
  XNOR2X1 U1242 ( .A(n330), .B(n2982), .Y(n2277) );
  XNOR2X1 U1243 ( .A(n330), .B(n2961), .Y(n2278) );
  XNOR2X1 U1244 ( .A(n330), .B(n2975), .Y(n2279) );
  XNOR2X1 U1245 ( .A(n330), .B(n2991), .Y(n2280) );
  XNOR2X1 U1246 ( .A(n330), .B(n2964), .Y(n2281) );
  XNOR2X1 U1247 ( .A(n330), .B(n2978), .Y(n2282) );
  XNOR2X1 U1248 ( .A(n330), .B(n2971), .Y(n2283) );
  XNOR2X1 U1249 ( .A(n329), .B(n2973), .Y(n2284) );
  XNOR2X1 U1250 ( .A(n329), .B(n2993), .Y(n2285) );
  XNOR2X1 U1251 ( .A(n329), .B(n2959), .Y(n2286) );
  XNOR2X1 U1252 ( .A(n329), .B(n2940), .Y(n2287) );
  XNOR2X1 U1253 ( .A(n329), .B(n2996), .Y(n2288) );
  XNOR2X1 U1254 ( .A(n329), .B(n2980), .Y(n2289) );
  XNOR2X1 U1255 ( .A(n329), .B(n439), .Y(n2290) );
  XNOR2X1 U1256 ( .A(n329), .B(n2911), .Y(n2291) );
  XNOR2X1 U1257 ( .A(n329), .B(n2944), .Y(n2292) );
  OAI22X1 U1258 ( .A(n376), .B(n2316), .C(n2798), .D(n426), .Y(n1745) );
  OAI22X1 U1259 ( .A(n2294), .B(n375), .C(n2295), .D(n425), .Y(n1806) );
  OAI22X1 U1260 ( .A(n2295), .B(n375), .C(n2296), .D(n425), .Y(n1807) );
  OAI22X1 U1261 ( .A(n2296), .B(n375), .C(n2297), .D(n425), .Y(n1808) );
  OAI22X1 U1262 ( .A(n2297), .B(n375), .C(n2298), .D(n425), .Y(n1809) );
  OAI22X1 U1263 ( .A(n2298), .B(n375), .C(n2299), .D(n425), .Y(n1810) );
  OAI22X1 U1264 ( .A(n2299), .B(n375), .C(n2300), .D(n425), .Y(n1811) );
  OAI22X1 U1265 ( .A(n2300), .B(n375), .C(n2301), .D(n425), .Y(n1812) );
  OAI22X1 U1266 ( .A(n2301), .B(n375), .C(n2302), .D(n425), .Y(n1813) );
  OAI22X1 U1267 ( .A(n2302), .B(n375), .C(n2303), .D(n425), .Y(n1814) );
  OAI22X1 U1268 ( .A(n2303), .B(n375), .C(n2304), .D(n425), .Y(n1815) );
  OAI22X1 U1269 ( .A(n2304), .B(n374), .C(n2305), .D(n425), .Y(n1816) );
  OAI22X1 U1270 ( .A(n2305), .B(n374), .C(n2306), .D(n424), .Y(n1817) );
  OAI22X1 U1271 ( .A(n2306), .B(n374), .C(n2307), .D(n424), .Y(n1818) );
  OAI22X1 U1272 ( .A(n2307), .B(n374), .C(n2308), .D(n424), .Y(n1819) );
  OAI22X1 U1273 ( .A(n2308), .B(n374), .C(n2309), .D(n424), .Y(n1820) );
  OAI22X1 U1274 ( .A(n2309), .B(n374), .C(n2310), .D(n424), .Y(n1821) );
  OAI22X1 U1275 ( .A(n2310), .B(n374), .C(n2311), .D(n424), .Y(n1822) );
  OAI22X1 U1276 ( .A(n2311), .B(n374), .C(n2312), .D(n424), .Y(n1823) );
  OAI22X1 U1277 ( .A(n2312), .B(n374), .C(n2313), .D(n424), .Y(n1824) );
  OAI22X1 U1278 ( .A(n2313), .B(n374), .C(n2314), .D(n424), .Y(n1825) );
  OAI22X1 U1279 ( .A(n2314), .B(n374), .C(n2315), .D(n424), .Y(n1826) );
  XNOR2X1 U1280 ( .A(n328), .B(n477), .Y(n2294) );
  XNOR2X1 U1281 ( .A(n327), .B(n475), .Y(n2295) );
  XNOR2X1 U1282 ( .A(n327), .B(n473), .Y(n2296) );
  XNOR2X1 U1283 ( .A(n327), .B(n471), .Y(n2297) );
  XNOR2X1 U1284 ( .A(n327), .B(n469), .Y(n2298) );
  XNOR2X1 U1285 ( .A(n327), .B(n467), .Y(n2299) );
  XNOR2X1 U1286 ( .A(n327), .B(n2983), .Y(n2300) );
  XNOR2X1 U1287 ( .A(n327), .B(n2962), .Y(n2301) );
  XNOR2X1 U1288 ( .A(n327), .B(n2976), .Y(n2302) );
  XNOR2X1 U1289 ( .A(n327), .B(n2991), .Y(n2303) );
  XNOR2X1 U1290 ( .A(n327), .B(n2965), .Y(n2304) );
  XNOR2X1 U1291 ( .A(n327), .B(n2978), .Y(n2305) );
  XNOR2X1 U1292 ( .A(n327), .B(n2971), .Y(n2306) );
  XNOR2X1 U1293 ( .A(n326), .B(n2973), .Y(n2307) );
  XNOR2X1 U1294 ( .A(n326), .B(n2994), .Y(n2308) );
  XNOR2X1 U1295 ( .A(n326), .B(n2960), .Y(n2309) );
  XNOR2X1 U1296 ( .A(n326), .B(n2968), .Y(n2310) );
  XNOR2X1 U1297 ( .A(n326), .B(n2996), .Y(n2311) );
  XNOR2X1 U1298 ( .A(n326), .B(n2981), .Y(n2312) );
  XNOR2X1 U1299 ( .A(n326), .B(n439), .Y(n2313) );
  XNOR2X1 U1300 ( .A(n326), .B(n2911), .Y(n2314) );
  XNOR2X1 U1301 ( .A(n326), .B(n2913), .Y(n2315) );
  OAI22X1 U1302 ( .A(n373), .B(n2341), .C(n2799), .D(n423), .Y(n1746) );
  OAI22X1 U1303 ( .A(n2317), .B(n372), .C(n2318), .D(n423), .Y(n1828) );
  OAI22X1 U1304 ( .A(n2318), .B(n372), .C(n2319), .D(n422), .Y(n1829) );
  OAI22X1 U1305 ( .A(n2319), .B(n372), .C(n2320), .D(n422), .Y(n1830) );
  OAI22X1 U1306 ( .A(n2320), .B(n372), .C(n2321), .D(n422), .Y(n1831) );
  OAI22X1 U1307 ( .A(n2321), .B(n372), .C(n2322), .D(n422), .Y(n1832) );
  OAI22X1 U1308 ( .A(n2322), .B(n372), .C(n2323), .D(n422), .Y(n1833) );
  OAI22X1 U1309 ( .A(n2323), .B(n372), .C(n2324), .D(n422), .Y(n1834) );
  OAI22X1 U1310 ( .A(n2324), .B(n372), .C(n2325), .D(n422), .Y(n1835) );
  OAI22X1 U1311 ( .A(n2325), .B(n372), .C(n2326), .D(n422), .Y(n1836) );
  OAI22X1 U1312 ( .A(n2326), .B(n372), .C(n2327), .D(n422), .Y(n1837) );
  OAI22X1 U1313 ( .A(n2327), .B(n372), .C(n2328), .D(n422), .Y(n1838) );
  OAI22X1 U1314 ( .A(n2328), .B(n372), .C(n2329), .D(n422), .Y(n1839) );
  OAI22X1 U1315 ( .A(n2329), .B(n371), .C(n2330), .D(n422), .Y(n1840) );
  OAI22X1 U1316 ( .A(n2330), .B(n371), .C(n2331), .D(n421), .Y(n1841) );
  OAI22X1 U1317 ( .A(n2331), .B(n371), .C(n2332), .D(n421), .Y(n1842) );
  OAI22X1 U1318 ( .A(n2332), .B(n371), .C(n2333), .D(n421), .Y(n1843) );
  OAI22X1 U1319 ( .A(n2333), .B(n371), .C(n2334), .D(n421), .Y(n1844) );
  OAI22X1 U1320 ( .A(n2334), .B(n371), .C(n2335), .D(n421), .Y(n1845) );
  OAI22X1 U1321 ( .A(n2335), .B(n371), .C(n2336), .D(n421), .Y(n1846) );
  OAI22X1 U1322 ( .A(n2336), .B(n371), .C(n2337), .D(n421), .Y(n1847) );
  OAI22X1 U1323 ( .A(n2337), .B(n371), .C(n2338), .D(n421), .Y(n1848) );
  OAI22X1 U1324 ( .A(n2338), .B(n371), .C(n2339), .D(n421), .Y(n1849) );
  OAI22X1 U1325 ( .A(n2339), .B(n371), .C(n2340), .D(n421), .Y(n1850) );
  XNOR2X1 U1326 ( .A(n325), .B(n481), .Y(n2317) );
  XNOR2X1 U1327 ( .A(n325), .B(n479), .Y(n2318) );
  XNOR2X1 U1328 ( .A(n325), .B(n477), .Y(n2319) );
  XNOR2X1 U1329 ( .A(n324), .B(n475), .Y(n2320) );
  XNOR2X1 U1330 ( .A(n324), .B(n473), .Y(n2321) );
  XNOR2X1 U1331 ( .A(n324), .B(n471), .Y(n2322) );
  XNOR2X1 U1332 ( .A(n324), .B(n469), .Y(n2323) );
  XNOR2X1 U1333 ( .A(n324), .B(n467), .Y(n2324) );
  XNOR2X1 U1334 ( .A(n324), .B(n2982), .Y(n2325) );
  XNOR2X1 U1335 ( .A(n324), .B(n2961), .Y(n2326) );
  XNOR2X1 U1336 ( .A(n324), .B(n2975), .Y(n2327) );
  XNOR2X1 U1337 ( .A(n324), .B(n2991), .Y(n2328) );
  XNOR2X1 U1338 ( .A(n324), .B(n2964), .Y(n2329) );
  XNOR2X1 U1339 ( .A(n324), .B(n2978), .Y(n2330) );
  XNOR2X1 U1340 ( .A(n324), .B(n2970), .Y(n2331) );
  XNOR2X1 U1341 ( .A(n323), .B(n2973), .Y(n2332) );
  XNOR2X1 U1342 ( .A(n323), .B(n2993), .Y(n2333) );
  XNOR2X1 U1343 ( .A(n323), .B(n2959), .Y(n2334) );
  XNOR2X1 U1344 ( .A(n323), .B(n2968), .Y(n2335) );
  XNOR2X1 U1345 ( .A(n323), .B(n2996), .Y(n2336) );
  XNOR2X1 U1346 ( .A(n323), .B(n2980), .Y(n2337) );
  XNOR2X1 U1347 ( .A(n323), .B(n439), .Y(n2338) );
  XNOR2X1 U1348 ( .A(n323), .B(n2911), .Y(n2339) );
  XNOR2X1 U1349 ( .A(n323), .B(n2941), .Y(n2340) );
  OAI22X1 U1350 ( .A(n370), .B(n2368), .C(n2800), .D(n420), .Y(n1747) );
  OAI22X1 U1351 ( .A(n2342), .B(n370), .C(n2343), .D(n420), .Y(n1852) );
  OAI22X1 U1352 ( .A(n2343), .B(n370), .C(n2344), .D(n420), .Y(n1853) );
  OAI22X1 U1353 ( .A(n2344), .B(n369), .C(n2345), .D(n420), .Y(n1854) );
  OAI22X1 U1354 ( .A(n2345), .B(n369), .C(n2346), .D(n419), .Y(n1855) );
  OAI22X1 U1355 ( .A(n2346), .B(n369), .C(n2347), .D(n419), .Y(n1856) );
  OAI22X1 U1356 ( .A(n2347), .B(n369), .C(n2348), .D(n419), .Y(n1857) );
  OAI22X1 U1357 ( .A(n2348), .B(n369), .C(n2349), .D(n419), .Y(n1858) );
  OAI22X1 U1358 ( .A(n2349), .B(n369), .C(n2350), .D(n419), .Y(n1859) );
  OAI22X1 U1359 ( .A(n2350), .B(n369), .C(n2351), .D(n419), .Y(n1860) );
  OAI22X1 U1360 ( .A(n2351), .B(n369), .C(n2352), .D(n419), .Y(n1861) );
  OAI22X1 U1361 ( .A(n2352), .B(n369), .C(n2353), .D(n419), .Y(n1862) );
  OAI22X1 U1362 ( .A(n2353), .B(n369), .C(n2354), .D(n419), .Y(n1863) );
  OAI22X1 U1363 ( .A(n2354), .B(n369), .C(n2355), .D(n419), .Y(n1864) );
  OAI22X1 U1364 ( .A(n2355), .B(n369), .C(n2356), .D(n419), .Y(n1865) );
  OAI22X1 U1365 ( .A(n2356), .B(n368), .C(n2357), .D(n419), .Y(n1866) );
  OAI22X1 U1366 ( .A(n2357), .B(n368), .C(n2358), .D(n418), .Y(n1867) );
  OAI22X1 U1367 ( .A(n2358), .B(n368), .C(n2359), .D(n418), .Y(n1868) );
  OAI22X1 U1368 ( .A(n2359), .B(n368), .C(n2360), .D(n418), .Y(n1869) );
  OAI22X1 U1369 ( .A(n2360), .B(n368), .C(n2361), .D(n418), .Y(n1870) );
  OAI22X1 U1370 ( .A(n2361), .B(n368), .C(n2362), .D(n418), .Y(n1871) );
  OAI22X1 U1371 ( .A(n2362), .B(n368), .C(n2363), .D(n418), .Y(n1872) );
  OAI22X1 U1372 ( .A(n2363), .B(n368), .C(n2364), .D(n418), .Y(n1873) );
  OAI22X1 U1373 ( .A(n2364), .B(n368), .C(n2365), .D(n418), .Y(n1874) );
  OAI22X1 U1374 ( .A(n2365), .B(n368), .C(n2366), .D(n418), .Y(n1875) );
  OAI22X1 U1375 ( .A(n2366), .B(n368), .C(n2367), .D(n418), .Y(n1876) );
  XNOR2X1 U1376 ( .A(n322), .B(n485), .Y(n2342) );
  XNOR2X1 U1377 ( .A(n322), .B(n483), .Y(n2343) );
  XNOR2X1 U1378 ( .A(n322), .B(n481), .Y(n2344) );
  XNOR2X1 U1379 ( .A(n322), .B(n479), .Y(n2345) );
  XNOR2X1 U1380 ( .A(n322), .B(n477), .Y(n2346) );
  XNOR2X1 U1381 ( .A(n321), .B(n475), .Y(n2347) );
  XNOR2X1 U1382 ( .A(n321), .B(n473), .Y(n2348) );
  XNOR2X1 U1383 ( .A(n321), .B(n471), .Y(n2349) );
  XNOR2X1 U1384 ( .A(n321), .B(n469), .Y(n2350) );
  XNOR2X1 U1385 ( .A(n321), .B(n467), .Y(n2351) );
  XNOR2X1 U1386 ( .A(n321), .B(n2983), .Y(n2352) );
  XNOR2X1 U1387 ( .A(n321), .B(n2962), .Y(n2353) );
  XNOR2X1 U1388 ( .A(n321), .B(n2976), .Y(n2354) );
  XNOR2X1 U1389 ( .A(n321), .B(n2991), .Y(n2355) );
  XNOR2X1 U1390 ( .A(n321), .B(n2965), .Y(n2356) );
  XNOR2X1 U1391 ( .A(n321), .B(n2978), .Y(n2357) );
  XNOR2X1 U1392 ( .A(n321), .B(n2971), .Y(n2358) );
  XNOR2X1 U1393 ( .A(n320), .B(n2973), .Y(n2359) );
  XNOR2X1 U1394 ( .A(n320), .B(n2994), .Y(n2360) );
  XNOR2X1 U1395 ( .A(n320), .B(n2960), .Y(n2361) );
  XNOR2X1 U1396 ( .A(n320), .B(n2940), .Y(n2362) );
  XNOR2X1 U1397 ( .A(n320), .B(n2996), .Y(n2363) );
  XNOR2X1 U1398 ( .A(n320), .B(n2981), .Y(n2364) );
  XNOR2X1 U1399 ( .A(n320), .B(n439), .Y(n2365) );
  XNOR2X1 U1400 ( .A(n320), .B(n2911), .Y(n2366) );
  XNOR2X1 U1401 ( .A(n320), .B(n2998), .Y(n2367) );
  OAI22X1 U1402 ( .A(n367), .B(n2397), .C(n2801), .D(n417), .Y(n1748) );
  OAI22X1 U1403 ( .A(n2369), .B(n367), .C(n2370), .D(n417), .Y(n1878) );
  OAI22X1 U1404 ( .A(n2370), .B(n367), .C(n2371), .D(n417), .Y(n1879) );
  OAI22X1 U1405 ( .A(n2371), .B(n367), .C(n2372), .D(n417), .Y(n1880) );
  OAI22X1 U1406 ( .A(n2372), .B(n367), .C(n2373), .D(n417), .Y(n1881) );
  OAI22X1 U1407 ( .A(n2373), .B(n366), .C(n2374), .D(n417), .Y(n1882) );
  OAI22X1 U1408 ( .A(n2374), .B(n366), .C(n2375), .D(n416), .Y(n1883) );
  OAI22X1 U1409 ( .A(n2375), .B(n366), .C(n2376), .D(n416), .Y(n1884) );
  OAI22X1 U1410 ( .A(n2376), .B(n366), .C(n2377), .D(n416), .Y(n1885) );
  OAI22X1 U1411 ( .A(n2377), .B(n366), .C(n2378), .D(n416), .Y(n1886) );
  OAI22X1 U1412 ( .A(n2378), .B(n366), .C(n2379), .D(n416), .Y(n1887) );
  OAI22X1 U1413 ( .A(n2379), .B(n366), .C(n2380), .D(n416), .Y(n1888) );
  OAI22X1 U1414 ( .A(n2380), .B(n366), .C(n2381), .D(n416), .Y(n1889) );
  OAI22X1 U1415 ( .A(n2381), .B(n366), .C(n2382), .D(n416), .Y(n1890) );
  OAI22X1 U1416 ( .A(n2382), .B(n366), .C(n2383), .D(n416), .Y(n1891) );
  OAI22X1 U1417 ( .A(n2383), .B(n366), .C(n2384), .D(n416), .Y(n1892) );
  OAI22X1 U1418 ( .A(n2384), .B(n366), .C(n2385), .D(n416), .Y(n1893) );
  OAI22X1 U1419 ( .A(n2385), .B(n365), .C(n2386), .D(n416), .Y(n1894) );
  OAI22X1 U1420 ( .A(n2386), .B(n365), .C(n2387), .D(n415), .Y(n1895) );
  OAI22X1 U1421 ( .A(n2387), .B(n365), .C(n2388), .D(n415), .Y(n1896) );
  OAI22X1 U1422 ( .A(n2388), .B(n365), .C(n2389), .D(n415), .Y(n1897) );
  OAI22X1 U1423 ( .A(n2389), .B(n365), .C(n2390), .D(n415), .Y(n1898) );
  OAI22X1 U1424 ( .A(n2390), .B(n365), .C(n2391), .D(n415), .Y(n1899) );
  OAI22X1 U1425 ( .A(n2391), .B(n365), .C(n2392), .D(n415), .Y(n1900) );
  OAI22X1 U1426 ( .A(n2392), .B(n365), .C(n2393), .D(n415), .Y(n1901) );
  OAI22X1 U1427 ( .A(n2393), .B(n365), .C(n2394), .D(n415), .Y(n1902) );
  OAI22X1 U1428 ( .A(n2394), .B(n365), .C(n2395), .D(n415), .Y(n1903) );
  OAI22X1 U1429 ( .A(n2395), .B(n365), .C(n2396), .D(n415), .Y(n1904) );
  XNOR2X1 U1430 ( .A(n319), .B(b[27]), .Y(n2369) );
  XNOR2X1 U1431 ( .A(n319), .B(b[26]), .Y(n2370) );
  XNOR2X1 U1432 ( .A(n319), .B(n485), .Y(n2371) );
  XNOR2X1 U1433 ( .A(n319), .B(n483), .Y(n2372) );
  XNOR2X1 U1434 ( .A(n319), .B(n481), .Y(n2373) );
  XNOR2X1 U1435 ( .A(n319), .B(n479), .Y(n2374) );
  XNOR2X1 U1436 ( .A(n319), .B(n477), .Y(n2375) );
  XNOR2X1 U1437 ( .A(n318), .B(n475), .Y(n2376) );
  XNOR2X1 U1438 ( .A(n318), .B(n473), .Y(n2377) );
  XNOR2X1 U1439 ( .A(n318), .B(n471), .Y(n2378) );
  XNOR2X1 U1440 ( .A(n318), .B(n469), .Y(n2379) );
  XNOR2X1 U1441 ( .A(n318), .B(n467), .Y(n2380) );
  XNOR2X1 U1442 ( .A(n318), .B(n2982), .Y(n2381) );
  XNOR2X1 U1443 ( .A(n318), .B(n2961), .Y(n2382) );
  XNOR2X1 U1444 ( .A(n318), .B(n2975), .Y(n2383) );
  XNOR2X1 U1445 ( .A(n318), .B(n2991), .Y(n2384) );
  XNOR2X1 U1446 ( .A(n318), .B(n2964), .Y(n2385) );
  XNOR2X1 U1447 ( .A(n318), .B(n2978), .Y(n2386) );
  XNOR2X1 U1448 ( .A(n318), .B(n2970), .Y(n2387) );
  XNOR2X1 U1449 ( .A(n317), .B(n2973), .Y(n2388) );
  XNOR2X1 U1450 ( .A(n317), .B(n2993), .Y(n2389) );
  XNOR2X1 U1451 ( .A(n317), .B(n2959), .Y(n2390) );
  XNOR2X1 U1452 ( .A(n317), .B(n2968), .Y(n2391) );
  XNOR2X1 U1453 ( .A(n317), .B(n2996), .Y(n2392) );
  XNOR2X1 U1454 ( .A(n317), .B(n2980), .Y(n2393) );
  XNOR2X1 U1455 ( .A(n317), .B(n439), .Y(n2394) );
  XNOR2X1 U1456 ( .A(n317), .B(n2911), .Y(n2395) );
  XNOR2X1 U1457 ( .A(n317), .B(n2944), .Y(n2396) );
  OAI22X1 U1458 ( .A(n364), .B(n2428), .C(n2802), .D(n414), .Y(n1749) );
  OAI22X1 U1459 ( .A(n2398), .B(n364), .C(n2399), .D(n414), .Y(n1906) );
  OAI22X1 U1460 ( .A(n2399), .B(n364), .C(n2400), .D(n414), .Y(n1907) );
  OAI22X1 U1461 ( .A(n2400), .B(n364), .C(n2401), .D(n414), .Y(n1908) );
  OAI22X1 U1462 ( .A(n2401), .B(n364), .C(n2402), .D(n414), .Y(n1909) );
  OAI22X1 U1463 ( .A(n2402), .B(n364), .C(n2403), .D(n414), .Y(n1910) );
  OAI22X1 U1464 ( .A(n2403), .B(n364), .C(n2404), .D(n414), .Y(n1911) );
  OAI22X1 U1465 ( .A(n2404), .B(n363), .C(n2405), .D(n414), .Y(n1912) );
  OAI22X1 U1466 ( .A(n2405), .B(n363), .C(n2406), .D(n413), .Y(n1913) );
  OAI22X1 U1467 ( .A(n2406), .B(n363), .C(n2407), .D(n413), .Y(n1914) );
  OAI22X1 U1468 ( .A(n2407), .B(n363), .C(n2408), .D(n413), .Y(n1915) );
  OAI22X1 U1469 ( .A(n2408), .B(n363), .C(n2409), .D(n413), .Y(n1916) );
  OAI22X1 U1470 ( .A(n2409), .B(n363), .C(n2410), .D(n413), .Y(n1917) );
  OAI22X1 U1471 ( .A(n2410), .B(n363), .C(n2411), .D(n413), .Y(n1918) );
  OAI22X1 U1472 ( .A(n2411), .B(n363), .C(n2412), .D(n413), .Y(n1919) );
  OAI22X1 U1473 ( .A(n2412), .B(n363), .C(n2413), .D(n413), .Y(n1920) );
  OAI22X1 U1474 ( .A(n2413), .B(n363), .C(n2414), .D(n413), .Y(n1921) );
  OAI22X1 U1475 ( .A(n2414), .B(n363), .C(n2415), .D(n413), .Y(n1922) );
  OAI22X1 U1476 ( .A(n2415), .B(n363), .C(n2416), .D(n413), .Y(n1923) );
  OAI22X1 U1477 ( .A(n2416), .B(n362), .C(n2417), .D(n413), .Y(n1924) );
  OAI22X1 U1478 ( .A(n2417), .B(n362), .C(n2418), .D(n412), .Y(n1925) );
  OAI22X1 U1479 ( .A(n2418), .B(n362), .C(n2419), .D(n412), .Y(n1926) );
  OAI22X1 U1480 ( .A(n2419), .B(n362), .C(n2420), .D(n412), .Y(n1927) );
  OAI22X1 U1481 ( .A(n2420), .B(n362), .C(n2421), .D(n412), .Y(n1928) );
  OAI22X1 U1482 ( .A(n2421), .B(n362), .C(n2422), .D(n412), .Y(n1929) );
  OAI22X1 U1483 ( .A(n2422), .B(n362), .C(n2423), .D(n412), .Y(n1930) );
  OAI22X1 U1484 ( .A(n2423), .B(n362), .C(n2424), .D(n412), .Y(n1931) );
  OAI22X1 U1485 ( .A(n2424), .B(n362), .C(n2425), .D(n412), .Y(n1932) );
  OAI22X1 U1486 ( .A(n2425), .B(n362), .C(n2426), .D(n412), .Y(n1933) );
  OAI22X1 U1487 ( .A(n2426), .B(n362), .C(n2427), .D(n412), .Y(n1934) );
  XNOR2X1 U1488 ( .A(n316), .B(b[29]), .Y(n2398) );
  XNOR2X1 U1489 ( .A(n316), .B(b[28]), .Y(n2399) );
  XNOR2X1 U1490 ( .A(n316), .B(b[27]), .Y(n2400) );
  XNOR2X1 U1491 ( .A(n316), .B(b[26]), .Y(n2401) );
  XNOR2X1 U1492 ( .A(n316), .B(n485), .Y(n2402) );
  XNOR2X1 U1493 ( .A(n316), .B(n483), .Y(n2403) );
  XNOR2X1 U1494 ( .A(n316), .B(n481), .Y(n2404) );
  XNOR2X1 U1495 ( .A(n316), .B(n479), .Y(n2405) );
  XNOR2X1 U1496 ( .A(n316), .B(n477), .Y(n2406) );
  XNOR2X1 U1497 ( .A(n315), .B(n475), .Y(n2407) );
  XNOR2X1 U1498 ( .A(n315), .B(n473), .Y(n2408) );
  XNOR2X1 U1499 ( .A(n315), .B(n471), .Y(n2409) );
  XNOR2X1 U1500 ( .A(n315), .B(n469), .Y(n2410) );
  XNOR2X1 U1501 ( .A(n315), .B(n467), .Y(n2411) );
  XNOR2X1 U1502 ( .A(n315), .B(n2983), .Y(n2412) );
  XNOR2X1 U1503 ( .A(n315), .B(n2962), .Y(n2413) );
  XNOR2X1 U1504 ( .A(n315), .B(n2976), .Y(n2414) );
  XNOR2X1 U1505 ( .A(n315), .B(n2991), .Y(n2415) );
  XNOR2X1 U1506 ( .A(n315), .B(n2965), .Y(n2416) );
  XNOR2X1 U1507 ( .A(n315), .B(n2978), .Y(n2417) );
  XNOR2X1 U1508 ( .A(n315), .B(n2971), .Y(n2418) );
  XNOR2X1 U1509 ( .A(n314), .B(n2973), .Y(n2419) );
  XNOR2X1 U1510 ( .A(n314), .B(n2994), .Y(n2420) );
  XNOR2X1 U1511 ( .A(n314), .B(n2960), .Y(n2421) );
  XNOR2X1 U1512 ( .A(n314), .B(n2968), .Y(n2422) );
  XNOR2X1 U1513 ( .A(n314), .B(n2996), .Y(n2423) );
  XNOR2X1 U1514 ( .A(n314), .B(n2981), .Y(n2424) );
  XNOR2X1 U1515 ( .A(n314), .B(n439), .Y(n2425) );
  XNOR2X1 U1516 ( .A(n314), .B(n2911), .Y(n2426) );
  XNOR2X1 U1517 ( .A(n314), .B(n2913), .Y(n2427) );
  OAI22X1 U1518 ( .A(n361), .B(n2461), .C(n2803), .D(n411), .Y(n1750) );
  OAI22X1 U1519 ( .A(n2429), .B(n361), .C(n2430), .D(n411), .Y(n1936) );
  OAI22X1 U1520 ( .A(n2430), .B(n361), .C(n2431), .D(n411), .Y(n1937) );
  OAI22X1 U1521 ( .A(n2431), .B(n361), .C(n2432), .D(n411), .Y(n1938) );
  OAI22X1 U1522 ( .A(n2432), .B(n361), .C(n2433), .D(n411), .Y(n1939) );
  OAI22X1 U1523 ( .A(n2433), .B(n361), .C(n2434), .D(n411), .Y(n1940) );
  OAI22X1 U1524 ( .A(n2434), .B(n361), .C(n2435), .D(n411), .Y(n1941) );
  OAI22X1 U1525 ( .A(n2435), .B(n361), .C(n2436), .D(n411), .Y(n1942) );
  OAI22X1 U1526 ( .A(n2436), .B(n361), .C(n2437), .D(n411), .Y(n1943) );
  OAI22X1 U1527 ( .A(n2437), .B(n360), .C(n2438), .D(n411), .Y(n1944) );
  OAI22X1 U1528 ( .A(n2438), .B(n360), .C(n2439), .D(n410), .Y(n1945) );
  OAI22X1 U1529 ( .A(n2439), .B(n360), .C(n2440), .D(n410), .Y(n1946) );
  OAI22X1 U1530 ( .A(n2440), .B(n360), .C(n2441), .D(n410), .Y(n1947) );
  OAI22X1 U1531 ( .A(n2441), .B(n360), .C(n2442), .D(n410), .Y(n1948) );
  OAI22X1 U1532 ( .A(n2442), .B(n360), .C(n2443), .D(n410), .Y(n1949) );
  OAI22X1 U1533 ( .A(n2443), .B(n360), .C(n2444), .D(n410), .Y(n1950) );
  OAI22X1 U1534 ( .A(n2444), .B(n360), .C(n2445), .D(n410), .Y(n1951) );
  OAI22X1 U1535 ( .A(n2445), .B(n360), .C(n2446), .D(n410), .Y(n1952) );
  OAI22X1 U1536 ( .A(n2446), .B(n360), .C(n2447), .D(n410), .Y(n1953) );
  OAI22X1 U1537 ( .A(n2447), .B(n360), .C(n2448), .D(n410), .Y(n1954) );
  OAI22X1 U1538 ( .A(n2448), .B(n360), .C(n2449), .D(n410), .Y(n1955) );
  OAI22X1 U1539 ( .A(n2449), .B(n359), .C(n2450), .D(n410), .Y(n1956) );
  OAI22X1 U1540 ( .A(n2450), .B(n359), .C(n2451), .D(n409), .Y(n1957) );
  OAI22X1 U1541 ( .A(n2451), .B(n359), .C(n2452), .D(n409), .Y(n1958) );
  OAI22X1 U1542 ( .A(n2452), .B(n359), .C(n2453), .D(n409), .Y(n1959) );
  OAI22X1 U1543 ( .A(n2453), .B(n359), .C(n2454), .D(n409), .Y(n1960) );
  OAI22X1 U1544 ( .A(n2454), .B(n359), .C(n2455), .D(n409), .Y(n1961) );
  OAI22X1 U1545 ( .A(n2455), .B(n359), .C(n2456), .D(n409), .Y(n1962) );
  OAI22X1 U1546 ( .A(n2456), .B(n359), .C(n2457), .D(n409), .Y(n1963) );
  OAI22X1 U1547 ( .A(n2457), .B(n359), .C(n2458), .D(n409), .Y(n1964) );
  OAI22X1 U1548 ( .A(n2458), .B(n359), .C(n2459), .D(n409), .Y(n1965) );
  OAI22X1 U1549 ( .A(n2459), .B(n359), .C(n2460), .D(n409), .Y(n1966) );
  XNOR2X1 U1550 ( .A(n313), .B(b[31]), .Y(n2429) );
  XNOR2X1 U1551 ( .A(n313), .B(b[30]), .Y(n2430) );
  XNOR2X1 U1552 ( .A(n313), .B(b[29]), .Y(n2431) );
  XNOR2X1 U1553 ( .A(n313), .B(b[28]), .Y(n2432) );
  XNOR2X1 U1554 ( .A(n313), .B(b[27]), .Y(n2433) );
  XNOR2X1 U1555 ( .A(n313), .B(b[26]), .Y(n2434) );
  XNOR2X1 U1556 ( .A(n313), .B(n485), .Y(n2435) );
  XNOR2X1 U1557 ( .A(n313), .B(n483), .Y(n2436) );
  XNOR2X1 U1558 ( .A(n313), .B(n481), .Y(n2437) );
  XNOR2X1 U1559 ( .A(n313), .B(n479), .Y(n2438) );
  XNOR2X1 U1560 ( .A(n313), .B(n477), .Y(n2439) );
  XNOR2X1 U1561 ( .A(n312), .B(n475), .Y(n2440) );
  XNOR2X1 U1562 ( .A(n312), .B(n473), .Y(n2441) );
  XNOR2X1 U1563 ( .A(n312), .B(n471), .Y(n2442) );
  XNOR2X1 U1564 ( .A(n312), .B(n469), .Y(n2443) );
  XNOR2X1 U1565 ( .A(n312), .B(n467), .Y(n2444) );
  XNOR2X1 U1566 ( .A(n312), .B(n2982), .Y(n2445) );
  XNOR2X1 U1567 ( .A(n312), .B(n2961), .Y(n2446) );
  XNOR2X1 U1568 ( .A(n312), .B(n2975), .Y(n2447) );
  XNOR2X1 U1569 ( .A(n312), .B(n2991), .Y(n2448) );
  XNOR2X1 U1570 ( .A(n312), .B(n2964), .Y(n2449) );
  XNOR2X1 U1571 ( .A(n312), .B(n2978), .Y(n2450) );
  XNOR2X1 U1572 ( .A(n312), .B(n2970), .Y(n2451) );
  XNOR2X1 U1573 ( .A(n311), .B(n2973), .Y(n2452) );
  XNOR2X1 U1574 ( .A(n311), .B(n2993), .Y(n2453) );
  XNOR2X1 U1575 ( .A(n311), .B(n2959), .Y(n2454) );
  XNOR2X1 U1576 ( .A(n311), .B(n2940), .Y(n2455) );
  XNOR2X1 U1577 ( .A(n311), .B(n2996), .Y(n2456) );
  XNOR2X1 U1578 ( .A(n311), .B(n2980), .Y(n2457) );
  XNOR2X1 U1579 ( .A(n311), .B(n439), .Y(n2458) );
  XNOR2X1 U1580 ( .A(n311), .B(n2911), .Y(n2459) );
  XNOR2X1 U1581 ( .A(n311), .B(n2944), .Y(n2460) );
  OAI22X1 U1582 ( .A(n358), .B(n2494), .C(n2804), .D(n408), .Y(n1751) );
  OAI22X1 U1583 ( .A(n2804), .B(n358), .C(n2462), .D(n408), .Y(n1969) );
  OAI22X1 U1584 ( .A(n2462), .B(n358), .C(n2463), .D(n408), .Y(n1970) );
  OAI22X1 U1585 ( .A(n2463), .B(n358), .C(n2464), .D(n408), .Y(n1971) );
  OAI22X1 U1586 ( .A(n2464), .B(n358), .C(n2465), .D(n408), .Y(n1972) );
  OAI22X1 U1587 ( .A(n2465), .B(n358), .C(n2466), .D(n408), .Y(n1973) );
  OAI22X1 U1588 ( .A(n2466), .B(n358), .C(n2467), .D(n408), .Y(n1974) );
  OAI22X1 U1589 ( .A(n2467), .B(n358), .C(n2468), .D(n408), .Y(n1975) );
  OAI22X1 U1590 ( .A(n2468), .B(n358), .C(n2469), .D(n408), .Y(n1976) );
  OAI22X1 U1591 ( .A(n2469), .B(n358), .C(n2470), .D(n408), .Y(n1977) );
  OAI22X1 U1592 ( .A(n2470), .B(n357), .C(n2471), .D(n408), .Y(n1978) );
  OAI22X1 U1593 ( .A(n2471), .B(n357), .C(n2472), .D(n407), .Y(n1979) );
  OAI22X1 U1594 ( .A(n2472), .B(n357), .C(n2473), .D(n407), .Y(n1980) );
  OAI22X1 U1595 ( .A(n2473), .B(n357), .C(n2474), .D(n407), .Y(n1981) );
  OAI22X1 U1596 ( .A(n2474), .B(n357), .C(n2475), .D(n407), .Y(n1982) );
  OAI22X1 U1597 ( .A(n2475), .B(n357), .C(n2476), .D(n407), .Y(n1983) );
  OAI22X1 U1598 ( .A(n2476), .B(n357), .C(n2477), .D(n407), .Y(n1984) );
  OAI22X1 U1599 ( .A(n2477), .B(n357), .C(n2478), .D(n407), .Y(n1985) );
  OAI22X1 U1600 ( .A(n2478), .B(n357), .C(n2479), .D(n407), .Y(n1986) );
  OAI22X1 U1601 ( .A(n2479), .B(n357), .C(n2480), .D(n407), .Y(n1987) );
  OAI22X1 U1602 ( .A(n2480), .B(n357), .C(n2481), .D(n407), .Y(n1988) );
  OAI22X1 U1603 ( .A(n2481), .B(n357), .C(n2482), .D(n407), .Y(n1989) );
  OAI22X1 U1604 ( .A(n2482), .B(n356), .C(n2483), .D(n407), .Y(n1990) );
  OAI22X1 U1605 ( .A(n2483), .B(n356), .C(n2484), .D(n406), .Y(n1991) );
  OAI22X1 U1606 ( .A(n2484), .B(n356), .C(n2485), .D(n406), .Y(n1992) );
  OAI22X1 U1607 ( .A(n2485), .B(n356), .C(n2486), .D(n406), .Y(n1993) );
  OAI22X1 U1608 ( .A(n2486), .B(n356), .C(n2487), .D(n406), .Y(n1994) );
  OAI22X1 U1609 ( .A(n2487), .B(n356), .C(n2488), .D(n406), .Y(n1995) );
  OAI22X1 U1610 ( .A(n2488), .B(n356), .C(n2489), .D(n406), .Y(n1996) );
  OAI22X1 U1611 ( .A(n2489), .B(n356), .C(n2490), .D(n406), .Y(n1997) );
  OAI22X1 U1612 ( .A(n2490), .B(n356), .C(n2491), .D(n406), .Y(n1998) );
  OAI22X1 U1613 ( .A(n2491), .B(n356), .C(n2492), .D(n406), .Y(n1999) );
  OAI22X1 U1614 ( .A(n2492), .B(n356), .C(n2493), .D(n406), .Y(n2000) );
  XNOR2X1 U1615 ( .A(n310), .B(n497), .Y(n2462) );
  XNOR2X1 U1616 ( .A(n310), .B(n495), .Y(n2463) );
  XNOR2X1 U1617 ( .A(n310), .B(n493), .Y(n2464) );
  XNOR2X1 U1618 ( .A(n310), .B(n491), .Y(n2465) );
  XNOR2X1 U1619 ( .A(n310), .B(n489), .Y(n2466) );
  XNOR2X1 U1620 ( .A(n310), .B(n487), .Y(n2467) );
  XNOR2X1 U1621 ( .A(n310), .B(n485), .Y(n2468) );
  XNOR2X1 U1622 ( .A(n310), .B(n483), .Y(n2469) );
  XNOR2X1 U1623 ( .A(n310), .B(n481), .Y(n2470) );
  XNOR2X1 U1624 ( .A(n310), .B(n479), .Y(n2471) );
  XNOR2X1 U1625 ( .A(n310), .B(n477), .Y(n2472) );
  XNOR2X1 U1626 ( .A(n309), .B(n475), .Y(n2473) );
  XNOR2X1 U1627 ( .A(n309), .B(n473), .Y(n2474) );
  XNOR2X1 U1628 ( .A(n309), .B(n471), .Y(n2475) );
  XNOR2X1 U1629 ( .A(n309), .B(n469), .Y(n2476) );
  XNOR2X1 U1630 ( .A(n309), .B(n467), .Y(n2477) );
  XNOR2X1 U1631 ( .A(n309), .B(n2983), .Y(n2478) );
  XNOR2X1 U1632 ( .A(n309), .B(n2962), .Y(n2479) );
  XNOR2X1 U1633 ( .A(n309), .B(n2976), .Y(n2480) );
  XNOR2X1 U1634 ( .A(n309), .B(n2991), .Y(n2481) );
  XNOR2X1 U1635 ( .A(n309), .B(n2965), .Y(n2482) );
  XNOR2X1 U1636 ( .A(n309), .B(n2978), .Y(n2483) );
  XNOR2X1 U1637 ( .A(n309), .B(n2971), .Y(n2484) );
  XNOR2X1 U1638 ( .A(n308), .B(n2973), .Y(n2485) );
  XNOR2X1 U1639 ( .A(n308), .B(n2994), .Y(n2486) );
  XNOR2X1 U1640 ( .A(n308), .B(n2960), .Y(n2487) );
  XNOR2X1 U1641 ( .A(n308), .B(n2968), .Y(n2488) );
  XNOR2X1 U1642 ( .A(n308), .B(n2996), .Y(n2489) );
  XNOR2X1 U1643 ( .A(n308), .B(n2981), .Y(n2490) );
  XNOR2X1 U1644 ( .A(n308), .B(n439), .Y(n2491) );
  XNOR2X1 U1645 ( .A(n308), .B(n2911), .Y(n2492) );
  XNOR2X1 U1646 ( .A(n308), .B(n2998), .Y(n2493) );
  OAI22X1 U1647 ( .A(n355), .B(n2527), .C(n2805), .D(n405), .Y(n1752) );
  OAI22X1 U1648 ( .A(n2805), .B(n355), .C(n2495), .D(n405), .Y(n2003) );
  OAI22X1 U1649 ( .A(n2495), .B(n355), .C(n2496), .D(n405), .Y(n2004) );
  OAI22X1 U1650 ( .A(n2496), .B(n355), .C(n2497), .D(n405), .Y(n2005) );
  OAI22X1 U1651 ( .A(n2497), .B(n355), .C(n2498), .D(n405), .Y(n2006) );
  OAI22X1 U1652 ( .A(n2498), .B(n355), .C(n2499), .D(n405), .Y(n2007) );
  OAI22X1 U1653 ( .A(n2499), .B(n355), .C(n2500), .D(n405), .Y(n2008) );
  OAI22X1 U1654 ( .A(n2500), .B(n355), .C(n2501), .D(n405), .Y(n2009) );
  OAI22X1 U1655 ( .A(n2501), .B(n355), .C(n2502), .D(n405), .Y(n2010) );
  OAI22X1 U1656 ( .A(n2502), .B(n355), .C(n2503), .D(n405), .Y(n2011) );
  OAI22X1 U1657 ( .A(n2503), .B(n354), .C(n2504), .D(n405), .Y(n2012) );
  OAI22X1 U1658 ( .A(n2504), .B(n354), .C(n2505), .D(n404), .Y(n2013) );
  OAI22X1 U1659 ( .A(n2505), .B(n354), .C(n2506), .D(n404), .Y(n2014) );
  OAI22X1 U1660 ( .A(n2506), .B(n354), .C(n2507), .D(n404), .Y(n2015) );
  OAI22X1 U1661 ( .A(n2507), .B(n354), .C(n2508), .D(n404), .Y(n2016) );
  OAI22X1 U1662 ( .A(n2508), .B(n354), .C(n2509), .D(n404), .Y(n2017) );
  OAI22X1 U1663 ( .A(n2509), .B(n354), .C(n2510), .D(n404), .Y(n2018) );
  OAI22X1 U1664 ( .A(n2510), .B(n354), .C(n2511), .D(n404), .Y(n2019) );
  OAI22X1 U1665 ( .A(n2511), .B(n354), .C(n2512), .D(n404), .Y(n2020) );
  OAI22X1 U1666 ( .A(n2512), .B(n354), .C(n2513), .D(n404), .Y(n2021) );
  OAI22X1 U1667 ( .A(n2513), .B(n354), .C(n2514), .D(n404), .Y(n2022) );
  OAI22X1 U1668 ( .A(n2514), .B(n354), .C(n2515), .D(n404), .Y(n2023) );
  OAI22X1 U1669 ( .A(n2515), .B(n353), .C(n2516), .D(n404), .Y(n2024) );
  OAI22X1 U1670 ( .A(n2516), .B(n353), .C(n2517), .D(n403), .Y(n2025) );
  OAI22X1 U1671 ( .A(n2517), .B(n353), .C(n2518), .D(n403), .Y(n2026) );
  OAI22X1 U1672 ( .A(n2518), .B(n353), .C(n2519), .D(n403), .Y(n2027) );
  OAI22X1 U1673 ( .A(n2519), .B(n353), .C(n2520), .D(n403), .Y(n2028) );
  OAI22X1 U1674 ( .A(n2520), .B(n353), .C(n2521), .D(n403), .Y(n2029) );
  OAI22X1 U1675 ( .A(n2521), .B(n353), .C(n2522), .D(n403), .Y(n2030) );
  OAI22X1 U1676 ( .A(n2522), .B(n353), .C(n2523), .D(n403), .Y(n2031) );
  OAI22X1 U1677 ( .A(n2523), .B(n353), .C(n2524), .D(n403), .Y(n2032) );
  OAI22X1 U1678 ( .A(n2524), .B(n353), .C(n2525), .D(n403), .Y(n2033) );
  OAI22X1 U1679 ( .A(n2525), .B(n353), .C(n2526), .D(n403), .Y(n2034) );
  XNOR2X1 U1680 ( .A(n307), .B(n497), .Y(n2495) );
  XNOR2X1 U1681 ( .A(n307), .B(n495), .Y(n2496) );
  XNOR2X1 U1682 ( .A(n307), .B(n493), .Y(n2497) );
  XNOR2X1 U1683 ( .A(n307), .B(n491), .Y(n2498) );
  XNOR2X1 U1684 ( .A(n307), .B(n489), .Y(n2499) );
  XNOR2X1 U1685 ( .A(n307), .B(n487), .Y(n2500) );
  XNOR2X1 U1686 ( .A(n307), .B(n485), .Y(n2501) );
  XNOR2X1 U1687 ( .A(n307), .B(n483), .Y(n2502) );
  XNOR2X1 U1688 ( .A(n307), .B(n481), .Y(n2503) );
  XNOR2X1 U1689 ( .A(n307), .B(n479), .Y(n2504) );
  XNOR2X1 U1690 ( .A(n307), .B(n477), .Y(n2505) );
  XNOR2X1 U1691 ( .A(n306), .B(n475), .Y(n2506) );
  XNOR2X1 U1692 ( .A(n306), .B(n473), .Y(n2507) );
  XNOR2X1 U1693 ( .A(n306), .B(n471), .Y(n2508) );
  XNOR2X1 U1694 ( .A(n306), .B(n469), .Y(n2509) );
  XNOR2X1 U1695 ( .A(n306), .B(n467), .Y(n2510) );
  XNOR2X1 U1696 ( .A(n306), .B(n2982), .Y(n2511) );
  XNOR2X1 U1697 ( .A(n306), .B(n2961), .Y(n2512) );
  XNOR2X1 U1698 ( .A(n306), .B(n2975), .Y(n2513) );
  XNOR2X1 U1699 ( .A(n306), .B(n2991), .Y(n2514) );
  XNOR2X1 U1700 ( .A(n306), .B(n2964), .Y(n2515) );
  XNOR2X1 U1701 ( .A(n306), .B(n2978), .Y(n2516) );
  XNOR2X1 U1702 ( .A(n306), .B(n2970), .Y(n2517) );
  XNOR2X1 U1703 ( .A(n305), .B(n2973), .Y(n2518) );
  XNOR2X1 U1704 ( .A(n305), .B(n2993), .Y(n2519) );
  XNOR2X1 U1705 ( .A(n305), .B(n2959), .Y(n2520) );
  XNOR2X1 U1706 ( .A(n305), .B(n2968), .Y(n2521) );
  XNOR2X1 U1707 ( .A(n305), .B(n2996), .Y(n2522) );
  XNOR2X1 U1708 ( .A(n305), .B(n2980), .Y(n2523) );
  XNOR2X1 U1709 ( .A(n305), .B(n2915), .Y(n2524) );
  XNOR2X1 U1710 ( .A(n305), .B(n2911), .Y(n2525) );
  XNOR2X1 U1711 ( .A(n305), .B(n2998), .Y(n2526) );
  OAI22X1 U1712 ( .A(n352), .B(n2560), .C(n2806), .D(n402), .Y(n1753) );
  OAI22X1 U1713 ( .A(n2806), .B(n352), .C(n2528), .D(n402), .Y(n2037) );
  OAI22X1 U1714 ( .A(n2528), .B(n352), .C(n2529), .D(n402), .Y(n2038) );
  OAI22X1 U1715 ( .A(n2529), .B(n352), .C(n2530), .D(n402), .Y(n2039) );
  OAI22X1 U1716 ( .A(n2530), .B(n352), .C(n2531), .D(n402), .Y(n2040) );
  OAI22X1 U1717 ( .A(n2531), .B(n352), .C(n2532), .D(n402), .Y(n2041) );
  OAI22X1 U1718 ( .A(n2532), .B(n352), .C(n2533), .D(n402), .Y(n2042) );
  OAI22X1 U1719 ( .A(n2533), .B(n352), .C(n2534), .D(n402), .Y(n2043) );
  OAI22X1 U1720 ( .A(n2534), .B(n352), .C(n2535), .D(n402), .Y(n2044) );
  OAI22X1 U1721 ( .A(n2535), .B(n352), .C(n2536), .D(n402), .Y(n2045) );
  OAI22X1 U1722 ( .A(n2536), .B(n351), .C(n2537), .D(n402), .Y(n2046) );
  OAI22X1 U1723 ( .A(n2537), .B(n351), .C(n2538), .D(n401), .Y(n2047) );
  OAI22X1 U1724 ( .A(n2538), .B(n351), .C(n2539), .D(n401), .Y(n2048) );
  OAI22X1 U1725 ( .A(n2539), .B(n351), .C(n2540), .D(n401), .Y(n2049) );
  OAI22X1 U1726 ( .A(n2540), .B(n351), .C(n2541), .D(n401), .Y(n2050) );
  OAI22X1 U1727 ( .A(n2541), .B(n351), .C(n2542), .D(n401), .Y(n2051) );
  OAI22X1 U1728 ( .A(n2542), .B(n351), .C(n2543), .D(n401), .Y(n2052) );
  OAI22X1 U1729 ( .A(n2543), .B(n351), .C(n2544), .D(n401), .Y(n2053) );
  OAI22X1 U1730 ( .A(n2544), .B(n351), .C(n2545), .D(n401), .Y(n2054) );
  OAI22X1 U1731 ( .A(n2545), .B(n351), .C(n2546), .D(n401), .Y(n2055) );
  OAI22X1 U1732 ( .A(n2546), .B(n351), .C(n2547), .D(n401), .Y(n2056) );
  OAI22X1 U1733 ( .A(n2547), .B(n351), .C(n2548), .D(n401), .Y(n2057) );
  OAI22X1 U1734 ( .A(n2548), .B(n350), .C(n2549), .D(n401), .Y(n2058) );
  OAI22X1 U1735 ( .A(n2549), .B(n350), .C(n2550), .D(n400), .Y(n2059) );
  OAI22X1 U1736 ( .A(n2550), .B(n350), .C(n2551), .D(n400), .Y(n2060) );
  OAI22X1 U1737 ( .A(n2551), .B(n350), .C(n2552), .D(n400), .Y(n2061) );
  OAI22X1 U1738 ( .A(n2552), .B(n350), .C(n2553), .D(n400), .Y(n2062) );
  OAI22X1 U1739 ( .A(n2553), .B(n350), .C(n2554), .D(n400), .Y(n2063) );
  OAI22X1 U1740 ( .A(n2554), .B(n350), .C(n2555), .D(n400), .Y(n2064) );
  OAI22X1 U1741 ( .A(n2555), .B(n350), .C(n2556), .D(n400), .Y(n2065) );
  OAI22X1 U1742 ( .A(n2556), .B(n350), .C(n2557), .D(n400), .Y(n2066) );
  OAI22X1 U1743 ( .A(n2557), .B(n350), .C(n2558), .D(n400), .Y(n2067) );
  OAI22X1 U1744 ( .A(n2558), .B(n350), .C(n2559), .D(n400), .Y(n2068) );
  XNOR2X1 U1745 ( .A(n304), .B(n497), .Y(n2528) );
  XNOR2X1 U1746 ( .A(n304), .B(n495), .Y(n2529) );
  XNOR2X1 U1747 ( .A(n304), .B(n493), .Y(n2530) );
  XNOR2X1 U1748 ( .A(n304), .B(n491), .Y(n2531) );
  XNOR2X1 U1749 ( .A(n304), .B(n489), .Y(n2532) );
  XNOR2X1 U1750 ( .A(n304), .B(n487), .Y(n2533) );
  XNOR2X1 U1751 ( .A(n304), .B(n485), .Y(n2534) );
  XNOR2X1 U1752 ( .A(n304), .B(n483), .Y(n2535) );
  XNOR2X1 U1753 ( .A(n304), .B(n481), .Y(n2536) );
  XNOR2X1 U1754 ( .A(n304), .B(n479), .Y(n2537) );
  XNOR2X1 U1755 ( .A(n304), .B(n477), .Y(n2538) );
  XNOR2X1 U1756 ( .A(n303), .B(n475), .Y(n2539) );
  XNOR2X1 U1757 ( .A(n303), .B(n473), .Y(n2540) );
  XNOR2X1 U1758 ( .A(n303), .B(n471), .Y(n2541) );
  XNOR2X1 U1759 ( .A(n303), .B(n469), .Y(n2542) );
  XNOR2X1 U1760 ( .A(n303), .B(n467), .Y(n2543) );
  XNOR2X1 U1761 ( .A(n303), .B(n2983), .Y(n2544) );
  XNOR2X1 U1762 ( .A(n303), .B(n2962), .Y(n2545) );
  XNOR2X1 U1763 ( .A(n303), .B(n2976), .Y(n2546) );
  XNOR2X1 U1764 ( .A(n303), .B(n2991), .Y(n2547) );
  XNOR2X1 U1765 ( .A(n303), .B(n2965), .Y(n2548) );
  XNOR2X1 U1766 ( .A(n303), .B(n2978), .Y(n2549) );
  XNOR2X1 U1767 ( .A(n303), .B(n2971), .Y(n2550) );
  XNOR2X1 U1768 ( .A(n302), .B(n2973), .Y(n2551) );
  XNOR2X1 U1769 ( .A(n302), .B(n2994), .Y(n2552) );
  XNOR2X1 U1770 ( .A(n302), .B(n2960), .Y(n2553) );
  XNOR2X1 U1771 ( .A(n302), .B(n2940), .Y(n2554) );
  XNOR2X1 U1772 ( .A(n302), .B(n2996), .Y(n2555) );
  XNOR2X1 U1773 ( .A(n302), .B(n2979), .Y(n2556) );
  XNOR2X1 U1774 ( .A(n302), .B(n2915), .Y(n2557) );
  XNOR2X1 U1775 ( .A(n302), .B(n2985), .Y(n2558) );
  XNOR2X1 U1776 ( .A(n302), .B(n2997), .Y(n2559) );
  OAI22X1 U1777 ( .A(n349), .B(n2593), .C(n2807), .D(n399), .Y(n1754) );
  OAI22X1 U1778 ( .A(n2807), .B(n349), .C(n2561), .D(n399), .Y(n2071) );
  OAI22X1 U1779 ( .A(n2561), .B(n349), .C(n2562), .D(n399), .Y(n2072) );
  OAI22X1 U1780 ( .A(n2562), .B(n349), .C(n2563), .D(n399), .Y(n2073) );
  OAI22X1 U1781 ( .A(n2563), .B(n349), .C(n2564), .D(n399), .Y(n2074) );
  OAI22X1 U1782 ( .A(n2564), .B(n349), .C(n2565), .D(n399), .Y(n2075) );
  OAI22X1 U1783 ( .A(n2565), .B(n349), .C(n2566), .D(n399), .Y(n2076) );
  OAI22X1 U1784 ( .A(n2566), .B(n349), .C(n2567), .D(n399), .Y(n2077) );
  OAI22X1 U1785 ( .A(n2567), .B(n349), .C(n2568), .D(n399), .Y(n2078) );
  OAI22X1 U1786 ( .A(n2568), .B(n349), .C(n2569), .D(n399), .Y(n2079) );
  OAI22X1 U1787 ( .A(n2569), .B(n348), .C(n2570), .D(n399), .Y(n2080) );
  OAI22X1 U1788 ( .A(n2570), .B(n348), .C(n2571), .D(n398), .Y(n2081) );
  OAI22X1 U1789 ( .A(n2571), .B(n348), .C(n2572), .D(n398), .Y(n2082) );
  OAI22X1 U1790 ( .A(n2572), .B(n348), .C(n2573), .D(n398), .Y(n2083) );
  OAI22X1 U1791 ( .A(n2573), .B(n348), .C(n2574), .D(n398), .Y(n2084) );
  OAI22X1 U1792 ( .A(n2574), .B(n348), .C(n2575), .D(n398), .Y(n2085) );
  OAI22X1 U1793 ( .A(n2575), .B(n348), .C(n2576), .D(n398), .Y(n2086) );
  OAI22X1 U1794 ( .A(n2576), .B(n348), .C(n2577), .D(n398), .Y(n2087) );
  OAI22X1 U1795 ( .A(n2577), .B(n348), .C(n2578), .D(n398), .Y(n2088) );
  OAI22X1 U1796 ( .A(n2578), .B(n348), .C(n2579), .D(n398), .Y(n2089) );
  OAI22X1 U1797 ( .A(n2579), .B(n348), .C(n2580), .D(n398), .Y(n2090) );
  OAI22X1 U1798 ( .A(n2580), .B(n348), .C(n2581), .D(n398), .Y(n2091) );
  OAI22X1 U1799 ( .A(n2581), .B(n347), .C(n2582), .D(n398), .Y(n2092) );
  OAI22X1 U1800 ( .A(n2582), .B(n347), .C(n2583), .D(n397), .Y(n2093) );
  OAI22X1 U1801 ( .A(n2583), .B(n347), .C(n2584), .D(n397), .Y(n2094) );
  OAI22X1 U1802 ( .A(n2584), .B(n347), .C(n2585), .D(n397), .Y(n2095) );
  OAI22X1 U1803 ( .A(n2585), .B(n347), .C(n2586), .D(n397), .Y(n2096) );
  OAI22X1 U1804 ( .A(n2586), .B(n347), .C(n2587), .D(n397), .Y(n2097) );
  OAI22X1 U1805 ( .A(n2587), .B(n347), .C(n2588), .D(n397), .Y(n2098) );
  OAI22X1 U1806 ( .A(n2588), .B(n347), .C(n2589), .D(n397), .Y(n2099) );
  OAI22X1 U1807 ( .A(n2589), .B(n347), .C(n2590), .D(n397), .Y(n2100) );
  OAI22X1 U1808 ( .A(n2590), .B(n347), .C(n2591), .D(n397), .Y(n2101) );
  OAI22X1 U1809 ( .A(n2591), .B(n347), .C(n2592), .D(n397), .Y(n2102) );
  XNOR2X1 U1810 ( .A(n301), .B(n497), .Y(n2561) );
  XNOR2X1 U1811 ( .A(n301), .B(n495), .Y(n2562) );
  XNOR2X1 U1812 ( .A(n301), .B(n493), .Y(n2563) );
  XNOR2X1 U1813 ( .A(n301), .B(n491), .Y(n2564) );
  XNOR2X1 U1814 ( .A(n301), .B(n489), .Y(n2565) );
  XNOR2X1 U1815 ( .A(n301), .B(n487), .Y(n2566) );
  XNOR2X1 U1816 ( .A(n301), .B(n485), .Y(n2567) );
  XNOR2X1 U1817 ( .A(n301), .B(n483), .Y(n2568) );
  XNOR2X1 U1818 ( .A(n301), .B(n481), .Y(n2569) );
  XNOR2X1 U1819 ( .A(n301), .B(n479), .Y(n2570) );
  XNOR2X1 U1820 ( .A(n301), .B(n477), .Y(n2571) );
  XNOR2X1 U1821 ( .A(n300), .B(n475), .Y(n2572) );
  XNOR2X1 U1822 ( .A(n300), .B(n473), .Y(n2573) );
  XNOR2X1 U1823 ( .A(n300), .B(n471), .Y(n2574) );
  XNOR2X1 U1824 ( .A(n300), .B(n469), .Y(n2575) );
  XNOR2X1 U1825 ( .A(n300), .B(n467), .Y(n2576) );
  XNOR2X1 U1826 ( .A(n300), .B(n2982), .Y(n2577) );
  XNOR2X1 U1827 ( .A(n300), .B(n2961), .Y(n2578) );
  XNOR2X1 U1828 ( .A(n300), .B(n2975), .Y(n2579) );
  XNOR2X1 U1829 ( .A(n300), .B(n459), .Y(n2580) );
  XNOR2X1 U1830 ( .A(n300), .B(n2964), .Y(n2581) );
  XNOR2X1 U1831 ( .A(n300), .B(n2978), .Y(n2582) );
  XNOR2X1 U1832 ( .A(n300), .B(n2970), .Y(n2583) );
  XNOR2X1 U1833 ( .A(n299), .B(n2973), .Y(n2584) );
  XNOR2X1 U1834 ( .A(n299), .B(n2993), .Y(n2585) );
  XNOR2X1 U1835 ( .A(n299), .B(n2959), .Y(n2586) );
  XNOR2X1 U1836 ( .A(n299), .B(n2968), .Y(n2587) );
  XNOR2X1 U1837 ( .A(n299), .B(b[4]), .Y(n2588) );
  XNOR2X1 U1838 ( .A(n299), .B(n2979), .Y(n2589) );
  XNOR2X1 U1839 ( .A(n299), .B(n2915), .Y(n2590) );
  XNOR2X1 U1840 ( .A(n299), .B(n2910), .Y(n2591) );
  XNOR2X1 U1841 ( .A(n299), .B(n2941), .Y(n2592) );
  OAI22X1 U1842 ( .A(n346), .B(n2626), .C(n2808), .D(n396), .Y(n1755) );
  OAI22X1 U1843 ( .A(n2808), .B(n346), .C(n2594), .D(n396), .Y(n2105) );
  OAI22X1 U1844 ( .A(n2594), .B(n346), .C(n2595), .D(n396), .Y(n2106) );
  OAI22X1 U1845 ( .A(n2595), .B(n346), .C(n2596), .D(n396), .Y(n2107) );
  OAI22X1 U1846 ( .A(n2596), .B(n346), .C(n2597), .D(n396), .Y(n2108) );
  OAI22X1 U1847 ( .A(n2597), .B(n346), .C(n2598), .D(n396), .Y(n2109) );
  OAI22X1 U1848 ( .A(n2598), .B(n346), .C(n2599), .D(n396), .Y(n2110) );
  OAI22X1 U1849 ( .A(n2599), .B(n346), .C(n2600), .D(n396), .Y(n2111) );
  OAI22X1 U1850 ( .A(n2600), .B(n346), .C(n2601), .D(n396), .Y(n2112) );
  OAI22X1 U1851 ( .A(n2601), .B(n346), .C(n2602), .D(n396), .Y(n2113) );
  OAI22X1 U1852 ( .A(n2602), .B(n345), .C(n2603), .D(n396), .Y(n2114) );
  OAI22X1 U1853 ( .A(n2603), .B(n345), .C(n2604), .D(n395), .Y(n2115) );
  OAI22X1 U1854 ( .A(n2604), .B(n345), .C(n2605), .D(n395), .Y(n2116) );
  OAI22X1 U1855 ( .A(n2605), .B(n345), .C(n2606), .D(n395), .Y(n2117) );
  OAI22X1 U1856 ( .A(n2606), .B(n345), .C(n2607), .D(n395), .Y(n2118) );
  OAI22X1 U1857 ( .A(n2607), .B(n345), .C(n2608), .D(n395), .Y(n2119) );
  OAI22X1 U1858 ( .A(n2608), .B(n345), .C(n2609), .D(n395), .Y(n2120) );
  OAI22X1 U1859 ( .A(n2609), .B(n345), .C(n2610), .D(n395), .Y(n2121) );
  OAI22X1 U1860 ( .A(n2610), .B(n345), .C(n2611), .D(n395), .Y(n2122) );
  OAI22X1 U1861 ( .A(n2611), .B(n345), .C(n2612), .D(n395), .Y(n2123) );
  OAI22X1 U1862 ( .A(n2612), .B(n345), .C(n2613), .D(n395), .Y(n2124) );
  OAI22X1 U1863 ( .A(n2613), .B(n345), .C(n2614), .D(n395), .Y(n2125) );
  OAI22X1 U1864 ( .A(n2614), .B(n344), .C(n2615), .D(n395), .Y(n2126) );
  OAI22X1 U1865 ( .A(n2615), .B(n344), .C(n2616), .D(n394), .Y(n2127) );
  OAI22X1 U1866 ( .A(n2616), .B(n344), .C(n2617), .D(n394), .Y(n2128) );
  OAI22X1 U1867 ( .A(n2617), .B(n344), .C(n2618), .D(n394), .Y(n2129) );
  OAI22X1 U1868 ( .A(n2618), .B(n344), .C(n2619), .D(n394), .Y(n2130) );
  OAI22X1 U1869 ( .A(n2619), .B(n344), .C(n2620), .D(n394), .Y(n2131) );
  OAI22X1 U1870 ( .A(n2620), .B(n344), .C(n2621), .D(n394), .Y(n2132) );
  OAI22X1 U1871 ( .A(n2621), .B(n344), .C(n2622), .D(n394), .Y(n2133) );
  OAI22X1 U1872 ( .A(n2622), .B(n344), .C(n2623), .D(n394), .Y(n2134) );
  OAI22X1 U1873 ( .A(n2623), .B(n344), .C(n2624), .D(n394), .Y(n2135) );
  OAI22X1 U1874 ( .A(n2624), .B(n344), .C(n2625), .D(n394), .Y(n2136) );
  XNOR2X1 U1875 ( .A(n298), .B(n497), .Y(n2594) );
  XNOR2X1 U1876 ( .A(n298), .B(n495), .Y(n2595) );
  XNOR2X1 U1877 ( .A(n298), .B(n493), .Y(n2596) );
  XNOR2X1 U1878 ( .A(n298), .B(n491), .Y(n2597) );
  XNOR2X1 U1879 ( .A(n298), .B(n489), .Y(n2598) );
  XNOR2X1 U1880 ( .A(n298), .B(n487), .Y(n2599) );
  XNOR2X1 U1881 ( .A(n298), .B(n485), .Y(n2600) );
  XNOR2X1 U1882 ( .A(n298), .B(n483), .Y(n2601) );
  XNOR2X1 U1883 ( .A(n298), .B(n481), .Y(n2602) );
  XNOR2X1 U1884 ( .A(n298), .B(n479), .Y(n2603) );
  XNOR2X1 U1885 ( .A(n298), .B(n477), .Y(n2604) );
  XNOR2X1 U1886 ( .A(n297), .B(n475), .Y(n2605) );
  XNOR2X1 U1887 ( .A(n297), .B(n473), .Y(n2606) );
  XNOR2X1 U1888 ( .A(n297), .B(n471), .Y(n2607) );
  XNOR2X1 U1889 ( .A(n297), .B(n469), .Y(n2608) );
  XNOR2X1 U1890 ( .A(n297), .B(n467), .Y(n2609) );
  XNOR2X1 U1891 ( .A(n297), .B(n2983), .Y(n2610) );
  XNOR2X1 U1892 ( .A(n297), .B(n2962), .Y(n2611) );
  XNOR2X1 U1893 ( .A(n297), .B(n2976), .Y(n2612) );
  XNOR2X1 U1894 ( .A(n297), .B(n459), .Y(n2613) );
  XNOR2X1 U1895 ( .A(n297), .B(n2965), .Y(n2614) );
  XNOR2X1 U1896 ( .A(n297), .B(n2978), .Y(n2615) );
  XNOR2X1 U1897 ( .A(n297), .B(n2971), .Y(n2616) );
  XNOR2X1 U1898 ( .A(n296), .B(b[8]), .Y(n2617) );
  XNOR2X1 U1899 ( .A(n296), .B(b[7]), .Y(n2618) );
  XNOR2X1 U1900 ( .A(n296), .B(n2959), .Y(n2619) );
  XNOR2X1 U1901 ( .A(n296), .B(n2967), .Y(n2620) );
  XNOR2X1 U1902 ( .A(n296), .B(b[4]), .Y(n2621) );
  XNOR2X1 U1903 ( .A(n296), .B(n2995), .Y(n2622) );
  XNOR2X1 U1904 ( .A(n296), .B(n2915), .Y(n2623) );
  XNOR2X1 U1905 ( .A(n296), .B(n2985), .Y(n2624) );
  XNOR2X1 U1906 ( .A(n296), .B(n2997), .Y(n2625) );
  OAI22X1 U1907 ( .A(n343), .B(n2659), .C(n2809), .D(n393), .Y(n1756) );
  OAI22X1 U1908 ( .A(n2809), .B(n343), .C(n2627), .D(n393), .Y(n2139) );
  OAI22X1 U1909 ( .A(n2627), .B(n343), .C(n2628), .D(n393), .Y(n2140) );
  OAI22X1 U1910 ( .A(n2628), .B(n343), .C(n2629), .D(n393), .Y(n2141) );
  OAI22X1 U1911 ( .A(n2629), .B(n343), .C(n2630), .D(n393), .Y(n2142) );
  OAI22X1 U1912 ( .A(n2630), .B(n343), .C(n2631), .D(n393), .Y(n2143) );
  OAI22X1 U1913 ( .A(n2631), .B(n343), .C(n2632), .D(n393), .Y(n2144) );
  OAI22X1 U1914 ( .A(n2632), .B(n343), .C(n2633), .D(n393), .Y(n2145) );
  OAI22X1 U1915 ( .A(n2633), .B(n343), .C(n2634), .D(n393), .Y(n2146) );
  OAI22X1 U1916 ( .A(n2634), .B(n343), .C(n2635), .D(n393), .Y(n2147) );
  OAI22X1 U1917 ( .A(n2635), .B(n342), .C(n2636), .D(n393), .Y(n2148) );
  OAI22X1 U1918 ( .A(n2636), .B(n342), .C(n2637), .D(n392), .Y(n2149) );
  OAI22X1 U1919 ( .A(n2637), .B(n342), .C(n2638), .D(n392), .Y(n2150) );
  OAI22X1 U1920 ( .A(n2638), .B(n342), .C(n2639), .D(n392), .Y(n2151) );
  OAI22X1 U1921 ( .A(n2639), .B(n342), .C(n2640), .D(n392), .Y(n2152) );
  OAI22X1 U1922 ( .A(n2640), .B(n342), .C(n2641), .D(n392), .Y(n2153) );
  OAI22X1 U1923 ( .A(n2641), .B(n342), .C(n2642), .D(n392), .Y(n2154) );
  OAI22X1 U1924 ( .A(n2642), .B(n342), .C(n2643), .D(n392), .Y(n2155) );
  OAI22X1 U1925 ( .A(n2643), .B(n342), .C(n2644), .D(n392), .Y(n2156) );
  OAI22X1 U1926 ( .A(n2644), .B(n342), .C(n2645), .D(n392), .Y(n2157) );
  OAI22X1 U1927 ( .A(n2645), .B(n342), .C(n2646), .D(n392), .Y(n2158) );
  OAI22X1 U1928 ( .A(n2646), .B(n342), .C(n2647), .D(n392), .Y(n2159) );
  OAI22X1 U1929 ( .A(n2647), .B(n341), .C(n2648), .D(n392), .Y(n2160) );
  OAI22X1 U1930 ( .A(n2648), .B(n341), .C(n2649), .D(n391), .Y(n2161) );
  OAI22X1 U1931 ( .A(n2649), .B(n341), .C(n2650), .D(n391), .Y(n2162) );
  OAI22X1 U1932 ( .A(n2650), .B(n341), .C(n2651), .D(n391), .Y(n2163) );
  OAI22X1 U1933 ( .A(n2651), .B(n341), .C(n2652), .D(n391), .Y(n2164) );
  OAI22X1 U1934 ( .A(n2652), .B(n341), .C(n2653), .D(n391), .Y(n2165) );
  OAI22X1 U1935 ( .A(n2653), .B(n341), .C(n2654), .D(n391), .Y(n2166) );
  OAI22X1 U1936 ( .A(n2654), .B(n341), .C(n2655), .D(n391), .Y(n2167) );
  OAI22X1 U1937 ( .A(n2655), .B(n341), .C(n2656), .D(n391), .Y(n2168) );
  OAI22X1 U1938 ( .A(n2656), .B(n341), .C(n2657), .D(n391), .Y(n2169) );
  OAI22X1 U1939 ( .A(n2657), .B(n341), .C(n2658), .D(n391), .Y(n2170) );
  XNOR2X1 U1940 ( .A(n295), .B(n497), .Y(n2627) );
  XNOR2X1 U1941 ( .A(n295), .B(n495), .Y(n2628) );
  XNOR2X1 U1942 ( .A(n295), .B(n493), .Y(n2629) );
  XNOR2X1 U1943 ( .A(n295), .B(n491), .Y(n2630) );
  XNOR2X1 U1944 ( .A(n295), .B(n489), .Y(n2631) );
  XNOR2X1 U1945 ( .A(n295), .B(n487), .Y(n2632) );
  XNOR2X1 U1946 ( .A(n295), .B(n485), .Y(n2633) );
  XNOR2X1 U1947 ( .A(n295), .B(n483), .Y(n2634) );
  XNOR2X1 U1948 ( .A(n295), .B(n481), .Y(n2635) );
  XNOR2X1 U1949 ( .A(n295), .B(n479), .Y(n2636) );
  XNOR2X1 U1950 ( .A(n295), .B(n477), .Y(n2637) );
  XNOR2X1 U1951 ( .A(n294), .B(n475), .Y(n2638) );
  XNOR2X1 U1952 ( .A(n294), .B(n473), .Y(n2639) );
  XNOR2X1 U1953 ( .A(n294), .B(n471), .Y(n2640) );
  XNOR2X1 U1954 ( .A(n294), .B(n469), .Y(n2641) );
  XNOR2X1 U1955 ( .A(n294), .B(n467), .Y(n2642) );
  XNOR2X1 U1956 ( .A(n294), .B(n2982), .Y(n2643) );
  XNOR2X1 U1957 ( .A(n294), .B(n2961), .Y(n2644) );
  XNOR2X1 U1958 ( .A(n294), .B(n2975), .Y(n2645) );
  XNOR2X1 U1959 ( .A(n294), .B(n459), .Y(n2646) );
  XNOR2X1 U1960 ( .A(n294), .B(n2964), .Y(n2647) );
  XNOR2X1 U1961 ( .A(n294), .B(n2978), .Y(n2648) );
  XNOR2X1 U1962 ( .A(n294), .B(n2970), .Y(n2649) );
  XNOR2X1 U1963 ( .A(n293), .B(b[8]), .Y(n2650) );
  XNOR2X1 U1964 ( .A(n293), .B(b[7]), .Y(n2651) );
  XNOR2X1 U1965 ( .A(n293), .B(n2960), .Y(n2652) );
  XNOR2X1 U1966 ( .A(n293), .B(n2968), .Y(n2653) );
  XNOR2X1 U1967 ( .A(n293), .B(b[4]), .Y(n2654) );
  XNOR2X1 U1968 ( .A(n293), .B(n441), .Y(n2655) );
  XNOR2X1 U1969 ( .A(n2914), .B(n293), .Y(n2656) );
  XNOR2X1 U1970 ( .A(n293), .B(n2910), .Y(n2657) );
  XNOR2X1 U1971 ( .A(n293), .B(n2944), .Y(n2658) );
  OAI22X1 U1972 ( .A(n340), .B(n2692), .C(n2810), .D(n390), .Y(n1757) );
  OAI22X1 U1973 ( .A(n2810), .B(n340), .C(n2660), .D(n390), .Y(n2173) );
  OAI22X1 U1974 ( .A(n2660), .B(n340), .C(n2661), .D(n390), .Y(n2174) );
  OAI22X1 U1975 ( .A(n2661), .B(n340), .C(n2662), .D(n390), .Y(n2175) );
  OAI22X1 U1976 ( .A(n2662), .B(n340), .C(n2663), .D(n390), .Y(n2176) );
  OAI22X1 U1977 ( .A(n2663), .B(n340), .C(n2664), .D(n390), .Y(n2177) );
  OAI22X1 U1978 ( .A(n2664), .B(n340), .C(n2665), .D(n390), .Y(n2178) );
  OAI22X1 U1979 ( .A(n2665), .B(n340), .C(n2666), .D(n390), .Y(n2179) );
  OAI22X1 U1980 ( .A(n2666), .B(n340), .C(n2667), .D(n390), .Y(n2180) );
  OAI22X1 U1981 ( .A(n2667), .B(n340), .C(n2668), .D(n390), .Y(n2181) );
  OAI22X1 U1982 ( .A(n2668), .B(n339), .C(n2669), .D(n390), .Y(n2182) );
  OAI22X1 U1983 ( .A(n2669), .B(n339), .C(n2670), .D(n389), .Y(n2183) );
  OAI22X1 U1984 ( .A(n2670), .B(n339), .C(n2671), .D(n389), .Y(n2184) );
  OAI22X1 U1985 ( .A(n2671), .B(n339), .C(n2672), .D(n389), .Y(n2185) );
  OAI22X1 U1986 ( .A(n2672), .B(n339), .C(n2673), .D(n389), .Y(n2186) );
  OAI22X1 U1987 ( .A(n2673), .B(n339), .C(n2674), .D(n389), .Y(n2187) );
  OAI22X1 U1988 ( .A(n2674), .B(n339), .C(n2675), .D(n389), .Y(n2188) );
  OAI22X1 U1989 ( .A(n2675), .B(n339), .C(n2676), .D(n389), .Y(n2189) );
  OAI22X1 U1990 ( .A(n2676), .B(n339), .C(n2677), .D(n389), .Y(n2190) );
  OAI22X1 U1991 ( .A(n2677), .B(n339), .C(n2678), .D(n389), .Y(n2191) );
  OAI22X1 U1992 ( .A(n2678), .B(n339), .C(n2679), .D(n389), .Y(n2192) );
  OAI22X1 U1993 ( .A(n2679), .B(n339), .C(n2680), .D(n389), .Y(n2193) );
  OAI22X1 U1994 ( .A(n2680), .B(n338), .C(n2681), .D(n389), .Y(n2194) );
  OAI22X1 U1995 ( .A(n2681), .B(n338), .C(n2682), .D(n388), .Y(n2195) );
  OAI22X1 U1996 ( .A(n2682), .B(n338), .C(n2683), .D(n388), .Y(n2196) );
  OAI22X1 U1997 ( .A(n2683), .B(n338), .C(n2684), .D(n388), .Y(n2197) );
  OAI22X1 U1998 ( .A(n2684), .B(n338), .C(n2685), .D(n388), .Y(n2198) );
  OAI22X1 U1999 ( .A(n2685), .B(n338), .C(n2686), .D(n388), .Y(n2199) );
  OAI22X1 U2000 ( .A(n2686), .B(n338), .C(n2687), .D(n388), .Y(n2200) );
  OAI22X1 U2001 ( .A(n2687), .B(n338), .C(n2688), .D(n388), .Y(n2201) );
  OAI22X1 U2002 ( .A(n2688), .B(n338), .C(n2689), .D(n388), .Y(n2202) );
  OAI22X1 U2003 ( .A(n2689), .B(n338), .C(n2690), .D(n388), .Y(n2203) );
  OAI22X1 U2004 ( .A(n2690), .B(n338), .C(n2691), .D(n388), .Y(n2204) );
  XNOR2X1 U2005 ( .A(n292), .B(n497), .Y(n2660) );
  XNOR2X1 U2006 ( .A(n292), .B(n495), .Y(n2661) );
  XNOR2X1 U2007 ( .A(n292), .B(n493), .Y(n2662) );
  XNOR2X1 U2008 ( .A(n292), .B(n491), .Y(n2663) );
  XNOR2X1 U2009 ( .A(n292), .B(n489), .Y(n2664) );
  XNOR2X1 U2010 ( .A(n292), .B(n487), .Y(n2665) );
  XNOR2X1 U2011 ( .A(n292), .B(n485), .Y(n2666) );
  XNOR2X1 U2012 ( .A(n292), .B(n483), .Y(n2667) );
  XNOR2X1 U2013 ( .A(n292), .B(n481), .Y(n2668) );
  XNOR2X1 U2014 ( .A(n292), .B(n479), .Y(n2669) );
  XNOR2X1 U2015 ( .A(n292), .B(n477), .Y(n2670) );
  XNOR2X1 U2016 ( .A(n291), .B(n475), .Y(n2671) );
  XNOR2X1 U2017 ( .A(n291), .B(n473), .Y(n2672) );
  XNOR2X1 U2018 ( .A(n291), .B(n471), .Y(n2673) );
  XNOR2X1 U2019 ( .A(n291), .B(n469), .Y(n2674) );
  XNOR2X1 U2020 ( .A(n291), .B(n467), .Y(n2675) );
  XNOR2X1 U2021 ( .A(n291), .B(n2983), .Y(n2676) );
  XNOR2X1 U2022 ( .A(n291), .B(n2962), .Y(n2677) );
  XNOR2X1 U2023 ( .A(n291), .B(n2976), .Y(n2678) );
  XNOR2X1 U2024 ( .A(n291), .B(n459), .Y(n2679) );
  XNOR2X1 U2025 ( .A(n291), .B(b[11]), .Y(n2680) );
  XNOR2X1 U2026 ( .A(n291), .B(b[10]), .Y(n2681) );
  XNOR2X1 U2027 ( .A(n291), .B(n2969), .Y(n2682) );
  XNOR2X1 U2028 ( .A(n290), .B(b[8]), .Y(n2683) );
  XNOR2X1 U2029 ( .A(n290), .B(b[7]), .Y(n2684) );
  XNOR2X1 U2030 ( .A(n290), .B(n2958), .Y(n2685) );
  XNOR2X1 U2031 ( .A(n290), .B(n2967), .Y(n2686) );
  XNOR2X1 U2032 ( .A(n290), .B(b[4]), .Y(n2687) );
  XNOR2X1 U2033 ( .A(n290), .B(n2943), .Y(n2688) );
  XNOR2X1 U2034 ( .A(n290), .B(n2915), .Y(n2689) );
  XNOR2X1 U2035 ( .A(n290), .B(n2910), .Y(n2690) );
  XNOR2X1 U2036 ( .A(n290), .B(n2912), .Y(n2691) );
  OAI22X1 U2037 ( .A(n337), .B(n2725), .C(n2811), .D(n387), .Y(n1758) );
  OAI22X1 U2038 ( .A(n337), .B(n2811), .C(n2693), .D(n387), .Y(n2207) );
  OAI22X1 U2039 ( .A(n337), .B(n2693), .C(n2694), .D(n387), .Y(n2208) );
  OAI22X1 U2040 ( .A(n337), .B(n2694), .C(n2695), .D(n387), .Y(n2209) );
  OAI22X1 U2041 ( .A(n337), .B(n2695), .C(n2696), .D(n387), .Y(n2210) );
  OAI22X1 U2042 ( .A(n337), .B(n2696), .C(n2697), .D(n387), .Y(n2211) );
  OAI22X1 U2043 ( .A(n337), .B(n2697), .C(n2698), .D(n387), .Y(n2212) );
  OAI22X1 U2044 ( .A(n337), .B(n2698), .C(n2699), .D(n387), .Y(n2213) );
  OAI22X1 U2045 ( .A(n337), .B(n2699), .C(n2700), .D(n387), .Y(n2214) );
  OAI22X1 U2046 ( .A(n337), .B(n2700), .C(n2701), .D(n387), .Y(n2215) );
  OAI22X1 U2047 ( .A(n336), .B(n2701), .C(n2702), .D(n387), .Y(n2216) );
  OAI22X1 U2048 ( .A(n336), .B(n2702), .C(n2703), .D(n386), .Y(n2217) );
  OAI22X1 U2049 ( .A(n336), .B(n2703), .C(n2704), .D(n386), .Y(n2218) );
  OAI22X1 U2050 ( .A(n336), .B(n2704), .C(n2705), .D(n386), .Y(n2219) );
  OAI22X1 U2051 ( .A(n336), .B(n2705), .C(n2706), .D(n386), .Y(n2220) );
  OAI22X1 U2052 ( .A(n336), .B(n2706), .C(n2707), .D(n386), .Y(n2221) );
  OAI22X1 U2053 ( .A(n336), .B(n2707), .C(n2708), .D(n386), .Y(n2222) );
  OAI22X1 U2054 ( .A(n336), .B(n2708), .C(n2709), .D(n386), .Y(n2223) );
  OAI22X1 U2055 ( .A(n336), .B(n2709), .C(n2710), .D(n386), .Y(n2224) );
  OAI22X1 U2056 ( .A(n336), .B(n2710), .C(n2711), .D(n386), .Y(n2225) );
  OAI22X1 U2057 ( .A(n2987), .B(n336), .C(n2712), .D(n386), .Y(n2226) );
  OAI22X1 U2058 ( .A(n336), .B(n2712), .C(n2713), .D(n386), .Y(n2227) );
  OAI22X1 U2059 ( .A(n335), .B(n2713), .C(n2988), .D(n386), .Y(n2228) );
  OAI22X1 U2060 ( .A(n335), .B(n2714), .C(n2715), .D(n385), .Y(n2229) );
  OAI22X1 U2061 ( .A(n335), .B(n2715), .C(n2716), .D(n385), .Y(n2230) );
  OAI22X1 U2062 ( .A(n335), .B(n2716), .C(n2717), .D(n385), .Y(n2231) );
  OAI22X1 U2063 ( .A(n335), .B(n2717), .C(n2718), .D(n385), .Y(n2232) );
  OAI22X1 U2064 ( .A(n335), .B(n2718), .C(n2719), .D(n385), .Y(n2233) );
  OAI22X1 U2065 ( .A(n335), .B(n2719), .C(n2720), .D(n385), .Y(n2234) );
  OAI22X1 U2066 ( .A(n335), .B(n2720), .C(n2721), .D(n385), .Y(n2235) );
  OAI22X1 U2067 ( .A(n335), .B(n2721), .C(n2722), .D(n385), .Y(n2236) );
  OAI22X1 U2068 ( .A(n335), .B(n2722), .C(n2723), .D(n385), .Y(n2237) );
  OAI22X1 U2069 ( .A(n335), .B(n2723), .C(n2724), .D(n385), .Y(n2238) );
  XNOR2X1 U2070 ( .A(n289), .B(n497), .Y(n2693) );
  XNOR2X1 U2071 ( .A(n289), .B(n495), .Y(n2694) );
  XNOR2X1 U2072 ( .A(n289), .B(n493), .Y(n2695) );
  XNOR2X1 U2073 ( .A(n289), .B(n491), .Y(n2696) );
  XNOR2X1 U2074 ( .A(n289), .B(n489), .Y(n2697) );
  XNOR2X1 U2075 ( .A(n289), .B(n487), .Y(n2698) );
  XNOR2X1 U2076 ( .A(n289), .B(n485), .Y(n2699) );
  XNOR2X1 U2077 ( .A(n289), .B(n483), .Y(n2700) );
  XNOR2X1 U2078 ( .A(n289), .B(n481), .Y(n2701) );
  XNOR2X1 U2079 ( .A(n289), .B(n479), .Y(n2702) );
  XNOR2X1 U2080 ( .A(n289), .B(n477), .Y(n2703) );
  XNOR2X1 U2081 ( .A(n288), .B(n475), .Y(n2704) );
  XNOR2X1 U2082 ( .A(n288), .B(n473), .Y(n2705) );
  XNOR2X1 U2083 ( .A(n288), .B(n471), .Y(n2706) );
  XNOR2X1 U2084 ( .A(n288), .B(n469), .Y(n2707) );
  XNOR2X1 U2085 ( .A(n288), .B(n467), .Y(n2708) );
  XNOR2X1 U2088 ( .A(n288), .B(n2974), .Y(n2711) );
  XNOR2X1 U2089 ( .A(n288), .B(n459), .Y(n2712) );
  XNOR2X1 U2090 ( .A(n288), .B(b[11]), .Y(n2713) );
  XNOR2X1 U2091 ( .A(n288), .B(b[10]), .Y(n2714) );
  XNOR2X1 U2092 ( .A(n288), .B(n2969), .Y(n2715) );
  XNOR2X1 U2093 ( .A(n287), .B(b[8]), .Y(n2716) );
  XNOR2X1 U2094 ( .A(n287), .B(b[7]), .Y(n2717) );
  XNOR2X1 U2095 ( .A(n287), .B(n2958), .Y(n2718) );
  XNOR2X1 U2096 ( .A(n287), .B(n2940), .Y(n2719) );
  XNOR2X1 U2097 ( .A(n287), .B(b[4]), .Y(n2720) );
  XNOR2X1 U2098 ( .A(n287), .B(n2995), .Y(n2721) );
  XNOR2X1 U2099 ( .A(n2915), .B(n287), .Y(n2722) );
  XNOR2X1 U2100 ( .A(n287), .B(n2910), .Y(n2723) );
  XNOR2X1 U2101 ( .A(n287), .B(n2944), .Y(n2724) );
  INVX2 U2102 ( .A(n332), .Y(n2796) );
  INVX2 U2104 ( .A(n329), .Y(n2797) );
  INVX2 U2106 ( .A(n326), .Y(n2798) );
  INVX2 U2108 ( .A(n323), .Y(n2799) );
  INVX2 U2110 ( .A(n320), .Y(n2800) );
  INVX2 U2112 ( .A(n317), .Y(n2801) );
  INVX2 U2114 ( .A(n314), .Y(n2802) );
  INVX2 U2116 ( .A(n311), .Y(n2803) );
  INVX2 U2118 ( .A(n308), .Y(n2804) );
  INVX2 U2120 ( .A(n305), .Y(n2805) );
  INVX2 U2122 ( .A(n302), .Y(n2806) );
  INVX2 U2124 ( .A(n299), .Y(n2807) );
  INVX2 U2126 ( .A(n296), .Y(n2808) );
  INVX2 U2128 ( .A(n293), .Y(n2809) );
  INVX2 U2130 ( .A(n290), .Y(n2810) );
  INVX2 U2132 ( .A(n287), .Y(n2811) );
  NAND2X1 U2135 ( .A(n2752), .B(n2780), .Y(n432) );
  XOR2X1 U2136 ( .A(a[30]), .B(a[31]), .Y(n2752) );
  XNOR2X1 U2137 ( .A(a[30]), .B(a[29]), .Y(n2780) );
  NAND2X1 U2138 ( .A(n2753), .B(n2781), .Y(n429) );
  XOR2X1 U2139 ( .A(a[28]), .B(a[29]), .Y(n2753) );
  XNOR2X1 U2140 ( .A(a[28]), .B(a[27]), .Y(n2781) );
  NAND2X1 U2141 ( .A(n2754), .B(n2782), .Y(n426) );
  XOR2X1 U2142 ( .A(a[26]), .B(a[27]), .Y(n2754) );
  XNOR2X1 U2143 ( .A(a[26]), .B(a[25]), .Y(n2782) );
  NAND2X1 U2144 ( .A(n2755), .B(n2783), .Y(n423) );
  XOR2X1 U2145 ( .A(a[24]), .B(a[25]), .Y(n2755) );
  XNOR2X1 U2146 ( .A(a[24]), .B(a[23]), .Y(n2783) );
  NAND2X1 U2147 ( .A(n2756), .B(n2784), .Y(n2768) );
  XOR2X1 U2148 ( .A(a[22]), .B(a[23]), .Y(n2756) );
  XNOR2X1 U2149 ( .A(a[22]), .B(a[21]), .Y(n2784) );
  NAND2X1 U2150 ( .A(n2757), .B(n2785), .Y(n2769) );
  XOR2X1 U2151 ( .A(a[20]), .B(a[21]), .Y(n2757) );
  XNOR2X1 U2152 ( .A(a[20]), .B(a[19]), .Y(n2785) );
  NAND2X1 U2153 ( .A(n2758), .B(n2786), .Y(n2770) );
  XOR2X1 U2154 ( .A(a[18]), .B(a[19]), .Y(n2758) );
  XNOR2X1 U2155 ( .A(a[18]), .B(a[17]), .Y(n2786) );
  NAND2X1 U2156 ( .A(n2759), .B(n2787), .Y(n2771) );
  XOR2X1 U2157 ( .A(a[16]), .B(a[17]), .Y(n2759) );
  XNOR2X1 U2158 ( .A(a[16]), .B(a[15]), .Y(n2787) );
  NAND2X1 U2159 ( .A(n2760), .B(n2788), .Y(n2772) );
  XOR2X1 U2160 ( .A(a[14]), .B(a[15]), .Y(n2760) );
  XNOR2X1 U2161 ( .A(a[14]), .B(a[13]), .Y(n2788) );
  NAND2X1 U2162 ( .A(n2761), .B(n2789), .Y(n2773) );
  XOR2X1 U2163 ( .A(a[12]), .B(a[13]), .Y(n2761) );
  XNOR2X1 U2164 ( .A(a[12]), .B(a[11]), .Y(n2789) );
  NAND2X1 U2165 ( .A(n2762), .B(n2790), .Y(n2774) );
  XOR2X1 U2166 ( .A(a[10]), .B(a[11]), .Y(n2762) );
  XNOR2X1 U2167 ( .A(a[10]), .B(a[9]), .Y(n2790) );
  NAND2X1 U2168 ( .A(n2763), .B(n2791), .Y(n2775) );
  XOR2X1 U2169 ( .A(a[8]), .B(a[9]), .Y(n2763) );
  XNOR2X1 U2170 ( .A(a[8]), .B(a[7]), .Y(n2791) );
  NAND2X1 U2171 ( .A(n2764), .B(n2792), .Y(n2776) );
  XOR2X1 U2172 ( .A(a[6]), .B(a[7]), .Y(n2764) );
  XNOR2X1 U2173 ( .A(a[6]), .B(a[5]), .Y(n2792) );
  NAND2X1 U2174 ( .A(n2765), .B(n2793), .Y(n2777) );
  XOR2X1 U2175 ( .A(a[4]), .B(a[5]), .Y(n2765) );
  XNOR2X1 U2176 ( .A(a[4]), .B(a[3]), .Y(n2793) );
  NAND2X1 U2177 ( .A(n2766), .B(n2794), .Y(n2778) );
  XOR2X1 U2178 ( .A(a[2]), .B(a[3]), .Y(n2766) );
  XNOR2X1 U2179 ( .A(a[2]), .B(a[1]), .Y(n2794) );
  NAND2X1 U2180 ( .A(n2795), .B(n2767), .Y(n2779) );
  XOR2X1 U2181 ( .A(a[0]), .B(a[1]), .Y(n2767) );
  INVX2 U2182 ( .A(a[0]), .Y(n2795) );
  INVX1 U2185 ( .A(n789), .Y(n878) );
  BUFX4 U2186 ( .A(b[6]), .Y(n2959) );
  BUFX4 U2187 ( .A(b[17]), .Y(n469) );
  INVX4 U2188 ( .A(n2966), .Y(n2940) );
  INVX4 U2189 ( .A(b[5]), .Y(n2966) );
  INVX8 U2190 ( .A(n2986), .Y(n2909) );
  INVX8 U2191 ( .A(n2909), .Y(n2910) );
  INVX8 U2192 ( .A(n2909), .Y(n2911) );
  INVX2 U2193 ( .A(n2984), .Y(n2985) );
  INVX2 U2194 ( .A(n2966), .Y(n2967) );
  INVX2 U2195 ( .A(b[1]), .Y(n2984) );
  INVX4 U2196 ( .A(n2984), .Y(n2986) );
  BUFX2 U2197 ( .A(n461), .Y(n2976) );
  BUFX2 U2198 ( .A(n2945), .Y(n2912) );
  BUFX2 U2199 ( .A(n2945), .Y(n2913) );
  INVX1 U2200 ( .A(n2999), .Y(n2945) );
  BUFX2 U2201 ( .A(b[2]), .Y(n2914) );
  BUFX4 U2202 ( .A(b[2]), .Y(n2915) );
  OR2X2 U2203 ( .A(n1615), .B(n1600), .Y(n2916) );
  OR2X2 U2204 ( .A(n1431), .B(n1406), .Y(n2917) );
  INVX2 U2205 ( .A(b[10]), .Y(n2977) );
  OR2X2 U2206 ( .A(n1631), .B(n1616), .Y(n2918) );
  OR2X2 U2207 ( .A(n1741), .B(n1740), .Y(n2919) );
  OR2X2 U2208 ( .A(n1719), .B(n1712), .Y(n2920) );
  OR2X2 U2209 ( .A(n1703), .B(n1694), .Y(n2921) );
  OR2X2 U2210 ( .A(n2237), .B(n2954), .Y(n2922) );
  OR2X2 U2211 ( .A(n1479), .B(n1456), .Y(n2923) );
  OR2X2 U2212 ( .A(n1455), .B(n1432), .Y(n2924) );
  OR2X2 U2213 ( .A(n920), .B(n901), .Y(n2925) );
  INVX2 U2214 ( .A(b[11]), .Y(n2963) );
  AND2X2 U2215 ( .A(n2998), .B(n152), .Y(n2926) );
  AND2X2 U2216 ( .A(n2944), .B(n125), .Y(n2927) );
  AND2X2 U2217 ( .A(n2944), .B(a[0]), .Y(product[0]) );
  OR2X2 U2218 ( .A(n1758), .B(n2238), .Y(n2929) );
  AND2X2 U2219 ( .A(n2941), .B(n98), .Y(n2930) );
  INVX2 U2220 ( .A(b[7]), .Y(n2992) );
  INVX2 U2221 ( .A(n2972), .Y(n2973) );
  INVX2 U2222 ( .A(b[8]), .Y(n2972) );
  OR2X2 U2223 ( .A(n900), .B(n891), .Y(n2931) );
  XOR2X1 U2224 ( .A(n1691), .B(n1689), .Y(n2932) );
  XOR2X1 U2225 ( .A(n1682), .B(n2932), .Y(n1676) );
  NAND2X1 U2226 ( .A(n1682), .B(n1691), .Y(n2933) );
  NAND2X1 U2227 ( .A(n1682), .B(n1689), .Y(n2934) );
  NAND2X1 U2228 ( .A(n1691), .B(n1689), .Y(n2935) );
  NAND3X1 U2229 ( .A(n2933), .B(n2934), .C(n2935), .Y(n1675) );
  XOR2X1 U2230 ( .A(n1656), .B(n1667), .Y(n2936) );
  XOR2X1 U2231 ( .A(n1654), .B(n2936), .Y(n1650) );
  NAND2X1 U2232 ( .A(n1654), .B(n1656), .Y(n2937) );
  NAND2X1 U2233 ( .A(n1654), .B(n1667), .Y(n2938) );
  NAND2X1 U2234 ( .A(n1656), .B(n1667), .Y(n2939) );
  NAND3X1 U2235 ( .A(n2937), .B(n2938), .C(n2939), .Y(n1649) );
  BUFX4 U2236 ( .A(b[9]), .Y(n453) );
  INVX2 U2237 ( .A(n2999), .Y(n2941) );
  BUFX2 U2238 ( .A(b[3]), .Y(n2995) );
  BUFX4 U2239 ( .A(n433), .Y(n2944) );
  INVX8 U2240 ( .A(n433), .Y(n2999) );
  INVX4 U2241 ( .A(n2999), .Y(n2997) );
  XNOR2X1 U2242 ( .A(n780), .B(n2942), .Y(product[15]) );
  AND2X2 U2243 ( .A(n779), .B(n876), .Y(n2942) );
  BUFX4 U2244 ( .A(b[12]), .Y(n459) );
  BUFX4 U2245 ( .A(b[3]), .Y(n441) );
  INVX4 U2246 ( .A(n2977), .Y(n2978) );
  BUFX4 U2247 ( .A(n441), .Y(n2979) );
  BUFX2 U2248 ( .A(b[3]), .Y(n2943) );
  BUFX4 U2249 ( .A(b[0]), .Y(n433) );
  INVX1 U2250 ( .A(n2992), .Y(n2994) );
  INVX4 U2251 ( .A(n2966), .Y(n2968) );
  INVX1 U2252 ( .A(n745), .Y(n743) );
  INVX1 U2253 ( .A(n746), .Y(n744) );
  INVX1 U2254 ( .A(n2918), .Y(n761) );
  BUFX4 U2255 ( .A(n453), .Y(n2970) );
  AND2X2 U2256 ( .A(n2941), .B(n143), .Y(n2948) );
  XNOR2X1 U2257 ( .A(n288), .B(n465), .Y(n2709) );
  XNOR2X1 U2258 ( .A(n288), .B(n463), .Y(n2710) );
  AND2X2 U2259 ( .A(n2941), .B(n178), .Y(n2950) );
  AND2X2 U2260 ( .A(n2998), .B(n226), .Y(n2953) );
  AND2X2 U2261 ( .A(n2941), .B(n258), .Y(n2954) );
  AND2X2 U2262 ( .A(n843), .B(n2929), .Y(product[1]) );
  INVX2 U2263 ( .A(n601), .Y(n595) );
  INVX2 U2264 ( .A(n581), .Y(n579) );
  INVX2 U2265 ( .A(n677), .Y(n676) );
  INVX2 U2266 ( .A(n698), .Y(n697) );
  INVX2 U2267 ( .A(n649), .Y(n647) );
  INVX2 U2268 ( .A(n634), .Y(n632) );
  INVX2 U2269 ( .A(n633), .Y(n631) );
  INVX2 U2270 ( .A(n669), .Y(n663) );
  INVX2 U2271 ( .A(n602), .Y(n600) );
  INVX2 U2272 ( .A(n582), .Y(n580) );
  OR2X2 U2273 ( .A(n554), .B(n581), .Y(n2946) );
  INVX2 U2274 ( .A(n727), .Y(n726) );
  INVX2 U2275 ( .A(n748), .Y(n747) );
  INVX2 U2276 ( .A(n695), .Y(n693) );
  INVX2 U2277 ( .A(n696), .Y(n694) );
  INVX2 U2278 ( .A(n650), .Y(n648) );
  INVX2 U2279 ( .A(n642), .Y(n640) );
  INVX2 U2280 ( .A(n643), .Y(n641) );
  INVX2 U2281 ( .A(n670), .Y(n668) );
  BUFX2 U2282 ( .A(n608), .Y(n499) );
  INVX2 U2283 ( .A(n592), .Y(n590) );
  INVX2 U2284 ( .A(n574), .Y(n572) );
  INVX2 U2285 ( .A(n593), .Y(n591) );
  INVX2 U2286 ( .A(n575), .Y(n573) );
  INVX1 U2287 ( .A(n759), .Y(n757) );
  INVX2 U2288 ( .A(n718), .Y(n716) );
  INVX2 U2289 ( .A(n768), .Y(n767) );
  INVX2 U2290 ( .A(n786), .Y(n785) );
  INVX2 U2291 ( .A(n725), .Y(n723) );
  INVX2 U2292 ( .A(n711), .Y(n709) );
  INVX2 U2293 ( .A(n706), .Y(n704) );
  INVX2 U2294 ( .A(n660), .Y(n658) );
  INVX2 U2295 ( .A(n661), .Y(n659) );
  INVX2 U2296 ( .A(n553), .Y(n551) );
  INVX2 U2297 ( .A(n559), .Y(n557) );
  INVX2 U2298 ( .A(n2242), .Y(n2991) );
  INVX1 U2299 ( .A(n774), .Y(n772) );
  INVX2 U2300 ( .A(n2999), .Y(n2998) );
  INVX1 U2301 ( .A(n766), .Y(n764) );
  INVX1 U2302 ( .A(n783), .Y(n781) );
  INVX1 U2303 ( .A(n784), .Y(n782) );
  INVX2 U2304 ( .A(n773), .Y(n771) );
  INVX1 U2305 ( .A(n801), .Y(n799) );
  BUFX2 U2306 ( .A(n463), .Y(n2962) );
  BUFX2 U2307 ( .A(n461), .Y(n2975) );
  BUFX2 U2308 ( .A(b[6]), .Y(n2960) );
  INVX4 U2309 ( .A(n2250), .Y(n2996) );
  BUFX2 U2310 ( .A(n2943), .Y(n2980) );
  BUFX2 U2311 ( .A(n2943), .Y(n2981) );
  INVX1 U2312 ( .A(n812), .Y(n810) );
  INVX2 U2313 ( .A(n2963), .Y(n2964) );
  INVX2 U2314 ( .A(n2963), .Y(n2965) );
  INVX2 U2315 ( .A(n2992), .Y(n2993) );
  BUFX2 U2316 ( .A(b[6]), .Y(n2958) );
  BUFX2 U2317 ( .A(n453), .Y(n2969) );
  BUFX4 U2318 ( .A(b[16]), .Y(n467) );
  BUFX2 U2319 ( .A(b[19]), .Y(n473) );
  BUFX4 U2320 ( .A(b[18]), .Y(n471) );
  BUFX2 U2321 ( .A(b[20]), .Y(n475) );
  BUFX2 U2322 ( .A(b[21]), .Y(n477) );
  BUFX2 U2323 ( .A(b[23]), .Y(n481) );
  BUFX2 U2324 ( .A(b[22]), .Y(n479) );
  BUFX2 U2325 ( .A(b[24]), .Y(n483) );
  INVX1 U2326 ( .A(n832), .Y(n830) );
  INVX1 U2327 ( .A(n840), .Y(n838) );
  INVX2 U2328 ( .A(n843), .Y(n841) );
  BUFX2 U2329 ( .A(b[15]), .Y(n465) );
  BUFX2 U2330 ( .A(b[27]), .Y(n489) );
  BUFX2 U2331 ( .A(b[26]), .Y(n487) );
  BUFX2 U2332 ( .A(b[30]), .Y(n495) );
  BUFX2 U2333 ( .A(b[28]), .Y(n491) );
  AND2X1 U2334 ( .A(n2913), .B(n134), .Y(n2947) );
  AND2X1 U2335 ( .A(n2941), .B(n168), .Y(n2949) );
  AND2X1 U2336 ( .A(n2944), .B(n216), .Y(n2951) );
  AND2X1 U2337 ( .A(n2944), .B(n116), .Y(n2952) );
  AND2X1 U2338 ( .A(n2913), .B(n89), .Y(n2955) );
  AND2X1 U2339 ( .A(n2941), .B(n107), .Y(n2956) );
  BUFX2 U2340 ( .A(n334), .Y(n332) );
  BUFX2 U2341 ( .A(n2796), .Y(n383) );
  BUFX2 U2342 ( .A(n334), .Y(n333) );
  BUFX2 U2343 ( .A(n2817), .Y(n310) );
  BUFX2 U2344 ( .A(n2816), .Y(n313) );
  BUFX2 U2345 ( .A(n2816), .Y(n311) );
  BUFX2 U2346 ( .A(n2814), .Y(n317) );
  BUFX2 U2347 ( .A(n2815), .Y(n314) );
  BUFX2 U2348 ( .A(n2817), .Y(n308) );
  BUFX2 U2349 ( .A(n2818), .Y(n305) );
  BUFX2 U2350 ( .A(n2813), .Y(n320) );
  BUFX2 U2351 ( .A(n2815), .Y(n316) );
  BUFX2 U2352 ( .A(n2814), .Y(n319) );
  BUFX2 U2353 ( .A(n2773), .Y(n405) );
  BUFX2 U2354 ( .A(n2772), .Y(n408) );
  BUFX2 U2355 ( .A(n2787), .Y(n359) );
  BUFX2 U2356 ( .A(n2773), .Y(n403) );
  BUFX2 U2357 ( .A(n2772), .Y(n406) );
  BUFX2 U2358 ( .A(n2771), .Y(n409) );
  BUFX2 U2359 ( .A(n2770), .Y(n412) );
  BUFX2 U2360 ( .A(n2769), .Y(n415) );
  BUFX2 U2361 ( .A(n2771), .Y(n411) );
  BUFX2 U2362 ( .A(n2813), .Y(n322) );
  BUFX2 U2363 ( .A(n2770), .Y(n414) );
  BUFX2 U2364 ( .A(n2769), .Y(n417) );
  BUFX2 U2365 ( .A(n2768), .Y(n420) );
  BUFX2 U2366 ( .A(n2821), .Y(n297) );
  BUFX2 U2367 ( .A(n2820), .Y(n300) );
  BUFX2 U2368 ( .A(n2818), .Y(n306) );
  BUFX2 U2369 ( .A(n2818), .Y(n307) );
  BUFX2 U2370 ( .A(n2821), .Y(n298) );
  BUFX2 U2371 ( .A(n2820), .Y(n301) );
  BUFX2 U2372 ( .A(n2819), .Y(n304) );
  BUFX2 U2373 ( .A(n331), .Y(n329) );
  BUFX2 U2374 ( .A(n2820), .Y(n299) );
  BUFX2 U2375 ( .A(n2822), .Y(n293) );
  BUFX2 U2376 ( .A(n2821), .Y(n296) );
  BUFX2 U2377 ( .A(n2819), .Y(n302) );
  BUFX2 U2378 ( .A(n2812), .Y(n323) );
  BUFX2 U2379 ( .A(n328), .Y(n326) );
  BUFX2 U2380 ( .A(n2776), .Y(n396) );
  BUFX2 U2381 ( .A(n2775), .Y(n399) );
  BUFX2 U2382 ( .A(n2774), .Y(n402) );
  BUFX2 U2383 ( .A(n2792), .Y(n346) );
  BUFX2 U2384 ( .A(n2791), .Y(n349) );
  BUFX2 U2385 ( .A(n2790), .Y(n352) );
  BUFX2 U2386 ( .A(n2789), .Y(n355) );
  BUFX2 U2387 ( .A(n2788), .Y(n358) );
  BUFX2 U2388 ( .A(n2792), .Y(n344) );
  BUFX2 U2389 ( .A(n2791), .Y(n347) );
  BUFX2 U2390 ( .A(n2790), .Y(n350) );
  BUFX2 U2391 ( .A(n2789), .Y(n353) );
  BUFX2 U2392 ( .A(n2788), .Y(n356) );
  BUFX2 U2393 ( .A(n2786), .Y(n362) );
  BUFX2 U2394 ( .A(n2785), .Y(n365) );
  BUFX2 U2395 ( .A(n2784), .Y(n368) );
  BUFX2 U2396 ( .A(n2783), .Y(n371) );
  BUFX2 U2397 ( .A(n2782), .Y(n374) );
  BUFX2 U2398 ( .A(n2781), .Y(n377) );
  BUFX2 U2399 ( .A(n2780), .Y(n380) );
  BUFX2 U2400 ( .A(n2777), .Y(n391) );
  BUFX2 U2401 ( .A(n2776), .Y(n394) );
  BUFX2 U2402 ( .A(n2775), .Y(n397) );
  BUFX2 U2403 ( .A(n2774), .Y(n400) );
  BUFX2 U2404 ( .A(n2768), .Y(n418) );
  BUFX2 U2405 ( .A(n423), .Y(n421) );
  BUFX2 U2406 ( .A(n426), .Y(n424) );
  BUFX2 U2407 ( .A(n429), .Y(n427) );
  BUFX2 U2408 ( .A(n432), .Y(n430) );
  BUFX2 U2409 ( .A(n2787), .Y(n361) );
  BUFX2 U2410 ( .A(n2786), .Y(n364) );
  BUFX2 U2411 ( .A(n2785), .Y(n367) );
  BUFX2 U2412 ( .A(n2812), .Y(n325) );
  BUFX2 U2413 ( .A(a[31]), .Y(n334) );
  BUFX2 U2414 ( .A(n2784), .Y(n370) );
  BUFX2 U2415 ( .A(n2783), .Y(n373) );
  BUFX2 U2416 ( .A(n2782), .Y(n376) );
  BUFX2 U2417 ( .A(n2781), .Y(n379) );
  BUFX2 U2418 ( .A(n2780), .Y(n382) );
  BUFX2 U2419 ( .A(n2824), .Y(n288) );
  BUFX2 U2420 ( .A(n2822), .Y(n294) );
  BUFX2 U2421 ( .A(n2823), .Y(n291) );
  BUFX2 U2422 ( .A(n2819), .Y(n303) );
  BUFX2 U2423 ( .A(n2817), .Y(n309) );
  BUFX2 U2424 ( .A(n2816), .Y(n312) );
  BUFX2 U2425 ( .A(n2815), .Y(n315) );
  BUFX2 U2426 ( .A(n2813), .Y(n321) );
  BUFX2 U2427 ( .A(n2814), .Y(n318) );
  BUFX2 U2428 ( .A(n2812), .Y(n324) );
  BUFX2 U2429 ( .A(n328), .Y(n327) );
  BUFX2 U2430 ( .A(n2822), .Y(n295) );
  BUFX2 U2431 ( .A(n2824), .Y(n289) );
  BUFX2 U2432 ( .A(n2823), .Y(n292) );
  BUFX2 U2433 ( .A(n331), .Y(n330) );
  BUFX2 U2434 ( .A(n2824), .Y(n287) );
  BUFX2 U2435 ( .A(n2823), .Y(n290) );
  BUFX2 U2436 ( .A(n2778), .Y(n390) );
  BUFX2 U2437 ( .A(n2777), .Y(n393) );
  BUFX2 U2438 ( .A(n2778), .Y(n389) );
  BUFX2 U2439 ( .A(n2777), .Y(n392) );
  BUFX2 U2440 ( .A(n2776), .Y(n395) );
  BUFX2 U2441 ( .A(n2775), .Y(n398) );
  BUFX2 U2442 ( .A(n2774), .Y(n401) );
  BUFX2 U2443 ( .A(n2773), .Y(n404) );
  BUFX2 U2444 ( .A(n2772), .Y(n407) );
  BUFX2 U2445 ( .A(n2771), .Y(n410) );
  BUFX2 U2446 ( .A(n2770), .Y(n413) );
  BUFX2 U2447 ( .A(n2769), .Y(n416) );
  BUFX2 U2448 ( .A(n2768), .Y(n419) );
  BUFX2 U2449 ( .A(n423), .Y(n422) );
  BUFX2 U2450 ( .A(n2794), .Y(n339) );
  BUFX2 U2451 ( .A(n2792), .Y(n345) );
  BUFX2 U2452 ( .A(n2793), .Y(n342) );
  BUFX2 U2453 ( .A(n2791), .Y(n348) );
  BUFX2 U2454 ( .A(n2790), .Y(n351) );
  BUFX2 U2455 ( .A(n2789), .Y(n354) );
  BUFX2 U2456 ( .A(n2794), .Y(n340) );
  BUFX2 U2457 ( .A(n2793), .Y(n343) );
  BUFX2 U2458 ( .A(n2793), .Y(n341) );
  BUFX2 U2459 ( .A(n2794), .Y(n338) );
  BUFX2 U2460 ( .A(n2778), .Y(n388) );
  BUFX2 U2461 ( .A(n2788), .Y(n357) );
  BUFX2 U2462 ( .A(n2787), .Y(n360) );
  BUFX2 U2463 ( .A(n2786), .Y(n363) );
  BUFX2 U2464 ( .A(n2785), .Y(n366) );
  BUFX2 U2465 ( .A(n2784), .Y(n369) );
  BUFX2 U2466 ( .A(n2783), .Y(n372) );
  BUFX2 U2467 ( .A(n426), .Y(n425) );
  BUFX2 U2468 ( .A(n2782), .Y(n375) );
  BUFX2 U2469 ( .A(n429), .Y(n428) );
  BUFX2 U2470 ( .A(n432), .Y(n431) );
  BUFX2 U2471 ( .A(n2781), .Y(n378) );
  BUFX2 U2472 ( .A(n2780), .Y(n381) );
  BUFX2 U2473 ( .A(a[21]), .Y(n2814) );
  BUFX2 U2474 ( .A(a[23]), .Y(n2813) );
  BUFX2 U2475 ( .A(a[15]), .Y(n2817) );
  BUFX2 U2476 ( .A(a[13]), .Y(n2818) );
  BUFX2 U2477 ( .A(a[17]), .Y(n2816) );
  BUFX2 U2478 ( .A(a[19]), .Y(n2815) );
  BUFX2 U2479 ( .A(a[27]), .Y(n328) );
  BUFX2 U2480 ( .A(a[25]), .Y(n2812) );
  BUFX2 U2481 ( .A(a[5]), .Y(n2822) );
  BUFX2 U2482 ( .A(a[7]), .Y(n2821) );
  BUFX2 U2483 ( .A(a[9]), .Y(n2820) );
  BUFX2 U2484 ( .A(a[11]), .Y(n2819) );
  BUFX2 U2485 ( .A(a[29]), .Y(n331) );
  BUFX2 U2486 ( .A(n2779), .Y(n387) );
  BUFX2 U2487 ( .A(n2779), .Y(n386) );
  BUFX2 U2488 ( .A(n2795), .Y(n337) );
  BUFX2 U2489 ( .A(n2795), .Y(n336) );
  BUFX2 U2490 ( .A(n2795), .Y(n335) );
  BUFX2 U2491 ( .A(n2779), .Y(n385) );
  BUFX2 U2492 ( .A(a[1]), .Y(n2824) );
  BUFX2 U2493 ( .A(a[3]), .Y(n2823) );
  BUFX2 U2494 ( .A(n463), .Y(n2961) );
  BUFX2 U2495 ( .A(b[14]), .Y(n463) );
  BUFX2 U2496 ( .A(n453), .Y(n2971) );
  BUFX2 U2497 ( .A(b[31]), .Y(n497) );
  BUFX2 U2498 ( .A(n461), .Y(n2974) );
  BUFX2 U2499 ( .A(b[13]), .Y(n461) );
  BUFX2 U2500 ( .A(n465), .Y(n2982) );
  BUFX2 U2501 ( .A(n465), .Y(n2983) );
  INVX1 U2502 ( .A(n2982), .Y(n2239) );
  XNOR2X1 U2503 ( .A(n288), .B(n2974), .Y(n2987) );
  INVX1 U2504 ( .A(n2961), .Y(n2240) );
  XNOR2X1 U2505 ( .A(n288), .B(b[10]), .Y(n2988) );
  INVX1 U2506 ( .A(n2975), .Y(n2241) );
  INVX1 U2507 ( .A(n778), .Y(n876) );
  BUFX2 U2508 ( .A(b[25]), .Y(n485) );
  INVX2 U2509 ( .A(n806), .Y(n804) );
  BUFX2 U2510 ( .A(n823), .Y(n2989) );
  INVX1 U2511 ( .A(n885), .Y(n2990) );
  INVX1 U2512 ( .A(n459), .Y(n2242) );
  INVX2 U2513 ( .A(n805), .Y(n803) );
  INVX1 U2514 ( .A(n2978), .Y(n2244) );
  INVX1 U2515 ( .A(n2959), .Y(n2248) );
  INVX1 U2516 ( .A(n2970), .Y(n2245) );
  BUFX2 U2517 ( .A(n2915), .Y(n439) );
  INVX1 U2518 ( .A(n2964), .Y(n2243) );
  INVX1 U2519 ( .A(n792), .Y(n879) );
  INVX1 U2520 ( .A(n825), .Y(n824) );
  INVX1 U2521 ( .A(n822), .Y(n885) );
  INVX1 U2522 ( .A(n2980), .Y(n2251) );
  INVX1 U2523 ( .A(n433), .Y(n3000) );
  BUFX2 U2524 ( .A(b[29]), .Y(n493) );
  INVX1 U2525 ( .A(n808), .Y(n807) );
  INVX1 U2526 ( .A(n795), .Y(n794) );
  INVX1 U2527 ( .A(n819), .Y(n884) );
endmodule


module poly5_DW_mult_uns_49 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n68, n72, n76, n80, n95, n103, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n150, n151, n152, n154, n155, n157, n159, n160, n161, n162, n163,
         n164, n166, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n180, n181, n182, n183, n184, n185, n186, n187, n189,
         n191, n192, n193, n194, n195, n196, n197, n198, n202, n204, n205,
         n206, n207, n208, n209, n210, n211, n213, n216, n217, n218, n219,
         n220, n221, n222, n225, n226, n227, n228, n229, n231, n232, n233,
         n234, n235, n236, n237, n238, n241, n242, n243, n244, n245, n246,
         n247, n249, n250, n251, n252, n253, n254, n255, n256, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n280, n281, n282, n283, n284, n285, n288,
         n289, n290, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n302, n304, n305, n306, n307, n311, n313, n314, n315, n316, n317,
         n318, n322, n324, n325, n326, n327, n332, n333, n334, n335, n337,
         n339, n340, n341, n342, n343, n344, n345, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n360, n362, n363,
         n364, n365, n367, n370, n371, n372, n373, n375, n377, n378, n380,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n419, n420, n421, n422, n427, n428, n429, n430,
         n435, n436, n437, n438, n446, n448, n450, n451, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n468, n470, n471,
         n472, n474, n477, n478, n479, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1675, n1705, n1783, n1784, n1785,
         n1786, n1787, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1878, n1879, n1880, n1881, n1882, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004;

  NAND2X1 U85 ( .A(n154), .B(n1884), .Y(n121) );
  NAND2X1 U88 ( .A(n486), .B(n479), .Y(n154) );
  XNOR2X1 U89 ( .A(n162), .B(n122), .Y(product[46]) );
  OAI21X1 U90 ( .A(n1890), .B(n1913), .C(n157), .Y(n155) );
  OAI21X1 U94 ( .A(n160), .B(n164), .C(n161), .Y(n159) );
  NAND2X1 U95 ( .A(n161), .B(n448), .Y(n122) );
  NOR2X1 U97 ( .A(n502), .B(n487), .Y(n160) );
  NAND2X1 U98 ( .A(n502), .B(n487), .Y(n161) );
  XNOR2X1 U99 ( .A(n169), .B(n123), .Y(product[45]) );
  OAI21X1 U100 ( .A(n163), .B(n1913), .C(n164), .Y(n162) );
  NAND2X1 U101 ( .A(n1894), .B(n172), .Y(n163) );
  AOI21X1 U102 ( .A(n1894), .B(n173), .C(n166), .Y(n164) );
  NAND2X1 U105 ( .A(n168), .B(n1894), .Y(n123) );
  NAND2X1 U108 ( .A(n518), .B(n503), .Y(n168) );
  XNOR2X1 U109 ( .A(n176), .B(n124), .Y(product[44]) );
  OAI21X1 U110 ( .A(n170), .B(n1913), .C(n171), .Y(n169) );
  NOR2X1 U113 ( .A(n174), .B(n177), .Y(n172) );
  OAI21X1 U114 ( .A(n178), .B(n174), .C(n175), .Y(n173) );
  NAND2X1 U115 ( .A(n175), .B(n450), .Y(n124) );
  NOR2X1 U117 ( .A(n536), .B(n519), .Y(n174) );
  NAND2X1 U118 ( .A(n536), .B(n519), .Y(n175) );
  XOR2X1 U119 ( .A(n1913), .B(n125), .Y(product[43]) );
  OAI21X1 U120 ( .A(n177), .B(n1913), .C(n178), .Y(n176) );
  NAND2X1 U121 ( .A(n178), .B(n451), .Y(n125) );
  NOR2X1 U123 ( .A(n554), .B(n537), .Y(n177) );
  NAND2X1 U124 ( .A(n554), .B(n537), .Y(n178) );
  XNOR2X1 U125 ( .A(n192), .B(n126), .Y(product[42]) );
  AOI21X1 U126 ( .A(n267), .B(n180), .C(n181), .Y(n120) );
  NOR2X1 U127 ( .A(n182), .B(n235), .Y(n180) );
  OAI21X1 U128 ( .A(n182), .B(n236), .C(n183), .Y(n181) );
  NAND2X1 U129 ( .A(n184), .B(n219), .Y(n182) );
  AOI21X1 U130 ( .A(n220), .B(n184), .C(n185), .Y(n183) );
  NOR2X1 U131 ( .A(n210), .B(n186), .Y(n184) );
  OAI21X1 U132 ( .A(n211), .B(n186), .C(n187), .Y(n185) );
  NAND2X1 U133 ( .A(n1895), .B(n1891), .Y(n186) );
  AOI21X1 U134 ( .A(n1895), .B(n202), .C(n189), .Y(n187) );
  NAND2X1 U137 ( .A(n191), .B(n1895), .Y(n126) );
  NAND2X1 U140 ( .A(n574), .B(n555), .Y(n191) );
  XNOR2X1 U141 ( .A(n205), .B(n127), .Y(product[41]) );
  OAI21X1 U142 ( .A(n266), .B(n193), .C(n194), .Y(n192) );
  NAND2X1 U143 ( .A(n195), .B(n237), .Y(n193) );
  AOI21X1 U144 ( .A(n195), .B(n238), .C(n196), .Y(n194) );
  NOR2X1 U145 ( .A(n197), .B(n221), .Y(n195) );
  OAI21X1 U146 ( .A(n197), .B(n222), .C(n198), .Y(n196) );
  NAND2X1 U147 ( .A(n1891), .B(n454), .Y(n197) );
  AOI21X1 U148 ( .A(n1891), .B(n213), .C(n202), .Y(n198) );
  NAND2X1 U153 ( .A(n204), .B(n1891), .Y(n127) );
  NAND2X1 U156 ( .A(n575), .B(n594), .Y(n204) );
  XNOR2X1 U157 ( .A(n216), .B(n128), .Y(product[40]) );
  OAI21X1 U158 ( .A(n266), .B(n206), .C(n207), .Y(n205) );
  NAND2X1 U159 ( .A(n208), .B(n237), .Y(n206) );
  AOI21X1 U160 ( .A(n238), .B(n208), .C(n209), .Y(n207) );
  NOR2X1 U161 ( .A(n210), .B(n221), .Y(n208) );
  OAI21X1 U162 ( .A(n210), .B(n222), .C(n211), .Y(n209) );
  NAND2X1 U167 ( .A(n211), .B(n454), .Y(n128) );
  NOR2X1 U169 ( .A(n616), .B(n595), .Y(n210) );
  NAND2X1 U170 ( .A(n616), .B(n595), .Y(n211) );
  XNOR2X1 U171 ( .A(n227), .B(n129), .Y(product[39]) );
  OAI21X1 U172 ( .A(n266), .B(n217), .C(n218), .Y(n216) );
  NAND2X1 U173 ( .A(n219), .B(n237), .Y(n217) );
  AOI21X1 U174 ( .A(n219), .B(n238), .C(n220), .Y(n218) );
  NOR2X1 U179 ( .A(n225), .B(n232), .Y(n219) );
  OAI21X1 U180 ( .A(n233), .B(n225), .C(n226), .Y(n220) );
  NAND2X1 U181 ( .A(n226), .B(n455), .Y(n129) );
  NOR2X1 U183 ( .A(n638), .B(n617), .Y(n225) );
  NAND2X1 U184 ( .A(n638), .B(n617), .Y(n226) );
  XNOR2X1 U185 ( .A(n234), .B(n130), .Y(product[38]) );
  OAI21X1 U186 ( .A(n266), .B(n228), .C(n229), .Y(n227) );
  NAND2X1 U187 ( .A(n456), .B(n237), .Y(n228) );
  AOI21X1 U188 ( .A(n456), .B(n238), .C(n231), .Y(n229) );
  NAND2X1 U191 ( .A(n233), .B(n456), .Y(n130) );
  NOR2X1 U193 ( .A(n662), .B(n639), .Y(n232) );
  NAND2X1 U194 ( .A(n662), .B(n639), .Y(n233) );
  XNOR2X1 U195 ( .A(n245), .B(n131), .Y(product[37]) );
  OAI21X1 U196 ( .A(n235), .B(n266), .C(n236), .Y(n234) );
  NAND2X1 U201 ( .A(n241), .B(n255), .Y(n235) );
  AOI21X1 U202 ( .A(n241), .B(n256), .C(n242), .Y(n236) );
  NOR2X1 U203 ( .A(n243), .B(n250), .Y(n241) );
  OAI21X1 U204 ( .A(n251), .B(n243), .C(n244), .Y(n242) );
  NAND2X1 U205 ( .A(n244), .B(n457), .Y(n131) );
  NOR2X1 U207 ( .A(n686), .B(n663), .Y(n243) );
  NAND2X1 U208 ( .A(n686), .B(n663), .Y(n244) );
  XNOR2X1 U209 ( .A(n252), .B(n132), .Y(product[36]) );
  OAI21X1 U210 ( .A(n246), .B(n266), .C(n247), .Y(n245) );
  NAND2X1 U211 ( .A(n458), .B(n255), .Y(n246) );
  AOI21X1 U212 ( .A(n458), .B(n256), .C(n249), .Y(n247) );
  NAND2X1 U215 ( .A(n251), .B(n458), .Y(n132) );
  NOR2X1 U217 ( .A(n712), .B(n687), .Y(n250) );
  NAND2X1 U218 ( .A(n712), .B(n687), .Y(n251) );
  XNOR2X1 U219 ( .A(n263), .B(n133), .Y(product[35]) );
  OAI21X1 U220 ( .A(n253), .B(n266), .C(n254), .Y(n252) );
  NOR2X1 U227 ( .A(n264), .B(n261), .Y(n255) );
  OAI21X1 U228 ( .A(n265), .B(n261), .C(n262), .Y(n256) );
  NAND2X1 U229 ( .A(n262), .B(n459), .Y(n133) );
  NOR2X1 U231 ( .A(n738), .B(n713), .Y(n261) );
  NAND2X1 U232 ( .A(n738), .B(n713), .Y(n262) );
  XOR2X1 U233 ( .A(n266), .B(n134), .Y(product[34]) );
  OAI21X1 U234 ( .A(n264), .B(n266), .C(n265), .Y(n263) );
  NAND2X1 U235 ( .A(n265), .B(n460), .Y(n134) );
  NOR2X1 U237 ( .A(n766), .B(n739), .Y(n264) );
  NAND2X1 U238 ( .A(n766), .B(n739), .Y(n265) );
  XOR2X1 U239 ( .A(n274), .B(n135), .Y(product[33]) );
  OAI21X1 U241 ( .A(n296), .B(n268), .C(n269), .Y(n267) );
  NAND2X1 U242 ( .A(n282), .B(n270), .Y(n268) );
  AOI21X1 U243 ( .A(n283), .B(n270), .C(n271), .Y(n269) );
  NOR2X1 U244 ( .A(n277), .B(n272), .Y(n270) );
  OAI21X1 U245 ( .A(n280), .B(n272), .C(n273), .Y(n271) );
  NAND2X1 U246 ( .A(n273), .B(n461), .Y(n135) );
  NOR2X1 U248 ( .A(n794), .B(n767), .Y(n272) );
  NAND2X1 U249 ( .A(n794), .B(n767), .Y(n273) );
  XOR2X1 U250 ( .A(n281), .B(n136), .Y(product[32]) );
  AOI21X1 U251 ( .A(n275), .B(n295), .C(n276), .Y(n274) );
  NOR2X1 U252 ( .A(n277), .B(n284), .Y(n275) );
  OAI21X1 U253 ( .A(n277), .B(n285), .C(n280), .Y(n276) );
  NAND2X1 U256 ( .A(n280), .B(n462), .Y(n136) );
  NOR2X1 U258 ( .A(n824), .B(n795), .Y(n277) );
  NAND2X1 U259 ( .A(n824), .B(n795), .Y(n280) );
  AOI21X1 U261 ( .A(n282), .B(n295), .C(n283), .Y(n281) );
  NOR2X1 U266 ( .A(n293), .B(n288), .Y(n282) );
  OAI21X1 U267 ( .A(n294), .B(n288), .C(n289), .Y(n283) );
  NOR2X1 U270 ( .A(n852), .B(n825), .Y(n288) );
  NAND2X1 U271 ( .A(n852), .B(n825), .Y(n289) );
  XNOR2X1 U272 ( .A(n295), .B(n138), .Y(product[30]) );
  AOI21X1 U273 ( .A(n464), .B(n295), .C(n292), .Y(n290) );
  NAND2X1 U276 ( .A(n294), .B(n464), .Y(n138) );
  NOR2X1 U278 ( .A(n880), .B(n853), .Y(n293) );
  NAND2X1 U279 ( .A(n880), .B(n853), .Y(n294) );
  XNOR2X1 U280 ( .A(n305), .B(n139), .Y(product[29]) );
  AOI21X1 U282 ( .A(n333), .B(n297), .C(n298), .Y(n296) );
  NOR2X1 U283 ( .A(n315), .B(n299), .Y(n297) );
  OAI21X1 U284 ( .A(n316), .B(n299), .C(n300), .Y(n298) );
  NAND2X1 U285 ( .A(n1887), .B(n1888), .Y(n299) );
  AOI21X1 U286 ( .A(n311), .B(n1888), .C(n302), .Y(n300) );
  NAND2X1 U289 ( .A(n304), .B(n1888), .Y(n139) );
  NAND2X1 U292 ( .A(n906), .B(n881), .Y(n304) );
  XNOR2X1 U293 ( .A(n314), .B(n140), .Y(product[28]) );
  OAI21X1 U294 ( .A(n306), .B(n332), .C(n307), .Y(n305) );
  NAND2X1 U295 ( .A(n1887), .B(n317), .Y(n306) );
  AOI21X1 U296 ( .A(n1887), .B(n318), .C(n311), .Y(n307) );
  NAND2X1 U301 ( .A(n313), .B(n1887), .Y(n140) );
  NAND2X1 U304 ( .A(n932), .B(n907), .Y(n313) );
  XNOR2X1 U305 ( .A(n325), .B(n141), .Y(product[27]) );
  OAI21X1 U306 ( .A(n315), .B(n332), .C(n316), .Y(n314) );
  NAND2X1 U311 ( .A(n468), .B(n1892), .Y(n315) );
  AOI21X1 U312 ( .A(n1804), .B(n1892), .C(n322), .Y(n316) );
  NAND2X1 U315 ( .A(n324), .B(n1892), .Y(n141) );
  NAND2X1 U318 ( .A(n956), .B(n933), .Y(n324) );
  XOR2X1 U319 ( .A(n332), .B(n142), .Y(product[26]) );
  OAI21X1 U320 ( .A(n326), .B(n332), .C(n327), .Y(n325) );
  NAND2X1 U325 ( .A(n327), .B(n468), .Y(n142) );
  NOR2X1 U327 ( .A(n980), .B(n957), .Y(n326) );
  XOR2X1 U329 ( .A(n340), .B(n143), .Y(product[25]) );
  OAI21X1 U331 ( .A(n334), .B(n351), .C(n335), .Y(n333) );
  NAND2X1 U332 ( .A(n1896), .B(n341), .Y(n334) );
  AOI21X1 U333 ( .A(n1896), .B(n342), .C(n337), .Y(n335) );
  NAND2X1 U336 ( .A(n339), .B(n1896), .Y(n143) );
  NAND2X1 U339 ( .A(n1002), .B(n981), .Y(n339) );
  XOR2X1 U340 ( .A(n345), .B(n144), .Y(product[24]) );
  AOI21X1 U341 ( .A(n341), .B(n350), .C(n342), .Y(n340) );
  NOR2X1 U342 ( .A(n348), .B(n343), .Y(n341) );
  OAI21X1 U343 ( .A(n349), .B(n343), .C(n344), .Y(n342) );
  NAND2X1 U344 ( .A(n344), .B(n470), .Y(n144) );
  NOR2X1 U346 ( .A(n1024), .B(n1003), .Y(n343) );
  NAND2X1 U347 ( .A(n1024), .B(n1003), .Y(n344) );
  XNOR2X1 U348 ( .A(n350), .B(n145), .Y(product[23]) );
  AOI21X1 U349 ( .A(n471), .B(n350), .C(n347), .Y(n345) );
  NAND2X1 U352 ( .A(n349), .B(n471), .Y(n145) );
  NOR2X1 U354 ( .A(n1044), .B(n1025), .Y(n348) );
  NAND2X1 U355 ( .A(n1044), .B(n1025), .Y(n349) );
  XNOR2X1 U356 ( .A(n356), .B(n146), .Y(product[22]) );
  AOI21X1 U358 ( .A(n371), .B(n352), .C(n353), .Y(n351) );
  NOR2X1 U359 ( .A(n354), .B(n357), .Y(n352) );
  OAI21X1 U360 ( .A(n354), .B(n358), .C(n355), .Y(n353) );
  NAND2X1 U361 ( .A(n355), .B(n472), .Y(n146) );
  NOR2X1 U363 ( .A(n1064), .B(n1045), .Y(n354) );
  NAND2X1 U364 ( .A(n1064), .B(n1045), .Y(n355) );
  XNOR2X1 U365 ( .A(n363), .B(n147), .Y(product[21]) );
  OAI21X1 U366 ( .A(n357), .B(n370), .C(n358), .Y(n356) );
  NAND2X1 U367 ( .A(n474), .B(n1893), .Y(n357) );
  AOI21X1 U368 ( .A(n367), .B(n1893), .C(n360), .Y(n358) );
  NAND2X1 U371 ( .A(n362), .B(n1847), .Y(n147) );
  NAND2X1 U374 ( .A(n1082), .B(n1065), .Y(n362) );
  XOR2X1 U375 ( .A(n370), .B(n148), .Y(product[20]) );
  OAI21X1 U376 ( .A(n364), .B(n370), .C(n365), .Y(n363) );
  NAND2X1 U381 ( .A(n365), .B(n474), .Y(n148) );
  NOR2X1 U383 ( .A(n1100), .B(n1083), .Y(n364) );
  NAND2X1 U384 ( .A(n1100), .B(n1083), .Y(n365) );
  OAI21X1 U387 ( .A(n372), .B(n384), .C(n373), .Y(n371) );
  NAND2X1 U388 ( .A(n1900), .B(n1899), .Y(n372) );
  AOI21X1 U389 ( .A(n380), .B(n1899), .C(n375), .Y(n373) );
  NAND2X1 U395 ( .A(n1116), .B(n1101), .Y(n377) );
  XNOR2X1 U396 ( .A(n383), .B(n150), .Y(product[18]) );
  AOI21X1 U397 ( .A(n1900), .B(n383), .C(n380), .Y(n378) );
  NAND2X1 U400 ( .A(n382), .B(n1900), .Y(n150) );
  NAND2X1 U403 ( .A(n1132), .B(n1117), .Y(n382) );
  XNOR2X1 U404 ( .A(n389), .B(n151), .Y(product[17]) );
  AOI21X1 U406 ( .A(n385), .B(n393), .C(n386), .Y(n384) );
  NOR2X1 U407 ( .A(n390), .B(n387), .Y(n385) );
  OAI21X1 U408 ( .A(n391), .B(n387), .C(n388), .Y(n386) );
  NAND2X1 U409 ( .A(n388), .B(n477), .Y(n151) );
  NOR2X1 U411 ( .A(n1146), .B(n1133), .Y(n387) );
  NAND2X1 U412 ( .A(n1146), .B(n1133), .Y(n388) );
  XOR2X1 U413 ( .A(n392), .B(n152), .Y(product[16]) );
  OAI21X1 U414 ( .A(n390), .B(n392), .C(n391), .Y(n389) );
  NAND2X1 U415 ( .A(n391), .B(n478), .Y(n152) );
  NOR2X1 U417 ( .A(n1160), .B(n1147), .Y(n390) );
  NAND2X1 U418 ( .A(n1160), .B(n1147), .Y(n391) );
  OAI21X1 U420 ( .A(n404), .B(n394), .C(n395), .Y(n393) );
  NAND2X1 U421 ( .A(n1906), .B(n1901), .Y(n394) );
  AOI21X1 U422 ( .A(n1903), .B(n1901), .C(n1905), .Y(n395) );
  AOI21X1 U431 ( .A(n411), .B(n405), .C(n406), .Y(n404) );
  NOR2X1 U432 ( .A(n409), .B(n407), .Y(n405) );
  OAI21X1 U433 ( .A(n410), .B(n407), .C(n408), .Y(n406) );
  NOR2X1 U434 ( .A(n1194), .B(n1185), .Y(n407) );
  NAND2X1 U435 ( .A(n1194), .B(n1185), .Y(n408) );
  NOR2X1 U436 ( .A(n1204), .B(n1195), .Y(n409) );
  NAND2X1 U437 ( .A(n1204), .B(n1195), .Y(n410) );
  OAI21X1 U438 ( .A(n412), .B(n414), .C(n413), .Y(n411) );
  NOR2X1 U439 ( .A(n1212), .B(n1205), .Y(n412) );
  NAND2X1 U440 ( .A(n1212), .B(n1205), .Y(n413) );
  AOI21X1 U441 ( .A(n1902), .B(n419), .C(n1904), .Y(n414) );
  OAI21X1 U446 ( .A(n420), .B(n422), .C(n421), .Y(n419) );
  NOR2X1 U447 ( .A(n1226), .B(n1221), .Y(n420) );
  NAND2X1 U448 ( .A(n1226), .B(n1221), .Y(n421) );
  AOI21X1 U449 ( .A(n427), .B(n1898), .C(n1897), .Y(n422) );
  OAI21X1 U454 ( .A(n428), .B(n430), .C(n429), .Y(n427) );
  NOR2X1 U455 ( .A(n1236), .B(n1233), .Y(n428) );
  NAND2X1 U456 ( .A(n1236), .B(n1233), .Y(n429) );
  AOI21X1 U457 ( .A(n435), .B(n1909), .C(n1910), .Y(n430) );
  OAI21X1 U462 ( .A(n436), .B(n438), .C(n437), .Y(n435) );
  NOR2X1 U463 ( .A(n1242), .B(n1241), .Y(n436) );
  NAND2X1 U464 ( .A(n1242), .B(n1241), .Y(n437) );
  AOI21X1 U465 ( .A(n1911), .B(n1907), .C(n1908), .Y(n438) );
  NAND2X1 U473 ( .A(n1675), .B(a[1]), .Y(n446) );
  FAX1 U474 ( .A(n491), .B(n504), .C(n489), .YC(n486), .YS(n487) );
  FAX1 U475 ( .A(n508), .B(n493), .C(n506), .YC(n488), .YS(n489) );
  FAX1 U476 ( .A(n497), .B(n510), .C(n495), .YC(n490), .YS(n491) );
  FAX1 U477 ( .A(n512), .B(n501), .C(n499), .YC(n492), .YS(n493) );
  FAX1 U478 ( .A(n1335), .B(n516), .C(n514), .YC(n494), .YS(n495) );
  FAX1 U479 ( .A(a[23]), .B(n1278), .C(n1315), .YC(n496), .YS(n497) );
  FAX1 U480 ( .A(n1400), .B(n1261), .C(n1296), .YC(n498), .YS(n499) );
  FAX1 U481 ( .A(n1245), .B(n1378), .C(n1356), .YC(n500), .YS(n501) );
  FAX1 U482 ( .A(n507), .B(n520), .C(n505), .YC(n502), .YS(n503) );
  FAX1 U483 ( .A(n509), .B(n524), .C(n522), .YC(n504), .YS(n505) );
  FAX1 U484 ( .A(n528), .B(n526), .C(n511), .YC(n506), .YS(n507) );
  FAX1 U485 ( .A(n517), .B(n515), .C(n513), .YC(n508), .YS(n509) );
  FAX1 U486 ( .A(n534), .B(n532), .C(n530), .YC(n510), .YS(n511) );
  FAX1 U487 ( .A(n1279), .B(n1336), .C(n1316), .YC(n512), .YS(n513) );
  FAX1 U488 ( .A(n1401), .B(n1262), .C(n1297), .YC(n514), .YS(n515) );
  FAX1 U489 ( .A(n1246), .B(n1379), .C(n1357), .YC(n516), .YS(n517) );
  FAX1 U490 ( .A(n523), .B(n538), .C(n521), .YC(n518), .YS(n519) );
  FAX1 U491 ( .A(n542), .B(n525), .C(n540), .YC(n520), .YS(n521) );
  FAX1 U492 ( .A(n544), .B(n529), .C(n527), .YC(n522), .YS(n523) );
  FAX1 U493 ( .A(n533), .B(n531), .C(n546), .YC(n524), .YS(n525) );
  FAX1 U494 ( .A(n550), .B(n548), .C(n535), .YC(n526), .YS(n527) );
  FAX1 U495 ( .A(n1280), .B(n1337), .C(n552), .YC(n528), .YS(n529) );
  FAX1 U496 ( .A(n1263), .B(a[22]), .C(n1317), .YC(n530), .YS(n531) );
  FAX1 U497 ( .A(n1423), .B(n1402), .C(n1298), .YC(n532), .YS(n533) );
  FAX1 U498 ( .A(n1247), .B(n1380), .C(n1358), .YC(n534), .YS(n535) );
  FAX1 U499 ( .A(n541), .B(n556), .C(n539), .YC(n536), .YS(n537) );
  FAX1 U500 ( .A(n560), .B(n543), .C(n558), .YC(n538), .YS(n539) );
  FAX1 U501 ( .A(n547), .B(n562), .C(n545), .YC(n540), .YS(n541) );
  FAX1 U502 ( .A(n551), .B(n549), .C(n564), .YC(n542), .YS(n543) );
  FAX1 U503 ( .A(n568), .B(n566), .C(n553), .YC(n544), .YS(n545) );
  FAX1 U504 ( .A(n1338), .B(n572), .C(n570), .YC(n546), .YS(n547) );
  FAX1 U505 ( .A(n1264), .B(n1281), .C(n1318), .YC(n548), .YS(n549) );
  FAX1 U506 ( .A(n1424), .B(n1403), .C(n1299), .YC(n550), .YS(n551) );
  FAX1 U507 ( .A(n1248), .B(n1381), .C(n1359), .YC(n552), .YS(n553) );
  FAX1 U508 ( .A(n559), .B(n576), .C(n557), .YC(n554), .YS(n555) );
  FAX1 U509 ( .A(n580), .B(n561), .C(n578), .YC(n556), .YS(n557) );
  FAX1 U510 ( .A(n582), .B(n565), .C(n563), .YC(n558), .YS(n559) );
  FAX1 U511 ( .A(n569), .B(n586), .C(n584), .YC(n560), .YS(n561) );
  FAX1 U512 ( .A(n573), .B(n571), .C(n567), .YC(n562), .YS(n563) );
  FAX1 U513 ( .A(n592), .B(n590), .C(n588), .YC(n564), .YS(n565) );
  FAX1 U514 ( .A(a[21]), .B(n1300), .C(n1339), .YC(n566), .YS(n567) );
  FAX1 U515 ( .A(n1445), .B(n1265), .C(n1319), .YC(n568), .YS(n569) );
  FAX1 U516 ( .A(n1425), .B(n1404), .C(n1282), .YC(n570), .YS(n571) );
  FAX1 U517 ( .A(n1249), .B(n1360), .C(n1382), .YC(n572), .YS(n573) );
  FAX1 U518 ( .A(n579), .B(n596), .C(n577), .YC(n574), .YS(n575) );
  FAX1 U519 ( .A(n600), .B(n581), .C(n598), .YC(n576), .YS(n577) );
  FAX1 U520 ( .A(n602), .B(n585), .C(n583), .YC(n578), .YS(n579) );
  FAX1 U521 ( .A(n606), .B(n587), .C(n604), .YC(n580), .YS(n581) );
  FAX1 U522 ( .A(n593), .B(n591), .C(n589), .YC(n582), .YS(n583) );
  FAX1 U523 ( .A(n612), .B(n610), .C(n608), .YC(n584), .YS(n585) );
  FAX1 U524 ( .A(n1301), .B(n1340), .C(n614), .YC(n586), .YS(n587) );
  FAX1 U525 ( .A(n1446), .B(n1266), .C(n1320), .YC(n588), .YS(n589) );
  FAX1 U526 ( .A(n1426), .B(n1405), .C(n1283), .YC(n590), .YS(n591) );
  FAX1 U527 ( .A(n1250), .B(n1383), .C(n1361), .YC(n592), .YS(n593) );
  FAX1 U528 ( .A(n620), .B(n597), .C(n618), .YC(n594), .YS(n595) );
  FAX1 U529 ( .A(n622), .B(n601), .C(n599), .YC(n596), .YS(n597) );
  FAX1 U530 ( .A(n605), .B(n603), .C(n624), .YC(n598), .YS(n599) );
  FAX1 U531 ( .A(n628), .B(n626), .C(n607), .YC(n600), .YS(n601) );
  FAX1 U532 ( .A(n613), .B(n611), .C(n609), .YC(n602), .YS(n603) );
  FAX1 U533 ( .A(n632), .B(n630), .C(n615), .YC(n604), .YS(n605) );
  FAX1 U534 ( .A(n1302), .B(n636), .C(n634), .YC(n606), .YS(n607) );
  FAX1 U535 ( .A(n1267), .B(a[20]), .C(n1321), .YC(n608), .YS(n609) );
  FAX1 U536 ( .A(n1466), .B(n1447), .C(n1341), .YC(n610), .YS(n611) );
  FAX1 U537 ( .A(n1406), .B(n1427), .C(n1284), .YC(n612), .YS(n613) );
  FAX1 U538 ( .A(n1251), .B(n1384), .C(n1362), .YC(n614), .YS(n615) );
  FAX1 U539 ( .A(n621), .B(n640), .C(n619), .YC(n616), .YS(n617) );
  FAX1 U540 ( .A(n644), .B(n623), .C(n642), .YC(n618), .YS(n619) );
  FAX1 U541 ( .A(n627), .B(n625), .C(n646), .YC(n620), .YS(n621) );
  FAX1 U542 ( .A(n650), .B(n648), .C(n629), .YC(n622), .YS(n623) );
  FAX1 U543 ( .A(n633), .B(n631), .C(n652), .YC(n624), .YS(n625) );
  FAX1 U544 ( .A(n656), .B(n637), .C(n635), .YC(n626), .YS(n627) );
  FAX1 U545 ( .A(n660), .B(n658), .C(n654), .YC(n628), .YS(n629) );
  FAX1 U546 ( .A(n1268), .B(n1303), .C(n1342), .YC(n630), .YS(n631) );
  FAX1 U547 ( .A(n1467), .B(n1448), .C(n1322), .YC(n632), .YS(n633) );
  FAX1 U548 ( .A(n1428), .B(n1407), .C(n1285), .YC(n634), .YS(n635) );
  FAX1 U549 ( .A(n1252), .B(n1385), .C(n1363), .YC(n636), .YS(n637) );
  FAX1 U550 ( .A(n643), .B(n664), .C(n641), .YC(n638), .YS(n639) );
  FAX1 U551 ( .A(n668), .B(n645), .C(n666), .YC(n640), .YS(n641) );
  FAX1 U552 ( .A(n649), .B(n670), .C(n647), .YC(n642), .YS(n643) );
  FAX1 U553 ( .A(n653), .B(n672), .C(n651), .YC(n644), .YS(n645) );
  FAX1 U554 ( .A(n657), .B(n676), .C(n674), .YC(n646), .YS(n647) );
  FAX1 U555 ( .A(n661), .B(n659), .C(n655), .YC(n648), .YS(n649) );
  FAX1 U556 ( .A(n682), .B(n680), .C(n678), .YC(n650), .YS(n651) );
  FAX1 U557 ( .A(a[19]), .B(n1343), .C(n684), .YC(n652), .YS(n653) );
  FAX1 U558 ( .A(n1468), .B(n1269), .C(n1323), .YC(n654), .YS(n655) );
  FAX1 U559 ( .A(n1449), .B(n1486), .C(n1286), .YC(n656), .YS(n657) );
  FAX1 U560 ( .A(n1408), .B(n1429), .C(n1304), .YC(n658), .YS(n659) );
  FAX1 U561 ( .A(n1253), .B(n1386), .C(n1364), .YC(n660), .YS(n661) );
  FAX1 U562 ( .A(n667), .B(n688), .C(n665), .YC(n662), .YS(n663) );
  FAX1 U563 ( .A(n692), .B(n669), .C(n690), .YC(n664), .YS(n665) );
  FAX1 U564 ( .A(n673), .B(n694), .C(n671), .YC(n666), .YS(n667) );
  FAX1 U565 ( .A(n698), .B(n696), .C(n675), .YC(n668), .YS(n669) );
  FAX1 U566 ( .A(n681), .B(n700), .C(n677), .YC(n670), .YS(n671) );
  FAX1 U567 ( .A(n685), .B(n683), .C(n679), .YC(n672), .YS(n673) );
  FAX1 U568 ( .A(n706), .B(n704), .C(n702), .YC(n674), .YS(n675) );
  FAX1 U569 ( .A(n1344), .B(n710), .C(n708), .YC(n676), .YS(n677) );
  FAX1 U570 ( .A(n1487), .B(n1270), .C(n1324), .YC(n678), .YS(n679) );
  FAX1 U571 ( .A(n1450), .B(n1469), .C(n1287), .YC(n680), .YS(n681) );
  FAX1 U572 ( .A(n1409), .B(n1430), .C(n1305), .YC(n682), .YS(n683) );
  FAX1 U573 ( .A(n1254), .B(n1387), .C(n1365), .YC(n684), .YS(n685) );
  FAX1 U574 ( .A(n691), .B(n714), .C(n689), .YC(n686), .YS(n687) );
  FAX1 U575 ( .A(n718), .B(n693), .C(n716), .YC(n688), .YS(n689) );
  FAX1 U576 ( .A(n722), .B(n720), .C(n695), .YC(n690), .YS(n691) );
  FAX1 U577 ( .A(n701), .B(n699), .C(n697), .YC(n692), .YS(n693) );
  FAX1 U578 ( .A(n728), .B(n726), .C(n724), .YC(n694), .YS(n695) );
  FAX1 U579 ( .A(n707), .B(n705), .C(n703), .YC(n696), .YS(n697) );
  FAX1 U580 ( .A(n732), .B(n711), .C(n709), .YC(n698), .YS(n699) );
  FAX1 U581 ( .A(n736), .B(n734), .C(n730), .YC(n700), .YS(n701) );
  FAX1 U582 ( .A(n1505), .B(n1345), .C(n1325), .YC(n702), .YS(n703) );
  FAX1 U583 ( .A(n1470), .B(n1271), .C(a[18]), .YC(n704), .YS(n705) );
  FAX1 U584 ( .A(n1488), .B(n1451), .C(n1288), .YC(n706), .YS(n707) );
  FAX1 U585 ( .A(n1431), .B(n1410), .C(n1306), .YC(n708), .YS(n709) );
  FAX1 U586 ( .A(n1255), .B(n1388), .C(n1366), .YC(n710), .YS(n711) );
  FAX1 U587 ( .A(n717), .B(n740), .C(n715), .YC(n712), .YS(n713) );
  FAX1 U589 ( .A(n723), .B(n746), .C(n721), .YC(n716), .YS(n717) );
  FAX1 U591 ( .A(n752), .B(n729), .C(n750), .YC(n720), .YS(n721) );
  FAX1 U592 ( .A(n733), .B(n731), .C(n754), .YC(n722), .YS(n723) );
  FAX1 U593 ( .A(n758), .B(n737), .C(n735), .YC(n724), .YS(n725) );
  FAX1 U594 ( .A(n762), .B(n760), .C(n756), .YC(n726), .YS(n727) );
  FAX1 U595 ( .A(n1346), .B(n1326), .C(n764), .YC(n728), .YS(n729) );
  FAX1 U596 ( .A(n1452), .B(n1506), .C(n1272), .YC(n730), .YS(n731) );
  FAX1 U597 ( .A(n1471), .B(n1489), .C(n1289), .YC(n732), .YS(n733) );
  FAX1 U598 ( .A(n1411), .B(n1432), .C(n1307), .YC(n734), .YS(n735) );
  FAX1 U599 ( .A(n1256), .B(n1389), .C(n1367), .YC(n736), .YS(n737) );
  FAX1 U600 ( .A(n743), .B(n768), .C(n741), .YC(n738), .YS(n739) );
  FAX1 U601 ( .A(n747), .B(n745), .C(n770), .YC(n740), .YS(n741) );
  FAX1 U602 ( .A(n749), .B(n774), .C(n772), .YC(n742), .YS(n743) );
  FAX1 U603 ( .A(n753), .B(n751), .C(n776), .YC(n744), .YS(n745) );
  FAX1 U604 ( .A(n780), .B(n755), .C(n778), .YC(n746), .YS(n747) );
  FAX1 U606 ( .A(n765), .B(n763), .C(n757), .YC(n750), .YS(n751) );
  FAX1 U607 ( .A(n788), .B(n786), .C(n784), .YC(n752), .YS(n753) );
  FAX1 U608 ( .A(n1327), .B(n792), .C(n790), .YC(n754), .YS(n755) );
  FAX1 U609 ( .A(n1507), .B(n1273), .C(n1347), .YC(n756), .YS(n757) );
  FAX1 U610 ( .A(n1472), .B(n1523), .C(a[17]), .YC(n758), .YS(n759) );
  FAX1 U611 ( .A(n1453), .B(n1490), .C(n1290), .YC(n760), .YS(n761) );
  FAX1 U612 ( .A(n1433), .B(n1412), .C(n1308), .YC(n762), .YS(n763) );
  FAX1 U613 ( .A(n1257), .B(n1390), .C(n1368), .YC(n764), .YS(n765) );
  FAX1 U616 ( .A(n777), .B(n802), .C(n800), .YC(n770), .YS(n771) );
  FAX1 U617 ( .A(n781), .B(n804), .C(n779), .YC(n772), .YS(n773) );
  FAX1 U618 ( .A(n808), .B(n783), .C(n806), .YC(n774), .YS(n775) );
  FAX1 U619 ( .A(n789), .B(n785), .C(n810), .YC(n776), .YS(n777) );
  FAX1 U620 ( .A(n793), .B(n791), .C(n787), .YC(n778), .YS(n779) );
  FAX1 U621 ( .A(n816), .B(n814), .C(n812), .YC(n780), .YS(n781) );
  FAX1 U622 ( .A(n822), .B(n820), .C(n818), .YC(n782), .YS(n783) );
  FAX1 U623 ( .A(n1508), .B(n1348), .C(n1328), .YC(n784), .YS(n785) );
  FAX1 U624 ( .A(n1473), .B(n1524), .C(n1274), .YC(n786), .YS(n787) );
  FAX1 U625 ( .A(n1491), .B(n1454), .C(n1291), .YC(n788), .YS(n789) );
  FAX1 U626 ( .A(n1413), .B(n1434), .C(n1309), .YC(n790), .YS(n791) );
  FAX1 U627 ( .A(n1258), .B(n1391), .C(n1369), .YC(n792), .YS(n793) );
  FAX1 U628 ( .A(n799), .B(n826), .C(n797), .YC(n794), .YS(n795) );
  FAX1 U629 ( .A(n803), .B(n801), .C(n828), .YC(n796), .YS(n797) );
  FAX1 U630 ( .A(n805), .B(n832), .C(n830), .YC(n798), .YS(n799) );
  FAX1 U631 ( .A(n834), .B(n809), .C(n807), .YC(n800), .YS(n801) );
  FAX1 U632 ( .A(n838), .B(n811), .C(n836), .YC(n802), .YS(n803) );
  FAX1 U633 ( .A(n817), .B(n813), .C(n840), .YC(n804), .YS(n805) );
  FAX1 U634 ( .A(n819), .B(n821), .C(n815), .YC(n806), .YS(n807) );
  FAX1 U635 ( .A(n842), .B(n846), .C(n844), .YC(n808), .YS(n809) );
  FAX1 U636 ( .A(n823), .B(n850), .C(n848), .YC(n810), .YS(n811) );
  FAX1 U637 ( .A(n1509), .B(n1349), .C(n1329), .YC(n812), .YS(n813) );
  FAX1 U638 ( .A(n1474), .B(n1525), .C(n1275), .YC(n814), .YS(n815) );
  FAX1 U639 ( .A(n1492), .B(n1455), .C(n1292), .YC(n816), .YS(n817) );
  FAX1 U641 ( .A(a[16]), .B(n1392), .C(n1370), .YC(n820), .YS(n821) );
  HAX1 U642 ( .A(n1259), .B(n1540), .YC(n822), .YS(n823) );
  FAX1 U643 ( .A(n829), .B(n854), .C(n827), .YC(n824), .YS(n825) );
  FAX1 U644 ( .A(n833), .B(n831), .C(n856), .YC(n826), .YS(n827) );
  FAX1 U645 ( .A(n835), .B(n860), .C(n858), .YC(n828), .YS(n829) );
  FAX1 U646 ( .A(n839), .B(n862), .C(n837), .YC(n830), .YS(n831) );
  FAX1 U647 ( .A(n841), .B(n866), .C(n864), .YC(n832), .YS(n833) );
  FAX1 U648 ( .A(n847), .B(n845), .C(n843), .YC(n834), .YS(n835) );
  FAX1 U649 ( .A(n872), .B(n868), .C(n849), .YC(n836), .YS(n837) );
  FAX1 U650 ( .A(n876), .B(n874), .C(n870), .YC(n838), .YS(n839) );
  FAX1 U651 ( .A(n1330), .B(n878), .C(n851), .YC(n840), .YS(n841) );
  FAX1 U652 ( .A(n1526), .B(n1510), .C(n1350), .YC(n842), .YS(n843) );
  FAX1 U653 ( .A(n1456), .B(n1475), .C(n1276), .YC(n844), .YS(n845) );
  FAX1 U654 ( .A(n1436), .B(n1493), .C(n1311), .YC(n846), .YS(n847) );
  FAX1 U655 ( .A(n1371), .B(n1415), .C(n1293), .YC(n848), .YS(n849) );
  HAX1 U656 ( .A(n1541), .B(n1393), .YC(n850), .YS(n851) );
  FAX1 U657 ( .A(n857), .B(n882), .C(n855), .YC(n852), .YS(n853) );
  FAX1 U658 ( .A(n886), .B(n859), .C(n884), .YC(n854), .YS(n855) );
  FAX1 U659 ( .A(n863), .B(n888), .C(n861), .YC(n856), .YS(n857) );
  FAX1 U660 ( .A(n867), .B(n890), .C(n865), .YC(n858), .YS(n859) );
  FAX1 U661 ( .A(n869), .B(n894), .C(n892), .YC(n860), .YS(n861) );
  FAX1 U663 ( .A(n898), .B(n896), .C(n877), .YC(n864), .YS(n865) );
  FAX1 U664 ( .A(n879), .B(n902), .C(n900), .YC(n866), .YS(n867) );
  FAX1 U665 ( .A(n1351), .B(n1331), .C(n904), .YC(n868), .YS(n869) );
  FAX1 U666 ( .A(n1476), .B(n1527), .C(n1511), .YC(n870), .YS(n871) );
  FAX1 U667 ( .A(n1494), .B(n1457), .C(n1294), .YC(n872), .YS(n873) );
  FAX1 U668 ( .A(n1416), .B(n1437), .C(n1312), .YC(n874), .YS(n875) );
  FAX1 U669 ( .A(a[15]), .B(n1394), .C(n1372), .YC(n876), .YS(n877) );
  HAX1 U670 ( .A(n1542), .B(n1556), .YC(n878), .YS(n879) );
  FAX1 U671 ( .A(n885), .B(n908), .C(n883), .YC(n880), .YS(n881) );
  FAX1 U672 ( .A(n912), .B(n887), .C(n910), .YC(n882), .YS(n883) );
  FAX1 U673 ( .A(n914), .B(n891), .C(n889), .YC(n884), .YS(n885) );
  FAX1 U674 ( .A(n918), .B(n916), .C(n893), .YC(n886), .YS(n887) );
  FAX1 U675 ( .A(n899), .B(n897), .C(n895), .YC(n888), .YS(n889) );
  FAX1 U676 ( .A(n903), .B(n901), .C(n920), .YC(n890), .YS(n891) );
  FAX1 U677 ( .A(n924), .B(n926), .C(n922), .YC(n892), .YS(n893) );
  FAX1 U678 ( .A(n930), .B(n905), .C(n928), .YC(n894), .YS(n895) );
  FAX1 U679 ( .A(n1458), .B(n1352), .C(n1332), .YC(n896), .YS(n897) );
  FAX1 U681 ( .A(n1438), .B(n1417), .C(n1528), .YC(n900), .YS(n901) );
  FAX1 U682 ( .A(n1395), .B(n1373), .C(n1313), .YC(n902), .YS(n903) );
  HAX1 U683 ( .A(n1543), .B(n1557), .YC(n904), .YS(n905) );
  FAX1 U686 ( .A(n940), .B(n917), .C(n915), .YC(n910), .YS(n911) );
  FAX1 U687 ( .A(n944), .B(n942), .C(n919), .YC(n912), .YS(n913) );
  FAX1 U688 ( .A(n925), .B(n923), .C(n921), .YC(n914), .YS(n915) );
  FAX1 U689 ( .A(n946), .B(n948), .C(n927), .YC(n916), .YS(n917) );
  FAX1 U690 ( .A(n952), .B(n950), .C(n929), .YC(n918), .YS(n919) );
  FAX1 U691 ( .A(n1333), .B(n954), .C(n931), .YC(n920), .YS(n921) );
  FAX1 U692 ( .A(n1496), .B(n1459), .C(n1353), .YC(n922), .YS(n923) );
  FAX1 U693 ( .A(n1418), .B(n1478), .C(n1513), .YC(n924), .YS(n925) );
  FAX1 U694 ( .A(n1374), .B(n1439), .C(n1529), .YC(n926), .YS(n927) );
  FAX1 U695 ( .A(n1558), .B(a[14]), .C(n1396), .YC(n928), .YS(n929) );
  HAX1 U696 ( .A(n1544), .B(n1571), .YC(n930), .YS(n931) );
  FAX1 U699 ( .A(n964), .B(n943), .C(n941), .YC(n936), .YS(n937) );
  FAX1 U700 ( .A(n968), .B(n966), .C(n945), .YC(n938), .YS(n939) );
  FAX1 U701 ( .A(n951), .B(n949), .C(n947), .YC(n940), .YS(n941) );
  FAX1 U702 ( .A(n972), .B(n970), .C(n953), .YC(n942), .YS(n943) );
  FAX1 U703 ( .A(n955), .B(n976), .C(n974), .YC(n944), .YS(n945) );
  FAX1 U705 ( .A(n1514), .B(n1497), .C(n1479), .YC(n948), .YS(n949) );
  FAX1 U706 ( .A(n1440), .B(n1419), .C(n1530), .YC(n950), .YS(n951) );
  FAX1 U707 ( .A(n1572), .B(n1397), .C(n1375), .YC(n952), .YS(n953) );
  HAX1 U708 ( .A(n1545), .B(n1559), .YC(n954), .YS(n955) );
  FAX1 U710 ( .A(n986), .B(n963), .C(n984), .YC(n958), .YS(n959) );
  FAX1 U711 ( .A(n988), .B(n967), .C(n965), .YC(n960), .YS(n961) );
  FAX1 U712 ( .A(n971), .B(n969), .C(n990), .YC(n962), .YS(n963) );
  FAX1 U713 ( .A(n975), .B(n973), .C(n992), .YC(n964), .YS(n965) );
  FAX1 U715 ( .A(n1000), .B(n979), .C(n998), .YC(n968), .YS(n969) );
  FAX1 U716 ( .A(n1498), .B(n1461), .C(n1480), .YC(n970), .YS(n971) );
  FAX1 U717 ( .A(n1420), .B(n1441), .C(n1531), .YC(n972), .YS(n973) );
  FAX1 U718 ( .A(n1398), .B(n1376), .C(n1515), .YC(n974), .YS(n975) );
  FAX1 U719 ( .A(n1560), .B(n1573), .C(a[13]), .YC(n976), .YS(n977) );
  FAX1 U721 ( .A(n985), .B(n1004), .C(n983), .YC(n980), .YS(n981) );
  FAX1 U722 ( .A(n1008), .B(n987), .C(n1006), .YC(n982), .YS(n983) );
  FAX1 U723 ( .A(n1010), .B(n991), .C(n989), .YC(n984), .YS(n985) );
  FAX1 U724 ( .A(n995), .B(n993), .C(n1012), .YC(n986), .YS(n987) );
  FAX1 U725 ( .A(n999), .B(n1014), .C(n997), .YC(n988), .YS(n989) );
  FAX1 U726 ( .A(n1020), .B(n1018), .C(n1016), .YC(n990), .YS(n991) );
  FAX1 U727 ( .A(n1499), .B(n1022), .C(n1001), .YC(n992), .YS(n993) );
  FAX1 U728 ( .A(n1516), .B(n1462), .C(n1481), .YC(n994), .YS(n995) );
  FAX1 U729 ( .A(n1442), .B(n1421), .C(n1532), .YC(n996), .YS(n997) );
  FAX1 U730 ( .A(n1586), .B(n1574), .C(n1399), .YC(n998), .YS(n999) );
  HAX1 U731 ( .A(n1547), .B(n1561), .YC(n1000), .YS(n1001) );
  FAX1 U732 ( .A(n1007), .B(n1026), .C(n1005), .YC(n1002), .YS(n1003) );
  FAX1 U734 ( .A(n1032), .B(n1013), .C(n1030), .YC(n1006), .YS(n1007) );
  FAX1 U735 ( .A(n1017), .B(n1015), .C(n1034), .YC(n1008), .YS(n1009) );
  FAX1 U736 ( .A(n1038), .B(n1036), .C(n1019), .YC(n1010), .YS(n1011) );
  FAX1 U737 ( .A(n1023), .B(n1040), .C(n1021), .YC(n1012), .YS(n1013) );
  FAX1 U739 ( .A(n1500), .B(n1463), .C(n1517), .YC(n1016), .YS(n1017) );
  FAX1 U740 ( .A(n1575), .B(n1443), .C(n1422), .YC(n1018), .YS(n1019) );
  FAX1 U741 ( .A(n1562), .B(n1587), .C(a[12]), .YC(n1020), .YS(n1021) );
  HAX1 U742 ( .A(n1548), .B(n1598), .YC(n1022), .YS(n1023) );
  FAX1 U743 ( .A(n1029), .B(n1046), .C(n1027), .YC(n1024), .YS(n1025) );
  FAX1 U744 ( .A(n1033), .B(n1031), .C(n1048), .YC(n1026), .YS(n1027) );
  FAX1 U746 ( .A(n1039), .B(n1037), .C(n1054), .YC(n1030), .YS(n1031) );
  FAX1 U747 ( .A(n1058), .B(n1041), .C(n1056), .YC(n1032), .YS(n1033) );
  FAX1 U748 ( .A(n1062), .B(n1043), .C(n1060), .YC(n1034), .YS(n1035) );
  FAX1 U749 ( .A(n1501), .B(n1483), .C(n1534), .YC(n1036), .YS(n1037) );
  FAX1 U750 ( .A(n1444), .B(n1464), .C(n1518), .YC(n1038), .YS(n1039) );
  FAX1 U751 ( .A(n1563), .B(n1576), .C(n1599), .YC(n1040), .YS(n1041) );
  HAX1 U752 ( .A(n1549), .B(n1588), .YC(n1042), .YS(n1043) );
  FAX1 U753 ( .A(n1049), .B(n1066), .C(n1047), .YC(n1044), .YS(n1045) );
  FAX1 U754 ( .A(n1053), .B(n1051), .C(n1068), .YC(n1046), .YS(n1047) );
  FAX1 U755 ( .A(n1055), .B(n1072), .C(n1070), .YC(n1048), .YS(n1049) );
  FAX1 U756 ( .A(n1059), .B(n1074), .C(n1057), .YC(n1050), .YS(n1051) );
  FAX1 U757 ( .A(n1078), .B(n1061), .C(n1076), .YC(n1052), .YS(n1053) );
  FAX1 U758 ( .A(n1535), .B(n1080), .C(n1063), .YC(n1054), .YS(n1055) );
  FAX1 U759 ( .A(n1502), .B(n1484), .C(n1519), .YC(n1056), .YS(n1057) );
  FAX1 U760 ( .A(n1589), .B(n1610), .C(n1465), .YC(n1058), .YS(n1059) );
  FAX1 U761 ( .A(n1564), .B(n1577), .C(a[11]), .YC(n1060), .YS(n1061) );
  HAX1 U762 ( .A(n1550), .B(n1600), .YC(n1062), .YS(n1063) );
  FAX1 U763 ( .A(n1069), .B(n1084), .C(n1067), .YC(n1064), .YS(n1065) );
  FAX1 U764 ( .A(n1073), .B(n1071), .C(n1086), .YC(n1066), .YS(n1067) );
  FAX1 U765 ( .A(n1075), .B(n1090), .C(n1088), .YC(n1068), .YS(n1069) );
  FAX1 U766 ( .A(n1079), .B(n1092), .C(n1077), .YC(n1070), .YS(n1071) );
  FAX1 U767 ( .A(n1081), .B(n1096), .C(n1094), .YC(n1072), .YS(n1073) );
  FAX1 U768 ( .A(n1536), .B(n1520), .C(n1098), .YC(n1074), .YS(n1075) );
  FAX1 U769 ( .A(n1578), .B(n1485), .C(n1503), .YC(n1076), .YS(n1077) );
  FAX1 U770 ( .A(n1601), .B(n1590), .C(n1565), .YC(n1078), .YS(n1079) );
  HAX1 U771 ( .A(n1551), .B(n1611), .YC(n1080), .YS(n1081) );
  FAX1 U772 ( .A(n1087), .B(n1102), .C(n1085), .YC(n1082), .YS(n1083) );
  FAX1 U773 ( .A(n1091), .B(n1089), .C(n1104), .YC(n1084), .YS(n1085) );
  FAX1 U775 ( .A(n1110), .B(n1097), .C(n1095), .YC(n1088), .YS(n1089) );
  FAX1 U776 ( .A(n1114), .B(n1099), .C(n1112), .YC(n1090), .YS(n1091) );
  FAX1 U777 ( .A(n1504), .B(n1537), .C(n1521), .YC(n1092), .YS(n1093) );
  FAX1 U778 ( .A(n1591), .B(n1579), .C(n1566), .YC(n1094), .YS(n1095) );
  FAX1 U779 ( .A(n1612), .B(n1602), .C(a[10]), .YC(n1096), .YS(n1097) );
  HAX1 U780 ( .A(n1552), .B(n1621), .YC(n1098), .YS(n1099) );
  FAX1 U781 ( .A(n1105), .B(n1118), .C(n1103), .YC(n1100), .YS(n1101) );
  FAX1 U782 ( .A(n1122), .B(n1107), .C(n1120), .YC(n1102), .YS(n1103) );
  FAX1 U783 ( .A(n1124), .B(n1111), .C(n1109), .YC(n1104), .YS(n1105) );
  FAX1 U784 ( .A(n1128), .B(n1126), .C(n1113), .YC(n1106), .YS(n1107) );
  FAX1 U785 ( .A(n1522), .B(n1130), .C(n1115), .YC(n1108), .YS(n1109) );
  FAX1 U786 ( .A(n1603), .B(n1580), .C(n1538), .YC(n1110), .YS(n1111) );
  FAX1 U787 ( .A(n1622), .B(n1613), .C(n1592), .YC(n1112), .YS(n1113) );
  HAX1 U788 ( .A(n1553), .B(n1567), .YC(n1114), .YS(n1115) );
  FAX1 U789 ( .A(n1121), .B(n1134), .C(n1119), .YC(n1116), .YS(n1117) );
  FAX1 U790 ( .A(n1138), .B(n1136), .C(n1123), .YC(n1118), .YS(n1119) );
  FAX1 U791 ( .A(n1127), .B(n1129), .C(n1125), .YC(n1120), .YS(n1121) );
  FAX1 U792 ( .A(n1131), .B(n1142), .C(n1140), .YC(n1122), .YS(n1123) );
  FAX1 U793 ( .A(n1593), .B(n1539), .C(n1144), .YC(n1124), .YS(n1125) );
  FAX1 U794 ( .A(n1604), .B(n1623), .C(n1568), .YC(n1126), .YS(n1127) );
  FAX1 U795 ( .A(n1631), .B(n1614), .C(a[9]), .YC(n1128), .YS(n1129) );
  HAX1 U796 ( .A(n1554), .B(n1581), .YC(n1130), .YS(n1131) );
  FAX1 U797 ( .A(n1137), .B(n1148), .C(n1135), .YC(n1132), .YS(n1133) );
  FAX1 U798 ( .A(n1152), .B(n1150), .C(n1139), .YC(n1134), .YS(n1135) );
  FAX1 U799 ( .A(n1154), .B(n1141), .C(n1143), .YC(n1136), .YS(n1137) );
  FAX1 U800 ( .A(n1158), .B(n1145), .C(n1156), .YC(n1138), .YS(n1139) );
  FAX1 U801 ( .A(n1624), .B(n1615), .C(n1594), .YC(n1140), .YS(n1141) );
  FAX1 U802 ( .A(n1605), .B(n1632), .C(n1582), .YC(n1142), .YS(n1143) );
  HAX1 U803 ( .A(n1555), .B(n1569), .YC(n1144), .YS(n1145) );
  FAX1 U804 ( .A(n1151), .B(n1162), .C(n1149), .YC(n1146), .YS(n1147) );
  FAX1 U805 ( .A(n1157), .B(n1153), .C(n1164), .YC(n1148), .YS(n1149) );
  FAX1 U806 ( .A(n1168), .B(n1166), .C(n1155), .YC(n1150), .YS(n1151) );
  FAX1 U807 ( .A(n1595), .B(n1159), .C(n1170), .YC(n1152), .YS(n1153) );
  FAX1 U809 ( .A(n1606), .B(n1616), .C(n1570), .YC(n1156), .YS(n1157) );
  HAX1 U810 ( .A(n1640), .B(a[8]), .YC(n1158), .YS(n1159) );
  FAX1 U811 ( .A(n1174), .B(n1165), .C(n1163), .YC(n1160), .YS(n1161) );
  FAX1 U812 ( .A(n1169), .B(n1167), .C(n1176), .YC(n1162), .YS(n1163) );
  FAX1 U813 ( .A(n1171), .B(n1180), .C(n1178), .YC(n1164), .YS(n1165) );
  FAX1 U814 ( .A(n1607), .B(n1596), .C(n1584), .YC(n1166), .YS(n1167) );
  FAX1 U815 ( .A(n1626), .B(n1617), .C(n1182), .YC(n1168), .YS(n1169) );
  HAX1 U816 ( .A(n1641), .B(n1634), .YC(n1170), .YS(n1171) );
  FAX1 U817 ( .A(n1186), .B(n1177), .C(n1175), .YC(n1172), .YS(n1173) );
  FAX1 U818 ( .A(n1188), .B(n1181), .C(n1179), .YC(n1174), .YS(n1175) );
  FAX1 U819 ( .A(n1192), .B(n1183), .C(n1190), .YC(n1176), .YS(n1177) );
  FAX1 U820 ( .A(n1618), .B(n1627), .C(n1597), .YC(n1178), .YS(n1179) );
  FAX1 U821 ( .A(n1642), .B(n1635), .C(n1608), .YC(n1180), .YS(n1181) );
  HAX1 U822 ( .A(n1648), .B(a[7]), .YC(n1182), .YS(n1183) );
  FAX1 U823 ( .A(n1189), .B(n1196), .C(n1187), .YC(n1184), .YS(n1185) );
  FAX1 U824 ( .A(n1200), .B(n1198), .C(n1191), .YC(n1186), .YS(n1187) );
  FAX1 U825 ( .A(n1628), .B(n1609), .C(n1193), .YC(n1188), .YS(n1189) );
  FAX1 U826 ( .A(n1619), .B(n1636), .C(n1202), .YC(n1190), .YS(n1191) );
  HAX1 U827 ( .A(n1649), .B(n1643), .YC(n1192), .YS(n1193) );
  FAX1 U828 ( .A(n1199), .B(n1206), .C(n1197), .YC(n1194), .YS(n1195) );
  FAX1 U829 ( .A(n1203), .B(n1208), .C(n1201), .YC(n1196), .YS(n1197) );
  FAX1 U830 ( .A(n1637), .B(n1629), .C(n1210), .YC(n1198), .YS(n1199) );
  FAX1 U831 ( .A(n1655), .B(n1644), .C(n1620), .YC(n1200), .YS(n1201) );
  HAX1 U832 ( .A(n1650), .B(a[6]), .YC(n1202), .YS(n1203) );
  FAX1 U833 ( .A(n1214), .B(n1209), .C(n1207), .YC(n1204), .YS(n1205) );
  FAX1 U834 ( .A(n1218), .B(n1211), .C(n1216), .YC(n1206), .YS(n1207) );
  FAX1 U835 ( .A(n1645), .B(n1638), .C(n1630), .YC(n1208), .YS(n1209) );
  HAX1 U836 ( .A(n1656), .B(n1651), .YC(n1210), .YS(n1211) );
  FAX1 U837 ( .A(n1222), .B(n1217), .C(n1215), .YC(n1212), .YS(n1213) );
  FAX1 U838 ( .A(n1639), .B(n1224), .C(n1219), .YC(n1214), .YS(n1215) );
  FAX1 U839 ( .A(n1657), .B(a[5]), .C(n1646), .YC(n1216), .YS(n1217) );
  HAX1 U840 ( .A(n1661), .B(n1652), .YC(n1218), .YS(n1219) );
  FAX1 U841 ( .A(n1225), .B(n1228), .C(n1223), .YC(n1220), .YS(n1221) );
  FAX1 U842 ( .A(n1658), .B(n1647), .C(n1230), .YC(n1222), .YS(n1223) );
  HAX1 U843 ( .A(n1662), .B(n1653), .YC(n1224), .YS(n1225) );
  FAX1 U844 ( .A(n1231), .B(n1234), .C(n1229), .YC(n1226), .YS(n1227) );
  FAX1 U845 ( .A(n1663), .B(n1659), .C(n1654), .YC(n1228), .YS(n1229) );
  HAX1 U846 ( .A(n1666), .B(a[4]), .YC(n1230), .YS(n1231) );
  FAX1 U847 ( .A(n1660), .B(n1238), .C(n1235), .YC(n1232), .YS(n1233) );
  HAX1 U848 ( .A(n1667), .B(n1664), .YC(n1234), .YS(n1235) );
  FAX1 U849 ( .A(a[3]), .B(n1665), .C(n1240), .YC(n1236), .YS(n1237) );
  HAX1 U850 ( .A(n1670), .B(n1668), .YC(n1238), .YS(n1239) );
  HAX1 U851 ( .A(n1671), .B(n1669), .YC(n1240), .YS(n1241) );
  HAX1 U852 ( .A(n1673), .B(a[2]), .YC(n1242), .YS(n1243) );
  NOR2X1 U853 ( .A(n1940), .B(n1784), .Y(n1244) );
  NOR2X1 U854 ( .A(n1940), .B(n1917), .Y(n1245) );
  NOR2X1 U855 ( .A(n1940), .B(n1964), .Y(n1246) );
  NOR2X1 U856 ( .A(n1939), .B(n1914), .Y(n1247) );
  NOR2X1 U857 ( .A(n1939), .B(n1968), .Y(n1248) );
  NOR2X1 U858 ( .A(n1939), .B(n1925), .Y(n1249) );
  NOR2X1 U859 ( .A(n1939), .B(n1970), .Y(n1250) );
  NOR2X1 U860 ( .A(n1939), .B(n1928), .Y(n1251) );
  NOR2X1 U861 ( .A(n1939), .B(n1974), .Y(n1252) );
  NOR2X1 U862 ( .A(n1939), .B(n1930), .Y(n1253) );
  NOR2X1 U863 ( .A(n1939), .B(n1978), .Y(n1254) );
  NOR2X1 U864 ( .A(n1933), .B(n1939), .Y(n1255) );
  NOR2X1 U865 ( .A(n1984), .B(n1939), .Y(n1256) );
  NOR2X1 U866 ( .A(n1936), .B(n1939), .Y(n1257) );
  NOR2X1 U867 ( .A(n1987), .B(n1939), .Y(n1258) );
  NOR2X1 U868 ( .A(n1992), .B(n1939), .Y(n1259) );
  NOR2X1 U869 ( .A(n1923), .B(n80), .Y(n1260) );
  NOR2X1 U870 ( .A(n1961), .B(n80), .Y(n1261) );
  NOR2X1 U871 ( .A(n1918), .B(n80), .Y(n1262) );
  NOR2X1 U872 ( .A(n1964), .B(n80), .Y(n1263) );
  NOR2X1 U873 ( .A(n1915), .B(n80), .Y(n1264) );
  NOR2X1 U874 ( .A(n1968), .B(n80), .Y(n1265) );
  NOR2X1 U875 ( .A(n1926), .B(n80), .Y(n1266) );
  NOR2X1 U876 ( .A(n1972), .B(n80), .Y(n1267) );
  NOR2X1 U877 ( .A(n1928), .B(n80), .Y(n1268) );
  NOR2X1 U878 ( .A(n1975), .B(n80), .Y(n1269) );
  NOR2X1 U879 ( .A(n1930), .B(n80), .Y(n1270) );
  NOR2X1 U880 ( .A(n1978), .B(n80), .Y(n1271) );
  NOR2X1 U881 ( .A(n1933), .B(n80), .Y(n1272) );
  NOR2X1 U882 ( .A(n1984), .B(n80), .Y(n1273) );
  NOR2X1 U883 ( .A(n1936), .B(n80), .Y(n1274) );
  NOR2X1 U884 ( .A(n1987), .B(n80), .Y(n1275) );
  NOR2X1 U885 ( .A(n1992), .B(n80), .Y(n1276) );
  NOR2X1 U886 ( .A(n1956), .B(n1942), .Y(n1277) );
  NOR2X1 U887 ( .A(n1923), .B(n1942), .Y(n1278) );
  NOR2X1 U888 ( .A(n1961), .B(n1941), .Y(n1279) );
  NOR2X1 U889 ( .A(n1917), .B(n1941), .Y(n1280) );
  NOR2X1 U890 ( .A(n1964), .B(n1941), .Y(n1281) );
  NOR2X1 U891 ( .A(n1914), .B(n1941), .Y(n1282) );
  NOR2X1 U892 ( .A(n1969), .B(n1941), .Y(n1283) );
  NOR2X1 U893 ( .A(n1925), .B(n1941), .Y(n1284) );
  NOR2X1 U894 ( .A(n1972), .B(n1941), .Y(n1285) );
  NOR2X1 U895 ( .A(n1928), .B(n1941), .Y(n1286) );
  NOR2X1 U896 ( .A(n1974), .B(n1941), .Y(n1287) );
  NOR2X1 U897 ( .A(n1932), .B(n1941), .Y(n1288) );
  NOR2X1 U898 ( .A(n1978), .B(n1941), .Y(n1289) );
  NOR2X1 U899 ( .A(n1933), .B(n1941), .Y(n1290) );
  NOR2X1 U900 ( .A(n1984), .B(n1942), .Y(n1291) );
  NOR2X1 U901 ( .A(n1936), .B(n1942), .Y(n1292) );
  NOR2X1 U902 ( .A(n1987), .B(n1942), .Y(n1293) );
  NOR2X1 U903 ( .A(n1992), .B(n1942), .Y(n1294) );
  NOR2X1 U904 ( .A(n1938), .B(n76), .Y(n1295) );
  NOR2X1 U905 ( .A(n1956), .B(n76), .Y(n1296) );
  NOR2X1 U906 ( .A(n1923), .B(n76), .Y(n1297) );
  NOR2X1 U907 ( .A(n1961), .B(n76), .Y(n1298) );
  NOR2X1 U908 ( .A(n1918), .B(n76), .Y(n1299) );
  NOR2X1 U909 ( .A(n1964), .B(n76), .Y(n1300) );
  NOR2X1 U910 ( .A(n1915), .B(n76), .Y(n1301) );
  NOR2X1 U911 ( .A(n1969), .B(n76), .Y(n1302) );
  NOR2X1 U912 ( .A(n1925), .B(n76), .Y(n1303) );
  NOR2X1 U913 ( .A(n1972), .B(n76), .Y(n1304) );
  NOR2X1 U914 ( .A(n1928), .B(n76), .Y(n1305) );
  NOR2X1 U915 ( .A(n1975), .B(n76), .Y(n1306) );
  NOR2X1 U916 ( .A(n1932), .B(n76), .Y(n1307) );
  NOR2X1 U917 ( .A(n1979), .B(n76), .Y(n1308) );
  NOR2X1 U918 ( .A(n1933), .B(n76), .Y(n1309) );
  NOR2X1 U919 ( .A(n1984), .B(n76), .Y(n1310) );
  NOR2X1 U920 ( .A(n1936), .B(n76), .Y(n1311) );
  NOR2X1 U923 ( .A(n1953), .B(n1944), .Y(n1314) );
  NOR2X1 U924 ( .A(n1938), .B(n1944), .Y(n1315) );
  NOR2X1 U925 ( .A(n1956), .B(n1944), .Y(n1316) );
  NOR2X1 U926 ( .A(n1923), .B(n1944), .Y(n1317) );
  NOR2X1 U927 ( .A(n1961), .B(n1943), .Y(n1318) );
  NOR2X1 U928 ( .A(n1918), .B(n1943), .Y(n1319) );
  NOR2X1 U929 ( .A(n1964), .B(n1943), .Y(n1320) );
  NOR2X1 U930 ( .A(n1915), .B(n1943), .Y(n1321) );
  NOR2X1 U931 ( .A(n1968), .B(n1943), .Y(n1322) );
  NOR2X1 U932 ( .A(n1925), .B(n1943), .Y(n1323) );
  NOR2X1 U933 ( .A(n1972), .B(n1943), .Y(n1324) );
  NOR2X1 U934 ( .A(n1928), .B(n1943), .Y(n1325) );
  NOR2X1 U935 ( .A(n1974), .B(n1943), .Y(n1326) );
  NOR2X1 U936 ( .A(n1932), .B(n1943), .Y(n1327) );
  NOR2X1 U937 ( .A(n1978), .B(n1943), .Y(n1328) );
  NOR2X1 U938 ( .A(n1933), .B(n1943), .Y(n1329) );
  NOR2X1 U939 ( .A(n1984), .B(n1944), .Y(n1330) );
  NOR2X1 U940 ( .A(n1936), .B(n1944), .Y(n1331) );
  NOR2X1 U941 ( .A(n1987), .B(n1944), .Y(n1332) );
  NOR2X1 U942 ( .A(n1992), .B(n1944), .Y(n1333) );
  NOR2X1 U943 ( .A(n1921), .B(n1882), .Y(n1334) );
  NOR2X1 U944 ( .A(n1952), .B(n1882), .Y(n1335) );
  NOR2X1 U945 ( .A(n1938), .B(n1882), .Y(n1336) );
  NOR2X1 U946 ( .A(n1956), .B(n1882), .Y(n1337) );
  NOR2X1 U947 ( .A(n1923), .B(n1882), .Y(n1338) );
  NOR2X1 U948 ( .A(n1961), .B(n72), .Y(n1339) );
  NOR2X1 U949 ( .A(n1918), .B(n72), .Y(n1340) );
  NOR2X1 U950 ( .A(n1964), .B(n72), .Y(n1341) );
  NOR2X1 U951 ( .A(n1915), .B(n72), .Y(n1342) );
  NOR2X1 U952 ( .A(n1968), .B(n72), .Y(n1343) );
  NOR2X1 U953 ( .A(n1925), .B(n72), .Y(n1344) );
  NOR2X1 U954 ( .A(n1972), .B(n72), .Y(n1345) );
  NOR2X1 U955 ( .A(n1928), .B(n72), .Y(n1346) );
  NOR2X1 U956 ( .A(n1974), .B(n72), .Y(n1347) );
  NOR2X1 U957 ( .A(n1932), .B(n72), .Y(n1348) );
  NOR2X1 U958 ( .A(n1978), .B(n72), .Y(n1349) );
  NOR2X1 U959 ( .A(n1934), .B(n72), .Y(n1350) );
  NOR2X1 U960 ( .A(n1983), .B(n72), .Y(n1351) );
  NOR2X1 U961 ( .A(n1935), .B(n72), .Y(n1352) );
  NOR2X1 U962 ( .A(n1986), .B(n72), .Y(n1353) );
  NOR2X1 U963 ( .A(n1992), .B(n72), .Y(n1354) );
  NOR2X1 U964 ( .A(n1946), .B(n1950), .Y(n1355) );
  NOR2X1 U965 ( .A(n1946), .B(n1921), .Y(n1356) );
  NOR2X1 U966 ( .A(n1946), .B(n1952), .Y(n1357) );
  NOR2X1 U967 ( .A(n1946), .B(n1938), .Y(n1358) );
  NOR2X1 U968 ( .A(n1946), .B(n1956), .Y(n1359) );
  NOR2X1 U969 ( .A(n1923), .B(n1946), .Y(n1360) );
  NOR2X1 U970 ( .A(n1786), .B(n1945), .Y(n1361) );
  NOR2X1 U971 ( .A(n1918), .B(n1945), .Y(n1362) );
  NOR2X1 U972 ( .A(n1964), .B(n1945), .Y(n1363) );
  NOR2X1 U973 ( .A(n1915), .B(n1945), .Y(n1364) );
  NOR2X1 U974 ( .A(n1968), .B(n1945), .Y(n1365) );
  NOR2X1 U975 ( .A(n1926), .B(n1945), .Y(n1366) );
  NOR2X1 U976 ( .A(n1971), .B(n1945), .Y(n1367) );
  NOR2X1 U977 ( .A(n1929), .B(n1945), .Y(n1368) );
  NOR2X1 U978 ( .A(n1974), .B(n1945), .Y(n1369) );
  NOR2X1 U979 ( .A(n1932), .B(n1945), .Y(n1370) );
  NOR2X1 U980 ( .A(n1979), .B(n1945), .Y(n1371) );
  NOR2X1 U981 ( .A(n1934), .B(n1945), .Y(n1372) );
  NOR2X1 U982 ( .A(n1983), .B(n1946), .Y(n1373) );
  NOR2X1 U983 ( .A(n1935), .B(n1946), .Y(n1374) );
  NOR2X1 U984 ( .A(n1986), .B(n1946), .Y(n1375) );
  NOR2X1 U985 ( .A(n1992), .B(n1946), .Y(n1376) );
  NOR2X1 U986 ( .A(n68), .B(n1937), .Y(n1377) );
  NOR2X1 U987 ( .A(n68), .B(n1950), .Y(n1378) );
  NOR2X1 U988 ( .A(n68), .B(n1921), .Y(n1379) );
  NOR2X1 U989 ( .A(n68), .B(n1952), .Y(n1380) );
  NOR2X1 U990 ( .A(n68), .B(n1938), .Y(n1381) );
  NOR2X1 U991 ( .A(n68), .B(n1955), .Y(n1382) );
  NOR2X1 U992 ( .A(n1924), .B(n68), .Y(n1383) );
  NOR2X1 U993 ( .A(n1787), .B(n68), .Y(n1384) );
  NOR2X1 U994 ( .A(n1918), .B(n68), .Y(n1385) );
  NOR2X1 U995 ( .A(n1966), .B(n68), .Y(n1386) );
  NOR2X1 U996 ( .A(n1915), .B(n68), .Y(n1387) );
  NOR2X1 U997 ( .A(n1968), .B(n68), .Y(n1388) );
  NOR2X1 U998 ( .A(n1925), .B(n68), .Y(n1389) );
  NOR2X1 U999 ( .A(n1971), .B(n68), .Y(n1390) );
  NOR2X1 U1000 ( .A(n1928), .B(n68), .Y(n1391) );
  NOR2X1 U1001 ( .A(n1975), .B(n68), .Y(n1392) );
  NOR2X1 U1002 ( .A(n1931), .B(n68), .Y(n1393) );
  NOR2X1 U1003 ( .A(n1978), .B(n68), .Y(n1394) );
  NOR2X1 U1004 ( .A(n1934), .B(n68), .Y(n1395) );
  NOR2X1 U1005 ( .A(n1983), .B(n68), .Y(n1396) );
  NOR2X1 U1006 ( .A(n1935), .B(n68), .Y(n1397) );
  NOR2X1 U1007 ( .A(n1986), .B(n68), .Y(n1398) );
  NOR2X1 U1008 ( .A(n1991), .B(n68), .Y(n1399) );
  NOR2X1 U1009 ( .A(n1948), .B(n1937), .Y(n1400) );
  NOR2X1 U1010 ( .A(n1948), .B(n1950), .Y(n1401) );
  NOR2X1 U1011 ( .A(n1921), .B(n1948), .Y(n1402) );
  NOR2X1 U1012 ( .A(n1948), .B(n1952), .Y(n1403) );
  NOR2X1 U1013 ( .A(n1948), .B(n1938), .Y(n1404) );
  NOR2X1 U1014 ( .A(n1948), .B(n1955), .Y(n1405) );
  NOR2X1 U1015 ( .A(n1923), .B(n1948), .Y(n1406) );
  NOR2X1 U1016 ( .A(n1787), .B(n1947), .Y(n1407) );
  NOR2X1 U1017 ( .A(n1918), .B(n1947), .Y(n1408) );
  NOR2X1 U1018 ( .A(n1964), .B(n1947), .Y(n1409) );
  NOR2X1 U1019 ( .A(n1915), .B(n1947), .Y(n1410) );
  NOR2X1 U1020 ( .A(n1968), .B(n1947), .Y(n1411) );
  NOR2X1 U1021 ( .A(n1926), .B(n1947), .Y(n1412) );
  NOR2X1 U1022 ( .A(n1971), .B(n1947), .Y(n1413) );
  NOR2X1 U1023 ( .A(n1929), .B(n1947), .Y(n1414) );
  NOR2X1 U1024 ( .A(n1975), .B(n1947), .Y(n1415) );
  NOR2X1 U1025 ( .A(n1931), .B(n1947), .Y(n1416) );
  NOR2X1 U1026 ( .A(n1979), .B(n1947), .Y(n1417) );
  NOR2X1 U1027 ( .A(n1934), .B(n1947), .Y(n1418) );
  NOR2X1 U1028 ( .A(n1983), .B(n1948), .Y(n1419) );
  NOR2X1 U1029 ( .A(n1935), .B(n1948), .Y(n1420) );
  NOR2X1 U1030 ( .A(n1986), .B(n1948), .Y(n1421) );
  NOR2X1 U1031 ( .A(n1991), .B(n1948), .Y(n1422) );
  NOR2X1 U1032 ( .A(n1937), .B(n1949), .Y(n1423) );
  NOR2X1 U1033 ( .A(n1937), .B(n1921), .Y(n1424) );
  NOR2X1 U1034 ( .A(n1937), .B(n1952), .Y(n1425) );
  NOR2X1 U1035 ( .A(n1937), .B(n1938), .Y(n1426) );
  NOR2X1 U1036 ( .A(n1937), .B(n1955), .Y(n1427) );
  NOR2X1 U1037 ( .A(n1923), .B(n1937), .Y(n1428) );
  NOR2X1 U1038 ( .A(n1786), .B(n1937), .Y(n1429) );
  NOR2X1 U1039 ( .A(n1918), .B(n1937), .Y(n1430) );
  NOR2X1 U1040 ( .A(n1964), .B(n1937), .Y(n1431) );
  NOR2X1 U1041 ( .A(n1915), .B(n1937), .Y(n1432) );
  NOR2X1 U1042 ( .A(n1969), .B(n1937), .Y(n1433) );
  NOR2X1 U1043 ( .A(n1926), .B(n1937), .Y(n1434) );
  NOR2X1 U1044 ( .A(n1971), .B(n1937), .Y(n1435) );
  NOR2X1 U1045 ( .A(n1929), .B(n1937), .Y(n1436) );
  NOR2X1 U1050 ( .A(n1983), .B(n1937), .Y(n1441) );
  NOR2X1 U1052 ( .A(n1986), .B(n1937), .Y(n1443) );
  NOR2X1 U1053 ( .A(n1991), .B(n1937), .Y(n1444) );
  NOR2X1 U1054 ( .A(n1950), .B(n1921), .Y(n1445) );
  NOR2X1 U1055 ( .A(n1950), .B(n1952), .Y(n1446) );
  NOR2X1 U1056 ( .A(n1950), .B(n1938), .Y(n1447) );
  NOR2X1 U1057 ( .A(n1950), .B(n1955), .Y(n1448) );
  NOR2X1 U1058 ( .A(n1923), .B(n1950), .Y(n1449) );
  NOR2X1 U1059 ( .A(n1787), .B(n1950), .Y(n1450) );
  NOR2X1 U1060 ( .A(n1918), .B(n1949), .Y(n1451) );
  NOR2X1 U1061 ( .A(n1964), .B(n1949), .Y(n1452) );
  NOR2X1 U1062 ( .A(n1915), .B(n1949), .Y(n1453) );
  NOR2X1 U1063 ( .A(n1968), .B(n1949), .Y(n1454) );
  NOR2X1 U1064 ( .A(n1926), .B(n1949), .Y(n1455) );
  NOR2X1 U1065 ( .A(n1972), .B(n1949), .Y(n1456) );
  NOR2X1 U1066 ( .A(n1929), .B(n1949), .Y(n1457) );
  NOR2X1 U1067 ( .A(n1975), .B(n1949), .Y(n1458) );
  NOR2X1 U1068 ( .A(n1931), .B(n1949), .Y(n1459) );
  NOR2X1 U1069 ( .A(n1979), .B(n1949), .Y(n1460) );
  NOR2X1 U1070 ( .A(n1934), .B(n1949), .Y(n1461) );
  NOR2X1 U1071 ( .A(n1983), .B(n1950), .Y(n1462) );
  NOR2X1 U1072 ( .A(n1935), .B(n1950), .Y(n1463) );
  NOR2X1 U1073 ( .A(n1986), .B(n1950), .Y(n1464) );
  NOR2X1 U1074 ( .A(n1991), .B(n1950), .Y(n1465) );
  NOR2X1 U1075 ( .A(n1921), .B(n1952), .Y(n1466) );
  NOR2X1 U1076 ( .A(n1921), .B(n1938), .Y(n1467) );
  NOR2X1 U1077 ( .A(n1921), .B(n1955), .Y(n1468) );
  NOR2X1 U1078 ( .A(n1923), .B(n1921), .Y(n1469) );
  NOR2X1 U1079 ( .A(n1787), .B(n1921), .Y(n1470) );
  NOR2X1 U1080 ( .A(n1918), .B(n1920), .Y(n1471) );
  NOR2X1 U1081 ( .A(n1964), .B(n1921), .Y(n1472) );
  NOR2X1 U1082 ( .A(n1915), .B(n1921), .Y(n1473) );
  NOR2X1 U1083 ( .A(n1968), .B(n1921), .Y(n1474) );
  NOR2X1 U1084 ( .A(n1926), .B(n1921), .Y(n1475) );
  NOR2X1 U1085 ( .A(n1971), .B(n1921), .Y(n1476) );
  NOR2X1 U1086 ( .A(n1929), .B(n1920), .Y(n1477) );
  NOR2X1 U1088 ( .A(n1931), .B(n1920), .Y(n1479) );
  NOR2X1 U1089 ( .A(n1979), .B(n1920), .Y(n1480) );
  NOR2X1 U1090 ( .A(n1934), .B(n1921), .Y(n1481) );
  NOR2X1 U1091 ( .A(n1983), .B(n1921), .Y(n1482) );
  NOR2X1 U1092 ( .A(n1935), .B(n1921), .Y(n1483) );
  NOR2X1 U1093 ( .A(n1986), .B(n1920), .Y(n1484) );
  NOR2X1 U1094 ( .A(n1991), .B(n1920), .Y(n1485) );
  NOR2X1 U1095 ( .A(n1952), .B(n1938), .Y(n1486) );
  NOR2X1 U1096 ( .A(n1953), .B(n1955), .Y(n1487) );
  NOR2X1 U1097 ( .A(n1923), .B(n1951), .Y(n1488) );
  NOR2X1 U1098 ( .A(n1786), .B(n1951), .Y(n1489) );
  NOR2X1 U1099 ( .A(n1918), .B(n1951), .Y(n1490) );
  NOR2X1 U1100 ( .A(n1964), .B(n1951), .Y(n1491) );
  NOR2X1 U1101 ( .A(n1915), .B(n1952), .Y(n1492) );
  NOR2X1 U1102 ( .A(n1968), .B(n1951), .Y(n1493) );
  NOR2X1 U1103 ( .A(n1926), .B(n1951), .Y(n1494) );
  NOR2X1 U1104 ( .A(n1971), .B(n1951), .Y(n1495) );
  NOR2X1 U1105 ( .A(n1929), .B(n1951), .Y(n1496) );
  NOR2X1 U1106 ( .A(n1974), .B(n1951), .Y(n1497) );
  NOR2X1 U1108 ( .A(n1979), .B(n1951), .Y(n1499) );
  NOR2X1 U1109 ( .A(n1934), .B(n1951), .Y(n1500) );
  NOR2X1 U1110 ( .A(n1983), .B(n1952), .Y(n1501) );
  NOR2X1 U1111 ( .A(n1935), .B(n1952), .Y(n1502) );
  NOR2X1 U1112 ( .A(n1986), .B(n1952), .Y(n1503) );
  NOR2X1 U1113 ( .A(n1991), .B(n1952), .Y(n1504) );
  NOR2X1 U1114 ( .A(n1938), .B(n1955), .Y(n1505) );
  NOR2X1 U1115 ( .A(n1923), .B(n1938), .Y(n1506) );
  NOR2X1 U1116 ( .A(n1786), .B(n1938), .Y(n1507) );
  NOR2X1 U1117 ( .A(n1918), .B(n1938), .Y(n1508) );
  NOR2X1 U1118 ( .A(n1964), .B(n1938), .Y(n1509) );
  NOR2X1 U1119 ( .A(n1915), .B(n1938), .Y(n1510) );
  NOR2X1 U1120 ( .A(n1968), .B(n1938), .Y(n1511) );
  NOR2X1 U1121 ( .A(n1926), .B(n1938), .Y(n1512) );
  NOR2X1 U1122 ( .A(n1971), .B(n1938), .Y(n1513) );
  NOR2X1 U1123 ( .A(n1929), .B(n1938), .Y(n1514) );
  NOR2X1 U1124 ( .A(n1974), .B(n1938), .Y(n1515) );
  NOR2X1 U1125 ( .A(n1931), .B(n1938), .Y(n1516) );
  NOR2X1 U1126 ( .A(n1979), .B(n1938), .Y(n1517) );
  NOR2X1 U1127 ( .A(n1934), .B(n1938), .Y(n1518) );
  NOR2X1 U1128 ( .A(n1983), .B(n1938), .Y(n1519) );
  NOR2X1 U1129 ( .A(n1935), .B(n1938), .Y(n1520) );
  NOR2X1 U1130 ( .A(n1986), .B(n1938), .Y(n1521) );
  NOR2X1 U1131 ( .A(n1991), .B(n1938), .Y(n1522) );
  NOR2X1 U1132 ( .A(n1923), .B(n1954), .Y(n1523) );
  NOR2X1 U1133 ( .A(n1786), .B(n1954), .Y(n1524) );
  NOR2X1 U1134 ( .A(n1918), .B(n1954), .Y(n1525) );
  NOR2X1 U1135 ( .A(n1964), .B(n1954), .Y(n1526) );
  NOR2X1 U1136 ( .A(n1915), .B(n1954), .Y(n1527) );
  NOR2X1 U1139 ( .A(n1971), .B(n1954), .Y(n1530) );
  NOR2X1 U1140 ( .A(n1929), .B(n1954), .Y(n1531) );
  NOR2X1 U1141 ( .A(n1975), .B(n1954), .Y(n1532) );
  NOR2X1 U1143 ( .A(n1979), .B(n1954), .Y(n1534) );
  NOR2X1 U1144 ( .A(n1934), .B(n1955), .Y(n1535) );
  NOR2X1 U1145 ( .A(n1983), .B(n1955), .Y(n1536) );
  NOR2X1 U1147 ( .A(n1986), .B(n1955), .Y(n1538) );
  NOR2X1 U1148 ( .A(n1991), .B(n1955), .Y(n1539) );
  NOR2X1 U1149 ( .A(n1923), .B(n1784), .Y(n1540) );
  NOR2X1 U1150 ( .A(n1923), .B(n1917), .Y(n1541) );
  NOR2X1 U1151 ( .A(n1922), .B(n1965), .Y(n1542) );
  NOR2X1 U1152 ( .A(n1922), .B(n1914), .Y(n1543) );
  NOR2X1 U1153 ( .A(n1922), .B(n1967), .Y(n1544) );
  NOR2X1 U1154 ( .A(n1922), .B(n1926), .Y(n1545) );
  NOR2X1 U1156 ( .A(n1929), .B(n1923), .Y(n1547) );
  NOR2X1 U1157 ( .A(n1974), .B(n1923), .Y(n1548) );
  NOR2X1 U1158 ( .A(n1931), .B(n1923), .Y(n1549) );
  NOR2X1 U1159 ( .A(n1979), .B(n1923), .Y(n1550) );
  NOR2X1 U1160 ( .A(n1934), .B(n1924), .Y(n1551) );
  NOR2X1 U1161 ( .A(n1983), .B(n1922), .Y(n1552) );
  NOR2X1 U1162 ( .A(n1935), .B(n1923), .Y(n1553) );
  NOR2X1 U1163 ( .A(n1986), .B(n1923), .Y(n1554) );
  NOR2X1 U1164 ( .A(n1991), .B(n1923), .Y(n1555) );
  NOR2X1 U1165 ( .A(n1961), .B(n1917), .Y(n1556) );
  NOR2X1 U1166 ( .A(n1786), .B(n1965), .Y(n1557) );
  NOR2X1 U1167 ( .A(n1916), .B(n1787), .Y(n1558) );
  NOR2X1 U1168 ( .A(n1967), .B(n1785), .Y(n1559) );
  NOR2X1 U1169 ( .A(n1926), .B(n1787), .Y(n1560) );
  NOR2X1 U1170 ( .A(n1971), .B(n1784), .Y(n1561) );
  NOR2X1 U1171 ( .A(n1928), .B(n1784), .Y(n1562) );
  NOR2X1 U1172 ( .A(n1974), .B(n1784), .Y(n1563) );
  NOR2X1 U1173 ( .A(n1930), .B(n1783), .Y(n1564) );
  NOR2X1 U1174 ( .A(n1978), .B(n1783), .Y(n1565) );
  NOR2X1 U1175 ( .A(n1933), .B(n1784), .Y(n1566) );
  NOR2X1 U1176 ( .A(n1982), .B(n1783), .Y(n1567) );
  NOR2X1 U1177 ( .A(n1936), .B(n1784), .Y(n1568) );
  NOR2X1 U1178 ( .A(n1985), .B(n1784), .Y(n1569) );
  NOR2X1 U1179 ( .A(n1990), .B(n1784), .Y(n1570) );
  NOR2X1 U1180 ( .A(n1705), .B(n1965), .Y(n1571) );
  NOR2X1 U1181 ( .A(n1916), .B(n1918), .Y(n1572) );
  NOR2X1 U1182 ( .A(n1967), .B(n1918), .Y(n1573) );
  NOR2X1 U1183 ( .A(n1926), .B(n1918), .Y(n1574) );
  NOR2X1 U1184 ( .A(n1971), .B(n1918), .Y(n1575) );
  NOR2X1 U1185 ( .A(n1928), .B(n1917), .Y(n1576) );
  NOR2X1 U1186 ( .A(n1974), .B(n1917), .Y(n1577) );
  NOR2X1 U1187 ( .A(n1930), .B(n1917), .Y(n1578) );
  NOR2X1 U1188 ( .A(n1978), .B(n1917), .Y(n1579) );
  NOR2X1 U1189 ( .A(n1933), .B(n1917), .Y(n1580) );
  NOR2X1 U1190 ( .A(n1982), .B(n1917), .Y(n1581) );
  NOR2X1 U1191 ( .A(n1936), .B(n1917), .Y(n1582) );
  NOR2X1 U1192 ( .A(n1985), .B(n1917), .Y(n1583) );
  NOR2X1 U1193 ( .A(n1990), .B(n1917), .Y(n1584) );
  NOR2X1 U1195 ( .A(n1967), .B(n1965), .Y(n1586) );
  NOR2X1 U1196 ( .A(n1926), .B(n1964), .Y(n1587) );
  NOR2X1 U1197 ( .A(n1971), .B(n1964), .Y(n1588) );
  NOR2X1 U1198 ( .A(n1928), .B(n1966), .Y(n1589) );
  NOR2X1 U1199 ( .A(n1975), .B(n1965), .Y(n1590) );
  NOR2X1 U1200 ( .A(n1930), .B(n1964), .Y(n1591) );
  NOR2X1 U1201 ( .A(n1978), .B(n1965), .Y(n1592) );
  NOR2X1 U1202 ( .A(n1933), .B(n1964), .Y(n1593) );
  NOR2X1 U1203 ( .A(n1982), .B(n1966), .Y(n1594) );
  NOR2X1 U1204 ( .A(n1936), .B(n1964), .Y(n1595) );
  NOR2X1 U1205 ( .A(n1985), .B(n1964), .Y(n1596) );
  NOR2X1 U1206 ( .A(n1990), .B(n1964), .Y(n1597) );
  NOR2X1 U1207 ( .A(n1916), .B(n1969), .Y(n1598) );
  NOR2X1 U1208 ( .A(n1916), .B(n1925), .Y(n1599) );
  NOR2X1 U1209 ( .A(n1916), .B(n1970), .Y(n1600) );
  NOR2X1 U1210 ( .A(n1929), .B(n1914), .Y(n1601) );
  NOR2X1 U1211 ( .A(n1974), .B(n1914), .Y(n1602) );
  NOR2X1 U1212 ( .A(n1930), .B(n1914), .Y(n1603) );
  NOR2X1 U1213 ( .A(n1978), .B(n1914), .Y(n1604) );
  NOR2X1 U1214 ( .A(n1933), .B(n1914), .Y(n1605) );
  NOR2X1 U1215 ( .A(n1982), .B(n1914), .Y(n1606) );
  NOR2X1 U1216 ( .A(n1936), .B(n1914), .Y(n1607) );
  NOR2X1 U1217 ( .A(n1985), .B(n1914), .Y(n1608) );
  NOR2X1 U1218 ( .A(n1990), .B(n1914), .Y(n1609) );
  NOR2X1 U1219 ( .A(n1968), .B(n1925), .Y(n1610) );
  NOR2X1 U1220 ( .A(n1969), .B(n1970), .Y(n1611) );
  NOR2X1 U1221 ( .A(n1929), .B(n1968), .Y(n1612) );
  NOR2X1 U1222 ( .A(n1974), .B(n1967), .Y(n1613) );
  NOR2X1 U1223 ( .A(n1930), .B(n1967), .Y(n1614) );
  NOR2X1 U1224 ( .A(n1978), .B(n1968), .Y(n1615) );
  NOR2X1 U1225 ( .A(n1933), .B(n1968), .Y(n1616) );
  NOR2X1 U1226 ( .A(n1982), .B(n1968), .Y(n1617) );
  NOR2X1 U1227 ( .A(n1936), .B(n1968), .Y(n1618) );
  NOR2X1 U1228 ( .A(n1985), .B(n1969), .Y(n1619) );
  NOR2X1 U1229 ( .A(n1990), .B(n1969), .Y(n1620) );
  NOR2X1 U1230 ( .A(n1925), .B(n1970), .Y(n1621) );
  NOR2X1 U1231 ( .A(n1929), .B(n1925), .Y(n1622) );
  NOR2X1 U1232 ( .A(n1975), .B(n1925), .Y(n1623) );
  NOR2X1 U1233 ( .A(n1930), .B(n1925), .Y(n1624) );
  NOR2X1 U1234 ( .A(n1979), .B(n1925), .Y(n1625) );
  NOR2X1 U1235 ( .A(n1933), .B(n1925), .Y(n1626) );
  NOR2X1 U1236 ( .A(n1982), .B(n1925), .Y(n1627) );
  NOR2X1 U1237 ( .A(n1936), .B(n1925), .Y(n1628) );
  NOR2X1 U1238 ( .A(n1985), .B(n1925), .Y(n1629) );
  NOR2X1 U1239 ( .A(n1990), .B(n1925), .Y(n1630) );
  NOR2X1 U1241 ( .A(n1974), .B(n1970), .Y(n1632) );
  NOR2X1 U1242 ( .A(n1931), .B(n1971), .Y(n1633) );
  NOR2X1 U1243 ( .A(n1979), .B(n1971), .Y(n1634) );
  NOR2X1 U1244 ( .A(n1933), .B(n1970), .Y(n1635) );
  NOR2X1 U1245 ( .A(n1982), .B(n1970), .Y(n1636) );
  NOR2X1 U1246 ( .A(n1936), .B(n1970), .Y(n1637) );
  NOR2X1 U1247 ( .A(n1985), .B(n1970), .Y(n1638) );
  NOR2X1 U1248 ( .A(n1990), .B(n1970), .Y(n1639) );
  NOR2X1 U1249 ( .A(n1974), .B(n1928), .Y(n1640) );
  NOR2X1 U1250 ( .A(n1931), .B(n1928), .Y(n1641) );
  NOR2X1 U1251 ( .A(n1979), .B(n1928), .Y(n1642) );
  NOR2X1 U1252 ( .A(n1933), .B(n1928), .Y(n1643) );
  NOR2X1 U1253 ( .A(n1982), .B(n1928), .Y(n1644) );
  NOR2X1 U1254 ( .A(n1936), .B(n1928), .Y(n1645) );
  NOR2X1 U1255 ( .A(n1985), .B(n1928), .Y(n1646) );
  NOR2X1 U1256 ( .A(n1990), .B(n1928), .Y(n1647) );
  NOR2X1 U1257 ( .A(n95), .B(n1973), .Y(n1648) );
  NOR2X1 U1258 ( .A(n1979), .B(n1974), .Y(n1649) );
  NOR2X1 U1259 ( .A(n1933), .B(n1973), .Y(n1650) );
  NOR2X1 U1260 ( .A(n1982), .B(n1974), .Y(n1651) );
  NOR2X1 U1261 ( .A(n1936), .B(n1974), .Y(n1652) );
  NOR2X1 U1262 ( .A(n1985), .B(n1974), .Y(n1653) );
  NOR2X1 U1263 ( .A(n1990), .B(n1975), .Y(n1654) );
  NOR2X1 U1264 ( .A(n1931), .B(n1978), .Y(n1655) );
  NOR2X1 U1265 ( .A(n1934), .B(n1930), .Y(n1656) );
  NOR2X1 U1266 ( .A(n1982), .B(n1930), .Y(n1657) );
  NOR2X1 U1267 ( .A(n1935), .B(n1930), .Y(n1658) );
  NOR2X1 U1268 ( .A(n1985), .B(n1930), .Y(n1659) );
  NOR2X1 U1269 ( .A(n1990), .B(n1930), .Y(n1660) );
  NOR2X1 U1270 ( .A(n1934), .B(n1978), .Y(n1661) );
  NOR2X1 U1271 ( .A(n1983), .B(n1978), .Y(n1662) );
  NOR2X1 U1272 ( .A(n1936), .B(n1978), .Y(n1663) );
  NOR2X1 U1273 ( .A(n1985), .B(n1978), .Y(n1664) );
  NOR2X1 U1274 ( .A(n1990), .B(n1978), .Y(n1665) );
  NOR2X1 U1275 ( .A(n1983), .B(n1933), .Y(n1666) );
  NOR2X1 U1276 ( .A(n1935), .B(n1933), .Y(n1667) );
  NOR2X1 U1277 ( .A(n1985), .B(n1933), .Y(n1668) );
  NOR2X1 U1278 ( .A(n1990), .B(n1933), .Y(n1669) );
  NOR2X1 U1279 ( .A(n1935), .B(n1982), .Y(n1670) );
  NOR2X1 U1280 ( .A(n1986), .B(n1982), .Y(n1671) );
  NOR2X1 U1281 ( .A(n1991), .B(n1982), .Y(n1672) );
  NOR2X1 U1282 ( .A(n1986), .B(n1936), .Y(n1673) );
  NOR2X1 U1284 ( .A(n1991), .B(n1985), .Y(n1675) );
  INVX8 U1341 ( .A(b[29]), .Y(n1942) );
  BUFX2 U1342 ( .A(n1959), .Y(n1783) );
  BUFX4 U1343 ( .A(n1959), .Y(n1784) );
  INVX1 U1344 ( .A(n1957), .Y(n1959) );
  INVX4 U1345 ( .A(b[26]), .Y(n72) );
  INVX4 U1346 ( .A(n103), .Y(n1927) );
  BUFX2 U1347 ( .A(n1960), .Y(n1785) );
  BUFX4 U1348 ( .A(n1960), .Y(n1786) );
  BUFX4 U1349 ( .A(n1960), .Y(n1787) );
  INVX2 U1350 ( .A(b[7]), .Y(n1973) );
  INVX4 U1351 ( .A(n1981), .Y(n1980) );
  INVX2 U1352 ( .A(b[3]), .Y(n1981) );
  INVX4 U1353 ( .A(b[27]), .Y(n1944) );
  INVX2 U1354 ( .A(n1980), .Y(n1982) );
  INVX2 U1355 ( .A(a[12]), .Y(n1916) );
  INVX2 U1356 ( .A(n1962), .Y(n1965) );
  INVX2 U1357 ( .A(b[16]), .Y(n1922) );
  INVX2 U1358 ( .A(a[28]), .Y(n1800) );
  INVX2 U1359 ( .A(b[0]), .Y(n1989) );
  INVX2 U1360 ( .A(b[10]), .Y(n103) );
  INVX2 U1361 ( .A(b[14]), .Y(n1705) );
  INVX2 U1362 ( .A(b[20]), .Y(n1920) );
  INVX4 U1363 ( .A(n1976), .Y(n1979) );
  INVX4 U1364 ( .A(n1976), .Y(n1978) );
  INVX2 U1365 ( .A(n1980), .Y(n1983) );
  INVX2 U1366 ( .A(n1957), .Y(n1960) );
  INVX4 U1367 ( .A(n1927), .Y(n1926) );
  INVX4 U1368 ( .A(n1927), .Y(n1925) );
  INVX2 U1369 ( .A(n1705), .Y(n1919) );
  INVX2 U1370 ( .A(n1963), .Y(n1962) );
  INVX2 U1371 ( .A(b[13]), .Y(n1963) );
  INVX2 U1372 ( .A(b[19]), .Y(n1951) );
  INVX2 U1373 ( .A(a[12]), .Y(n1915) );
  INVX4 U1374 ( .A(b[12]), .Y(n1914) );
  INVX2 U1375 ( .A(b[31]), .Y(n1939) );
  INVX4 U1376 ( .A(n1958), .Y(n1957) );
  INVX2 U1377 ( .A(b[15]), .Y(n1958) );
  INVX4 U1378 ( .A(n1919), .Y(n1917) );
  INVX4 U1379 ( .A(n1919), .Y(n1918) );
  INVX4 U1380 ( .A(n1962), .Y(n1964) );
  INVX4 U1381 ( .A(a[20]), .Y(n1921) );
  INVX2 U1382 ( .A(b[19]), .Y(n1952) );
  INVX2 U1383 ( .A(n1957), .Y(n1961) );
  INVX4 U1384 ( .A(b[18]), .Y(n1938) );
  INVX4 U1385 ( .A(a[16]), .Y(n1923) );
  INVX2 U1386 ( .A(n1989), .Y(n1988) );
  INVX2 U1387 ( .A(n1988), .Y(n1991) );
  INVX4 U1388 ( .A(a[4]), .Y(n1933) );
  XNOR2X1 U1389 ( .A(n290), .B(n1886), .Y(product[31]) );
  INVX2 U1390 ( .A(b[6]), .Y(n95) );
  INVX4 U1391 ( .A(b[8]), .Y(n1929) );
  XOR2X1 U1392 ( .A(n1625), .B(n1583), .Y(n1789) );
  XOR2X1 U1393 ( .A(n1633), .B(n1789), .Y(n1155) );
  NAND2X1 U1394 ( .A(n1633), .B(n1625), .Y(n1790) );
  NAND2X1 U1395 ( .A(n1633), .B(n1583), .Y(n1791) );
  NAND2X1 U1396 ( .A(n1625), .B(n1583), .Y(n1792) );
  NAND3X1 U1397 ( .A(n1790), .B(n1791), .C(n1792), .Y(n1154) );
  XOR2X1 U1398 ( .A(n982), .B(n961), .Y(n1793) );
  XOR2X1 U1399 ( .A(n1793), .B(n959), .Y(n957) );
  NAND2X1 U1400 ( .A(n959), .B(n982), .Y(n1794) );
  NAND2X1 U1401 ( .A(n959), .B(n961), .Y(n1795) );
  NAND2X1 U1402 ( .A(n982), .B(n961), .Y(n1796) );
  NAND3X1 U1403 ( .A(n1794), .B(n1795), .C(n1796), .Y(n956) );
  BUFX2 U1404 ( .A(n719), .Y(n1797) );
  AND2X2 U1405 ( .A(a[6]), .B(a[17]), .Y(n1533) );
  INVX2 U1406 ( .A(a[6]), .Y(n1931) );
  INVX1 U1407 ( .A(n958), .Y(n1798) );
  INVX2 U1408 ( .A(n1798), .Y(n1799) );
  NOR2X1 U1409 ( .A(n1991), .B(n1800), .Y(n1313) );
  AND2X2 U1410 ( .A(a[12]), .B(n1962), .Y(n1585) );
  AND2X2 U1411 ( .A(n1546), .B(n1585), .Y(n1801) );
  BUFX2 U1412 ( .A(n934), .Y(n1802) );
  BUFX2 U1413 ( .A(n1435), .Y(n1803) );
  AND2X2 U1414 ( .A(n980), .B(n957), .Y(n1804) );
  INVX1 U1415 ( .A(n1804), .Y(n327) );
  AND2X2 U1416 ( .A(a[2]), .B(a[17]), .Y(n1537) );
  XOR2X1 U1417 ( .A(n962), .B(n939), .Y(n1805) );
  XOR2X1 U1418 ( .A(n1805), .B(n960), .Y(n935) );
  XOR2X1 U1419 ( .A(n937), .B(n958), .Y(n1806) );
  XOR2X1 U1420 ( .A(n1806), .B(n935), .Y(n933) );
  NAND2X1 U1421 ( .A(n962), .B(n939), .Y(n1807) );
  NAND2X1 U1422 ( .A(n962), .B(n960), .Y(n1808) );
  NAND2X1 U1423 ( .A(n939), .B(n960), .Y(n1809) );
  NAND3X1 U1424 ( .A(n1807), .B(n1808), .C(n1809), .Y(n934) );
  NAND2X1 U1425 ( .A(n937), .B(n1799), .Y(n1810) );
  NAND2X1 U1426 ( .A(n937), .B(n935), .Y(n1811) );
  NAND2X1 U1427 ( .A(n1799), .B(n935), .Y(n1812) );
  NAND3X1 U1428 ( .A(n1810), .B(n1811), .C(n1812), .Y(n932) );
  XOR2X1 U1429 ( .A(n1435), .B(n1414), .Y(n1813) );
  XOR2X1 U1430 ( .A(n1310), .B(n1813), .Y(n819) );
  NAND2X1 U1431 ( .A(n1310), .B(n1803), .Y(n1814) );
  NAND2X1 U1432 ( .A(n1310), .B(n1414), .Y(n1815) );
  NAND2X1 U1433 ( .A(n1803), .B(n1414), .Y(n1816) );
  NAND3X1 U1434 ( .A(n1814), .B(n1815), .C(n1816), .Y(n818) );
  AND2X2 U1435 ( .A(n1927), .B(a[17]), .Y(n1529) );
  XOR2X1 U1436 ( .A(n761), .B(n759), .Y(n1817) );
  XOR2X1 U1437 ( .A(n1817), .B(n782), .Y(n749) );
  NAND2X1 U1438 ( .A(n761), .B(n759), .Y(n1818) );
  NAND2X1 U1439 ( .A(n761), .B(n782), .Y(n1819) );
  NAND2X1 U1440 ( .A(n759), .B(n782), .Y(n1820) );
  NAND3X1 U1441 ( .A(n1818), .B(n1819), .C(n1820), .Y(n748) );
  XOR2X1 U1442 ( .A(n727), .B(n725), .Y(n1821) );
  XOR2X1 U1443 ( .A(n1821), .B(n748), .Y(n719) );
  NAND2X1 U1444 ( .A(n727), .B(n725), .Y(n1822) );
  NAND2X1 U1445 ( .A(n727), .B(n748), .Y(n1823) );
  NAND2X1 U1446 ( .A(n725), .B(n748), .Y(n1824) );
  NAND3X1 U1447 ( .A(n1822), .B(n1823), .C(n1824), .Y(n718) );
  XOR2X1 U1448 ( .A(n1477), .B(n1495), .Y(n1825) );
  XOR2X1 U1449 ( .A(n1512), .B(n1825), .Y(n899) );
  NAND2X1 U1450 ( .A(n1512), .B(n1477), .Y(n1826) );
  NAND2X1 U1451 ( .A(n1512), .B(n1495), .Y(n1827) );
  NAND2X1 U1452 ( .A(n1477), .B(n1495), .Y(n1828) );
  NAND3X1 U1453 ( .A(n1826), .B(n1827), .C(n1828), .Y(n898) );
  INVX1 U1454 ( .A(n393), .Y(n392) );
  XOR2X1 U1455 ( .A(n938), .B(n913), .Y(n1829) );
  XOR2X1 U1456 ( .A(n1829), .B(n936), .Y(n909) );
  XOR2X1 U1457 ( .A(n911), .B(n934), .Y(n1830) );
  XOR2X1 U1458 ( .A(n1830), .B(n909), .Y(n907) );
  NAND2X1 U1459 ( .A(n938), .B(n913), .Y(n1831) );
  NAND2X1 U1460 ( .A(n938), .B(n936), .Y(n1832) );
  NAND2X1 U1461 ( .A(n913), .B(n936), .Y(n1833) );
  NAND3X1 U1462 ( .A(n1831), .B(n1832), .C(n1833), .Y(n908) );
  NAND2X1 U1463 ( .A(n911), .B(n1802), .Y(n1834) );
  NAND2X1 U1464 ( .A(n911), .B(n909), .Y(n1835) );
  NAND2X1 U1465 ( .A(n1802), .B(n909), .Y(n1836) );
  NAND3X1 U1466 ( .A(n1834), .B(n1835), .C(n1836), .Y(n906) );
  XOR2X1 U1467 ( .A(n1093), .B(n1108), .Y(n1837) );
  XOR2X1 U1468 ( .A(n1841), .B(n1837), .Y(n1087) );
  NAND2X1 U1469 ( .A(n1106), .B(n1093), .Y(n1838) );
  NAND2X1 U1470 ( .A(n1106), .B(n1108), .Y(n1839) );
  NAND2X1 U1471 ( .A(n1093), .B(n1108), .Y(n1840) );
  NAND3X1 U1472 ( .A(n1838), .B(n1839), .C(n1840), .Y(n1086) );
  BUFX2 U1473 ( .A(n1106), .Y(n1841) );
  XOR2X1 U1474 ( .A(n996), .B(n977), .Y(n1842) );
  XOR2X1 U1475 ( .A(n994), .B(n1842), .Y(n967) );
  NAND2X1 U1476 ( .A(n994), .B(n996), .Y(n1843) );
  NAND2X1 U1477 ( .A(n994), .B(n977), .Y(n1844) );
  NAND2X1 U1478 ( .A(n996), .B(n977), .Y(n1845) );
  NAND3X1 U1479 ( .A(n1843), .B(n1844), .C(n1845), .Y(n966) );
  AND2X2 U1480 ( .A(a[11]), .B(b[17]), .Y(n1528) );
  INVX1 U1481 ( .A(n1893), .Y(n1846) );
  INVX2 U1482 ( .A(n1846), .Y(n1847) );
  AND2X2 U1483 ( .A(b[16]), .B(a[9]), .Y(n1546) );
  XOR2X1 U1484 ( .A(n1482), .B(n1533), .Y(n1848) );
  XOR2X1 U1485 ( .A(n1042), .B(n1848), .Y(n1015) );
  NAND2X1 U1486 ( .A(n1042), .B(n1482), .Y(n1849) );
  NAND2X1 U1487 ( .A(n1042), .B(n1533), .Y(n1850) );
  NAND2X1 U1488 ( .A(n1482), .B(n1533), .Y(n1851) );
  NAND3X1 U1489 ( .A(n1849), .B(n1850), .C(n1851), .Y(n1014) );
  BUFX2 U1490 ( .A(n1009), .Y(n1852) );
  XOR2X1 U1491 ( .A(n1035), .B(n1052), .Y(n1853) );
  XOR2X1 U1492 ( .A(n1853), .B(n1050), .Y(n1029) );
  NAND2X1 U1493 ( .A(n1035), .B(n1052), .Y(n1854) );
  NAND2X1 U1494 ( .A(n1035), .B(n1050), .Y(n1855) );
  NAND2X1 U1495 ( .A(n1052), .B(n1050), .Y(n1856) );
  NAND3X1 U1496 ( .A(n1854), .B(n1855), .C(n1856), .Y(n1028) );
  XOR2X1 U1497 ( .A(n1011), .B(n1009), .Y(n1857) );
  XOR2X1 U1498 ( .A(n1857), .B(n1028), .Y(n1005) );
  NAND2X1 U1499 ( .A(n1011), .B(n1852), .Y(n1858) );
  NAND2X1 U1500 ( .A(n1011), .B(n1028), .Y(n1859) );
  NAND2X1 U1501 ( .A(n1852), .B(n1028), .Y(n1860) );
  NAND3X1 U1502 ( .A(n1858), .B(n1859), .C(n1860), .Y(n1004) );
  XOR2X1 U1503 ( .A(n719), .B(n744), .Y(n1861) );
  XOR2X1 U1504 ( .A(n742), .B(n1861), .Y(n715) );
  NAND2X1 U1505 ( .A(n742), .B(n1797), .Y(n1862) );
  NAND2X1 U1506 ( .A(n742), .B(n744), .Y(n1863) );
  NAND2X1 U1507 ( .A(n1797), .B(n744), .Y(n1864) );
  NAND3X1 U1508 ( .A(n1862), .B(n1863), .C(n1864), .Y(n714) );
  XOR2X1 U1509 ( .A(n775), .B(n773), .Y(n1865) );
  XOR2X1 U1510 ( .A(n1865), .B(n798), .Y(n769) );
  XOR2X1 U1511 ( .A(n771), .B(n796), .Y(n1866) );
  XOR2X1 U1512 ( .A(n1866), .B(n769), .Y(n767) );
  NAND2X1 U1513 ( .A(n775), .B(n773), .Y(n1867) );
  NAND2X1 U1514 ( .A(n775), .B(n798), .Y(n1868) );
  NAND2X1 U1515 ( .A(n773), .B(n798), .Y(n1869) );
  NAND3X1 U1516 ( .A(n1867), .B(n1868), .C(n1869), .Y(n768) );
  NAND2X1 U1517 ( .A(n771), .B(n796), .Y(n1870) );
  NAND2X1 U1518 ( .A(n771), .B(n769), .Y(n1871) );
  NAND2X1 U1519 ( .A(n796), .B(n769), .Y(n1872) );
  NAND3X1 U1520 ( .A(n1870), .B(n1871), .C(n1872), .Y(n766) );
  AND2X2 U1521 ( .A(a[7]), .B(a[22]), .Y(n1437) );
  AND2X2 U1522 ( .A(a[6]), .B(b[19]), .Y(n1498) );
  AND2X2 U1523 ( .A(a[1]), .B(b[28]), .Y(n1312) );
  XOR2X1 U1524 ( .A(n873), .B(n871), .Y(n1873) );
  XOR2X1 U1525 ( .A(n1873), .B(n875), .Y(n863) );
  NAND2X1 U1526 ( .A(n875), .B(n873), .Y(n1874) );
  NAND2X1 U1527 ( .A(n875), .B(n871), .Y(n1875) );
  NAND2X1 U1528 ( .A(n873), .B(n871), .Y(n1876) );
  NAND3X1 U1529 ( .A(n1874), .B(n1875), .C(n1876), .Y(n862) );
  AND2X2 U1530 ( .A(a[8]), .B(a[9]), .Y(n1631) );
  AND2X2 U1531 ( .A(n1976), .B(a[22]), .Y(n1439) );
  XOR2X1 U1532 ( .A(n1546), .B(n1585), .Y(n979) );
  INVX1 U1533 ( .A(n343), .Y(n470) );
  AND2X2 U1534 ( .A(a[2]), .B(a[22]), .Y(n1442) );
  INVX2 U1535 ( .A(b[2]), .Y(n1935) );
  INVX1 U1536 ( .A(n384), .Y(n383) );
  INVX1 U1537 ( .A(n387), .Y(n477) );
  AND2X2 U1538 ( .A(a[7]), .B(a[20]), .Y(n1478) );
  AND2X2 U1539 ( .A(a[6]), .B(a[22]), .Y(n1438) );
  AND2X2 U1540 ( .A(a[4]), .B(a[22]), .Y(n1440) );
  INVX2 U1541 ( .A(b[4]), .Y(n1934) );
  INVX8 U1542 ( .A(a[9]), .Y(n1971) );
  INVX2 U1543 ( .A(n1988), .Y(n1992) );
  XOR2X1 U1544 ( .A(n1460), .B(n1354), .Y(n1878) );
  XOR2X1 U1545 ( .A(n1801), .B(n1878), .Y(n947) );
  NAND2X1 U1546 ( .A(n1801), .B(n1460), .Y(n1879) );
  NAND2X1 U1547 ( .A(n1801), .B(n1354), .Y(n1880) );
  NAND2X1 U1548 ( .A(n1460), .B(n1354), .Y(n1881) );
  NAND3X1 U1549 ( .A(n1881), .B(n1880), .C(n1879), .Y(n946) );
  INVX4 U1550 ( .A(a[8]), .Y(n1928) );
  INVX2 U1551 ( .A(a[1]), .Y(n1987) );
  BUFX2 U1552 ( .A(n72), .Y(n1882) );
  OR2X1 U1553 ( .A(n160), .B(n163), .Y(n1890) );
  INVX1 U1554 ( .A(n159), .Y(n157) );
  XNOR2X1 U1555 ( .A(n155), .B(n121), .Y(product[47]) );
  AND2X2 U1556 ( .A(n1172), .B(n1161), .Y(n1905) );
  OR2X1 U1557 ( .A(n1232), .B(n1227), .Y(n1898) );
  OR2X1 U1558 ( .A(n1220), .B(n1213), .Y(n1902) );
  OR2X1 U1559 ( .A(n1184), .B(n1173), .Y(n1906) );
  OR2X1 U1560 ( .A(n486), .B(n479), .Y(n1884) );
  INVX2 U1561 ( .A(a[2]), .Y(n1936) );
  XNOR2X1 U1562 ( .A(n1885), .B(n1994), .Y(n1993) );
  XNOR2X1 U1563 ( .A(n1997), .B(n1377), .Y(n1885) );
  OR2X1 U1564 ( .A(n1672), .B(n1243), .Y(n1907) );
  INVX2 U1565 ( .A(b[9]), .Y(n1972) );
  INVX4 U1566 ( .A(a[7]), .Y(n1975) );
  INVX2 U1567 ( .A(n1980), .Y(n1984) );
  INVX8 U1568 ( .A(a[11]), .Y(n1968) );
  INVX8 U1569 ( .A(a[1]), .Y(n1986) );
  INVX8 U1570 ( .A(b[22]), .Y(n1937) );
  OR2X1 U1571 ( .A(n1239), .B(n1237), .Y(n1909) );
  AND2X2 U1572 ( .A(n1239), .B(n1237), .Y(n1910) );
  INVX8 U1573 ( .A(b[29]), .Y(n1941) );
  INVX8 U1574 ( .A(b[25]), .Y(n1945) );
  AND2X2 U1575 ( .A(n289), .B(n463), .Y(n1886) );
  OR2X2 U1576 ( .A(n932), .B(n907), .Y(n1887) );
  OR2X2 U1577 ( .A(n906), .B(n881), .Y(n1888) );
  XNOR2X1 U1578 ( .A(n378), .B(n1889), .Y(product[19]) );
  AND2X2 U1579 ( .A(n377), .B(n1899), .Y(n1889) );
  OR2X2 U1580 ( .A(n575), .B(n594), .Y(n1891) );
  OR2X2 U1581 ( .A(n956), .B(n933), .Y(n1892) );
  OR2X2 U1582 ( .A(n1082), .B(n1065), .Y(n1893) );
  OR2X2 U1583 ( .A(n518), .B(n503), .Y(n1894) );
  OR2X2 U1584 ( .A(n574), .B(n555), .Y(n1895) );
  OR2X2 U1585 ( .A(n1002), .B(n981), .Y(n1896) );
  AND2X1 U1586 ( .A(n1232), .B(n1227), .Y(n1897) );
  OR2X2 U1587 ( .A(n1116), .B(n1101), .Y(n1899) );
  OR2X2 U1588 ( .A(n1132), .B(n1117), .Y(n1900) );
  OR2X2 U1589 ( .A(n1172), .B(n1161), .Y(n1901) );
  AND2X1 U1590 ( .A(n1184), .B(n1173), .Y(n1903) );
  AND2X1 U1591 ( .A(n1220), .B(n1213), .Y(n1904) );
  INVX4 U1592 ( .A(n1988), .Y(n1990) );
  INVX1 U1593 ( .A(b[31]), .Y(n1940) );
  AND2X1 U1594 ( .A(n1672), .B(n1243), .Y(n1908) );
  INVX4 U1595 ( .A(a[6]), .Y(n1930) );
  INVX1 U1596 ( .A(n1962), .Y(n1966) );
  INVX4 U1597 ( .A(a[11]), .Y(n1969) );
  INVX1 U1598 ( .A(a[6]), .Y(n1932) );
  INVX1 U1599 ( .A(a[17]), .Y(n1956) );
  INVX1 U1600 ( .A(a[16]), .Y(n1924) );
  NOR2X1 U1601 ( .A(n446), .B(n1912), .Y(n1911) );
  OR2X2 U1602 ( .A(n1991), .B(n1936), .Y(n1912) );
  INVX1 U1603 ( .A(b[19]), .Y(n1953) );
  INVX4 U1604 ( .A(b[21]), .Y(n1950) );
  INVX1 U1605 ( .A(n351), .Y(n350) );
  INVX1 U1606 ( .A(n272), .Y(n461) );
  INVX1 U1607 ( .A(n315), .Y(n317) );
  INVX1 U1608 ( .A(n288), .Y(n463) );
  INVX1 U1609 ( .A(n316), .Y(n318) );
  INVX1 U1610 ( .A(n256), .Y(n254) );
  INVX1 U1611 ( .A(n283), .Y(n285) );
  BUFX4 U1612 ( .A(n120), .Y(n1913) );
  INVX1 U1613 ( .A(n261), .Y(n459) );
  INVX1 U1614 ( .A(n277), .Y(n462) );
  INVX8 U1615 ( .A(b[30]), .Y(n80) );
  INVX8 U1616 ( .A(b[28]), .Y(n76) );
  INVX8 U1617 ( .A(b[24]), .Y(n68) );
  INVX4 U1618 ( .A(n267), .Y(n266) );
  INVX8 U1619 ( .A(b[27]), .Y(n1943) );
  INVX8 U1620 ( .A(b[25]), .Y(n1946) );
  INVX8 U1621 ( .A(b[23]), .Y(n1947) );
  INVX8 U1622 ( .A(b[23]), .Y(n1948) );
  INVX8 U1623 ( .A(b[21]), .Y(n1949) );
  INVX8 U1624 ( .A(a[17]), .Y(n1954) );
  INVX8 U1625 ( .A(a[17]), .Y(n1955) );
  INVX8 U1626 ( .A(b[11]), .Y(n1967) );
  INVX8 U1627 ( .A(a[9]), .Y(n1970) );
  INVX8 U1628 ( .A(b[7]), .Y(n1974) );
  INVX8 U1629 ( .A(n1977), .Y(n1976) );
  INVX8 U1630 ( .A(b[5]), .Y(n1977) );
  INVX8 U1631 ( .A(b[1]), .Y(n1985) );
  XOR2X1 U1632 ( .A(n488), .B(n1993), .Y(n479) );
  XOR2X1 U1633 ( .A(n490), .B(n1995), .Y(n1994) );
  XOR2X1 U1634 ( .A(n492), .B(n1996), .Y(n1995) );
  XOR2X1 U1635 ( .A(n498), .B(n496), .Y(n1996) );
  XOR2X1 U1636 ( .A(n494), .B(n1998), .Y(n1997) );
  XOR2X1 U1637 ( .A(n1999), .B(n1355), .Y(n1998) );
  XOR2X1 U1638 ( .A(n2000), .B(n2001), .Y(n1999) );
  XOR2X1 U1639 ( .A(n2002), .B(n1295), .Y(n2001) );
  XOR2X1 U1640 ( .A(n2003), .B(n1277), .Y(n2002) );
  XOR2X1 U1641 ( .A(n1260), .B(n1244), .Y(n2003) );
  XOR2X1 U1642 ( .A(n500), .B(n2004), .Y(n2000) );
  XOR2X1 U1643 ( .A(n1334), .B(n1314), .Y(n2004) );
  INVX2 U1644 ( .A(n390), .Y(n478) );
  INVX2 U1645 ( .A(n354), .Y(n472) );
  INVX2 U1646 ( .A(n264), .Y(n460) );
  INVX2 U1647 ( .A(n243), .Y(n457) );
  INVX2 U1648 ( .A(n225), .Y(n455) );
  INVX2 U1649 ( .A(n177), .Y(n451) );
  INVX2 U1650 ( .A(n174), .Y(n450) );
  INVX2 U1651 ( .A(n160), .Y(n448) );
  INVX2 U1652 ( .A(n382), .Y(n380) );
  INVX2 U1653 ( .A(n377), .Y(n375) );
  INVX2 U1654 ( .A(n371), .Y(n370) );
  INVX2 U1655 ( .A(n365), .Y(n367) );
  INVX2 U1656 ( .A(n364), .Y(n474) );
  INVX2 U1657 ( .A(n362), .Y(n360) );
  INVX2 U1658 ( .A(n349), .Y(n347) );
  INVX2 U1659 ( .A(n348), .Y(n471) );
  INVX2 U1660 ( .A(n339), .Y(n337) );
  INVX2 U1661 ( .A(n333), .Y(n332) );
  INVX2 U1662 ( .A(n326), .Y(n468) );
  INVX2 U1663 ( .A(n324), .Y(n322) );
  INVX2 U1664 ( .A(n313), .Y(n311) );
  INVX2 U1665 ( .A(n304), .Y(n302) );
  INVX2 U1666 ( .A(n296), .Y(n295) );
  INVX2 U1667 ( .A(n294), .Y(n292) );
  INVX2 U1668 ( .A(n293), .Y(n464) );
  INVX2 U1669 ( .A(n282), .Y(n284) );
  INVX2 U1670 ( .A(n255), .Y(n253) );
  INVX2 U1671 ( .A(n251), .Y(n249) );
  INVX2 U1672 ( .A(n250), .Y(n458) );
  INVX2 U1673 ( .A(n236), .Y(n238) );
  INVX2 U1674 ( .A(n235), .Y(n237) );
  INVX2 U1675 ( .A(n233), .Y(n231) );
  INVX2 U1676 ( .A(n232), .Y(n456) );
  INVX2 U1677 ( .A(n220), .Y(n222) );
  INVX2 U1678 ( .A(n219), .Y(n221) );
  INVX2 U1679 ( .A(n211), .Y(n213) );
  INVX2 U1680 ( .A(n210), .Y(n454) );
  INVX2 U1681 ( .A(n204), .Y(n202) );
  INVX2 U1682 ( .A(n191), .Y(n189) );
  INVX2 U1683 ( .A(n173), .Y(n171) );
  INVX2 U1684 ( .A(n172), .Y(n170) );
  INVX2 U1685 ( .A(n168), .Y(n166) );
endmodule


module poly5_DW01_sub_78 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n18,
         n19, n20, n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n68, n69, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, \B[0] , n193, n194;
  assign n52 = B[15];
  assign n69 = B[9];
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR2X1 U1 ( .A(n2), .B(B[31]), .Y(DIFF[31]) );
  XNOR2X1 U2 ( .A(n5), .B(B[30]), .Y(DIFF[30]) );
  NOR2X1 U3 ( .A(n194), .B(n1), .Y(n2) );
  XOR2X1 U6 ( .A(n1), .B(B[29]), .Y(DIFF[29]) );
  NOR2X1 U7 ( .A(B[29]), .B(n1), .Y(n5) );
  XNOR2X1 U8 ( .A(n9), .B(B[28]), .Y(DIFF[28]) );
  NAND2X1 U9 ( .A(n27), .B(n6), .Y(n1) );
  NOR2X1 U10 ( .A(n7), .B(n13), .Y(n6) );
  NAND2X1 U11 ( .A(n11), .B(n8), .Y(n7) );
  XNOR2X1 U13 ( .A(n12), .B(B[27]), .Y(DIFF[27]) );
  NOR2X1 U14 ( .A(n26), .B(n10), .Y(n9) );
  NAND2X1 U15 ( .A(n11), .B(n14), .Y(n10) );
  XNOR2X1 U17 ( .A(n17), .B(B[26]), .Y(DIFF[26]) );
  NOR2X1 U18 ( .A(n13), .B(n26), .Y(n12) );
  NAND2X1 U21 ( .A(n16), .B(n22), .Y(n13) );
  NOR2X1 U22 ( .A(B[25]), .B(B[26]), .Y(n16) );
  XNOR2X1 U23 ( .A(n20), .B(B[25]), .Y(DIFF[25]) );
  NOR2X1 U24 ( .A(n18), .B(n26), .Y(n17) );
  NAND2X1 U25 ( .A(n19), .B(n22), .Y(n18) );
  XNOR2X1 U27 ( .A(n25), .B(B[24]), .Y(DIFF[24]) );
  NOR2X1 U28 ( .A(n21), .B(n26), .Y(n20) );
  NOR2X1 U32 ( .A(B[23]), .B(B[24]), .Y(n22) );
  XOR2X1 U33 ( .A(n26), .B(B[23]), .Y(DIFF[23]) );
  NOR2X1 U34 ( .A(B[23]), .B(n26), .Y(n25) );
  XOR2X1 U35 ( .A(n30), .B(B[22]), .Y(DIFF[22]) );
  NOR2X1 U37 ( .A(n39), .B(n28), .Y(n27) );
  NAND2X1 U38 ( .A(n29), .B(n33), .Y(n28) );
  NOR2X1 U39 ( .A(B[21]), .B(B[22]), .Y(n29) );
  XOR2X1 U40 ( .A(n32), .B(B[21]), .Y(DIFF[21]) );
  NAND2X1 U41 ( .A(n38), .B(n31), .Y(n30) );
  NOR2X1 U42 ( .A(B[21]), .B(n34), .Y(n31) );
  XOR2X1 U43 ( .A(n36), .B(B[20]), .Y(DIFF[20]) );
  NAND2X1 U44 ( .A(n33), .B(n38), .Y(n32) );
  NOR2X1 U47 ( .A(B[19]), .B(B[20]), .Y(n33) );
  XNOR2X1 U48 ( .A(n38), .B(B[19]), .Y(DIFF[19]) );
  NAND2X1 U49 ( .A(n37), .B(n38), .Y(n36) );
  XNOR2X1 U51 ( .A(n43), .B(B[18]), .Y(DIFF[18]) );
  NAND2X1 U53 ( .A(n55), .B(n40), .Y(n39) );
  NOR2X1 U54 ( .A(n47), .B(n41), .Y(n40) );
  NAND2X1 U55 ( .A(n45), .B(n42), .Y(n41) );
  XNOR2X1 U57 ( .A(n46), .B(B[17]), .Y(DIFF[17]) );
  NOR2X1 U58 ( .A(n54), .B(n44), .Y(n43) );
  NAND2X1 U59 ( .A(n45), .B(n48), .Y(n44) );
  XNOR2X1 U61 ( .A(n51), .B(B[16]), .Y(DIFF[16]) );
  NOR2X1 U62 ( .A(n47), .B(n54), .Y(n46) );
  NAND2X1 U65 ( .A(n53), .B(n50), .Y(n47) );
  XOR2X1 U67 ( .A(n54), .B(n193), .Y(DIFF[15]) );
  NOR2X1 U68 ( .A(n52), .B(n54), .Y(n51) );
  XOR2X1 U71 ( .A(n58), .B(B[14]), .Y(DIFF[14]) );
  NOR2X1 U73 ( .A(n63), .B(n56), .Y(n55) );
  NAND2X1 U74 ( .A(n57), .B(n59), .Y(n56) );
  XOR2X1 U76 ( .A(n60), .B(B[13]), .Y(DIFF[13]) );
  NAND2X1 U77 ( .A(n59), .B(n62), .Y(n58) );
  NOR2X1 U78 ( .A(B[13]), .B(B[12]), .Y(n59) );
  XNOR2X1 U79 ( .A(n62), .B(B[12]), .Y(DIFF[12]) );
  NAND2X1 U80 ( .A(n61), .B(n62), .Y(n60) );
  XNOR2X1 U82 ( .A(n65), .B(B[11]), .Y(DIFF[11]) );
  NAND2X1 U84 ( .A(n72), .B(n64), .Y(n63) );
  NOR2X1 U85 ( .A(B[11]), .B(n66), .Y(n64) );
  XNOR2X1 U86 ( .A(n68), .B(B[10]), .Y(DIFF[10]) );
  NOR2X1 U87 ( .A(n66), .B(n71), .Y(n65) );
  XOR2X1 U90 ( .A(n71), .B(n69), .Y(DIFF[9]) );
  NOR2X1 U91 ( .A(n69), .B(n71), .Y(n68) );
  XOR2X1 U94 ( .A(n75), .B(B[8]), .Y(DIFF[8]) );
  NOR2X1 U96 ( .A(n78), .B(n73), .Y(n72) );
  NAND2X1 U97 ( .A(n76), .B(n74), .Y(n73) );
  XNOR2X1 U99 ( .A(n77), .B(B[7]), .Y(DIFF[7]) );
  NAND2X1 U100 ( .A(n76), .B(n77), .Y(n75) );
  XNOR2X1 U102 ( .A(n80), .B(B[6]), .Y(DIFF[6]) );
  NAND2X1 U104 ( .A(n79), .B(n82), .Y(n78) );
  NOR2X1 U105 ( .A(B[5]), .B(B[6]), .Y(n79) );
  XOR2X1 U106 ( .A(n81), .B(B[5]), .Y(DIFF[5]) );
  NOR2X1 U107 ( .A(B[5]), .B(n81), .Y(n80) );
  XOR2X1 U108 ( .A(n85), .B(B[4]), .Y(DIFF[4]) );
  NOR2X1 U110 ( .A(n88), .B(n83), .Y(n82) );
  NAND2X1 U111 ( .A(n86), .B(n84), .Y(n83) );
  XNOR2X1 U113 ( .A(B[3]), .B(n87), .Y(DIFF[3]) );
  NAND2X1 U114 ( .A(n86), .B(n87), .Y(n85) );
  XNOR2X1 U116 ( .A(B[2]), .B(n90), .Y(DIFF[2]) );
  NAND2X1 U118 ( .A(n89), .B(n90), .Y(n88) );
  XOR2X1 U120 ( .A(B[1]), .B(\B[0] ), .Y(DIFF[1]) );
  NOR2X1 U121 ( .A(\B[0] ), .B(B[1]), .Y(n90) );
  INVX2 U125 ( .A(n53), .Y(n193) );
  INVX4 U126 ( .A(n27), .Y(n26) );
  INVX1 U127 ( .A(B[25]), .Y(n19) );
  OR2X2 U128 ( .A(B[29]), .B(B[30]), .Y(n194) );
  INVX1 U129 ( .A(n63), .Y(n62) );
  INVX1 U130 ( .A(B[19]), .Y(n37) );
  OR2X1 U131 ( .A(n69), .B(B[10]), .Y(n66) );
  INVX1 U132 ( .A(n47), .Y(n48) );
  INVX1 U133 ( .A(n33), .Y(n34) );
  INVX1 U134 ( .A(n22), .Y(n21) );
  INVX1 U135 ( .A(n13), .Y(n14) );
  INVX2 U136 ( .A(B[2]), .Y(n89) );
  INVX2 U137 ( .A(n88), .Y(n87) );
  INVX2 U138 ( .A(B[3]), .Y(n86) );
  INVX2 U139 ( .A(B[4]), .Y(n84) );
  INVX2 U140 ( .A(n82), .Y(n81) );
  INVX2 U141 ( .A(B[28]), .Y(n8) );
  INVX2 U142 ( .A(n78), .Y(n77) );
  INVX2 U143 ( .A(B[7]), .Y(n76) );
  INVX2 U144 ( .A(B[8]), .Y(n74) );
  INVX2 U145 ( .A(n72), .Y(n71) );
  INVX2 U146 ( .A(B[12]), .Y(n61) );
  INVX2 U147 ( .A(B[14]), .Y(n57) );
  INVX2 U148 ( .A(n55), .Y(n54) );
  INVX2 U149 ( .A(n52), .Y(n53) );
  INVX2 U150 ( .A(B[16]), .Y(n50) );
  INVX2 U151 ( .A(B[17]), .Y(n45) );
  INVX2 U152 ( .A(B[18]), .Y(n42) );
  INVX2 U153 ( .A(n39), .Y(n38) );
  INVX2 U154 ( .A(B[27]), .Y(n11) );
endmodule


module poly5_DW_mult_uns_57 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n289, n292, n295, n298, n301, n304, n307, n310, n313, n316, n319,
         n322, n325, n328, n330, n333, n433, n437, n439, n441, n443, n445,
         n447, n449, n451, n453, n455, n457, n459, n461, n463, n465, n467,
         n469, n471, n473, n475, n477, n479, n481, n483, n485, n487, n489,
         n491, n493, n495, n497, n499, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n547, n548, n549, n551, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n569, n571, n572, n573, n574, n578, n580, n581, n582, n583,
         n584, n585, n586, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n617, n618, n619, n620, n621,
         n622, n623, n624, n627, n628, n629, n630, n631, n633, n634, n635,
         n636, n637, n638, n639, n640, n643, n644, n645, n646, n647, n648,
         n649, n651, n652, n653, n654, n655, n656, n657, n658, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n682, n683, n684, n685, n686, n687, n690,
         n691, n692, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n704, n706, n707, n708, n709, n713, n715, n716, n717, n718, n719,
         n720, n724, n726, n727, n728, n729, n731, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n748, n749, n750,
         n751, n752, n753, n756, n757, n758, n760, n761, n762, n764, n765,
         n766, n767, n768, n769, n770, n771, n773, n775, n776, n777, n778,
         n780, n783, n784, n785, n786, n788, n790, n791, n793, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n810, n812, n813, n815, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n833, n835,
         n836, n837, n838, n839, n841, n843, n844, n845, n846, n847, n849,
         n851, n852, n853, n854, n856, n858, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n879,
         n880, n881, n882, n883, n884, n886, n889, n890, n893, n894, n895,
         n897, n899, n901, n903, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2764, n2765, n2766, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n3179, n3178, n3177, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176;
  assign n289 = b[1];
  assign n292 = b[3];
  assign n295 = b[5];
  assign n298 = b[7];
  assign n301 = b[9];
  assign n304 = b[11];
  assign n307 = b[13];
  assign n310 = b[15];
  assign n313 = b[17];
  assign n316 = b[19];
  assign n319 = b[21];
  assign n322 = b[23];
  assign n325 = b[25];
  assign n328 = b[27];
  assign n330 = b[29];
  assign n333 = b[31];
  assign n433 = a[0];
  assign n437 = a[1];
  assign n439 = a[2];
  assign n441 = a[3];
  assign n443 = a[4];
  assign n445 = a[5];
  assign n447 = a[6];
  assign n449 = a[7];
  assign n451 = a[8];
  assign n453 = a[9];
  assign n455 = a[10];
  assign n457 = a[11];
  assign n459 = a[12];
  assign n461 = a[13];
  assign n463 = a[14];
  assign n465 = a[15];
  assign n467 = a[16];
  assign n469 = a[17];
  assign n471 = a[18];
  assign n473 = a[19];
  assign n475 = a[20];
  assign n477 = a[21];
  assign n479 = a[22];
  assign n481 = a[23];
  assign n483 = a[24];
  assign n485 = a[25];
  assign n487 = a[26];
  assign n489 = a[27];
  assign n491 = a[28];
  assign n493 = a[29];
  assign n495 = a[30];
  assign n497 = a[31];

  XNOR2X1 U294 ( .A(n554), .B(n501), .Y(product[46]) );
  OAI21X1 U295 ( .A(n548), .B(n3020), .C(n549), .Y(n547) );
  NAND2X1 U296 ( .A(n2932), .B(n557), .Y(n548) );
  AOI21X1 U297 ( .A(n2932), .B(n558), .C(n551), .Y(n549) );
  NAND2X1 U300 ( .A(n553), .B(n2932), .Y(n501) );
  NAND2X1 U303 ( .A(n932), .B(n913), .Y(n553) );
  XNOR2X1 U304 ( .A(n561), .B(n502), .Y(product[45]) );
  OAI21X1 U305 ( .A(n555), .B(n3020), .C(n556), .Y(n554) );
  NOR2X1 U308 ( .A(n559), .B(n562), .Y(n557) );
  OAI21X1 U309 ( .A(n559), .B(n563), .C(n560), .Y(n558) );
  NAND2X1 U310 ( .A(n560), .B(n858), .Y(n502) );
  NOR2X1 U312 ( .A(n952), .B(n933), .Y(n559) );
  NAND2X1 U313 ( .A(n952), .B(n933), .Y(n560) );
  XNOR2X1 U314 ( .A(n572), .B(n503), .Y(n3177) );
  OAI21X1 U315 ( .A(n562), .B(n3020), .C(n563), .Y(n561) );
  NAND2X1 U316 ( .A(n593), .B(n564), .Y(n562) );
  AOI21X1 U317 ( .A(n594), .B(n564), .C(n565), .Y(n563) );
  NOR2X1 U318 ( .A(n586), .B(n566), .Y(n564) );
  OAI21X1 U319 ( .A(n589), .B(n566), .C(n567), .Y(n565) );
  NAND2X1 U320 ( .A(n2983), .B(n2979), .Y(n566) );
  AOI21X1 U321 ( .A(n578), .B(n2983), .C(n569), .Y(n567) );
  NAND2X1 U324 ( .A(n571), .B(n2983), .Y(n503) );
  NAND2X1 U327 ( .A(n974), .B(n953), .Y(n571) );
  XNOR2X1 U328 ( .A(n581), .B(n504), .Y(product[43]) );
  OAI21X1 U329 ( .A(n573), .B(n3020), .C(n574), .Y(n572) );
  NAND2X1 U330 ( .A(n2979), .B(n584), .Y(n573) );
  AOI21X1 U331 ( .A(n2979), .B(n585), .C(n578), .Y(n574) );
  NAND2X1 U336 ( .A(n580), .B(n2979), .Y(n504) );
  NAND2X1 U339 ( .A(n996), .B(n975), .Y(n580) );
  XNOR2X1 U340 ( .A(n590), .B(n505), .Y(product[42]) );
  OAI21X1 U341 ( .A(n582), .B(n3019), .C(n583), .Y(n581) );
  NOR2X1 U344 ( .A(n586), .B(n591), .Y(n584) );
  OAI21X1 U345 ( .A(n586), .B(n592), .C(n589), .Y(n585) );
  NAND2X1 U348 ( .A(n589), .B(n861), .Y(n505) );
  NOR2X1 U350 ( .A(n1020), .B(n997), .Y(n586) );
  NAND2X1 U351 ( .A(n1020), .B(n997), .Y(n589) );
  XNOR2X1 U352 ( .A(n597), .B(n506), .Y(product[41]) );
  OAI21X1 U353 ( .A(n591), .B(n3019), .C(n592), .Y(n590) );
  NOR2X1 U356 ( .A(n595), .B(n598), .Y(n593) );
  OAI21X1 U357 ( .A(n599), .B(n595), .C(n596), .Y(n594) );
  NAND2X1 U358 ( .A(n596), .B(n862), .Y(n506) );
  NOR2X1 U360 ( .A(n1044), .B(n1021), .Y(n595) );
  NAND2X1 U361 ( .A(n1044), .B(n1021), .Y(n596) );
  XOR2X1 U362 ( .A(n3020), .B(n507), .Y(product[40]) );
  OAI21X1 U363 ( .A(n598), .B(n3019), .C(n599), .Y(n597) );
  NAND2X1 U364 ( .A(n599), .B(n863), .Y(n507) );
  NOR2X1 U366 ( .A(n1070), .B(n1045), .Y(n598) );
  NAND2X1 U367 ( .A(n1070), .B(n1045), .Y(n599) );
  XNOR2X1 U368 ( .A(n609), .B(n508), .Y(product[39]) );
  AOI21X1 U369 ( .A(n669), .B(n601), .C(n602), .Y(n499) );
  NOR2X1 U370 ( .A(n603), .B(n637), .Y(n601) );
  OAI21X1 U371 ( .A(n603), .B(n638), .C(n604), .Y(n602) );
  NAND2X1 U372 ( .A(n605), .B(n621), .Y(n603) );
  AOI21X1 U373 ( .A(n605), .B(n622), .C(n606), .Y(n604) );
  NOR2X1 U374 ( .A(n607), .B(n614), .Y(n605) );
  OAI21X1 U375 ( .A(n617), .B(n607), .C(n608), .Y(n606) );
  NAND2X1 U376 ( .A(n608), .B(n864), .Y(n508) );
  NOR2X1 U378 ( .A(n1096), .B(n1071), .Y(n607) );
  NAND2X1 U379 ( .A(n1096), .B(n1071), .Y(n608) );
  XNOR2X1 U380 ( .A(n618), .B(n509), .Y(product[38]) );
  OAI21X1 U381 ( .A(n3017), .B(n610), .C(n611), .Y(n609) );
  NAND2X1 U382 ( .A(n639), .B(n612), .Y(n610) );
  AOI21X1 U383 ( .A(n640), .B(n612), .C(n613), .Y(n611) );
  NOR2X1 U384 ( .A(n614), .B(n623), .Y(n612) );
  OAI21X1 U385 ( .A(n614), .B(n624), .C(n617), .Y(n613) );
  NAND2X1 U388 ( .A(n617), .B(n865), .Y(n509) );
  NOR2X1 U390 ( .A(n1124), .B(n1097), .Y(n614) );
  NAND2X1 U391 ( .A(n1124), .B(n1097), .Y(n617) );
  XNOR2X1 U392 ( .A(n629), .B(n510), .Y(product[37]) );
  OAI21X1 U393 ( .A(n3018), .B(n619), .C(n620), .Y(n618) );
  NAND2X1 U394 ( .A(n621), .B(n639), .Y(n619) );
  AOI21X1 U395 ( .A(n621), .B(n640), .C(n622), .Y(n620) );
  NOR2X1 U400 ( .A(n627), .B(n634), .Y(n621) );
  OAI21X1 U401 ( .A(n635), .B(n627), .C(n628), .Y(n622) );
  NAND2X1 U402 ( .A(n628), .B(n866), .Y(n510) );
  NOR2X1 U404 ( .A(n1152), .B(n1125), .Y(n627) );
  NAND2X1 U405 ( .A(n1152), .B(n1125), .Y(n628) );
  XNOR2X1 U406 ( .A(n636), .B(n511), .Y(product[36]) );
  OAI21X1 U407 ( .A(n3017), .B(n630), .C(n631), .Y(n629) );
  NAND2X1 U408 ( .A(n867), .B(n639), .Y(n630) );
  AOI21X1 U409 ( .A(n867), .B(n640), .C(n633), .Y(n631) );
  NAND2X1 U412 ( .A(n635), .B(n867), .Y(n511) );
  NOR2X1 U414 ( .A(n1182), .B(n1153), .Y(n634) );
  NAND2X1 U415 ( .A(n1182), .B(n1153), .Y(n635) );
  XNOR2X1 U416 ( .A(n647), .B(n512), .Y(product[35]) );
  OAI21X1 U417 ( .A(n637), .B(n3018), .C(n638), .Y(n636) );
  NAND2X1 U422 ( .A(n657), .B(n643), .Y(n637) );
  AOI21X1 U423 ( .A(n658), .B(n643), .C(n644), .Y(n638) );
  NOR2X1 U424 ( .A(n645), .B(n652), .Y(n643) );
  OAI21X1 U425 ( .A(n653), .B(n645), .C(n646), .Y(n644) );
  NAND2X1 U426 ( .A(n646), .B(n868), .Y(n512) );
  NOR2X1 U428 ( .A(n1212), .B(n1183), .Y(n645) );
  NAND2X1 U429 ( .A(n1212), .B(n1183), .Y(n646) );
  XNOR2X1 U430 ( .A(n654), .B(n513), .Y(product[34]) );
  OAI21X1 U431 ( .A(n648), .B(n3017), .C(n649), .Y(n647) );
  NAND2X1 U432 ( .A(n869), .B(n657), .Y(n648) );
  AOI21X1 U433 ( .A(n869), .B(n658), .C(n651), .Y(n649) );
  NAND2X1 U436 ( .A(n653), .B(n869), .Y(n513) );
  NOR2X1 U438 ( .A(n1244), .B(n1213), .Y(n652) );
  NAND2X1 U439 ( .A(n1244), .B(n1213), .Y(n653) );
  XNOR2X1 U440 ( .A(n665), .B(n514), .Y(product[33]) );
  OAI21X1 U441 ( .A(n655), .B(n3018), .C(n656), .Y(n654) );
  NOR2X1 U448 ( .A(n666), .B(n663), .Y(n657) );
  OAI21X1 U449 ( .A(n667), .B(n663), .C(n664), .Y(n658) );
  NAND2X1 U450 ( .A(n664), .B(n870), .Y(n514) );
  NOR2X1 U452 ( .A(n1275), .B(n1245), .Y(n663) );
  NAND2X1 U453 ( .A(n1275), .B(n1245), .Y(n664) );
  XOR2X1 U454 ( .A(n3017), .B(n515), .Y(product[32]) );
  OAI21X1 U455 ( .A(n666), .B(n3017), .C(n667), .Y(n665) );
  NAND2X1 U456 ( .A(n667), .B(n871), .Y(n515) );
  NOR2X1 U458 ( .A(n1305), .B(n1276), .Y(n666) );
  NAND2X1 U459 ( .A(n1305), .B(n1276), .Y(n667) );
  XOR2X1 U460 ( .A(n676), .B(n516), .Y(product[31]) );
  OAI21X1 U462 ( .A(n670), .B(n698), .C(n671), .Y(n669) );
  NAND2X1 U463 ( .A(n684), .B(n672), .Y(n670) );
  AOI21X1 U464 ( .A(n685), .B(n672), .C(n673), .Y(n671) );
  NOR2X1 U465 ( .A(n679), .B(n674), .Y(n672) );
  OAI21X1 U466 ( .A(n682), .B(n674), .C(n675), .Y(n673) );
  NAND2X1 U467 ( .A(n675), .B(n872), .Y(n516) );
  NOR2X1 U469 ( .A(n1335), .B(n1306), .Y(n674) );
  NAND2X1 U470 ( .A(n1335), .B(n1306), .Y(n675) );
  XOR2X1 U471 ( .A(n683), .B(n517), .Y(product[30]) );
  AOI21X1 U472 ( .A(n677), .B(n697), .C(n678), .Y(n676) );
  NOR2X1 U473 ( .A(n679), .B(n686), .Y(n677) );
  OAI21X1 U474 ( .A(n679), .B(n687), .C(n682), .Y(n678) );
  NAND2X1 U477 ( .A(n682), .B(n873), .Y(n517) );
  NOR2X1 U479 ( .A(n1363), .B(n1336), .Y(n679) );
  NAND2X1 U480 ( .A(n1363), .B(n1336), .Y(n682) );
  AOI21X1 U482 ( .A(n684), .B(n697), .C(n685), .Y(n683) );
  NOR2X1 U487 ( .A(n695), .B(n690), .Y(n684) );
  OAI21X1 U488 ( .A(n696), .B(n690), .C(n691), .Y(n685) );
  NOR2X1 U491 ( .A(n1391), .B(n1364), .Y(n690) );
  NAND2X1 U492 ( .A(n1391), .B(n1364), .Y(n691) );
  XNOR2X1 U493 ( .A(n697), .B(n519), .Y(n3178) );
  AOI21X1 U494 ( .A(n875), .B(n3022), .C(n694), .Y(n692) );
  NAND2X1 U497 ( .A(n696), .B(n875), .Y(n519) );
  NOR2X1 U499 ( .A(n1417), .B(n1392), .Y(n695) );
  NAND2X1 U500 ( .A(n1417), .B(n1392), .Y(n696) );
  XNOR2X1 U501 ( .A(n707), .B(n520), .Y(product[27]) );
  AOI21X1 U503 ( .A(n735), .B(n699), .C(n700), .Y(n698) );
  NOR2X1 U504 ( .A(n717), .B(n701), .Y(n699) );
  OAI21X1 U505 ( .A(n718), .B(n701), .C(n702), .Y(n700) );
  NAND2X1 U506 ( .A(n2980), .B(n2981), .Y(n701) );
  AOI21X1 U507 ( .A(n713), .B(n2981), .C(n704), .Y(n702) );
  NAND2X1 U510 ( .A(n706), .B(n2981), .Y(n520) );
  NAND2X1 U513 ( .A(n1443), .B(n1418), .Y(n706) );
  XNOR2X1 U514 ( .A(n716), .B(n521), .Y(product[26]) );
  OAI21X1 U515 ( .A(n708), .B(n734), .C(n709), .Y(n707) );
  NAND2X1 U516 ( .A(n2980), .B(n719), .Y(n708) );
  AOI21X1 U517 ( .A(n2980), .B(n720), .C(n713), .Y(n709) );
  NAND2X1 U522 ( .A(n715), .B(n2980), .Y(n521) );
  NAND2X1 U525 ( .A(n1467), .B(n1444), .Y(n715) );
  OAI21X1 U527 ( .A(n717), .B(n734), .C(n718), .Y(n716) );
  NAND2X1 U532 ( .A(n879), .B(n2982), .Y(n717) );
  AOI21X1 U533 ( .A(n731), .B(n2982), .C(n724), .Y(n718) );
  NAND2X1 U536 ( .A(n726), .B(n2982), .Y(n522) );
  NAND2X1 U539 ( .A(n1491), .B(n1468), .Y(n726) );
  XOR2X1 U540 ( .A(n734), .B(n523), .Y(product[24]) );
  OAI21X1 U541 ( .A(n728), .B(n734), .C(n729), .Y(n727) );
  NAND2X1 U546 ( .A(n729), .B(n879), .Y(n523) );
  NOR2X1 U548 ( .A(n1513), .B(n1492), .Y(n728) );
  NAND2X1 U549 ( .A(n1513), .B(n1492), .Y(n729) );
  XOR2X1 U550 ( .A(n742), .B(n524), .Y(product[23]) );
  OAI21X1 U552 ( .A(n764), .B(n736), .C(n737), .Y(n735) );
  NAND2X1 U553 ( .A(n750), .B(n738), .Y(n736) );
  AOI21X1 U554 ( .A(n751), .B(n738), .C(n739), .Y(n737) );
  NOR2X1 U555 ( .A(n745), .B(n740), .Y(n738) );
  OAI21X1 U556 ( .A(n748), .B(n740), .C(n741), .Y(n739) );
  NAND2X1 U557 ( .A(n741), .B(n880), .Y(n524) );
  NOR2X1 U559 ( .A(n1535), .B(n1514), .Y(n740) );
  NAND2X1 U560 ( .A(n1535), .B(n1514), .Y(n741) );
  XOR2X1 U561 ( .A(n749), .B(n525), .Y(n3179) );
  AOI21X1 U562 ( .A(n2942), .B(n743), .C(n744), .Y(n742) );
  NOR2X1 U563 ( .A(n745), .B(n752), .Y(n743) );
  OAI21X1 U564 ( .A(n745), .B(n753), .C(n748), .Y(n744) );
  NAND2X1 U567 ( .A(n748), .B(n881), .Y(n525) );
  NOR2X1 U569 ( .A(n1555), .B(n1536), .Y(n745) );
  NAND2X1 U570 ( .A(n1555), .B(n1536), .Y(n748) );
  XOR2X1 U571 ( .A(n758), .B(n526), .Y(product[21]) );
  AOI21X1 U572 ( .A(n750), .B(n2942), .C(n751), .Y(n749) );
  NOR2X1 U577 ( .A(n761), .B(n756), .Y(n750) );
  OAI21X1 U578 ( .A(n762), .B(n756), .C(n757), .Y(n751) );
  NAND2X1 U579 ( .A(n757), .B(n882), .Y(n526) );
  NOR2X1 U581 ( .A(n1575), .B(n1556), .Y(n756) );
  NAND2X1 U582 ( .A(n1575), .B(n1556), .Y(n757) );
  XNOR2X1 U583 ( .A(n2942), .B(n527), .Y(product[20]) );
  AOI21X1 U584 ( .A(n883), .B(n2942), .C(n760), .Y(n758) );
  NAND2X1 U587 ( .A(n762), .B(n883), .Y(n527) );
  NOR2X1 U589 ( .A(n1593), .B(n1576), .Y(n761) );
  NAND2X1 U590 ( .A(n1593), .B(n1576), .Y(n762) );
  XNOR2X1 U591 ( .A(n769), .B(n528), .Y(product[19]) );
  AOI21X1 U593 ( .A(n784), .B(n765), .C(n766), .Y(n764) );
  NOR2X1 U594 ( .A(n767), .B(n770), .Y(n765) );
  OAI21X1 U595 ( .A(n767), .B(n771), .C(n768), .Y(n766) );
  NAND2X1 U596 ( .A(n768), .B(n884), .Y(n528) );
  NOR2X1 U598 ( .A(n1611), .B(n1594), .Y(n767) );
  NAND2X1 U599 ( .A(n1611), .B(n1594), .Y(n768) );
  XNOR2X1 U600 ( .A(n776), .B(n529), .Y(product[18]) );
  OAI21X1 U601 ( .A(n770), .B(n783), .C(n771), .Y(n769) );
  NAND2X1 U602 ( .A(n886), .B(n2985), .Y(n770) );
  AOI21X1 U603 ( .A(n780), .B(n2985), .C(n773), .Y(n771) );
  NAND2X1 U606 ( .A(n775), .B(n2985), .Y(n529) );
  NAND2X1 U609 ( .A(n1627), .B(n1612), .Y(n775) );
  XOR2X1 U610 ( .A(n783), .B(n530), .Y(product[17]) );
  OAI21X1 U611 ( .A(n777), .B(n783), .C(n778), .Y(n776) );
  NAND2X1 U616 ( .A(n778), .B(n886), .Y(n530) );
  NOR2X1 U618 ( .A(n1643), .B(n1628), .Y(n777) );
  NAND2X1 U619 ( .A(n1643), .B(n1628), .Y(n778) );
  OAI21X1 U622 ( .A(n785), .B(n797), .C(n786), .Y(n784) );
  NAND2X1 U623 ( .A(n2987), .B(n2986), .Y(n785) );
  AOI21X1 U624 ( .A(n793), .B(n2986), .C(n788), .Y(n786) );
  NAND2X1 U630 ( .A(n1657), .B(n1644), .Y(n790) );
  XNOR2X1 U631 ( .A(n796), .B(n532), .Y(product[15]) );
  AOI21X1 U632 ( .A(n2987), .B(n796), .C(n793), .Y(n791) );
  NAND2X1 U635 ( .A(n795), .B(n2987), .Y(n532) );
  NAND2X1 U638 ( .A(n1671), .B(n1658), .Y(n795) );
  XNOR2X1 U639 ( .A(n802), .B(n533), .Y(product[14]) );
  AOI21X1 U641 ( .A(n806), .B(n798), .C(n799), .Y(n797) );
  NOR2X1 U642 ( .A(n803), .B(n800), .Y(n798) );
  OAI21X1 U643 ( .A(n804), .B(n800), .C(n801), .Y(n799) );
  NAND2X1 U644 ( .A(n801), .B(n889), .Y(n533) );
  NOR2X1 U646 ( .A(n1683), .B(n1672), .Y(n800) );
  NAND2X1 U647 ( .A(n1683), .B(n1672), .Y(n801) );
  XOR2X1 U648 ( .A(n805), .B(n534), .Y(product[13]) );
  OAI21X1 U649 ( .A(n803), .B(n805), .C(n804), .Y(n802) );
  NAND2X1 U650 ( .A(n804), .B(n890), .Y(n534) );
  NOR2X1 U652 ( .A(n1695), .B(n1684), .Y(n803) );
  NAND2X1 U653 ( .A(n1695), .B(n1684), .Y(n804) );
  XOR2X1 U654 ( .A(n813), .B(n535), .Y(product[12]) );
  OAI21X1 U656 ( .A(n807), .B(n819), .C(n808), .Y(n806) );
  NAND2X1 U657 ( .A(n2989), .B(n2988), .Y(n807) );
  AOI21X1 U658 ( .A(n815), .B(n2988), .C(n810), .Y(n808) );
  NAND2X1 U661 ( .A(n812), .B(n2988), .Y(n535) );
  NAND2X1 U664 ( .A(n1705), .B(n1696), .Y(n812) );
  XNOR2X1 U665 ( .A(n818), .B(n536), .Y(product[11]) );
  AOI21X1 U666 ( .A(n2989), .B(n818), .C(n815), .Y(n813) );
  NAND2X1 U669 ( .A(n817), .B(n2989), .Y(n536) );
  NAND2X1 U672 ( .A(n1715), .B(n1706), .Y(n817) );
  XNOR2X1 U673 ( .A(n824), .B(n537), .Y(product[10]) );
  AOI21X1 U675 ( .A(n828), .B(n820), .C(n821), .Y(n819) );
  NOR2X1 U676 ( .A(n825), .B(n822), .Y(n820) );
  OAI21X1 U677 ( .A(n826), .B(n822), .C(n823), .Y(n821) );
  NAND2X1 U678 ( .A(n823), .B(n893), .Y(n537) );
  NOR2X1 U680 ( .A(n1723), .B(n1716), .Y(n822) );
  NAND2X1 U681 ( .A(n1723), .B(n1716), .Y(n823) );
  XOR2X1 U682 ( .A(n827), .B(n538), .Y(product[9]) );
  OAI21X1 U683 ( .A(n825), .B(n827), .C(n826), .Y(n824) );
  NAND2X1 U684 ( .A(n826), .B(n894), .Y(n538) );
  NOR2X1 U686 ( .A(n1731), .B(n1724), .Y(n825) );
  NAND2X1 U687 ( .A(n1731), .B(n1724), .Y(n826) );
  XOR2X1 U688 ( .A(n831), .B(n539), .Y(product[8]) );
  OAI21X1 U690 ( .A(n829), .B(n831), .C(n830), .Y(n828) );
  NAND2X1 U691 ( .A(n830), .B(n895), .Y(n539) );
  NOR2X1 U693 ( .A(n1737), .B(n1732), .Y(n829) );
  NAND2X1 U694 ( .A(n1737), .B(n1732), .Y(n830) );
  XNOR2X1 U695 ( .A(n836), .B(n540), .Y(product[7]) );
  AOI21X1 U696 ( .A(n2991), .B(n836), .C(n833), .Y(n831) );
  NAND2X1 U699 ( .A(n835), .B(n2991), .Y(n540) );
  NAND2X1 U702 ( .A(n1743), .B(n1738), .Y(n835) );
  XOR2X1 U703 ( .A(n541), .B(n839), .Y(product[6]) );
  OAI21X1 U704 ( .A(n839), .B(n837), .C(n838), .Y(n836) );
  NAND2X1 U705 ( .A(n838), .B(n897), .Y(n541) );
  NOR2X1 U707 ( .A(n1747), .B(n1744), .Y(n837) );
  NAND2X1 U708 ( .A(n1747), .B(n1744), .Y(n838) );
  XNOR2X1 U709 ( .A(n542), .B(n844), .Y(product[5]) );
  AOI21X1 U710 ( .A(n844), .B(n2990), .C(n841), .Y(n839) );
  NAND2X1 U713 ( .A(n843), .B(n2990), .Y(n542) );
  NAND2X1 U716 ( .A(n1751), .B(n1748), .Y(n843) );
  XOR2X1 U717 ( .A(n543), .B(n847), .Y(product[4]) );
  OAI21X1 U718 ( .A(n847), .B(n845), .C(n846), .Y(n844) );
  NAND2X1 U719 ( .A(n846), .B(n899), .Y(n543) );
  NOR2X1 U721 ( .A(n1753), .B(n1752), .Y(n845) );
  NAND2X1 U722 ( .A(n1753), .B(n1752), .Y(n846) );
  XNOR2X1 U723 ( .A(n544), .B(n852), .Y(product[3]) );
  AOI21X1 U724 ( .A(n852), .B(n3021), .C(n849), .Y(n847) );
  NAND2X1 U727 ( .A(n851), .B(n3021), .Y(n544) );
  NAND2X1 U730 ( .A(n1769), .B(n1754), .Y(n851) );
  XOR2X1 U731 ( .A(n545), .B(n856), .Y(product[2]) );
  OAI21X1 U732 ( .A(n856), .B(n853), .C(n854), .Y(n852) );
  NAND2X1 U733 ( .A(n854), .B(n901), .Y(n545) );
  NOR2X1 U735 ( .A(n2218), .B(n2249), .Y(n853) );
  NAND2X1 U736 ( .A(n2218), .B(n2249), .Y(n854) );
  NAND2X1 U741 ( .A(n2250), .B(n1770), .Y(n856) );
  FAX1 U742 ( .A(n917), .B(n934), .C(n915), .YC(n912), .YS(n913) );
  FAX1 U743 ( .A(n938), .B(n919), .C(n936), .YC(n914), .YS(n915) );
  FAX1 U744 ( .A(n923), .B(n940), .C(n921), .YC(n916), .YS(n917) );
  FAX1 U745 ( .A(n944), .B(n925), .C(n942), .YC(n918), .YS(n919) );
  FAX1 U746 ( .A(n929), .B(n927), .C(n946), .YC(n920), .YS(n921) );
  FAX1 U747 ( .A(n1892), .B(n1920), .C(n948), .YC(n922), .YS(n923) );
  FAX1 U748 ( .A(n950), .B(n1866), .C(n1950), .YC(n924), .YS(n925) );
  FAX1 U749 ( .A(n1782), .B(n1820), .C(n1842), .YC(n926), .YS(n927) );
  FAX1 U750 ( .A(n931), .B(n1982), .C(n1800), .YC(n928), .YS(n929) );
  FAX1 U752 ( .A(n937), .B(n954), .C(n935), .YC(n932), .YS(n933) );
  FAX1 U753 ( .A(n958), .B(n939), .C(n956), .YC(n934), .YS(n935) );
  FAX1 U754 ( .A(n943), .B(n960), .C(n941), .YC(n936), .YS(n937) );
  FAX1 U755 ( .A(n947), .B(n945), .C(n962), .YC(n938), .YS(n939) );
  FAX1 U756 ( .A(n949), .B(n966), .C(n964), .YC(n940), .YS(n941) );
  FAX1 U757 ( .A(n1893), .B(n970), .C(n968), .YC(n942), .YS(n943) );
  FAX1 U758 ( .A(n1983), .B(n1921), .C(n951), .YC(n944), .YS(n945) );
  FAX1 U759 ( .A(n1843), .B(n1867), .C(n1951), .YC(n946), .YS(n947) );
  FAX1 U760 ( .A(n1801), .B(n1821), .C(n1783), .YC(n948), .YS(n949) );
  FAX1 U761 ( .A(n2015), .B(n972), .C(n1772), .YC(n950), .YS(n951) );
  FAX1 U762 ( .A(n957), .B(n976), .C(n955), .YC(n952), .YS(n953) );
  FAX1 U763 ( .A(n980), .B(n959), .C(n978), .YC(n954), .YS(n955) );
  FAX1 U764 ( .A(n963), .B(n982), .C(n961), .YC(n956), .YS(n957) );
  FAX1 U765 ( .A(n986), .B(n965), .C(n984), .YC(n958), .YS(n959) );
  FAX1 U766 ( .A(n969), .B(n988), .C(n967), .YC(n960), .YS(n961) );
  FAX1 U767 ( .A(n992), .B(n971), .C(n990), .YC(n962), .YS(n963) );
  FAX1 U768 ( .A(n1984), .B(n1922), .C(n1952), .YC(n964), .YS(n965) );
  FAX1 U769 ( .A(n1868), .B(n994), .C(n1894), .YC(n966), .YS(n967) );
  FAX1 U770 ( .A(n1802), .B(n1784), .C(n1844), .YC(n968), .YS(n969) );
  FAX1 U771 ( .A(n973), .B(n2016), .C(n1822), .YC(n970), .YS(n971) );
  FAX1 U773 ( .A(n979), .B(n998), .C(n977), .YC(n974), .YS(n975) );
  FAX1 U774 ( .A(n1002), .B(n981), .C(n1000), .YC(n976), .YS(n977) );
  FAX1 U775 ( .A(n985), .B(n1004), .C(n983), .YC(n978), .YS(n979) );
  FAX1 U776 ( .A(n1008), .B(n987), .C(n1006), .YC(n980), .YS(n981) );
  FAX1 U777 ( .A(n991), .B(n1010), .C(n989), .YC(n982), .YS(n983) );
  FAX1 U778 ( .A(n1014), .B(n993), .C(n1012), .YC(n984), .YS(n985) );
  FAX1 U779 ( .A(n1953), .B(n1923), .C(n1016), .YC(n986), .YS(n987) );
  FAX1 U780 ( .A(n1985), .B(n2017), .C(n995), .YC(n988), .YS(n989) );
  FAX1 U781 ( .A(n1785), .B(n1869), .C(n1895), .YC(n990), .YS(n991) );
  FAX1 U782 ( .A(n1823), .B(n1845), .C(n1803), .YC(n992), .YS(n993) );
  FAX1 U783 ( .A(n2049), .B(n1018), .C(n1773), .YC(n994), .YS(n995) );
  FAX1 U784 ( .A(n1001), .B(n1022), .C(n999), .YC(n996), .YS(n997) );
  FAX1 U785 ( .A(n1026), .B(n1003), .C(n1024), .YC(n998), .YS(n999) );
  FAX1 U786 ( .A(n1007), .B(n1028), .C(n1005), .YC(n1000), .YS(n1001) );
  FAX1 U787 ( .A(n1032), .B(n1009), .C(n1030), .YC(n1002), .YS(n1003) );
  FAX1 U788 ( .A(n1036), .B(n1034), .C(n1011), .YC(n1004), .YS(n1005) );
  FAX1 U789 ( .A(n1017), .B(n1015), .C(n1013), .YC(n1006), .YS(n1007) );
  FAX1 U790 ( .A(n1954), .B(n1040), .C(n1038), .YC(n1008), .YS(n1009) );
  FAX1 U791 ( .A(n1924), .B(n2018), .C(n1986), .YC(n1010), .YS(n1011) );
  FAX1 U792 ( .A(n1870), .B(n1896), .C(n1042), .YC(n1012), .YS(n1013) );
  FAX1 U793 ( .A(n1846), .B(n1804), .C(n1786), .YC(n1014), .YS(n1015) );
  FAX1 U794 ( .A(n1019), .B(n2050), .C(n1824), .YC(n1016), .YS(n1017) );
  FAX1 U796 ( .A(n1025), .B(n1046), .C(n1023), .YC(n1020), .YS(n1021) );
  FAX1 U797 ( .A(n1050), .B(n1027), .C(n1048), .YC(n1022), .YS(n1023) );
  FAX1 U798 ( .A(n1031), .B(n1052), .C(n1029), .YC(n1024), .YS(n1025) );
  FAX1 U799 ( .A(n1056), .B(n1033), .C(n1054), .YC(n1026), .YS(n1027) );
  FAX1 U800 ( .A(n1058), .B(n1037), .C(n1035), .YC(n1028), .YS(n1029) );
  FAX1 U801 ( .A(n1041), .B(n1039), .C(n1060), .YC(n1030), .YS(n1031) );
  FAX1 U802 ( .A(n1066), .B(n1064), .C(n1062), .YC(n1032), .YS(n1033) );
  FAX1 U803 ( .A(n1987), .B(n1955), .C(n1043), .YC(n1034), .YS(n1035) );
  FAX1 U804 ( .A(n1925), .B(n2019), .C(n2051), .YC(n1036), .YS(n1037) );
  FAX1 U805 ( .A(n1805), .B(n1825), .C(n1897), .YC(n1038), .YS(n1039) );
  FAX1 U806 ( .A(n1847), .B(n1871), .C(n1787), .YC(n1040), .YS(n1041) );
  FAX1 U807 ( .A(n2083), .B(n1068), .C(n1774), .YC(n1042), .YS(n1043) );
  FAX1 U808 ( .A(n1049), .B(n1072), .C(n1047), .YC(n1044), .YS(n1045) );
  FAX1 U809 ( .A(n1076), .B(n1051), .C(n1074), .YC(n1046), .YS(n1047) );
  FAX1 U810 ( .A(n1055), .B(n1078), .C(n1053), .YC(n1048), .YS(n1049) );
  FAX1 U811 ( .A(n1082), .B(n1057), .C(n1080), .YC(n1050), .YS(n1051) );
  FAX1 U812 ( .A(n1061), .B(n1084), .C(n1059), .YC(n1052), .YS(n1053) );
  FAX1 U813 ( .A(n1063), .B(n1088), .C(n1086), .YC(n1054), .YS(n1055) );
  FAX1 U814 ( .A(n1090), .B(n1067), .C(n1065), .YC(n1056), .YS(n1057) );
  FAX1 U815 ( .A(n1988), .B(n2020), .C(n1092), .YC(n1058), .YS(n1059) );
  FAX1 U816 ( .A(n1094), .B(n1956), .C(n2052), .YC(n1060), .YS(n1061) );
  FAX1 U817 ( .A(n1788), .B(n1898), .C(n1926), .YC(n1062), .YS(n1063) );
  FAX1 U818 ( .A(n1872), .B(n1806), .C(n1826), .YC(n1064), .YS(n1065) );
  FAX1 U819 ( .A(n1069), .B(n2084), .C(n1848), .YC(n1066), .YS(n1067) );
  FAX1 U821 ( .A(n1075), .B(n1098), .C(n1073), .YC(n1070), .YS(n1071) );
  FAX1 U822 ( .A(n1102), .B(n1077), .C(n1100), .YC(n1072), .YS(n1073) );
  FAX1 U823 ( .A(n1081), .B(n1104), .C(n1079), .YC(n1074), .YS(n1075) );
  FAX1 U824 ( .A(n1108), .B(n1083), .C(n1106), .YC(n1076), .YS(n1077) );
  FAX1 U825 ( .A(n1087), .B(n1110), .C(n1085), .YC(n1078), .YS(n1079) );
  FAX1 U826 ( .A(n1114), .B(n1112), .C(n1089), .YC(n1080), .YS(n1081) );
  FAX1 U827 ( .A(n1116), .B(n1093), .C(n1091), .YC(n1082), .YS(n1083) );
  FAX1 U828 ( .A(n1989), .B(n1120), .C(n1118), .YC(n1084), .YS(n1085) );
  FAX1 U829 ( .A(n2085), .B(n2021), .C(n1095), .YC(n1086), .YS(n1087) );
  FAX1 U830 ( .A(n1927), .B(n1957), .C(n2053), .YC(n1088), .YS(n1089) );
  FAX1 U831 ( .A(n1849), .B(n1827), .C(n1789), .YC(n1090), .YS(n1091) );
  FAX1 U832 ( .A(n1899), .B(n1873), .C(n1807), .YC(n1092), .YS(n1093) );
  FAX1 U833 ( .A(n2117), .B(n1122), .C(n1775), .YC(n1094), .YS(n1095) );
  FAX1 U834 ( .A(n1101), .B(n1126), .C(n1099), .YC(n1096), .YS(n1097) );
  FAX1 U835 ( .A(n1130), .B(n1103), .C(n1128), .YC(n1098), .YS(n1099) );
  FAX1 U836 ( .A(n1107), .B(n1132), .C(n1105), .YC(n1100), .YS(n1101) );
  FAX1 U837 ( .A(n1136), .B(n1109), .C(n1134), .YC(n1102), .YS(n1103) );
  FAX1 U838 ( .A(n1113), .B(n1138), .C(n1111), .YC(n1104), .YS(n1105) );
  FAX1 U839 ( .A(n1142), .B(n1115), .C(n1140), .YC(n1106), .YS(n1107) );
  FAX1 U840 ( .A(n1144), .B(n1119), .C(n1117), .YC(n1108), .YS(n1109) );
  FAX1 U841 ( .A(n1148), .B(n1146), .C(n1121), .YC(n1110), .YS(n1111) );
  FAX1 U842 ( .A(n2086), .B(n2022), .C(n2054), .YC(n1112), .YS(n1113) );
  FAX1 U843 ( .A(n1958), .B(n1150), .C(n1990), .YC(n1114), .YS(n1115) );
  FAX1 U844 ( .A(n1850), .B(n1808), .C(n1928), .YC(n1116), .YS(n1117) );
  FAX1 U845 ( .A(n1900), .B(n1828), .C(n1790), .YC(n1118), .YS(n1119) );
  FAX1 U846 ( .A(n1123), .B(n2118), .C(n1874), .YC(n1120), .YS(n1121) );
  FAX1 U848 ( .A(n1129), .B(n1154), .C(n1127), .YC(n1124), .YS(n1125) );
  FAX1 U849 ( .A(n1158), .B(n1131), .C(n1156), .YC(n1126), .YS(n1127) );
  FAX1 U850 ( .A(n1135), .B(n1160), .C(n1133), .YC(n1128), .YS(n1129) );
  FAX1 U851 ( .A(n1164), .B(n1137), .C(n1162), .YC(n1130), .YS(n1131) );
  FAX1 U852 ( .A(n1141), .B(n1166), .C(n1139), .YC(n1132), .YS(n1133) );
  FAX1 U853 ( .A(n1170), .B(n1143), .C(n1168), .YC(n1134), .YS(n1135) );
  FAX1 U854 ( .A(n1172), .B(n1147), .C(n1145), .YC(n1136), .YS(n1137) );
  FAX1 U855 ( .A(n1176), .B(n1174), .C(n1149), .YC(n1138), .YS(n1139) );
  FAX1 U856 ( .A(n2055), .B(n2023), .C(n1178), .YC(n1140), .YS(n1141) );
  FAX1 U857 ( .A(n2087), .B(n2119), .C(n1151), .YC(n1142), .YS(n1143) );
  FAX1 U858 ( .A(n1851), .B(n1959), .C(n1991), .YC(n1144), .YS(n1145) );
  FAX1 U859 ( .A(n1875), .B(n1809), .C(n1829), .YC(n1146), .YS(n1147) );
  FAX1 U860 ( .A(n1929), .B(n1901), .C(n1791), .YC(n1148), .YS(n1149) );
  FAX1 U861 ( .A(n2151), .B(n1180), .C(n1776), .YC(n1150), .YS(n1151) );
  FAX1 U862 ( .A(n1157), .B(n1184), .C(n1155), .YC(n1152), .YS(n1153) );
  FAX1 U863 ( .A(n1188), .B(n1159), .C(n1186), .YC(n1154), .YS(n1155) );
  FAX1 U864 ( .A(n1163), .B(n1190), .C(n1161), .YC(n1156), .YS(n1157) );
  FAX1 U865 ( .A(n1194), .B(n1165), .C(n1192), .YC(n1158), .YS(n1159) );
  FAX1 U866 ( .A(n1196), .B(n1169), .C(n1167), .YC(n1160), .YS(n1161) );
  FAX1 U867 ( .A(n1200), .B(n1171), .C(n1198), .YC(n1162), .YS(n1163) );
  FAX1 U868 ( .A(n1175), .B(n1173), .C(n1202), .YC(n1164), .YS(n1165) );
  FAX1 U869 ( .A(n1204), .B(n1179), .C(n1177), .YC(n1166), .YS(n1167) );
  FAX1 U870 ( .A(n2056), .B(n1208), .C(n1206), .YC(n1168), .YS(n1169) );
  FAX1 U871 ( .A(n2024), .B(n2120), .C(n2088), .YC(n1170), .YS(n1171) );
  FAX1 U872 ( .A(n1960), .B(n1992), .C(n1210), .YC(n1172), .YS(n1173) );
  FAX1 U873 ( .A(n1876), .B(n1810), .C(n1852), .YC(n1174), .YS(n1175) );
  FAX1 U874 ( .A(n1902), .B(n1792), .C(n1830), .YC(n1176), .YS(n1177) );
  FAX1 U875 ( .A(n1181), .B(n1930), .C(n2152), .YC(n1178), .YS(n1179) );
  FAX1 U878 ( .A(n1218), .B(n1189), .C(n1216), .YC(n1184), .YS(n1185) );
  FAX1 U879 ( .A(n1193), .B(n1220), .C(n1191), .YC(n1186), .YS(n1187) );
  FAX1 U880 ( .A(n1224), .B(n1195), .C(n1222), .YC(n1188), .YS(n1189) );
  FAX1 U881 ( .A(n1226), .B(n1199), .C(n1197), .YC(n1190), .YS(n1191) );
  FAX1 U882 ( .A(n1203), .B(n1201), .C(n1228), .YC(n1192), .YS(n1193) );
  FAX1 U883 ( .A(n1205), .B(n1232), .C(n1230), .YC(n1194), .YS(n1195) );
  FAX1 U884 ( .A(n1234), .B(n1209), .C(n1207), .YC(n1196), .YS(n1197) );
  FAX1 U885 ( .A(n2057), .B(n1238), .C(n1236), .YC(n1198), .YS(n1199) );
  FAX1 U886 ( .A(n2153), .B(n2089), .C(n1240), .YC(n1200), .YS(n1201) );
  FAX1 U887 ( .A(n2025), .B(n1211), .C(n2121), .YC(n1202), .YS(n1203) );
  FAX1 U888 ( .A(n1853), .B(n1877), .C(n1993), .YC(n1204), .YS(n1205) );
  FAX1 U889 ( .A(n1903), .B(n1811), .C(n1831), .YC(n1206), .YS(n1207) );
  FAX1 U890 ( .A(n1931), .B(n1961), .C(n1793), .YC(n1208), .YS(n1209) );
  FAX1 U891 ( .A(n1242), .B(n2185), .C(n1777), .YC(n1210), .YS(n1211) );
  FAX1 U892 ( .A(n1217), .B(n1246), .C(n1215), .YC(n1212), .YS(n1213) );
  FAX1 U893 ( .A(n1250), .B(n1219), .C(n1248), .YC(n1214), .YS(n1215) );
  FAX1 U894 ( .A(n1223), .B(n1252), .C(n1221), .YC(n1216), .YS(n1217) );
  FAX1 U895 ( .A(n1256), .B(n1225), .C(n1254), .YC(n1218), .YS(n1219) );
  FAX1 U896 ( .A(n1258), .B(n1229), .C(n1227), .YC(n1220), .YS(n1221) );
  FAX1 U897 ( .A(n1233), .B(n1231), .C(n1260), .YC(n1222), .YS(n1223) );
  FAX1 U898 ( .A(n1235), .B(n1264), .C(n1262), .YC(n1224), .YS(n1225) );
  FAX1 U899 ( .A(n1241), .B(n1239), .C(n1237), .YC(n1226), .YS(n1227) );
  FAX1 U900 ( .A(n1270), .B(n1268), .C(n1266), .YC(n1228), .YS(n1229) );
  FAX1 U901 ( .A(n2090), .B(n2122), .C(n1272), .YC(n1230), .YS(n1231) );
  FAX1 U902 ( .A(n2026), .B(n2058), .C(n2154), .YC(n1232), .YS(n1233) );
  FAX1 U903 ( .A(n1854), .B(n1878), .C(n1994), .YC(n1234), .YS(n1235) );
  FAX1 U904 ( .A(n1904), .B(n1812), .C(n1832), .YC(n1236), .YS(n1237) );
  FAX1 U905 ( .A(n1962), .B(n1932), .C(n1794), .YC(n1238), .YS(n1239) );
  FAX1 U906 ( .A(n1274), .B(n1778), .C(n2186), .YC(n1240), .YS(n1241) );
  FAX1 U908 ( .A(n1249), .B(n1277), .C(n1247), .YC(n1244), .YS(n1245) );
  FAX1 U909 ( .A(n1281), .B(n1251), .C(n1279), .YC(n1246), .YS(n1247) );
  FAX1 U910 ( .A(n1255), .B(n1283), .C(n1253), .YC(n1248), .YS(n1249) );
  FAX1 U911 ( .A(n1287), .B(n1257), .C(n1285), .YC(n1250), .YS(n1251) );
  FAX1 U912 ( .A(n1289), .B(n1261), .C(n1259), .YC(n1252), .YS(n1253) );
  FAX1 U913 ( .A(n1265), .B(n1291), .C(n1263), .YC(n1254), .YS(n1255) );
  FAX1 U914 ( .A(n1267), .B(n1295), .C(n1293), .YC(n1256), .YS(n1257) );
  FAX1 U915 ( .A(n1297), .B(n1271), .C(n1269), .YC(n1258), .YS(n1259) );
  FAX1 U916 ( .A(n1301), .B(n1299), .C(n1273), .YC(n1260), .YS(n1261) );
  FAX1 U917 ( .A(n2123), .B(n2091), .C(n1303), .YC(n1262), .YS(n1263) );
  FAX1 U918 ( .A(n2059), .B(n2155), .C(n2187), .YC(n1264), .YS(n1265) );
  FAX1 U919 ( .A(n1855), .B(n1879), .C(n2027), .YC(n1266), .YS(n1267) );
  FAX1 U920 ( .A(n1905), .B(n1833), .C(n1813), .YC(n1268), .YS(n1269) );
  FAX1 U921 ( .A(n1963), .B(n1933), .C(n1795), .YC(n1270), .YS(n1271) );
  FAX1 U922 ( .A(n1274), .B(n1779), .C(n1995), .YC(n1272), .YS(n1273) );
  FAX1 U924 ( .A(n1280), .B(n1307), .C(n1278), .YC(n1275), .YS(n1276) );
  FAX1 U925 ( .A(n1311), .B(n1282), .C(n1309), .YC(n1277), .YS(n1278) );
  FAX1 U926 ( .A(n1286), .B(n1313), .C(n1284), .YC(n1279), .YS(n1280) );
  FAX1 U927 ( .A(n1290), .B(n1288), .C(n1315), .YC(n1281), .YS(n1282) );
  FAX1 U928 ( .A(n1319), .B(n1292), .C(n1317), .YC(n1283), .YS(n1284) );
  FAX1 U929 ( .A(n1296), .B(n1294), .C(n1321), .YC(n1285), .YS(n1286) );
  FAX1 U930 ( .A(n1300), .B(n1325), .C(n1323), .YC(n1287), .YS(n1288) );
  FAX1 U931 ( .A(n1304), .B(n1302), .C(n1298), .YC(n1289), .YS(n1290) );
  FAX1 U932 ( .A(n1331), .B(n1329), .C(n1327), .YC(n1291), .YS(n1292) );
  FAX1 U933 ( .A(n2188), .B(n2124), .C(n2156), .YC(n1293), .YS(n1294) );
  FAX1 U934 ( .A(n2060), .B(n1333), .C(n2092), .YC(n1295), .YS(n1296) );
  FAX1 U935 ( .A(n1856), .B(n1880), .C(n2028), .YC(n1297), .YS(n1298) );
  FAX1 U936 ( .A(n1906), .B(n1834), .C(n1814), .YC(n1299), .YS(n1300) );
  FAX1 U937 ( .A(n1996), .B(n1934), .C(n1796), .YC(n1301), .YS(n1302) );
  FAX1 U939 ( .A(n1310), .B(n1337), .C(n1308), .YC(n1305), .YS(n1306) );
  FAX1 U940 ( .A(n1341), .B(n1312), .C(n1339), .YC(n1307), .YS(n1308) );
  FAX1 U941 ( .A(n1316), .B(n1343), .C(n1314), .YC(n1309), .YS(n1310) );
  FAX1 U942 ( .A(n1320), .B(n1345), .C(n1318), .YC(n1311), .YS(n1312) );
  FAX1 U943 ( .A(n1349), .B(n1322), .C(n1347), .YC(n1313), .YS(n1314) );
  FAX1 U944 ( .A(n1326), .B(n1351), .C(n1324), .YC(n1315), .YS(n1316) );
  FAX1 U945 ( .A(n1330), .B(n1328), .C(n1353), .YC(n1317), .YS(n1318) );
  FAX1 U946 ( .A(n1357), .B(n1355), .C(n1332), .YC(n1319), .YS(n1320) );
  FAX1 U947 ( .A(n2125), .B(n1361), .C(n1359), .YC(n1321), .YS(n1322) );
  FAX1 U948 ( .A(n2220), .B(n2157), .C(n1334), .YC(n1323), .YS(n1324) );
  FAX1 U949 ( .A(n2061), .B(n2093), .C(n2189), .YC(n1325), .YS(n1326) );
  FAX1 U950 ( .A(n1857), .B(n1881), .C(n1755), .YC(n1327), .YS(n1328) );
  FAX1 U951 ( .A(n1907), .B(n1835), .C(n1815), .YC(n1329), .YS(n1330) );
  FAX1 U952 ( .A(n1997), .B(n1965), .C(n1797), .YC(n1331), .YS(n1332) );
  HAX1 U953 ( .A(n2029), .B(n1935), .YC(n1333), .YS(n1334) );
  FAX1 U954 ( .A(n1340), .B(n1365), .C(n1338), .YC(n1335), .YS(n1336) );
  FAX1 U955 ( .A(n1369), .B(n1342), .C(n1367), .YC(n1337), .YS(n1338) );
  FAX1 U956 ( .A(n1346), .B(n1371), .C(n1344), .YC(n1339), .YS(n1340) );
  FAX1 U957 ( .A(n1350), .B(n1348), .C(n1373), .YC(n1341), .YS(n1342) );
  FAX1 U958 ( .A(n1377), .B(n1352), .C(n1375), .YC(n1343), .YS(n1344) );
  FAX1 U959 ( .A(n1381), .B(n1379), .C(n1354), .YC(n1345), .YS(n1346) );
  FAX1 U960 ( .A(n1358), .B(n1360), .C(n1356), .YC(n1347), .YS(n1348) );
  FAX1 U961 ( .A(n1385), .B(n1383), .C(n1362), .YC(n1349), .YS(n1350) );
  FAX1 U962 ( .A(n2221), .B(n2158), .C(n1387), .YC(n1351), .YS(n1352) );
  FAX1 U963 ( .A(n1389), .B(n2126), .C(n2190), .YC(n1353), .YS(n1354) );
  FAX1 U964 ( .A(n1936), .B(n2062), .C(n2094), .YC(n1355), .YS(n1356) );
  FAX1 U965 ( .A(n1908), .B(n1836), .C(n1882), .YC(n1357), .YS(n1358) );
  FAX1 U966 ( .A(n1966), .B(n1858), .C(n1816), .YC(n1359), .YS(n1360) );
  FAX1 U967 ( .A(n1798), .B(n1998), .C(n2030), .YC(n1361), .YS(n1362) );
  FAX1 U968 ( .A(n1368), .B(n1393), .C(n1366), .YC(n1363), .YS(n1364) );
  FAX1 U969 ( .A(n1372), .B(n1370), .C(n1395), .YC(n1365), .YS(n1366) );
  FAX1 U970 ( .A(n1399), .B(n1374), .C(n1397), .YC(n1367), .YS(n1368) );
  FAX1 U971 ( .A(n1378), .B(n1401), .C(n1376), .YC(n1369), .YS(n1370) );
  FAX1 U972 ( .A(n1380), .B(n1405), .C(n1403), .YC(n1371), .YS(n1372) );
  FAX1 U973 ( .A(n1386), .B(n1407), .C(n1382), .YC(n1373), .YS(n1374) );
  FAX1 U974 ( .A(n1409), .B(n1388), .C(n1384), .YC(n1375), .YS(n1376) );
  FAX1 U975 ( .A(n1415), .B(n1413), .C(n1411), .YC(n1377), .YS(n1378) );
  FAX1 U976 ( .A(n2191), .B(n2159), .C(n1390), .YC(n1379), .YS(n1380) );
  FAX1 U977 ( .A(n2095), .B(n2127), .C(n2222), .YC(n1381), .YS(n1382) );
  FAX1 U978 ( .A(n1883), .B(n1909), .C(n1756), .YC(n1383), .YS(n1384) );
  FAX1 U979 ( .A(n1999), .B(n1837), .C(n1859), .YC(n1385), .YS(n1386) );
  FAX1 U980 ( .A(n2031), .B(n1937), .C(n1817), .YC(n1387), .YS(n1388) );
  HAX1 U981 ( .A(n2063), .B(n1967), .YC(n1389), .YS(n1390) );
  FAX1 U982 ( .A(n1396), .B(n1419), .C(n1394), .YC(n1391), .YS(n1392) );
  FAX1 U983 ( .A(n1423), .B(n1398), .C(n1421), .YC(n1393), .YS(n1394) );
  FAX1 U984 ( .A(n1402), .B(n1425), .C(n1400), .YC(n1395), .YS(n1396) );
  FAX1 U985 ( .A(n1406), .B(n1427), .C(n1404), .YC(n1397), .YS(n1398) );
  FAX1 U986 ( .A(n1431), .B(n1408), .C(n1429), .YC(n1399), .YS(n1400) );
  FAX1 U987 ( .A(n1412), .B(n1410), .C(n1433), .YC(n1401), .YS(n1402) );
  FAX1 U988 ( .A(n1435), .B(n1416), .C(n1414), .YC(n1403), .YS(n1404) );
  FAX1 U989 ( .A(n2192), .B(n1439), .C(n1437), .YC(n1405), .YS(n1406) );
  FAX1 U990 ( .A(n1441), .B(n2160), .C(n2223), .YC(n1407), .YS(n1408) );
  FAX1 U991 ( .A(n1938), .B(n2096), .C(n2128), .YC(n1409), .YS(n1410) );
  FAX1 U992 ( .A(n1968), .B(n1884), .C(n1910), .YC(n1411), .YS(n1412) );
  FAX1 U993 ( .A(n2000), .B(n1860), .C(n1838), .YC(n1413), .YS(n1414) );
  FAX1 U994 ( .A(n1818), .B(n2064), .C(n2032), .YC(n1415), .YS(n1416) );
  FAX1 U995 ( .A(n1422), .B(n1445), .C(n1420), .YC(n1417), .YS(n1418) );
  FAX1 U996 ( .A(n1449), .B(n1424), .C(n1447), .YC(n1419), .YS(n1420) );
  FAX1 U997 ( .A(n1428), .B(n1451), .C(n1426), .YC(n1421), .YS(n1422) );
  FAX1 U998 ( .A(n1432), .B(n1453), .C(n1430), .YC(n1423), .YS(n1424) );
  FAX1 U999 ( .A(n1457), .B(n1434), .C(n1455), .YC(n1425), .YS(n1426) );
  FAX1 U1000 ( .A(n1440), .B(n1438), .C(n1436), .YC(n1427), .YS(n1428) );
  FAX1 U1001 ( .A(n1463), .B(n1461), .C(n1459), .YC(n1429), .YS(n1430) );
  FAX1 U1002 ( .A(n2193), .B(n1442), .C(n1465), .YC(n1431), .YS(n1432) );
  FAX1 U1003 ( .A(n2129), .B(n2161), .C(n2224), .YC(n1433), .YS(n1434) );
  FAX1 U1004 ( .A(n1861), .B(n1885), .C(n1757), .YC(n1435), .YS(n1436) );
  FAX1 U1005 ( .A(n1939), .B(n2033), .C(n1911), .YC(n1437), .YS(n1438) );
  FAX1 U1006 ( .A(n2097), .B(n2001), .C(n1839), .YC(n1439), .YS(n1440) );
  HAX1 U1007 ( .A(n2065), .B(n1969), .YC(n1441), .YS(n1442) );
  FAX1 U1009 ( .A(n1473), .B(n1450), .C(n1471), .YC(n1445), .YS(n1446) );
  FAX1 U1010 ( .A(n1454), .B(n1475), .C(n1452), .YC(n1447), .YS(n1448) );
  FAX1 U1011 ( .A(n1479), .B(n1477), .C(n1456), .YC(n1449), .YS(n1450) );
  FAX1 U1012 ( .A(n1460), .B(n1481), .C(n1458), .YC(n1451), .YS(n1452) );
  FAX1 U1013 ( .A(n1466), .B(n1464), .C(n1462), .YC(n1453), .YS(n1454) );
  FAX1 U1014 ( .A(n1487), .B(n1485), .C(n1483), .YC(n1455), .YS(n1456) );
  FAX1 U1015 ( .A(n1489), .B(n2194), .C(n2225), .YC(n1457), .YS(n1458) );
  FAX1 U1016 ( .A(n1912), .B(n2130), .C(n2162), .YC(n1459), .YS(n1460) );
  FAX1 U1017 ( .A(n1940), .B(n1886), .C(n1970), .YC(n1461), .YS(n1462) );
  FAX1 U1018 ( .A(n2002), .B(n2034), .C(n1862), .YC(n1463), .YS(n1464) );
  FAX1 U1019 ( .A(n1840), .B(n2098), .C(n2066), .YC(n1465), .YS(n1466) );
  FAX1 U1020 ( .A(n1472), .B(n1493), .C(n1470), .YC(n1467), .YS(n1468) );
  FAX1 U1021 ( .A(n1497), .B(n1474), .C(n1495), .YC(n1469), .YS(n1470) );
  FAX1 U1022 ( .A(n1499), .B(n1478), .C(n1476), .YC(n1471), .YS(n1472) );
  FAX1 U1023 ( .A(n1503), .B(n1501), .C(n1480), .YC(n1473), .YS(n1474) );
  FAX1 U1024 ( .A(n1486), .B(n1484), .C(n1482), .YC(n1475), .YS(n1476) );
  FAX1 U1025 ( .A(n1507), .B(n1505), .C(n1488), .YC(n1477), .YS(n1478) );
  FAX1 U1026 ( .A(n1490), .B(n1511), .C(n1509), .YC(n1479), .YS(n1480) );
  FAX1 U1027 ( .A(n2163), .B(n2195), .C(n2226), .YC(n1481), .YS(n1482) );
  FAX1 U1028 ( .A(n1887), .B(n2035), .C(n1758), .YC(n1483), .YS(n1484) );
  FAX1 U1029 ( .A(n1941), .B(n2067), .C(n1913), .YC(n1485), .YS(n1486) );
  FAX1 U1030 ( .A(n2131), .B(n2003), .C(n1863), .YC(n1487), .YS(n1488) );
  HAX1 U1031 ( .A(n2099), .B(n1971), .YC(n1489), .YS(n1490) );
  FAX1 U1032 ( .A(n1496), .B(n1515), .C(n1494), .YC(n1491), .YS(n1492) );
  FAX1 U1033 ( .A(n1519), .B(n1498), .C(n1517), .YC(n1493), .YS(n1494) );
  FAX1 U1034 ( .A(n1521), .B(n1502), .C(n1500), .YC(n1495), .YS(n1496) );
  FAX1 U1035 ( .A(n1525), .B(n1523), .C(n1504), .YC(n1497), .YS(n1498) );
  FAX1 U1036 ( .A(n1510), .B(n1508), .C(n1506), .YC(n1499), .YS(n1500) );
  FAX1 U1037 ( .A(n1529), .B(n1527), .C(n1512), .YC(n1501), .YS(n1502) );
  FAX1 U1038 ( .A(n1533), .B(n2227), .C(n1531), .YC(n1503), .YS(n1504) );
  FAX1 U1039 ( .A(n1942), .B(n2164), .C(n2196), .YC(n1505), .YS(n1506) );
  FAX1 U1040 ( .A(n2036), .B(n2068), .C(n1972), .YC(n1507), .YS(n1508) );
  FAX1 U1041 ( .A(n2004), .B(n1914), .C(n1888), .YC(n1509), .YS(n1510) );
  FAX1 U1042 ( .A(n1864), .B(n2100), .C(n2132), .YC(n1511), .YS(n1512) );
  FAX1 U1045 ( .A(n1543), .B(n1524), .C(n1522), .YC(n1517), .YS(n1518) );
  FAX1 U1046 ( .A(n1530), .B(n1526), .C(n1545), .YC(n1519), .YS(n1520) );
  FAX1 U1047 ( .A(n1547), .B(n1532), .C(n1528), .YC(n1521), .YS(n1522) );
  FAX1 U1048 ( .A(n1553), .B(n1551), .C(n1549), .YC(n1523), .YS(n1524) );
  FAX1 U1049 ( .A(n2197), .B(n2228), .C(n1534), .YC(n1525), .YS(n1526) );
  FAX1 U1050 ( .A(n2101), .B(n1915), .C(n1759), .YC(n1527), .YS(n1528) );
  FAX1 U1051 ( .A(n2037), .B(n2069), .C(n1943), .YC(n1529), .YS(n1530) );
  FAX1 U1052 ( .A(n2133), .B(n2005), .C(n1889), .YC(n1531), .YS(n1532) );
  HAX1 U1053 ( .A(n2165), .B(n1973), .YC(n1533), .YS(n1534) );
  FAX1 U1054 ( .A(n1540), .B(n1557), .C(n1538), .YC(n1535), .YS(n1536) );
  FAX1 U1055 ( .A(n1544), .B(n1542), .C(n1559), .YC(n1537), .YS(n1538) );
  FAX1 U1056 ( .A(n1563), .B(n1546), .C(n1561), .YC(n1539), .YS(n1540) );
  FAX1 U1057 ( .A(n1552), .B(n1548), .C(n1565), .YC(n1541), .YS(n1542) );
  FAX1 U1058 ( .A(n1567), .B(n1554), .C(n1550), .YC(n1543), .YS(n1544) );
  FAX1 U1059 ( .A(n1573), .B(n1571), .C(n1569), .YC(n1545), .YS(n1546) );
  FAX1 U1060 ( .A(n2070), .B(n2198), .C(n2229), .YC(n1547), .YS(n1548) );
  FAX1 U1061 ( .A(n2006), .B(n2102), .C(n1974), .YC(n1549), .YS(n1550) );
  FAX1 U1062 ( .A(n2038), .B(n1944), .C(n1916), .YC(n1551), .YS(n1552) );
  FAX1 U1063 ( .A(n1890), .B(n2134), .C(n2166), .YC(n1553), .YS(n1554) );
  FAX1 U1064 ( .A(n1560), .B(n1577), .C(n1558), .YC(n1555), .YS(n1556) );
  FAX1 U1065 ( .A(n1564), .B(n1562), .C(n1579), .YC(n1557), .YS(n1558) );
  FAX1 U1066 ( .A(n1583), .B(n1566), .C(n1581), .YC(n1559), .YS(n1560) );
  FAX1 U1067 ( .A(n1570), .B(n1568), .C(n1585), .YC(n1561), .YS(n1562) );
  FAX1 U1068 ( .A(n1589), .B(n1587), .C(n1572), .YC(n1563), .YS(n1564) );
  FAX1 U1069 ( .A(n2230), .B(n1574), .C(n1591), .YC(n1565), .YS(n1566) );
  FAX1 U1070 ( .A(n2135), .B(n2103), .C(n1760), .YC(n1567), .YS(n1568) );
  FAX1 U1071 ( .A(n2007), .B(n1945), .C(n2071), .YC(n1569), .YS(n1570) );
  FAX1 U1072 ( .A(n2167), .B(n2039), .C(n1917), .YC(n1571), .YS(n1572) );
  HAX1 U1073 ( .A(n2199), .B(n1975), .YC(n1573), .YS(n1574) );
  FAX1 U1074 ( .A(n1580), .B(n1595), .C(n1578), .YC(n1575), .YS(n1576) );
  FAX1 U1075 ( .A(n1584), .B(n1582), .C(n1597), .YC(n1577), .YS(n1578) );
  FAX1 U1076 ( .A(n1586), .B(n1601), .C(n1599), .YC(n1579), .YS(n1580) );
  FAX1 U1077 ( .A(n1592), .B(n1588), .C(n1590), .YC(n1581), .YS(n1582) );
  FAX1 U1078 ( .A(n1607), .B(n1605), .C(n1603), .YC(n1583), .YS(n1584) );
  FAX1 U1079 ( .A(n2136), .B(n2231), .C(n1609), .YC(n1585), .YS(n1586) );
  FAX1 U1080 ( .A(n2072), .B(n2104), .C(n2008), .YC(n1587), .YS(n1588) );
  FAX1 U1081 ( .A(n2040), .B(n1976), .C(n1946), .YC(n1589), .YS(n1590) );
  FAX1 U1082 ( .A(n1918), .B(n2200), .C(n2168), .YC(n1591), .YS(n1592) );
  FAX1 U1083 ( .A(n1598), .B(n1613), .C(n1596), .YC(n1593), .YS(n1594) );
  FAX1 U1084 ( .A(n1602), .B(n1600), .C(n1615), .YC(n1595), .YS(n1596) );
  FAX1 U1085 ( .A(n1604), .B(n1619), .C(n1617), .YC(n1597), .YS(n1598) );
  FAX1 U1086 ( .A(n1621), .B(n1608), .C(n1606), .YC(n1599), .YS(n1600) );
  FAX1 U1087 ( .A(n1610), .B(n1625), .C(n1623), .YC(n1601), .YS(n1602) );
  FAX1 U1088 ( .A(n2137), .B(n2105), .C(n1761), .YC(n1603), .YS(n1604) );
  FAX1 U1089 ( .A(n2073), .B(n2169), .C(n2009), .YC(n1605), .YS(n1606) );
  FAX1 U1090 ( .A(n2201), .B(n2041), .C(n1947), .YC(n1607), .YS(n1608) );
  HAX1 U1091 ( .A(n2232), .B(n1977), .YC(n1609), .YS(n1610) );
  FAX1 U1094 ( .A(n1624), .B(n1635), .C(n1633), .YC(n1615), .YS(n1616) );
  FAX1 U1095 ( .A(n1637), .B(n1626), .C(n1622), .YC(n1617), .YS(n1618) );
  FAX1 U1096 ( .A(n2106), .B(n1641), .C(n1639), .YC(n1619), .YS(n1620) );
  FAX1 U1097 ( .A(n2138), .B(n2042), .C(n2074), .YC(n1621), .YS(n1622) );
  FAX1 U1098 ( .A(n2170), .B(n2010), .C(n1978), .YC(n1623), .YS(n1624) );
  FAX1 U1099 ( .A(n1948), .B(n2233), .C(n2202), .YC(n1625), .YS(n1626) );
  FAX1 U1100 ( .A(n1632), .B(n1645), .C(n1630), .YC(n1627), .YS(n1628) );
  FAX1 U1101 ( .A(n1649), .B(n1647), .C(n1634), .YC(n1629), .YS(n1630) );
  FAX1 U1102 ( .A(n1638), .B(n1640), .C(n1636), .YC(n1631), .YS(n1632) );
  FAX1 U1103 ( .A(n1655), .B(n1653), .C(n1651), .YC(n1633), .YS(n1634) );
  FAX1 U1104 ( .A(n2139), .B(n1762), .C(n1642), .YC(n1635), .YS(n1636) );
  FAX1 U1105 ( .A(n2043), .B(n2171), .C(n2107), .YC(n1637), .YS(n1638) );
  FAX1 U1106 ( .A(n2075), .B(n2203), .C(n1979), .YC(n1639), .YS(n1640) );
  HAX1 U1107 ( .A(n2234), .B(n2011), .YC(n1641), .YS(n1642) );
  FAX1 U1108 ( .A(n1648), .B(n1659), .C(n1646), .YC(n1643), .YS(n1644) );
  FAX1 U1109 ( .A(n1663), .B(n1661), .C(n1650), .YC(n1645), .YS(n1646) );
  FAX1 U1110 ( .A(n1656), .B(n1652), .C(n1654), .YC(n1647), .YS(n1648) );
  FAX1 U1111 ( .A(n1669), .B(n1667), .C(n1665), .YC(n1649), .YS(n1650) );
  FAX1 U1112 ( .A(n2140), .B(n2076), .C(n2108), .YC(n1651), .YS(n1652) );
  FAX1 U1113 ( .A(n2172), .B(n2044), .C(n2012), .YC(n1653), .YS(n1654) );
  FAX1 U1114 ( .A(n1980), .B(n2235), .C(n2204), .YC(n1655), .YS(n1656) );
  FAX1 U1115 ( .A(n1662), .B(n1673), .C(n1660), .YC(n1657), .YS(n1658) );
  FAX1 U1116 ( .A(n1677), .B(n1675), .C(n1664), .YC(n1659), .YS(n1660) );
  FAX1 U1117 ( .A(n1679), .B(n1666), .C(n1668), .YC(n1661), .YS(n1662) );
  FAX1 U1118 ( .A(n1763), .B(n1670), .C(n1681), .YC(n1663), .YS(n1664) );
  FAX1 U1119 ( .A(n2173), .B(n2077), .C(n2141), .YC(n1665), .YS(n1666) );
  FAX1 U1120 ( .A(n2109), .B(n2205), .C(n2013), .YC(n1667), .YS(n1668) );
  HAX1 U1121 ( .A(n2236), .B(n2045), .YC(n1669), .YS(n1670) );
  FAX1 U1122 ( .A(n1676), .B(n1685), .C(n1674), .YC(n1671), .YS(n1672) );
  FAX1 U1123 ( .A(n1680), .B(n1678), .C(n1687), .YC(n1673), .YS(n1674) );
  FAX1 U1124 ( .A(n1691), .B(n1689), .C(n1682), .YC(n1675), .YS(n1676) );
  FAX1 U1125 ( .A(n2142), .B(n2110), .C(n1693), .YC(n1677), .YS(n1678) );
  FAX1 U1126 ( .A(n2174), .B(n2078), .C(n2046), .YC(n1679), .YS(n1680) );
  FAX1 U1127 ( .A(n2014), .B(n2237), .C(n2206), .YC(n1681), .YS(n1682) );
  FAX1 U1128 ( .A(n1688), .B(n1697), .C(n1686), .YC(n1683), .YS(n1684) );
  FAX1 U1129 ( .A(n1692), .B(n1690), .C(n1699), .YC(n1685), .YS(n1686) );
  FAX1 U1130 ( .A(n1694), .B(n1703), .C(n1701), .YC(n1687), .YS(n1688) );
  FAX1 U1131 ( .A(n2175), .B(n2143), .C(n1764), .YC(n1689), .YS(n1690) );
  FAX1 U1132 ( .A(n2111), .B(n2207), .C(n2047), .YC(n1691), .YS(n1692) );
  HAX1 U1133 ( .A(n2238), .B(n2079), .YC(n1693), .YS(n1694) );
  FAX1 U1134 ( .A(n1707), .B(n1700), .C(n1698), .YC(n1695), .YS(n1696) );
  FAX1 U1135 ( .A(n1704), .B(n1702), .C(n1709), .YC(n1697), .YS(n1698) );
  FAX1 U1136 ( .A(n2144), .B(n1713), .C(n1711), .YC(n1699), .YS(n1700) );
  FAX1 U1137 ( .A(n2176), .B(n2112), .C(n2080), .YC(n1701), .YS(n1702) );
  FAX1 U1138 ( .A(n2048), .B(n2239), .C(n2208), .YC(n1703), .YS(n1704) );
  FAX1 U1139 ( .A(n1710), .B(n1717), .C(n1708), .YC(n1705), .YS(n1706) );
  FAX1 U1140 ( .A(n1721), .B(n1719), .C(n1712), .YC(n1707), .YS(n1708) );
  FAX1 U1141 ( .A(n2209), .B(n1765), .C(n1714), .YC(n1709), .YS(n1710) );
  FAX1 U1142 ( .A(n2145), .B(n2177), .C(n2081), .YC(n1711), .YS(n1712) );
  HAX1 U1143 ( .A(n2240), .B(n2113), .YC(n1713), .YS(n1714) );
  FAX1 U1144 ( .A(n1720), .B(n1725), .C(n1718), .YC(n1715), .YS(n1716) );
  FAX1 U1145 ( .A(n1729), .B(n1727), .C(n1722), .YC(n1717), .YS(n1718) );
  FAX1 U1146 ( .A(n2178), .B(n2146), .C(n2114), .YC(n1719), .YS(n1720) );
  FAX1 U1147 ( .A(n2082), .B(n2241), .C(n2210), .YC(n1721), .YS(n1722) );
  FAX1 U1148 ( .A(n1728), .B(n1733), .C(n1726), .YC(n1723), .YS(n1724) );
  FAX1 U1149 ( .A(n1766), .B(n1730), .C(n1735), .YC(n1725), .YS(n1726) );
  FAX1 U1150 ( .A(n2211), .B(n2179), .C(n2115), .YC(n1727), .YS(n1728) );
  HAX1 U1151 ( .A(n2242), .B(n2147), .YC(n1729), .YS(n1730) );
  FAX1 U1152 ( .A(n1739), .B(n1736), .C(n1734), .YC(n1731), .YS(n1732) );
  FAX1 U1153 ( .A(n2180), .B(n2148), .C(n1741), .YC(n1733), .YS(n1734) );
  FAX1 U1154 ( .A(n2116), .B(n2243), .C(n2212), .YC(n1735), .YS(n1736) );
  FAX1 U1155 ( .A(n1742), .B(n1745), .C(n1740), .YC(n1737), .YS(n1738) );
  FAX1 U1156 ( .A(n2213), .B(n2149), .C(n1767), .YC(n1739), .YS(n1740) );
  HAX1 U1157 ( .A(n2244), .B(n2181), .YC(n1741), .YS(n1742) );
  FAX1 U1158 ( .A(n2182), .B(n1749), .C(n1746), .YC(n1743), .YS(n1744) );
  FAX1 U1159 ( .A(n2150), .B(n2245), .C(n2214), .YC(n1745), .YS(n1746) );
  FAX1 U1160 ( .A(n2183), .B(n1768), .C(n1750), .YC(n1747), .YS(n1748) );
  HAX1 U1161 ( .A(n2246), .B(n2215), .YC(n1749), .YS(n1750) );
  FAX1 U1162 ( .A(n2184), .B(n2247), .C(n2216), .YC(n1751), .YS(n1752) );
  HAX1 U1163 ( .A(n2248), .B(n2217), .YC(n1753), .YS(n1754) );
  NOR2X1 U1164 ( .A(n3054), .B(n3093), .Y(n1771) );
  NOR2X1 U1165 ( .A(n3054), .B(n3090), .Y(n930) );
  NOR2X1 U1166 ( .A(n3054), .B(n3088), .Y(n1772) );
  NOR2X1 U1167 ( .A(n3054), .B(n3085), .Y(n972) );
  NOR2X1 U1168 ( .A(n3054), .B(n3083), .Y(n1773) );
  NOR2X1 U1169 ( .A(n3054), .B(n3081), .Y(n1018) );
  NOR2X1 U1170 ( .A(n3054), .B(n3079), .Y(n1774) );
  NOR2X1 U1171 ( .A(n3054), .B(n3077), .Y(n1068) );
  NOR2X1 U1172 ( .A(n3054), .B(n3075), .Y(n1775) );
  NOR2X1 U1173 ( .A(n3054), .B(n3073), .Y(n1122) );
  NOR2X1 U1174 ( .A(n3054), .B(n3071), .Y(n1776) );
  NOR2X1 U1175 ( .A(n3054), .B(n3068), .Y(n1180) );
  NOR2X1 U1176 ( .A(n3054), .B(n3065), .Y(n1777) );
  NOR2X1 U1177 ( .A(n3054), .B(n3063), .Y(n1778) );
  NOR2X1 U1178 ( .A(n3054), .B(n3060), .Y(n1779) );
  OAI22X1 U1194 ( .A(n3054), .B(n2931), .C(n2927), .D(n2284), .Y(n1755) );
  OAI22X1 U1195 ( .A(n2931), .B(n2267), .C(n2927), .D(n2266), .Y(n1781) );
  OAI22X1 U1196 ( .A(n2927), .B(n2267), .C(n2931), .D(n2268), .Y(n1782) );
  OAI22X1 U1197 ( .A(n2931), .B(n2269), .C(n2927), .D(n2268), .Y(n1783) );
  OAI22X1 U1198 ( .A(n2927), .B(n2269), .C(n2931), .D(n2270), .Y(n1784) );
  OAI22X1 U1199 ( .A(n2931), .B(n2271), .C(n2927), .D(n2270), .Y(n1785) );
  OAI22X1 U1200 ( .A(n2927), .B(n2271), .C(n2931), .D(n2272), .Y(n1786) );
  OAI22X1 U1201 ( .A(n2931), .B(n2273), .C(n2927), .D(n2272), .Y(n1787) );
  OAI22X1 U1202 ( .A(n2927), .B(n2273), .C(n2931), .D(n2274), .Y(n1788) );
  OAI22X1 U1203 ( .A(n2931), .B(n2275), .C(n2927), .D(n2274), .Y(n1789) );
  OAI22X1 U1204 ( .A(n2927), .B(n2275), .C(n2931), .D(n2276), .Y(n1790) );
  OAI22X1 U1205 ( .A(n2931), .B(n2277), .C(n2927), .D(n2276), .Y(n1791) );
  OAI22X1 U1206 ( .A(n2927), .B(n2277), .C(n2931), .D(n2278), .Y(n1792) );
  OAI22X1 U1207 ( .A(n2931), .B(n2279), .C(n2927), .D(n2278), .Y(n1793) );
  OAI22X1 U1208 ( .A(n2927), .B(n2279), .C(n2931), .D(n2280), .Y(n1794) );
  OAI22X1 U1209 ( .A(n2931), .B(n2281), .C(n2927), .D(n2280), .Y(n1795) );
  OAI22X1 U1210 ( .A(n2927), .B(n2281), .C(n2931), .D(n2282), .Y(n1796) );
  OAI22X1 U1211 ( .A(n2931), .B(n2283), .C(n2927), .D(n2282), .Y(n1797) );
  XNOR2X1 U1212 ( .A(n3097), .B(n3052), .Y(n2266) );
  XNOR2X1 U1213 ( .A(n3094), .B(n3052), .Y(n2267) );
  XNOR2X1 U1214 ( .A(n3091), .B(n3052), .Y(n2268) );
  XNOR2X1 U1215 ( .A(n3089), .B(n3052), .Y(n2269) );
  XNOR2X1 U1216 ( .A(n3086), .B(n3052), .Y(n2270) );
  XNOR2X1 U1217 ( .A(n3084), .B(n3052), .Y(n2271) );
  XNOR2X1 U1218 ( .A(n3082), .B(n3052), .Y(n2272) );
  XNOR2X1 U1219 ( .A(n3080), .B(n3052), .Y(n2273) );
  XNOR2X1 U1220 ( .A(n3078), .B(n3052), .Y(n2274) );
  XNOR2X1 U1221 ( .A(n3076), .B(n3052), .Y(n2275) );
  XNOR2X1 U1222 ( .A(n3074), .B(n3053), .Y(n2276) );
  XNOR2X1 U1223 ( .A(n3072), .B(n3053), .Y(n2277) );
  XNOR2X1 U1224 ( .A(n3070), .B(n3053), .Y(n2278) );
  XNOR2X1 U1225 ( .A(n3067), .B(n3053), .Y(n2279) );
  XNOR2X1 U1226 ( .A(n3064), .B(n3052), .Y(n2280) );
  XNOR2X1 U1227 ( .A(n3062), .B(n3053), .Y(n2281) );
  XNOR2X1 U1228 ( .A(n437), .B(n3053), .Y(n2282) );
  XNOR2X1 U1229 ( .A(n3055), .B(n3052), .Y(n2283) );
  OAI22X1 U1230 ( .A(n3114), .B(n2930), .C(n2926), .D(n2305), .Y(n1756) );
  OAI22X1 U1231 ( .A(n2930), .B(n2286), .C(n2926), .D(n2285), .Y(n1799) );
  OAI22X1 U1232 ( .A(n2926), .B(n2286), .C(n2930), .D(n2287), .Y(n1800) );
  OAI22X1 U1233 ( .A(n2930), .B(n2288), .C(n2926), .D(n2287), .Y(n1801) );
  OAI22X1 U1234 ( .A(n2926), .B(n2288), .C(n2930), .D(n2289), .Y(n1802) );
  OAI22X1 U1235 ( .A(n2930), .B(n2290), .C(n2926), .D(n2289), .Y(n1803) );
  OAI22X1 U1236 ( .A(n2926), .B(n2290), .C(n2930), .D(n2291), .Y(n1804) );
  OAI22X1 U1237 ( .A(n2930), .B(n2292), .C(n2926), .D(n2291), .Y(n1805) );
  OAI22X1 U1238 ( .A(n2926), .B(n2292), .C(n2930), .D(n2293), .Y(n1806) );
  OAI22X1 U1239 ( .A(n2930), .B(n2294), .C(n2926), .D(n2293), .Y(n1807) );
  OAI22X1 U1240 ( .A(n2926), .B(n2294), .C(n2930), .D(n2295), .Y(n1808) );
  OAI22X1 U1241 ( .A(n2930), .B(n2296), .C(n2926), .D(n2295), .Y(n1809) );
  OAI22X1 U1242 ( .A(n2926), .B(n2296), .C(n2930), .D(n2297), .Y(n1810) );
  OAI22X1 U1243 ( .A(n2930), .B(n2298), .C(n2926), .D(n2297), .Y(n1811) );
  OAI22X1 U1244 ( .A(n2926), .B(n2298), .C(n2930), .D(n2299), .Y(n1812) );
  OAI22X1 U1245 ( .A(n2930), .B(n2300), .C(n2926), .D(n2299), .Y(n1813) );
  OAI22X1 U1246 ( .A(n2926), .B(n2300), .C(n2930), .D(n2301), .Y(n1814) );
  OAI22X1 U1247 ( .A(n2930), .B(n2302), .C(n2926), .D(n2301), .Y(n1815) );
  OAI22X1 U1248 ( .A(n2926), .B(n2302), .C(n2930), .D(n2303), .Y(n1816) );
  OAI22X1 U1249 ( .A(n2930), .B(n2304), .C(n2926), .D(n2303), .Y(n1817) );
  XNOR2X1 U1250 ( .A(n3101), .B(n3112), .Y(n2285) );
  XNOR2X1 U1251 ( .A(n3099), .B(n3112), .Y(n2286) );
  XNOR2X1 U1252 ( .A(n2964), .B(n3112), .Y(n2287) );
  XNOR2X1 U1253 ( .A(n3094), .B(n3112), .Y(n2288) );
  XNOR2X1 U1254 ( .A(n3091), .B(n3112), .Y(n2289) );
  XNOR2X1 U1255 ( .A(n3089), .B(n3112), .Y(n2290) );
  XNOR2X1 U1256 ( .A(n3086), .B(n3112), .Y(n2291) );
  XNOR2X1 U1257 ( .A(n3084), .B(n3112), .Y(n2292) );
  XNOR2X1 U1258 ( .A(n3082), .B(n3112), .Y(n2293) );
  XNOR2X1 U1259 ( .A(n3080), .B(n3112), .Y(n2294) );
  XNOR2X1 U1260 ( .A(n3078), .B(n3112), .Y(n2295) );
  XNOR2X1 U1261 ( .A(n3076), .B(n3112), .Y(n2296) );
  XNOR2X1 U1262 ( .A(n3074), .B(n3113), .Y(n2297) );
  XNOR2X1 U1263 ( .A(n3072), .B(n3113), .Y(n2298) );
  XNOR2X1 U1264 ( .A(n2962), .B(n3113), .Y(n2299) );
  XNOR2X1 U1265 ( .A(n3067), .B(n3113), .Y(n2300) );
  XNOR2X1 U1266 ( .A(n3064), .B(n3113), .Y(n2301) );
  XNOR2X1 U1267 ( .A(n3062), .B(n3113), .Y(n2302) );
  XNOR2X1 U1268 ( .A(n437), .B(n3113), .Y(n2303) );
  XNOR2X1 U1269 ( .A(n3055), .B(n3113), .Y(n2304) );
  OAI22X1 U1270 ( .A(n3117), .B(n2928), .C(n2925), .D(n2328), .Y(n1757) );
  OAI22X1 U1271 ( .A(n2928), .B(n2307), .C(n2925), .D(n2306), .Y(n1819) );
  OAI22X1 U1272 ( .A(n2928), .B(n2308), .C(n2925), .D(n2307), .Y(n1820) );
  OAI22X1 U1273 ( .A(n2928), .B(n2309), .C(n2925), .D(n2308), .Y(n1821) );
  OAI22X1 U1274 ( .A(n2925), .B(n2309), .C(n2928), .D(n2310), .Y(n1822) );
  OAI22X1 U1275 ( .A(n2928), .B(n2311), .C(n2925), .D(n2310), .Y(n1823) );
  OAI22X1 U1276 ( .A(n2925), .B(n2311), .C(n2928), .D(n2312), .Y(n1824) );
  OAI22X1 U1277 ( .A(n2928), .B(n2313), .C(n2925), .D(n2312), .Y(n1825) );
  OAI22X1 U1278 ( .A(n2925), .B(n2313), .C(n2928), .D(n2314), .Y(n1826) );
  OAI22X1 U1279 ( .A(n2928), .B(n2315), .C(n2925), .D(n2314), .Y(n1827) );
  OAI22X1 U1280 ( .A(n2925), .B(n2315), .C(n2928), .D(n2316), .Y(n1828) );
  OAI22X1 U1281 ( .A(n2928), .B(n2317), .C(n2925), .D(n2316), .Y(n1829) );
  OAI22X1 U1282 ( .A(n2925), .B(n2317), .C(n2928), .D(n2318), .Y(n1830) );
  OAI22X1 U1283 ( .A(n2928), .B(n2319), .C(n2925), .D(n2318), .Y(n1831) );
  OAI22X1 U1284 ( .A(n2925), .B(n2319), .C(n2928), .D(n2320), .Y(n1832) );
  OAI22X1 U1285 ( .A(n2928), .B(n2321), .C(n2925), .D(n2320), .Y(n1833) );
  OAI22X1 U1286 ( .A(n2925), .B(n2321), .C(n2928), .D(n2322), .Y(n1834) );
  OAI22X1 U1287 ( .A(n2928), .B(n2323), .C(n2925), .D(n2322), .Y(n1835) );
  OAI22X1 U1288 ( .A(n2925), .B(n2323), .C(n2928), .D(n2324), .Y(n1836) );
  OAI22X1 U1289 ( .A(n2928), .B(n2325), .C(n2925), .D(n2324), .Y(n1837) );
  OAI22X1 U1290 ( .A(n2925), .B(n2325), .C(n2928), .D(n2326), .Y(n1838) );
  OAI22X1 U1291 ( .A(n2928), .B(n2327), .C(n2925), .D(n2326), .Y(n1839) );
  XNOR2X1 U1292 ( .A(n3106), .B(n3115), .Y(n2306) );
  XNOR2X1 U1293 ( .A(n3104), .B(n3115), .Y(n2307) );
  XNOR2X1 U1294 ( .A(n3102), .B(n3116), .Y(n2308) );
  XNOR2X1 U1295 ( .A(n3099), .B(n3116), .Y(n2309) );
  XNOR2X1 U1296 ( .A(n2965), .B(n3116), .Y(n2310) );
  XNOR2X1 U1297 ( .A(n3094), .B(n3116), .Y(n2311) );
  XNOR2X1 U1298 ( .A(n3091), .B(n3116), .Y(n2312) );
  XNOR2X1 U1299 ( .A(n3089), .B(n3116), .Y(n2313) );
  XNOR2X1 U1300 ( .A(n3086), .B(n3116), .Y(n2314) );
  XNOR2X1 U1301 ( .A(n3084), .B(n3116), .Y(n2315) );
  XNOR2X1 U1302 ( .A(n3082), .B(n3116), .Y(n2316) );
  XNOR2X1 U1303 ( .A(n3080), .B(n3116), .Y(n2317) );
  XNOR2X1 U1304 ( .A(n3078), .B(n3115), .Y(n2318) );
  XNOR2X1 U1305 ( .A(n3076), .B(n3115), .Y(n2319) );
  XNOR2X1 U1306 ( .A(n3074), .B(n3115), .Y(n2320) );
  XNOR2X1 U1307 ( .A(n3072), .B(n3115), .Y(n2321) );
  XNOR2X1 U1308 ( .A(n2962), .B(n3115), .Y(n2322) );
  XNOR2X1 U1309 ( .A(n3067), .B(n3115), .Y(n2323) );
  XNOR2X1 U1310 ( .A(n3064), .B(n3115), .Y(n2324) );
  XNOR2X1 U1311 ( .A(n3062), .B(n3115), .Y(n2325) );
  XNOR2X1 U1312 ( .A(n437), .B(n3115), .Y(n2326) );
  XNOR2X1 U1313 ( .A(n3055), .B(n3115), .Y(n2327) );
  OAI22X1 U1314 ( .A(n3120), .B(n2929), .C(n3040), .D(n2353), .Y(n1758) );
  OAI22X1 U1315 ( .A(n2929), .B(n2330), .C(n3040), .D(n2329), .Y(n1841) );
  OAI22X1 U1316 ( .A(n3040), .B(n2330), .C(n2929), .D(n2331), .Y(n1842) );
  OAI22X1 U1317 ( .A(n2929), .B(n2332), .C(n3040), .D(n2331), .Y(n1843) );
  OAI22X1 U1318 ( .A(n2929), .B(n2333), .C(n3040), .D(n2332), .Y(n1844) );
  OAI22X1 U1319 ( .A(n2929), .B(n2334), .C(n3040), .D(n2333), .Y(n1845) );
  OAI22X1 U1320 ( .A(n3040), .B(n2334), .C(n2929), .D(n2335), .Y(n1846) );
  OAI22X1 U1321 ( .A(n2929), .B(n2336), .C(n3040), .D(n2335), .Y(n1847) );
  OAI22X1 U1322 ( .A(n3040), .B(n2336), .C(n2929), .D(n2337), .Y(n1848) );
  OAI22X1 U1323 ( .A(n2929), .B(n2338), .C(n3040), .D(n2337), .Y(n1849) );
  OAI22X1 U1324 ( .A(n3040), .B(n2338), .C(n2929), .D(n2339), .Y(n1850) );
  OAI22X1 U1325 ( .A(n2929), .B(n2340), .C(n3040), .D(n2339), .Y(n1851) );
  OAI22X1 U1326 ( .A(n3040), .B(n2340), .C(n2929), .D(n2341), .Y(n1852) );
  OAI22X1 U1327 ( .A(n2929), .B(n2342), .C(n3040), .D(n2341), .Y(n1853) );
  OAI22X1 U1328 ( .A(n3040), .B(n2342), .C(n2929), .D(n2343), .Y(n1854) );
  OAI22X1 U1329 ( .A(n2929), .B(n2344), .C(n3040), .D(n2343), .Y(n1855) );
  OAI22X1 U1330 ( .A(n3040), .B(n2344), .C(n2929), .D(n2345), .Y(n1856) );
  OAI22X1 U1331 ( .A(n2929), .B(n2346), .C(n3040), .D(n2345), .Y(n1857) );
  OAI22X1 U1332 ( .A(n3040), .B(n2346), .C(n2929), .D(n2347), .Y(n1858) );
  OAI22X1 U1333 ( .A(n2929), .B(n2348), .C(n3040), .D(n2347), .Y(n1859) );
  OAI22X1 U1334 ( .A(n3040), .B(n2348), .C(n2929), .D(n2349), .Y(n1860) );
  OAI22X1 U1335 ( .A(n2929), .B(n2350), .C(n3040), .D(n2349), .Y(n1861) );
  OAI22X1 U1336 ( .A(n3040), .B(n2350), .C(n2929), .D(n2351), .Y(n1862) );
  OAI22X1 U1337 ( .A(n2929), .B(n2352), .C(n3040), .D(n2351), .Y(n1863) );
  XNOR2X1 U1338 ( .A(n3110), .B(n3119), .Y(n2329) );
  XNOR2X1 U1340 ( .A(n3106), .B(n3118), .Y(n2331) );
  XNOR2X1 U1341 ( .A(n3104), .B(n3118), .Y(n2332) );
  XNOR2X1 U1342 ( .A(n3101), .B(n3119), .Y(n2333) );
  XNOR2X1 U1343 ( .A(n3099), .B(n3118), .Y(n2334) );
  XNOR2X1 U1344 ( .A(n2976), .B(n3119), .Y(n2335) );
  XNOR2X1 U1345 ( .A(n3094), .B(n3119), .Y(n2336) );
  XNOR2X1 U1346 ( .A(n3091), .B(n3119), .Y(n2337) );
  XNOR2X1 U1347 ( .A(n3089), .B(n3119), .Y(n2338) );
  XNOR2X1 U1348 ( .A(n3086), .B(n3119), .Y(n2339) );
  XNOR2X1 U1349 ( .A(n3084), .B(n3119), .Y(n2340) );
  XNOR2X1 U1350 ( .A(n3082), .B(n3119), .Y(n2341) );
  XNOR2X1 U1351 ( .A(n3080), .B(n3119), .Y(n2342) );
  XNOR2X1 U1352 ( .A(n3078), .B(n3119), .Y(n2343) );
  XNOR2X1 U1353 ( .A(n3076), .B(n3118), .Y(n2344) );
  XNOR2X1 U1354 ( .A(n3074), .B(n3118), .Y(n2345) );
  XNOR2X1 U1355 ( .A(n3072), .B(n3118), .Y(n2346) );
  XNOR2X1 U1356 ( .A(n3070), .B(n3118), .Y(n2347) );
  XNOR2X1 U1357 ( .A(n3067), .B(n3118), .Y(n2348) );
  XNOR2X1 U1358 ( .A(n3064), .B(n3118), .Y(n2349) );
  XNOR2X1 U1359 ( .A(n3061), .B(n3118), .Y(n2350) );
  XNOR2X1 U1360 ( .A(n437), .B(n3118), .Y(n2351) );
  XNOR2X1 U1361 ( .A(n3055), .B(n3118), .Y(n2352) );
  OAI22X1 U1362 ( .A(n3124), .B(n2924), .C(n3041), .D(n2380), .Y(n1759) );
  OAI22X1 U1363 ( .A(n2924), .B(n2355), .C(n3041), .D(n2354), .Y(n1865) );
  OAI22X1 U1364 ( .A(n2924), .B(n2356), .C(n3041), .D(n2355), .Y(n1866) );
  OAI22X1 U1365 ( .A(n2924), .B(n2357), .C(n3041), .D(n2356), .Y(n1867) );
  OAI22X1 U1366 ( .A(n3041), .B(n2357), .C(n2924), .D(n2358), .Y(n1868) );
  OAI22X1 U1367 ( .A(n2924), .B(n2359), .C(n3041), .D(n2358), .Y(n1869) );
  OAI22X1 U1368 ( .A(n2924), .B(n2360), .C(n3041), .D(n2359), .Y(n1870) );
  OAI22X1 U1369 ( .A(n2924), .B(n2361), .C(n3041), .D(n2360), .Y(n1871) );
  OAI22X1 U1370 ( .A(n3041), .B(n2361), .C(n2924), .D(n2362), .Y(n1872) );
  OAI22X1 U1371 ( .A(n2924), .B(n2363), .C(n3041), .D(n2362), .Y(n1873) );
  OAI22X1 U1372 ( .A(n3041), .B(n2363), .C(n2924), .D(n2364), .Y(n1874) );
  OAI22X1 U1373 ( .A(n2924), .B(n2365), .C(n3041), .D(n2364), .Y(n1875) );
  OAI22X1 U1374 ( .A(n3041), .B(n2365), .C(n2924), .D(n2366), .Y(n1876) );
  OAI22X1 U1375 ( .A(n2924), .B(n2367), .C(n3041), .D(n2366), .Y(n1877) );
  OAI22X1 U1376 ( .A(n3041), .B(n2367), .C(n2924), .D(n2368), .Y(n1878) );
  OAI22X1 U1377 ( .A(n2924), .B(n2369), .C(n3041), .D(n2368), .Y(n1879) );
  OAI22X1 U1378 ( .A(n3041), .B(n2369), .C(n2924), .D(n2370), .Y(n1880) );
  OAI22X1 U1379 ( .A(n2924), .B(n2371), .C(n3041), .D(n2370), .Y(n1881) );
  OAI22X1 U1380 ( .A(n3041), .B(n2371), .C(n2924), .D(n2372), .Y(n1882) );
  OAI22X1 U1381 ( .A(n2924), .B(n2373), .C(n3041), .D(n2372), .Y(n1883) );
  OAI22X1 U1382 ( .A(n3041), .B(n2373), .C(n2924), .D(n2374), .Y(n1884) );
  OAI22X1 U1383 ( .A(n2924), .B(n2375), .C(n3041), .D(n2374), .Y(n1885) );
  OAI22X1 U1384 ( .A(n3041), .B(n2375), .C(n2924), .D(n2376), .Y(n1886) );
  OAI22X1 U1385 ( .A(n2924), .B(n2377), .C(n3041), .D(n2376), .Y(n1887) );
  OAI22X1 U1386 ( .A(n3041), .B(n2377), .C(n2924), .D(n2378), .Y(n1888) );
  OAI22X1 U1387 ( .A(n2924), .B(n2379), .C(n3041), .D(n2378), .Y(n1889) );
  XNOR2X1 U1388 ( .A(n485), .B(n3122), .Y(n2354) );
  XNOR2X1 U1389 ( .A(n3028), .B(n3121), .Y(n2355) );
  XNOR2X1 U1390 ( .A(n3110), .B(n3121), .Y(n2356) );
  XNOR2X1 U1391 ( .A(n3108), .B(n3121), .Y(n2357) );
  XNOR2X1 U1392 ( .A(n3106), .B(n3121), .Y(n2358) );
  XNOR2X1 U1393 ( .A(n3104), .B(n3121), .Y(n2359) );
  XNOR2X1 U1394 ( .A(n3102), .B(n3122), .Y(n2360) );
  XNOR2X1 U1395 ( .A(n471), .B(n3123), .Y(n2361) );
  XNOR2X1 U1396 ( .A(n3097), .B(n3123), .Y(n2362) );
  XNOR2X1 U1397 ( .A(n467), .B(n3122), .Y(n2363) );
  XNOR2X1 U1398 ( .A(n3091), .B(n3122), .Y(n2364) );
  XNOR2X1 U1399 ( .A(n3089), .B(n3122), .Y(n2365) );
  XNOR2X1 U1400 ( .A(n3086), .B(n3122), .Y(n2366) );
  XNOR2X1 U1401 ( .A(n3084), .B(n3122), .Y(n2367) );
  XNOR2X1 U1402 ( .A(n3082), .B(n3122), .Y(n2368) );
  XNOR2X1 U1403 ( .A(n3080), .B(n3122), .Y(n2369) );
  XNOR2X1 U1404 ( .A(n3078), .B(n3122), .Y(n2370) );
  XNOR2X1 U1405 ( .A(n3076), .B(n3121), .Y(n2371) );
  XNOR2X1 U1406 ( .A(n3074), .B(n3121), .Y(n2372) );
  XNOR2X1 U1407 ( .A(n3072), .B(n3121), .Y(n2373) );
  XNOR2X1 U1408 ( .A(n3070), .B(n3121), .Y(n2374) );
  XNOR2X1 U1409 ( .A(n3067), .B(n3121), .Y(n2375) );
  XNOR2X1 U1410 ( .A(n3064), .B(n3121), .Y(n2376) );
  XNOR2X1 U1411 ( .A(n3062), .B(n3121), .Y(n2377) );
  XNOR2X1 U1412 ( .A(n437), .B(n3122), .Y(n2378) );
  XNOR2X1 U1413 ( .A(n3055), .B(n3122), .Y(n2379) );
  OAI22X1 U1414 ( .A(n3127), .B(n2923), .C(n3042), .D(n2409), .Y(n1760) );
  OAI22X1 U1415 ( .A(n2923), .B(n2382), .C(n3042), .D(n2381), .Y(n1891) );
  OAI22X1 U1416 ( .A(n3042), .B(n2382), .C(n2923), .D(n2383), .Y(n1892) );
  OAI22X1 U1417 ( .A(n2923), .B(n2384), .C(n3042), .D(n2383), .Y(n1893) );
  OAI22X1 U1418 ( .A(n2923), .B(n2385), .C(n3042), .D(n2384), .Y(n1894) );
  OAI22X1 U1419 ( .A(n2923), .B(n2386), .C(n3042), .D(n2385), .Y(n1895) );
  OAI22X1 U1420 ( .A(n3042), .B(n2386), .C(n2923), .D(n2387), .Y(n1896) );
  OAI22X1 U1421 ( .A(n2923), .B(n2388), .C(n3042), .D(n2387), .Y(n1897) );
  OAI22X1 U1422 ( .A(n2923), .B(n2389), .C(n3042), .D(n2388), .Y(n1898) );
  OAI22X1 U1423 ( .A(n2923), .B(n2390), .C(n3042), .D(n2389), .Y(n1899) );
  OAI22X1 U1424 ( .A(n3042), .B(n2390), .C(n2923), .D(n2391), .Y(n1900) );
  OAI22X1 U1425 ( .A(n2923), .B(n2392), .C(n3042), .D(n2391), .Y(n1901) );
  OAI22X1 U1426 ( .A(n3042), .B(n2392), .C(n2923), .D(n2393), .Y(n1902) );
  OAI22X1 U1427 ( .A(n2923), .B(n2394), .C(n3042), .D(n2393), .Y(n1903) );
  OAI22X1 U1428 ( .A(n3042), .B(n2394), .C(n2923), .D(n2395), .Y(n1904) );
  OAI22X1 U1429 ( .A(n2923), .B(n2396), .C(n3042), .D(n2395), .Y(n1905) );
  OAI22X1 U1430 ( .A(n3042), .B(n2396), .C(n2923), .D(n2397), .Y(n1906) );
  OAI22X1 U1431 ( .A(n2923), .B(n2398), .C(n3042), .D(n2397), .Y(n1907) );
  OAI22X1 U1432 ( .A(n3042), .B(n2398), .C(n2923), .D(n2399), .Y(n1908) );
  OAI22X1 U1433 ( .A(n2923), .B(n2400), .C(n3042), .D(n2399), .Y(n1909) );
  OAI22X1 U1434 ( .A(n3042), .B(n2400), .C(n2923), .D(n2401), .Y(n1910) );
  OAI22X1 U1435 ( .A(n2923), .B(n2402), .C(n3042), .D(n2401), .Y(n1911) );
  OAI22X1 U1436 ( .A(n3042), .B(n2402), .C(n2923), .D(n2403), .Y(n1912) );
  OAI22X1 U1437 ( .A(n2923), .B(n2404), .C(n3042), .D(n2403), .Y(n1913) );
  OAI22X1 U1438 ( .A(n3042), .B(n2404), .C(n2923), .D(n2405), .Y(n1914) );
  OAI22X1 U1439 ( .A(n2923), .B(n2406), .C(n3042), .D(n2405), .Y(n1915) );
  OAI22X1 U1440 ( .A(n3042), .B(n2406), .C(n2923), .D(n2407), .Y(n1916) );
  OAI22X1 U1441 ( .A(n2923), .B(n2408), .C(n3042), .D(n2407), .Y(n1917) );
  XNOR2X1 U1442 ( .A(n489), .B(n3125), .Y(n2381) );
  XNOR2X1 U1443 ( .A(n487), .B(n3125), .Y(n2382) );
  XNOR2X1 U1444 ( .A(n485), .B(n3125), .Y(n2383) );
  XNOR2X1 U1445 ( .A(n3029), .B(n3125), .Y(n2384) );
  XNOR2X1 U1446 ( .A(n3110), .B(n3125), .Y(n2385) );
  XNOR2X1 U1447 ( .A(n3108), .B(n3125), .Y(n2386) );
  XNOR2X1 U1448 ( .A(n3106), .B(n3125), .Y(n2387) );
  XNOR2X1 U1449 ( .A(n3104), .B(n3125), .Y(n2388) );
  XNOR2X1 U1450 ( .A(n3101), .B(n3125), .Y(n2389) );
  XNOR2X1 U1451 ( .A(n3099), .B(n3126), .Y(n2390) );
  XNOR2X1 U1452 ( .A(n2964), .B(n3126), .Y(n2391) );
  XNOR2X1 U1453 ( .A(n467), .B(n3126), .Y(n2392) );
  XNOR2X1 U1454 ( .A(n3091), .B(n3126), .Y(n2393) );
  XNOR2X1 U1455 ( .A(n3089), .B(n3125), .Y(n2394) );
  XNOR2X1 U1456 ( .A(n3086), .B(n3125), .Y(n2395) );
  XNOR2X1 U1457 ( .A(n3084), .B(n3125), .Y(n2396) );
  XNOR2X1 U1458 ( .A(n3082), .B(n3125), .Y(n2397) );
  XNOR2X1 U1459 ( .A(n3080), .B(n3125), .Y(n2398) );
  XNOR2X1 U1460 ( .A(n3078), .B(n3125), .Y(n2399) );
  XNOR2X1 U1461 ( .A(n3076), .B(n3125), .Y(n2400) );
  XNOR2X1 U1462 ( .A(n3074), .B(n3125), .Y(n2401) );
  XNOR2X1 U1463 ( .A(n3072), .B(n3125), .Y(n2402) );
  XNOR2X1 U1464 ( .A(n2963), .B(n3125), .Y(n2403) );
  XNOR2X1 U1465 ( .A(n3067), .B(n3125), .Y(n2404) );
  XNOR2X1 U1466 ( .A(n3064), .B(n3125), .Y(n2405) );
  XNOR2X1 U1467 ( .A(n3062), .B(n3125), .Y(n2406) );
  XNOR2X1 U1468 ( .A(n437), .B(n3125), .Y(n2407) );
  XNOR2X1 U1469 ( .A(n3056), .B(n3125), .Y(n2408) );
  OAI22X1 U1470 ( .A(n3130), .B(n3030), .C(n3043), .D(n2440), .Y(n1761) );
  OAI22X1 U1471 ( .A(n3043), .B(n2410), .C(n3030), .D(n2411), .Y(n1919) );
  OAI22X1 U1472 ( .A(n3043), .B(n2411), .C(n3030), .D(n2412), .Y(n1920) );
  OAI22X1 U1473 ( .A(n3030), .B(n2413), .C(n3043), .D(n2412), .Y(n1921) );
  OAI22X1 U1474 ( .A(n3043), .B(n2413), .C(n3030), .D(n2414), .Y(n1922) );
  OAI22X1 U1475 ( .A(n3030), .B(n2415), .C(n3043), .D(n2414), .Y(n1923) );
  OAI22X1 U1476 ( .A(n3030), .B(n2416), .C(n3043), .D(n2415), .Y(n1924) );
  OAI22X1 U1477 ( .A(n3030), .B(n2417), .C(n3043), .D(n2416), .Y(n1925) );
  OAI22X1 U1478 ( .A(n3043), .B(n2417), .C(n3030), .D(n2418), .Y(n1926) );
  OAI22X1 U1479 ( .A(n3030), .B(n2419), .C(n3043), .D(n2418), .Y(n1927) );
  OAI22X1 U1480 ( .A(n3030), .B(n2420), .C(n3043), .D(n2419), .Y(n1928) );
  OAI22X1 U1481 ( .A(n3030), .B(n2421), .C(n3043), .D(n2420), .Y(n1929) );
  OAI22X1 U1482 ( .A(n3043), .B(n2421), .C(n3030), .D(n2422), .Y(n1930) );
  OAI22X1 U1483 ( .A(n3030), .B(n2423), .C(n3043), .D(n2422), .Y(n1931) );
  OAI22X1 U1484 ( .A(n3043), .B(n2423), .C(n3030), .D(n2424), .Y(n1932) );
  OAI22X1 U1485 ( .A(n3030), .B(n2425), .C(n3043), .D(n2424), .Y(n1933) );
  OAI22X1 U1486 ( .A(n3043), .B(n2425), .C(n3030), .D(n2426), .Y(n1934) );
  OAI22X1 U1487 ( .A(n3030), .B(n2427), .C(n3043), .D(n2426), .Y(n1935) );
  OAI22X1 U1488 ( .A(n3043), .B(n2427), .C(n3030), .D(n2428), .Y(n1936) );
  OAI22X1 U1489 ( .A(n3030), .B(n2429), .C(n3043), .D(n2428), .Y(n1937) );
  OAI22X1 U1490 ( .A(n3043), .B(n2429), .C(n3030), .D(n2430), .Y(n1938) );
  OAI22X1 U1491 ( .A(n3030), .B(n2431), .C(n3043), .D(n2430), .Y(n1939) );
  OAI22X1 U1492 ( .A(n3043), .B(n2431), .C(n3030), .D(n2432), .Y(n1940) );
  OAI22X1 U1493 ( .A(n3030), .B(n2433), .C(n3043), .D(n2432), .Y(n1941) );
  OAI22X1 U1494 ( .A(n3043), .B(n2433), .C(n3030), .D(n2434), .Y(n1942) );
  OAI22X1 U1495 ( .A(n3030), .B(n2435), .C(n3043), .D(n2434), .Y(n1943) );
  OAI22X1 U1496 ( .A(n3043), .B(n2435), .C(n3030), .D(n2436), .Y(n1944) );
  OAI22X1 U1497 ( .A(n3030), .B(n2437), .C(n3043), .D(n2436), .Y(n1945) );
  OAI22X1 U1498 ( .A(n3043), .B(n2437), .C(n3030), .D(n2438), .Y(n1946) );
  OAI22X1 U1499 ( .A(n3030), .B(n2439), .C(n3043), .D(n2438), .Y(n1947) );
  XNOR2X1 U1500 ( .A(n493), .B(n3128), .Y(n2410) );
  XNOR2X1 U1501 ( .A(n491), .B(n3128), .Y(n2411) );
  XNOR2X1 U1502 ( .A(n489), .B(n3128), .Y(n2412) );
  XNOR2X1 U1503 ( .A(n487), .B(n3128), .Y(n2413) );
  XNOR2X1 U1504 ( .A(n485), .B(n3128), .Y(n2414) );
  XNOR2X1 U1505 ( .A(n3028), .B(n3128), .Y(n2415) );
  XNOR2X1 U1506 ( .A(n3110), .B(n3128), .Y(n2416) );
  XNOR2X1 U1507 ( .A(n3108), .B(n3128), .Y(n2417) );
  XNOR2X1 U1508 ( .A(n3106), .B(n3128), .Y(n2418) );
  XNOR2X1 U1509 ( .A(n3104), .B(n3128), .Y(n2419) );
  XNOR2X1 U1510 ( .A(n3101), .B(n3129), .Y(n2420) );
  XNOR2X1 U1511 ( .A(n471), .B(n3129), .Y(n2421) );
  XNOR2X1 U1512 ( .A(n2965), .B(n3129), .Y(n2422) );
  XNOR2X1 U1513 ( .A(n467), .B(n3129), .Y(n2423) );
  XNOR2X1 U1514 ( .A(n3091), .B(n3129), .Y(n2424) );
  XNOR2X1 U1515 ( .A(n3089), .B(n3129), .Y(n2425) );
  XNOR2X1 U1516 ( .A(n3086), .B(n3128), .Y(n2426) );
  XNOR2X1 U1517 ( .A(n3084), .B(n3128), .Y(n2427) );
  XNOR2X1 U1518 ( .A(n3082), .B(n3128), .Y(n2428) );
  XNOR2X1 U1519 ( .A(n3080), .B(n3128), .Y(n2429) );
  XNOR2X1 U1520 ( .A(n3078), .B(n3128), .Y(n2430) );
  XNOR2X1 U1521 ( .A(n3076), .B(n3128), .Y(n2431) );
  XNOR2X1 U1522 ( .A(n3074), .B(n3128), .Y(n2432) );
  XNOR2X1 U1523 ( .A(n3072), .B(n3128), .Y(n2433) );
  XNOR2X1 U1524 ( .A(n2963), .B(n3128), .Y(n2434) );
  XNOR2X1 U1525 ( .A(n3067), .B(n3128), .Y(n2435) );
  XNOR2X1 U1526 ( .A(n3064), .B(n3128), .Y(n2436) );
  XNOR2X1 U1527 ( .A(n3061), .B(n3128), .Y(n2437) );
  XNOR2X1 U1528 ( .A(n437), .B(n3128), .Y(n2438) );
  XNOR2X1 U1529 ( .A(n3056), .B(n3128), .Y(n2439) );
  OAI22X1 U1530 ( .A(n3133), .B(n3031), .C(n3044), .D(n2473), .Y(n1762) );
  OAI22X1 U1531 ( .A(n3044), .B(n2441), .C(n3031), .D(n2442), .Y(n1949) );
  OAI22X1 U1532 ( .A(n3031), .B(n2443), .C(n3044), .D(n2442), .Y(n1950) );
  OAI22X1 U1533 ( .A(n3044), .B(n2443), .C(n3031), .D(n2444), .Y(n1951) );
  OAI22X1 U1534 ( .A(n3044), .B(n2444), .C(n3031), .D(n2445), .Y(n1952) );
  OAI22X1 U1535 ( .A(n3031), .B(n2446), .C(n3044), .D(n2445), .Y(n1953) );
  OAI22X1 U1536 ( .A(n3044), .B(n2446), .C(n3031), .D(n2447), .Y(n1954) );
  OAI22X1 U1537 ( .A(n3031), .B(n2448), .C(n3044), .D(n2447), .Y(n1955) );
  OAI22X1 U1538 ( .A(n3031), .B(n2449), .C(n3044), .D(n2448), .Y(n1956) );
  OAI22X1 U1539 ( .A(n3031), .B(n2450), .C(n3044), .D(n2449), .Y(n1957) );
  OAI22X1 U1540 ( .A(n3044), .B(n2450), .C(n3031), .D(n2451), .Y(n1958) );
  OAI22X1 U1541 ( .A(n3031), .B(n2452), .C(n3044), .D(n2451), .Y(n1959) );
  OAI22X1 U1542 ( .A(n3031), .B(n2453), .C(n3044), .D(n2452), .Y(n1960) );
  OAI22X1 U1543 ( .A(n3031), .B(n2454), .C(n3044), .D(n2453), .Y(n1961) );
  OAI22X1 U1544 ( .A(n3044), .B(n2454), .C(n3031), .D(n2455), .Y(n1962) );
  OAI22X1 U1545 ( .A(n3031), .B(n2456), .C(n3044), .D(n2455), .Y(n1963) );
  OAI22X1 U1546 ( .A(n3044), .B(n2456), .C(n3031), .D(n2457), .Y(n1964) );
  OAI22X1 U1547 ( .A(n3031), .B(n2458), .C(n3044), .D(n2457), .Y(n1965) );
  OAI22X1 U1548 ( .A(n3044), .B(n2458), .C(n3031), .D(n2459), .Y(n1966) );
  OAI22X1 U1549 ( .A(n3031), .B(n2460), .C(n3044), .D(n2459), .Y(n1967) );
  OAI22X1 U1550 ( .A(n3044), .B(n2460), .C(n3031), .D(n2461), .Y(n1968) );
  OAI22X1 U1551 ( .A(n3031), .B(n2462), .C(n3044), .D(n2461), .Y(n1969) );
  OAI22X1 U1552 ( .A(n3044), .B(n2462), .C(n3031), .D(n2463), .Y(n1970) );
  OAI22X1 U1553 ( .A(n3031), .B(n2464), .C(n3044), .D(n2463), .Y(n1971) );
  OAI22X1 U1554 ( .A(n3044), .B(n2464), .C(n3031), .D(n2465), .Y(n1972) );
  OAI22X1 U1555 ( .A(n3031), .B(n2466), .C(n3044), .D(n2465), .Y(n1973) );
  OAI22X1 U1556 ( .A(n3044), .B(n2466), .C(n3031), .D(n2467), .Y(n1974) );
  OAI22X1 U1557 ( .A(n3031), .B(n2468), .C(n3044), .D(n2467), .Y(n1975) );
  OAI22X1 U1558 ( .A(n3044), .B(n2468), .C(n3031), .D(n2469), .Y(n1976) );
  OAI22X1 U1559 ( .A(n3031), .B(n2470), .C(n3044), .D(n2469), .Y(n1977) );
  OAI22X1 U1560 ( .A(n3044), .B(n2470), .C(n3031), .D(n2471), .Y(n1978) );
  OAI22X1 U1561 ( .A(n3031), .B(n2472), .C(n3044), .D(n2471), .Y(n1979) );
  XNOR2X1 U1562 ( .A(n497), .B(n3132), .Y(n2441) );
  XNOR2X1 U1563 ( .A(n495), .B(n3131), .Y(n2442) );
  XNOR2X1 U1564 ( .A(n493), .B(n3131), .Y(n2443) );
  XNOR2X1 U1565 ( .A(n491), .B(n3131), .Y(n2444) );
  XNOR2X1 U1566 ( .A(n489), .B(n3131), .Y(n2445) );
  XNOR2X1 U1567 ( .A(n487), .B(n3131), .Y(n2446) );
  XNOR2X1 U1568 ( .A(n485), .B(n3131), .Y(n2447) );
  XNOR2X1 U1569 ( .A(n3029), .B(n3131), .Y(n2448) );
  XNOR2X1 U1570 ( .A(n3110), .B(n3131), .Y(n2449) );
  XNOR2X1 U1571 ( .A(n3108), .B(n3131), .Y(n2450) );
  XNOR2X1 U1572 ( .A(n3106), .B(n3131), .Y(n2451) );
  XNOR2X1 U1573 ( .A(n3104), .B(n3131), .Y(n2452) );
  XNOR2X1 U1574 ( .A(n3101), .B(n3131), .Y(n2453) );
  XNOR2X1 U1575 ( .A(n471), .B(n3131), .Y(n2454) );
  XNOR2X1 U1576 ( .A(n2965), .B(n3131), .Y(n2455) );
  XNOR2X1 U1577 ( .A(n467), .B(n3131), .Y(n2456) );
  XNOR2X1 U1578 ( .A(n3091), .B(n3131), .Y(n2457) );
  XNOR2X1 U1579 ( .A(n3089), .B(n3131), .Y(n2458) );
  XNOR2X1 U1580 ( .A(n3086), .B(n3131), .Y(n2459) );
  XNOR2X1 U1581 ( .A(n3084), .B(n3131), .Y(n2460) );
  XNOR2X1 U1582 ( .A(n3082), .B(n3131), .Y(n2461) );
  XNOR2X1 U1583 ( .A(n3080), .B(n3132), .Y(n2462) );
  XNOR2X1 U1584 ( .A(n3078), .B(n3132), .Y(n2463) );
  XNOR2X1 U1585 ( .A(n3076), .B(n3131), .Y(n2464) );
  XNOR2X1 U1586 ( .A(n3074), .B(n3132), .Y(n2465) );
  XNOR2X1 U1587 ( .A(n3072), .B(n3132), .Y(n2466) );
  XNOR2X1 U1588 ( .A(n3069), .B(n3132), .Y(n2467) );
  XNOR2X1 U1589 ( .A(n3067), .B(n3132), .Y(n2468) );
  XNOR2X1 U1590 ( .A(n3064), .B(n3132), .Y(n2469) );
  XNOR2X1 U1591 ( .A(n3061), .B(n3132), .Y(n2470) );
  XNOR2X1 U1592 ( .A(n437), .B(n3132), .Y(n2471) );
  XNOR2X1 U1593 ( .A(n3056), .B(n3132), .Y(n2472) );
  OAI22X1 U1594 ( .A(n3136), .B(n3032), .C(n3045), .D(n2506), .Y(n1763) );
  OAI22X1 U1595 ( .A(n3136), .B(n3045), .C(n3032), .D(n2474), .Y(n1982) );
  OAI22X1 U1596 ( .A(n3045), .B(n2474), .C(n3032), .D(n2475), .Y(n1983) );
  OAI22X1 U1597 ( .A(n3032), .B(n2476), .C(n3045), .D(n2475), .Y(n1984) );
  OAI22X1 U1598 ( .A(n3045), .B(n2476), .C(n3032), .D(n2477), .Y(n1985) );
  OAI22X1 U1599 ( .A(n3045), .B(n2477), .C(n3032), .D(n2478), .Y(n1986) );
  OAI22X1 U1600 ( .A(n3032), .B(n2479), .C(n3045), .D(n2478), .Y(n1987) );
  OAI22X1 U1601 ( .A(n3045), .B(n2479), .C(n3032), .D(n2480), .Y(n1988) );
  OAI22X1 U1602 ( .A(n3032), .B(n2481), .C(n3045), .D(n2480), .Y(n1989) );
  OAI22X1 U1603 ( .A(n3032), .B(n2482), .C(n3045), .D(n2481), .Y(n1990) );
  OAI22X1 U1604 ( .A(n3032), .B(n2483), .C(n3045), .D(n2482), .Y(n1991) );
  OAI22X1 U1605 ( .A(n3045), .B(n2483), .C(n3032), .D(n2484), .Y(n1992) );
  OAI22X1 U1606 ( .A(n3032), .B(n2485), .C(n3045), .D(n2484), .Y(n1993) );
  OAI22X1 U1607 ( .A(n3032), .B(n2486), .C(n3045), .D(n2485), .Y(n1994) );
  OAI22X1 U1608 ( .A(n3032), .B(n2487), .C(n3045), .D(n2486), .Y(n1995) );
  OAI22X1 U1609 ( .A(n3045), .B(n2487), .C(n3032), .D(n2488), .Y(n1996) );
  OAI22X1 U1610 ( .A(n3032), .B(n2489), .C(n3045), .D(n2488), .Y(n1997) );
  OAI22X1 U1611 ( .A(n3045), .B(n2489), .C(n3032), .D(n2490), .Y(n1998) );
  OAI22X1 U1612 ( .A(n3032), .B(n2491), .C(n3045), .D(n2490), .Y(n1999) );
  OAI22X1 U1613 ( .A(n3045), .B(n2491), .C(n3032), .D(n2492), .Y(n2000) );
  OAI22X1 U1614 ( .A(n3032), .B(n2493), .C(n3045), .D(n2492), .Y(n2001) );
  OAI22X1 U1615 ( .A(n3045), .B(n2493), .C(n3032), .D(n2494), .Y(n2002) );
  OAI22X1 U1616 ( .A(n3032), .B(n2495), .C(n3045), .D(n2494), .Y(n2003) );
  OAI22X1 U1617 ( .A(n3045), .B(n2495), .C(n3032), .D(n2496), .Y(n2004) );
  OAI22X1 U1618 ( .A(n3032), .B(n2497), .C(n3045), .D(n2496), .Y(n2005) );
  OAI22X1 U1619 ( .A(n3045), .B(n2497), .C(n3032), .D(n2498), .Y(n2006) );
  OAI22X1 U1620 ( .A(n3032), .B(n2499), .C(n3045), .D(n2498), .Y(n2007) );
  OAI22X1 U1621 ( .A(n3045), .B(n2499), .C(n3032), .D(n2500), .Y(n2008) );
  OAI22X1 U1622 ( .A(n3032), .B(n2501), .C(n3045), .D(n2500), .Y(n2009) );
  OAI22X1 U1623 ( .A(n3045), .B(n2501), .C(n3032), .D(n2502), .Y(n2010) );
  OAI22X1 U1624 ( .A(n3032), .B(n2503), .C(n3045), .D(n2502), .Y(n2011) );
  OAI22X1 U1625 ( .A(n3045), .B(n2503), .C(n3032), .D(n2504), .Y(n2012) );
  OAI22X1 U1626 ( .A(n3032), .B(n2505), .C(n3045), .D(n2504), .Y(n2013) );
  XNOR2X1 U1627 ( .A(n497), .B(n3134), .Y(n2474) );
  XNOR2X1 U1628 ( .A(n495), .B(n3134), .Y(n2475) );
  XNOR2X1 U1629 ( .A(n493), .B(n3134), .Y(n2476) );
  XNOR2X1 U1630 ( .A(n491), .B(n3134), .Y(n2477) );
  XNOR2X1 U1631 ( .A(n489), .B(n3134), .Y(n2478) );
  XNOR2X1 U1632 ( .A(n487), .B(n3134), .Y(n2479) );
  XNOR2X1 U1633 ( .A(n485), .B(n3134), .Y(n2480) );
  XNOR2X1 U1634 ( .A(n3029), .B(n3134), .Y(n2481) );
  XNOR2X1 U1635 ( .A(n3110), .B(n3134), .Y(n2482) );
  XNOR2X1 U1636 ( .A(n3108), .B(n3134), .Y(n2483) );
  XNOR2X1 U1637 ( .A(n3106), .B(n3134), .Y(n2484) );
  XNOR2X1 U1638 ( .A(n3104), .B(n3134), .Y(n2485) );
  XNOR2X1 U1639 ( .A(n3102), .B(n3135), .Y(n2486) );
  XNOR2X1 U1640 ( .A(n471), .B(n3135), .Y(n2487) );
  XNOR2X1 U1641 ( .A(n3097), .B(n3135), .Y(n2488) );
  XNOR2X1 U1642 ( .A(n467), .B(n3135), .Y(n2489) );
  XNOR2X1 U1643 ( .A(n3092), .B(n3135), .Y(n2490) );
  XNOR2X1 U1644 ( .A(n3089), .B(n3135), .Y(n2491) );
  XNOR2X1 U1645 ( .A(n3087), .B(n3135), .Y(n2492) );
  XNOR2X1 U1646 ( .A(n2968), .B(n3134), .Y(n2493) );
  XNOR2X1 U1647 ( .A(n2960), .B(n3135), .Y(n2494) );
  XNOR2X1 U1648 ( .A(n2967), .B(n3134), .Y(n2495) );
  XNOR2X1 U1649 ( .A(n2961), .B(n3134), .Y(n2496) );
  XNOR2X1 U1650 ( .A(n3076), .B(n3134), .Y(n2497) );
  XNOR2X1 U1651 ( .A(n2974), .B(n3134), .Y(n2498) );
  XNOR2X1 U1652 ( .A(n2975), .B(n3134), .Y(n2499) );
  XNOR2X1 U1653 ( .A(n3069), .B(n3134), .Y(n2500) );
  XNOR2X1 U1654 ( .A(n3067), .B(n3134), .Y(n2501) );
  XNOR2X1 U1655 ( .A(n2973), .B(n3134), .Y(n2502) );
  XNOR2X1 U1656 ( .A(n3061), .B(n3134), .Y(n2503) );
  XNOR2X1 U1657 ( .A(n437), .B(n3134), .Y(n2504) );
  XNOR2X1 U1658 ( .A(n3056), .B(n3134), .Y(n2505) );
  OAI22X1 U1659 ( .A(n3139), .B(n3033), .C(n3046), .D(n2539), .Y(n1764) );
  OAI22X1 U1660 ( .A(n3139), .B(n3046), .C(n3033), .D(n2507), .Y(n2016) );
  OAI22X1 U1661 ( .A(n3046), .B(n2507), .C(n3033), .D(n2508), .Y(n2017) );
  OAI22X1 U1662 ( .A(n3033), .B(n2509), .C(n3046), .D(n2508), .Y(n2018) );
  OAI22X1 U1663 ( .A(n3046), .B(n2509), .C(n3033), .D(n2510), .Y(n2019) );
  OAI22X1 U1664 ( .A(n3046), .B(n2510), .C(n3033), .D(n2511), .Y(n2020) );
  OAI22X1 U1665 ( .A(n3033), .B(n2512), .C(n3046), .D(n2511), .Y(n2021) );
  OAI22X1 U1666 ( .A(n3046), .B(n2512), .C(n3033), .D(n2513), .Y(n2022) );
  OAI22X1 U1667 ( .A(n3033), .B(n2514), .C(n3046), .D(n2513), .Y(n2023) );
  OAI22X1 U1668 ( .A(n3033), .B(n2515), .C(n3046), .D(n2514), .Y(n2024) );
  OAI22X1 U1669 ( .A(n3033), .B(n2516), .C(n3046), .D(n2515), .Y(n2025) );
  OAI22X1 U1670 ( .A(n3046), .B(n2516), .C(n3033), .D(n2517), .Y(n2026) );
  OAI22X1 U1671 ( .A(n3033), .B(n2518), .C(n3046), .D(n2517), .Y(n2027) );
  OAI22X1 U1672 ( .A(n3033), .B(n2519), .C(n3046), .D(n2518), .Y(n2028) );
  OAI22X1 U1673 ( .A(n3033), .B(n2520), .C(n3046), .D(n2519), .Y(n2029) );
  OAI22X1 U1674 ( .A(n3046), .B(n2520), .C(n3033), .D(n2521), .Y(n2030) );
  OAI22X1 U1675 ( .A(n3033), .B(n2522), .C(n3046), .D(n2521), .Y(n2031) );
  OAI22X1 U1676 ( .A(n3046), .B(n2522), .C(n3033), .D(n2523), .Y(n2032) );
  OAI22X1 U1677 ( .A(n3033), .B(n2524), .C(n3046), .D(n2523), .Y(n2033) );
  OAI22X1 U1678 ( .A(n3046), .B(n2524), .C(n3033), .D(n2525), .Y(n2034) );
  OAI22X1 U1679 ( .A(n3033), .B(n2526), .C(n3046), .D(n2525), .Y(n2035) );
  OAI22X1 U1680 ( .A(n3046), .B(n2526), .C(n3033), .D(n2527), .Y(n2036) );
  OAI22X1 U1681 ( .A(n3033), .B(n2528), .C(n3046), .D(n2527), .Y(n2037) );
  OAI22X1 U1682 ( .A(n3046), .B(n2528), .C(n3033), .D(n2529), .Y(n2038) );
  OAI22X1 U1683 ( .A(n3033), .B(n2530), .C(n3046), .D(n2529), .Y(n2039) );
  OAI22X1 U1684 ( .A(n3046), .B(n2530), .C(n3033), .D(n2531), .Y(n2040) );
  OAI22X1 U1685 ( .A(n3033), .B(n2532), .C(n3046), .D(n2531), .Y(n2041) );
  OAI22X1 U1686 ( .A(n3046), .B(n2532), .C(n3033), .D(n2533), .Y(n2042) );
  OAI22X1 U1687 ( .A(n3033), .B(n2534), .C(n3046), .D(n2533), .Y(n2043) );
  OAI22X1 U1688 ( .A(n3046), .B(n2534), .C(n3033), .D(n2535), .Y(n2044) );
  OAI22X1 U1689 ( .A(n3033), .B(n2536), .C(n3046), .D(n2535), .Y(n2045) );
  OAI22X1 U1690 ( .A(n3046), .B(n2536), .C(n3033), .D(n2537), .Y(n2046) );
  OAI22X1 U1691 ( .A(n3033), .B(n2538), .C(n3046), .D(n2537), .Y(n2047) );
  XNOR2X1 U1692 ( .A(n497), .B(n3137), .Y(n2507) );
  XNOR2X1 U1693 ( .A(n495), .B(n3138), .Y(n2508) );
  XNOR2X1 U1694 ( .A(n493), .B(n3138), .Y(n2509) );
  XNOR2X1 U1695 ( .A(n491), .B(n3138), .Y(n2510) );
  XNOR2X1 U1696 ( .A(n489), .B(n3138), .Y(n2511) );
  XNOR2X1 U1697 ( .A(n487), .B(n3138), .Y(n2512) );
  XNOR2X1 U1698 ( .A(n485), .B(n3138), .Y(n2513) );
  XNOR2X1 U1699 ( .A(n3028), .B(n3138), .Y(n2514) );
  XNOR2X1 U1700 ( .A(n3110), .B(n3138), .Y(n2515) );
  XNOR2X1 U1701 ( .A(n3108), .B(n3138), .Y(n2516) );
  XNOR2X1 U1702 ( .A(n3106), .B(n3138), .Y(n2517) );
  XNOR2X1 U1703 ( .A(n3104), .B(n3138), .Y(n2518) );
  XNOR2X1 U1704 ( .A(n3102), .B(n3138), .Y(n2519) );
  XNOR2X1 U1705 ( .A(n471), .B(n3138), .Y(n2520) );
  XNOR2X1 U1706 ( .A(n2964), .B(n3138), .Y(n2521) );
  XNOR2X1 U1707 ( .A(n467), .B(n3138), .Y(n2522) );
  XNOR2X1 U1708 ( .A(n3092), .B(n3138), .Y(n2523) );
  XNOR2X1 U1709 ( .A(n3089), .B(n3138), .Y(n2524) );
  XNOR2X1 U1710 ( .A(n3087), .B(n3138), .Y(n2525) );
  XNOR2X1 U1711 ( .A(n2968), .B(n3137), .Y(n2526) );
  XNOR2X1 U1712 ( .A(n2960), .B(n3138), .Y(n2527) );
  XNOR2X1 U1713 ( .A(n2967), .B(n3138), .Y(n2528) );
  XNOR2X1 U1714 ( .A(n2961), .B(n3137), .Y(n2529) );
  XNOR2X1 U1715 ( .A(n3076), .B(n3138), .Y(n2530) );
  XNOR2X1 U1716 ( .A(n2974), .B(n3137), .Y(n2531) );
  XNOR2X1 U1717 ( .A(n2975), .B(n3137), .Y(n2532) );
  XNOR2X1 U1718 ( .A(n3069), .B(n3137), .Y(n2533) );
  XNOR2X1 U1719 ( .A(n3067), .B(n3137), .Y(n2534) );
  XNOR2X1 U1720 ( .A(n2973), .B(n3137), .Y(n2535) );
  XNOR2X1 U1721 ( .A(n3062), .B(n3137), .Y(n2536) );
  XNOR2X1 U1722 ( .A(n437), .B(n3137), .Y(n2537) );
  XNOR2X1 U1723 ( .A(n3055), .B(n3137), .Y(n2538) );
  OAI22X1 U1724 ( .A(n3142), .B(n3034), .C(n3047), .D(n2572), .Y(n1765) );
  OAI22X1 U1725 ( .A(n3142), .B(n3047), .C(n3034), .D(n2540), .Y(n2050) );
  OAI22X1 U1726 ( .A(n3047), .B(n2540), .C(n3034), .D(n2541), .Y(n2051) );
  OAI22X1 U1727 ( .A(n3034), .B(n2542), .C(n3047), .D(n2541), .Y(n2052) );
  OAI22X1 U1728 ( .A(n3047), .B(n2542), .C(n3034), .D(n2543), .Y(n2053) );
  OAI22X1 U1729 ( .A(n3047), .B(n2543), .C(n3034), .D(n2544), .Y(n2054) );
  OAI22X1 U1730 ( .A(n3034), .B(n2545), .C(n3047), .D(n2544), .Y(n2055) );
  OAI22X1 U1731 ( .A(n3047), .B(n2545), .C(n3034), .D(n2546), .Y(n2056) );
  OAI22X1 U1732 ( .A(n3034), .B(n2547), .C(n3047), .D(n2546), .Y(n2057) );
  OAI22X1 U1733 ( .A(n3034), .B(n2548), .C(n3047), .D(n2547), .Y(n2058) );
  OAI22X1 U1734 ( .A(n3034), .B(n2549), .C(n3047), .D(n2548), .Y(n2059) );
  OAI22X1 U1735 ( .A(n3047), .B(n2549), .C(n3034), .D(n2550), .Y(n2060) );
  OAI22X1 U1736 ( .A(n3034), .B(n2551), .C(n3047), .D(n2550), .Y(n2061) );
  OAI22X1 U1737 ( .A(n3034), .B(n2552), .C(n3047), .D(n2551), .Y(n2062) );
  OAI22X1 U1738 ( .A(n3034), .B(n2553), .C(n3047), .D(n2552), .Y(n2063) );
  OAI22X1 U1739 ( .A(n3047), .B(n2553), .C(n3034), .D(n2554), .Y(n2064) );
  OAI22X1 U1740 ( .A(n3034), .B(n2555), .C(n3047), .D(n2554), .Y(n2065) );
  OAI22X1 U1741 ( .A(n3047), .B(n2555), .C(n3034), .D(n2556), .Y(n2066) );
  OAI22X1 U1742 ( .A(n3034), .B(n2557), .C(n3047), .D(n2556), .Y(n2067) );
  OAI22X1 U1743 ( .A(n3047), .B(n2557), .C(n3034), .D(n2558), .Y(n2068) );
  OAI22X1 U1744 ( .A(n3034), .B(n2559), .C(n3047), .D(n2558), .Y(n2069) );
  OAI22X1 U1745 ( .A(n3047), .B(n2559), .C(n3034), .D(n2560), .Y(n2070) );
  OAI22X1 U1746 ( .A(n3034), .B(n2561), .C(n3047), .D(n2560), .Y(n2071) );
  OAI22X1 U1747 ( .A(n3047), .B(n2561), .C(n3034), .D(n2562), .Y(n2072) );
  OAI22X1 U1748 ( .A(n3034), .B(n2563), .C(n3047), .D(n2562), .Y(n2073) );
  OAI22X1 U1749 ( .A(n3047), .B(n2563), .C(n3034), .D(n2564), .Y(n2074) );
  OAI22X1 U1750 ( .A(n3034), .B(n2565), .C(n3047), .D(n2564), .Y(n2075) );
  OAI22X1 U1751 ( .A(n3047), .B(n2565), .C(n3034), .D(n2566), .Y(n2076) );
  OAI22X1 U1752 ( .A(n3034), .B(n2567), .C(n3047), .D(n2566), .Y(n2077) );
  OAI22X1 U1753 ( .A(n3047), .B(n2567), .C(n3034), .D(n2568), .Y(n2078) );
  OAI22X1 U1754 ( .A(n3034), .B(n2569), .C(n3047), .D(n2568), .Y(n2079) );
  OAI22X1 U1755 ( .A(n3047), .B(n2569), .C(n3034), .D(n2570), .Y(n2080) );
  OAI22X1 U1756 ( .A(n3034), .B(n2571), .C(n3047), .D(n2570), .Y(n2081) );
  XNOR2X1 U1757 ( .A(n497), .B(n3141), .Y(n2540) );
  XNOR2X1 U1758 ( .A(n495), .B(n3140), .Y(n2541) );
  XNOR2X1 U1759 ( .A(n493), .B(n3140), .Y(n2542) );
  XNOR2X1 U1760 ( .A(n491), .B(n3140), .Y(n2543) );
  XNOR2X1 U1761 ( .A(n489), .B(n3140), .Y(n2544) );
  XNOR2X1 U1762 ( .A(n487), .B(n3140), .Y(n2545) );
  XNOR2X1 U1763 ( .A(n485), .B(n3140), .Y(n2546) );
  XNOR2X1 U1764 ( .A(n3029), .B(n3140), .Y(n2547) );
  XNOR2X1 U1765 ( .A(n3110), .B(n3140), .Y(n2548) );
  XNOR2X1 U1766 ( .A(n3108), .B(n3140), .Y(n2549) );
  XNOR2X1 U1767 ( .A(n3106), .B(n3140), .Y(n2550) );
  XNOR2X1 U1768 ( .A(n3104), .B(n3140), .Y(n2551) );
  XNOR2X1 U1769 ( .A(n3102), .B(n3140), .Y(n2552) );
  XNOR2X1 U1770 ( .A(n471), .B(n3140), .Y(n2553) );
  XNOR2X1 U1771 ( .A(n2976), .B(n3140), .Y(n2554) );
  XNOR2X1 U1772 ( .A(n467), .B(n3140), .Y(n2555) );
  XNOR2X1 U1773 ( .A(n3092), .B(n3140), .Y(n2556) );
  XNOR2X1 U1774 ( .A(n3089), .B(n3140), .Y(n2557) );
  XNOR2X1 U1775 ( .A(n3087), .B(n3140), .Y(n2558) );
  XNOR2X1 U1776 ( .A(n2968), .B(n3141), .Y(n2559) );
  XNOR2X1 U1777 ( .A(n2960), .B(n3140), .Y(n2560) );
  XNOR2X1 U1778 ( .A(n2967), .B(n3140), .Y(n2561) );
  XNOR2X1 U1779 ( .A(n2961), .B(n3141), .Y(n2562) );
  XNOR2X1 U1780 ( .A(n3076), .B(n3140), .Y(n2563) );
  XNOR2X1 U1781 ( .A(n2974), .B(n3141), .Y(n2564) );
  XNOR2X1 U1782 ( .A(n2975), .B(n3141), .Y(n2565) );
  XNOR2X1 U1783 ( .A(n3069), .B(n3141), .Y(n2566) );
  XNOR2X1 U1784 ( .A(n3067), .B(n3141), .Y(n2567) );
  XNOR2X1 U1785 ( .A(n2973), .B(n3141), .Y(n2568) );
  XNOR2X1 U1786 ( .A(n3062), .B(n3141), .Y(n2569) );
  XNOR2X1 U1787 ( .A(n437), .B(n3141), .Y(n2570) );
  XNOR2X1 U1788 ( .A(n3055), .B(n3141), .Y(n2571) );
  OAI22X1 U1789 ( .A(n3145), .B(n3035), .C(n3048), .D(n2605), .Y(n1766) );
  OAI22X1 U1790 ( .A(n3048), .B(n3145), .C(n3035), .D(n2573), .Y(n2084) );
  OAI22X1 U1791 ( .A(n3048), .B(n2573), .C(n3035), .D(n2574), .Y(n2085) );
  OAI22X1 U1792 ( .A(n3035), .B(n2575), .C(n3048), .D(n2574), .Y(n2086) );
  OAI22X1 U1793 ( .A(n3048), .B(n2575), .C(n3035), .D(n2576), .Y(n2087) );
  OAI22X1 U1794 ( .A(n3048), .B(n2576), .C(n3035), .D(n2577), .Y(n2088) );
  OAI22X1 U1795 ( .A(n3035), .B(n2578), .C(n3048), .D(n2577), .Y(n2089) );
  OAI22X1 U1796 ( .A(n3048), .B(n2578), .C(n3035), .D(n2579), .Y(n2090) );
  OAI22X1 U1797 ( .A(n3035), .B(n2580), .C(n3048), .D(n2579), .Y(n2091) );
  OAI22X1 U1798 ( .A(n3035), .B(n2581), .C(n3048), .D(n2580), .Y(n2092) );
  OAI22X1 U1799 ( .A(n3035), .B(n2582), .C(n3048), .D(n2581), .Y(n2093) );
  OAI22X1 U1800 ( .A(n3048), .B(n2582), .C(n3035), .D(n2583), .Y(n2094) );
  OAI22X1 U1801 ( .A(n3035), .B(n2584), .C(n3048), .D(n2583), .Y(n2095) );
  OAI22X1 U1802 ( .A(n3035), .B(n2585), .C(n3048), .D(n2584), .Y(n2096) );
  OAI22X1 U1803 ( .A(n3035), .B(n2586), .C(n3048), .D(n2585), .Y(n2097) );
  OAI22X1 U1804 ( .A(n3048), .B(n2586), .C(n3035), .D(n2587), .Y(n2098) );
  OAI22X1 U1805 ( .A(n3035), .B(n2588), .C(n3048), .D(n2587), .Y(n2099) );
  OAI22X1 U1806 ( .A(n3048), .B(n2588), .C(n3035), .D(n2589), .Y(n2100) );
  OAI22X1 U1807 ( .A(n3035), .B(n2590), .C(n3048), .D(n2589), .Y(n2101) );
  OAI22X1 U1808 ( .A(n3048), .B(n2590), .C(n3035), .D(n2591), .Y(n2102) );
  OAI22X1 U1809 ( .A(n3035), .B(n2592), .C(n3048), .D(n2591), .Y(n2103) );
  OAI22X1 U1810 ( .A(n3048), .B(n2592), .C(n3035), .D(n2593), .Y(n2104) );
  OAI22X1 U1811 ( .A(n3035), .B(n2594), .C(n3048), .D(n2593), .Y(n2105) );
  OAI22X1 U1812 ( .A(n3048), .B(n2594), .C(n3035), .D(n2595), .Y(n2106) );
  OAI22X1 U1813 ( .A(n3035), .B(n2596), .C(n3048), .D(n2595), .Y(n2107) );
  OAI22X1 U1814 ( .A(n3048), .B(n2596), .C(n3035), .D(n2597), .Y(n2108) );
  OAI22X1 U1815 ( .A(n3035), .B(n2598), .C(n3048), .D(n2597), .Y(n2109) );
  OAI22X1 U1816 ( .A(n3048), .B(n2598), .C(n3035), .D(n2599), .Y(n2110) );
  OAI22X1 U1817 ( .A(n3035), .B(n2600), .C(n3048), .D(n2599), .Y(n2111) );
  OAI22X1 U1818 ( .A(n3048), .B(n2600), .C(n3035), .D(n2601), .Y(n2112) );
  OAI22X1 U1819 ( .A(n3035), .B(n2602), .C(n3048), .D(n2601), .Y(n2113) );
  OAI22X1 U1820 ( .A(n3048), .B(n2602), .C(n3035), .D(n2603), .Y(n2114) );
  OAI22X1 U1821 ( .A(n3035), .B(n2604), .C(n3048), .D(n2603), .Y(n2115) );
  XNOR2X1 U1822 ( .A(n497), .B(n3144), .Y(n2573) );
  XNOR2X1 U1823 ( .A(n495), .B(n3143), .Y(n2574) );
  XNOR2X1 U1824 ( .A(n493), .B(n3143), .Y(n2575) );
  XNOR2X1 U1825 ( .A(n491), .B(n3143), .Y(n2576) );
  XNOR2X1 U1826 ( .A(n489), .B(n3143), .Y(n2577) );
  XNOR2X1 U1827 ( .A(n487), .B(n3143), .Y(n2578) );
  XNOR2X1 U1828 ( .A(n485), .B(n3143), .Y(n2579) );
  XNOR2X1 U1829 ( .A(n3028), .B(n3143), .Y(n2580) );
  XNOR2X1 U1830 ( .A(n3110), .B(n3143), .Y(n2581) );
  XNOR2X1 U1831 ( .A(n3108), .B(n3143), .Y(n2582) );
  XNOR2X1 U1832 ( .A(n3106), .B(n3143), .Y(n2583) );
  XNOR2X1 U1833 ( .A(n3104), .B(n3143), .Y(n2584) );
  XNOR2X1 U1834 ( .A(n3101), .B(n3143), .Y(n2585) );
  XNOR2X1 U1835 ( .A(n471), .B(n3143), .Y(n2586) );
  XNOR2X1 U1836 ( .A(n2964), .B(n3143), .Y(n2587) );
  XNOR2X1 U1837 ( .A(n467), .B(n3143), .Y(n2588) );
  XNOR2X1 U1838 ( .A(n3092), .B(n3143), .Y(n2589) );
  XNOR2X1 U1839 ( .A(n3089), .B(n3143), .Y(n2590) );
  XNOR2X1 U1840 ( .A(n3087), .B(n3143), .Y(n2591) );
  XNOR2X1 U1841 ( .A(n2968), .B(n3144), .Y(n2592) );
  XNOR2X1 U1842 ( .A(n2960), .B(n3143), .Y(n2593) );
  XNOR2X1 U1843 ( .A(n2967), .B(n3143), .Y(n2594) );
  XNOR2X1 U1844 ( .A(n2961), .B(n3144), .Y(n2595) );
  XNOR2X1 U1845 ( .A(n3076), .B(n3143), .Y(n2596) );
  XNOR2X1 U1846 ( .A(n2974), .B(n3144), .Y(n2597) );
  XNOR2X1 U1847 ( .A(n2975), .B(n3144), .Y(n2598) );
  XNOR2X1 U1848 ( .A(n2962), .B(n3144), .Y(n2599) );
  XNOR2X1 U1849 ( .A(n3067), .B(n3144), .Y(n2600) );
  XNOR2X1 U1850 ( .A(n2973), .B(n3144), .Y(n2601) );
  XNOR2X1 U1851 ( .A(n3062), .B(n3144), .Y(n2602) );
  XNOR2X1 U1852 ( .A(n437), .B(n3144), .Y(n2603) );
  XNOR2X1 U1853 ( .A(n3055), .B(n3144), .Y(n2604) );
  OAI22X1 U1854 ( .A(n3148), .B(n3036), .C(n3049), .D(n2638), .Y(n1767) );
  OAI22X1 U1855 ( .A(n3148), .B(n3049), .C(n3036), .D(n2606), .Y(n2118) );
  OAI22X1 U1856 ( .A(n3049), .B(n2606), .C(n3036), .D(n2607), .Y(n2119) );
  OAI22X1 U1857 ( .A(n3036), .B(n2608), .C(n3049), .D(n2607), .Y(n2120) );
  OAI22X1 U1858 ( .A(n3049), .B(n2608), .C(n3036), .D(n2609), .Y(n2121) );
  OAI22X1 U1859 ( .A(n3049), .B(n2609), .C(n3036), .D(n2610), .Y(n2122) );
  OAI22X1 U1860 ( .A(n3036), .B(n2611), .C(n3049), .D(n2610), .Y(n2123) );
  OAI22X1 U1861 ( .A(n3049), .B(n2611), .C(n3036), .D(n2612), .Y(n2124) );
  OAI22X1 U1862 ( .A(n3036), .B(n2613), .C(n3049), .D(n2612), .Y(n2125) );
  OAI22X1 U1863 ( .A(n3036), .B(n2614), .C(n3049), .D(n2613), .Y(n2126) );
  OAI22X1 U1864 ( .A(n3036), .B(n2615), .C(n3049), .D(n2614), .Y(n2127) );
  OAI22X1 U1865 ( .A(n3049), .B(n2615), .C(n3036), .D(n2616), .Y(n2128) );
  OAI22X1 U1866 ( .A(n3036), .B(n2617), .C(n3049), .D(n2616), .Y(n2129) );
  OAI22X1 U1867 ( .A(n3036), .B(n2618), .C(n3049), .D(n2617), .Y(n2130) );
  OAI22X1 U1868 ( .A(n3036), .B(n2619), .C(n3049), .D(n2618), .Y(n2131) );
  OAI22X1 U1869 ( .A(n3049), .B(n2619), .C(n3036), .D(n2620), .Y(n2132) );
  OAI22X1 U1870 ( .A(n3036), .B(n2621), .C(n3049), .D(n2620), .Y(n2133) );
  OAI22X1 U1871 ( .A(n3049), .B(n2621), .C(n3036), .D(n2622), .Y(n2134) );
  OAI22X1 U1872 ( .A(n3036), .B(n2623), .C(n3049), .D(n2622), .Y(n2135) );
  OAI22X1 U1873 ( .A(n3049), .B(n2623), .C(n3036), .D(n2624), .Y(n2136) );
  OAI22X1 U1874 ( .A(n3036), .B(n2625), .C(n3049), .D(n2624), .Y(n2137) );
  OAI22X1 U1875 ( .A(n3049), .B(n2625), .C(n3036), .D(n2626), .Y(n2138) );
  OAI22X1 U1876 ( .A(n3036), .B(n2627), .C(n3049), .D(n2626), .Y(n2139) );
  OAI22X1 U1877 ( .A(n3049), .B(n2627), .C(n3036), .D(n2628), .Y(n2140) );
  OAI22X1 U1878 ( .A(n3036), .B(n2629), .C(n3049), .D(n2628), .Y(n2141) );
  OAI22X1 U1879 ( .A(n3049), .B(n2629), .C(n3036), .D(n2630), .Y(n2142) );
  OAI22X1 U1880 ( .A(n3036), .B(n2631), .C(n3049), .D(n2630), .Y(n2143) );
  OAI22X1 U1881 ( .A(n3049), .B(n2631), .C(n3036), .D(n2632), .Y(n2144) );
  OAI22X1 U1882 ( .A(n3036), .B(n2633), .C(n3049), .D(n2632), .Y(n2145) );
  OAI22X1 U1883 ( .A(n3049), .B(n2633), .C(n3036), .D(n2634), .Y(n2146) );
  OAI22X1 U1884 ( .A(n3036), .B(n2635), .C(n3049), .D(n2634), .Y(n2147) );
  OAI22X1 U1885 ( .A(n3049), .B(n2635), .C(n3036), .D(n2636), .Y(n2148) );
  OAI22X1 U1886 ( .A(n3036), .B(n2637), .C(n3049), .D(n2636), .Y(n2149) );
  XNOR2X1 U1887 ( .A(n497), .B(n3147), .Y(n2606) );
  XNOR2X1 U1888 ( .A(n495), .B(n3146), .Y(n2607) );
  XNOR2X1 U1889 ( .A(n493), .B(n3146), .Y(n2608) );
  XNOR2X1 U1890 ( .A(n491), .B(n3146), .Y(n2609) );
  XNOR2X1 U1891 ( .A(n489), .B(n3146), .Y(n2610) );
  XNOR2X1 U1892 ( .A(n487), .B(n3146), .Y(n2611) );
  XNOR2X1 U1893 ( .A(n485), .B(n3146), .Y(n2612) );
  XNOR2X1 U1894 ( .A(n3029), .B(n3146), .Y(n2613) );
  XNOR2X1 U1895 ( .A(n481), .B(n3146), .Y(n2614) );
  XNOR2X1 U1896 ( .A(n3108), .B(n3146), .Y(n2615) );
  XNOR2X1 U1897 ( .A(n3106), .B(n3146), .Y(n2616) );
  XNOR2X1 U1898 ( .A(n3104), .B(n3146), .Y(n2617) );
  XNOR2X1 U1899 ( .A(n3102), .B(n3146), .Y(n2618) );
  XNOR2X1 U1900 ( .A(n471), .B(n3146), .Y(n2619) );
  XNOR2X1 U1901 ( .A(n3097), .B(n3146), .Y(n2620) );
  XNOR2X1 U1902 ( .A(n467), .B(n3146), .Y(n2621) );
  XNOR2X1 U1903 ( .A(n3091), .B(n3146), .Y(n2622) );
  XNOR2X1 U1904 ( .A(n3089), .B(n3146), .Y(n2623) );
  XNOR2X1 U1905 ( .A(n3086), .B(n3146), .Y(n2624) );
  XNOR2X1 U1906 ( .A(n3084), .B(n3147), .Y(n2625) );
  XNOR2X1 U1907 ( .A(n3082), .B(n3146), .Y(n2626) );
  XNOR2X1 U1908 ( .A(n3080), .B(n3146), .Y(n2627) );
  XNOR2X1 U1909 ( .A(n3078), .B(n3147), .Y(n2628) );
  XNOR2X1 U1910 ( .A(n3076), .B(n3146), .Y(n2629) );
  XNOR2X1 U1911 ( .A(n3074), .B(n3147), .Y(n2630) );
  XNOR2X1 U1912 ( .A(n3072), .B(n3147), .Y(n2631) );
  XNOR2X1 U1913 ( .A(n3069), .B(n3147), .Y(n2632) );
  XNOR2X1 U1914 ( .A(n3067), .B(n3147), .Y(n2633) );
  XNOR2X1 U1915 ( .A(n3064), .B(n3147), .Y(n2634) );
  XNOR2X1 U1916 ( .A(n3062), .B(n3147), .Y(n2635) );
  XNOR2X1 U1917 ( .A(n437), .B(n3147), .Y(n2636) );
  XNOR2X1 U1918 ( .A(n3055), .B(n3147), .Y(n2637) );
  OAI22X1 U1919 ( .A(n3151), .B(n3037), .C(n3050), .D(n2671), .Y(n1768) );
  OAI22X1 U1920 ( .A(n3151), .B(n3050), .C(n3037), .D(n2639), .Y(n2152) );
  OAI22X1 U1921 ( .A(n3050), .B(n2639), .C(n3037), .D(n2640), .Y(n2153) );
  OAI22X1 U1922 ( .A(n3037), .B(n2641), .C(n3050), .D(n2640), .Y(n2154) );
  OAI22X1 U1923 ( .A(n3050), .B(n2641), .C(n3037), .D(n2642), .Y(n2155) );
  OAI22X1 U1924 ( .A(n3050), .B(n2642), .C(n3037), .D(n2643), .Y(n2156) );
  OAI22X1 U1925 ( .A(n3037), .B(n2644), .C(n3050), .D(n2643), .Y(n2157) );
  OAI22X1 U1926 ( .A(n3050), .B(n2644), .C(n3037), .D(n2645), .Y(n2158) );
  OAI22X1 U1927 ( .A(n3037), .B(n2646), .C(n3050), .D(n2645), .Y(n2159) );
  OAI22X1 U1928 ( .A(n3037), .B(n2647), .C(n3050), .D(n2646), .Y(n2160) );
  OAI22X1 U1929 ( .A(n3037), .B(n2648), .C(n3050), .D(n2647), .Y(n2161) );
  OAI22X1 U1930 ( .A(n3050), .B(n2648), .C(n3037), .D(n2649), .Y(n2162) );
  OAI22X1 U1931 ( .A(n3037), .B(n2650), .C(n3050), .D(n2649), .Y(n2163) );
  OAI22X1 U1932 ( .A(n3037), .B(n2651), .C(n3050), .D(n2650), .Y(n2164) );
  OAI22X1 U1933 ( .A(n3037), .B(n2652), .C(n3050), .D(n2651), .Y(n2165) );
  OAI22X1 U1934 ( .A(n3050), .B(n2652), .C(n3037), .D(n2653), .Y(n2166) );
  OAI22X1 U1935 ( .A(n3037), .B(n2654), .C(n3050), .D(n2653), .Y(n2167) );
  OAI22X1 U1936 ( .A(n3050), .B(n2654), .C(n3037), .D(n2655), .Y(n2168) );
  OAI22X1 U1937 ( .A(n3037), .B(n2656), .C(n3050), .D(n2655), .Y(n2169) );
  OAI22X1 U1938 ( .A(n3050), .B(n2656), .C(n3037), .D(n2657), .Y(n2170) );
  OAI22X1 U1939 ( .A(n3037), .B(n2658), .C(n3050), .D(n2657), .Y(n2171) );
  OAI22X1 U1940 ( .A(n3050), .B(n2658), .C(n3037), .D(n2659), .Y(n2172) );
  OAI22X1 U1941 ( .A(n3037), .B(n2660), .C(n3050), .D(n2659), .Y(n2173) );
  OAI22X1 U1942 ( .A(n3050), .B(n2660), .C(n3037), .D(n2661), .Y(n2174) );
  OAI22X1 U1943 ( .A(n3037), .B(n2662), .C(n3050), .D(n2661), .Y(n2175) );
  OAI22X1 U1944 ( .A(n3050), .B(n2662), .C(n3037), .D(n2663), .Y(n2176) );
  OAI22X1 U1945 ( .A(n3037), .B(n2664), .C(n3050), .D(n2663), .Y(n2177) );
  OAI22X1 U1946 ( .A(n3050), .B(n2664), .C(n3037), .D(n2665), .Y(n2178) );
  OAI22X1 U1947 ( .A(n3037), .B(n2666), .C(n3050), .D(n2665), .Y(n2179) );
  OAI22X1 U1948 ( .A(n3050), .B(n2666), .C(n3037), .D(n2667), .Y(n2180) );
  OAI22X1 U1949 ( .A(n3037), .B(n2668), .C(n3050), .D(n2667), .Y(n2181) );
  OAI22X1 U1950 ( .A(n3050), .B(n2668), .C(n3037), .D(n2669), .Y(n2182) );
  OAI22X1 U1951 ( .A(n3037), .B(n2670), .C(n3050), .D(n2669), .Y(n2183) );
  XNOR2X1 U1952 ( .A(n497), .B(n3149), .Y(n2639) );
  XNOR2X1 U1953 ( .A(n495), .B(n3149), .Y(n2640) );
  XNOR2X1 U1954 ( .A(n493), .B(n3149), .Y(n2641) );
  XNOR2X1 U1955 ( .A(n491), .B(n3149), .Y(n2642) );
  XNOR2X1 U1956 ( .A(n489), .B(n3149), .Y(n2643) );
  XNOR2X1 U1957 ( .A(n487), .B(n3149), .Y(n2644) );
  XNOR2X1 U1958 ( .A(n485), .B(n3149), .Y(n2645) );
  XNOR2X1 U1959 ( .A(n3028), .B(n3149), .Y(n2646) );
  XNOR2X1 U1960 ( .A(n481), .B(n3149), .Y(n2647) );
  XNOR2X1 U1961 ( .A(n3108), .B(n3149), .Y(n2648) );
  XNOR2X1 U1962 ( .A(n3106), .B(n3149), .Y(n2649) );
  XNOR2X1 U1963 ( .A(n3104), .B(n3149), .Y(n2650) );
  XNOR2X1 U1964 ( .A(n3101), .B(n3150), .Y(n2651) );
  XNOR2X1 U1965 ( .A(n471), .B(n3150), .Y(n2652) );
  XNOR2X1 U1966 ( .A(n2965), .B(n3150), .Y(n2653) );
  XNOR2X1 U1967 ( .A(n467), .B(n3150), .Y(n2654) );
  XNOR2X1 U1968 ( .A(n3091), .B(n3150), .Y(n2655) );
  XNOR2X1 U1969 ( .A(n3089), .B(n3150), .Y(n2656) );
  XNOR2X1 U1970 ( .A(n3086), .B(n3150), .Y(n2657) );
  XNOR2X1 U1971 ( .A(n3084), .B(n3149), .Y(n2658) );
  XNOR2X1 U1972 ( .A(n3082), .B(n3150), .Y(n2659) );
  XNOR2X1 U1973 ( .A(n3080), .B(n3149), .Y(n2660) );
  XNOR2X1 U1974 ( .A(n3078), .B(n3149), .Y(n2661) );
  XNOR2X1 U1975 ( .A(n3076), .B(n3149), .Y(n2662) );
  XNOR2X1 U1976 ( .A(n3074), .B(n3149), .Y(n2663) );
  XNOR2X1 U1977 ( .A(n3072), .B(n3149), .Y(n2664) );
  XNOR2X1 U1978 ( .A(n3069), .B(n3149), .Y(n2665) );
  XNOR2X1 U1979 ( .A(n3067), .B(n3149), .Y(n2666) );
  XNOR2X1 U1980 ( .A(n3064), .B(n3149), .Y(n2667) );
  XNOR2X1 U1981 ( .A(n3062), .B(n3149), .Y(n2668) );
  XNOR2X1 U1982 ( .A(n437), .B(n3149), .Y(n2669) );
  XNOR2X1 U1983 ( .A(n3055), .B(n3149), .Y(n2670) );
  OAI22X1 U1984 ( .A(n3154), .B(n3038), .C(n3051), .D(n2704), .Y(n1769) );
  OAI22X1 U1985 ( .A(n3051), .B(n3154), .C(n3038), .D(n2672), .Y(n2186) );
  OAI22X1 U1986 ( .A(n3051), .B(n2672), .C(n3038), .D(n2673), .Y(n2187) );
  OAI22X1 U1987 ( .A(n3038), .B(n2674), .C(n3051), .D(n2673), .Y(n2188) );
  OAI22X1 U1988 ( .A(n3051), .B(n2674), .C(n3038), .D(n2675), .Y(n2189) );
  OAI22X1 U1989 ( .A(n3051), .B(n2675), .C(n3038), .D(n2676), .Y(n2190) );
  OAI22X1 U1990 ( .A(n3038), .B(n2677), .C(n3051), .D(n2676), .Y(n2191) );
  OAI22X1 U1991 ( .A(n3051), .B(n2677), .C(n3038), .D(n2678), .Y(n2192) );
  OAI22X1 U1992 ( .A(n3038), .B(n2679), .C(n3051), .D(n2678), .Y(n2193) );
  OAI22X1 U1993 ( .A(n3038), .B(n2680), .C(n3051), .D(n2679), .Y(n2194) );
  OAI22X1 U1994 ( .A(n3038), .B(n2681), .C(n3051), .D(n2680), .Y(n2195) );
  OAI22X1 U1995 ( .A(n3051), .B(n2681), .C(n3038), .D(n2682), .Y(n2196) );
  OAI22X1 U1996 ( .A(n3038), .B(n2683), .C(n3051), .D(n2682), .Y(n2197) );
  OAI22X1 U1997 ( .A(n3038), .B(n2684), .C(n3051), .D(n2683), .Y(n2198) );
  OAI22X1 U1998 ( .A(n3038), .B(n2685), .C(n3051), .D(n2684), .Y(n2199) );
  OAI22X1 U1999 ( .A(n3051), .B(n2685), .C(n3038), .D(n2686), .Y(n2200) );
  OAI22X1 U2000 ( .A(n3038), .B(n2687), .C(n3051), .D(n2686), .Y(n2201) );
  OAI22X1 U2001 ( .A(n3051), .B(n2687), .C(n3038), .D(n2688), .Y(n2202) );
  OAI22X1 U2002 ( .A(n3038), .B(n2689), .C(n3051), .D(n2688), .Y(n2203) );
  OAI22X1 U2003 ( .A(n3051), .B(n2689), .C(n3038), .D(n2690), .Y(n2204) );
  OAI22X1 U2004 ( .A(n3038), .B(n2691), .C(n3051), .D(n2690), .Y(n2205) );
  OAI22X1 U2005 ( .A(n3051), .B(n2691), .C(n3038), .D(n2692), .Y(n2206) );
  OAI22X1 U2006 ( .A(n3038), .B(n2693), .C(n3051), .D(n2692), .Y(n2207) );
  OAI22X1 U2007 ( .A(n3051), .B(n2693), .C(n3038), .D(n2694), .Y(n2208) );
  OAI22X1 U2008 ( .A(n3038), .B(n2695), .C(n3051), .D(n2694), .Y(n2209) );
  OAI22X1 U2009 ( .A(n3051), .B(n2695), .C(n3038), .D(n2696), .Y(n2210) );
  OAI22X1 U2010 ( .A(n3038), .B(n2697), .C(n3051), .D(n2696), .Y(n2211) );
  OAI22X1 U2011 ( .A(n3051), .B(n2697), .C(n3038), .D(n2698), .Y(n2212) );
  OAI22X1 U2012 ( .A(n3038), .B(n2699), .C(n3051), .D(n2698), .Y(n2213) );
  OAI22X1 U2013 ( .A(n3051), .B(n2699), .C(n3038), .D(n2700), .Y(n2214) );
  OAI22X1 U2014 ( .A(n3038), .B(n2701), .C(n3051), .D(n2700), .Y(n2215) );
  OAI22X1 U2015 ( .A(n3051), .B(n2701), .C(n3038), .D(n2702), .Y(n2216) );
  OAI22X1 U2016 ( .A(n3038), .B(n2703), .C(n3051), .D(n2702), .Y(n2217) );
  XNOR2X1 U2017 ( .A(n497), .B(n3153), .Y(n2672) );
  XNOR2X1 U2018 ( .A(n495), .B(n3152), .Y(n2673) );
  XNOR2X1 U2019 ( .A(n493), .B(n3152), .Y(n2674) );
  XNOR2X1 U2020 ( .A(n491), .B(n3152), .Y(n2675) );
  XNOR2X1 U2021 ( .A(n489), .B(n3152), .Y(n2676) );
  XNOR2X1 U2022 ( .A(n487), .B(n3152), .Y(n2677) );
  XNOR2X1 U2023 ( .A(n485), .B(n3152), .Y(n2678) );
  XNOR2X1 U2024 ( .A(n3029), .B(n3152), .Y(n2679) );
  XNOR2X1 U2025 ( .A(n481), .B(n3152), .Y(n2680) );
  XNOR2X1 U2026 ( .A(n3108), .B(n3152), .Y(n2681) );
  XNOR2X1 U2027 ( .A(n3106), .B(n3152), .Y(n2682) );
  XNOR2X1 U2028 ( .A(n3104), .B(n3152), .Y(n2683) );
  XNOR2X1 U2029 ( .A(n3102), .B(n3152), .Y(n2684) );
  XNOR2X1 U2030 ( .A(n471), .B(n3152), .Y(n2685) );
  XNOR2X1 U2031 ( .A(n3096), .B(n3152), .Y(n2686) );
  XNOR2X1 U2032 ( .A(n467), .B(n3152), .Y(n2687) );
  XNOR2X1 U2033 ( .A(n3091), .B(n3152), .Y(n2688) );
  XNOR2X1 U2034 ( .A(n3089), .B(n3152), .Y(n2689) );
  XNOR2X1 U2035 ( .A(n3086), .B(n3152), .Y(n2690) );
  XNOR2X1 U2036 ( .A(n3084), .B(n3153), .Y(n2691) );
  XNOR2X1 U2037 ( .A(n3082), .B(n3152), .Y(n2692) );
  XNOR2X1 U2038 ( .A(n3080), .B(n3152), .Y(n2693) );
  XNOR2X1 U2039 ( .A(n3078), .B(n3153), .Y(n2694) );
  XNOR2X1 U2040 ( .A(n3076), .B(n3152), .Y(n2695) );
  XNOR2X1 U2041 ( .A(n3074), .B(n3153), .Y(n2696) );
  XNOR2X1 U2042 ( .A(n3072), .B(n3153), .Y(n2697) );
  XNOR2X1 U2043 ( .A(n2963), .B(n3153), .Y(n2698) );
  XNOR2X1 U2044 ( .A(n3067), .B(n3153), .Y(n2699) );
  XNOR2X1 U2045 ( .A(n2973), .B(n3153), .Y(n2700) );
  XNOR2X1 U2046 ( .A(n3061), .B(n3153), .Y(n2701) );
  XNOR2X1 U2047 ( .A(n437), .B(n3153), .Y(n2702) );
  XNOR2X1 U2048 ( .A(n3055), .B(n3153), .Y(n2703) );
  OAI22X1 U2049 ( .A(n3157), .B(n3039), .C(n3158), .D(n2737), .Y(n1770) );
  OAI22X1 U2050 ( .A(n3158), .B(n3157), .C(n3039), .D(n2705), .Y(n2219) );
  OAI22X1 U2051 ( .A(n3158), .B(n2705), .C(n3039), .D(n2706), .Y(n2220) );
  OAI22X1 U2052 ( .A(n3039), .B(n2707), .C(n3158), .D(n2706), .Y(n2221) );
  OAI22X1 U2053 ( .A(n3158), .B(n2707), .C(n3039), .D(n2708), .Y(n2222) );
  OAI22X1 U2054 ( .A(n3158), .B(n2708), .C(n3039), .D(n2709), .Y(n2223) );
  OAI22X1 U2055 ( .A(n3039), .B(n2710), .C(n3158), .D(n2709), .Y(n2224) );
  OAI22X1 U2056 ( .A(n3158), .B(n2710), .C(n3039), .D(n2711), .Y(n2225) );
  OAI22X1 U2057 ( .A(n3039), .B(n2712), .C(n3158), .D(n2711), .Y(n2226) );
  OAI22X1 U2058 ( .A(n3039), .B(n2713), .C(n3158), .D(n2712), .Y(n2227) );
  OAI22X1 U2059 ( .A(n3039), .B(n2714), .C(n3158), .D(n2713), .Y(n2228) );
  OAI22X1 U2060 ( .A(n3158), .B(n2714), .C(n3039), .D(n2715), .Y(n2229) );
  OAI22X1 U2061 ( .A(n3039), .B(n2716), .C(n3158), .D(n2715), .Y(n2230) );
  OAI22X1 U2062 ( .A(n3039), .B(n2717), .C(n3158), .D(n2716), .Y(n2231) );
  OAI22X1 U2063 ( .A(n3039), .B(n2718), .C(n3158), .D(n2717), .Y(n2232) );
  OAI22X1 U2064 ( .A(n3158), .B(n2718), .C(n3039), .D(n2719), .Y(n2233) );
  OAI22X1 U2065 ( .A(n3039), .B(n2720), .C(n3158), .D(n2719), .Y(n2234) );
  OAI22X1 U2066 ( .A(n3158), .B(n2720), .C(n3039), .D(n2721), .Y(n2235) );
  OAI22X1 U2067 ( .A(n3039), .B(n2722), .C(n3158), .D(n2721), .Y(n2236) );
  OAI22X1 U2068 ( .A(n3158), .B(n2722), .C(n3039), .D(n2723), .Y(n2237) );
  OAI22X1 U2069 ( .A(n3039), .B(n2724), .C(n3158), .D(n2723), .Y(n2238) );
  OAI22X1 U2070 ( .A(n3158), .B(n2724), .C(n3039), .D(n2725), .Y(n2239) );
  OAI22X1 U2071 ( .A(n3039), .B(n2726), .C(n3158), .D(n2725), .Y(n2240) );
  OAI22X1 U2072 ( .A(n3158), .B(n2726), .C(n3039), .D(n2727), .Y(n2241) );
  OAI22X1 U2073 ( .A(n3039), .B(n2728), .C(n3158), .D(n2727), .Y(n2242) );
  OAI22X1 U2074 ( .A(n3158), .B(n2728), .C(n3039), .D(n2729), .Y(n2243) );
  OAI22X1 U2075 ( .A(n3039), .B(n2730), .C(n3158), .D(n2729), .Y(n2244) );
  OAI22X1 U2076 ( .A(n3158), .B(n2730), .C(n3039), .D(n2731), .Y(n2245) );
  OAI22X1 U2077 ( .A(n3039), .B(n2732), .C(n3158), .D(n2731), .Y(n2246) );
  OAI22X1 U2078 ( .A(n3158), .B(n2732), .C(n3039), .D(n2733), .Y(n2247) );
  OAI22X1 U2079 ( .A(n3039), .B(n2734), .C(n3158), .D(n2733), .Y(n2248) );
  OAI22X1 U2080 ( .A(n3158), .B(n2734), .C(n3039), .D(n2735), .Y(n2249) );
  OAI22X1 U2081 ( .A(n3039), .B(n2736), .C(n3158), .D(n2735), .Y(n2250) );
  XNOR2X1 U2082 ( .A(n497), .B(n3155), .Y(n2705) );
  XNOR2X1 U2083 ( .A(n495), .B(n3156), .Y(n2706) );
  XNOR2X1 U2084 ( .A(n493), .B(n3156), .Y(n2707) );
  XNOR2X1 U2085 ( .A(n491), .B(n3156), .Y(n2708) );
  XNOR2X1 U2086 ( .A(n489), .B(n3156), .Y(n2709) );
  XNOR2X1 U2087 ( .A(n487), .B(n3156), .Y(n2710) );
  XNOR2X1 U2088 ( .A(n485), .B(n3156), .Y(n2711) );
  XNOR2X1 U2089 ( .A(n3028), .B(n3156), .Y(n2712) );
  XNOR2X1 U2090 ( .A(n481), .B(n3156), .Y(n2713) );
  XNOR2X1 U2091 ( .A(n3108), .B(n3156), .Y(n2714) );
  XNOR2X1 U2092 ( .A(n3106), .B(n3156), .Y(n2715) );
  XNOR2X1 U2093 ( .A(n3104), .B(n3156), .Y(n2716) );
  XNOR2X1 U2094 ( .A(n3101), .B(n3156), .Y(n2717) );
  XNOR2X1 U2095 ( .A(n471), .B(n3156), .Y(n2718) );
  XNOR2X1 U2096 ( .A(n3096), .B(n3156), .Y(n2719) );
  XNOR2X1 U2097 ( .A(n467), .B(n3156), .Y(n2720) );
  XNOR2X1 U2098 ( .A(n3091), .B(n3156), .Y(n2721) );
  XNOR2X1 U2099 ( .A(n3089), .B(n3156), .Y(n2722) );
  XNOR2X1 U2100 ( .A(n3086), .B(n3156), .Y(n2723) );
  XNOR2X1 U2101 ( .A(n3084), .B(n3155), .Y(n2724) );
  XNOR2X1 U2102 ( .A(n3082), .B(n3156), .Y(n2725) );
  XNOR2X1 U2103 ( .A(n3080), .B(n3156), .Y(n2726) );
  XNOR2X1 U2104 ( .A(n3078), .B(n3155), .Y(n2727) );
  XNOR2X1 U2105 ( .A(n3076), .B(n3156), .Y(n2728) );
  XNOR2X1 U2106 ( .A(n3074), .B(n3155), .Y(n2729) );
  XNOR2X1 U2107 ( .A(n3072), .B(n3155), .Y(n2730) );
  XNOR2X1 U2108 ( .A(n3069), .B(n3155), .Y(n2731) );
  XNOR2X1 U2109 ( .A(n3066), .B(n3155), .Y(n2732) );
  XNOR2X1 U2110 ( .A(n2973), .B(n3155), .Y(n2733) );
  XNOR2X1 U2111 ( .A(n3061), .B(n3155), .Y(n2734) );
  XNOR2X1 U2112 ( .A(n437), .B(n3155), .Y(n2735) );
  XNOR2X1 U2113 ( .A(n3055), .B(n3155), .Y(n2736) );
  XOR2X1 U2148 ( .A(b[30]), .B(n3053), .Y(n2764) );
  XOR2X1 U2151 ( .A(b[28]), .B(n3113), .Y(n2765) );
  XOR2X1 U2154 ( .A(b[26]), .B(n3116), .Y(n2766) );
  XOR2X1 U2160 ( .A(n3123), .B(b[22]), .Y(n2768) );
  XOR2X1 U2163 ( .A(n3126), .B(b[20]), .Y(n2769) );
  XOR2X1 U2166 ( .A(n3129), .B(b[18]), .Y(n2770) );
  XOR2X1 U2169 ( .A(n3131), .B(b[16]), .Y(n2771) );
  XOR2X1 U2172 ( .A(n3135), .B(b[14]), .Y(n2772) );
  XOR2X1 U2175 ( .A(n3138), .B(b[12]), .Y(n2773) );
  XOR2X1 U2178 ( .A(b[10]), .B(n3140), .Y(n2774) );
  XOR2X1 U2181 ( .A(n3143), .B(b[8]), .Y(n2775) );
  XOR2X1 U2184 ( .A(n3146), .B(b[6]), .Y(n2776) );
  XOR2X1 U2187 ( .A(n3150), .B(b[4]), .Y(n2777) );
  XOR2X1 U2190 ( .A(n3152), .B(b[2]), .Y(n2778) );
  XOR2X1 U2193 ( .A(n3156), .B(b[0]), .Y(n2779) );
  INVX4 U2197 ( .A(n735), .Y(n734) );
  INVX8 U2198 ( .A(n3083), .Y(n3082) );
  INVX8 U2199 ( .A(n3085), .Y(n3084) );
  INVX8 U2200 ( .A(n3079), .Y(n3078) );
  INVX8 U2201 ( .A(n3075), .Y(n3074) );
  INVX8 U2202 ( .A(n3107), .Y(n3106) );
  INVX8 U2203 ( .A(n3073), .Y(n3072) );
  INVX8 U2204 ( .A(n3081), .Y(n3080) );
  INVX4 U2205 ( .A(n455), .Y(n3081) );
  INVX8 U2206 ( .A(n3109), .Y(n3108) );
  INVX4 U2207 ( .A(n479), .Y(n3109) );
  INVX8 U2208 ( .A(n3105), .Y(n3104) );
  INVX4 U2209 ( .A(n475), .Y(n3105) );
  BUFX4 U2210 ( .A(n3178), .Y(product[28]) );
  INVX4 U2211 ( .A(n3027), .Y(n3028) );
  INVX4 U2212 ( .A(n483), .Y(n3027) );
  INVX4 U2213 ( .A(n3063), .Y(n3062) );
  INVX4 U2214 ( .A(n439), .Y(n3063) );
  INVX8 U2215 ( .A(n3088), .Y(n3086) );
  INVX4 U2216 ( .A(n461), .Y(n3088) );
  INVX2 U2217 ( .A(n451), .Y(n3077) );
  INVX2 U2218 ( .A(n445), .Y(n3071) );
  INVX4 U2219 ( .A(n3071), .Y(n3069) );
  INVX2 U2220 ( .A(n3093), .Y(n3092) );
  INVX4 U2221 ( .A(n3065), .Y(n3064) );
  INVX2 U2222 ( .A(n473), .Y(n3103) );
  INVX2 U2223 ( .A(n465), .Y(n3093) );
  INVX4 U2224 ( .A(n3103), .Y(n3101) );
  INVX4 U2225 ( .A(n3063), .Y(n3061) );
  INVX2 U2226 ( .A(n477), .Y(n3107) );
  INVX2 U2227 ( .A(n3111), .Y(n3110) );
  INVX1 U2228 ( .A(n698), .Y(n697) );
  BUFX4 U2229 ( .A(n3179), .Y(product[22]) );
  NAND2X1 U2230 ( .A(n2769), .B(n3042), .Y(n2923) );
  NAND2X1 U2231 ( .A(n2768), .B(n3041), .Y(n2924) );
  XNOR2X1 U2232 ( .A(b[26]), .B(n3119), .Y(n2925) );
  XNOR2X1 U2233 ( .A(n3116), .B(b[28]), .Y(n2926) );
  XNOR2X1 U2234 ( .A(n3113), .B(b[30]), .Y(n2927) );
  INVX2 U2235 ( .A(b[0]), .Y(n3158) );
  NAND2X1 U2236 ( .A(n2925), .B(n2766), .Y(n2928) );
  OR2X2 U2237 ( .A(n3016), .B(n3015), .Y(n2929) );
  NAND2X1 U2238 ( .A(n2765), .B(n2926), .Y(n2930) );
  NAND2X1 U2239 ( .A(n2764), .B(n2927), .Y(n2931) );
  INVX1 U2240 ( .A(n437), .Y(n3060) );
  INVX2 U2241 ( .A(n471), .Y(n3100) );
  INVX2 U2242 ( .A(n467), .Y(n3095) );
  INVX2 U2243 ( .A(n443), .Y(n3068) );
  INVX2 U2244 ( .A(n463), .Y(n3090) );
  INVX2 U2245 ( .A(n764), .Y(n2942) );
  INVX2 U2246 ( .A(n784), .Y(n783) );
  OR2X2 U2247 ( .A(n932), .B(n913), .Y(n2932) );
  AND2X2 U2248 ( .A(n691), .B(n874), .Y(n2933) );
  XOR2X1 U2249 ( .A(n1620), .B(n1618), .Y(n2934) );
  XOR2X1 U2250 ( .A(n2934), .B(n1631), .Y(n1614) );
  XOR2X1 U2251 ( .A(n1616), .B(n1629), .Y(n2935) );
  XOR2X1 U2252 ( .A(n2935), .B(n1614), .Y(n1612) );
  NAND2X1 U2253 ( .A(n1620), .B(n1618), .Y(n2936) );
  NAND2X1 U2254 ( .A(n1620), .B(n1631), .Y(n2937) );
  NAND2X1 U2255 ( .A(n1618), .B(n1631), .Y(n2938) );
  NAND3X1 U2256 ( .A(n2936), .B(n2937), .C(n2938), .Y(n1613) );
  NAND2X1 U2257 ( .A(n1616), .B(n1629), .Y(n2939) );
  NAND2X1 U2258 ( .A(n1616), .B(n1614), .Y(n2940) );
  NAND2X1 U2259 ( .A(n1629), .B(n1614), .Y(n2941) );
  NAND3X1 U2260 ( .A(n2939), .B(n2940), .C(n2941), .Y(n1611) );
  BUFX2 U2261 ( .A(n1214), .Y(n2943) );
  XOR2X1 U2262 ( .A(n1964), .B(n1780), .Y(n2944) );
  XOR2X1 U2263 ( .A(n2219), .B(n2944), .Y(n1304) );
  NAND2X1 U2264 ( .A(n2219), .B(n1964), .Y(n2945) );
  NAND2X1 U2265 ( .A(n2219), .B(n1780), .Y(n2946) );
  NAND2X1 U2266 ( .A(n1964), .B(n1780), .Y(n2947) );
  NAND3X1 U2267 ( .A(n2945), .B(n2946), .C(n2947), .Y(n1303) );
  XOR2X1 U2268 ( .A(n1541), .B(n1520), .Y(n2948) );
  XOR2X1 U2269 ( .A(n2948), .B(n1539), .Y(n1516) );
  XOR2X1 U2270 ( .A(n1518), .B(n1537), .Y(n2949) );
  XOR2X1 U2271 ( .A(n2949), .B(n1516), .Y(n1514) );
  NAND2X1 U2272 ( .A(n1541), .B(n1520), .Y(n2950) );
  NAND2X1 U2273 ( .A(n1541), .B(n1539), .Y(n2951) );
  NAND2X1 U2274 ( .A(n1520), .B(n1539), .Y(n2952) );
  NAND3X1 U2275 ( .A(n2950), .B(n2951), .C(n2952), .Y(n1515) );
  NAND2X1 U2276 ( .A(n1518), .B(n1537), .Y(n2953) );
  NAND2X1 U2277 ( .A(n1518), .B(n1516), .Y(n2954) );
  NAND2X1 U2278 ( .A(n1537), .B(n1516), .Y(n2955) );
  NAND3X1 U2279 ( .A(n2953), .B(n2954), .C(n2955), .Y(n1513) );
  INVX1 U2280 ( .A(n797), .Y(n796) );
  INVX8 U2281 ( .A(n3068), .Y(n3067) );
  XNOR2X1 U2282 ( .A(n2956), .B(n1185), .Y(n1183) );
  XNOR2X1 U2283 ( .A(n1214), .B(n1187), .Y(n2956) );
  NAND2X1 U2284 ( .A(n1185), .B(n2943), .Y(n2957) );
  NAND2X1 U2285 ( .A(n1185), .B(n1187), .Y(n2958) );
  NAND2X1 U2286 ( .A(n2943), .B(n1187), .Y(n2959) );
  NAND3X1 U2287 ( .A(n2957), .B(n2958), .C(n2959), .Y(n1182) );
  BUFX4 U2288 ( .A(n441), .Y(n2973) );
  INVX1 U2289 ( .A(n685), .Y(n687) );
  INVX1 U2290 ( .A(n690), .Y(n874) );
  XNOR2X1 U2291 ( .A(n692), .B(n2933), .Y(product[29]) );
  BUFX4 U2292 ( .A(n499), .Y(n3020) );
  INVX2 U2293 ( .A(n638), .Y(n640) );
  INVX2 U2294 ( .A(n698), .Y(n3022) );
  INVX4 U2295 ( .A(n3027), .Y(n3029) );
  BUFX2 U2296 ( .A(n457), .Y(n2960) );
  BUFX2 U2297 ( .A(n453), .Y(n2961) );
  INVX1 U2298 ( .A(n3071), .Y(n2962) );
  INVX1 U2299 ( .A(n3071), .Y(n2963) );
  INVX2 U2300 ( .A(n3098), .Y(n2964) );
  INVX2 U2301 ( .A(n3098), .Y(n2965) );
  BUFX4 U2302 ( .A(n3177), .Y(product[44]) );
  BUFX2 U2303 ( .A(n455), .Y(n2967) );
  BUFX2 U2304 ( .A(n459), .Y(n2968) );
  INVX8 U2305 ( .A(n3093), .Y(n3091) );
  INVX8 U2306 ( .A(n3090), .Y(n3089) );
  INVX1 U2307 ( .A(n3071), .Y(n3070) );
  INVX2 U2308 ( .A(n3088), .Y(n3087) );
  BUFX4 U2309 ( .A(n449), .Y(n2974) );
  BUFX4 U2310 ( .A(n447), .Y(n2975) );
  INVX1 U2311 ( .A(n3068), .Y(n3066) );
  INVX2 U2312 ( .A(n441), .Y(n3065) );
  NAND2X1 U2313 ( .A(n727), .B(n522), .Y(n2971) );
  NAND2X1 U2314 ( .A(n2969), .B(n2970), .Y(n2972) );
  NAND2X1 U2315 ( .A(n2971), .B(n2972), .Y(product[25]) );
  INVX1 U2316 ( .A(n727), .Y(n2969) );
  INVX1 U2317 ( .A(n522), .Y(n2970) );
  INVX8 U2318 ( .A(n3077), .Y(n3076) );
  INVX4 U2319 ( .A(n469), .Y(n3098) );
  INVX2 U2320 ( .A(n3098), .Y(n3096) );
  INVX1 U2321 ( .A(n3098), .Y(n2976) );
  INVX2 U2322 ( .A(n481), .Y(n3111) );
  XOR2X1 U2323 ( .A(n791), .B(n2978), .Y(product[16]) );
  NAND2X1 U2324 ( .A(n790), .B(n2986), .Y(n2978) );
  AND2X2 U2325 ( .A(n856), .B(n2993), .Y(product[1]) );
  OR2X1 U2326 ( .A(n2250), .B(n1770), .Y(n2993) );
  INVX2 U2327 ( .A(n3057), .Y(n3056) );
  INVX4 U2328 ( .A(n3103), .Y(n3102) );
  INVX2 U2329 ( .A(n3098), .Y(n3097) );
  INVX1 U2330 ( .A(n3095), .Y(n3094) );
  INVX1 U2331 ( .A(n3100), .Y(n3099) );
  INVX4 U2332 ( .A(n453), .Y(n3079) );
  INVX4 U2333 ( .A(n459), .Y(n3085) );
  INVX4 U2334 ( .A(n449), .Y(n3075) );
  INVX4 U2335 ( .A(n447), .Y(n3073) );
  INVX4 U2336 ( .A(n457), .Y(n3083) );
  OR2X2 U2337 ( .A(n996), .B(n975), .Y(n2979) );
  OR2X2 U2338 ( .A(n1467), .B(n1444), .Y(n2980) );
  OR2X2 U2339 ( .A(n1443), .B(n1418), .Y(n2981) );
  OR2X2 U2340 ( .A(n1491), .B(n1468), .Y(n2982) );
  OR2X2 U2341 ( .A(n974), .B(n953), .Y(n2983) );
  XNOR2X1 U2342 ( .A(n547), .B(n2984), .Y(product[47]) );
  XNOR2X1 U2343 ( .A(n903), .B(n912), .Y(n2984) );
  OR2X2 U2344 ( .A(n1627), .B(n1612), .Y(n2985) );
  OR2X2 U2345 ( .A(n1657), .B(n1644), .Y(n2986) );
  OR2X2 U2346 ( .A(n1671), .B(n1658), .Y(n2987) );
  OR2X2 U2347 ( .A(n1705), .B(n1696), .Y(n2988) );
  OR2X2 U2348 ( .A(n1715), .B(n1706), .Y(n2989) );
  OR2X2 U2349 ( .A(n1751), .B(n1748), .Y(n2990) );
  OR2X2 U2350 ( .A(n1743), .B(n1738), .Y(n2991) );
  INVX2 U2351 ( .A(n3054), .Y(n3052) );
  INVX2 U2352 ( .A(n3054), .Y(n3053) );
  XOR2X1 U2353 ( .A(n3109), .B(n3118), .Y(n2330) );
  INVX2 U2354 ( .A(n3151), .Y(n3150) );
  INVX1 U2355 ( .A(n333), .Y(n3054) );
  INVX2 U2356 ( .A(n2996), .Y(n3050) );
  INVX2 U2357 ( .A(n3000), .Y(n3039) );
  INVX2 U2358 ( .A(n3001), .Y(n3038) );
  INVX2 U2359 ( .A(n2994), .Y(n3035) );
  INVX2 U2360 ( .A(n2995), .Y(n3037) );
  INVX2 U2361 ( .A(n2998), .Y(n3051) );
  INVX2 U2362 ( .A(n3002), .Y(n3032) );
  INVX2 U2363 ( .A(n2997), .Y(n3048) );
  INVX2 U2364 ( .A(n2999), .Y(n3045) );
  INVX2 U2365 ( .A(n3133), .Y(n3132) );
  INVX2 U2366 ( .A(n3130), .Y(n3129) );
  INVX2 U2367 ( .A(n3005), .Y(n3030) );
  INVX2 U2368 ( .A(n3133), .Y(n3131) );
  INVX2 U2369 ( .A(n3130), .Y(n3128) );
  AND2X1 U2370 ( .A(n3048), .B(n2775), .Y(n2994) );
  AND2X1 U2371 ( .A(n3050), .B(n2777), .Y(n2995) );
  INVX2 U2372 ( .A(n3145), .Y(n3143) );
  INVX2 U2373 ( .A(n3139), .Y(n3138) );
  INVX2 U2374 ( .A(n3136), .Y(n3135) );
  INVX2 U2375 ( .A(n3127), .Y(n3125) );
  INVX2 U2376 ( .A(n3117), .Y(n3116) );
  INVX2 U2377 ( .A(n3124), .Y(n3122) );
  INVX2 U2378 ( .A(n3124), .Y(n3121) );
  INVX2 U2379 ( .A(n3114), .Y(n3112) );
  INVX2 U2380 ( .A(n3120), .Y(n3118) );
  INVX2 U2381 ( .A(n3120), .Y(n3119) );
  INVX2 U2382 ( .A(n3117), .Y(n3115) );
  INVX2 U2383 ( .A(n3151), .Y(n3149) );
  INVX2 U2384 ( .A(n3114), .Y(n3113) );
  XOR2X1 U2385 ( .A(b[4]), .B(n3153), .Y(n2996) );
  XOR2X1 U2386 ( .A(b[8]), .B(n3147), .Y(n2997) );
  XOR2X1 U2387 ( .A(b[2]), .B(n3155), .Y(n2998) );
  XOR2X1 U2388 ( .A(b[14]), .B(n3137), .Y(n2999) );
  AND2X1 U2389 ( .A(n3158), .B(n2779), .Y(n3000) );
  AND2X1 U2390 ( .A(n3051), .B(n2778), .Y(n3001) );
  AND2X1 U2391 ( .A(n3045), .B(n2772), .Y(n3002) );
  INVX2 U2392 ( .A(n3012), .Y(n3046) );
  INVX2 U2393 ( .A(n3011), .Y(n3047) );
  INVX2 U2394 ( .A(n3010), .Y(n3049) );
  INVX2 U2395 ( .A(n3009), .Y(n3033) );
  INVX2 U2396 ( .A(n3008), .Y(n3036) );
  INVX2 U2397 ( .A(n3006), .Y(n3031) );
  INVX1 U2398 ( .A(n295), .Y(n3151) );
  INVX2 U2399 ( .A(n3013), .Y(n3041) );
  INVX2 U2400 ( .A(n3007), .Y(n3034) );
  INVX2 U2401 ( .A(n3015), .Y(n3040) );
  INVX2 U2402 ( .A(n3003), .Y(n3042) );
  INVX2 U2403 ( .A(n3004), .Y(n3043) );
  INVX2 U2404 ( .A(n3127), .Y(n3126) );
  INVX2 U2405 ( .A(n3014), .Y(n3044) );
  INVX2 U2406 ( .A(n3124), .Y(n3123) );
  INVX2 U2407 ( .A(n3154), .Y(n3152) );
  XOR2X1 U2408 ( .A(n3129), .B(b[20]), .Y(n3003) );
  XOR2X1 U2409 ( .A(b[18]), .B(n3132), .Y(n3004) );
  AND2X1 U2410 ( .A(n2770), .B(n3043), .Y(n3005) );
  AND2X1 U2411 ( .A(n3044), .B(n2771), .Y(n3006) );
  AND2X1 U2412 ( .A(n2774), .B(n3047), .Y(n3007) );
  AND2X1 U2413 ( .A(n2776), .B(n3049), .Y(n3008) );
  AND2X1 U2414 ( .A(n2773), .B(n3046), .Y(n3009) );
  INVX2 U2415 ( .A(n3136), .Y(n3134) );
  INVX2 U2416 ( .A(n3142), .Y(n3141) );
  INVX2 U2417 ( .A(n3139), .Y(n3137) );
  INVX2 U2418 ( .A(n3142), .Y(n3140) );
  INVX2 U2419 ( .A(n3145), .Y(n3144) );
  INVX2 U2420 ( .A(n3148), .Y(n3146) );
  INVX2 U2421 ( .A(n3148), .Y(n3147) );
  INVX2 U2422 ( .A(n3157), .Y(n3155) );
  INVX2 U2423 ( .A(n3154), .Y(n3153) );
  INVX1 U2424 ( .A(n292), .Y(n3154) );
  INVX2 U2425 ( .A(n3157), .Y(n3156) );
  XOR2X1 U2426 ( .A(n3150), .B(b[6]), .Y(n3010) );
  XOR2X1 U2427 ( .A(b[10]), .B(n3144), .Y(n3011) );
  XOR2X1 U2428 ( .A(b[12]), .B(n3141), .Y(n3012) );
  XOR2X1 U2429 ( .A(n3126), .B(b[22]), .Y(n3013) );
  XOR2X1 U2430 ( .A(n3135), .B(b[16]), .Y(n3014) );
  XOR2X1 U2431 ( .A(n3123), .B(b[24]), .Y(n3015) );
  INVX1 U2432 ( .A(n319), .Y(n3127) );
  INVX1 U2433 ( .A(n322), .Y(n3124) );
  INVX1 U2434 ( .A(n325), .Y(n3120) );
  INVX1 U2435 ( .A(n330), .Y(n3114) );
  XNOR2X1 U2436 ( .A(n3118), .B(b[24]), .Y(n3016) );
  INVX1 U2437 ( .A(n328), .Y(n3117) );
  INVX1 U2438 ( .A(n289), .Y(n3157) );
  INVX1 U2439 ( .A(n313), .Y(n3133) );
  INVX1 U2440 ( .A(n745), .Y(n881) );
  INVX1 U2441 ( .A(n298), .Y(n3148) );
  INVX1 U2442 ( .A(n304), .Y(n3142) );
  INVX1 U2443 ( .A(n307), .Y(n3139) );
  INVX2 U2444 ( .A(n433), .Y(n3059) );
  INVX2 U2445 ( .A(n433), .Y(n3058) );
  INVX1 U2446 ( .A(n301), .Y(n3145) );
  INVX1 U2447 ( .A(n310), .Y(n3136) );
  INVX1 U2448 ( .A(n316), .Y(n3130) );
  BUFX4 U2449 ( .A(n668), .Y(n3017) );
  BUFX2 U2450 ( .A(n668), .Y(n3018) );
  INVX2 U2451 ( .A(n669), .Y(n668) );
  BUFX2 U2452 ( .A(n499), .Y(n3019) );
  INVX1 U2453 ( .A(n751), .Y(n753) );
  OR2X2 U2454 ( .A(n1769), .B(n1754), .Y(n3021) );
  XOR2X1 U2455 ( .A(n1448), .B(n1469), .Y(n3023) );
  XOR2X1 U2456 ( .A(n1446), .B(n3023), .Y(n1444) );
  NAND2X1 U2457 ( .A(n1446), .B(n1448), .Y(n3024) );
  NAND2X1 U2458 ( .A(n1446), .B(n1469), .Y(n3025) );
  NAND2X1 U2459 ( .A(n1448), .B(n1469), .Y(n3026) );
  NAND3X1 U2460 ( .A(n3024), .B(n3025), .C(n3026), .Y(n1443) );
  INVX1 U2461 ( .A(n740), .Y(n880) );
  INVX1 U2462 ( .A(n819), .Y(n818) );
  INVX1 U2463 ( .A(n828), .Y(n827) );
  INVX1 U2464 ( .A(n806), .Y(n805) );
  INVX1 U2465 ( .A(n627), .Y(n866) );
  INVX1 U2466 ( .A(n663), .Y(n870) );
  INVX1 U2467 ( .A(n658), .Y(n656) );
  INVX8 U2468 ( .A(n3057), .Y(n3055) );
  INVX8 U2469 ( .A(n433), .Y(n3057) );
  NOR2X1 U2470 ( .A(n3158), .B(n3058), .Y(product[0]) );
  INVX2 U2471 ( .A(n972), .Y(n973) );
  INVX2 U2472 ( .A(n930), .Y(n931) );
  XOR2X1 U2473 ( .A(n3159), .B(n914), .Y(n903) );
  XOR2X1 U2474 ( .A(n3160), .B(n3161), .Y(n3159) );
  XOR2X1 U2475 ( .A(n3162), .B(n916), .Y(n3161) );
  XOR2X1 U2476 ( .A(n3163), .B(n3164), .Y(n3162) );
  XOR2X1 U2477 ( .A(n3165), .B(n1949), .Y(n3164) );
  XOR2X1 U2478 ( .A(n930), .B(n920), .Y(n3165) );
  XOR2X1 U2479 ( .A(n3166), .B(n3167), .Y(n3163) );
  XOR2X1 U2480 ( .A(n3168), .B(n3169), .Y(n3167) );
  XOR2X1 U2481 ( .A(n1919), .B(n1891), .Y(n3169) );
  XOR2X1 U2482 ( .A(n3170), .B(n3171), .Y(n3168) );
  XNOR2X1 U2483 ( .A(n1865), .B(n1819), .Y(n3171) );
  XOR2X1 U2484 ( .A(n3172), .B(n1781), .Y(n3170) );
  XOR2X1 U2485 ( .A(n3173), .B(n1799), .Y(n3172) );
  XOR2X1 U2486 ( .A(n3174), .B(n1771), .Y(n3173) );
  OAI21X1 U2487 ( .A(n3002), .B(n2999), .C(n3135), .Y(n3174) );
  XOR2X1 U2488 ( .A(n1841), .B(n3175), .Y(n3166) );
  XOR2X1 U2489 ( .A(n928), .B(n926), .Y(n3175) );
  XOR2X1 U2490 ( .A(n3176), .B(n918), .Y(n3160) );
  XNOR2X1 U2491 ( .A(n924), .B(n922), .Y(n3176) );
  INVX2 U2492 ( .A(n853), .Y(n901) );
  INVX2 U2493 ( .A(n845), .Y(n899) );
  INVX2 U2494 ( .A(n837), .Y(n897) );
  INVX2 U2495 ( .A(n829), .Y(n895) );
  INVX2 U2496 ( .A(n825), .Y(n894) );
  INVX2 U2497 ( .A(n822), .Y(n893) );
  INVX2 U2498 ( .A(n803), .Y(n890) );
  INVX2 U2499 ( .A(n800), .Y(n889) );
  INVX2 U2500 ( .A(n767), .Y(n884) );
  INVX2 U2501 ( .A(n756), .Y(n882) );
  INVX2 U2502 ( .A(n679), .Y(n873) );
  INVX2 U2503 ( .A(n674), .Y(n872) );
  INVX2 U2504 ( .A(n666), .Y(n871) );
  INVX2 U2505 ( .A(n645), .Y(n868) );
  INVX2 U2506 ( .A(n614), .Y(n865) );
  INVX2 U2507 ( .A(n607), .Y(n864) );
  INVX2 U2508 ( .A(n598), .Y(n863) );
  INVX2 U2509 ( .A(n595), .Y(n862) );
  INVX2 U2510 ( .A(n586), .Y(n861) );
  INVX2 U2511 ( .A(n559), .Y(n858) );
  INVX2 U2512 ( .A(n851), .Y(n849) );
  INVX2 U2513 ( .A(n843), .Y(n841) );
  INVX2 U2514 ( .A(n835), .Y(n833) );
  INVX2 U2515 ( .A(n817), .Y(n815) );
  INVX2 U2516 ( .A(n812), .Y(n810) );
  INVX2 U2517 ( .A(n795), .Y(n793) );
  INVX2 U2518 ( .A(n790), .Y(n788) );
  INVX2 U2519 ( .A(n778), .Y(n780) );
  INVX2 U2520 ( .A(n777), .Y(n886) );
  INVX2 U2521 ( .A(n775), .Y(n773) );
  INVX2 U2522 ( .A(n762), .Y(n760) );
  INVX2 U2523 ( .A(n761), .Y(n883) );
  INVX2 U2524 ( .A(n750), .Y(n752) );
  INVX2 U2525 ( .A(n729), .Y(n731) );
  INVX2 U2526 ( .A(n728), .Y(n879) );
  INVX2 U2527 ( .A(n726), .Y(n724) );
  INVX2 U2528 ( .A(n718), .Y(n720) );
  INVX2 U2529 ( .A(n717), .Y(n719) );
  INVX2 U2530 ( .A(n715), .Y(n713) );
  INVX2 U2531 ( .A(n706), .Y(n704) );
  INVX2 U2532 ( .A(n696), .Y(n694) );
  INVX2 U2533 ( .A(n695), .Y(n875) );
  INVX2 U2534 ( .A(n684), .Y(n686) );
  INVX2 U2535 ( .A(n657), .Y(n655) );
  INVX2 U2536 ( .A(n653), .Y(n651) );
  INVX2 U2537 ( .A(n652), .Y(n869) );
  INVX2 U2538 ( .A(n637), .Y(n639) );
  INVX2 U2539 ( .A(n635), .Y(n633) );
  INVX2 U2540 ( .A(n634), .Y(n867) );
  INVX2 U2541 ( .A(n622), .Y(n624) );
  INVX2 U2542 ( .A(n621), .Y(n623) );
  INVX2 U2543 ( .A(n594), .Y(n592) );
  INVX2 U2544 ( .A(n593), .Y(n591) );
  INVX2 U2545 ( .A(n585), .Y(n583) );
  INVX2 U2546 ( .A(n584), .Y(n582) );
  INVX2 U2547 ( .A(n580), .Y(n578) );
  INVX2 U2548 ( .A(n571), .Y(n569) );
  INVX2 U2549 ( .A(n558), .Y(n556) );
  INVX2 U2550 ( .A(n557), .Y(n555) );
  INVX2 U2551 ( .A(n553), .Y(n551) );
  NAND2X1 U2552 ( .A(n3156), .B(n3059), .Y(n2737) );
  NAND2X1 U2553 ( .A(n3152), .B(n3059), .Y(n2704) );
  NAND2X1 U2554 ( .A(n3150), .B(n3059), .Y(n2671) );
  NAND2X1 U2555 ( .A(n3146), .B(n3059), .Y(n2638) );
  NAND2X1 U2556 ( .A(n3143), .B(n3059), .Y(n2605) );
  NAND2X1 U2557 ( .A(n3140), .B(n3059), .Y(n2572) );
  NAND2X1 U2558 ( .A(n3138), .B(n3059), .Y(n2539) );
  NAND2X1 U2559 ( .A(n3135), .B(n3059), .Y(n2506) );
  NAND2X1 U2560 ( .A(n3131), .B(n3059), .Y(n2473) );
  NAND2X1 U2561 ( .A(n3129), .B(n3059), .Y(n2440) );
  NAND2X1 U2562 ( .A(n3126), .B(n3059), .Y(n2409) );
  NAND2X1 U2563 ( .A(n3123), .B(n3059), .Y(n2380) );
  NAND2X1 U2564 ( .A(n3118), .B(n3058), .Y(n2353) );
  NAND2X1 U2565 ( .A(n3116), .B(n3058), .Y(n2328) );
  NAND2X1 U2566 ( .A(n3113), .B(n3058), .Y(n2305) );
  NAND2X1 U2567 ( .A(n3053), .B(n3058), .Y(n2284) );
  NOR2X1 U2568 ( .A(n3051), .B(n3057), .Y(n2218) );
  OAI21X1 U2569 ( .A(n3001), .B(n2998), .C(n3152), .Y(n2185) );
  NOR2X1 U2570 ( .A(n3050), .B(n3057), .Y(n2184) );
  OAI21X1 U2571 ( .A(n2995), .B(n2996), .C(n3150), .Y(n2151) );
  NOR2X1 U2572 ( .A(n3049), .B(n3057), .Y(n2150) );
  OAI21X1 U2573 ( .A(n3008), .B(n3010), .C(n3146), .Y(n2117) );
  NOR2X1 U2574 ( .A(n3048), .B(n3057), .Y(n2116) );
  OAI21X1 U2575 ( .A(n2994), .B(n2997), .C(n3143), .Y(n2083) );
  NOR2X1 U2576 ( .A(n3047), .B(n3058), .Y(n2082) );
  OAI21X1 U2577 ( .A(n3007), .B(n3011), .C(n3140), .Y(n2049) );
  NOR2X1 U2578 ( .A(n3046), .B(n3058), .Y(n2048) );
  OAI21X1 U2579 ( .A(n3009), .B(n3012), .C(n3138), .Y(n2015) );
  NOR2X1 U2580 ( .A(n3045), .B(n3058), .Y(n2014) );
  NOR2X1 U2581 ( .A(n3044), .B(n3058), .Y(n1980) );
  NOR2X1 U2582 ( .A(n3043), .B(n3058), .Y(n1948) );
  NOR2X1 U2583 ( .A(n3042), .B(n3058), .Y(n1918) );
  NOR2X1 U2584 ( .A(n3041), .B(n3058), .Y(n1890) );
  NOR2X1 U2585 ( .A(n3040), .B(n3058), .Y(n1864) );
  NOR2X1 U2586 ( .A(n2925), .B(n3058), .Y(n1840) );
  NOR2X1 U2587 ( .A(n2926), .B(n3058), .Y(n1818) );
  NOR2X1 U2588 ( .A(n2927), .B(n3058), .Y(n1798) );
  NOR2X1 U2589 ( .A(n3054), .B(n3057), .Y(n1780) );
  INVX2 U2590 ( .A(n1242), .Y(n1274) );
  OAI21X1 U2591 ( .A(b[0]), .B(n3000), .C(n3156), .Y(n1242) );
  INVX2 U2592 ( .A(n1180), .Y(n1181) );
  INVX2 U2593 ( .A(n1122), .Y(n1123) );
  INVX2 U2594 ( .A(n1068), .Y(n1069) );
  INVX2 U2595 ( .A(n1018), .Y(n1019) );
endmodule


module poly5 ( clk, rst, pushin, opin, datain, pushout, dataout );
  input [3:0] opin;
  input [31:0] datain;
  output [31:0] dataout;
  input clk, rst, pushin;
  output pushout;
  wire   pushdata, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500,
         N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511,
         N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, N668, N669, N670, N671, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686,
         N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697,
         N698, N699, N701, N702, N703, N704, N705, N706, N707, N708, N709,
         N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720,
         N721, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731,
         N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742,
         N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753,
         N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N798,
         N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809,
         N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820,
         N821, N822, N823, N824, N825, N826, N827, N829, N830, N831, N832,
         N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843,
         N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854,
         N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865,
         N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876,
         N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889,
         N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900,
         N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N912,
         N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N946, N947, N949, N951, N952, N953, N954, N955, N956, N957, N958,
         N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969,
         N970, N971, N972, N973, N974, N1040, N1041, N1042, N1043, N1044,
         N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054,
         N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064,
         N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074,
         N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084,
         N1085, N1086, N1087, N1090, N1091, N1092, N1093, N1094, N1095, N1096,
         N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106,
         N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116,
         N1117, N1118, N1119, N1120, N1121, N1123, N1124, N1125, N1126, N1127,
         N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137,
         N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147,
         N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157,
         N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167,
         N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177,
         N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1188,
         N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198,
         N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208,
         N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218,
         N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226, N1227, N1228,
         N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238,
         N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248,
         N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258,
         N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268,
         N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278,
         N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288,
         N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298,
         N1299, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310,
         N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320,
         N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330,
         N1331, N1332, N1333, N1335, N1336, N1337, N1338, N1339, N1340, N1341,
         N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351,
         N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361,
         N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371,
         N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381,
         N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391,
         N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1463, N1464, N1465,
         N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473, N1474, N1475,
         N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483, N1484, N1485,
         N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493, N1494, N1495,
         N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503, N1504, N1505,
         N1506, N1507, N1508, N1509, N1510, N1513, N1514, N1515, N1516, N1517,
         N1518, N1519, N1520, N1521, N1522, N1523, N1524, N1525, N1526, N1527,
         N1528, N1529, N1530, N1531, N1532, N1533, N1534, N1535, N1536, N1537,
         N1538, N1539, N1540, N1541, N1542, N1543, N1544, N1546, N1547, N1548,
         N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556, N1557, N1558,
         N1559, N1560, N1561, N1562, N1563, N1564, N1565, N1566, N1567, N1568,
         N1569, N1570, N1571, N1572, N1573, N1574, N1575, N1576, N1577, N1578,
         N1579, N1580, N1581, N1582, N1583, N1584, N1585, N1586, N1587, N1588,
         N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598,
         N1599, N1600, N1601, N1602, N1603, N1604, N1605, N1606, N1607, N1608,
         N1609, N1674, N1675, N1676, N1677, N1678, N1679, N1680, N1681, N1682,
         N1683, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692,
         N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702,
         N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712,
         N1713, N1714, N1715, N1716, N1717, N1718, N1719, N1720, N1721, N1724,
         N1725, N1726, N1727, N1728, N1729, N1730, N1731, N1732, N1733, N1734,
         N1735, N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1743, N1744,
         N1745, N1746, N1747, N1748, N1749, N1750, N1751, N1752, N1753, N1754,
         N1755, N1757, N1758, N1759, N1760, N1761, N1762, N1763, N1764, N1765,
         N1766, N1767, N1768, N1769, N1770, N1771, N1772, N1773, N1774, N1775,
         N1776, N1777, N1778, N1779, N1780, N1781, N1782, N1783, N1784, N1785,
         N1786, N1787, N1788, N1789, N1790, N1791, N1792, N1793, N1794, N1795,
         N1796, N1797, N1798, N1799, N1800, N1801, N1802, N1803, N1804, N1805,
         N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813, N1814, N1815,
         N1816, N1817, N1818, N1819, N1820, N1885, N1886, N1887, N1888, N1889,
         N1890, N1891, N1892, N1893, N1894, N1895, N1896, N1897, N1898, N1899,
         N1900, N1901, N1902, N1903, N1904, N1905, N1906, N1907, N1908, N1909,
         N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917, N1918, N1919,
         N1920, N1921, N1922, N1923, N1924, N1925, N1926, N1927, N1928, N1929,
         N1930, N1931, N1932, N1935, N1936, N1937, N1938, N1939, N1940, N1941,
         N1942, N1943, N1944, N1945, N1946, N1947, N1948, N1949, N1950, N1951,
         N1952, N1953, N1954, N1955, N1956, N1957, N1958, N1959, N1960, N1961,
         N1962, N1963, N1964, N1965, N1966, N1968, N1969, N1970, N1971, N1972,
         N1973, N1974, N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1982,
         N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991, N1992,
         N1993, N1994, N1995, N1996, N1997, N1998, N1999, N2000, N2001, N2002,
         N2003, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012,
         N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022,
         N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2031, N2096,
         N2097, N2098, N2099, N2100, N2101, N2102, N2103, N2104, N2105, N2106,
         N2107, N2108, N2109, N2110, N2111, N2112, N2113, N2114, N2115, N2116,
         N2117, N2118, N2119, N2120, N2121, N2122, N2123, N2124, N2125, N2126,
         N2127, N2128, N2129, N2130, N2131, N2132, N2133, N2134, N2135, N2136,
         N2137, N2138, N2139, N2140, N2141, N2142, N2143, N2146, N2147, N2148,
         N2149, N2150, N2151, N2152, N2153, N2154, N2155, N2156, N2157, N2158,
         N2159, N2160, N2161, N2162, N2163, N2164, N2165, N2166, N2167, N2168,
         N2169, N2170, N2171, N2172, N2173, N2174, N2175, N2176, N2177, n229,
         n230, n268, n307, n510, n511, n513, n577, n610, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n709, n710,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n1219, n1380,
         n1413, n1606, n1607, n1608, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, N2305, N2304, N2303, N2302, N2301, N2300, N2299,
         N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289,
         N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279,
         N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269,
         N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259,
         N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249,
         N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239,
         N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229,
         N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219,
         N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209,
         N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199,
         N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189,
         N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179,
         N2178, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258;
  wire   [31:0] a0;
  wire   [31:0] a1;
  wire   [31:0] a2;
  wire   [31:0] a3;
  wire   [31:0] a4;
  wire   [31:0] a5;
  wire   [31:0] x;
  wire   [31:0] res;
  wire   [31:0] t1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287;

  DFFSR \a4_reg[31]  ( .D(n1380), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[31])
         );
  DFFSR \a4_reg[30]  ( .D(n1828), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[30])
         );
  DFFSR \a4_reg[29]  ( .D(n1827), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[29])
         );
  DFFSR \a4_reg[28]  ( .D(n1826), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[28])
         );
  DFFSR \a4_reg[27]  ( .D(n1825), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[27])
         );
  DFFSR \a4_reg[26]  ( .D(n1824), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[26])
         );
  DFFSR \a4_reg[25]  ( .D(n1823), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[25])
         );
  DFFSR \a4_reg[24]  ( .D(n1822), .CLK(clk), .R(n1945), .S(1'b1), .Q(a4[24])
         );
  DFFSR \a4_reg[23]  ( .D(n1821), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[23])
         );
  DFFSR \a4_reg[22]  ( .D(n1820), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[22])
         );
  DFFSR \a4_reg[21]  ( .D(n1819), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[21])
         );
  DFFSR \a4_reg[20]  ( .D(n1818), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[20])
         );
  DFFSR \a4_reg[19]  ( .D(n1817), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[19])
         );
  DFFSR \a4_reg[18]  ( .D(n1816), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[18])
         );
  DFFSR \a4_reg[17]  ( .D(n1815), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[17])
         );
  DFFSR \a4_reg[16]  ( .D(n1814), .CLK(clk), .R(1'b1), .S(n1956), .Q(a4[16])
         );
  DFFSR \a4_reg[15]  ( .D(n1813), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[15])
         );
  DFFSR \a4_reg[14]  ( .D(n1812), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[14])
         );
  DFFSR \a4_reg[13]  ( .D(n1811), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[13])
         );
  DFFSR \a4_reg[12]  ( .D(n1810), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[12])
         );
  DFFSR \a4_reg[11]  ( .D(n1809), .CLK(clk), .R(n1944), .S(1'b1), .Q(a4[11])
         );
  DFFSR \a4_reg[10]  ( .D(n1808), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[10])
         );
  DFFSR \a4_reg[9]  ( .D(n1807), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[9]) );
  DFFSR \a4_reg[8]  ( .D(n1806), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[8]) );
  DFFSR \a4_reg[7]  ( .D(n1805), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[7]) );
  DFFSR \a4_reg[6]  ( .D(n1804), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[6]) );
  DFFSR \a4_reg[5]  ( .D(n1803), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[5]) );
  DFFSR \a4_reg[4]  ( .D(n1802), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[4]) );
  DFFSR \a4_reg[3]  ( .D(n1801), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[3]) );
  DFFSR \a4_reg[2]  ( .D(n1800), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[2]) );
  DFFSR \a4_reg[1]  ( .D(n1799), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[1]) );
  DFFSR \a4_reg[0]  ( .D(n1798), .CLK(clk), .R(n1943), .S(1'b1), .Q(a4[0]) );
  DFFSR \a5_reg[31]  ( .D(n1413), .CLK(clk), .R(n1943), .S(1'b1), .Q(a5[31])
         );
  DFFSR \a5_reg[30]  ( .D(n1797), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[30])
         );
  DFFSR \a5_reg[29]  ( .D(n1796), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[29])
         );
  DFFSR \a5_reg[28]  ( .D(n1795), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[28])
         );
  DFFSR \a5_reg[27]  ( .D(n1794), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[27])
         );
  DFFSR \a5_reg[26]  ( .D(n1793), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[26])
         );
  DFFSR \a5_reg[25]  ( .D(n1792), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[25])
         );
  DFFSR \a5_reg[24]  ( .D(n1791), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[24])
         );
  DFFSR \a5_reg[23]  ( .D(n1790), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[23])
         );
  DFFSR \a5_reg[22]  ( .D(n1789), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[22])
         );
  DFFSR \a5_reg[21]  ( .D(n1788), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[21])
         );
  DFFSR \a5_reg[20]  ( .D(n1787), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[20])
         );
  DFFSR \a5_reg[19]  ( .D(n1786), .CLK(clk), .R(n1942), .S(1'b1), .Q(a5[19])
         );
  DFFSR \a5_reg[18]  ( .D(n1785), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[18])
         );
  DFFSR \a5_reg[17]  ( .D(n1784), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[17])
         );
  DFFSR \a5_reg[16]  ( .D(n1783), .CLK(clk), .R(1'b1), .S(n1956), .Q(a5[16])
         );
  DFFSR \a5_reg[15]  ( .D(n1782), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[15])
         );
  DFFSR \a5_reg[14]  ( .D(n1781), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[14])
         );
  DFFSR \a5_reg[13]  ( .D(n1780), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[13])
         );
  DFFSR \a5_reg[12]  ( .D(n1779), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[12])
         );
  DFFSR \a5_reg[11]  ( .D(n1778), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[11])
         );
  DFFSR \a5_reg[10]  ( .D(n1777), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[10])
         );
  DFFSR \a5_reg[9]  ( .D(n1776), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[9]) );
  DFFSR \a5_reg[8]  ( .D(n1775), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[8]) );
  DFFSR \a5_reg[7]  ( .D(n1774), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[7]) );
  DFFSR \a5_reg[6]  ( .D(n1773), .CLK(clk), .R(n1941), .S(1'b1), .Q(a5[6]) );
  DFFSR \a5_reg[5]  ( .D(n1772), .CLK(clk), .R(n1940), .S(1'b1), .Q(a5[5]) );
  DFFSR \a5_reg[4]  ( .D(n1771), .CLK(clk), .R(n1940), .S(1'b1), .Q(a5[4]) );
  DFFSR \a5_reg[3]  ( .D(n1770), .CLK(clk), .R(n1940), .S(1'b1), .Q(a5[3]) );
  DFFSR \a5_reg[2]  ( .D(n1769), .CLK(clk), .R(n1940), .S(1'b1), .Q(a5[2]) );
  DFFSR \a5_reg[1]  ( .D(n1768), .CLK(clk), .R(n1940), .S(1'b1), .Q(a5[1]) );
  DFFSR \a5_reg[0]  ( .D(n1767), .CLK(clk), .R(n1940), .S(1'b1), .Q(a5[0]) );
  DFFSR \resq_reg[31]  ( .D(res[31]), .CLK(clk), .R(n1940), .S(1'b1), .Q(
        dataout[31]) );
  DFFSR \resq_reg[30]  ( .D(res[30]), .CLK(clk), .R(n1940), .S(1'b1), .Q(
        dataout[30]) );
  DFFSR \resq_reg[29]  ( .D(res[29]), .CLK(clk), .R(n1940), .S(1'b1), .Q(
        dataout[29]) );
  DFFSR \resq_reg[28]  ( .D(res[28]), .CLK(clk), .R(n1940), .S(1'b1), .Q(
        dataout[28]) );
  DFFSR \resq_reg[27]  ( .D(res[27]), .CLK(clk), .R(n1940), .S(1'b1), .Q(
        dataout[27]) );
  DFFSR \resq_reg[26]  ( .D(res[26]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[26]) );
  DFFSR \resq_reg[25]  ( .D(res[25]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[25]) );
  DFFSR \resq_reg[24]  ( .D(res[24]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[24]) );
  DFFSR \resq_reg[23]  ( .D(res[23]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[23]) );
  DFFSR \resq_reg[22]  ( .D(res[22]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[22]) );
  DFFSR \resq_reg[21]  ( .D(res[21]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[21]) );
  DFFSR \resq_reg[20]  ( .D(res[20]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[20]) );
  DFFSR \resq_reg[19]  ( .D(res[19]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[19]) );
  DFFSR \resq_reg[18]  ( .D(res[18]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[18]) );
  DFFSR \resq_reg[17]  ( .D(res[17]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[17]) );
  DFFSR \resq_reg[16]  ( .D(res[16]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[16]) );
  DFFSR \resq_reg[15]  ( .D(res[15]), .CLK(clk), .R(n1939), .S(1'b1), .Q(
        dataout[15]) );
  DFFSR \resq_reg[14]  ( .D(res[14]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[14]) );
  DFFSR \resq_reg[13]  ( .D(res[13]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[13]) );
  DFFSR \resq_reg[12]  ( .D(res[12]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[12]) );
  DFFSR \resq_reg[11]  ( .D(res[11]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[11]) );
  DFFSR \resq_reg[10]  ( .D(res[10]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[10]) );
  DFFSR \resq_reg[9]  ( .D(res[9]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[9]) );
  DFFSR \resq_reg[8]  ( .D(res[8]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[8]) );
  DFFSR \resq_reg[7]  ( .D(res[7]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[7]) );
  DFFSR \resq_reg[6]  ( .D(res[6]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[6]) );
  DFFSR \resq_reg[5]  ( .D(res[5]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[5]) );
  DFFSR \resq_reg[4]  ( .D(res[4]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[4]) );
  DFFSR \resq_reg[3]  ( .D(res[3]), .CLK(clk), .R(n1938), .S(1'b1), .Q(
        dataout[3]) );
  DFFSR \resq_reg[2]  ( .D(res[2]), .CLK(clk), .R(n1937), .S(1'b1), .Q(
        dataout[2]) );
  DFFSR \resq_reg[1]  ( .D(res[1]), .CLK(clk), .R(n1937), .S(1'b1), .Q(
        dataout[1]) );
  DFFSR \resq_reg[0]  ( .D(res[0]), .CLK(clk), .R(n1937), .S(1'b1), .Q(
        dataout[0]) );
  DFFSR \x_reg[31]  ( .D(n1766), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[31]) );
  DFFSR \x_reg[30]  ( .D(n1765), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[30]) );
  DFFSR \x_reg[29]  ( .D(n1764), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[29]) );
  DFFSR \x_reg[28]  ( .D(n1763), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[28]) );
  DFFSR \x_reg[27]  ( .D(n1762), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[27]) );
  DFFSR \x_reg[26]  ( .D(n1761), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[26]) );
  DFFSR \x_reg[25]  ( .D(n1760), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[25]) );
  DFFSR \x_reg[24]  ( .D(n1759), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[24]) );
  DFFSR \x_reg[23]  ( .D(n1758), .CLK(clk), .R(n1937), .S(1'b1), .Q(x[23]) );
  DFFSR \x_reg[22]  ( .D(n1757), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[22]) );
  DFFSR \x_reg[21]  ( .D(n1756), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[21]) );
  DFFSR \x_reg[20]  ( .D(n1755), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[20]) );
  DFFSR \x_reg[19]  ( .D(n1754), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[19]) );
  DFFSR \x_reg[18]  ( .D(n1753), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[18]) );
  DFFSR \x_reg[17]  ( .D(n1752), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[17]) );
  DFFSR \x_reg[16]  ( .D(n1751), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[16]) );
  DFFSR \x_reg[15]  ( .D(n1750), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[15]) );
  DFFSR \x_reg[14]  ( .D(n1749), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[14]) );
  DFFSR \x_reg[13]  ( .D(n1748), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[13]) );
  DFFSR \x_reg[12]  ( .D(n1747), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[12]) );
  DFFSR \x_reg[11]  ( .D(n1746), .CLK(clk), .R(n1936), .S(1'b1), .Q(x[11]) );
  DFFSR \x_reg[10]  ( .D(n1745), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[10]) );
  DFFSR \x_reg[9]  ( .D(n1744), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[9]) );
  DFFSR \x_reg[8]  ( .D(n1743), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[8]) );
  DFFSR \x_reg[7]  ( .D(n1742), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[7]) );
  DFFSR \x_reg[6]  ( .D(n1741), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[6]) );
  DFFSR \x_reg[5]  ( .D(n1740), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[5]) );
  DFFSR \x_reg[4]  ( .D(n1739), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[4]) );
  DFFSR \x_reg[3]  ( .D(n1738), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[3]) );
  DFFSR \x_reg[2]  ( .D(n1737), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[2]) );
  DFFSR \x_reg[1]  ( .D(n1736), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[1]) );
  DFFSR \x_reg[0]  ( .D(n1735), .CLK(clk), .R(n1935), .S(1'b1), .Q(x[0]) );
  DFFPOSX1 pushdata_reg ( .D(n1850), .CLK(clk), .Q(pushdata) );
  DFFSR pushdataq_reg ( .D(n1847), .CLK(clk), .R(n1940), .S(1'b1), .Q(pushout)
         );
  DFFSR \a0_reg[31]  ( .D(n1734), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[31])
         );
  DFFSR \a0_reg[30]  ( .D(n1733), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[30])
         );
  DFFSR \a0_reg[29]  ( .D(n1732), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[29])
         );
  DFFSR \a0_reg[28]  ( .D(n1731), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[28])
         );
  DFFSR \a0_reg[27]  ( .D(n1730), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[27])
         );
  DFFSR \a0_reg[26]  ( .D(n1729), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[26])
         );
  DFFSR \a0_reg[25]  ( .D(n1728), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[25])
         );
  DFFSR \a0_reg[24]  ( .D(n1727), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[24])
         );
  DFFSR \a0_reg[23]  ( .D(n1726), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[23])
         );
  DFFSR \a0_reg[22]  ( .D(n1725), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[22])
         );
  DFFSR \a0_reg[21]  ( .D(n1724), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[21])
         );
  DFFSR \a0_reg[20]  ( .D(n1723), .CLK(clk), .R(n1955), .S(1'b1), .Q(a0[20])
         );
  DFFSR \a0_reg[19]  ( .D(n1722), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[19])
         );
  DFFSR \a0_reg[18]  ( .D(n1721), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[18])
         );
  DFFSR \a0_reg[17]  ( .D(n1720), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[17])
         );
  DFFSR \a0_reg[16]  ( .D(n1719), .CLK(clk), .R(1'b1), .S(n1956), .Q(a0[16])
         );
  DFFSR \a0_reg[15]  ( .D(n1718), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[15])
         );
  DFFSR \a0_reg[14]  ( .D(n1717), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[14])
         );
  DFFSR \a0_reg[13]  ( .D(n1716), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[13])
         );
  DFFSR \a0_reg[12]  ( .D(n1715), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[12])
         );
  DFFSR \a0_reg[11]  ( .D(n1714), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[11])
         );
  DFFSR \a0_reg[10]  ( .D(n1713), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[10])
         );
  DFFSR \a0_reg[9]  ( .D(n1712), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[9]) );
  DFFSR \a0_reg[8]  ( .D(n1711), .CLK(clk), .R(n1954), .S(1'b1), .Q(a0[8]) );
  DFFSR \a0_reg[7]  ( .D(n1710), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[7]) );
  DFFSR \a0_reg[6]  ( .D(n1709), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[6]) );
  DFFSR \a0_reg[5]  ( .D(n1708), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[5]) );
  DFFSR \a0_reg[4]  ( .D(n1707), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[4]) );
  DFFSR \a0_reg[3]  ( .D(n1706), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[3]) );
  DFFSR \a0_reg[2]  ( .D(n1705), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[2]) );
  DFFSR \a0_reg[1]  ( .D(n1704), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[1]) );
  DFFSR \a0_reg[0]  ( .D(n1703), .CLK(clk), .R(n1953), .S(1'b1), .Q(a0[0]) );
  DFFSR \a1_reg[31]  ( .D(n1606), .CLK(clk), .R(n1953), .S(1'b1), .Q(a1[31])
         );
  DFFSR \a1_reg[30]  ( .D(n1702), .CLK(clk), .R(n1953), .S(1'b1), .Q(a1[30])
         );
  DFFSR \a1_reg[29]  ( .D(n1701), .CLK(clk), .R(n1953), .S(1'b1), .Q(a1[29])
         );
  DFFSR \a1_reg[28]  ( .D(n1700), .CLK(clk), .R(n1953), .S(1'b1), .Q(a1[28])
         );
  DFFSR \a1_reg[27]  ( .D(n1699), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[27])
         );
  DFFSR \a1_reg[26]  ( .D(n1698), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[26])
         );
  DFFSR \a1_reg[25]  ( .D(n1697), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[25])
         );
  DFFSR \a1_reg[24]  ( .D(n1696), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[24])
         );
  DFFSR \a1_reg[23]  ( .D(n1695), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[23])
         );
  DFFSR \a1_reg[22]  ( .D(n1694), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[22])
         );
  DFFSR \a1_reg[21]  ( .D(n1693), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[21])
         );
  DFFSR \a1_reg[20]  ( .D(n1692), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[20])
         );
  DFFSR \a1_reg[19]  ( .D(n1691), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[19])
         );
  DFFSR \a1_reg[18]  ( .D(n1690), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[18])
         );
  DFFSR \a1_reg[17]  ( .D(n1689), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[17])
         );
  DFFSR \a1_reg[16]  ( .D(n1688), .CLK(clk), .R(1'b1), .S(n1955), .Q(a1[16])
         );
  DFFSR \a1_reg[15]  ( .D(n1687), .CLK(clk), .R(n1952), .S(1'b1), .Q(a1[15])
         );
  DFFSR \a1_reg[14]  ( .D(n1686), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[14])
         );
  DFFSR \a1_reg[13]  ( .D(n1685), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[13])
         );
  DFFSR \a1_reg[12]  ( .D(n1684), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[12])
         );
  DFFSR \a1_reg[11]  ( .D(n1683), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[11])
         );
  DFFSR \a1_reg[10]  ( .D(n1682), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[10])
         );
  DFFSR \a1_reg[9]  ( .D(n1681), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[9]) );
  DFFSR \a1_reg[8]  ( .D(n1680), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[8]) );
  DFFSR \a1_reg[7]  ( .D(n1679), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[7]) );
  DFFSR \a1_reg[6]  ( .D(n1678), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[6]) );
  DFFSR \a1_reg[5]  ( .D(n1677), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[5]) );
  DFFSR \a1_reg[4]  ( .D(n1676), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[4]) );
  DFFSR \a1_reg[3]  ( .D(n1675), .CLK(clk), .R(n1951), .S(1'b1), .Q(a1[3]) );
  DFFSR \a1_reg[2]  ( .D(n1674), .CLK(clk), .R(n1950), .S(1'b1), .Q(a1[2]) );
  DFFSR \a1_reg[1]  ( .D(n1673), .CLK(clk), .R(n1950), .S(1'b1), .Q(a1[1]) );
  DFFSR \a1_reg[0]  ( .D(n1672), .CLK(clk), .R(n1950), .S(1'b1), .Q(a1[0]) );
  DFFSR \a2_reg[31]  ( .D(n1607), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[31])
         );
  DFFSR \a2_reg[30]  ( .D(n1671), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[30])
         );
  DFFSR \a2_reg[29]  ( .D(n1670), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[29])
         );
  DFFSR \a2_reg[28]  ( .D(n1669), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[28])
         );
  DFFSR \a2_reg[27]  ( .D(n1668), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[27])
         );
  DFFSR \a2_reg[26]  ( .D(n1667), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[26])
         );
  DFFSR \a2_reg[25]  ( .D(n1666), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[25])
         );
  DFFSR \a2_reg[24]  ( .D(n1665), .CLK(clk), .R(n1950), .S(1'b1), .Q(a2[24])
         );
  DFFSR \a2_reg[23]  ( .D(n1664), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[23])
         );
  DFFSR \a2_reg[22]  ( .D(n1663), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[22])
         );
  DFFSR \a2_reg[21]  ( .D(n1662), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[21])
         );
  DFFSR \a2_reg[20]  ( .D(n1661), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[20])
         );
  DFFSR \a2_reg[19]  ( .D(n1660), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[19])
         );
  DFFSR \a2_reg[18]  ( .D(n1659), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[18])
         );
  DFFSR \a2_reg[17]  ( .D(n1658), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[17])
         );
  DFFSR \a2_reg[16]  ( .D(n1657), .CLK(clk), .R(1'b1), .S(n1955), .Q(a2[16])
         );
  DFFSR \a2_reg[15]  ( .D(n1656), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[15])
         );
  DFFSR \a2_reg[14]  ( .D(n1655), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[14])
         );
  DFFSR \a2_reg[13]  ( .D(n1654), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[13])
         );
  DFFSR \a2_reg[12]  ( .D(n1653), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[12])
         );
  DFFSR \a2_reg[11]  ( .D(n1652), .CLK(clk), .R(n1949), .S(1'b1), .Q(a2[11])
         );
  DFFSR \a2_reg[10]  ( .D(n1651), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[10])
         );
  DFFSR \a2_reg[9]  ( .D(n1650), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[9]) );
  DFFSR \a2_reg[8]  ( .D(n1649), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[8]) );
  DFFSR \a2_reg[7]  ( .D(n1648), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[7]) );
  DFFSR \a2_reg[6]  ( .D(n1647), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[6]) );
  DFFSR \a2_reg[5]  ( .D(n1646), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[5]) );
  DFFSR \a2_reg[4]  ( .D(n1645), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[4]) );
  DFFSR \a2_reg[3]  ( .D(n1644), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[3]) );
  DFFSR \a2_reg[2]  ( .D(n1643), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[2]) );
  DFFSR \a2_reg[1]  ( .D(n1642), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[1]) );
  DFFSR \a2_reg[0]  ( .D(n1641), .CLK(clk), .R(n1948), .S(1'b1), .Q(a2[0]) );
  DFFSR \a3_reg[31]  ( .D(n1608), .CLK(clk), .R(n1948), .S(1'b1), .Q(a3[31])
         );
  DFFSR \a3_reg[30]  ( .D(n1640), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[30])
         );
  DFFSR \a3_reg[29]  ( .D(n1639), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[29])
         );
  DFFSR \a3_reg[28]  ( .D(n1638), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[28])
         );
  DFFSR \a3_reg[27]  ( .D(n1637), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[27])
         );
  DFFSR \a3_reg[26]  ( .D(n1636), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[26])
         );
  DFFSR \a3_reg[25]  ( .D(n1635), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[25])
         );
  DFFSR \a3_reg[24]  ( .D(n1634), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[24])
         );
  DFFSR \a3_reg[23]  ( .D(n1633), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[23])
         );
  DFFSR \a3_reg[22]  ( .D(n1632), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[22])
         );
  DFFSR \a3_reg[21]  ( .D(n1631), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[21])
         );
  DFFSR \a3_reg[20]  ( .D(n1630), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[20])
         );
  DFFSR \a3_reg[19]  ( .D(n1629), .CLK(clk), .R(n1947), .S(1'b1), .Q(a3[19])
         );
  DFFSR \a3_reg[18]  ( .D(n1628), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[18])
         );
  DFFSR \a3_reg[17]  ( .D(n1627), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[17])
         );
  DFFSR \a3_reg[16]  ( .D(n1626), .CLK(clk), .R(1'b1), .S(n1956), .Q(a3[16])
         );
  DFFSR \a3_reg[15]  ( .D(n1625), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[15])
         );
  DFFSR \a3_reg[14]  ( .D(n1624), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[14])
         );
  DFFSR \a3_reg[13]  ( .D(n1623), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[13])
         );
  DFFSR \a3_reg[12]  ( .D(n1622), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[12])
         );
  DFFSR \a3_reg[11]  ( .D(n1621), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[11])
         );
  DFFSR \a3_reg[10]  ( .D(n1620), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[10])
         );
  DFFSR \a3_reg[9]  ( .D(n1619), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[9]) );
  DFFSR \a3_reg[8]  ( .D(n1618), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[8]) );
  DFFSR \a3_reg[7]  ( .D(n1617), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[7]) );
  DFFSR \a3_reg[6]  ( .D(n1616), .CLK(clk), .R(n1946), .S(1'b1), .Q(a3[6]) );
  DFFSR \a3_reg[5]  ( .D(n1615), .CLK(clk), .R(n1945), .S(1'b1), .Q(a3[5]) );
  DFFSR \a3_reg[4]  ( .D(n1614), .CLK(clk), .R(n1945), .S(1'b1), .Q(a3[4]) );
  DFFSR \a3_reg[3]  ( .D(n1613), .CLK(clk), .R(n1945), .S(1'b1), .Q(a3[3]) );
  DFFSR \a3_reg[2]  ( .D(n1612), .CLK(clk), .R(n1945), .S(1'b1), .Q(a3[2]) );
  DFFSR \a3_reg[1]  ( .D(n1611), .CLK(clk), .R(n1950), .S(1'b1), .Q(a3[1]) );
  DFFSR \a3_reg[0]  ( .D(n1610), .CLK(clk), .R(n1935), .S(1'b1), .Q(a3[0]) );
  OAI21X1 U3 ( .A(n1849), .B(n1998), .C(n230), .Y(n1219) );
  NAND2X1 U4 ( .A(pushdata), .B(n1849), .Y(n230) );
  OAI22X1 U89 ( .A(n1995), .B(n2040), .C(n268), .D(n3072), .Y(n1380) );
  OAI22X1 U157 ( .A(n1987), .B(n2038), .C(n3072), .D(n1981), .Y(n1413) );
  OAI22X1 U450 ( .A(n1979), .B(n2045), .C(n3072), .D(n1973), .Y(n1606) );
  OAI22X1 U452 ( .A(n1972), .B(n2044), .C(n3072), .D(n1966), .Y(n1607) );
  OAI22X1 U454 ( .A(n1965), .B(n2042), .C(n3072), .D(n1959), .Y(n1608) );
  OAI22X1 U457 ( .A(n1965), .B(n3258), .C(n1959), .D(n3103), .Y(n1610) );
  OAI22X1 U458 ( .A(n1965), .B(n3257), .C(n1959), .D(n3102), .Y(n1611) );
  OAI22X1 U459 ( .A(n1965), .B(n3256), .C(n1959), .D(n3101), .Y(n1612) );
  OAI22X1 U460 ( .A(n1964), .B(n3255), .C(n1959), .D(n3100), .Y(n1613) );
  OAI22X1 U461 ( .A(n1964), .B(n3254), .C(n1959), .D(n3099), .Y(n1614) );
  OAI22X1 U462 ( .A(n1964), .B(n3253), .C(n1959), .D(n3098), .Y(n1615) );
  OAI22X1 U463 ( .A(n1964), .B(n3252), .C(n1959), .D(n3097), .Y(n1616) );
  OAI22X1 U464 ( .A(n1964), .B(n3251), .C(n1959), .D(n3096), .Y(n1617) );
  OAI22X1 U465 ( .A(n1964), .B(n3250), .C(n1959), .D(n3095), .Y(n1618) );
  OAI22X1 U466 ( .A(n1964), .B(n3249), .C(n1959), .D(n3094), .Y(n1619) );
  OAI22X1 U467 ( .A(n1964), .B(n3248), .C(n1959), .D(n3093), .Y(n1620) );
  OAI22X1 U468 ( .A(n1963), .B(n3247), .C(n1959), .D(n3092), .Y(n1621) );
  OAI22X1 U469 ( .A(n1963), .B(n3246), .C(n1959), .D(n3091), .Y(n1622) );
  OAI22X1 U470 ( .A(n1963), .B(n3245), .C(n1959), .D(n3090), .Y(n1623) );
  OAI22X1 U471 ( .A(n1963), .B(n3244), .C(n1959), .D(n3089), .Y(n1624) );
  OAI22X1 U472 ( .A(n1963), .B(n3243), .C(n1959), .D(n3088), .Y(n1625) );
  OAI22X1 U473 ( .A(n1963), .B(n3242), .C(n1959), .D(n3087), .Y(n1626) );
  OAI22X1 U474 ( .A(n1963), .B(n3241), .C(n1959), .D(n3086), .Y(n1627) );
  OAI22X1 U475 ( .A(n1963), .B(n3240), .C(n1959), .D(n3085), .Y(n1628) );
  OAI22X1 U476 ( .A(n1962), .B(n3239), .C(n1959), .D(n3084), .Y(n1629) );
  OAI22X1 U477 ( .A(n1962), .B(n3238), .C(n1959), .D(n3083), .Y(n1630) );
  OAI22X1 U478 ( .A(n1962), .B(n3237), .C(n1959), .D(n3082), .Y(n1631) );
  OAI22X1 U479 ( .A(n1962), .B(n3236), .C(n1959), .D(n3081), .Y(n1632) );
  OAI22X1 U480 ( .A(n1961), .B(n3235), .C(n1959), .D(n3080), .Y(n1633) );
  OAI22X1 U481 ( .A(n1961), .B(n3234), .C(n1959), .D(n3079), .Y(n1634) );
  OAI22X1 U482 ( .A(n1961), .B(n3233), .C(n1959), .D(n3078), .Y(n1635) );
  OAI22X1 U483 ( .A(n1961), .B(n3232), .C(n1959), .D(n3077), .Y(n1636) );
  OAI22X1 U484 ( .A(n1960), .B(n3231), .C(n1959), .D(n3076), .Y(n1637) );
  OAI22X1 U485 ( .A(n1960), .B(n3230), .C(n1959), .D(n3075), .Y(n1638) );
  OAI22X1 U486 ( .A(n1960), .B(n3229), .C(n1959), .D(n3074), .Y(n1639) );
  OAI22X1 U487 ( .A(n1960), .B(n3228), .C(n1959), .D(n3073), .Y(n1640) );
  NOR2X1 U489 ( .A(n577), .B(n3071), .Y(n513) );
  OAI22X1 U490 ( .A(n1972), .B(n3227), .C(n1966), .D(n3103), .Y(n1641) );
  OAI22X1 U491 ( .A(n1972), .B(n3226), .C(n1966), .D(n3102), .Y(n1642) );
  OAI22X1 U492 ( .A(n1972), .B(n3225), .C(n1966), .D(n3101), .Y(n1643) );
  OAI22X1 U493 ( .A(n1971), .B(n3224), .C(n1966), .D(n3100), .Y(n1644) );
  OAI22X1 U494 ( .A(n1971), .B(n3223), .C(n1966), .D(n3099), .Y(n1645) );
  OAI22X1 U495 ( .A(n1971), .B(n3222), .C(n1966), .D(n3098), .Y(n1646) );
  OAI22X1 U496 ( .A(n1971), .B(n3221), .C(n1966), .D(n3097), .Y(n1647) );
  OAI22X1 U497 ( .A(n1971), .B(n3220), .C(n1966), .D(n3096), .Y(n1648) );
  OAI22X1 U498 ( .A(n1971), .B(n3219), .C(n1966), .D(n3095), .Y(n1649) );
  OAI22X1 U499 ( .A(n1971), .B(n3218), .C(n1966), .D(n3094), .Y(n1650) );
  OAI22X1 U500 ( .A(n1971), .B(n3217), .C(n1966), .D(n3093), .Y(n1651) );
  OAI22X1 U501 ( .A(n1970), .B(n3216), .C(n1966), .D(n3092), .Y(n1652) );
  OAI22X1 U502 ( .A(n1970), .B(n3215), .C(n1966), .D(n3091), .Y(n1653) );
  OAI22X1 U503 ( .A(n1970), .B(n3214), .C(n1966), .D(n3090), .Y(n1654) );
  OAI22X1 U504 ( .A(n1970), .B(n3213), .C(n1966), .D(n3089), .Y(n1655) );
  OAI22X1 U505 ( .A(n1970), .B(n3212), .C(n1966), .D(n3088), .Y(n1656) );
  OAI22X1 U506 ( .A(n1970), .B(n3211), .C(n1966), .D(n3087), .Y(n1657) );
  OAI22X1 U507 ( .A(n1970), .B(n3210), .C(n1966), .D(n3086), .Y(n1658) );
  OAI22X1 U508 ( .A(n1970), .B(n3209), .C(n1966), .D(n3085), .Y(n1659) );
  OAI22X1 U509 ( .A(n1969), .B(n3208), .C(n1966), .D(n3084), .Y(n1660) );
  OAI22X1 U510 ( .A(n1969), .B(n3207), .C(n1966), .D(n3083), .Y(n1661) );
  OAI22X1 U511 ( .A(n1969), .B(n3206), .C(n1966), .D(n3082), .Y(n1662) );
  OAI22X1 U512 ( .A(n1969), .B(n3205), .C(n1966), .D(n3081), .Y(n1663) );
  OAI22X1 U513 ( .A(n1968), .B(n3204), .C(n1966), .D(n3080), .Y(n1664) );
  OAI22X1 U514 ( .A(n1968), .B(n3203), .C(n1966), .D(n3079), .Y(n1665) );
  OAI22X1 U515 ( .A(n1968), .B(n3202), .C(n1966), .D(n3078), .Y(n1666) );
  OAI22X1 U516 ( .A(n1968), .B(n3201), .C(n1966), .D(n3077), .Y(n1667) );
  OAI22X1 U517 ( .A(n1967), .B(n3200), .C(n1966), .D(n3076), .Y(n1668) );
  OAI22X1 U518 ( .A(n1967), .B(n3199), .C(n1966), .D(n3075), .Y(n1669) );
  OAI22X1 U519 ( .A(n1967), .B(n3198), .C(n1966), .D(n3074), .Y(n1670) );
  OAI22X1 U520 ( .A(n1967), .B(n3197), .C(n1966), .D(n3073), .Y(n1671) );
  NOR2X1 U522 ( .A(n577), .B(opin[0]), .Y(n511) );
  NAND3X1 U523 ( .A(pushin), .B(opin[1]), .C(n610), .Y(n577) );
  NOR2X1 U524 ( .A(opin[3]), .B(opin[2]), .Y(n610) );
  OAI22X1 U525 ( .A(n1979), .B(n3196), .C(n1973), .D(n3103), .Y(n1672) );
  OAI22X1 U526 ( .A(n1979), .B(n3195), .C(n1973), .D(n3102), .Y(n1673) );
  OAI22X1 U527 ( .A(n1979), .B(n3194), .C(n1973), .D(n3101), .Y(n1674) );
  OAI22X1 U528 ( .A(n1978), .B(n3193), .C(n1973), .D(n3100), .Y(n1675) );
  OAI22X1 U529 ( .A(n1978), .B(n3192), .C(n1973), .D(n3099), .Y(n1676) );
  OAI22X1 U530 ( .A(n1978), .B(n3191), .C(n1973), .D(n3098), .Y(n1677) );
  OAI22X1 U531 ( .A(n1978), .B(n3190), .C(n1973), .D(n3097), .Y(n1678) );
  OAI22X1 U532 ( .A(n1978), .B(n3189), .C(n1973), .D(n3096), .Y(n1679) );
  OAI22X1 U533 ( .A(n1978), .B(n3188), .C(n1973), .D(n3095), .Y(n1680) );
  OAI22X1 U534 ( .A(n1978), .B(n3187), .C(n1973), .D(n3094), .Y(n1681) );
  OAI22X1 U535 ( .A(n1978), .B(n3186), .C(n1973), .D(n3093), .Y(n1682) );
  OAI22X1 U536 ( .A(n1977), .B(n3185), .C(n1973), .D(n3092), .Y(n1683) );
  OAI22X1 U537 ( .A(n1977), .B(n3184), .C(n510), .D(n3091), .Y(n1684) );
  OAI22X1 U538 ( .A(n1977), .B(n3183), .C(n510), .D(n3090), .Y(n1685) );
  OAI22X1 U539 ( .A(n1977), .B(n3182), .C(n510), .D(n3089), .Y(n1686) );
  OAI22X1 U540 ( .A(n1977), .B(n3181), .C(n510), .D(n3088), .Y(n1687) );
  OAI22X1 U541 ( .A(n1977), .B(n3180), .C(n510), .D(n3087), .Y(n1688) );
  OAI22X1 U542 ( .A(n1977), .B(n3179), .C(n510), .D(n3086), .Y(n1689) );
  OAI22X1 U543 ( .A(n1977), .B(n3178), .C(n510), .D(n3085), .Y(n1690) );
  OAI22X1 U544 ( .A(n1976), .B(n3177), .C(n510), .D(n3084), .Y(n1691) );
  OAI22X1 U545 ( .A(n1976), .B(n3176), .C(n510), .D(n3083), .Y(n1692) );
  OAI22X1 U546 ( .A(n1976), .B(n3175), .C(n510), .D(n3082), .Y(n1693) );
  OAI22X1 U547 ( .A(n1976), .B(n3174), .C(n510), .D(n3081), .Y(n1694) );
  OAI22X1 U548 ( .A(n1975), .B(n3173), .C(n510), .D(n3080), .Y(n1695) );
  OAI22X1 U549 ( .A(n1975), .B(n3172), .C(n510), .D(n3079), .Y(n1696) );
  OAI22X1 U550 ( .A(n1975), .B(n3171), .C(n510), .D(n3078), .Y(n1697) );
  OAI22X1 U551 ( .A(n1975), .B(n3170), .C(n510), .D(n3077), .Y(n1698) );
  OAI22X1 U552 ( .A(n1974), .B(n3169), .C(n1973), .D(n3076), .Y(n1699) );
  OAI22X1 U553 ( .A(n1974), .B(n3168), .C(n510), .D(n3075), .Y(n1700) );
  OAI22X1 U554 ( .A(n1974), .B(n3167), .C(n1973), .D(n3074), .Y(n1701) );
  OAI22X1 U555 ( .A(n1974), .B(n3166), .C(n1973), .D(n3073), .Y(n1702) );
  NAND3X1 U557 ( .A(opin[0]), .B(n3070), .C(n643), .Y(n510) );
  OAI21X1 U558 ( .A(n3103), .B(n1957), .C(n645), .Y(n1703) );
  NAND2X1 U559 ( .A(a0[0]), .B(n1957), .Y(n645) );
  OAI21X1 U560 ( .A(n3102), .B(n1957), .C(n646), .Y(n1704) );
  NAND2X1 U561 ( .A(a0[1]), .B(n644), .Y(n646) );
  OAI21X1 U562 ( .A(n3101), .B(n1957), .C(n647), .Y(n1705) );
  NAND2X1 U563 ( .A(a0[2]), .B(n1957), .Y(n647) );
  OAI21X1 U564 ( .A(n3100), .B(n1957), .C(n648), .Y(n1706) );
  NAND2X1 U565 ( .A(a0[3]), .B(n644), .Y(n648) );
  OAI21X1 U566 ( .A(n3099), .B(n1957), .C(n649), .Y(n1707) );
  NAND2X1 U567 ( .A(a0[4]), .B(n644), .Y(n649) );
  OAI21X1 U568 ( .A(n3098), .B(n1957), .C(n650), .Y(n1708) );
  NAND2X1 U569 ( .A(a0[5]), .B(n644), .Y(n650) );
  OAI21X1 U570 ( .A(n3097), .B(n1957), .C(n651), .Y(n1709) );
  NAND2X1 U571 ( .A(a0[6]), .B(n644), .Y(n651) );
  OAI21X1 U572 ( .A(n3096), .B(n1957), .C(n652), .Y(n1710) );
  NAND2X1 U573 ( .A(a0[7]), .B(n644), .Y(n652) );
  OAI21X1 U574 ( .A(n3095), .B(n1957), .C(n653), .Y(n1711) );
  NAND2X1 U575 ( .A(a0[8]), .B(n644), .Y(n653) );
  OAI21X1 U576 ( .A(n3094), .B(n1957), .C(n654), .Y(n1712) );
  NAND2X1 U577 ( .A(a0[9]), .B(n644), .Y(n654) );
  OAI21X1 U578 ( .A(n3093), .B(n1957), .C(n655), .Y(n1713) );
  NAND2X1 U579 ( .A(a0[10]), .B(n644), .Y(n655) );
  OAI21X1 U580 ( .A(n3092), .B(n1957), .C(n656), .Y(n1714) );
  NAND2X1 U581 ( .A(a0[11]), .B(n644), .Y(n656) );
  OAI21X1 U582 ( .A(n3091), .B(n1957), .C(n657), .Y(n1715) );
  NAND2X1 U583 ( .A(a0[12]), .B(n644), .Y(n657) );
  OAI21X1 U584 ( .A(n3090), .B(n1957), .C(n658), .Y(n1716) );
  NAND2X1 U585 ( .A(a0[13]), .B(n644), .Y(n658) );
  OAI21X1 U586 ( .A(n3089), .B(n1957), .C(n659), .Y(n1717) );
  NAND2X1 U587 ( .A(a0[14]), .B(n644), .Y(n659) );
  OAI21X1 U588 ( .A(n3088), .B(n1957), .C(n660), .Y(n1718) );
  NAND2X1 U589 ( .A(a0[15]), .B(n644), .Y(n660) );
  OAI21X1 U590 ( .A(n3087), .B(n1957), .C(n661), .Y(n1719) );
  NAND2X1 U591 ( .A(a0[16]), .B(n644), .Y(n661) );
  OAI21X1 U592 ( .A(n3086), .B(n1957), .C(n662), .Y(n1720) );
  NAND2X1 U593 ( .A(a0[17]), .B(n644), .Y(n662) );
  OAI21X1 U594 ( .A(n3085), .B(n1957), .C(n663), .Y(n1721) );
  NAND2X1 U595 ( .A(a0[18]), .B(n644), .Y(n663) );
  OAI21X1 U596 ( .A(n3084), .B(n1957), .C(n664), .Y(n1722) );
  NAND2X1 U597 ( .A(a0[19]), .B(n644), .Y(n664) );
  OAI21X1 U598 ( .A(n3083), .B(n1957), .C(n665), .Y(n1723) );
  NAND2X1 U599 ( .A(a0[20]), .B(n644), .Y(n665) );
  OAI21X1 U600 ( .A(n3082), .B(n1957), .C(n666), .Y(n1724) );
  NAND2X1 U601 ( .A(a0[21]), .B(n1957), .Y(n666) );
  OAI21X1 U602 ( .A(n3081), .B(n1957), .C(n667), .Y(n1725) );
  NAND2X1 U603 ( .A(a0[22]), .B(n644), .Y(n667) );
  OAI21X1 U604 ( .A(n3080), .B(n644), .C(n668), .Y(n1726) );
  NAND2X1 U605 ( .A(a0[23]), .B(n1957), .Y(n668) );
  OAI21X1 U606 ( .A(n3079), .B(n1957), .C(n669), .Y(n1727) );
  NAND2X1 U607 ( .A(a0[24]), .B(n644), .Y(n669) );
  OAI21X1 U608 ( .A(n3078), .B(n644), .C(n670), .Y(n1728) );
  NAND2X1 U609 ( .A(a0[25]), .B(n644), .Y(n670) );
  OAI21X1 U610 ( .A(n3077), .B(n644), .C(n671), .Y(n1729) );
  NAND2X1 U611 ( .A(a0[26]), .B(n644), .Y(n671) );
  OAI21X1 U612 ( .A(n3076), .B(n1957), .C(n672), .Y(n1730) );
  NAND2X1 U613 ( .A(a0[27]), .B(n644), .Y(n672) );
  OAI21X1 U614 ( .A(n3075), .B(n644), .C(n673), .Y(n1731) );
  NAND2X1 U615 ( .A(a0[28]), .B(n644), .Y(n673) );
  OAI21X1 U616 ( .A(n3074), .B(n644), .C(n674), .Y(n1732) );
  NAND2X1 U617 ( .A(a0[29]), .B(n1957), .Y(n674) );
  OAI21X1 U618 ( .A(n3073), .B(n644), .C(n675), .Y(n1733) );
  NAND2X1 U619 ( .A(a0[30]), .B(n1957), .Y(n675) );
  OAI21X1 U620 ( .A(n3072), .B(n644), .C(n676), .Y(n1734) );
  NAND2X1 U621 ( .A(a0[31]), .B(n644), .Y(n676) );
  NAND3X1 U622 ( .A(n3071), .B(n3070), .C(n643), .Y(n644) );
  NAND3X1 U657 ( .A(pushin), .B(opin[3]), .C(n709), .Y(n229) );
  NOR2X1 U658 ( .A(n3070), .B(n710), .Y(n709) );
  NAND2X1 U659 ( .A(opin[1]), .B(opin[0]), .Y(n710) );
  OAI22X1 U661 ( .A(n1987), .B(n3165), .C(n1981), .D(n3103), .Y(n1767) );
  OAI22X1 U662 ( .A(n1987), .B(n3164), .C(n1981), .D(n3102), .Y(n1768) );
  OAI22X1 U663 ( .A(n1987), .B(n3163), .C(n1981), .D(n3101), .Y(n1769) );
  OAI22X1 U664 ( .A(n1986), .B(n3162), .C(n1981), .D(n3100), .Y(n1770) );
  OAI22X1 U665 ( .A(n1986), .B(n3161), .C(n1981), .D(n3099), .Y(n1771) );
  OAI22X1 U666 ( .A(n1986), .B(n3160), .C(n1981), .D(n3098), .Y(n1772) );
  OAI22X1 U667 ( .A(n1986), .B(n3159), .C(n1981), .D(n3097), .Y(n1773) );
  OAI22X1 U668 ( .A(n1986), .B(n3158), .C(n1981), .D(n3096), .Y(n1774) );
  OAI22X1 U669 ( .A(n1986), .B(n3157), .C(n1981), .D(n3095), .Y(n1775) );
  OAI22X1 U670 ( .A(n1986), .B(n3156), .C(n1981), .D(n3094), .Y(n1776) );
  OAI22X1 U671 ( .A(n1986), .B(n3155), .C(n1981), .D(n3093), .Y(n1777) );
  OAI22X1 U672 ( .A(n1985), .B(n3154), .C(n1981), .D(n3092), .Y(n1778) );
  OAI22X1 U673 ( .A(n1985), .B(n3153), .C(n307), .D(n3091), .Y(n1779) );
  OAI22X1 U674 ( .A(n1985), .B(n3152), .C(n307), .D(n3090), .Y(n1780) );
  OAI22X1 U675 ( .A(n1985), .B(n3151), .C(n307), .D(n3089), .Y(n1781) );
  OAI22X1 U676 ( .A(n1985), .B(n3150), .C(n307), .D(n3088), .Y(n1782) );
  OAI22X1 U677 ( .A(n1985), .B(n3149), .C(n307), .D(n3087), .Y(n1783) );
  OAI22X1 U678 ( .A(n1985), .B(n3148), .C(n307), .D(n3086), .Y(n1784) );
  OAI22X1 U679 ( .A(n1985), .B(n3147), .C(n307), .D(n3085), .Y(n1785) );
  OAI22X1 U680 ( .A(n1984), .B(n3146), .C(n307), .D(n3084), .Y(n1786) );
  OAI22X1 U681 ( .A(n1984), .B(n3145), .C(n307), .D(n3083), .Y(n1787) );
  OAI22X1 U682 ( .A(n1984), .B(n3144), .C(n307), .D(n3082), .Y(n1788) );
  OAI22X1 U683 ( .A(n1984), .B(n3143), .C(n307), .D(n3081), .Y(n1789) );
  OAI22X1 U684 ( .A(n1983), .B(n3142), .C(n307), .D(n3080), .Y(n1790) );
  OAI22X1 U685 ( .A(n1983), .B(n3141), .C(n307), .D(n3079), .Y(n1791) );
  OAI22X1 U686 ( .A(n1983), .B(n3140), .C(n307), .D(n3078), .Y(n1792) );
  OAI22X1 U687 ( .A(n1983), .B(n3139), .C(n307), .D(n3077), .Y(n1793) );
  OAI22X1 U688 ( .A(n1982), .B(n3138), .C(n1981), .D(n3076), .Y(n1794) );
  OAI22X1 U689 ( .A(n1982), .B(n3137), .C(n307), .D(n3075), .Y(n1795) );
  OAI22X1 U690 ( .A(n1982), .B(n3136), .C(n1981), .D(n3074), .Y(n1796) );
  OAI22X1 U691 ( .A(n1982), .B(n3135), .C(n1981), .D(n3073), .Y(n1797) );
  NAND3X1 U693 ( .A(opin[2]), .B(opin[0]), .C(n643), .Y(n307) );
  OAI22X1 U694 ( .A(n1995), .B(n3134), .C(n1989), .D(n3103), .Y(n1798) );
  OAI22X1 U696 ( .A(n1995), .B(n3133), .C(n1989), .D(n3102), .Y(n1799) );
  OAI22X1 U698 ( .A(n1995), .B(n3132), .C(n268), .D(n3101), .Y(n1800) );
  OAI22X1 U700 ( .A(n1994), .B(n3131), .C(n268), .D(n3100), .Y(n1801) );
  OAI22X1 U702 ( .A(n1994), .B(n3130), .C(n1989), .D(n3099), .Y(n1802) );
  OAI22X1 U704 ( .A(n1994), .B(n3129), .C(n268), .D(n3098), .Y(n1803) );
  OAI22X1 U706 ( .A(n1994), .B(n3128), .C(n1989), .D(n3097), .Y(n1804) );
  OAI22X1 U708 ( .A(n1994), .B(n3127), .C(n268), .D(n3096), .Y(n1805) );
  OAI22X1 U710 ( .A(n1994), .B(n3126), .C(n268), .D(n3095), .Y(n1806) );
  OAI22X1 U712 ( .A(n1994), .B(n3125), .C(n268), .D(n3094), .Y(n1807) );
  OAI22X1 U714 ( .A(n1994), .B(n3124), .C(n268), .D(n3093), .Y(n1808) );
  OAI22X1 U716 ( .A(n1993), .B(n3123), .C(n268), .D(n3092), .Y(n1809) );
  OAI22X1 U718 ( .A(n1993), .B(n3122), .C(n268), .D(n3091), .Y(n1810) );
  OAI22X1 U720 ( .A(n1993), .B(n3121), .C(n268), .D(n3090), .Y(n1811) );
  OAI22X1 U722 ( .A(n1993), .B(n3120), .C(n268), .D(n3089), .Y(n1812) );
  OAI22X1 U724 ( .A(n1993), .B(n3119), .C(n268), .D(n3088), .Y(n1813) );
  OAI22X1 U726 ( .A(n1993), .B(n3118), .C(n268), .D(n3087), .Y(n1814) );
  OAI22X1 U728 ( .A(n1993), .B(n3117), .C(n268), .D(n3086), .Y(n1815) );
  OAI22X1 U730 ( .A(n1993), .B(n3116), .C(n268), .D(n3085), .Y(n1816) );
  OAI22X1 U732 ( .A(n1992), .B(n3115), .C(n1989), .D(n3084), .Y(n1817) );
  OAI22X1 U734 ( .A(n1992), .B(n3114), .C(n1989), .D(n3083), .Y(n1818) );
  OAI22X1 U736 ( .A(n1992), .B(n3113), .C(n1989), .D(n3082), .Y(n1819) );
  OAI22X1 U738 ( .A(n1992), .B(n3112), .C(n1989), .D(n3081), .Y(n1820) );
  OAI22X1 U740 ( .A(n1991), .B(n3111), .C(n1989), .D(n3080), .Y(n1821) );
  OAI22X1 U742 ( .A(n1991), .B(n3110), .C(n1989), .D(n3079), .Y(n1822) );
  OAI22X1 U744 ( .A(n1991), .B(n3109), .C(n1989), .D(n3078), .Y(n1823) );
  OAI22X1 U746 ( .A(n1991), .B(n3108), .C(n1989), .D(n3077), .Y(n1824) );
  OAI22X1 U748 ( .A(n1990), .B(n3107), .C(n1989), .D(n3076), .Y(n1825) );
  OAI22X1 U750 ( .A(n1990), .B(n3106), .C(n1989), .D(n3075), .Y(n1826) );
  OAI22X1 U752 ( .A(n1990), .B(n3105), .C(n1989), .D(n3074), .Y(n1827) );
  OAI22X1 U754 ( .A(n1990), .B(n3104), .C(n1989), .D(n3073), .Y(n1828) );
  NAND3X1 U757 ( .A(opin[2]), .B(n3071), .C(n643), .Y(n268) );
  NOR3X1 U758 ( .A(opin[1]), .B(opin[3]), .C(n3069), .Y(n643) );
  OAI21X1 U1110 ( .A(n1911), .B(n3166), .C(n902), .Y(N2030) );
  NAND2X1 U1111 ( .A(N1998), .B(a1[31]), .Y(n902) );
  OAI21X1 U1113 ( .A(n1911), .B(n3167), .C(n903), .Y(N2029) );
  NAND2X1 U1114 ( .A(N1997), .B(a1[31]), .Y(n903) );
  OAI21X1 U1116 ( .A(n1911), .B(n3168), .C(n904), .Y(N2028) );
  NAND2X1 U1117 ( .A(N1996), .B(a1[31]), .Y(n904) );
  OAI21X1 U1119 ( .A(n1911), .B(n3169), .C(n905), .Y(N2027) );
  NAND2X1 U1120 ( .A(N1995), .B(a1[31]), .Y(n905) );
  OAI21X1 U1122 ( .A(n1911), .B(n3170), .C(n906), .Y(N2026) );
  NAND2X1 U1123 ( .A(N1994), .B(a1[31]), .Y(n906) );
  OAI21X1 U1125 ( .A(n1911), .B(n3171), .C(n907), .Y(N2025) );
  NAND2X1 U1126 ( .A(N1993), .B(a1[31]), .Y(n907) );
  OAI21X1 U1128 ( .A(n1911), .B(n3172), .C(n908), .Y(N2024) );
  NAND2X1 U1129 ( .A(N1992), .B(a1[31]), .Y(n908) );
  OAI21X1 U1131 ( .A(n1911), .B(n3173), .C(n909), .Y(N2023) );
  NAND2X1 U1132 ( .A(N1991), .B(a1[31]), .Y(n909) );
  OAI21X1 U1134 ( .A(n1911), .B(n3174), .C(n910), .Y(N2022) );
  NAND2X1 U1135 ( .A(N1990), .B(a1[31]), .Y(n910) );
  OAI21X1 U1137 ( .A(n1911), .B(n3175), .C(n911), .Y(N2021) );
  NAND2X1 U1138 ( .A(N1989), .B(n1911), .Y(n911) );
  OAI21X1 U1140 ( .A(n1911), .B(n3176), .C(n912), .Y(N2020) );
  NAND2X1 U1141 ( .A(N1988), .B(n1911), .Y(n912) );
  OAI21X1 U1143 ( .A(a1[31]), .B(n3177), .C(n913), .Y(N2019) );
  NAND2X1 U1144 ( .A(N1987), .B(n1911), .Y(n913) );
  OAI21X1 U1146 ( .A(a1[31]), .B(n3178), .C(n914), .Y(N2018) );
  NAND2X1 U1147 ( .A(N1986), .B(n1911), .Y(n914) );
  OAI21X1 U1149 ( .A(a1[31]), .B(n3179), .C(n915), .Y(N2017) );
  NAND2X1 U1150 ( .A(N1985), .B(n1911), .Y(n915) );
  OAI21X1 U1152 ( .A(a1[31]), .B(n3180), .C(n916), .Y(N2016) );
  NAND2X1 U1153 ( .A(N1984), .B(n1911), .Y(n916) );
  OAI21X1 U1155 ( .A(a1[31]), .B(n3181), .C(n917), .Y(N2015) );
  NAND2X1 U1156 ( .A(N1983), .B(n1911), .Y(n917) );
  OAI21X1 U1158 ( .A(a1[31]), .B(n3182), .C(n918), .Y(N2014) );
  NAND2X1 U1159 ( .A(N1982), .B(n1911), .Y(n918) );
  OAI21X1 U1161 ( .A(a1[31]), .B(n3183), .C(n919), .Y(N2013) );
  NAND2X1 U1162 ( .A(N1981), .B(n1911), .Y(n919) );
  OAI21X1 U1164 ( .A(a1[31]), .B(n3184), .C(n920), .Y(N2012) );
  NAND2X1 U1165 ( .A(N1980), .B(n1911), .Y(n920) );
  OAI21X1 U1167 ( .A(a1[31]), .B(n3185), .C(n921), .Y(N2011) );
  NAND2X1 U1168 ( .A(N1979), .B(a1[31]), .Y(n921) );
  OAI21X1 U1170 ( .A(n1911), .B(n3186), .C(n922), .Y(N2010) );
  NAND2X1 U1171 ( .A(N1978), .B(n1911), .Y(n922) );
  OAI21X1 U1173 ( .A(a1[31]), .B(n3187), .C(n923), .Y(N2009) );
  NAND2X1 U1174 ( .A(N1977), .B(a1[31]), .Y(n923) );
  OAI21X1 U1176 ( .A(n1911), .B(n3188), .C(n924), .Y(N2008) );
  NAND2X1 U1177 ( .A(N1976), .B(a1[31]), .Y(n924) );
  OAI21X1 U1179 ( .A(a1[31]), .B(n3189), .C(n925), .Y(N2007) );
  NAND2X1 U1180 ( .A(N1975), .B(n1911), .Y(n925) );
  OAI21X1 U1182 ( .A(n1911), .B(n3190), .C(n926), .Y(N2006) );
  NAND2X1 U1183 ( .A(N1974), .B(a1[31]), .Y(n926) );
  OAI21X1 U1185 ( .A(n1911), .B(n3191), .C(n927), .Y(N2005) );
  NAND2X1 U1186 ( .A(N1973), .B(n1911), .Y(n927) );
  OAI21X1 U1188 ( .A(a1[31]), .B(n3192), .C(n928), .Y(N2004) );
  NAND2X1 U1189 ( .A(N1972), .B(n1911), .Y(n928) );
  OAI21X1 U1191 ( .A(n1911), .B(n3193), .C(n929), .Y(N2003) );
  NAND2X1 U1192 ( .A(N1971), .B(n1911), .Y(n929) );
  OAI21X1 U1194 ( .A(n1911), .B(n3194), .C(n930), .Y(N2002) );
  NAND2X1 U1195 ( .A(N1970), .B(a1[31]), .Y(n930) );
  OAI21X1 U1197 ( .A(a1[31]), .B(n3195), .C(n931), .Y(N2001) );
  NAND2X1 U1198 ( .A(N1969), .B(n1911), .Y(n931) );
  OAI21X1 U1200 ( .A(n1911), .B(n3196), .C(n932), .Y(N2000) );
  NAND2X1 U1201 ( .A(N1968), .B(n1911), .Y(n932) );
  AND2X2 U1109 ( .A(N1999), .B(a1[31]), .Y(N2031) );
  poly5_DW01_sub_0 sub_45_S2_C88 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N2143, N2142, N2141, N2140, 
        N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, 
        N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, 
        N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, 
        N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, 
        N2099, N2098, N2097, N2096}), .CI(1'b0), .DIFF({N2177, N2176, N2175, 
        N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, 
        N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, 
        N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15}) );
  poly5_DW01_sub_1 sub_31_C88 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B(a1), .CI(1'b0), .DIFF({N1999, N1998, N1997, N1996, N1995, 
        N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, 
        N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, 
        N1974, N1973, N1972, N1971, N1970, N1969, N1968}) );
  poly5_DW01_sub_2 sub_45_S2_C87 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N1932, N1931, N1930, N1929, 
        N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, 
        N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, 
        N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, 
        N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, 
        N1888, N1887, N1886, N1885}), .CI(1'b0), .DIFF({N1966, N1965, N1964, 
        N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, 
        N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, 
        N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31}) );
  poly5_DW01_sub_3 sub_31_C87 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n2043, a2[30:0]}), .CI(1'b0), .DIFF({N1788, N1787, N1786, 
        N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, 
        N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, 
        N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757}) );
  poly5_DW01_sub_4 sub_45_S2_C86 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N1721, N1720, N1719, N1718, 
        N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, 
        N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, 
        N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, 
        N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, 
        N1677, N1676, N1675, N1674}), .CI(1'b0), .DIFF({N1755, N1754, N1753, 
        N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, 
        N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, 
        N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47}) );
  poly5_DW01_sub_5 sub_31_C86 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n2041, a3[30:0]}), .CI(1'b0), .DIFF({N1577, N1576, N1575, 
        N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, 
        N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, 
        N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546}) );
  poly5_DW01_sub_6 sub_45_S2_C85 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N1510, N1509, N1508, N1507, 
        N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, 
        N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, 
        N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, 
        N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, 
        N1466, N1465, N1464, N1463}), .CI(1'b0), .DIFF({N1544, N1543, N1542, 
        N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, 
        N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, 
        N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63}) );
  poly5_DW01_sub_7 sub_31_C85 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n2039, a4[30:0]}), .CI(1'b0), .DIFF({N1366, N1365, N1364, 
        N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, 
        N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, 
        N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335}) );
  poly5_DW01_sub_10 sub_31_C84 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n2037, a5[30:0]}), .CI(1'b0), .DIFF({N1154, N1153, N1152, 
        N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, 
        N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, 
        N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123}) );
  poly5_DW01_add_4 add_4_root_add_0_root_add_89_5 ( .A(a0), .B({n3064, n3063, 
        n3062, n3061, n3060, n3059, n3058, n3057, n3056, n3055, n3054, n3053, 
        n3052, n3051, n3050, n3049, n3048, n3047, n3046, n3045, n3044, n3043, 
        n3042, n3041, n3040, n3039, n3038, n3037, n3036, n3035, n3034, n3033}), 
        .CI(1'b0), .SUM({N2241, N2240, N2239, N2238, N2237, N2236, N2235, 
        N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, 
        N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, 
        N2214, N2213, N2212, N2211, N2210}) );
  poly5_DW01_add_3 add_3_root_add_0_root_add_89_5 ( .A({N2241, N2240, N2239, 
        N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, 
        N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, 
        N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210}), .B({
        n3002, n3001, n3000, n2999, n2998, n2997, n2996, n2995, n2994, n2993, 
        n2992, n2991, n2990, n2989, n2988, n2987, n2986, n2985, n2984, n2983, 
        n2982, n2981, n2980, n2979, n2978, n2977, n2976, n2975, n2974, n2973, 
        n2972, n2971}), .CI(1'b0), .SUM({N2209, N2208, N2207, N2206, N2205, 
        N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, 
        N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, 
        N2184, N2183, N2182, N2181, N2180, N2179, N2178}) );
  poly5_DW01_add_2 add_2_root_add_0_root_add_89_5 ( .A({N2209, N2208, N2207, 
        N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, 
        N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, 
        N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178}), .B({
        n2939, n2938, n2937, n2936, n2935, n2934, n2933, n2932, n2931, n2930, 
        n2929, n2928, n2927, n2926, n2925, n2924, n2923, n2922, n2921, n2920, 
        n2919, n2918, n2917, n2916, n2915, n2914, n2913, n2912, n2911, n2910, 
        n2909, n2908}), .CI(1'b0), .SUM({N2305, N2304, N2303, N2302, N2301, 
        N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, 
        N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, 
        N2280, N2279, N2278, N2277, N2276, N2275, N2274}) );
  poly5_DW01_add_1 add_1_root_add_0_root_add_89_5 ( .A({N2305, N2304, N2303, 
        N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, 
        N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, 
        N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274}), .B({
        n2876, n2875, n2874, n2873, n2872, n2871, n2870, n2869, n2868, n2867, 
        n2866, n2865, n2864, n2863, n2862, n2861, n2860, n2859, n2858, n2857, 
        n2856, n2855, n2854, n2853, n2852, n2851, n2850, n2849, n2848, n2847, 
        n2846, n2845}), .CI(1'b0), .SUM({N2273, N2272, N2271, N2270, N2269, 
        N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, 
        N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, 
        N2248, N2247, N2246, N2245, N2244, N2243, N2242}) );
  poly5_DW_mult_uns_4 mult_43_C86 ( .a({N1609, N1608, N1607, N1606, N1605, 
        N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, 
        N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, 
        N1584, N1583, N1582, N1581, N1580, N1579, N1578}), .b({n2781, N763, 
        N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, 
        N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, 
        N738, N737, N736, N735, N734, N733}), .product({
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, N1721, N1720, 
        N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, 
        N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, 
        N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, 
        N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, 
        N1679, N1678, N1677, N1676, N1675, N1674}) );
  poly5_DW_mult_uns_3 mult_43_C87 ( .a({N1820, N1819, N1818, N1817, N1816, 
        N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, 
        N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, 
        N1795, N1794, N1793, N1792, N1791, N1790, N1789}), .b({n1833, n3032, 
        n3031, n1835, n3029, n3028, n1861, n3026, n3025, n3024, n3023, n3022, 
        n3021, n3020, n3019, n3018, n3017, n3016, n3015, n3014, n3013, n3012, 
        n3011, n3010, n3009, n3008, n3007, n3006, n3005, n3004, n1921, n3003}), 
        .product({SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, N1932, N1931, 
        N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, 
        N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, 
        N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, 
        N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, 
        N1890, N1889, N1888, N1887, N1886, N1885}) );
  poly5_DW_mult_uns_0 mult_43_C88 ( .a({N2031, N2030, N2029, N2028, N2027, 
        N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, 
        N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, 
        N2006, N2005, N2004, N2003, N2002, N2001, N2000}), .b({n1845, n1830, 
        n2004, n1890, n2006, n1892, n2008, N821, n2010, N819, n2012, N817, 
        n2014, n1852, n2016, N813, n2018, n1891, n1853, N809, n2020, n1855, 
        n2022, N805, n2024, N803, n2026, N801, N800, N799, n2028, n2030}), 
        .product({SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, N2143, N2142, 
        N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, 
        N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, 
        N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, 
        N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, 
        N2101, N2100, N2099, N2098, N2097, N2096}) );
  poly5_DW01_sub_22 r371 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n2034, x[30:17], n1842, x[15:9], n1843, x[7:6], n1885, n1886, n1841, 
        n1884, x[1], n1897}), .CI(1'b0), .DIFF({N310, N309, N308, N307, N306, 
        N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, 
        N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, 
        N281, N280, N279}) );
  poly5_DW01_sub_39 sub_45_S2_C81 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N665, N664, N663, N662, N661, 
        N660, N659, N658, N657, N656, N655, N654, N653, n1864, n1887, N650, 
        N649, n1836, n1882, N646, N645, N644, n1837, N642, N641, N640, N639, 
        N638, N637, n1865, N635, N634, N633, N632, N631, N630, N629, N628, 
        N627, N626, N625, N624, N623, N622, N621, N620, N619, N618}), .CI(1'b0), .DIFF({N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, 
        N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, 
        N676, N675, N674, N673, N672, N671, N670, N669, N668, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127}) );
  poly5_DW01_sub_43 r377 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n1873, n2970, n2969, n2968, n2967, n2966, n2965, n2964, n2963, n2962, 
        n2961, n2960, n2959, n2958, n2957, n2956, n2955, n2954, n2953, n2952, 
        n2951, n2950, n2949, n2948, n2947, n2946, n2945, n2944, n2943, n2942, 
        n2941, n2940}), .CI(1'b0), .DIFF({N732, N731, N730, N729, N728, N727, 
        N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, 
        N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, 
        N702, N701}) );
  poly5_DW_mult_uns_35 mult_43_C82 ( .a({n2781, N763, N762, N761, N760, N759, 
        N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, 
        N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, 
        N734, N733}), .b({n1845, n1830, n2004, n1890, n2006, n1892, n2008, 
        N821, n2010, N819, n2012, N817, n2014, n1852, n2016, N813, n2018, 
        n1891, n1853, N809, n2020, n1855, n2022, N805, n2024, N803, n2026, 
        N801, N800, N799, n2028, n2030}), .product({SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, SYNOPSYS_UNCONNECTED__132, 
        SYNOPSYS_UNCONNECTED__133, SYNOPSYS_UNCONNECTED__134, 
        SYNOPSYS_UNCONNECTED__135, SYNOPSYS_UNCONNECTED__136, 
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, SYNOPSYS_UNCONNECTED__142, 
        SYNOPSYS_UNCONNECTED__143, N876, N875, N874, N873, N872, N871, N870, 
        N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, 
        N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, 
        N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, 
        N833, N832, N831, N830, N829}) );
  poly5_DW01_sub_49 sub_45_S2_C82 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N876, N875, N874, N873, N872, 
        N871, N870, N869, N868, N867, N866, N865, N864, N863, n1840, N861, 
        N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, 
        N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, 
        N836, N835, N834, N833, N832, N831, N830, N829}), .CI(1'b0), .DIFF({
        N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, 
        N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, 
        N886, N885, N884, N883, N882, N881, N880, N879, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159}) );
  poly5_DW01_sub_52 r380 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n1895, n2907, n2906, n2905, n2904, n2903, n2902, n2901, n2900, n2899, 
        n2898, n2897, n2896, n2895, n2894, n2893, n2892, n2891, n2890, n2889, 
        n2888, n2887, n2886, n2885, n2884, n2883, n2882, n2881, n2880, n2879, 
        n2878, n2877}), .CI(1'b0), .DIFF({N943, N942, N941, N940, N939, N938, 
        N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, 
        N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, 
        N913, N912}) );
  poly5_DW_mult_uns_41 mult_43_C83 ( .a({n2780, N974, N973, N972, N971, N970, 
        N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, 
        N957, N956, n1894, N954, N953, N952, N951, n1893, N949, n1854, N947, 
        N946, N945, N944}), .b({n1845, n1830, n2004, n1890, n2006, n1892, 
        n2008, N821, n2010, N819, n2012, N817, n2014, n1852, n2016, N813, 
        n2018, n1891, n1853, N809, n2020, n1855, n2022, N805, n2024, N803, 
        n2026, N801, N800, N799, n2028, n2030}), .product({
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, N1087, N1086, 
        N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, 
        N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, 
        N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, 
        N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, 
        N1045, N1044, N1043, N1042, N1041, N1040}) );
  poly5_DW01_sub_56 sub_45_S2_C83 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N1087, N1086, N1085, n1883, 
        N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, 
        n1844, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, 
        N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, 
        N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, 
        N1043, N1042, N1041, N1040}), .CI(1'b0), .DIFF({N1121, N1120, N1119, 
        N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, 
        N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, 
        N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191}) );
  poly5_DW_mult_uns_43 mult_43_C84 ( .a({N1186, N1185, N1184, N1183, N1182, 
        N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, 
        N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, 
        N1161, N1160, N1159, N1158, N1157, N1156, N1155}), .b({N1251, N1250, 
        N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, 
        N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, 
        N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220}), 
        .product({SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, N1299, N1298, 
        N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, 
        N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, 
        N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, 
        N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, 
        N1257, N1256, N1255, N1254, N1253, N1252}) );
  poly5_DW01_sub_59 sub_38_C84 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n1922, n2844, n2843, n2842, n2841, n2840, n2839, n2838, 
        n2837, n2836, n2835, n2834, n2833, n2832, n2831, n2830, n2829, n2828, 
        n2827, n2826, n2825, n2824, n2823, n2822, n2821, n2820, n2819, n2818, 
        n2817, n2816, n2815, n2814}), .CI(1'b0), .DIFF({N1219, N1218, N1217, 
        N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, 
        N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, 
        N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188}) );
  poly5_DW01_sub_60 sub_45_S2_C84 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N1299, N1298, N1297, N1296, 
        N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, 
        N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, 
        N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, 
        N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, 
        N1255, N1254, N1253, N1252}), .CI(1'b0), .DIFF({N1333, N1332, N1331, 
        N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, 
        N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, 
        N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223}) );
  poly5_DW01_add_19 add_0_root_add_0_root_add_89_5 ( .A({N2273, N2272, N2271, 
        N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, 
        N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, 
        N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242}), .B({
        n2813, n2812, n2811, n2810, n2809, n2808, n2807, n2806, n2805, n2804, 
        n2803, n2802, n2801, n2800, n2799, n2798, n2797, n2796, n2795, n2794, 
        n2793, n2792, n2791, n2790, n2789, n2788, n2787, n2786, n2785, n2784, 
        n2783, n2782}), .CI(1'b0), .SUM(res) );
  poly5_DW_mult_uns_44 mult_43_C85 ( .a({N1398, N1397, N1396, N1395, N1394, 
        N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, 
        N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, 
        N1373, N1372, N1371, N1370, N1369, N1368, N1367}), .b({n2780, N974, 
        N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, 
        N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, 
        n1893, N949, n1854, N947, n1851, N945, N944}), .product({
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, N1510, N1509, 
        N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, 
        N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, 
        N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, 
        N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, 
        N1468, N1467, N1466, N1465, N1464, N1463}) );
  poly5_DW_mult_uns_49 mult_43_C80 ( .a({n1845, n1830, n2004, n1890, n2006, 
        n1892, n2008, N821, n2010, N819, n2012, N817, n2014, n1852, n2016, 
        N813, n2018, n1891, n1853, N809, n2020, n1855, n2022, N805, n2024, 
        N803, n2026, N801, N800, N799, n2028, n2030}), .b({n1845, n1830, n2004, 
        n1890, n2006, N823, n2008, N821, n2010, N819, n2012, N817, N816, N815, 
        n2016, N813, N812, N811, N810, N809, n2020, N807, n2022, N805, n2024, 
        N803, n2026, N801, N800, N799, n2028, n2030}), .product({
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, t1, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271}) );
  poly5_DW01_sub_78 r374 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n2031, t1[30:24], n1881, t1[22:20], n1888, t1[18:0]}), .CI(1'b0), 
        .DIFF({N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, 
        N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, 
        N499, N498, N497, N496, N495, N494, N493, N492, N491, N490}) );
  poly5_DW_mult_uns_57 mult_43_C81 ( .a({n1833, n3032, n3031, n1835, n3029, 
        n3028, n3027, n3026, n3025, n3024, n3023, n3022, n3021, n3020, n3019, 
        n3018, n3017, n3016, n3015, n3014, n3013, n3012, n3011, n3010, n3009, 
        n3008, n3007, n3006, n3005, n3004, n1921, n3003}), .b({n1845, n1830, 
        n2004, n1890, n2006, n1892, n2008, N821, n2010, N819, n2012, N817, 
        n2014, n1852, n2016, N813, n2018, n1891, n1853, N809, n2020, n1855, 
        n2022, N805, n2024, N803, n2026, N801, N800, N799, n2028, n2030}), 
        .product({SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, N665, N664, N663, 
        N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, 
        N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, 
        N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, 
        N626, N625, N624, N623, N622, N621, N620, N619, N618}) );
  BUFX4 U1941 ( .A(t1[19]), .Y(n1888) );
  INVX8 U1942 ( .A(n2027), .Y(n2026) );
  INVX4 U1943 ( .A(N802), .Y(n2027) );
  INVX4 U1944 ( .A(N827), .Y(n1829) );
  INVX8 U1945 ( .A(n1829), .Y(n1830) );
  INVX2 U1946 ( .A(n2077), .Y(N827) );
  BUFX4 U1947 ( .A(n2204), .Y(n1831) );
  INVX4 U1948 ( .A(n1880), .Y(n1832) );
  INVX8 U1949 ( .A(n1832), .Y(n1833) );
  INVX2 U1950 ( .A(n1862), .Y(n1880) );
  INVX4 U1951 ( .A(n2547), .Y(n1893) );
  INVX4 U1952 ( .A(n3030), .Y(n1834) );
  INVX8 U1953 ( .A(n1834), .Y(n1835) );
  INVX2 U1954 ( .A(n2206), .Y(n3030) );
  BUFX4 U1955 ( .A(N648), .Y(n1836) );
  INVX4 U1956 ( .A(n2104), .Y(N800) );
  INVX2 U1957 ( .A(n2337), .Y(n2965) );
  INVX2 U1958 ( .A(n2088), .Y(N816) );
  INVX2 U1959 ( .A(n2101), .Y(N803) );
  INVX2 U1960 ( .A(n2103), .Y(N801) );
  INVX2 U1961 ( .A(n2099), .Y(N805) );
  INVX2 U1962 ( .A(n2544), .Y(N953) );
  INVX2 U1963 ( .A(n2548), .Y(N949) );
  INVX2 U1964 ( .A(n2552), .Y(N945) );
  INVX2 U1965 ( .A(n2357), .Y(n2945) );
  INVX2 U1966 ( .A(N798), .Y(n2029) );
  INVX4 U1967 ( .A(n2025), .Y(n2024) );
  INVX2 U1968 ( .A(N804), .Y(n2025) );
  INVX4 U1969 ( .A(n2023), .Y(n2022) );
  INVX2 U1970 ( .A(N806), .Y(n2023) );
  INVX2 U1971 ( .A(n2541), .Y(N956) );
  INVX2 U1972 ( .A(n2513), .Y(n2885) );
  BUFX2 U1973 ( .A(N636), .Y(n1865) );
  INVX4 U1974 ( .A(n2233), .Y(n1921) );
  INVX2 U1975 ( .A(n2228), .Y(n3008) );
  INVX2 U1976 ( .A(n2227), .Y(n3009) );
  INVX2 U1977 ( .A(n2231), .Y(n3005) );
  INVX2 U1978 ( .A(N808), .Y(n2021) );
  INVX2 U1979 ( .A(n2385), .Y(N742) );
  INVX2 U1980 ( .A(n2225), .Y(n3011) );
  INVX2 U1981 ( .A(n2224), .Y(n3012) );
  BUFX2 U1982 ( .A(N652), .Y(n1864) );
  BUFX2 U1983 ( .A(N862), .Y(n1840) );
  INVX2 U1984 ( .A(n2539), .Y(N958) );
  INVX2 U1985 ( .A(n2538), .Y(N959) );
  INVX2 U1986 ( .A(n2358), .Y(n2944) );
  INVX2 U1987 ( .A(n2354), .Y(n2948) );
  INVX2 U1988 ( .A(n2223), .Y(n3013) );
  INVX2 U1989 ( .A(n2222), .Y(n3014) );
  INVX2 U1990 ( .A(n2352), .Y(n2950) );
  INVX4 U1991 ( .A(n2013), .Y(n2012) );
  INVX2 U1992 ( .A(N818), .Y(n2013) );
  INVX4 U1993 ( .A(n2009), .Y(n2008) );
  INVX2 U1994 ( .A(N822), .Y(n2009) );
  INVX2 U1995 ( .A(n2530), .Y(N967) );
  INVX2 U1996 ( .A(n2532), .Y(N965) );
  INVX2 U1997 ( .A(n2334), .Y(n2968) );
  INVX2 U1998 ( .A(N820), .Y(n2011) );
  INVX2 U1999 ( .A(N814), .Y(n2017) );
  INVX2 U2000 ( .A(n2007), .Y(n2006) );
  INVX2 U2001 ( .A(N824), .Y(n2007) );
  INVX2 U2002 ( .A(n2347), .Y(n2955) );
  INVX2 U2003 ( .A(n2367), .Y(N760) );
  INVX2 U2004 ( .A(n2534), .Y(N963) );
  INVX2 U2005 ( .A(n2527), .Y(N970) );
  INVX2 U2006 ( .A(n2522), .Y(n2780) );
  INVX2 U2007 ( .A(n2369), .Y(N758) );
  INVX2 U2008 ( .A(n2365), .Y(N762) );
  INVX2 U2009 ( .A(n2364), .Y(N763) );
  INVX2 U2010 ( .A(N816), .Y(n2015) );
  BUFX2 U2011 ( .A(N1084), .Y(n1883) );
  BUFX2 U2012 ( .A(x[2]), .Y(n1884) );
  BUFX2 U2013 ( .A(x[3]), .Y(n1841) );
  BUFX2 U2014 ( .A(x[8]), .Y(n1843) );
  BUFX2 U2015 ( .A(x[16]), .Y(n1842) );
  BUFX4 U2016 ( .A(N643), .Y(n1837) );
  INVX2 U2017 ( .A(n2551), .Y(n1851) );
  INVX2 U2018 ( .A(n2208), .Y(n1838) );
  INVX4 U2019 ( .A(n1838), .Y(n1839) );
  INVX1 U2020 ( .A(x[6]), .Y(n2052) );
  INVX1 U2021 ( .A(x[1]), .Y(n2047) );
  BUFX4 U2022 ( .A(N1073), .Y(n1844) );
  INVX2 U2023 ( .A(n1878), .Y(n1872) );
  INVX1 U2024 ( .A(n1856), .Y(n1904) );
  INVX2 U2025 ( .A(n2490), .Y(n1876) );
  INVX2 U2026 ( .A(n1926), .Y(n1925) );
  AND2X2 U2027 ( .A(N310), .B(n2035), .Y(n1845) );
  INVX2 U2028 ( .A(n2490), .Y(n1877) );
  INVX2 U2029 ( .A(n2545), .Y(N952) );
  XOR2X1 U2030 ( .A(n3067), .B(n2036), .Y(n1846) );
  INVX4 U2031 ( .A(n2029), .Y(n2028) );
  INVX2 U2032 ( .A(n2393), .Y(N734) );
  INVX2 U2033 ( .A(n1863), .Y(n1916) );
  INVX2 U2034 ( .A(n2107), .Y(n2030) );
  BUFX2 U2035 ( .A(n1848), .Y(n1847) );
  BUFX2 U2036 ( .A(pushdata), .Y(n1848) );
  BUFX4 U2037 ( .A(n1219), .Y(n1850) );
  BUFX2 U2038 ( .A(rst), .Y(n1849) );
  MUX2X1 U2039 ( .B(N924), .A(n2889), .S(n1900), .Y(n2541) );
  INVX1 U2040 ( .A(n1898), .Y(n1902) );
  MUX2X1 U2041 ( .B(n2881), .A(N916), .S(n1856), .Y(n2549) );
  BUFX4 U2042 ( .A(n3066), .Y(n1856) );
  INVX1 U2043 ( .A(N1290), .Y(n2735) );
  INVX1 U2044 ( .A(n2551), .Y(N946) );
  MUX2X1 U2045 ( .B(N289), .A(x[10]), .S(n2036), .Y(n2097) );
  MUX2X1 U2046 ( .B(N286), .A(x[7]), .S(n2036), .Y(n2100) );
  MUX2X1 U2047 ( .B(N285), .A(x[6]), .S(n2036), .Y(n2101) );
  BUFX2 U2048 ( .A(N815), .Y(n1852) );
  INVX2 U2049 ( .A(n2089), .Y(N815) );
  INVX2 U2050 ( .A(n2092), .Y(N812) );
  INVX1 U2051 ( .A(N812), .Y(n2019) );
  INVX2 U2052 ( .A(n2015), .Y(n2014) );
  MUX2X1 U2053 ( .B(N296), .A(x[17]), .S(n2036), .Y(n2090) );
  MUX2X1 U2054 ( .B(N298), .A(x[19]), .S(n2036), .Y(n2088) );
  BUFX2 U2055 ( .A(N810), .Y(n1853) );
  INVX2 U2056 ( .A(n2094), .Y(N810) );
  MUX2X1 U2057 ( .B(N299), .A(x[20]), .S(n2036), .Y(n2087) );
  INVX1 U2058 ( .A(n1904), .Y(n1908) );
  MUX2X1 U2059 ( .B(N291), .A(x[12]), .S(n2036), .Y(n2095) );
  MUX2X1 U2060 ( .B(N301), .A(x[22]), .S(n2036), .Y(n2085) );
  INVX4 U2061 ( .A(n2549), .Y(n1854) );
  MUX2X1 U2062 ( .B(N288), .A(x[9]), .S(n2036), .Y(n2098) );
  INVX2 U2063 ( .A(n2019), .Y(n2018) );
  BUFX2 U2064 ( .A(N647), .Y(n1882) );
  INVX1 U2065 ( .A(n1856), .Y(n1905) );
  INVX4 U2066 ( .A(n2526), .Y(N971) );
  INVX2 U2067 ( .A(n2543), .Y(N954) );
  INVX1 U2068 ( .A(N1319), .Y(n2744) );
  BUFX2 U2069 ( .A(N807), .Y(n1855) );
  INVX2 U2070 ( .A(n2097), .Y(N807) );
  INVX4 U2071 ( .A(n3066), .Y(n1926) );
  INVX4 U2072 ( .A(n2209), .Y(n3027) );
  INVX2 U2073 ( .A(n1877), .Y(n1857) );
  INVX1 U2074 ( .A(n1925), .Y(n1858) );
  INVX2 U2075 ( .A(n2046), .Y(n1859) );
  INVX1 U2076 ( .A(n3027), .Y(n1860) );
  INVX2 U2077 ( .A(n1860), .Y(n1861) );
  INVX4 U2078 ( .A(t1[31]), .Y(n2033) );
  INVX4 U2079 ( .A(n2036), .Y(n2034) );
  NAND2X1 U2080 ( .A(n2032), .B(N521), .Y(n1862) );
  INVX2 U2081 ( .A(n1924), .Y(n1923) );
  INVX1 U2082 ( .A(N1188), .Y(n2712) );
  INVX4 U2083 ( .A(n2205), .Y(n3031) );
  MUX2X1 U2084 ( .B(N717), .A(n2956), .S(n1857), .Y(n2378) );
  MUX2X1 U2085 ( .B(N730), .A(n2969), .S(n1857), .Y(n2365) );
  INVX2 U2086 ( .A(n2371), .Y(N756) );
  MUX2X1 U2087 ( .B(N939), .A(n2904), .S(n1899), .Y(n2526) );
  MUX2X1 U2088 ( .B(N929), .A(n2894), .S(n1906), .Y(n2536) );
  INVX2 U2089 ( .A(n2348), .Y(n2954) );
  MUX2X1 U2090 ( .B(N930), .A(n2895), .S(n1858), .Y(n2535) );
  MUX2X1 U2091 ( .B(N936), .A(n2901), .S(n1858), .Y(n2529) );
  MUX2X1 U2092 ( .B(N928), .A(n2893), .S(n1903), .Y(n2537) );
  MUX2X1 U2093 ( .B(N933), .A(n2898), .S(n1907), .Y(n2532) );
  MUX2X1 U2094 ( .B(N935), .A(n2900), .S(n1858), .Y(n2530) );
  INVX2 U2095 ( .A(n2528), .Y(N969) );
  INVX2 U2096 ( .A(n2540), .Y(N957) );
  INVX2 U2097 ( .A(n2687), .Y(n2827) );
  INVX2 U2098 ( .A(n2351), .Y(n2951) );
  MUX2X1 U2099 ( .B(N922), .A(n2887), .S(n1898), .Y(n2543) );
  MUX2X1 U2100 ( .B(n2891), .A(N926), .S(n1856), .Y(n2539) );
  INVX2 U2101 ( .A(n2512), .Y(n2886) );
  INVX2 U2102 ( .A(n2331), .Y(n1914) );
  INVX2 U2103 ( .A(n2235), .Y(n1913) );
  INVX2 U2104 ( .A(n1962), .Y(n1959) );
  INVX2 U2105 ( .A(n1976), .Y(n1973) );
  INVX2 U2106 ( .A(n1984), .Y(n1981) );
  INVX2 U2107 ( .A(n1992), .Y(n1989) );
  INVX2 U2108 ( .A(n1958), .Y(n1957) );
  INVX2 U2109 ( .A(n2554), .Y(n1918) );
  INVX2 U2110 ( .A(n1846), .Y(n1917) );
  INVX2 U2111 ( .A(n2651), .Y(n1919) );
  INVX2 U2112 ( .A(n2715), .Y(n1920) );
  INVX2 U2113 ( .A(n1916), .Y(n1915) );
  INVX2 U2114 ( .A(n2045), .Y(n1911) );
  INVX2 U2115 ( .A(n2108), .Y(n1912) );
  BUFX2 U2116 ( .A(n513), .Y(n1962) );
  BUFX2 U2117 ( .A(n513), .Y(n1961) );
  BUFX2 U2118 ( .A(n513), .Y(n1960) );
  BUFX2 U2119 ( .A(n1980), .Y(n1976) );
  BUFX2 U2120 ( .A(n1980), .Y(n1975) );
  BUFX2 U2121 ( .A(n1980), .Y(n1974) );
  BUFX2 U2122 ( .A(n1988), .Y(n1984) );
  BUFX2 U2123 ( .A(n1988), .Y(n1983) );
  BUFX2 U2124 ( .A(n1988), .Y(n1982) );
  BUFX2 U2125 ( .A(n1996), .Y(n1992) );
  BUFX2 U2126 ( .A(n1996), .Y(n1991) );
  BUFX2 U2127 ( .A(n1996), .Y(n1990) );
  BUFX2 U2128 ( .A(n513), .Y(n1964) );
  BUFX2 U2129 ( .A(n513), .Y(n1963) );
  BUFX2 U2130 ( .A(n1974), .Y(n1978) );
  BUFX2 U2131 ( .A(n1974), .Y(n1977) );
  BUFX2 U2132 ( .A(n1982), .Y(n1986) );
  BUFX2 U2133 ( .A(n1982), .Y(n1985) );
  BUFX2 U2134 ( .A(n1990), .Y(n1994) );
  BUFX2 U2135 ( .A(n1990), .Y(n1993) );
  INVX2 U2136 ( .A(n1969), .Y(n1966) );
  INVX2 U2137 ( .A(n2000), .Y(n1997) );
  INVX2 U2138 ( .A(n644), .Y(n1958) );
  BUFX2 U2139 ( .A(n513), .Y(n1965) );
  BUFX2 U2140 ( .A(n1974), .Y(n1979) );
  BUFX2 U2141 ( .A(n1982), .Y(n1987) );
  BUFX2 U2142 ( .A(n1990), .Y(n1995) );
  BUFX2 U2143 ( .A(n1933), .Y(n1955) );
  BUFX2 U2144 ( .A(n1930), .Y(n1946) );
  BUFX2 U2145 ( .A(n1931), .Y(n1947) );
  BUFX2 U2146 ( .A(n1931), .Y(n1948) );
  BUFX2 U2147 ( .A(n1931), .Y(n1949) );
  BUFX2 U2148 ( .A(n1932), .Y(n1950) );
  BUFX2 U2149 ( .A(n1932), .Y(n1951) );
  BUFX2 U2150 ( .A(n1932), .Y(n1952) );
  BUFX2 U2151 ( .A(n1933), .Y(n1953) );
  BUFX2 U2152 ( .A(n1933), .Y(n1954) );
  BUFX2 U2153 ( .A(n1927), .Y(n1935) );
  BUFX2 U2154 ( .A(n1927), .Y(n1936) );
  BUFX2 U2155 ( .A(n1927), .Y(n1937) );
  BUFX2 U2156 ( .A(n1928), .Y(n1938) );
  BUFX2 U2157 ( .A(n1928), .Y(n1939) );
  BUFX2 U2158 ( .A(n1928), .Y(n1940) );
  BUFX2 U2159 ( .A(n1929), .Y(n1941) );
  BUFX2 U2160 ( .A(n1929), .Y(n1942) );
  BUFX2 U2161 ( .A(n1929), .Y(n1943) );
  BUFX2 U2162 ( .A(n1930), .Y(n1944) );
  BUFX2 U2163 ( .A(n1930), .Y(n1945) );
  INVX2 U2164 ( .A(n2036), .Y(n2035) );
  XNOR2X1 U2165 ( .A(n3067), .B(n2042), .Y(n1863) );
  INVX2 U2166 ( .A(n2044), .Y(n2043) );
  INVX2 U2167 ( .A(n2042), .Y(n2041) );
  INVX2 U2168 ( .A(n2040), .Y(n2039) );
  INVX2 U2169 ( .A(n2038), .Y(n2037) );
  BUFX2 U2170 ( .A(n229), .Y(n1998) );
  BUFX2 U2171 ( .A(n229), .Y(n2000) );
  BUFX2 U2172 ( .A(n229), .Y(n1999) );
  BUFX2 U2173 ( .A(n511), .Y(n1969) );
  BUFX2 U2174 ( .A(n511), .Y(n1968) );
  BUFX2 U2175 ( .A(n511), .Y(n1967) );
  BUFX2 U2176 ( .A(n229), .Y(n2002) );
  BUFX2 U2177 ( .A(n229), .Y(n2001) );
  BUFX2 U2178 ( .A(n511), .Y(n1971) );
  BUFX2 U2179 ( .A(n511), .Y(n1970) );
  INVX2 U2180 ( .A(n510), .Y(n1980) );
  BUFX2 U2181 ( .A(n229), .Y(n2003) );
  INVX2 U2182 ( .A(n307), .Y(n1988) );
  INVX2 U2183 ( .A(n268), .Y(n1996) );
  BUFX2 U2184 ( .A(n511), .Y(n1972) );
  BUFX2 U2185 ( .A(n1934), .Y(n1956) );
  BUFX2 U2186 ( .A(n3068), .Y(n1934) );
  BUFX2 U2187 ( .A(n3068), .Y(n1931) );
  BUFX2 U2188 ( .A(n3068), .Y(n1932) );
  BUFX2 U2189 ( .A(n3068), .Y(n1933) );
  BUFX2 U2190 ( .A(n3068), .Y(n1927) );
  BUFX2 U2191 ( .A(n3068), .Y(n1928) );
  BUFX2 U2192 ( .A(n3068), .Y(n1929) );
  BUFX2 U2193 ( .A(n3068), .Y(n1930) );
  INVX4 U2194 ( .A(x[31]), .Y(n2036) );
  INVX2 U2195 ( .A(n2081), .Y(N823) );
  INVX4 U2196 ( .A(N826), .Y(n2005) );
  INVX2 U2197 ( .A(a1[31]), .Y(n2045) );
  INVX2 U2198 ( .A(a3[31]), .Y(n2042) );
  INVX2 U2199 ( .A(a2[31]), .Y(n2044) );
  INVX2 U2200 ( .A(a4[31]), .Y(n2040) );
  INVX2 U2201 ( .A(a5[31]), .Y(n2038) );
  INVX4 U2202 ( .A(n2524), .Y(N973) );
  INVX1 U2203 ( .A(x[13]), .Y(n2059) );
  INVX4 U2204 ( .A(n2218), .Y(n3018) );
  INVX1 U2205 ( .A(n1879), .Y(n1866) );
  INVX1 U2206 ( .A(n1879), .Y(n1867) );
  INVX1 U2207 ( .A(n1879), .Y(n1868) );
  INVX1 U2208 ( .A(n1879), .Y(n1869) );
  INVX1 U2209 ( .A(n1879), .Y(n1870) );
  INVX1 U2210 ( .A(n1879), .Y(n1871) );
  INVX1 U2211 ( .A(n1878), .Y(n1873) );
  INVX1 U2212 ( .A(n1878), .Y(n1874) );
  INVX1 U2213 ( .A(n1878), .Y(n1875) );
  INVX1 U2214 ( .A(n1857), .Y(n3067) );
  MUX2X1 U2215 ( .B(N665), .A(N699), .S(n1914), .Y(n1878) );
  MUX2X1 U2216 ( .B(N665), .A(N699), .S(n1914), .Y(n1879) );
  BUFX4 U2217 ( .A(t1[23]), .Y(n1881) );
  BUFX4 U2218 ( .A(x[5]), .Y(n1885) );
  BUFX4 U2219 ( .A(x[4]), .Y(n1886) );
  BUFX4 U2220 ( .A(N651), .Y(n1887) );
  INVX4 U2221 ( .A(n2083), .Y(N821) );
  INVX4 U2222 ( .A(n2085), .Y(N819) );
  INVX4 U2223 ( .A(n2091), .Y(N813) );
  INVX4 U2224 ( .A(n2087), .Y(N817) );
  INVX4 U2225 ( .A(N825), .Y(n1889) );
  INVX8 U2226 ( .A(n1889), .Y(n1890) );
  INVX4 U2227 ( .A(n2095), .Y(N809) );
  BUFX2 U2228 ( .A(N811), .Y(n1891) );
  BUFX2 U2229 ( .A(N823), .Y(n1892) );
  INVX1 U2230 ( .A(n1856), .Y(n1903) );
  INVX2 U2231 ( .A(n1907), .Y(n1910) );
  INVX2 U2232 ( .A(n3066), .Y(n1898) );
  MUX2X1 U2233 ( .B(N920), .A(n2885), .S(n1899), .Y(n2545) );
  INVX2 U2234 ( .A(n2542), .Y(n1894) );
  INVX2 U2235 ( .A(n2542), .Y(N955) );
  MUX2X1 U2236 ( .B(N918), .A(n2883), .S(n1926), .Y(n2547) );
  MUX2X1 U2237 ( .B(N921), .A(n2886), .S(n1898), .Y(n2544) );
  MUX2X1 U2238 ( .B(N912), .A(n2877), .S(n1926), .Y(n2553) );
  INVX1 U2239 ( .A(n1858), .Y(n1895) );
  INVX1 U2240 ( .A(N1214), .Y(n2660) );
  INVX4 U2241 ( .A(n2216), .Y(n3020) );
  MUX2X1 U2242 ( .B(N515), .A(t1[25]), .S(n2033), .Y(n2209) );
  INVX4 U2243 ( .A(n2207), .Y(n3029) );
  INVX1 U2244 ( .A(x[11]), .Y(n2057) );
  INVX1 U2245 ( .A(x[10]), .Y(n2056) );
  INVX2 U2246 ( .A(x[0]), .Y(n1896) );
  INVX4 U2247 ( .A(n1896), .Y(n1897) );
  INVX1 U2248 ( .A(x[12]), .Y(n2058) );
  INVX1 U2249 ( .A(x[17]), .Y(n2063) );
  INVX4 U2250 ( .A(n2363), .Y(n2781) );
  INVX4 U2251 ( .A(n2349), .Y(n2953) );
  INVX4 U2252 ( .A(n2550), .Y(N947) );
  INVX4 U2253 ( .A(n2508), .Y(n2890) );
  INVX1 U2254 ( .A(n3066), .Y(n1899) );
  INVX1 U2255 ( .A(n1925), .Y(n1900) );
  INVX2 U2256 ( .A(n1899), .Y(n1901) );
  INVX1 U2257 ( .A(n1856), .Y(n1906) );
  INVX1 U2258 ( .A(n1856), .Y(n1907) );
  INVX2 U2259 ( .A(n1905), .Y(n1909) );
  INVX1 U2260 ( .A(N1320), .Y(n2742) );
  INVX4 U2261 ( .A(n2234), .Y(n3003) );
  INVX4 U2262 ( .A(n2379), .Y(N748) );
  INVX4 U2263 ( .A(n2546), .Y(N951) );
  INVX1 U2264 ( .A(N1279), .Y(n2757) );
  INVX8 U2265 ( .A(n1831), .Y(n3032) );
  INVX1 U2266 ( .A(x[9]), .Y(n2055) );
  INVX4 U2267 ( .A(n2383), .Y(N744) );
  INVX1 U2268 ( .A(N1543), .Y(n2557) );
  INVX1 U2269 ( .A(n1886), .Y(n2050) );
  INVX1 U2270 ( .A(N1289), .Y(n2737) );
  INVX8 U2271 ( .A(n1839), .Y(n3028) );
  INVX1 U2272 ( .A(n1842), .Y(n2062) );
  INVX4 U2273 ( .A(n3065), .Y(n1924) );
  INVX1 U2274 ( .A(n1843), .Y(n2054) );
  INVX1 U2275 ( .A(N1285), .Y(n2745) );
  INVX1 U2276 ( .A(N1293), .Y(n2729) );
  INVX4 U2277 ( .A(n2650), .Y(n3066) );
  INVX1 U2278 ( .A(n1897), .Y(n2046) );
  INVX1 U2279 ( .A(N1283), .Y(n2749) );
  INVX8 U2280 ( .A(n1924), .Y(n1922) );
  INVX8 U2281 ( .A(n2005), .Y(n2004) );
  INVX8 U2282 ( .A(n2011), .Y(n2010) );
  INVX8 U2283 ( .A(n2017), .Y(n2016) );
  INVX8 U2284 ( .A(n2021), .Y(n2020) );
  INVX8 U2285 ( .A(n2033), .Y(n2031) );
  INVX8 U2286 ( .A(n2033), .Y(n2032) );
  INVX2 U2287 ( .A(a4[30]), .Y(n3104) );
  INVX2 U2288 ( .A(a4[29]), .Y(n3105) );
  INVX2 U2289 ( .A(a4[28]), .Y(n3106) );
  INVX2 U2290 ( .A(a4[27]), .Y(n3107) );
  INVX2 U2291 ( .A(a4[26]), .Y(n3108) );
  INVX2 U2292 ( .A(a4[25]), .Y(n3109) );
  INVX2 U2293 ( .A(a4[24]), .Y(n3110) );
  INVX2 U2294 ( .A(a4[23]), .Y(n3111) );
  INVX2 U2295 ( .A(a4[22]), .Y(n3112) );
  INVX2 U2296 ( .A(a4[21]), .Y(n3113) );
  INVX2 U2297 ( .A(a4[20]), .Y(n3114) );
  INVX2 U2298 ( .A(a4[19]), .Y(n3115) );
  INVX2 U2299 ( .A(a4[18]), .Y(n3116) );
  INVX2 U2300 ( .A(a4[17]), .Y(n3117) );
  INVX2 U2301 ( .A(a4[16]), .Y(n3118) );
  INVX2 U2302 ( .A(a4[15]), .Y(n3119) );
  INVX2 U2303 ( .A(a4[14]), .Y(n3120) );
  INVX2 U2304 ( .A(a4[13]), .Y(n3121) );
  INVX2 U2305 ( .A(a4[12]), .Y(n3122) );
  INVX2 U2306 ( .A(a4[11]), .Y(n3123) );
  INVX2 U2307 ( .A(a4[10]), .Y(n3124) );
  INVX2 U2308 ( .A(a4[9]), .Y(n3125) );
  INVX2 U2309 ( .A(a4[8]), .Y(n3126) );
  INVX2 U2310 ( .A(a4[7]), .Y(n3127) );
  INVX2 U2311 ( .A(a4[6]), .Y(n3128) );
  INVX2 U2312 ( .A(a4[5]), .Y(n3129) );
  INVX2 U2313 ( .A(a4[4]), .Y(n3130) );
  INVX2 U2314 ( .A(a4[3]), .Y(n3131) );
  INVX2 U2315 ( .A(a4[2]), .Y(n3132) );
  INVX2 U2316 ( .A(a4[1]), .Y(n3133) );
  INVX2 U2317 ( .A(a4[0]), .Y(n3134) );
  INVX2 U2318 ( .A(a5[30]), .Y(n3135) );
  INVX2 U2319 ( .A(a5[29]), .Y(n3136) );
  INVX2 U2320 ( .A(a5[28]), .Y(n3137) );
  INVX2 U2321 ( .A(a5[27]), .Y(n3138) );
  INVX2 U2322 ( .A(a5[26]), .Y(n3139) );
  INVX2 U2323 ( .A(a5[25]), .Y(n3140) );
  INVX2 U2324 ( .A(a5[24]), .Y(n3141) );
  INVX2 U2325 ( .A(a5[23]), .Y(n3142) );
  INVX2 U2326 ( .A(a5[22]), .Y(n3143) );
  INVX2 U2327 ( .A(a5[21]), .Y(n3144) );
  INVX2 U2328 ( .A(a5[20]), .Y(n3145) );
  INVX2 U2329 ( .A(a5[19]), .Y(n3146) );
  INVX2 U2330 ( .A(a5[18]), .Y(n3147) );
  INVX2 U2331 ( .A(a5[17]), .Y(n3148) );
  INVX2 U2332 ( .A(a5[16]), .Y(n3149) );
  INVX2 U2333 ( .A(a5[15]), .Y(n3150) );
  INVX2 U2334 ( .A(a5[14]), .Y(n3151) );
  INVX2 U2335 ( .A(a5[13]), .Y(n3152) );
  INVX2 U2336 ( .A(a5[12]), .Y(n3153) );
  INVX2 U2337 ( .A(a5[11]), .Y(n3154) );
  INVX2 U2338 ( .A(a5[10]), .Y(n3155) );
  INVX2 U2339 ( .A(a5[9]), .Y(n3156) );
  INVX2 U2340 ( .A(a5[8]), .Y(n3157) );
  INVX2 U2341 ( .A(a5[7]), .Y(n3158) );
  INVX2 U2342 ( .A(a5[6]), .Y(n3159) );
  INVX2 U2343 ( .A(a5[5]), .Y(n3160) );
  INVX2 U2344 ( .A(a5[4]), .Y(n3161) );
  INVX2 U2345 ( .A(a5[3]), .Y(n3162) );
  INVX2 U2346 ( .A(a5[2]), .Y(n3163) );
  INVX2 U2347 ( .A(a5[1]), .Y(n3164) );
  INVX2 U2348 ( .A(a5[0]), .Y(n3165) );
  INVX2 U2349 ( .A(a2[30]), .Y(n3197) );
  INVX2 U2350 ( .A(a2[29]), .Y(n3198) );
  INVX2 U2351 ( .A(a2[28]), .Y(n3199) );
  INVX2 U2352 ( .A(a2[27]), .Y(n3200) );
  INVX2 U2353 ( .A(a2[26]), .Y(n3201) );
  INVX2 U2354 ( .A(a2[25]), .Y(n3202) );
  INVX2 U2355 ( .A(a2[24]), .Y(n3203) );
  INVX2 U2356 ( .A(a2[23]), .Y(n3204) );
  INVX2 U2357 ( .A(a2[22]), .Y(n3205) );
  INVX2 U2358 ( .A(a2[21]), .Y(n3206) );
  INVX2 U2359 ( .A(a2[20]), .Y(n3207) );
  INVX2 U2360 ( .A(a2[19]), .Y(n3208) );
  INVX2 U2361 ( .A(a2[18]), .Y(n3209) );
  INVX2 U2362 ( .A(a2[17]), .Y(n3210) );
  INVX2 U2363 ( .A(a2[16]), .Y(n3211) );
  INVX2 U2364 ( .A(a2[15]), .Y(n3212) );
  INVX2 U2365 ( .A(a2[14]), .Y(n3213) );
  INVX2 U2366 ( .A(a2[13]), .Y(n3214) );
  INVX2 U2367 ( .A(a2[12]), .Y(n3215) );
  INVX2 U2368 ( .A(a2[11]), .Y(n3216) );
  INVX2 U2369 ( .A(a2[10]), .Y(n3217) );
  INVX2 U2370 ( .A(a2[9]), .Y(n3218) );
  INVX2 U2371 ( .A(a2[8]), .Y(n3219) );
  INVX2 U2372 ( .A(a2[7]), .Y(n3220) );
  INVX2 U2373 ( .A(a2[6]), .Y(n3221) );
  INVX2 U2374 ( .A(a2[5]), .Y(n3222) );
  INVX2 U2375 ( .A(a2[4]), .Y(n3223) );
  INVX2 U2376 ( .A(a2[3]), .Y(n3224) );
  INVX2 U2377 ( .A(a2[2]), .Y(n3225) );
  INVX2 U2378 ( .A(a2[1]), .Y(n3226) );
  INVX2 U2379 ( .A(a2[0]), .Y(n3227) );
  INVX2 U2380 ( .A(a3[30]), .Y(n3228) );
  INVX2 U2381 ( .A(a3[29]), .Y(n3229) );
  INVX2 U2382 ( .A(a3[28]), .Y(n3230) );
  INVX2 U2383 ( .A(a3[27]), .Y(n3231) );
  INVX2 U2384 ( .A(a3[26]), .Y(n3232) );
  INVX2 U2385 ( .A(a3[25]), .Y(n3233) );
  INVX2 U2386 ( .A(a3[24]), .Y(n3234) );
  INVX2 U2387 ( .A(a3[23]), .Y(n3235) );
  INVX2 U2388 ( .A(a3[22]), .Y(n3236) );
  INVX2 U2389 ( .A(a3[21]), .Y(n3237) );
  INVX2 U2390 ( .A(a3[20]), .Y(n3238) );
  INVX2 U2391 ( .A(a3[19]), .Y(n3239) );
  INVX2 U2392 ( .A(a3[18]), .Y(n3240) );
  INVX2 U2393 ( .A(a3[17]), .Y(n3241) );
  INVX2 U2394 ( .A(a3[16]), .Y(n3242) );
  INVX2 U2395 ( .A(a3[15]), .Y(n3243) );
  INVX2 U2396 ( .A(a3[14]), .Y(n3244) );
  INVX2 U2397 ( .A(a3[13]), .Y(n3245) );
  INVX2 U2398 ( .A(a3[12]), .Y(n3246) );
  INVX2 U2399 ( .A(a3[11]), .Y(n3247) );
  INVX2 U2400 ( .A(a3[10]), .Y(n3248) );
  INVX2 U2401 ( .A(a3[9]), .Y(n3249) );
  INVX2 U2402 ( .A(a3[8]), .Y(n3250) );
  INVX2 U2403 ( .A(a3[7]), .Y(n3251) );
  INVX2 U2404 ( .A(a3[6]), .Y(n3252) );
  INVX2 U2405 ( .A(a3[5]), .Y(n3253) );
  INVX2 U2406 ( .A(a3[4]), .Y(n3254) );
  INVX2 U2407 ( .A(a3[3]), .Y(n3255) );
  INVX2 U2408 ( .A(a3[2]), .Y(n3256) );
  INVX2 U2409 ( .A(a3[1]), .Y(n3257) );
  INVX2 U2410 ( .A(a3[0]), .Y(n3258) );
  OAI22X1 U2411 ( .A(n1998), .B(n3103), .C(n1997), .D(n2046), .Y(n1735) );
  OAI22X1 U2412 ( .A(n2003), .B(n3102), .C(n1997), .D(n2047), .Y(n1736) );
  INVX2 U2413 ( .A(n1884), .Y(n2048) );
  OAI22X1 U2414 ( .A(n2003), .B(n3101), .C(n1997), .D(n2048), .Y(n1737) );
  INVX2 U2415 ( .A(n1841), .Y(n2049) );
  OAI22X1 U2416 ( .A(n2003), .B(n3100), .C(n1997), .D(n2049), .Y(n1738) );
  OAI22X1 U2417 ( .A(n2003), .B(n3099), .C(n1997), .D(n2050), .Y(n1739) );
  INVX2 U2418 ( .A(n1885), .Y(n2051) );
  OAI22X1 U2419 ( .A(n2003), .B(n3098), .C(n1997), .D(n2051), .Y(n1740) );
  OAI22X1 U2420 ( .A(n2002), .B(n3097), .C(n1997), .D(n2052), .Y(n1741) );
  INVX2 U2421 ( .A(x[7]), .Y(n2053) );
  OAI22X1 U2422 ( .A(n2002), .B(n3096), .C(n1997), .D(n2053), .Y(n1742) );
  OAI22X1 U2423 ( .A(n2002), .B(n3095), .C(n1997), .D(n2054), .Y(n1743) );
  OAI22X1 U2424 ( .A(n2002), .B(n3094), .C(n1997), .D(n2055), .Y(n1744) );
  OAI22X1 U2425 ( .A(n2002), .B(n3093), .C(n1997), .D(n2056), .Y(n1745) );
  OAI22X1 U2426 ( .A(n2002), .B(n3092), .C(n1997), .D(n2057), .Y(n1746) );
  OAI22X1 U2427 ( .A(n2002), .B(n3091), .C(n1997), .D(n2058), .Y(n1747) );
  OAI22X1 U2428 ( .A(n2002), .B(n3090), .C(n1997), .D(n2059), .Y(n1748) );
  INVX2 U2429 ( .A(x[14]), .Y(n2060) );
  OAI22X1 U2430 ( .A(n2001), .B(n3089), .C(n1997), .D(n2060), .Y(n1749) );
  INVX2 U2431 ( .A(x[15]), .Y(n2061) );
  OAI22X1 U2432 ( .A(n2001), .B(n3088), .C(n1997), .D(n2061), .Y(n1750) );
  OAI22X1 U2433 ( .A(n2001), .B(n3087), .C(n1997), .D(n2062), .Y(n1751) );
  OAI22X1 U2434 ( .A(n2001), .B(n3086), .C(n1997), .D(n2063), .Y(n1752) );
  INVX2 U2435 ( .A(x[18]), .Y(n2064) );
  OAI22X1 U2436 ( .A(n2001), .B(n3085), .C(n1997), .D(n2064), .Y(n1753) );
  INVX2 U2437 ( .A(x[19]), .Y(n2065) );
  OAI22X1 U2438 ( .A(n2001), .B(n3084), .C(n1997), .D(n2065), .Y(n1754) );
  INVX2 U2439 ( .A(x[20]), .Y(n2066) );
  OAI22X1 U2440 ( .A(n2001), .B(n3083), .C(n1997), .D(n2066), .Y(n1755) );
  INVX2 U2441 ( .A(x[21]), .Y(n2067) );
  OAI22X1 U2442 ( .A(n2000), .B(n3082), .C(n1997), .D(n2067), .Y(n1756) );
  INVX2 U2443 ( .A(x[22]), .Y(n2068) );
  OAI22X1 U2444 ( .A(n2000), .B(n3081), .C(n1997), .D(n2068), .Y(n1757) );
  INVX2 U2445 ( .A(x[23]), .Y(n2069) );
  OAI22X1 U2446 ( .A(n2000), .B(n3080), .C(n1997), .D(n2069), .Y(n1758) );
  INVX2 U2447 ( .A(x[24]), .Y(n2070) );
  OAI22X1 U2448 ( .A(n2001), .B(n3079), .C(n1997), .D(n2070), .Y(n1759) );
  INVX2 U2449 ( .A(x[25]), .Y(n2071) );
  OAI22X1 U2450 ( .A(n2000), .B(n3078), .C(n1997), .D(n2071), .Y(n1760) );
  INVX2 U2451 ( .A(x[26]), .Y(n2072) );
  OAI22X1 U2452 ( .A(n1999), .B(n3077), .C(n1997), .D(n2072), .Y(n1761) );
  INVX2 U2453 ( .A(x[27]), .Y(n2073) );
  OAI22X1 U2454 ( .A(n1999), .B(n3076), .C(n1997), .D(n2073), .Y(n1762) );
  INVX2 U2455 ( .A(x[28]), .Y(n2074) );
  OAI22X1 U2456 ( .A(n1999), .B(n3075), .C(n1997), .D(n2074), .Y(n1763) );
  INVX2 U2457 ( .A(x[29]), .Y(n2075) );
  OAI22X1 U2458 ( .A(n1999), .B(n3074), .C(n1997), .D(n2075), .Y(n1764) );
  INVX2 U2459 ( .A(x[30]), .Y(n2076) );
  OAI22X1 U2460 ( .A(n1998), .B(n3073), .C(n1997), .D(n2076), .Y(n1765) );
  OAI22X1 U2461 ( .A(n1998), .B(n3072), .C(n1997), .D(n2036), .Y(n1766) );
  MUX2X1 U2462 ( .B(x[30]), .A(N309), .S(n2035), .Y(n2077) );
  MUX2X1 U2463 ( .B(x[29]), .A(N308), .S(n2035), .Y(n2078) );
  INVX2 U2464 ( .A(n2078), .Y(N826) );
  MUX2X1 U2465 ( .B(x[28]), .A(N307), .S(n2035), .Y(n2079) );
  INVX2 U2466 ( .A(n2079), .Y(N825) );
  MUX2X1 U2467 ( .B(x[27]), .A(N306), .S(n2035), .Y(n2080) );
  INVX2 U2468 ( .A(n2080), .Y(N824) );
  MUX2X1 U2469 ( .B(x[26]), .A(N305), .S(n2035), .Y(n2081) );
  MUX2X1 U2470 ( .B(x[25]), .A(N304), .S(n2035), .Y(n2082) );
  INVX2 U2471 ( .A(n2082), .Y(N822) );
  MUX2X1 U2472 ( .B(x[24]), .A(N303), .S(n2035), .Y(n2083) );
  MUX2X1 U2473 ( .B(x[23]), .A(N302), .S(n2035), .Y(n2084) );
  INVX2 U2474 ( .A(n2084), .Y(N820) );
  MUX2X1 U2475 ( .B(x[21]), .A(N300), .S(n2035), .Y(n2086) );
  INVX2 U2476 ( .A(n2086), .Y(N818) );
  MUX2X1 U2477 ( .B(x[18]), .A(N297), .S(n2035), .Y(n2089) );
  INVX2 U2478 ( .A(n2090), .Y(N814) );
  MUX2X1 U2479 ( .B(n1842), .A(N295), .S(n2035), .Y(n2091) );
  MUX2X1 U2480 ( .B(x[15]), .A(N294), .S(n2034), .Y(n2092) );
  MUX2X1 U2481 ( .B(x[14]), .A(N293), .S(n2034), .Y(n2093) );
  INVX2 U2482 ( .A(n2093), .Y(N811) );
  MUX2X1 U2483 ( .B(x[13]), .A(N292), .S(n2034), .Y(n2094) );
  MUX2X1 U2484 ( .B(x[11]), .A(N290), .S(n2034), .Y(n2096) );
  INVX2 U2485 ( .A(n2096), .Y(N808) );
  INVX2 U2486 ( .A(n2098), .Y(N806) );
  MUX2X1 U2487 ( .B(n1843), .A(N287), .S(n2034), .Y(n2099) );
  INVX2 U2488 ( .A(n2100), .Y(N804) );
  MUX2X1 U2489 ( .B(n1885), .A(N284), .S(n2034), .Y(n2102) );
  INVX2 U2490 ( .A(n2102), .Y(N802) );
  MUX2X1 U2491 ( .B(n1886), .A(N283), .S(n2034), .Y(n2103) );
  MUX2X1 U2492 ( .B(n1841), .A(N282), .S(n2034), .Y(n2104) );
  MUX2X1 U2493 ( .B(n1884), .A(N281), .S(n2034), .Y(n2105) );
  INVX2 U2494 ( .A(n2105), .Y(N799) );
  MUX2X1 U2495 ( .B(x[1]), .A(N280), .S(n2034), .Y(n2106) );
  INVX2 U2496 ( .A(n2106), .Y(N798) );
  MUX2X1 U2497 ( .B(n1859), .A(N279), .S(n2034), .Y(n2107) );
  INVX2 U2498 ( .A(N2177), .Y(n2110) );
  INVX2 U2499 ( .A(N2143), .Y(n2109) );
  XNOR2X1 U2500 ( .A(n2045), .B(n2034), .Y(n2108) );
  MUX2X1 U2501 ( .B(n2110), .A(n2109), .S(n1912), .Y(n3064) );
  INVX2 U2502 ( .A(N2176), .Y(n2112) );
  INVX2 U2503 ( .A(N2142), .Y(n2111) );
  MUX2X1 U2504 ( .B(n2112), .A(n2111), .S(n1912), .Y(n3063) );
  INVX2 U2505 ( .A(N2175), .Y(n2114) );
  INVX2 U2506 ( .A(N2141), .Y(n2113) );
  MUX2X1 U2507 ( .B(n2114), .A(n2113), .S(n1912), .Y(n3062) );
  INVX2 U2508 ( .A(N2174), .Y(n2116) );
  INVX2 U2509 ( .A(N2140), .Y(n2115) );
  MUX2X1 U2510 ( .B(n2116), .A(n2115), .S(n1912), .Y(n3061) );
  INVX2 U2511 ( .A(N2173), .Y(n2118) );
  INVX2 U2512 ( .A(N2139), .Y(n2117) );
  MUX2X1 U2513 ( .B(n2118), .A(n2117), .S(n1912), .Y(n3060) );
  INVX2 U2514 ( .A(N2172), .Y(n2120) );
  INVX2 U2515 ( .A(N2138), .Y(n2119) );
  MUX2X1 U2516 ( .B(n2120), .A(n2119), .S(n1912), .Y(n3059) );
  INVX2 U2517 ( .A(N2171), .Y(n2122) );
  INVX2 U2518 ( .A(N2137), .Y(n2121) );
  MUX2X1 U2519 ( .B(n2122), .A(n2121), .S(n1912), .Y(n3058) );
  INVX2 U2520 ( .A(N2170), .Y(n2124) );
  INVX2 U2521 ( .A(N2136), .Y(n2123) );
  MUX2X1 U2522 ( .B(n2124), .A(n2123), .S(n1912), .Y(n3057) );
  INVX2 U2523 ( .A(N2169), .Y(n2126) );
  INVX2 U2524 ( .A(N2135), .Y(n2125) );
  MUX2X1 U2525 ( .B(n2126), .A(n2125), .S(n1912), .Y(n3056) );
  INVX2 U2526 ( .A(N2168), .Y(n2128) );
  INVX2 U2527 ( .A(N2134), .Y(n2127) );
  MUX2X1 U2528 ( .B(n2128), .A(n2127), .S(n1912), .Y(n3055) );
  INVX2 U2529 ( .A(N2167), .Y(n2130) );
  INVX2 U2530 ( .A(N2133), .Y(n2129) );
  MUX2X1 U2531 ( .B(n2130), .A(n2129), .S(n1912), .Y(n3054) );
  INVX2 U2532 ( .A(N2166), .Y(n2132) );
  INVX2 U2533 ( .A(N2132), .Y(n2131) );
  MUX2X1 U2534 ( .B(n2132), .A(n2131), .S(n1912), .Y(n3053) );
  INVX2 U2535 ( .A(N2165), .Y(n2134) );
  INVX2 U2536 ( .A(N2131), .Y(n2133) );
  MUX2X1 U2537 ( .B(n2134), .A(n2133), .S(n1912), .Y(n3052) );
  INVX2 U2538 ( .A(N2164), .Y(n2136) );
  INVX2 U2539 ( .A(N2130), .Y(n2135) );
  MUX2X1 U2540 ( .B(n2136), .A(n2135), .S(n1912), .Y(n3051) );
  INVX2 U2541 ( .A(N2163), .Y(n2138) );
  INVX2 U2542 ( .A(N2129), .Y(n2137) );
  MUX2X1 U2543 ( .B(n2138), .A(n2137), .S(n1912), .Y(n3050) );
  INVX2 U2544 ( .A(N2162), .Y(n2140) );
  INVX2 U2545 ( .A(N2128), .Y(n2139) );
  MUX2X1 U2546 ( .B(n2140), .A(n2139), .S(n1912), .Y(n3049) );
  INVX2 U2547 ( .A(N2161), .Y(n2142) );
  INVX2 U2548 ( .A(N2127), .Y(n2141) );
  MUX2X1 U2549 ( .B(n2142), .A(n2141), .S(n1912), .Y(n3048) );
  INVX2 U2550 ( .A(N2160), .Y(n2144) );
  INVX2 U2551 ( .A(N2126), .Y(n2143) );
  MUX2X1 U2552 ( .B(n2144), .A(n2143), .S(n1912), .Y(n3047) );
  INVX2 U2553 ( .A(N2159), .Y(n2146) );
  INVX2 U2554 ( .A(N2125), .Y(n2145) );
  MUX2X1 U2555 ( .B(n2146), .A(n2145), .S(n1912), .Y(n3046) );
  INVX2 U2556 ( .A(N2158), .Y(n2148) );
  INVX2 U2557 ( .A(N2124), .Y(n2147) );
  MUX2X1 U2558 ( .B(n2148), .A(n2147), .S(n1912), .Y(n3045) );
  INVX2 U2559 ( .A(N2157), .Y(n2150) );
  INVX2 U2560 ( .A(N2123), .Y(n2149) );
  MUX2X1 U2561 ( .B(n2150), .A(n2149), .S(n1912), .Y(n3044) );
  INVX2 U2562 ( .A(N2156), .Y(n2152) );
  INVX2 U2563 ( .A(N2122), .Y(n2151) );
  MUX2X1 U2564 ( .B(n2152), .A(n2151), .S(n1912), .Y(n3043) );
  INVX2 U2565 ( .A(N2155), .Y(n2154) );
  INVX2 U2566 ( .A(N2121), .Y(n2153) );
  MUX2X1 U2567 ( .B(n2154), .A(n2153), .S(n1912), .Y(n3042) );
  INVX2 U2568 ( .A(N2154), .Y(n2156) );
  INVX2 U2569 ( .A(N2120), .Y(n2155) );
  MUX2X1 U2570 ( .B(n2156), .A(n2155), .S(n1912), .Y(n3041) );
  INVX2 U2571 ( .A(N2153), .Y(n2158) );
  INVX2 U2572 ( .A(N2119), .Y(n2157) );
  MUX2X1 U2573 ( .B(n2158), .A(n2157), .S(n1912), .Y(n3040) );
  INVX2 U2574 ( .A(N2152), .Y(n2160) );
  INVX2 U2575 ( .A(N2118), .Y(n2159) );
  MUX2X1 U2576 ( .B(n2160), .A(n2159), .S(n1912), .Y(n3039) );
  INVX2 U2577 ( .A(N2151), .Y(n2162) );
  INVX2 U2578 ( .A(N2117), .Y(n2161) );
  MUX2X1 U2579 ( .B(n2162), .A(n2161), .S(n1912), .Y(n3038) );
  INVX2 U2580 ( .A(N2150), .Y(n2164) );
  INVX2 U2581 ( .A(N2116), .Y(n2163) );
  MUX2X1 U2582 ( .B(n2164), .A(n2163), .S(n1912), .Y(n3037) );
  INVX2 U2583 ( .A(N2149), .Y(n2166) );
  INVX2 U2584 ( .A(N2115), .Y(n2165) );
  MUX2X1 U2585 ( .B(n2166), .A(n2165), .S(n1912), .Y(n3036) );
  INVX2 U2586 ( .A(N2148), .Y(n2168) );
  INVX2 U2587 ( .A(N2114), .Y(n2167) );
  MUX2X1 U2588 ( .B(n2168), .A(n2167), .S(n1912), .Y(n3035) );
  INVX2 U2589 ( .A(N2147), .Y(n2170) );
  INVX2 U2590 ( .A(N2113), .Y(n2169) );
  MUX2X1 U2591 ( .B(n2170), .A(n2169), .S(n1912), .Y(n3034) );
  INVX2 U2592 ( .A(N2146), .Y(n2172) );
  INVX2 U2593 ( .A(N2112), .Y(n2171) );
  MUX2X1 U2594 ( .B(n2172), .A(n2171), .S(n1912), .Y(n3033) );
  AND2X2 U2595 ( .A(N1788), .B(n2043), .Y(N1820) );
  INVX2 U2596 ( .A(N1787), .Y(n2173) );
  MUX2X1 U2597 ( .B(n3197), .A(n2173), .S(n2043), .Y(N1819) );
  INVX2 U2598 ( .A(N1786), .Y(n2174) );
  MUX2X1 U2599 ( .B(n3198), .A(n2174), .S(n2043), .Y(N1818) );
  INVX2 U2600 ( .A(N1785), .Y(n2175) );
  MUX2X1 U2601 ( .B(n3199), .A(n2175), .S(n2043), .Y(N1817) );
  INVX2 U2602 ( .A(N1784), .Y(n2176) );
  MUX2X1 U2603 ( .B(n3200), .A(n2176), .S(n2043), .Y(N1816) );
  INVX2 U2604 ( .A(N1783), .Y(n2177) );
  MUX2X1 U2605 ( .B(n3201), .A(n2177), .S(n2043), .Y(N1815) );
  INVX2 U2606 ( .A(N1782), .Y(n2178) );
  MUX2X1 U2607 ( .B(n3202), .A(n2178), .S(n2043), .Y(N1814) );
  INVX2 U2608 ( .A(N1781), .Y(n2179) );
  MUX2X1 U2609 ( .B(n3203), .A(n2179), .S(n2043), .Y(N1813) );
  INVX2 U2610 ( .A(N1780), .Y(n2180) );
  MUX2X1 U2611 ( .B(n3204), .A(n2180), .S(n2043), .Y(N1812) );
  INVX2 U2612 ( .A(N1779), .Y(n2181) );
  MUX2X1 U2613 ( .B(n3205), .A(n2181), .S(n2043), .Y(N1811) );
  INVX2 U2614 ( .A(N1778), .Y(n2182) );
  MUX2X1 U2615 ( .B(n3206), .A(n2182), .S(n2043), .Y(N1810) );
  INVX2 U2616 ( .A(N1777), .Y(n2183) );
  MUX2X1 U2617 ( .B(n3207), .A(n2183), .S(n2043), .Y(N1809) );
  INVX2 U2618 ( .A(N1776), .Y(n2184) );
  MUX2X1 U2619 ( .B(n3208), .A(n2184), .S(n2043), .Y(N1808) );
  INVX2 U2620 ( .A(N1775), .Y(n2185) );
  MUX2X1 U2621 ( .B(n3209), .A(n2185), .S(n2043), .Y(N1807) );
  INVX2 U2622 ( .A(N1774), .Y(n2186) );
  MUX2X1 U2623 ( .B(n3210), .A(n2186), .S(n2043), .Y(N1806) );
  INVX2 U2624 ( .A(N1773), .Y(n2187) );
  MUX2X1 U2625 ( .B(n3211), .A(n2187), .S(n2043), .Y(N1805) );
  INVX2 U2626 ( .A(N1772), .Y(n2188) );
  MUX2X1 U2627 ( .B(n3212), .A(n2188), .S(n2043), .Y(N1804) );
  INVX2 U2628 ( .A(N1771), .Y(n2189) );
  MUX2X1 U2629 ( .B(n3213), .A(n2189), .S(n2043), .Y(N1803) );
  INVX2 U2630 ( .A(N1770), .Y(n2190) );
  MUX2X1 U2631 ( .B(n3214), .A(n2190), .S(n2043), .Y(N1802) );
  INVX2 U2632 ( .A(N1769), .Y(n2191) );
  MUX2X1 U2633 ( .B(n3215), .A(n2191), .S(n2043), .Y(N1801) );
  INVX2 U2634 ( .A(N1768), .Y(n2192) );
  MUX2X1 U2635 ( .B(n3216), .A(n2192), .S(n2043), .Y(N1800) );
  INVX2 U2636 ( .A(N1767), .Y(n2193) );
  MUX2X1 U2637 ( .B(n3217), .A(n2193), .S(n2043), .Y(N1799) );
  INVX2 U2638 ( .A(N1766), .Y(n2194) );
  MUX2X1 U2639 ( .B(n3218), .A(n2194), .S(n2043), .Y(N1798) );
  INVX2 U2640 ( .A(N1765), .Y(n2195) );
  MUX2X1 U2641 ( .B(n3219), .A(n2195), .S(n2043), .Y(N1797) );
  INVX2 U2642 ( .A(N1764), .Y(n2196) );
  MUX2X1 U2643 ( .B(n3220), .A(n2196), .S(n2043), .Y(N1796) );
  INVX2 U2644 ( .A(N1763), .Y(n2197) );
  MUX2X1 U2645 ( .B(n3221), .A(n2197), .S(n2043), .Y(N1795) );
  INVX2 U2646 ( .A(N1762), .Y(n2198) );
  MUX2X1 U2647 ( .B(n3222), .A(n2198), .S(n2043), .Y(N1794) );
  INVX2 U2648 ( .A(N1761), .Y(n2199) );
  MUX2X1 U2649 ( .B(n3223), .A(n2199), .S(n2043), .Y(N1793) );
  INVX2 U2650 ( .A(N1760), .Y(n2200) );
  MUX2X1 U2651 ( .B(n3224), .A(n2200), .S(n2043), .Y(N1792) );
  INVX2 U2652 ( .A(N1759), .Y(n2201) );
  MUX2X1 U2653 ( .B(n3225), .A(n2201), .S(n2043), .Y(N1791) );
  INVX2 U2654 ( .A(N1758), .Y(n2202) );
  MUX2X1 U2655 ( .B(n3226), .A(n2202), .S(n2043), .Y(N1790) );
  INVX2 U2656 ( .A(N1757), .Y(n2203) );
  MUX2X1 U2657 ( .B(n3227), .A(n2203), .S(n2043), .Y(N1789) );
  MUX2X1 U2658 ( .B(t1[30]), .A(N520), .S(n2031), .Y(n2204) );
  MUX2X1 U2659 ( .B(t1[29]), .A(N519), .S(n2031), .Y(n2205) );
  MUX2X1 U2660 ( .B(t1[28]), .A(N518), .S(n2031), .Y(n2206) );
  MUX2X1 U2661 ( .B(t1[27]), .A(N517), .S(n2031), .Y(n2207) );
  MUX2X1 U2662 ( .B(t1[26]), .A(N516), .S(n2031), .Y(n2208) );
  MUX2X1 U2663 ( .B(t1[24]), .A(N514), .S(n2031), .Y(n2210) );
  INVX2 U2664 ( .A(n2210), .Y(n3026) );
  MUX2X1 U2665 ( .B(n1881), .A(N513), .S(n2031), .Y(n2211) );
  INVX2 U2666 ( .A(n2211), .Y(n3025) );
  MUX2X1 U2667 ( .B(t1[22]), .A(N512), .S(n2031), .Y(n2212) );
  INVX2 U2668 ( .A(n2212), .Y(n3024) );
  MUX2X1 U2669 ( .B(t1[21]), .A(N511), .S(n2031), .Y(n2213) );
  INVX2 U2670 ( .A(n2213), .Y(n3023) );
  MUX2X1 U2671 ( .B(t1[20]), .A(N510), .S(n2031), .Y(n2214) );
  INVX2 U2672 ( .A(n2214), .Y(n3022) );
  MUX2X1 U2673 ( .B(n1888), .A(N509), .S(n2031), .Y(n2215) );
  INVX2 U2674 ( .A(n2215), .Y(n3021) );
  MUX2X1 U2675 ( .B(t1[18]), .A(N508), .S(n2031), .Y(n2216) );
  MUX2X1 U2676 ( .B(t1[17]), .A(N507), .S(n2031), .Y(n2217) );
  INVX2 U2677 ( .A(n2217), .Y(n3019) );
  MUX2X1 U2678 ( .B(t1[16]), .A(N506), .S(n2031), .Y(n2218) );
  MUX2X1 U2679 ( .B(t1[15]), .A(N505), .S(n2032), .Y(n2219) );
  INVX2 U2680 ( .A(n2219), .Y(n3017) );
  MUX2X1 U2681 ( .B(t1[14]), .A(N504), .S(n2032), .Y(n2220) );
  INVX2 U2682 ( .A(n2220), .Y(n3016) );
  MUX2X1 U2683 ( .B(t1[13]), .A(N503), .S(n2032), .Y(n2221) );
  INVX2 U2684 ( .A(n2221), .Y(n3015) );
  MUX2X1 U2685 ( .B(t1[12]), .A(N502), .S(n2032), .Y(n2222) );
  MUX2X1 U2686 ( .B(t1[11]), .A(N501), .S(n2032), .Y(n2223) );
  MUX2X1 U2687 ( .B(t1[10]), .A(N500), .S(n2032), .Y(n2224) );
  MUX2X1 U2688 ( .B(t1[9]), .A(N499), .S(n2032), .Y(n2225) );
  MUX2X1 U2689 ( .B(t1[8]), .A(N498), .S(n2032), .Y(n2226) );
  INVX2 U2690 ( .A(n2226), .Y(n3010) );
  MUX2X1 U2691 ( .B(t1[7]), .A(N497), .S(n2032), .Y(n2227) );
  MUX2X1 U2692 ( .B(t1[6]), .A(N496), .S(n2032), .Y(n2228) );
  MUX2X1 U2693 ( .B(t1[5]), .A(N495), .S(n2032), .Y(n2229) );
  INVX2 U2694 ( .A(n2229), .Y(n3007) );
  MUX2X1 U2695 ( .B(t1[4]), .A(N494), .S(n2032), .Y(n2230) );
  INVX2 U2696 ( .A(n2230), .Y(n3006) );
  MUX2X1 U2697 ( .B(t1[3]), .A(N493), .S(n2032), .Y(n2231) );
  MUX2X1 U2698 ( .B(t1[2]), .A(N492), .S(n2032), .Y(n2232) );
  INVX2 U2699 ( .A(n2232), .Y(n3004) );
  MUX2X1 U2700 ( .B(t1[1]), .A(N491), .S(n2032), .Y(n2233) );
  MUX2X1 U2701 ( .B(t1[0]), .A(N490), .S(n2031), .Y(n2234) );
  INVX2 U2702 ( .A(N1932), .Y(n2237) );
  INVX2 U2703 ( .A(N1966), .Y(n2236) );
  XNOR2X1 U2704 ( .A(n2031), .B(n2043), .Y(n2235) );
  MUX2X1 U2705 ( .B(n2237), .A(n2236), .S(n1913), .Y(n3002) );
  INVX2 U2706 ( .A(N1931), .Y(n2239) );
  INVX2 U2707 ( .A(N1965), .Y(n2238) );
  MUX2X1 U2708 ( .B(n2239), .A(n2238), .S(n1913), .Y(n3001) );
  INVX2 U2709 ( .A(N1930), .Y(n2241) );
  INVX2 U2710 ( .A(N1964), .Y(n2240) );
  MUX2X1 U2711 ( .B(n2241), .A(n2240), .S(n1913), .Y(n3000) );
  INVX2 U2712 ( .A(N1929), .Y(n2243) );
  INVX2 U2713 ( .A(N1963), .Y(n2242) );
  MUX2X1 U2714 ( .B(n2243), .A(n2242), .S(n1913), .Y(n2999) );
  INVX2 U2715 ( .A(N1928), .Y(n2245) );
  INVX2 U2716 ( .A(N1962), .Y(n2244) );
  MUX2X1 U2717 ( .B(n2245), .A(n2244), .S(n1913), .Y(n2998) );
  INVX2 U2718 ( .A(N1927), .Y(n2247) );
  INVX2 U2719 ( .A(N1961), .Y(n2246) );
  MUX2X1 U2720 ( .B(n2247), .A(n2246), .S(n1913), .Y(n2997) );
  INVX2 U2721 ( .A(N1926), .Y(n2249) );
  INVX2 U2722 ( .A(N1960), .Y(n2248) );
  MUX2X1 U2723 ( .B(n2249), .A(n2248), .S(n1913), .Y(n2996) );
  INVX2 U2724 ( .A(N1925), .Y(n2251) );
  INVX2 U2725 ( .A(N1959), .Y(n2250) );
  MUX2X1 U2726 ( .B(n2251), .A(n2250), .S(n1913), .Y(n2995) );
  INVX2 U2727 ( .A(N1924), .Y(n2253) );
  INVX2 U2728 ( .A(N1958), .Y(n2252) );
  MUX2X1 U2729 ( .B(n2253), .A(n2252), .S(n1913), .Y(n2994) );
  INVX2 U2730 ( .A(N1923), .Y(n2255) );
  INVX2 U2731 ( .A(N1957), .Y(n2254) );
  MUX2X1 U2732 ( .B(n2255), .A(n2254), .S(n1913), .Y(n2993) );
  INVX2 U2733 ( .A(N1922), .Y(n2257) );
  INVX2 U2734 ( .A(N1956), .Y(n2256) );
  MUX2X1 U2735 ( .B(n2257), .A(n2256), .S(n1913), .Y(n2992) );
  INVX2 U2736 ( .A(N1921), .Y(n2259) );
  INVX2 U2737 ( .A(N1955), .Y(n2258) );
  MUX2X1 U2738 ( .B(n2259), .A(n2258), .S(n1913), .Y(n2991) );
  INVX2 U2739 ( .A(N1920), .Y(n2261) );
  INVX2 U2740 ( .A(N1954), .Y(n2260) );
  MUX2X1 U2741 ( .B(n2261), .A(n2260), .S(n1913), .Y(n2990) );
  INVX2 U2742 ( .A(N1919), .Y(n2263) );
  INVX2 U2743 ( .A(N1953), .Y(n2262) );
  MUX2X1 U2744 ( .B(n2263), .A(n2262), .S(n1913), .Y(n2989) );
  INVX2 U2745 ( .A(N1918), .Y(n2265) );
  INVX2 U2746 ( .A(N1952), .Y(n2264) );
  MUX2X1 U2747 ( .B(n2265), .A(n2264), .S(n1913), .Y(n2988) );
  INVX2 U2748 ( .A(N1917), .Y(n2267) );
  INVX2 U2749 ( .A(N1951), .Y(n2266) );
  MUX2X1 U2750 ( .B(n2267), .A(n2266), .S(n1913), .Y(n2987) );
  INVX2 U2751 ( .A(N1916), .Y(n2269) );
  INVX2 U2752 ( .A(N1950), .Y(n2268) );
  MUX2X1 U2753 ( .B(n2269), .A(n2268), .S(n1913), .Y(n2986) );
  INVX2 U2754 ( .A(N1915), .Y(n2271) );
  INVX2 U2755 ( .A(N1949), .Y(n2270) );
  MUX2X1 U2756 ( .B(n2271), .A(n2270), .S(n1913), .Y(n2985) );
  INVX2 U2757 ( .A(N1914), .Y(n2273) );
  INVX2 U2758 ( .A(N1948), .Y(n2272) );
  MUX2X1 U2759 ( .B(n2273), .A(n2272), .S(n1913), .Y(n2984) );
  INVX2 U2760 ( .A(N1913), .Y(n2275) );
  INVX2 U2761 ( .A(N1947), .Y(n2274) );
  MUX2X1 U2762 ( .B(n2275), .A(n2274), .S(n1913), .Y(n2983) );
  INVX2 U2763 ( .A(N1912), .Y(n2277) );
  INVX2 U2764 ( .A(N1946), .Y(n2276) );
  MUX2X1 U2765 ( .B(n2277), .A(n2276), .S(n1913), .Y(n2982) );
  INVX2 U2766 ( .A(N1911), .Y(n2279) );
  INVX2 U2767 ( .A(N1945), .Y(n2278) );
  MUX2X1 U2768 ( .B(n2279), .A(n2278), .S(n1913), .Y(n2981) );
  INVX2 U2769 ( .A(N1910), .Y(n2281) );
  INVX2 U2770 ( .A(N1944), .Y(n2280) );
  MUX2X1 U2771 ( .B(n2281), .A(n2280), .S(n1913), .Y(n2980) );
  INVX2 U2772 ( .A(N1909), .Y(n2283) );
  INVX2 U2773 ( .A(N1943), .Y(n2282) );
  MUX2X1 U2774 ( .B(n2283), .A(n2282), .S(n1913), .Y(n2979) );
  INVX2 U2775 ( .A(N1908), .Y(n2285) );
  INVX2 U2776 ( .A(N1942), .Y(n2284) );
  MUX2X1 U2777 ( .B(n2285), .A(n2284), .S(n1913), .Y(n2978) );
  INVX2 U2778 ( .A(N1907), .Y(n2287) );
  INVX2 U2779 ( .A(N1941), .Y(n2286) );
  MUX2X1 U2780 ( .B(n2287), .A(n2286), .S(n1913), .Y(n2977) );
  INVX2 U2781 ( .A(N1906), .Y(n2289) );
  INVX2 U2782 ( .A(N1940), .Y(n2288) );
  MUX2X1 U2783 ( .B(n2289), .A(n2288), .S(n1913), .Y(n2976) );
  INVX2 U2784 ( .A(N1905), .Y(n2291) );
  INVX2 U2785 ( .A(N1939), .Y(n2290) );
  MUX2X1 U2786 ( .B(n2291), .A(n2290), .S(n1913), .Y(n2975) );
  INVX2 U2787 ( .A(N1904), .Y(n2293) );
  INVX2 U2788 ( .A(N1938), .Y(n2292) );
  MUX2X1 U2789 ( .B(n2293), .A(n2292), .S(n1913), .Y(n2974) );
  INVX2 U2790 ( .A(N1903), .Y(n2295) );
  INVX2 U2791 ( .A(N1937), .Y(n2294) );
  MUX2X1 U2792 ( .B(n2295), .A(n2294), .S(n1913), .Y(n2973) );
  INVX2 U2793 ( .A(N1902), .Y(n2297) );
  INVX2 U2794 ( .A(N1936), .Y(n2296) );
  MUX2X1 U2795 ( .B(n2297), .A(n2296), .S(n1913), .Y(n2972) );
  INVX2 U2796 ( .A(N1901), .Y(n2299) );
  INVX2 U2797 ( .A(N1935), .Y(n2298) );
  MUX2X1 U2798 ( .B(n2299), .A(n2298), .S(n1913), .Y(n2971) );
  AND2X2 U2799 ( .A(N1577), .B(n2041), .Y(N1609) );
  INVX2 U2800 ( .A(N1576), .Y(n2300) );
  MUX2X1 U2801 ( .B(n3228), .A(n2300), .S(n2041), .Y(N1608) );
  INVX2 U2802 ( .A(N1575), .Y(n2301) );
  MUX2X1 U2803 ( .B(n3229), .A(n2301), .S(n2041), .Y(N1607) );
  INVX2 U2804 ( .A(N1574), .Y(n2302) );
  MUX2X1 U2805 ( .B(n3230), .A(n2302), .S(n2041), .Y(N1606) );
  INVX2 U2806 ( .A(N1573), .Y(n2303) );
  MUX2X1 U2807 ( .B(n3231), .A(n2303), .S(n2041), .Y(N1605) );
  INVX2 U2808 ( .A(N1572), .Y(n2304) );
  MUX2X1 U2809 ( .B(n3232), .A(n2304), .S(n2041), .Y(N1604) );
  INVX2 U2810 ( .A(N1571), .Y(n2305) );
  MUX2X1 U2811 ( .B(n3233), .A(n2305), .S(n2041), .Y(N1603) );
  INVX2 U2812 ( .A(N1570), .Y(n2306) );
  MUX2X1 U2813 ( .B(n3234), .A(n2306), .S(n2041), .Y(N1602) );
  INVX2 U2814 ( .A(N1569), .Y(n2307) );
  MUX2X1 U2815 ( .B(n3235), .A(n2307), .S(n2041), .Y(N1601) );
  INVX2 U2816 ( .A(N1568), .Y(n2308) );
  MUX2X1 U2817 ( .B(n3236), .A(n2308), .S(n2041), .Y(N1600) );
  INVX2 U2818 ( .A(N1567), .Y(n2309) );
  MUX2X1 U2819 ( .B(n3237), .A(n2309), .S(n2041), .Y(N1599) );
  INVX2 U2820 ( .A(N1566), .Y(n2310) );
  MUX2X1 U2821 ( .B(n3238), .A(n2310), .S(n2041), .Y(N1598) );
  INVX2 U2822 ( .A(N1565), .Y(n2311) );
  MUX2X1 U2823 ( .B(n3239), .A(n2311), .S(n2041), .Y(N1597) );
  INVX2 U2824 ( .A(N1564), .Y(n2312) );
  MUX2X1 U2825 ( .B(n3240), .A(n2312), .S(n2041), .Y(N1596) );
  INVX2 U2826 ( .A(N1563), .Y(n2313) );
  MUX2X1 U2827 ( .B(n3241), .A(n2313), .S(n2041), .Y(N1595) );
  INVX2 U2828 ( .A(N1562), .Y(n2314) );
  MUX2X1 U2829 ( .B(n3242), .A(n2314), .S(n2041), .Y(N1594) );
  INVX2 U2830 ( .A(N1561), .Y(n2315) );
  MUX2X1 U2831 ( .B(n3243), .A(n2315), .S(n2041), .Y(N1593) );
  INVX2 U2832 ( .A(N1560), .Y(n2316) );
  MUX2X1 U2833 ( .B(n3244), .A(n2316), .S(n2041), .Y(N1592) );
  INVX2 U2834 ( .A(N1559), .Y(n2317) );
  MUX2X1 U2835 ( .B(n3245), .A(n2317), .S(n2041), .Y(N1591) );
  INVX2 U2836 ( .A(N1558), .Y(n2318) );
  MUX2X1 U2837 ( .B(n3246), .A(n2318), .S(n2041), .Y(N1590) );
  INVX2 U2838 ( .A(N1557), .Y(n2319) );
  MUX2X1 U2839 ( .B(n3247), .A(n2319), .S(n2041), .Y(N1589) );
  INVX2 U2840 ( .A(N1556), .Y(n2320) );
  MUX2X1 U2841 ( .B(n3248), .A(n2320), .S(n2041), .Y(N1588) );
  INVX2 U2842 ( .A(N1555), .Y(n2321) );
  MUX2X1 U2843 ( .B(n3249), .A(n2321), .S(n2041), .Y(N1587) );
  INVX2 U2844 ( .A(N1554), .Y(n2322) );
  MUX2X1 U2845 ( .B(n3250), .A(n2322), .S(n2041), .Y(N1586) );
  INVX2 U2846 ( .A(N1553), .Y(n2323) );
  MUX2X1 U2847 ( .B(n3251), .A(n2323), .S(n2041), .Y(N1585) );
  INVX2 U2848 ( .A(N1552), .Y(n2324) );
  MUX2X1 U2849 ( .B(n3252), .A(n2324), .S(n2041), .Y(N1584) );
  INVX2 U2850 ( .A(N1551), .Y(n2325) );
  MUX2X1 U2851 ( .B(n3253), .A(n2325), .S(n2041), .Y(N1583) );
  INVX2 U2852 ( .A(N1550), .Y(n2326) );
  MUX2X1 U2853 ( .B(n3254), .A(n2326), .S(n2041), .Y(N1582) );
  INVX2 U2854 ( .A(N1549), .Y(n2327) );
  MUX2X1 U2855 ( .B(n3255), .A(n2327), .S(n2041), .Y(N1581) );
  INVX2 U2856 ( .A(N1548), .Y(n2328) );
  MUX2X1 U2857 ( .B(n3256), .A(n2328), .S(n2041), .Y(N1580) );
  INVX2 U2858 ( .A(N1547), .Y(n2329) );
  MUX2X1 U2859 ( .B(n3257), .A(n2329), .S(n2041), .Y(N1579) );
  INVX2 U2860 ( .A(N1546), .Y(n2330) );
  MUX2X1 U2861 ( .B(n3258), .A(n2330), .S(n2041), .Y(N1578) );
  XNOR2X1 U2862 ( .A(n2031), .B(n2034), .Y(n2331) );
  MUX2X1 U2863 ( .B(N665), .A(N699), .S(n1914), .Y(n2490) );
  MUX2X1 U2864 ( .B(N664), .A(N698), .S(n1914), .Y(n2332) );
  INVX2 U2865 ( .A(n2332), .Y(n2970) );
  MUX2X1 U2866 ( .B(N663), .A(N697), .S(n1914), .Y(n2333) );
  INVX2 U2867 ( .A(n2333), .Y(n2969) );
  MUX2X1 U2868 ( .B(N662), .A(N696), .S(n1914), .Y(n2334) );
  MUX2X1 U2869 ( .B(N661), .A(N695), .S(n1914), .Y(n2335) );
  INVX2 U2870 ( .A(n2335), .Y(n2967) );
  MUX2X1 U2871 ( .B(N660), .A(N694), .S(n1914), .Y(n2336) );
  INVX2 U2872 ( .A(n2336), .Y(n2966) );
  MUX2X1 U2873 ( .B(N659), .A(N693), .S(n1914), .Y(n2337) );
  MUX2X1 U2874 ( .B(N658), .A(N692), .S(n1914), .Y(n2338) );
  INVX2 U2875 ( .A(n2338), .Y(n2964) );
  MUX2X1 U2876 ( .B(N657), .A(N691), .S(n1914), .Y(n2339) );
  INVX2 U2877 ( .A(n2339), .Y(n2963) );
  MUX2X1 U2878 ( .B(N656), .A(N690), .S(n1914), .Y(n2340) );
  INVX2 U2879 ( .A(n2340), .Y(n2962) );
  MUX2X1 U2880 ( .B(N655), .A(N689), .S(n1914), .Y(n2341) );
  INVX2 U2881 ( .A(n2341), .Y(n2961) );
  MUX2X1 U2882 ( .B(N654), .A(N688), .S(n1914), .Y(n2342) );
  INVX2 U2883 ( .A(n2342), .Y(n2960) );
  MUX2X1 U2884 ( .B(N653), .A(N687), .S(n1914), .Y(n2343) );
  INVX2 U2885 ( .A(n2343), .Y(n2959) );
  MUX2X1 U2886 ( .B(n1864), .A(N686), .S(n1914), .Y(n2344) );
  INVX2 U2887 ( .A(n2344), .Y(n2958) );
  MUX2X1 U2888 ( .B(n1887), .A(N685), .S(n1914), .Y(n2345) );
  INVX2 U2889 ( .A(n2345), .Y(n2957) );
  MUX2X1 U2890 ( .B(N650), .A(N684), .S(n1914), .Y(n2346) );
  INVX2 U2891 ( .A(n2346), .Y(n2956) );
  MUX2X1 U2892 ( .B(N649), .A(N683), .S(n1914), .Y(n2347) );
  MUX2X1 U2893 ( .B(n1836), .A(N682), .S(n1914), .Y(n2348) );
  MUX2X1 U2894 ( .B(n1882), .A(N681), .S(n1914), .Y(n2349) );
  MUX2X1 U2895 ( .B(N646), .A(N680), .S(n1914), .Y(n2350) );
  INVX2 U2896 ( .A(n2350), .Y(n2952) );
  MUX2X1 U2897 ( .B(N645), .A(N679), .S(n1914), .Y(n2351) );
  MUX2X1 U2898 ( .B(N644), .A(N678), .S(n1914), .Y(n2352) );
  MUX2X1 U2899 ( .B(n1837), .A(N677), .S(n1914), .Y(n2353) );
  INVX2 U2900 ( .A(n2353), .Y(n2949) );
  MUX2X1 U2901 ( .B(N642), .A(N676), .S(n1914), .Y(n2354) );
  MUX2X1 U2902 ( .B(N641), .A(N675), .S(n1914), .Y(n2355) );
  INVX2 U2903 ( .A(n2355), .Y(n2947) );
  MUX2X1 U2904 ( .B(N640), .A(N674), .S(n1914), .Y(n2356) );
  INVX2 U2905 ( .A(n2356), .Y(n2946) );
  MUX2X1 U2906 ( .B(N639), .A(N673), .S(n1914), .Y(n2357) );
  MUX2X1 U2907 ( .B(N638), .A(N672), .S(n1914), .Y(n2358) );
  MUX2X1 U2908 ( .B(N637), .A(N671), .S(n1914), .Y(n2359) );
  INVX2 U2909 ( .A(n2359), .Y(n2943) );
  MUX2X1 U2910 ( .B(n1865), .A(N670), .S(n1914), .Y(n2360) );
  INVX2 U2911 ( .A(n2360), .Y(n2942) );
  MUX2X1 U2912 ( .B(N635), .A(N669), .S(n1914), .Y(n2361) );
  INVX2 U2913 ( .A(n2361), .Y(n2941) );
  MUX2X1 U2914 ( .B(N634), .A(N668), .S(n1914), .Y(n2362) );
  INVX2 U2915 ( .A(n2362), .Y(n2940) );
  NAND2X1 U2916 ( .A(N732), .B(n1868), .Y(n2363) );
  MUX2X1 U2917 ( .B(n2970), .A(N731), .S(n1867), .Y(n2364) );
  MUX2X1 U2918 ( .B(n2968), .A(N729), .S(n1874), .Y(n2366) );
  INVX2 U2919 ( .A(n2366), .Y(N761) );
  MUX2X1 U2920 ( .B(n2967), .A(N728), .S(n1869), .Y(n2367) );
  MUX2X1 U2921 ( .B(n2966), .A(N727), .S(n3067), .Y(n2368) );
  INVX2 U2922 ( .A(n2368), .Y(N759) );
  MUX2X1 U2923 ( .B(n2965), .A(N726), .S(n3067), .Y(n2369) );
  MUX2X1 U2924 ( .B(n2964), .A(N725), .S(n1870), .Y(n2370) );
  INVX2 U2925 ( .A(n2370), .Y(N757) );
  MUX2X1 U2926 ( .B(n2963), .A(N724), .S(n1872), .Y(n2371) );
  MUX2X1 U2927 ( .B(n2962), .A(N723), .S(n1871), .Y(n2372) );
  INVX2 U2928 ( .A(n2372), .Y(N755) );
  MUX2X1 U2929 ( .B(n2961), .A(N722), .S(n1867), .Y(n2373) );
  INVX2 U2930 ( .A(n2373), .Y(N754) );
  MUX2X1 U2931 ( .B(n2960), .A(N721), .S(n1875), .Y(n2374) );
  INVX2 U2932 ( .A(n2374), .Y(N753) );
  MUX2X1 U2933 ( .B(n2959), .A(N720), .S(n1867), .Y(n2375) );
  INVX2 U2934 ( .A(n2375), .Y(N752) );
  MUX2X1 U2935 ( .B(n2958), .A(N719), .S(n1867), .Y(n2376) );
  INVX2 U2936 ( .A(n2376), .Y(N751) );
  MUX2X1 U2937 ( .B(n2957), .A(N718), .S(n1866), .Y(n2377) );
  INVX2 U2938 ( .A(n2377), .Y(N750) );
  INVX2 U2939 ( .A(n2378), .Y(N749) );
  MUX2X1 U2940 ( .B(n2955), .A(N716), .S(n1875), .Y(n2379) );
  MUX2X1 U2941 ( .B(n2954), .A(N715), .S(n1877), .Y(n2380) );
  INVX2 U2942 ( .A(n2380), .Y(N747) );
  MUX2X1 U2943 ( .B(n2953), .A(N714), .S(n1876), .Y(n2381) );
  INVX2 U2944 ( .A(n2381), .Y(N746) );
  MUX2X1 U2945 ( .B(n2952), .A(N713), .S(n1872), .Y(n2382) );
  INVX2 U2946 ( .A(n2382), .Y(N745) );
  MUX2X1 U2947 ( .B(n2951), .A(N712), .S(n1870), .Y(n2383) );
  MUX2X1 U2948 ( .B(n2950), .A(N711), .S(n1872), .Y(n2384) );
  INVX2 U2949 ( .A(n2384), .Y(N743) );
  MUX2X1 U2950 ( .B(n2949), .A(N710), .S(n1874), .Y(n2385) );
  MUX2X1 U2951 ( .B(n2948), .A(N709), .S(n1876), .Y(n2386) );
  INVX2 U2952 ( .A(n2386), .Y(N741) );
  MUX2X1 U2953 ( .B(n2947), .A(N708), .S(n1877), .Y(n2387) );
  INVX2 U2954 ( .A(n2387), .Y(N740) );
  MUX2X1 U2955 ( .B(n2946), .A(N707), .S(n1871), .Y(n2388) );
  INVX2 U2956 ( .A(n2388), .Y(N739) );
  MUX2X1 U2957 ( .B(n2945), .A(N706), .S(n1869), .Y(n2389) );
  INVX2 U2958 ( .A(n2389), .Y(N738) );
  MUX2X1 U2959 ( .B(n2944), .A(N705), .S(n1876), .Y(n2390) );
  INVX2 U2960 ( .A(n2390), .Y(N737) );
  MUX2X1 U2961 ( .B(n2943), .A(N704), .S(n1873), .Y(n2391) );
  INVX2 U2962 ( .A(n2391), .Y(N736) );
  MUX2X1 U2963 ( .B(n2942), .A(N703), .S(n1866), .Y(n2392) );
  INVX2 U2964 ( .A(n2392), .Y(N735) );
  MUX2X1 U2965 ( .B(n2941), .A(N702), .S(n1868), .Y(n2393) );
  MUX2X1 U2966 ( .B(n2940), .A(N701), .S(n1876), .Y(n2394) );
  INVX2 U2967 ( .A(n2394), .Y(N733) );
  INVX2 U2968 ( .A(N1721), .Y(n2396) );
  INVX2 U2969 ( .A(N1755), .Y(n2395) );
  MUX2X1 U2970 ( .B(n2396), .A(n2395), .S(n1863), .Y(n2939) );
  INVX2 U2971 ( .A(N1720), .Y(n2398) );
  INVX2 U2972 ( .A(N1754), .Y(n2397) );
  MUX2X1 U2973 ( .B(n2398), .A(n2397), .S(n1863), .Y(n2938) );
  INVX2 U2974 ( .A(N1719), .Y(n2400) );
  INVX2 U2975 ( .A(N1753), .Y(n2399) );
  MUX2X1 U2976 ( .B(n2400), .A(n2399), .S(n1863), .Y(n2937) );
  INVX2 U2977 ( .A(N1718), .Y(n2402) );
  INVX2 U2978 ( .A(N1752), .Y(n2401) );
  MUX2X1 U2979 ( .B(n2402), .A(n2401), .S(n1863), .Y(n2936) );
  INVX2 U2980 ( .A(N1717), .Y(n2404) );
  INVX2 U2981 ( .A(N1751), .Y(n2403) );
  MUX2X1 U2982 ( .B(n2404), .A(n2403), .S(n1863), .Y(n2935) );
  INVX2 U2983 ( .A(N1716), .Y(n2406) );
  INVX2 U2984 ( .A(N1750), .Y(n2405) );
  MUX2X1 U2985 ( .B(n2406), .A(n2405), .S(n1863), .Y(n2934) );
  INVX2 U2986 ( .A(N1715), .Y(n2408) );
  INVX2 U2987 ( .A(N1749), .Y(n2407) );
  MUX2X1 U2988 ( .B(n2408), .A(n2407), .S(n1863), .Y(n2933) );
  INVX2 U2989 ( .A(N1714), .Y(n2410) );
  INVX2 U2990 ( .A(N1748), .Y(n2409) );
  MUX2X1 U2991 ( .B(n2410), .A(n2409), .S(n1863), .Y(n2932) );
  INVX2 U2992 ( .A(N1713), .Y(n2412) );
  INVX2 U2993 ( .A(N1747), .Y(n2411) );
  MUX2X1 U2994 ( .B(n2412), .A(n2411), .S(n1863), .Y(n2931) );
  INVX2 U2995 ( .A(N1712), .Y(n2414) );
  INVX2 U2996 ( .A(N1746), .Y(n2413) );
  MUX2X1 U2997 ( .B(n2414), .A(n2413), .S(n1863), .Y(n2930) );
  INVX2 U2998 ( .A(N1711), .Y(n2416) );
  INVX2 U2999 ( .A(N1745), .Y(n2415) );
  MUX2X1 U3000 ( .B(n2416), .A(n2415), .S(n1863), .Y(n2929) );
  INVX2 U3001 ( .A(N1710), .Y(n2418) );
  INVX2 U3002 ( .A(N1744), .Y(n2417) );
  MUX2X1 U3003 ( .B(n2418), .A(n2417), .S(n1863), .Y(n2928) );
  INVX2 U3004 ( .A(N1709), .Y(n2420) );
  INVX2 U3005 ( .A(N1743), .Y(n2419) );
  MUX2X1 U3006 ( .B(n2420), .A(n2419), .S(n1863), .Y(n2927) );
  INVX2 U3007 ( .A(N1708), .Y(n2422) );
  INVX2 U3008 ( .A(N1742), .Y(n2421) );
  MUX2X1 U3009 ( .B(n2422), .A(n2421), .S(n1863), .Y(n2926) );
  INVX2 U3010 ( .A(N1707), .Y(n2424) );
  INVX2 U3011 ( .A(N1741), .Y(n2423) );
  MUX2X1 U3012 ( .B(n2424), .A(n2423), .S(n1863), .Y(n2925) );
  INVX2 U3013 ( .A(N1706), .Y(n2426) );
  INVX2 U3014 ( .A(N1740), .Y(n2425) );
  MUX2X1 U3015 ( .B(n2426), .A(n2425), .S(n1863), .Y(n2924) );
  INVX2 U3016 ( .A(N1705), .Y(n2428) );
  INVX2 U3017 ( .A(N1739), .Y(n2427) );
  MUX2X1 U3018 ( .B(n2428), .A(n2427), .S(n1863), .Y(n2923) );
  INVX2 U3019 ( .A(N1704), .Y(n2430) );
  INVX2 U3020 ( .A(N1738), .Y(n2429) );
  MUX2X1 U3021 ( .B(n2430), .A(n2429), .S(n1863), .Y(n2922) );
  INVX2 U3022 ( .A(N1703), .Y(n2432) );
  INVX2 U3023 ( .A(N1737), .Y(n2431) );
  MUX2X1 U3024 ( .B(n2432), .A(n2431), .S(n1863), .Y(n2921) );
  INVX2 U3025 ( .A(N1702), .Y(n2434) );
  INVX2 U3026 ( .A(N1736), .Y(n2433) );
  MUX2X1 U3027 ( .B(n2434), .A(n2433), .S(n1915), .Y(n2920) );
  INVX2 U3028 ( .A(N1701), .Y(n2436) );
  INVX2 U3029 ( .A(N1735), .Y(n2435) );
  MUX2X1 U3030 ( .B(n2436), .A(n2435), .S(n1915), .Y(n2919) );
  INVX2 U3031 ( .A(N1700), .Y(n2438) );
  INVX2 U3032 ( .A(N1734), .Y(n2437) );
  MUX2X1 U3033 ( .B(n2438), .A(n2437), .S(n1915), .Y(n2918) );
  INVX2 U3034 ( .A(N1699), .Y(n2440) );
  INVX2 U3035 ( .A(N1733), .Y(n2439) );
  MUX2X1 U3036 ( .B(n2440), .A(n2439), .S(n1915), .Y(n2917) );
  INVX2 U3037 ( .A(N1698), .Y(n2442) );
  INVX2 U3038 ( .A(N1732), .Y(n2441) );
  MUX2X1 U3039 ( .B(n2442), .A(n2441), .S(n1915), .Y(n2916) );
  INVX2 U3040 ( .A(N1697), .Y(n2444) );
  INVX2 U3041 ( .A(N1731), .Y(n2443) );
  MUX2X1 U3042 ( .B(n2444), .A(n2443), .S(n1915), .Y(n2915) );
  INVX2 U3043 ( .A(N1696), .Y(n2446) );
  INVX2 U3044 ( .A(N1730), .Y(n2445) );
  MUX2X1 U3045 ( .B(n2446), .A(n2445), .S(n1915), .Y(n2914) );
  INVX2 U3046 ( .A(N1695), .Y(n2448) );
  INVX2 U3047 ( .A(N1729), .Y(n2447) );
  MUX2X1 U3048 ( .B(n2448), .A(n2447), .S(n1915), .Y(n2913) );
  INVX2 U3049 ( .A(N1694), .Y(n2450) );
  INVX2 U3050 ( .A(N1728), .Y(n2449) );
  MUX2X1 U3051 ( .B(n2450), .A(n2449), .S(n1915), .Y(n2912) );
  INVX2 U3052 ( .A(N1693), .Y(n2452) );
  INVX2 U3053 ( .A(N1727), .Y(n2451) );
  MUX2X1 U3054 ( .B(n2452), .A(n2451), .S(n1915), .Y(n2911) );
  INVX2 U3055 ( .A(N1692), .Y(n2454) );
  INVX2 U3056 ( .A(N1726), .Y(n2453) );
  MUX2X1 U3057 ( .B(n2454), .A(n2453), .S(n1915), .Y(n2910) );
  INVX2 U3058 ( .A(N1691), .Y(n2456) );
  INVX2 U3059 ( .A(N1725), .Y(n2455) );
  MUX2X1 U3060 ( .B(n2456), .A(n2455), .S(n1915), .Y(n2909) );
  INVX2 U3061 ( .A(N1690), .Y(n2458) );
  INVX2 U3062 ( .A(N1724), .Y(n2457) );
  MUX2X1 U3063 ( .B(n2458), .A(n2457), .S(n1915), .Y(n2908) );
  AND2X2 U3064 ( .A(N1366), .B(n2039), .Y(N1398) );
  INVX2 U3065 ( .A(N1365), .Y(n2459) );
  MUX2X1 U3066 ( .B(n3104), .A(n2459), .S(n2039), .Y(N1397) );
  INVX2 U3067 ( .A(N1364), .Y(n2460) );
  MUX2X1 U3068 ( .B(n3105), .A(n2460), .S(n2039), .Y(N1396) );
  INVX2 U3069 ( .A(N1363), .Y(n2461) );
  MUX2X1 U3070 ( .B(n3106), .A(n2461), .S(n2039), .Y(N1395) );
  INVX2 U3071 ( .A(N1362), .Y(n2462) );
  MUX2X1 U3072 ( .B(n3107), .A(n2462), .S(n2039), .Y(N1394) );
  INVX2 U3073 ( .A(N1361), .Y(n2463) );
  MUX2X1 U3074 ( .B(n3108), .A(n2463), .S(n2039), .Y(N1393) );
  INVX2 U3075 ( .A(N1360), .Y(n2464) );
  MUX2X1 U3076 ( .B(n3109), .A(n2464), .S(n2039), .Y(N1392) );
  INVX2 U3077 ( .A(N1359), .Y(n2465) );
  MUX2X1 U3078 ( .B(n3110), .A(n2465), .S(n2039), .Y(N1391) );
  INVX2 U3079 ( .A(N1358), .Y(n2466) );
  MUX2X1 U3080 ( .B(n3111), .A(n2466), .S(n2039), .Y(N1390) );
  INVX2 U3081 ( .A(N1357), .Y(n2467) );
  MUX2X1 U3082 ( .B(n3112), .A(n2467), .S(n2039), .Y(N1389) );
  INVX2 U3083 ( .A(N1356), .Y(n2468) );
  MUX2X1 U3084 ( .B(n3113), .A(n2468), .S(n2039), .Y(N1388) );
  INVX2 U3085 ( .A(N1355), .Y(n2469) );
  MUX2X1 U3086 ( .B(n3114), .A(n2469), .S(n2039), .Y(N1387) );
  INVX2 U3087 ( .A(N1354), .Y(n2470) );
  MUX2X1 U3088 ( .B(n3115), .A(n2470), .S(n2039), .Y(N1386) );
  INVX2 U3089 ( .A(N1353), .Y(n2471) );
  MUX2X1 U3090 ( .B(n3116), .A(n2471), .S(n2039), .Y(N1385) );
  INVX2 U3091 ( .A(N1352), .Y(n2472) );
  MUX2X1 U3092 ( .B(n3117), .A(n2472), .S(n2039), .Y(N1384) );
  INVX2 U3093 ( .A(N1351), .Y(n2473) );
  MUX2X1 U3094 ( .B(n3118), .A(n2473), .S(n2039), .Y(N1383) );
  INVX2 U3095 ( .A(N1350), .Y(n2474) );
  MUX2X1 U3096 ( .B(n3119), .A(n2474), .S(n2039), .Y(N1382) );
  INVX2 U3097 ( .A(N1349), .Y(n2475) );
  MUX2X1 U3098 ( .B(n3120), .A(n2475), .S(n2039), .Y(N1381) );
  INVX2 U3099 ( .A(N1348), .Y(n2476) );
  MUX2X1 U3100 ( .B(n3121), .A(n2476), .S(n2039), .Y(N1380) );
  INVX2 U3101 ( .A(N1347), .Y(n2477) );
  MUX2X1 U3102 ( .B(n3122), .A(n2477), .S(n2039), .Y(N1379) );
  INVX2 U3103 ( .A(N1346), .Y(n2478) );
  MUX2X1 U3104 ( .B(n3123), .A(n2478), .S(n2039), .Y(N1378) );
  INVX2 U3105 ( .A(N1345), .Y(n2479) );
  MUX2X1 U3106 ( .B(n3124), .A(n2479), .S(n2039), .Y(N1377) );
  INVX2 U3107 ( .A(N1344), .Y(n2480) );
  MUX2X1 U3108 ( .B(n3125), .A(n2480), .S(n2039), .Y(N1376) );
  INVX2 U3109 ( .A(N1343), .Y(n2481) );
  MUX2X1 U3110 ( .B(n3126), .A(n2481), .S(n2039), .Y(N1375) );
  INVX2 U3111 ( .A(N1342), .Y(n2482) );
  MUX2X1 U3112 ( .B(n3127), .A(n2482), .S(n2039), .Y(N1374) );
  INVX2 U3113 ( .A(N1341), .Y(n2483) );
  MUX2X1 U3114 ( .B(n3128), .A(n2483), .S(n2039), .Y(N1373) );
  INVX2 U3115 ( .A(N1340), .Y(n2484) );
  MUX2X1 U3116 ( .B(n3129), .A(n2484), .S(n2039), .Y(N1372) );
  INVX2 U3117 ( .A(N1339), .Y(n2485) );
  MUX2X1 U3118 ( .B(n3130), .A(n2485), .S(n2039), .Y(N1371) );
  INVX2 U3119 ( .A(N1338), .Y(n2486) );
  MUX2X1 U3120 ( .B(n3131), .A(n2486), .S(n2039), .Y(N1370) );
  INVX2 U3121 ( .A(N1337), .Y(n2487) );
  MUX2X1 U3122 ( .B(n3132), .A(n2487), .S(n2039), .Y(N1369) );
  INVX2 U3123 ( .A(N1336), .Y(n2488) );
  MUX2X1 U3124 ( .B(n3133), .A(n2488), .S(n2039), .Y(N1368) );
  INVX2 U3125 ( .A(N1335), .Y(n2489) );
  MUX2X1 U3126 ( .B(n3134), .A(n2489), .S(n2039), .Y(N1367) );
  MUX2X1 U3127 ( .B(N876), .A(N910), .S(n1917), .Y(n2650) );
  MUX2X1 U3128 ( .B(N875), .A(N909), .S(n1917), .Y(n2491) );
  INVX2 U3129 ( .A(n2491), .Y(n2907) );
  MUX2X1 U3130 ( .B(N874), .A(N908), .S(n1917), .Y(n2492) );
  INVX2 U3131 ( .A(n2492), .Y(n2906) );
  MUX2X1 U3132 ( .B(N873), .A(N907), .S(n1917), .Y(n2493) );
  INVX2 U3133 ( .A(n2493), .Y(n2905) );
  MUX2X1 U3134 ( .B(N872), .A(N906), .S(n1917), .Y(n2494) );
  INVX2 U3135 ( .A(n2494), .Y(n2904) );
  MUX2X1 U3136 ( .B(N871), .A(N905), .S(n1917), .Y(n2495) );
  INVX2 U3137 ( .A(n2495), .Y(n2903) );
  MUX2X1 U3138 ( .B(N870), .A(N904), .S(n1917), .Y(n2496) );
  INVX2 U3139 ( .A(n2496), .Y(n2902) );
  MUX2X1 U3140 ( .B(N869), .A(N903), .S(n1917), .Y(n2497) );
  INVX2 U3141 ( .A(n2497), .Y(n2901) );
  MUX2X1 U3142 ( .B(N868), .A(N902), .S(n1917), .Y(n2498) );
  INVX2 U3143 ( .A(n2498), .Y(n2900) );
  MUX2X1 U3144 ( .B(N867), .A(N901), .S(n1917), .Y(n2499) );
  INVX2 U3145 ( .A(n2499), .Y(n2899) );
  MUX2X1 U3146 ( .B(N866), .A(N900), .S(n1917), .Y(n2500) );
  INVX2 U3147 ( .A(n2500), .Y(n2898) );
  MUX2X1 U3148 ( .B(N865), .A(N899), .S(n1917), .Y(n2501) );
  INVX2 U3149 ( .A(n2501), .Y(n2897) );
  MUX2X1 U3150 ( .B(N864), .A(N898), .S(n1917), .Y(n2502) );
  INVX2 U3151 ( .A(n2502), .Y(n2896) );
  MUX2X1 U3152 ( .B(N863), .A(N897), .S(n1917), .Y(n2503) );
  INVX2 U3153 ( .A(n2503), .Y(n2895) );
  MUX2X1 U3154 ( .B(n1840), .A(N896), .S(n1917), .Y(n2504) );
  INVX2 U3155 ( .A(n2504), .Y(n2894) );
  MUX2X1 U3156 ( .B(N861), .A(N895), .S(n1917), .Y(n2505) );
  INVX2 U3157 ( .A(n2505), .Y(n2893) );
  MUX2X1 U3158 ( .B(N860), .A(N894), .S(n1917), .Y(n2506) );
  INVX2 U3159 ( .A(n2506), .Y(n2892) );
  MUX2X1 U3160 ( .B(N859), .A(N893), .S(n1917), .Y(n2507) );
  INVX2 U3161 ( .A(n2507), .Y(n2891) );
  MUX2X1 U3162 ( .B(N858), .A(N892), .S(n1917), .Y(n2508) );
  MUX2X1 U3163 ( .B(N857), .A(N891), .S(n1917), .Y(n2509) );
  INVX2 U3164 ( .A(n2509), .Y(n2889) );
  MUX2X1 U3165 ( .B(N856), .A(N890), .S(n1917), .Y(n2510) );
  INVX2 U3166 ( .A(n2510), .Y(n2888) );
  MUX2X1 U3167 ( .B(N855), .A(N889), .S(n1917), .Y(n2511) );
  INVX2 U3168 ( .A(n2511), .Y(n2887) );
  MUX2X1 U3169 ( .B(N854), .A(N888), .S(n1917), .Y(n2512) );
  MUX2X1 U3170 ( .B(N853), .A(N887), .S(n1917), .Y(n2513) );
  MUX2X1 U3171 ( .B(N852), .A(N886), .S(n1917), .Y(n2514) );
  INVX2 U3172 ( .A(n2514), .Y(n2884) );
  MUX2X1 U3173 ( .B(N851), .A(N885), .S(n1917), .Y(n2515) );
  INVX2 U3174 ( .A(n2515), .Y(n2883) );
  MUX2X1 U3175 ( .B(N850), .A(N884), .S(n1917), .Y(n2516) );
  INVX2 U3176 ( .A(n2516), .Y(n2882) );
  MUX2X1 U3177 ( .B(N849), .A(N883), .S(n1917), .Y(n2517) );
  INVX2 U3178 ( .A(n2517), .Y(n2881) );
  MUX2X1 U3179 ( .B(N848), .A(N882), .S(n1917), .Y(n2518) );
  INVX2 U3180 ( .A(n2518), .Y(n2880) );
  MUX2X1 U3181 ( .B(N847), .A(N881), .S(n1917), .Y(n2519) );
  INVX2 U3182 ( .A(n2519), .Y(n2879) );
  MUX2X1 U3183 ( .B(N846), .A(N880), .S(n1917), .Y(n2520) );
  INVX2 U3184 ( .A(n2520), .Y(n2878) );
  MUX2X1 U3185 ( .B(N845), .A(N879), .S(n1917), .Y(n2521) );
  INVX2 U3186 ( .A(n2521), .Y(n2877) );
  NAND2X1 U3187 ( .A(N943), .B(n1908), .Y(n2522) );
  MUX2X1 U3188 ( .B(n2907), .A(N942), .S(n1908), .Y(n2523) );
  INVX2 U3189 ( .A(n2523), .Y(N974) );
  MUX2X1 U3190 ( .B(n2906), .A(N941), .S(n1902), .Y(n2524) );
  MUX2X1 U3191 ( .B(n2905), .A(N940), .S(n1909), .Y(n2525) );
  INVX2 U3192 ( .A(n2525), .Y(N972) );
  MUX2X1 U3193 ( .B(n2903), .A(N938), .S(n1910), .Y(n2527) );
  MUX2X1 U3194 ( .B(n2902), .A(N937), .S(n1895), .Y(n2528) );
  INVX2 U3195 ( .A(n2529), .Y(N968) );
  MUX2X1 U3196 ( .B(n2899), .A(N934), .S(n1908), .Y(n2531) );
  INVX2 U3197 ( .A(n2531), .Y(N966) );
  MUX2X1 U3198 ( .B(n2897), .A(N932), .S(n1901), .Y(n2533) );
  INVX2 U3199 ( .A(n2533), .Y(N964) );
  MUX2X1 U3200 ( .B(n2896), .A(N931), .S(n1910), .Y(n2534) );
  INVX2 U3201 ( .A(n2535), .Y(N962) );
  INVX2 U3202 ( .A(n2536), .Y(N961) );
  INVX2 U3203 ( .A(n2537), .Y(N960) );
  MUX2X1 U3204 ( .B(n2892), .A(N927), .S(n1909), .Y(n2538) );
  MUX2X1 U3205 ( .B(n2890), .A(N925), .S(n1925), .Y(n2540) );
  MUX2X1 U3206 ( .B(n2888), .A(N923), .S(n1902), .Y(n2542) );
  MUX2X1 U3207 ( .B(n2884), .A(N919), .S(n1925), .Y(n2546) );
  MUX2X1 U3208 ( .B(n2882), .A(N917), .S(n3066), .Y(n2548) );
  MUX2X1 U3209 ( .B(n2880), .A(N915), .S(n1856), .Y(n2550) );
  MUX2X1 U3210 ( .B(n2879), .A(N914), .S(n1901), .Y(n2551) );
  MUX2X1 U3211 ( .B(n2878), .A(N913), .S(n3066), .Y(n2552) );
  INVX2 U3212 ( .A(n2553), .Y(N944) );
  INVX2 U3213 ( .A(N1510), .Y(n2556) );
  INVX2 U3214 ( .A(N1544), .Y(n2555) );
  XNOR2X1 U3215 ( .A(n1904), .B(n2040), .Y(n2554) );
  MUX2X1 U3216 ( .B(n2556), .A(n2555), .S(n1918), .Y(n2876) );
  INVX2 U3217 ( .A(N1509), .Y(n2558) );
  MUX2X1 U3218 ( .B(n2558), .A(n2557), .S(n1918), .Y(n2875) );
  INVX2 U3219 ( .A(N1508), .Y(n2560) );
  INVX2 U3220 ( .A(N1542), .Y(n2559) );
  MUX2X1 U3221 ( .B(n2560), .A(n2559), .S(n1918), .Y(n2874) );
  INVX2 U3222 ( .A(N1507), .Y(n2562) );
  INVX2 U3223 ( .A(N1541), .Y(n2561) );
  MUX2X1 U3224 ( .B(n2562), .A(n2561), .S(n1918), .Y(n2873) );
  INVX2 U3225 ( .A(N1506), .Y(n2564) );
  INVX2 U3226 ( .A(N1540), .Y(n2563) );
  MUX2X1 U3227 ( .B(n2564), .A(n2563), .S(n1918), .Y(n2872) );
  INVX2 U3228 ( .A(N1505), .Y(n2566) );
  INVX2 U3229 ( .A(N1539), .Y(n2565) );
  MUX2X1 U3230 ( .B(n2566), .A(n2565), .S(n1918), .Y(n2871) );
  INVX2 U3231 ( .A(N1504), .Y(n2568) );
  INVX2 U3232 ( .A(N1538), .Y(n2567) );
  MUX2X1 U3233 ( .B(n2568), .A(n2567), .S(n1918), .Y(n2870) );
  INVX2 U3234 ( .A(N1503), .Y(n2570) );
  INVX2 U3235 ( .A(N1537), .Y(n2569) );
  MUX2X1 U3236 ( .B(n2570), .A(n2569), .S(n1918), .Y(n2869) );
  INVX2 U3237 ( .A(N1502), .Y(n2572) );
  INVX2 U3238 ( .A(N1536), .Y(n2571) );
  MUX2X1 U3239 ( .B(n2572), .A(n2571), .S(n1918), .Y(n2868) );
  INVX2 U3240 ( .A(N1501), .Y(n2574) );
  INVX2 U3241 ( .A(N1535), .Y(n2573) );
  MUX2X1 U3242 ( .B(n2574), .A(n2573), .S(n1918), .Y(n2867) );
  INVX2 U3243 ( .A(N1500), .Y(n2576) );
  INVX2 U3244 ( .A(N1534), .Y(n2575) );
  MUX2X1 U3245 ( .B(n2576), .A(n2575), .S(n1918), .Y(n2866) );
  INVX2 U3246 ( .A(N1499), .Y(n2578) );
  INVX2 U3247 ( .A(N1533), .Y(n2577) );
  MUX2X1 U3248 ( .B(n2578), .A(n2577), .S(n1918), .Y(n2865) );
  INVX2 U3249 ( .A(N1498), .Y(n2580) );
  INVX2 U3250 ( .A(N1532), .Y(n2579) );
  MUX2X1 U3251 ( .B(n2580), .A(n2579), .S(n1918), .Y(n2864) );
  INVX2 U3252 ( .A(N1497), .Y(n2582) );
  INVX2 U3253 ( .A(N1531), .Y(n2581) );
  MUX2X1 U3254 ( .B(n2582), .A(n2581), .S(n1918), .Y(n2863) );
  INVX2 U3255 ( .A(N1496), .Y(n2584) );
  INVX2 U3256 ( .A(N1530), .Y(n2583) );
  MUX2X1 U3257 ( .B(n2584), .A(n2583), .S(n1918), .Y(n2862) );
  INVX2 U3258 ( .A(N1495), .Y(n2586) );
  INVX2 U3259 ( .A(N1529), .Y(n2585) );
  MUX2X1 U3260 ( .B(n2586), .A(n2585), .S(n1918), .Y(n2861) );
  INVX2 U3261 ( .A(N1494), .Y(n2588) );
  INVX2 U3262 ( .A(N1528), .Y(n2587) );
  MUX2X1 U3263 ( .B(n2588), .A(n2587), .S(n1918), .Y(n2860) );
  INVX2 U3264 ( .A(N1493), .Y(n2590) );
  INVX2 U3265 ( .A(N1527), .Y(n2589) );
  MUX2X1 U3266 ( .B(n2590), .A(n2589), .S(n1918), .Y(n2859) );
  INVX2 U3267 ( .A(N1492), .Y(n2592) );
  INVX2 U3268 ( .A(N1526), .Y(n2591) );
  MUX2X1 U3269 ( .B(n2592), .A(n2591), .S(n1918), .Y(n2858) );
  INVX2 U3270 ( .A(N1491), .Y(n2594) );
  INVX2 U3271 ( .A(N1525), .Y(n2593) );
  MUX2X1 U3272 ( .B(n2594), .A(n2593), .S(n1918), .Y(n2857) );
  INVX2 U3273 ( .A(N1490), .Y(n2596) );
  INVX2 U3274 ( .A(N1524), .Y(n2595) );
  MUX2X1 U3275 ( .B(n2596), .A(n2595), .S(n1918), .Y(n2856) );
  INVX2 U3276 ( .A(N1489), .Y(n2598) );
  INVX2 U3277 ( .A(N1523), .Y(n2597) );
  MUX2X1 U3278 ( .B(n2598), .A(n2597), .S(n1918), .Y(n2855) );
  INVX2 U3279 ( .A(N1488), .Y(n2600) );
  INVX2 U3280 ( .A(N1522), .Y(n2599) );
  MUX2X1 U3281 ( .B(n2600), .A(n2599), .S(n1918), .Y(n2854) );
  INVX2 U3282 ( .A(N1487), .Y(n2602) );
  INVX2 U3283 ( .A(N1521), .Y(n2601) );
  MUX2X1 U3284 ( .B(n2602), .A(n2601), .S(n1918), .Y(n2853) );
  INVX2 U3285 ( .A(N1486), .Y(n2604) );
  INVX2 U3286 ( .A(N1520), .Y(n2603) );
  MUX2X1 U3287 ( .B(n2604), .A(n2603), .S(n1918), .Y(n2852) );
  INVX2 U3288 ( .A(N1485), .Y(n2606) );
  INVX2 U3289 ( .A(N1519), .Y(n2605) );
  MUX2X1 U3290 ( .B(n2606), .A(n2605), .S(n1918), .Y(n2851) );
  INVX2 U3291 ( .A(N1484), .Y(n2608) );
  INVX2 U3292 ( .A(N1518), .Y(n2607) );
  MUX2X1 U3293 ( .B(n2608), .A(n2607), .S(n1918), .Y(n2850) );
  INVX2 U3294 ( .A(N1483), .Y(n2610) );
  INVX2 U3295 ( .A(N1517), .Y(n2609) );
  MUX2X1 U3296 ( .B(n2610), .A(n2609), .S(n1918), .Y(n2849) );
  INVX2 U3297 ( .A(N1482), .Y(n2612) );
  INVX2 U3298 ( .A(N1516), .Y(n2611) );
  MUX2X1 U3299 ( .B(n2612), .A(n2611), .S(n1918), .Y(n2848) );
  INVX2 U3300 ( .A(N1481), .Y(n2614) );
  INVX2 U3301 ( .A(N1515), .Y(n2613) );
  MUX2X1 U3302 ( .B(n2614), .A(n2613), .S(n1918), .Y(n2847) );
  INVX2 U3303 ( .A(N1480), .Y(n2616) );
  INVX2 U3304 ( .A(N1514), .Y(n2615) );
  MUX2X1 U3305 ( .B(n2616), .A(n2615), .S(n1918), .Y(n2846) );
  INVX2 U3306 ( .A(N1479), .Y(n2618) );
  INVX2 U3307 ( .A(N1513), .Y(n2617) );
  MUX2X1 U3308 ( .B(n2618), .A(n2617), .S(n1918), .Y(n2845) );
  AND2X2 U3309 ( .A(N1154), .B(n2037), .Y(N1186) );
  INVX2 U3310 ( .A(N1153), .Y(n2619) );
  MUX2X1 U3311 ( .B(n3135), .A(n2619), .S(n2037), .Y(N1185) );
  INVX2 U3312 ( .A(N1152), .Y(n2620) );
  MUX2X1 U3313 ( .B(n3136), .A(n2620), .S(n2037), .Y(N1184) );
  INVX2 U3314 ( .A(N1151), .Y(n2621) );
  MUX2X1 U3315 ( .B(n3137), .A(n2621), .S(n2037), .Y(N1183) );
  INVX2 U3316 ( .A(N1150), .Y(n2622) );
  MUX2X1 U3317 ( .B(n3138), .A(n2622), .S(n2037), .Y(N1182) );
  INVX2 U3318 ( .A(N1149), .Y(n2623) );
  MUX2X1 U3319 ( .B(n3139), .A(n2623), .S(n2037), .Y(N1181) );
  INVX2 U3320 ( .A(N1148), .Y(n2624) );
  MUX2X1 U3321 ( .B(n3140), .A(n2624), .S(n2037), .Y(N1180) );
  INVX2 U3322 ( .A(N1147), .Y(n2625) );
  MUX2X1 U3323 ( .B(n3141), .A(n2625), .S(n2037), .Y(N1179) );
  INVX2 U3324 ( .A(N1146), .Y(n2626) );
  MUX2X1 U3325 ( .B(n3142), .A(n2626), .S(n2037), .Y(N1178) );
  INVX2 U3326 ( .A(N1145), .Y(n2627) );
  MUX2X1 U3327 ( .B(n3143), .A(n2627), .S(n2037), .Y(N1177) );
  INVX2 U3328 ( .A(N1144), .Y(n2628) );
  MUX2X1 U3329 ( .B(n3144), .A(n2628), .S(n2037), .Y(N1176) );
  INVX2 U3330 ( .A(N1143), .Y(n2629) );
  MUX2X1 U3331 ( .B(n3145), .A(n2629), .S(n2037), .Y(N1175) );
  INVX2 U3332 ( .A(N1142), .Y(n2630) );
  MUX2X1 U3333 ( .B(n3146), .A(n2630), .S(n2037), .Y(N1174) );
  INVX2 U3334 ( .A(N1141), .Y(n2631) );
  MUX2X1 U3335 ( .B(n3147), .A(n2631), .S(n2037), .Y(N1173) );
  INVX2 U3336 ( .A(N1140), .Y(n2632) );
  MUX2X1 U3337 ( .B(n3148), .A(n2632), .S(n2037), .Y(N1172) );
  INVX2 U3338 ( .A(N1139), .Y(n2633) );
  MUX2X1 U3339 ( .B(n3149), .A(n2633), .S(n2037), .Y(N1171) );
  INVX2 U3340 ( .A(N1138), .Y(n2634) );
  MUX2X1 U3341 ( .B(n3150), .A(n2634), .S(n2037), .Y(N1170) );
  INVX2 U3342 ( .A(N1137), .Y(n2635) );
  MUX2X1 U3343 ( .B(n3151), .A(n2635), .S(n2037), .Y(N1169) );
  INVX2 U3344 ( .A(N1136), .Y(n2636) );
  MUX2X1 U3345 ( .B(n3152), .A(n2636), .S(n2037), .Y(N1168) );
  INVX2 U3346 ( .A(N1135), .Y(n2637) );
  MUX2X1 U3347 ( .B(n3153), .A(n2637), .S(n2037), .Y(N1167) );
  INVX2 U3348 ( .A(N1134), .Y(n2638) );
  MUX2X1 U3349 ( .B(n3154), .A(n2638), .S(n2037), .Y(N1166) );
  INVX2 U3350 ( .A(N1133), .Y(n2639) );
  MUX2X1 U3351 ( .B(n3155), .A(n2639), .S(n2037), .Y(N1165) );
  INVX2 U3352 ( .A(N1132), .Y(n2640) );
  MUX2X1 U3353 ( .B(n3156), .A(n2640), .S(n2037), .Y(N1164) );
  INVX2 U3354 ( .A(N1131), .Y(n2641) );
  MUX2X1 U3355 ( .B(n3157), .A(n2641), .S(n2037), .Y(N1163) );
  INVX2 U3356 ( .A(N1130), .Y(n2642) );
  MUX2X1 U3357 ( .B(n3158), .A(n2642), .S(n2037), .Y(N1162) );
  INVX2 U3358 ( .A(N1129), .Y(n2643) );
  MUX2X1 U3359 ( .B(n3159), .A(n2643), .S(n2037), .Y(N1161) );
  INVX2 U3360 ( .A(N1128), .Y(n2644) );
  MUX2X1 U3361 ( .B(n3160), .A(n2644), .S(n2037), .Y(N1160) );
  INVX2 U3362 ( .A(N1127), .Y(n2645) );
  MUX2X1 U3363 ( .B(n3161), .A(n2645), .S(n2037), .Y(N1159) );
  INVX2 U3364 ( .A(N1126), .Y(n2646) );
  MUX2X1 U3365 ( .B(n3162), .A(n2646), .S(n2037), .Y(N1158) );
  INVX2 U3366 ( .A(N1125), .Y(n2647) );
  MUX2X1 U3367 ( .B(n3163), .A(n2647), .S(n2037), .Y(N1157) );
  INVX2 U3368 ( .A(N1124), .Y(n2648) );
  MUX2X1 U3369 ( .B(n3164), .A(n2648), .S(n2037), .Y(N1156) );
  INVX2 U3370 ( .A(N1123), .Y(n2649) );
  MUX2X1 U3371 ( .B(n3165), .A(n2649), .S(n2037), .Y(N1155) );
  XNOR2X1 U3372 ( .A(n1904), .B(n2036), .Y(n2651) );
  MUX2X1 U3373 ( .B(N1087), .A(N1121), .S(n1919), .Y(n2714) );
  INVX2 U3374 ( .A(n2714), .Y(n3065) );
  MUX2X1 U3375 ( .B(N1086), .A(N1120), .S(n1919), .Y(n2653) );
  INVX2 U3376 ( .A(n2653), .Y(n2844) );
  MUX2X1 U3377 ( .B(N1085), .A(N1119), .S(n1919), .Y(n2655) );
  INVX2 U3378 ( .A(n2655), .Y(n2843) );
  MUX2X1 U3379 ( .B(n1883), .A(N1118), .S(n1919), .Y(n2657) );
  INVX2 U3380 ( .A(n2657), .Y(n2842) );
  MUX2X1 U3381 ( .B(N1083), .A(N1117), .S(n1919), .Y(n2659) );
  INVX2 U3382 ( .A(n2659), .Y(n2841) );
  MUX2X1 U3383 ( .B(N1082), .A(N1116), .S(n1919), .Y(n2661) );
  INVX2 U3384 ( .A(n2661), .Y(n2840) );
  MUX2X1 U3385 ( .B(N1081), .A(N1115), .S(n1919), .Y(n2663) );
  INVX2 U3386 ( .A(n2663), .Y(n2839) );
  MUX2X1 U3387 ( .B(N1080), .A(N1114), .S(n1919), .Y(n2665) );
  INVX2 U3388 ( .A(n2665), .Y(n2838) );
  MUX2X1 U3389 ( .B(N1079), .A(N1113), .S(n1919), .Y(n2667) );
  INVX2 U3390 ( .A(n2667), .Y(n2837) );
  MUX2X1 U3391 ( .B(N1078), .A(N1112), .S(n1919), .Y(n2669) );
  INVX2 U3392 ( .A(n2669), .Y(n2836) );
  MUX2X1 U3393 ( .B(N1077), .A(N1111), .S(n1919), .Y(n2671) );
  INVX2 U3394 ( .A(n2671), .Y(n2835) );
  MUX2X1 U3395 ( .B(N1076), .A(N1110), .S(n1919), .Y(n2673) );
  INVX2 U3396 ( .A(n2673), .Y(n2834) );
  MUX2X1 U3397 ( .B(N1075), .A(N1109), .S(n1919), .Y(n2675) );
  INVX2 U3398 ( .A(n2675), .Y(n2833) );
  MUX2X1 U3399 ( .B(N1074), .A(N1108), .S(n1919), .Y(n2677) );
  INVX2 U3400 ( .A(n2677), .Y(n2832) );
  MUX2X1 U3401 ( .B(n1844), .A(N1107), .S(n1919), .Y(n2679) );
  INVX2 U3402 ( .A(n2679), .Y(n2831) );
  MUX2X1 U3403 ( .B(N1072), .A(N1106), .S(n1919), .Y(n2681) );
  INVX2 U3404 ( .A(n2681), .Y(n2830) );
  MUX2X1 U3405 ( .B(N1071), .A(N1105), .S(n1919), .Y(n2683) );
  INVX2 U3406 ( .A(n2683), .Y(n2829) );
  MUX2X1 U3407 ( .B(N1070), .A(N1104), .S(n1919), .Y(n2685) );
  INVX2 U3408 ( .A(n2685), .Y(n2828) );
  MUX2X1 U3409 ( .B(N1069), .A(N1103), .S(n1919), .Y(n2687) );
  MUX2X1 U3410 ( .B(N1068), .A(N1102), .S(n1919), .Y(n2689) );
  INVX2 U3411 ( .A(n2689), .Y(n2826) );
  MUX2X1 U3412 ( .B(N1067), .A(N1101), .S(n1919), .Y(n2691) );
  INVX2 U3413 ( .A(n2691), .Y(n2825) );
  MUX2X1 U3414 ( .B(N1066), .A(N1100), .S(n1919), .Y(n2693) );
  INVX2 U3415 ( .A(n2693), .Y(n2824) );
  MUX2X1 U3416 ( .B(N1065), .A(N1099), .S(n1919), .Y(n2695) );
  INVX2 U3417 ( .A(n2695), .Y(n2823) );
  MUX2X1 U3418 ( .B(N1064), .A(N1098), .S(n1919), .Y(n2697) );
  INVX2 U3419 ( .A(n2697), .Y(n2822) );
  MUX2X1 U3420 ( .B(N1063), .A(N1097), .S(n1919), .Y(n2699) );
  INVX2 U3421 ( .A(n2699), .Y(n2821) );
  MUX2X1 U3422 ( .B(N1062), .A(N1096), .S(n1919), .Y(n2701) );
  INVX2 U3423 ( .A(n2701), .Y(n2820) );
  MUX2X1 U3424 ( .B(N1061), .A(N1095), .S(n1919), .Y(n2703) );
  INVX2 U3425 ( .A(n2703), .Y(n2819) );
  MUX2X1 U3426 ( .B(N1060), .A(N1094), .S(n1919), .Y(n2705) );
  INVX2 U3427 ( .A(n2705), .Y(n2818) );
  MUX2X1 U3428 ( .B(N1059), .A(N1093), .S(n1919), .Y(n2707) );
  INVX2 U3429 ( .A(n2707), .Y(n2817) );
  MUX2X1 U3430 ( .B(N1058), .A(N1092), .S(n1919), .Y(n2709) );
  INVX2 U3431 ( .A(n2709), .Y(n2816) );
  MUX2X1 U3432 ( .B(N1057), .A(N1091), .S(n1919), .Y(n2711) );
  INVX2 U3433 ( .A(n2711), .Y(n2815) );
  MUX2X1 U3434 ( .B(N1056), .A(N1090), .S(n1919), .Y(n2713) );
  INVX2 U3435 ( .A(n2713), .Y(n2814) );
  AND2X2 U3436 ( .A(N1219), .B(n1923), .Y(N1251) );
  INVX2 U3437 ( .A(N1218), .Y(n2652) );
  MUX2X1 U3438 ( .B(n2653), .A(n2652), .S(n1922), .Y(N1250) );
  INVX2 U3439 ( .A(N1217), .Y(n2654) );
  MUX2X1 U3440 ( .B(n2655), .A(n2654), .S(n1922), .Y(N1249) );
  INVX2 U3441 ( .A(N1216), .Y(n2656) );
  MUX2X1 U3442 ( .B(n2657), .A(n2656), .S(n1922), .Y(N1248) );
  INVX2 U3443 ( .A(N1215), .Y(n2658) );
  MUX2X1 U3444 ( .B(n2659), .A(n2658), .S(n1922), .Y(N1247) );
  MUX2X1 U3445 ( .B(n2661), .A(n2660), .S(n1922), .Y(N1246) );
  INVX2 U3446 ( .A(N1213), .Y(n2662) );
  MUX2X1 U3447 ( .B(n2663), .A(n2662), .S(n1922), .Y(N1245) );
  INVX2 U3448 ( .A(N1212), .Y(n2664) );
  MUX2X1 U3449 ( .B(n2665), .A(n2664), .S(n1922), .Y(N1244) );
  INVX2 U3450 ( .A(N1211), .Y(n2666) );
  MUX2X1 U3451 ( .B(n2667), .A(n2666), .S(n1922), .Y(N1243) );
  INVX2 U3452 ( .A(N1210), .Y(n2668) );
  MUX2X1 U3453 ( .B(n2669), .A(n2668), .S(n1922), .Y(N1242) );
  INVX2 U3454 ( .A(N1209), .Y(n2670) );
  MUX2X1 U3455 ( .B(n2671), .A(n2670), .S(n1922), .Y(N1241) );
  INVX2 U3456 ( .A(N1208), .Y(n2672) );
  MUX2X1 U3457 ( .B(n2673), .A(n2672), .S(n1922), .Y(N1240) );
  INVX2 U3458 ( .A(N1207), .Y(n2674) );
  MUX2X1 U3459 ( .B(n2675), .A(n2674), .S(n1922), .Y(N1239) );
  INVX2 U3460 ( .A(N1206), .Y(n2676) );
  MUX2X1 U3461 ( .B(n2677), .A(n2676), .S(n1922), .Y(N1238) );
  INVX2 U3462 ( .A(N1205), .Y(n2678) );
  MUX2X1 U3463 ( .B(n2679), .A(n2678), .S(n1922), .Y(N1237) );
  INVX2 U3464 ( .A(N1204), .Y(n2680) );
  MUX2X1 U3465 ( .B(n2681), .A(n2680), .S(n1922), .Y(N1236) );
  INVX2 U3466 ( .A(N1203), .Y(n2682) );
  MUX2X1 U3467 ( .B(n2683), .A(n2682), .S(n1922), .Y(N1235) );
  INVX2 U3468 ( .A(N1202), .Y(n2684) );
  MUX2X1 U3469 ( .B(n2685), .A(n2684), .S(n1922), .Y(N1234) );
  INVX2 U3470 ( .A(N1201), .Y(n2686) );
  MUX2X1 U3471 ( .B(n2687), .A(n2686), .S(n1922), .Y(N1233) );
  INVX2 U3472 ( .A(N1200), .Y(n2688) );
  MUX2X1 U3473 ( .B(n2689), .A(n2688), .S(n1923), .Y(N1232) );
  INVX2 U3474 ( .A(N1199), .Y(n2690) );
  MUX2X1 U3475 ( .B(n2691), .A(n2690), .S(n1923), .Y(N1231) );
  INVX2 U3476 ( .A(N1198), .Y(n2692) );
  MUX2X1 U3477 ( .B(n2693), .A(n2692), .S(n1923), .Y(N1230) );
  INVX2 U3478 ( .A(N1197), .Y(n2694) );
  MUX2X1 U3479 ( .B(n2695), .A(n2694), .S(n1923), .Y(N1229) );
  INVX2 U3480 ( .A(N1196), .Y(n2696) );
  MUX2X1 U3481 ( .B(n2697), .A(n2696), .S(n1923), .Y(N1228) );
  INVX2 U3482 ( .A(N1195), .Y(n2698) );
  MUX2X1 U3483 ( .B(n2699), .A(n2698), .S(n1923), .Y(N1227) );
  INVX2 U3484 ( .A(N1194), .Y(n2700) );
  MUX2X1 U3485 ( .B(n2701), .A(n2700), .S(n1923), .Y(N1226) );
  INVX2 U3486 ( .A(N1193), .Y(n2702) );
  MUX2X1 U3487 ( .B(n2703), .A(n2702), .S(n1923), .Y(N1225) );
  INVX2 U3488 ( .A(N1192), .Y(n2704) );
  MUX2X1 U3489 ( .B(n2705), .A(n2704), .S(n1923), .Y(N1224) );
  INVX2 U3490 ( .A(N1191), .Y(n2706) );
  MUX2X1 U3491 ( .B(n2707), .A(n2706), .S(n1923), .Y(N1223) );
  INVX2 U3492 ( .A(N1190), .Y(n2708) );
  MUX2X1 U3493 ( .B(n2709), .A(n2708), .S(n1923), .Y(N1222) );
  INVX2 U3494 ( .A(N1189), .Y(n2710) );
  MUX2X1 U3495 ( .B(n2711), .A(n2710), .S(n1923), .Y(N1221) );
  MUX2X1 U3496 ( .B(n2713), .A(n2712), .S(n1922), .Y(N1220) );
  INVX2 U3497 ( .A(N1299), .Y(n2717) );
  INVX2 U3498 ( .A(N1333), .Y(n2716) );
  XNOR2X1 U3499 ( .A(n2714), .B(n2038), .Y(n2715) );
  MUX2X1 U3500 ( .B(n2717), .A(n2716), .S(n1920), .Y(n2813) );
  INVX2 U3501 ( .A(N1298), .Y(n2719) );
  INVX2 U3502 ( .A(N1332), .Y(n2718) );
  MUX2X1 U3503 ( .B(n2719), .A(n2718), .S(n1920), .Y(n2812) );
  INVX2 U3504 ( .A(N1297), .Y(n2721) );
  INVX2 U3505 ( .A(N1331), .Y(n2720) );
  MUX2X1 U3506 ( .B(n2721), .A(n2720), .S(n1920), .Y(n2811) );
  INVX2 U3507 ( .A(N1296), .Y(n2723) );
  INVX2 U3508 ( .A(N1330), .Y(n2722) );
  MUX2X1 U3509 ( .B(n2723), .A(n2722), .S(n1920), .Y(n2810) );
  INVX2 U3510 ( .A(N1295), .Y(n2725) );
  INVX2 U3511 ( .A(N1329), .Y(n2724) );
  MUX2X1 U3512 ( .B(n2725), .A(n2724), .S(n1920), .Y(n2809) );
  INVX2 U3513 ( .A(N1294), .Y(n2727) );
  INVX2 U3514 ( .A(N1328), .Y(n2726) );
  MUX2X1 U3515 ( .B(n2727), .A(n2726), .S(n1920), .Y(n2808) );
  INVX2 U3516 ( .A(N1327), .Y(n2728) );
  MUX2X1 U3517 ( .B(n2729), .A(n2728), .S(n1920), .Y(n2807) );
  INVX2 U3518 ( .A(N1292), .Y(n2731) );
  INVX2 U3519 ( .A(N1326), .Y(n2730) );
  MUX2X1 U3520 ( .B(n2731), .A(n2730), .S(n1920), .Y(n2806) );
  INVX2 U3521 ( .A(N1291), .Y(n2733) );
  INVX2 U3522 ( .A(N1325), .Y(n2732) );
  MUX2X1 U3523 ( .B(n2733), .A(n2732), .S(n1920), .Y(n2805) );
  INVX2 U3524 ( .A(N1324), .Y(n2734) );
  MUX2X1 U3525 ( .B(n2735), .A(n2734), .S(n1920), .Y(n2804) );
  INVX2 U3526 ( .A(N1323), .Y(n2736) );
  MUX2X1 U3527 ( .B(n2737), .A(n2736), .S(n1920), .Y(n2803) );
  INVX2 U3528 ( .A(N1288), .Y(n2739) );
  INVX2 U3529 ( .A(N1322), .Y(n2738) );
  MUX2X1 U3530 ( .B(n2739), .A(n2738), .S(n1920), .Y(n2802) );
  INVX2 U3531 ( .A(N1287), .Y(n2741) );
  INVX2 U3532 ( .A(N1321), .Y(n2740) );
  MUX2X1 U3533 ( .B(n2741), .A(n2740), .S(n1920), .Y(n2801) );
  INVX2 U3534 ( .A(N1286), .Y(n2743) );
  MUX2X1 U3535 ( .B(n2743), .A(n2742), .S(n1920), .Y(n2800) );
  MUX2X1 U3536 ( .B(n2745), .A(n2744), .S(n1920), .Y(n2799) );
  INVX2 U3537 ( .A(N1284), .Y(n2747) );
  INVX2 U3538 ( .A(N1318), .Y(n2746) );
  MUX2X1 U3539 ( .B(n2747), .A(n2746), .S(n1920), .Y(n2798) );
  INVX2 U3540 ( .A(N1317), .Y(n2748) );
  MUX2X1 U3541 ( .B(n2749), .A(n2748), .S(n1920), .Y(n2797) );
  INVX2 U3542 ( .A(N1282), .Y(n2751) );
  INVX2 U3543 ( .A(N1316), .Y(n2750) );
  MUX2X1 U3544 ( .B(n2751), .A(n2750), .S(n1920), .Y(n2796) );
  INVX2 U3545 ( .A(N1281), .Y(n2753) );
  INVX2 U3546 ( .A(N1315), .Y(n2752) );
  MUX2X1 U3547 ( .B(n2753), .A(n2752), .S(n1920), .Y(n2795) );
  INVX2 U3548 ( .A(N1280), .Y(n2755) );
  INVX2 U3549 ( .A(N1314), .Y(n2754) );
  MUX2X1 U3550 ( .B(n2755), .A(n2754), .S(n1920), .Y(n2794) );
  INVX2 U3551 ( .A(N1313), .Y(n2756) );
  MUX2X1 U3552 ( .B(n2757), .A(n2756), .S(n1920), .Y(n2793) );
  INVX2 U3553 ( .A(N1278), .Y(n2759) );
  INVX2 U3554 ( .A(N1312), .Y(n2758) );
  MUX2X1 U3555 ( .B(n2759), .A(n2758), .S(n1920), .Y(n2792) );
  INVX2 U3556 ( .A(N1277), .Y(n2761) );
  INVX2 U3557 ( .A(N1311), .Y(n2760) );
  MUX2X1 U3558 ( .B(n2761), .A(n2760), .S(n1920), .Y(n2791) );
  INVX2 U3559 ( .A(N1276), .Y(n2763) );
  INVX2 U3560 ( .A(N1310), .Y(n2762) );
  MUX2X1 U3561 ( .B(n2763), .A(n2762), .S(n1920), .Y(n2790) );
  INVX2 U3562 ( .A(N1275), .Y(n2765) );
  INVX2 U3563 ( .A(N1309), .Y(n2764) );
  MUX2X1 U3564 ( .B(n2765), .A(n2764), .S(n1920), .Y(n2789) );
  INVX2 U3565 ( .A(N1274), .Y(n2767) );
  INVX2 U3566 ( .A(N1308), .Y(n2766) );
  MUX2X1 U3567 ( .B(n2767), .A(n2766), .S(n1920), .Y(n2788) );
  INVX2 U3568 ( .A(N1273), .Y(n2769) );
  INVX2 U3569 ( .A(N1307), .Y(n2768) );
  MUX2X1 U3570 ( .B(n2769), .A(n2768), .S(n1920), .Y(n2787) );
  INVX2 U3571 ( .A(N1272), .Y(n2771) );
  INVX2 U3572 ( .A(N1306), .Y(n2770) );
  MUX2X1 U3573 ( .B(n2771), .A(n2770), .S(n1920), .Y(n2786) );
  INVX2 U3574 ( .A(N1271), .Y(n2773) );
  INVX2 U3575 ( .A(N1305), .Y(n2772) );
  MUX2X1 U3576 ( .B(n2773), .A(n2772), .S(n1920), .Y(n2785) );
  INVX2 U3577 ( .A(N1270), .Y(n2775) );
  INVX2 U3578 ( .A(N1304), .Y(n2774) );
  MUX2X1 U3579 ( .B(n2775), .A(n2774), .S(n1920), .Y(n2784) );
  INVX2 U3580 ( .A(N1269), .Y(n2777) );
  INVX2 U3581 ( .A(N1303), .Y(n2776) );
  MUX2X1 U3582 ( .B(n2777), .A(n2776), .S(n1920), .Y(n2783) );
  INVX2 U3583 ( .A(N1268), .Y(n2779) );
  INVX2 U3584 ( .A(N1302), .Y(n2778) );
  MUX2X1 U3585 ( .B(n2779), .A(n2778), .S(n1920), .Y(n2782) );
  INVX2 U3586 ( .A(rst), .Y(n3068) );
  INVX2 U3587 ( .A(pushin), .Y(n3069) );
  INVX2 U3588 ( .A(opin[2]), .Y(n3070) );
  INVX2 U3589 ( .A(opin[0]), .Y(n3071) );
  INVX2 U3590 ( .A(datain[31]), .Y(n3072) );
  INVX2 U3591 ( .A(datain[30]), .Y(n3073) );
  INVX2 U3592 ( .A(datain[29]), .Y(n3074) );
  INVX2 U3593 ( .A(datain[28]), .Y(n3075) );
  INVX2 U3594 ( .A(datain[27]), .Y(n3076) );
  INVX2 U3595 ( .A(datain[26]), .Y(n3077) );
  INVX2 U3596 ( .A(datain[25]), .Y(n3078) );
  INVX2 U3597 ( .A(datain[24]), .Y(n3079) );
  INVX2 U3598 ( .A(datain[23]), .Y(n3080) );
  INVX2 U3599 ( .A(datain[22]), .Y(n3081) );
  INVX2 U3600 ( .A(datain[21]), .Y(n3082) );
  INVX2 U3601 ( .A(datain[20]), .Y(n3083) );
  INVX2 U3602 ( .A(datain[19]), .Y(n3084) );
  INVX2 U3603 ( .A(datain[18]), .Y(n3085) );
  INVX2 U3604 ( .A(datain[17]), .Y(n3086) );
  INVX2 U3605 ( .A(datain[16]), .Y(n3087) );
  INVX2 U3606 ( .A(datain[15]), .Y(n3088) );
  INVX2 U3607 ( .A(datain[14]), .Y(n3089) );
  INVX2 U3608 ( .A(datain[13]), .Y(n3090) );
  INVX2 U3609 ( .A(datain[12]), .Y(n3091) );
  INVX2 U3610 ( .A(datain[11]), .Y(n3092) );
  INVX2 U3611 ( .A(datain[10]), .Y(n3093) );
  INVX2 U3612 ( .A(datain[9]), .Y(n3094) );
  INVX2 U3613 ( .A(datain[8]), .Y(n3095) );
  INVX2 U3614 ( .A(datain[7]), .Y(n3096) );
  INVX2 U3615 ( .A(datain[6]), .Y(n3097) );
  INVX2 U3616 ( .A(datain[5]), .Y(n3098) );
  INVX2 U3617 ( .A(datain[4]), .Y(n3099) );
  INVX2 U3618 ( .A(datain[3]), .Y(n3100) );
  INVX2 U3619 ( .A(datain[2]), .Y(n3101) );
  INVX2 U3620 ( .A(datain[1]), .Y(n3102) );
  INVX2 U3621 ( .A(datain[0]), .Y(n3103) );
  INVX2 U3622 ( .A(a1[30]), .Y(n3166) );
  INVX2 U3623 ( .A(a1[29]), .Y(n3167) );
  INVX2 U3624 ( .A(a1[28]), .Y(n3168) );
  INVX2 U3625 ( .A(a1[27]), .Y(n3169) );
  INVX2 U3626 ( .A(a1[26]), .Y(n3170) );
  INVX2 U3627 ( .A(a1[25]), .Y(n3171) );
  INVX2 U3628 ( .A(a1[24]), .Y(n3172) );
  INVX2 U3629 ( .A(a1[23]), .Y(n3173) );
  INVX2 U3630 ( .A(a1[22]), .Y(n3174) );
  INVX2 U3631 ( .A(a1[21]), .Y(n3175) );
  INVX2 U3632 ( .A(a1[20]), .Y(n3176) );
  INVX2 U3633 ( .A(a1[19]), .Y(n3177) );
  INVX2 U3634 ( .A(a1[18]), .Y(n3178) );
  INVX2 U3635 ( .A(a1[17]), .Y(n3179) );
  INVX2 U3636 ( .A(a1[16]), .Y(n3180) );
  INVX2 U3637 ( .A(a1[15]), .Y(n3181) );
  INVX2 U3638 ( .A(a1[14]), .Y(n3182) );
  INVX2 U3639 ( .A(a1[13]), .Y(n3183) );
  INVX2 U3640 ( .A(a1[12]), .Y(n3184) );
  INVX2 U3641 ( .A(a1[11]), .Y(n3185) );
  INVX2 U3642 ( .A(a1[10]), .Y(n3186) );
  INVX2 U3643 ( .A(a1[9]), .Y(n3187) );
  INVX2 U3644 ( .A(a1[8]), .Y(n3188) );
  INVX2 U3645 ( .A(a1[7]), .Y(n3189) );
  INVX2 U3646 ( .A(a1[6]), .Y(n3190) );
  INVX2 U3647 ( .A(a1[5]), .Y(n3191) );
  INVX2 U3648 ( .A(a1[4]), .Y(n3192) );
  INVX2 U3649 ( .A(a1[3]), .Y(n3193) );
  INVX2 U3650 ( .A(a1[2]), .Y(n3194) );
  INVX2 U3651 ( .A(a1[1]), .Y(n3195) );
  INVX2 U3652 ( .A(a1[0]), .Y(n3196) );
endmodule

