
module sfilt_DW02_mult_3_stage_0 ( A, B, TC, CLK, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC, CLK;
  wire   n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695,
         \A_extended[32] , \B_extended[32] , \mult_97/n2953 , \mult_97/n2952 ,
         \mult_97/n2951 , \mult_97/n2950 , \mult_97/n2949 , \mult_97/n2948 ,
         \mult_97/n2947 , \mult_97/n2946 , \mult_97/n2945 , \mult_97/n2944 ,
         \mult_97/n2943 , \mult_97/n2942 , \mult_97/n2941 , \mult_97/n2940 ,
         \mult_97/n2939 , \mult_97/n2906 , \mult_97/n2905 , \mult_97/n2904 ,
         \mult_97/n2903 , \mult_97/n2902 , \mult_97/n2901 , \mult_97/n2900 ,
         \mult_97/n2899 , \mult_97/n2898 , \mult_97/n2897 , \mult_97/n2896 ,
         \mult_97/n2895 , \mult_97/n2894 , \mult_97/n2893 , \mult_97/n2892 ,
         \mult_97/n2891 , \mult_97/n2890 , \mult_97/n2889 , \mult_97/n2888 ,
         \mult_97/n2887 , \mult_97/n2886 , \mult_97/n2885 , \mult_97/n2884 ,
         \mult_97/n2883 , \mult_97/n2882 , \mult_97/n2881 , \mult_97/n2880 ,
         \mult_97/n2879 , \mult_97/n2878 , \mult_97/n2877 , \mult_97/n2876 ,
         \mult_97/n2875 , \mult_97/n2874 , \mult_97/n2873 , \mult_97/n2872 ,
         \mult_97/n2871 , \mult_97/n2870 , \mult_97/n2869 , \mult_97/n2868 ,
         \mult_97/n2867 , \mult_97/n2866 , \mult_97/n2865 , \mult_97/n2864 ,
         \mult_97/n2863 , \mult_97/n2862 , \mult_97/n2861 , \mult_97/n2860 ,
         \mult_97/n2859 , \mult_97/n2858 , \mult_97/n2857 , \mult_97/n2856 ,
         \mult_97/n2855 , \mult_97/n2854 , \mult_97/n2853 , \mult_97/n2852 ,
         \mult_97/n2851 , \mult_97/n2850 , \mult_97/n2849 , \mult_97/n2848 ,
         \mult_97/n2847 , \mult_97/n2846 , \mult_97/n2845 , \mult_97/n2844 ,
         \mult_97/n2843 , \mult_97/n2842 , \mult_97/n2841 , \mult_97/n2840 ,
         \mult_97/n2839 , \mult_97/n2838 , \mult_97/n2837 , \mult_97/n2836 ,
         \mult_97/n2835 , \mult_97/n2834 , \mult_97/n2833 , \mult_97/n2832 ,
         \mult_97/n2831 , \mult_97/n2830 , \mult_97/n2829 , \mult_97/n2828 ,
         \mult_97/n2827 , \mult_97/n2826 , \mult_97/n2825 , \mult_97/n2824 ,
         \mult_97/n2823 , \mult_97/n2822 , \mult_97/n2821 , \mult_97/n2820 ,
         \mult_97/n2819 , \mult_97/n2818 , \mult_97/n2817 , \mult_97/n2816 ,
         \mult_97/n2815 , \mult_97/n2814 , \mult_97/n2813 , \mult_97/n2812 ,
         \mult_97/n2811 , \mult_97/n2810 , \mult_97/n2809 , \mult_97/n2808 ,
         \mult_97/n2807 , \mult_97/n2806 , \mult_97/n2805 , \mult_97/n2804 ,
         \mult_97/n2803 , \mult_97/n2802 , \mult_97/n2801 , \mult_97/n2800 ,
         \mult_97/n2799 , \mult_97/n2798 , \mult_97/n2797 , \mult_97/n2796 ,
         \mult_97/n2795 , \mult_97/n2794 , \mult_97/n2793 , \mult_97/n2792 ,
         \mult_97/n2791 , \mult_97/n2790 , \mult_97/n2789 , \mult_97/n2788 ,
         \mult_97/n2787 , \mult_97/n2786 , \mult_97/n2785 , \mult_97/n2784 ,
         \mult_97/n2783 , \mult_97/n2782 , \mult_97/n2781 , \mult_97/n2780 ,
         \mult_97/n2779 , \mult_97/n2778 , \mult_97/n2777 , \mult_97/n2776 ,
         \mult_97/n2775 , \mult_97/n2774 , \mult_97/n2773 , \mult_97/n2772 ,
         \mult_97/n2771 , \mult_97/n2770 , \mult_97/n2769 , \mult_97/n2768 ,
         \mult_97/n2767 , \mult_97/n2766 , \mult_97/n2765 , \mult_97/n2764 ,
         \mult_97/n2763 , \mult_97/n2762 , \mult_97/n2761 , \mult_97/n2760 ,
         \mult_97/n2759 , \mult_97/n2758 , \mult_97/n2757 , \mult_97/n2756 ,
         \mult_97/n2755 , \mult_97/n2754 , \mult_97/n2753 , \mult_97/n2752 ,
         \mult_97/n2751 , \mult_97/n2750 , \mult_97/n2749 , \mult_97/n2748 ,
         \mult_97/n2747 , \mult_97/n2746 , \mult_97/n2745 , \mult_97/n2744 ,
         \mult_97/n2743 , \mult_97/n2742 , \mult_97/n2741 , \mult_97/n2740 ,
         \mult_97/n2739 , \mult_97/n2738 , \mult_97/n2737 , \mult_97/n2736 ,
         \mult_97/n2735 , \mult_97/n2734 , \mult_97/n2733 , \mult_97/n2732 ,
         \mult_97/n2731 , \mult_97/n2730 , \mult_97/n2729 , \mult_97/n2728 ,
         \mult_97/n2727 , \mult_97/n2726 , \mult_97/n2725 , \mult_97/n2724 ,
         \mult_97/n2723 , \mult_97/n2722 , \mult_97/n2721 , \mult_97/n2720 ,
         \mult_97/n2719 , \mult_97/n2718 , \mult_97/n2717 , \mult_97/n2716 ,
         \mult_97/n2715 , \mult_97/n2714 , \mult_97/n2713 , \mult_97/n2712 ,
         \mult_97/n2711 , \mult_97/n2710 , \mult_97/n2709 , \mult_97/n2708 ,
         \mult_97/n2707 , \mult_97/n2706 , \mult_97/n2705 , \mult_97/n2704 ,
         \mult_97/n2703 , \mult_97/n2702 , \mult_97/n2701 , \mult_97/n2700 ,
         \mult_97/n2699 , \mult_97/n2698 , \mult_97/n2697 , \mult_97/n2696 ,
         \mult_97/n2695 , \mult_97/n2694 , \mult_97/n2693 , \mult_97/n2692 ,
         \mult_97/n2691 , \mult_97/n2690 , \mult_97/n2689 , \mult_97/n2688 ,
         \mult_97/n2687 , \mult_97/n2686 , \mult_97/n2685 , \mult_97/n2684 ,
         \mult_97/n2683 , \mult_97/n2682 , \mult_97/n2681 , \mult_97/n2680 ,
         \mult_97/n2679 , \mult_97/n2678 , \mult_97/n2677 , \mult_97/n2676 ,
         \mult_97/n2675 , \mult_97/n2674 , \mult_97/n2673 , \mult_97/n2672 ,
         \mult_97/n2671 , \mult_97/n2670 , \mult_97/n2669 , \mult_97/n2668 ,
         \mult_97/n2667 , \mult_97/n2666 , \mult_97/n2665 , \mult_97/n2664 ,
         \mult_97/n2663 , \mult_97/n2662 , \mult_97/n2661 , \mult_97/n2660 ,
         \mult_97/n2659 , \mult_97/n2658 , \mult_97/n2657 , \mult_97/n2656 ,
         \mult_97/n2655 , \mult_97/n2654 , \mult_97/n2653 , \mult_97/n2652 ,
         \mult_97/n2651 , \mult_97/n2650 , \mult_97/n2649 , \mult_97/n2648 ,
         \mult_97/n2647 , \mult_97/n2646 , \mult_97/n2645 , \mult_97/n2644 ,
         \mult_97/n2643 , \mult_97/n2642 , \mult_97/n2641 , \mult_97/n2640 ,
         \mult_97/n2639 , \mult_97/n2638 , \mult_97/n2637 , \mult_97/n2636 ,
         \mult_97/n2635 , \mult_97/n2634 , \mult_97/n2633 , \mult_97/n2632 ,
         \mult_97/n2631 , \mult_97/n2630 , \mult_97/n2629 , \mult_97/n2628 ,
         \mult_97/n2627 , \mult_97/n2626 , \mult_97/n2625 , \mult_97/n2624 ,
         \mult_97/n2623 , \mult_97/n2622 , \mult_97/n2621 , \mult_97/n2620 ,
         \mult_97/n2619 , \mult_97/n2618 , \mult_97/n2617 , \mult_97/n2616 ,
         \mult_97/n2615 , \mult_97/n2614 , \mult_97/n2613 , \mult_97/n2612 ,
         \mult_97/n2611 , \mult_97/n2610 , \mult_97/n2609 , \mult_97/n2608 ,
         \mult_97/n2607 , \mult_97/n2606 , \mult_97/n2605 , \mult_97/n2604 ,
         \mult_97/n2603 , \mult_97/n2602 , \mult_97/n2601 , \mult_97/n2600 ,
         \mult_97/n2599 , \mult_97/n2598 , \mult_97/n2597 , \mult_97/n2596 ,
         \mult_97/n2595 , \mult_97/n2594 , \mult_97/n2593 , \mult_97/n2592 ,
         \mult_97/n2591 , \mult_97/n2590 , \mult_97/n2589 , \mult_97/n2588 ,
         \mult_97/n2587 , \mult_97/n2586 , \mult_97/n2585 , \mult_97/n2584 ,
         \mult_97/n2583 , \mult_97/n2582 , \mult_97/n2581 , \mult_97/n2580 ,
         \mult_97/n2579 , \mult_97/n2578 , \mult_97/n2577 , \mult_97/n2576 ,
         \mult_97/n2575 , \mult_97/n2574 , \mult_97/n2573 , \mult_97/n2572 ,
         \mult_97/n2571 , \mult_97/n2570 , \mult_97/n2569 , \mult_97/n2568 ,
         \mult_97/n2567 , \mult_97/n2566 , \mult_97/n2565 , \mult_97/n2564 ,
         \mult_97/n2563 , \mult_97/n2562 , \mult_97/n2561 , \mult_97/n2560 ,
         \mult_97/n2559 , \mult_97/n2558 , \mult_97/n2557 , \mult_97/n2556 ,
         \mult_97/n2555 , \mult_97/n2554 , \mult_97/n2553 , \mult_97/n2552 ,
         \mult_97/n2551 , \mult_97/n2550 , \mult_97/n2549 , \mult_97/n2548 ,
         \mult_97/n2547 , \mult_97/n2546 , \mult_97/n2545 , \mult_97/n2544 ,
         \mult_97/n2543 , \mult_97/n2542 , \mult_97/n2541 , \mult_97/n2540 ,
         \mult_97/n2539 , \mult_97/n2538 , \mult_97/n2537 , \mult_97/n2536 ,
         \mult_97/n2535 , \mult_97/n2534 , \mult_97/n2533 , \mult_97/n2532 ,
         \mult_97/n2531 , \mult_97/n2530 , \mult_97/n2529 , \mult_97/n2528 ,
         \mult_97/n2527 , \mult_97/n2526 , \mult_97/n2525 , \mult_97/n2524 ,
         \mult_97/n2523 , \mult_97/n2522 , \mult_97/n2521 , \mult_97/n2520 ,
         \mult_97/n2519 , \mult_97/n2518 , \mult_97/n2517 , \mult_97/n2516 ,
         \mult_97/n2515 , \mult_97/n2514 , \mult_97/n2513 , \mult_97/n2512 ,
         \mult_97/n2511 , \mult_97/n2510 , \mult_97/n2509 , \mult_97/n2508 ,
         \mult_97/n2507 , \mult_97/n2506 , \mult_97/n2505 , \mult_97/n2504 ,
         \mult_97/n2503 , \mult_97/n2502 , \mult_97/n2501 , \mult_97/n2500 ,
         \mult_97/n2499 , \mult_97/n2498 , \mult_97/n2497 , \mult_97/n2496 ,
         \mult_97/n2495 , \mult_97/n2494 , \mult_97/n2493 , \mult_97/n2492 ,
         \mult_97/n2491 , \mult_97/n2490 , \mult_97/n2489 , \mult_97/n2488 ,
         \mult_97/n2487 , \mult_97/n2486 , \mult_97/n2485 , \mult_97/n2484 ,
         \mult_97/n2483 , \mult_97/n2482 , \mult_97/n2481 , \mult_97/n2480 ,
         \mult_97/n2479 , \mult_97/n2478 , \mult_97/n2477 , \mult_97/n2476 ,
         \mult_97/n2475 , \mult_97/n2474 , \mult_97/n2473 , \mult_97/n2472 ,
         \mult_97/n2471 , \mult_97/n2470 , \mult_97/n2469 , \mult_97/n2468 ,
         \mult_97/n2467 , \mult_97/n2466 , \mult_97/n2465 , \mult_97/n2464 ,
         \mult_97/n2463 , \mult_97/n2462 , \mult_97/n2461 , \mult_97/n2460 ,
         \mult_97/n2459 , \mult_97/n2458 , \mult_97/n2457 , \mult_97/n2456 ,
         \mult_97/n2455 , \mult_97/n2454 , \mult_97/n2453 , \mult_97/n2452 ,
         \mult_97/n2451 , \mult_97/n2450 , \mult_97/n2449 , \mult_97/n2448 ,
         \mult_97/n2447 , \mult_97/n2446 , \mult_97/n2445 , \mult_97/n2444 ,
         \mult_97/n2443 , \mult_97/n2442 , \mult_97/n2441 , \mult_97/n2440 ,
         \mult_97/n2439 , \mult_97/n2438 , \mult_97/n2437 , \mult_97/n2436 ,
         \mult_97/n2435 , \mult_97/n2434 , \mult_97/n2433 , \mult_97/n2432 ,
         \mult_97/n2431 , \mult_97/n2430 , \mult_97/n2429 , \mult_97/n2428 ,
         \mult_97/n2427 , \mult_97/n2426 , \mult_97/n2425 , \mult_97/n2424 ,
         \mult_97/n2423 , \mult_97/n2422 , \mult_97/n2421 , \mult_97/n2420 ,
         \mult_97/n2419 , \mult_97/n2418 , \mult_97/n2417 , \mult_97/n2416 ,
         \mult_97/n2415 , \mult_97/n2414 , \mult_97/n2413 , \mult_97/n2412 ,
         \mult_97/n2411 , \mult_97/n2410 , \mult_97/n2409 , \mult_97/n2408 ,
         \mult_97/n2407 , \mult_97/n2406 , \mult_97/n2405 , \mult_97/n2404 ,
         \mult_97/n2403 , \mult_97/n2402 , \mult_97/n2401 , \mult_97/n2400 ,
         \mult_97/n2399 , \mult_97/n2398 , \mult_97/n2397 , \mult_97/n2396 ,
         \mult_97/n2395 , \mult_97/n2394 , \mult_97/n2393 , \mult_97/n2392 ,
         \mult_97/n2391 , \mult_97/n2390 , \mult_97/n2389 , \mult_97/n2388 ,
         \mult_97/n2387 , \mult_97/n2386 , \mult_97/n2385 , \mult_97/n2384 ,
         \mult_97/n2383 , \mult_97/n2382 , \mult_97/n2381 , \mult_97/n2380 ,
         \mult_97/n2379 , \mult_97/n2378 , \mult_97/n2377 , \mult_97/n2376 ,
         \mult_97/n2375 , \mult_97/n2374 , \mult_97/n2373 , \mult_97/n2372 ,
         \mult_97/n2371 , \mult_97/n2370 , \mult_97/n2369 , \mult_97/n2368 ,
         \mult_97/n2367 , \mult_97/n2366 , \mult_97/n2365 , \mult_97/n2364 ,
         \mult_97/n2363 , \mult_97/n2362 , \mult_97/n2361 , \mult_97/n2360 ,
         \mult_97/n2359 , \mult_97/n2358 , \mult_97/n2357 , \mult_97/n2356 ,
         \mult_97/n2355 , \mult_97/n2354 , \mult_97/n2353 , \mult_97/n2352 ,
         \mult_97/n2351 , \mult_97/n2350 , \mult_97/n2349 , \mult_97/n2348 ,
         \mult_97/n2347 , \mult_97/n2346 , \mult_97/n2345 , \mult_97/n2344 ,
         \mult_97/n2343 , \mult_97/n2342 , \mult_97/n2341 , \mult_97/n2340 ,
         \mult_97/n2339 , \mult_97/n2338 , \mult_97/n2337 , \mult_97/n2336 ,
         \mult_97/n2335 , \mult_97/n2334 , \mult_97/n2333 , \mult_97/n2332 ,
         \mult_97/n2331 , \mult_97/n2330 , \mult_97/n2329 , \mult_97/n2328 ,
         \mult_97/n2327 , \mult_97/n2326 , \mult_97/n2325 , \mult_97/n2324 ,
         \mult_97/n2323 , \mult_97/n2322 , \mult_97/n2321 , \mult_97/n2320 ,
         \mult_97/n2319 , \mult_97/n2318 , \mult_97/n2317 , \mult_97/n2316 ,
         \mult_97/n2315 , \mult_97/n2314 , \mult_97/n2313 , \mult_97/n2312 ,
         \mult_97/n2311 , \mult_97/n2310 , \mult_97/n2309 , \mult_97/n2308 ,
         \mult_97/n2307 , \mult_97/n2306 , \mult_97/n2305 , \mult_97/n2304 ,
         \mult_97/n2303 , \mult_97/n2302 , \mult_97/n2301 , \mult_97/n2300 ,
         \mult_97/n2299 , \mult_97/n2298 , \mult_97/n2297 , \mult_97/n2296 ,
         \mult_97/n2295 , \mult_97/n2294 , \mult_97/n2293 , \mult_97/n2292 ,
         \mult_97/n2291 , \mult_97/n2290 , \mult_97/n2289 , \mult_97/n2288 ,
         \mult_97/n2287 , \mult_97/n2286 , \mult_97/n2285 , \mult_97/n2284 ,
         \mult_97/n2283 , \mult_97/n2282 , \mult_97/n2281 , \mult_97/n2280 ,
         \mult_97/n2279 , \mult_97/n2278 , \mult_97/n2277 , \mult_97/n2276 ,
         \mult_97/n2275 , \mult_97/n2274 , \mult_97/n2273 , \mult_97/n2272 ,
         \mult_97/n2271 , \mult_97/n2270 , \mult_97/n2269 , \mult_97/n2268 ,
         \mult_97/n2267 , \mult_97/n2266 , \mult_97/n2265 , \mult_97/n2264 ,
         \mult_97/n2263 , \mult_97/n2262 , \mult_97/n2261 , \mult_97/n2260 ,
         \mult_97/n2259 , \mult_97/n2258 , \mult_97/n2257 , \mult_97/n2256 ,
         \mult_97/n2255 , \mult_97/n2254 , \mult_97/n2253 , \mult_97/n2252 ,
         \mult_97/n2251 , \mult_97/n2250 , \mult_97/n2249 , \mult_97/n2248 ,
         \mult_97/n2247 , \mult_97/n2246 , \mult_97/n2245 , \mult_97/n2244 ,
         \mult_97/n2243 , \mult_97/n2242 , \mult_97/n2241 , \mult_97/n2240 ,
         \mult_97/n2239 , \mult_97/n2238 , \mult_97/n2237 , \mult_97/n2236 ,
         \mult_97/n2235 , \mult_97/n2234 , \mult_97/n2233 , \mult_97/n2232 ,
         \mult_97/n2231 , \mult_97/n2230 , \mult_97/n2229 , \mult_97/n2228 ,
         \mult_97/n2227 , \mult_97/n2226 , \mult_97/n2225 , \mult_97/n2224 ,
         \mult_97/n2223 , \mult_97/n2222 , \mult_97/n2221 , \mult_97/n2220 ,
         \mult_97/n2219 , \mult_97/n2218 , \mult_97/n2217 , \mult_97/n2216 ,
         \mult_97/n2215 , \mult_97/n2214 , \mult_97/n2213 , \mult_97/n2212 ,
         \mult_97/n2211 , \mult_97/n2210 , \mult_97/n2209 , \mult_97/n2208 ,
         \mult_97/n2207 , \mult_97/n2206 , \mult_97/n2205 , \mult_97/n2204 ,
         \mult_97/n2203 , \mult_97/n2202 , \mult_97/n2201 , \mult_97/n2200 ,
         \mult_97/n2199 , \mult_97/n2198 , \mult_97/n2197 , \mult_97/n2196 ,
         \mult_97/n2195 , \mult_97/n2194 , \mult_97/n2193 , \mult_97/n2192 ,
         \mult_97/n2191 , \mult_97/n2190 , \mult_97/n2189 , \mult_97/n2188 ,
         \mult_97/n2187 , \mult_97/n2186 , \mult_97/n2185 , \mult_97/n2184 ,
         \mult_97/n2183 , \mult_97/n2182 , \mult_97/n2181 , \mult_97/n2180 ,
         \mult_97/n2179 , \mult_97/n2178 , \mult_97/n2177 , \mult_97/n2176 ,
         \mult_97/n2175 , \mult_97/n2174 , \mult_97/n2173 , \mult_97/n2172 ,
         \mult_97/n2171 , \mult_97/n2170 , \mult_97/n2169 , \mult_97/n2168 ,
         \mult_97/n2167 , \mult_97/n2166 , \mult_97/n2165 , \mult_97/n2164 ,
         \mult_97/n2163 , \mult_97/n2162 , \mult_97/n2161 , \mult_97/n2160 ,
         \mult_97/n2159 , \mult_97/n2158 , \mult_97/n2157 , \mult_97/n2156 ,
         \mult_97/n2155 , \mult_97/n2154 , \mult_97/n2153 , \mult_97/n2152 ,
         \mult_97/n2151 , \mult_97/n2150 , \mult_97/n2149 , \mult_97/n2148 ,
         \mult_97/n2147 , \mult_97/n2146 , \mult_97/n2145 , \mult_97/n2144 ,
         \mult_97/n2143 , \mult_97/n2142 , \mult_97/n2141 , \mult_97/n2140 ,
         \mult_97/n2139 , \mult_97/n2138 , \mult_97/n2137 , \mult_97/n2136 ,
         \mult_97/n2135 , \mult_97/n2134 , \mult_97/n2133 , \mult_97/n2132 ,
         \mult_97/n2131 , \mult_97/n2130 , \mult_97/n2129 , \mult_97/n2128 ,
         \mult_97/n2127 , \mult_97/n2126 , \mult_97/n2125 , \mult_97/n2124 ,
         \mult_97/n2123 , \mult_97/n2122 , \mult_97/n2121 , \mult_97/n2120 ,
         \mult_97/n2119 , \mult_97/n2118 , \mult_97/n2117 , \mult_97/n2116 ,
         \mult_97/n2115 , \mult_97/n2114 , \mult_97/n2113 , \mult_97/n2112 ,
         \mult_97/n2111 , \mult_97/n2110 , \mult_97/n2109 , \mult_97/n2108 ,
         \mult_97/n2107 , \mult_97/n2106 , \mult_97/n2105 , \mult_97/n2104 ,
         \mult_97/n2103 , \mult_97/n2102 , \mult_97/n2101 , \mult_97/n2100 ,
         \mult_97/n2099 , \mult_97/n2098 , \mult_97/n2097 , \mult_97/n2096 ,
         \mult_97/n2095 , \mult_97/n2094 , \mult_97/n2093 , \mult_97/n2092 ,
         \mult_97/n2091 , \mult_97/n2090 , \mult_97/n2089 , \mult_97/n2088 ,
         \mult_97/n2087 , \mult_97/n2086 , \mult_97/n2085 , \mult_97/n2084 ,
         \mult_97/n2083 , \mult_97/n2082 , \mult_97/n2081 , \mult_97/n2080 ,
         \mult_97/n2079 , \mult_97/n2078 , \mult_97/n2077 , \mult_97/n2076 ,
         \mult_97/n2075 , \mult_97/n2074 , \mult_97/n2073 , \mult_97/n2072 ,
         \mult_97/n2071 , \mult_97/n2070 , \mult_97/n2069 , \mult_97/n2068 ,
         \mult_97/n2067 , \mult_97/n2066 , \mult_97/n2065 , \mult_97/n2064 ,
         \mult_97/n2063 , \mult_97/n2062 , \mult_97/n2061 , \mult_97/n2060 ,
         \mult_97/n2059 , \mult_97/n2058 , \mult_97/n2057 , \mult_97/n2056 ,
         \mult_97/n2055 , \mult_97/n2054 , \mult_97/n2053 , \mult_97/n2052 ,
         \mult_97/n2051 , \mult_97/n2050 , \mult_97/n2049 , \mult_97/n2048 ,
         \mult_97/n2047 , \mult_97/n2046 , \mult_97/n2045 , \mult_97/n2044 ,
         \mult_97/n2043 , \mult_97/n2042 , \mult_97/n2041 , \mult_97/n2040 ,
         \mult_97/n2039 , \mult_97/n2038 , \mult_97/n2037 , \mult_97/n2036 ,
         \mult_97/n2035 , \mult_97/n2034 , \mult_97/n2033 , \mult_97/n2032 ,
         \mult_97/n2031 , \mult_97/n2030 , \mult_97/n2029 , \mult_97/n2028 ,
         \mult_97/n2027 , \mult_97/n2026 , \mult_97/n2025 , \mult_97/n2024 ,
         \mult_97/n2023 , \mult_97/n2022 , \mult_97/n2021 , \mult_97/n2020 ,
         \mult_97/n2019 , \mult_97/n2018 , \mult_97/n2017 , \mult_97/n2016 ,
         \mult_97/n2015 , \mult_97/n2014 , \mult_97/n2013 , \mult_97/n2012 ,
         \mult_97/n2011 , \mult_97/n2010 , \mult_97/n2009 , \mult_97/n2008 ,
         \mult_97/n2007 , \mult_97/n2006 , \mult_97/n2005 , \mult_97/n2004 ,
         \mult_97/n2003 , \mult_97/n2002 , \mult_97/n2001 , \mult_97/n2000 ,
         \mult_97/n1999 , \mult_97/n1998 , \mult_97/n1997 , \mult_97/n1996 ,
         \mult_97/n1995 , \mult_97/n1994 , \mult_97/n1993 , \mult_97/n1992 ,
         \mult_97/n1991 , \mult_97/n1990 , \mult_97/n1989 , \mult_97/n1988 ,
         \mult_97/n1987 , \mult_97/n1986 , \mult_97/n1985 , \mult_97/n1984 ,
         \mult_97/n1983 , \mult_97/n1982 , \mult_97/n1981 , \mult_97/n1980 ,
         \mult_97/n1979 , \mult_97/n1978 , \mult_97/n1977 , \mult_97/n1976 ,
         \mult_97/n1975 , \mult_97/n1974 , \mult_97/n1973 , \mult_97/n1972 ,
         \mult_97/n1971 , \mult_97/n1970 , \mult_97/n1969 , \mult_97/n1968 ,
         \mult_97/n1967 , \mult_97/n1966 , \mult_97/n1965 , \mult_97/n1964 ,
         \mult_97/n1963 , \mult_97/n1962 , \mult_97/n1961 , \mult_97/n1960 ,
         \mult_97/n1959 , \mult_97/n1958 , \mult_97/n1957 , \mult_97/n1956 ,
         \mult_97/n1955 , \mult_97/n1954 , \mult_97/n1953 , \mult_97/n1952 ,
         \mult_97/n1951 , \mult_97/n1950 , \mult_97/n1949 , \mult_97/n1948 ,
         \mult_97/n1947 , \mult_97/n1946 , \mult_97/n1945 , \mult_97/n1944 ,
         \mult_97/n1943 , \mult_97/n1942 , \mult_97/n1941 , \mult_97/n1940 ,
         \mult_97/n1939 , \mult_97/n1938 , \mult_97/n1937 , \mult_97/n1936 ,
         \mult_97/n1935 , \mult_97/n1934 , \mult_97/n1933 , \mult_97/n1932 ,
         \mult_97/n1931 , \mult_97/n1930 , \mult_97/n1929 , \mult_97/n1928 ,
         \mult_97/n1927 , \mult_97/n1926 , \mult_97/n1925 , \mult_97/n1924 ,
         \mult_97/n1923 , \mult_97/n1922 , \mult_97/n1921 , \mult_97/n1920 ,
         \mult_97/n1919 , \mult_97/n1918 , \mult_97/n1917 , \mult_97/n1916 ,
         \mult_97/n1915 , \mult_97/n1914 , \mult_97/n1913 , \mult_97/n1912 ,
         \mult_97/n1911 , \mult_97/n1910 , \mult_97/n1909 , \mult_97/n1908 ,
         \mult_97/n1907 , \mult_97/n1906 , \mult_97/n1905 , \mult_97/n1904 ,
         \mult_97/n1903 , \mult_97/n1902 , \mult_97/n1901 , \mult_97/n1900 ,
         \mult_97/n1899 , \mult_97/n1898 , \mult_97/n1897 , \mult_97/n1896 ,
         \mult_97/n1895 , \mult_97/n1894 , \mult_97/n1893 , \mult_97/n1892 ,
         \mult_97/n1891 , \mult_97/n1890 , \mult_97/n1889 , \mult_97/n1888 ,
         \mult_97/n1887 , \mult_97/n1886 , \mult_97/n1885 , \mult_97/n1884 ,
         \mult_97/n1883 , \mult_97/n1882 , \mult_97/n1881 , \mult_97/n1880 ,
         \mult_97/n1879 , \mult_97/n1878 , \mult_97/n1877 , \mult_97/n1876 ,
         \mult_97/n1875 , \mult_97/n1874 , \mult_97/n1873 , \mult_97/n1872 ,
         \mult_97/n1871 , \mult_97/n1870 , \mult_97/n1869 , \mult_97/n1868 ,
         \mult_97/n1867 , \mult_97/n1866 , \mult_97/n1865 , \mult_97/n1864 ,
         \mult_97/n1863 , \mult_97/n1862 , \mult_97/n1861 , \mult_97/n1860 ,
         \mult_97/n1859 , \mult_97/n1858 , \mult_97/n1857 , \mult_97/n1856 ,
         \mult_97/n1855 , \mult_97/n1854 , \mult_97/n1853 , \mult_97/n1852 ,
         \mult_97/n1851 , \mult_97/n1850 , \mult_97/n1849 , \mult_97/n1848 ,
         \mult_97/n1847 , \mult_97/n1846 , \mult_97/n1845 , \mult_97/n1844 ,
         \mult_97/n1843 , \mult_97/n1842 , \mult_97/n1841 , \mult_97/n1840 ,
         \mult_97/n1839 , \mult_97/n1838 , \mult_97/n1837 , \mult_97/n1836 ,
         \mult_97/n1835 , \mult_97/n1834 , \mult_97/n1833 , \mult_97/n1832 ,
         \mult_97/n1831 , \mult_97/n1830 , \mult_97/n1829 , \mult_97/n1828 ,
         \mult_97/n1827 , \mult_97/n1826 , \mult_97/n1825 , \mult_97/n1824 ,
         \mult_97/n1823 , \mult_97/n1822 , \mult_97/n1821 , \mult_97/n1820 ,
         \mult_97/n1819 , \mult_97/n1818 , \mult_97/n1817 , \mult_97/n1816 ,
         \mult_97/n1815 , \mult_97/n1814 , \mult_97/n1813 , \mult_97/n1812 ,
         \mult_97/n1811 , \mult_97/n1810 , \mult_97/n1809 , \mult_97/n1808 ,
         \mult_97/n1807 , \mult_97/n1806 , \mult_97/n1805 , \mult_97/n1804 ,
         \mult_97/n1803 , \mult_97/n1802 , \mult_97/n1801 , \mult_97/n1800 ,
         \mult_97/n1799 , \mult_97/n1798 , \mult_97/n1797 , \mult_97/n1796 ,
         \mult_97/n1795 , \mult_97/n1794 , \mult_97/n1793 , \mult_97/n1792 ,
         \mult_97/n1791 , \mult_97/n1790 , \mult_97/n1789 , \mult_97/n1788 ,
         \mult_97/n1787 , \mult_97/n1786 , \mult_97/n1785 , \mult_97/n1784 ,
         \mult_97/n1783 , \mult_97/n1782 , \mult_97/n1781 , \mult_97/n1780 ,
         \mult_97/n1779 , \mult_97/n1778 , \mult_97/n1777 , \mult_97/n1776 ,
         \mult_97/n1775 , \mult_97/n1774 , \mult_97/n1773 , \mult_97/n1772 ,
         \mult_97/n1771 , \mult_97/n1770 , \mult_97/n1769 , \mult_97/n1768 ,
         \mult_97/n1767 , \mult_97/n1766 , \mult_97/n1765 , \mult_97/n1764 ,
         \mult_97/n1763 , \mult_97/n1762 , \mult_97/n1761 , \mult_97/n1760 ,
         \mult_97/n1759 , \mult_97/n1758 , \mult_97/n1757 , \mult_97/n1756 ,
         \mult_97/n1755 , \mult_97/n1754 , \mult_97/n1753 , \mult_97/n1752 ,
         \mult_97/n1751 , \mult_97/n1750 , \mult_97/n1749 , \mult_97/n1748 ,
         \mult_97/n1747 , \mult_97/n1746 , \mult_97/n1745 , \mult_97/n1744 ,
         \mult_97/n1743 , \mult_97/n1742 , \mult_97/n1741 , \mult_97/n1740 ,
         \mult_97/n1739 , \mult_97/n1738 , \mult_97/n1737 , \mult_97/n1736 ,
         \mult_97/n1735 , \mult_97/n1734 , \mult_97/n1733 , \mult_97/n1732 ,
         \mult_97/n1731 , \mult_97/n1730 , \mult_97/n1729 , \mult_97/n1728 ,
         \mult_97/n1727 , \mult_97/n1726 , \mult_97/n1725 , \mult_97/n1724 ,
         \mult_97/n1723 , \mult_97/n1722 , \mult_97/n1721 , \mult_97/n1720 ,
         \mult_97/n1719 , \mult_97/n1718 , \mult_97/n1717 , \mult_97/n1716 ,
         \mult_97/n1715 , \mult_97/n1714 , \mult_97/n1713 , \mult_97/n1712 ,
         \mult_97/n1711 , \mult_97/n1710 , \mult_97/n1709 , \mult_97/n1708 ,
         \mult_97/n1707 , \mult_97/n1706 , \mult_97/n1705 , \mult_97/n1704 ,
         \mult_97/n1703 , \mult_97/n1702 , \mult_97/n1701 , \mult_97/n1700 ,
         \mult_97/n1699 , \mult_97/n1698 , \mult_97/n1697 , \mult_97/n1696 ,
         \mult_97/n1695 , \mult_97/n1694 , \mult_97/n1693 , \mult_97/n1692 ,
         \mult_97/n1691 , \mult_97/n1690 , \mult_97/n1689 , \mult_97/n1688 ,
         \mult_97/n1687 , \mult_97/n1686 , \mult_97/n1685 , \mult_97/n1684 ,
         \mult_97/n1683 , \mult_97/n1682 , \mult_97/n1681 , \mult_97/n1680 ,
         \mult_97/n1679 , \mult_97/n1678 , \mult_97/n1677 , \mult_97/n1676 ,
         \mult_97/n1675 , \mult_97/n1674 , \mult_97/n1673 , \mult_97/n1672 ,
         \mult_97/n1671 , \mult_97/n1670 , \mult_97/n1669 , \mult_97/n1668 ,
         \mult_97/n1667 , \mult_97/n1666 , \mult_97/n1665 , \mult_97/n1664 ,
         \mult_97/n1663 , \mult_97/n1662 , \mult_97/n1661 , \mult_97/n1660 ,
         \mult_97/n1659 , \mult_97/n1658 , \mult_97/n1657 , \mult_97/n1656 ,
         \mult_97/n1655 , \mult_97/n1654 , \mult_97/n1653 , \mult_97/n1652 ,
         \mult_97/n1651 , \mult_97/n1650 , \mult_97/n1649 , \mult_97/n1648 ,
         \mult_97/n1647 , \mult_97/n1646 , \mult_97/n1645 , \mult_97/n1644 ,
         \mult_97/n1643 , \mult_97/n1642 , \mult_97/n1641 , \mult_97/n1640 ,
         \mult_97/n1639 , \mult_97/n1638 , \mult_97/n1637 , \mult_97/n1636 ,
         \mult_97/n1635 , \mult_97/n1634 , \mult_97/n1633 , \mult_97/n1632 ,
         \mult_97/n1631 , \mult_97/n1630 , \mult_97/n1629 , \mult_97/n1628 ,
         \mult_97/n1627 , \mult_97/n1626 , \mult_97/n1625 , \mult_97/n1624 ,
         \mult_97/n1623 , \mult_97/n1622 , \mult_97/n1621 , \mult_97/n1620 ,
         \mult_97/n1619 , \mult_97/n1618 , \mult_97/n1617 , \mult_97/n1616 ,
         \mult_97/n1615 , \mult_97/n1614 , \mult_97/n1613 , \mult_97/n1612 ,
         \mult_97/n1611 , \mult_97/n1610 , \mult_97/n1609 , \mult_97/n1608 ,
         \mult_97/n1607 , \mult_97/n1606 , \mult_97/n1605 , \mult_97/n1604 ,
         \mult_97/n1603 , \mult_97/n1602 , \mult_97/n1601 , \mult_97/n1600 ,
         \mult_97/n1599 , \mult_97/n1598 , \mult_97/n1597 , \mult_97/n1596 ,
         \mult_97/n1595 , \mult_97/n1594 , \mult_97/n1593 , \mult_97/n1592 ,
         \mult_97/n1591 , \mult_97/n1590 , \mult_97/n1589 , \mult_97/n1588 ,
         \mult_97/n1587 , \mult_97/n1586 , \mult_97/n1585 , \mult_97/n1584 ,
         \mult_97/n1583 , \mult_97/n1582 , \mult_97/n1581 , \mult_97/n1580 ,
         \mult_97/n1579 , \mult_97/n1578 , \mult_97/n1577 , \mult_97/n1576 ,
         \mult_97/n1575 , \mult_97/n1574 , \mult_97/n1573 , \mult_97/n1572 ,
         \mult_97/n1571 , \mult_97/n1570 , \mult_97/n1569 , \mult_97/n1568 ,
         \mult_97/n1567 , \mult_97/n1566 , \mult_97/n1565 , \mult_97/n1564 ,
         \mult_97/n1563 , \mult_97/n1562 , \mult_97/n1561 , \mult_97/n1560 ,
         \mult_97/n1559 , \mult_97/n1558 , \mult_97/n1557 , \mult_97/n1556 ,
         \mult_97/n1555 , \mult_97/n1554 , \mult_97/n1553 , \mult_97/n1552 ,
         \mult_97/n1551 , \mult_97/n1550 , \mult_97/n1549 , \mult_97/n1548 ,
         \mult_97/n1547 , \mult_97/n1546 , \mult_97/n1545 , \mult_97/n1544 ,
         \mult_97/n1543 , \mult_97/n1542 , \mult_97/n1541 , \mult_97/n1540 ,
         \mult_97/n1539 , \mult_97/n1538 , \mult_97/n1537 , \mult_97/n1536 ,
         \mult_97/n1535 , \mult_97/n1534 , \mult_97/n1533 , \mult_97/n1532 ,
         \mult_97/n1531 , \mult_97/n1530 , \mult_97/n1529 , \mult_97/n1528 ,
         \mult_97/n1527 , \mult_97/n1526 , \mult_97/n1525 , \mult_97/n1524 ,
         \mult_97/n1523 , \mult_97/n1522 , \mult_97/n1521 , \mult_97/n1520 ,
         \mult_97/n1519 , \mult_97/n1518 , \mult_97/n1517 , \mult_97/n1516 ,
         \mult_97/n1515 , \mult_97/n1514 , \mult_97/n1513 , \mult_97/n1512 ,
         \mult_97/n1511 , \mult_97/n1510 , \mult_97/n1509 , \mult_97/n1508 ,
         \mult_97/n1507 , \mult_97/n1506 , \mult_97/n1505 , \mult_97/n1504 ,
         \mult_97/n1503 , \mult_97/n1502 , \mult_97/n1501 , \mult_97/n1500 ,
         \mult_97/n1499 , \mult_97/n1498 , \mult_97/n1497 , \mult_97/n1496 ,
         \mult_97/n1495 , \mult_97/n1494 , \mult_97/n1493 , \mult_97/n1492 ,
         \mult_97/n1491 , \mult_97/n1490 , \mult_97/n1489 , \mult_97/n1488 ,
         \mult_97/n1487 , \mult_97/n1486 , \mult_97/n1485 , \mult_97/n1484 ,
         \mult_97/n1483 , \mult_97/n1482 , \mult_97/n1481 , \mult_97/n1480 ,
         \mult_97/n1479 , \mult_97/n1478 , \mult_97/n1477 , \mult_97/n1476 ,
         \mult_97/n1475 , \mult_97/n1474 , \mult_97/n1473 , \mult_97/n1472 ,
         \mult_97/n1471 , \mult_97/n1470 , \mult_97/n1469 , \mult_97/n1468 ,
         \mult_97/n1467 , \mult_97/n1466 , \mult_97/n1465 , \mult_97/n1464 ,
         \mult_97/n1463 , \mult_97/n1462 , \mult_97/n1461 , \mult_97/n1460 ,
         \mult_97/n1459 , \mult_97/n1458 , \mult_97/n1457 , \mult_97/n1456 ,
         \mult_97/n1455 , \mult_97/n1454 , \mult_97/n1453 , \mult_97/n1452 ,
         \mult_97/n1451 , \mult_97/n1450 , \mult_97/n1449 , \mult_97/n1448 ,
         \mult_97/n1447 , \mult_97/n1446 , \mult_97/n1445 , \mult_97/n1444 ,
         \mult_97/n1443 , \mult_97/n1442 , \mult_97/n1441 , \mult_97/n1440 ,
         \mult_97/n1439 , \mult_97/n1438 , \mult_97/n1437 , \mult_97/n1436 ,
         \mult_97/n1435 , \mult_97/n1434 , \mult_97/n1433 , \mult_97/n1432 ,
         \mult_97/n1431 , \mult_97/n1430 , \mult_97/n1429 , \mult_97/n1428 ,
         \mult_97/n1427 , \mult_97/n1426 , \mult_97/n1425 , \mult_97/n1424 ,
         \mult_97/n1423 , \mult_97/n1422 , \mult_97/n1421 , \mult_97/n1420 ,
         \mult_97/n1419 , \mult_97/n1418 , \mult_97/n1417 , \mult_97/n1416 ,
         \mult_97/n1415 , \mult_97/n1414 , \mult_97/n1413 , \mult_97/n1412 ,
         \mult_97/n1411 , \mult_97/n1410 , \mult_97/n1409 , \mult_97/n1408 ,
         \mult_97/n1407 , \mult_97/n1406 , \mult_97/n1405 , \mult_97/n1404 ,
         \mult_97/n1403 , \mult_97/n1402 , \mult_97/n1401 , \mult_97/n1400 ,
         \mult_97/n1399 , \mult_97/n1398 , \mult_97/n1397 , \mult_97/n1396 ,
         \mult_97/n1395 , \mult_97/n1394 , \mult_97/n1393 , \mult_97/n1392 ,
         \mult_97/n1391 , \mult_97/n1390 , \mult_97/n1389 , \mult_97/n1388 ,
         \mult_97/n1387 , \mult_97/n1386 , \mult_97/n1385 , \mult_97/n1384 ,
         \mult_97/n1383 , \mult_97/n1382 , \mult_97/n1381 , \mult_97/n1380 ,
         \mult_97/n1379 , \mult_97/n1378 , \mult_97/n1377 , \mult_97/n1376 ,
         \mult_97/n1375 , \mult_97/n1374 , \mult_97/n1373 , \mult_97/n1372 ,
         \mult_97/n1371 , \mult_97/n1370 , \mult_97/n1369 , \mult_97/n1368 ,
         \mult_97/n1367 , \mult_97/n1366 , \mult_97/n1365 , \mult_97/n1364 ,
         \mult_97/n1363 , \mult_97/n1362 , \mult_97/n1361 , \mult_97/n1360 ,
         \mult_97/n1359 , \mult_97/n1358 , \mult_97/n1357 , \mult_97/n1356 ,
         \mult_97/n1355 , \mult_97/n1354 , \mult_97/n1353 , \mult_97/n1352 ,
         \mult_97/n1351 , \mult_97/n1350 , \mult_97/n1349 , \mult_97/n1348 ,
         \mult_97/n1347 , \mult_97/n1346 , \mult_97/n1345 , \mult_97/n1344 ,
         \mult_97/n1343 , \mult_97/n1342 , \mult_97/n1341 , \mult_97/n1340 ,
         \mult_97/n1339 , \mult_97/n1338 , \mult_97/n1337 , \mult_97/n1336 ,
         \mult_97/n1335 , \mult_97/n1334 , \mult_97/n1333 , \mult_97/n1332 ,
         \mult_97/n1331 , \mult_97/n1330 , \mult_97/n1329 , \mult_97/n1328 ,
         \mult_97/n1327 , \mult_97/n1326 , \mult_97/n1325 , \mult_97/n1324 ,
         \mult_97/n1323 , \mult_97/n1322 , \mult_97/n1321 , \mult_97/n1320 ,
         \mult_97/n1319 , \mult_97/n1318 , \mult_97/n1317 , \mult_97/n1316 ,
         \mult_97/n1315 , \mult_97/n1314 , \mult_97/n1313 , \mult_97/n1312 ,
         \mult_97/n1311 , \mult_97/n1310 , \mult_97/n1309 , \mult_97/n1308 ,
         \mult_97/n1307 , \mult_97/n1306 , \mult_97/n1305 , \mult_97/n1304 ,
         \mult_97/n1303 , \mult_97/n1302 , \mult_97/n1301 , \mult_97/n1300 ,
         \mult_97/n1299 , \mult_97/n1298 , \mult_97/n1297 , \mult_97/n1296 ,
         \mult_97/n1295 , \mult_97/n1294 , \mult_97/n1293 , \mult_97/n1292 ,
         \mult_97/n1291 , \mult_97/n1290 , \mult_97/n1289 , \mult_97/n1288 ,
         \mult_97/n1287 , \mult_97/n1286 , \mult_97/n1285 , \mult_97/n1284 ,
         \mult_97/n1283 , \mult_97/n1282 , \mult_97/n1281 , \mult_97/n1280 ,
         \mult_97/n1279 , \mult_97/n1278 , \mult_97/n1277 , \mult_97/n1276 ,
         \mult_97/n1275 , \mult_97/n1274 , \mult_97/n1273 , \mult_97/n1272 ,
         \mult_97/n1271 , \mult_97/n1270 , \mult_97/n1269 , \mult_97/n1268 ,
         \mult_97/n1267 , \mult_97/n1266 , \mult_97/n1265 , \mult_97/n1264 ,
         \mult_97/n1263 , \mult_97/n1262 , \mult_97/n1261 , \mult_97/n1260 ,
         \mult_97/n1259 , \mult_97/n1258 , \mult_97/n1257 , \mult_97/n1256 ,
         \mult_97/n1255 , \mult_97/n1254 , \mult_97/n1253 , \mult_97/n1252 ,
         \mult_97/n1251 , \mult_97/n1250 , \mult_97/n1249 , \mult_97/n1248 ,
         \mult_97/n1247 , \mult_97/n1246 , \mult_97/n1245 , \mult_97/n1244 ,
         \mult_97/n1243 , \mult_97/n1242 , \mult_97/n1241 , \mult_97/n1240 ,
         \mult_97/n1239 , \mult_97/n1238 , \mult_97/n1237 , \mult_97/n1236 ,
         \mult_97/n1235 , \mult_97/n1234 , \mult_97/n1233 , \mult_97/n1232 ,
         \mult_97/n1231 , \mult_97/n1230 , \mult_97/n1229 , \mult_97/n1228 ,
         \mult_97/n1227 , \mult_97/n1226 , \mult_97/n1225 , \mult_97/n1224 ,
         \mult_97/n1223 , \mult_97/n1222 , \mult_97/n1221 , \mult_97/n1220 ,
         \mult_97/n1219 , \mult_97/n1218 , \mult_97/n1217 , \mult_97/n1216 ,
         \mult_97/n1215 , \mult_97/n1214 , \mult_97/n1213 , \mult_97/n1212 ,
         \mult_97/n1211 , \mult_97/n1210 , \mult_97/n1209 , \mult_97/n1208 ,
         \mult_97/n1207 , \mult_97/n1206 , \mult_97/n1205 , \mult_97/n1204 ,
         \mult_97/n1203 , \mult_97/n1202 , \mult_97/n1201 , \mult_97/n1200 ,
         \mult_97/n1199 , \mult_97/n1198 , \mult_97/n1197 , \mult_97/n1196 ,
         \mult_97/n1195 , \mult_97/n1194 , \mult_97/n1193 , \mult_97/n1192 ,
         \mult_97/n1191 , \mult_97/n1190 , \mult_97/n1189 , \mult_97/n1188 ,
         \mult_97/n1187 , \mult_97/n1186 , \mult_97/n1185 , \mult_97/n1184 ,
         \mult_97/n1183 , \mult_97/n1182 , \mult_97/n1181 , \mult_97/n1180 ,
         \mult_97/n1179 , \mult_97/n1178 , \mult_97/n1177 , \mult_97/n1176 ,
         \mult_97/n1175 , \mult_97/n1174 , \mult_97/n1173 , \mult_97/n1172 ,
         \mult_97/n1171 , \mult_97/n1170 , \mult_97/n1169 , \mult_97/n1168 ,
         \mult_97/n1167 , \mult_97/n1166 , \mult_97/n1165 , \mult_97/n1164 ,
         \mult_97/n1163 , \mult_97/n1162 , \mult_97/n1161 , \mult_97/n1160 ,
         \mult_97/n1159 , \mult_97/n1158 , \mult_97/n1157 , \mult_97/n1156 ,
         \mult_97/n1155 , \mult_97/n1154 , \mult_97/n1153 , \mult_97/n1152 ,
         \mult_97/n1151 , \mult_97/n1150 , \mult_97/n1149 , \mult_97/n1148 ,
         \mult_97/n1147 , \mult_97/n1146 , \mult_97/n1145 , \mult_97/n1144 ,
         \mult_97/n1143 , \mult_97/n1142 , \mult_97/n1141 , \mult_97/n1140 ,
         \mult_97/n1139 , \mult_97/n1138 , \mult_97/n1137 , \mult_97/n1136 ,
         \mult_97/n1135 , \mult_97/n1134 , \mult_97/n1133 , \mult_97/n1132 ,
         \mult_97/n1131 , \mult_97/n1130 , \mult_97/n1129 , \mult_97/n1128 ,
         \mult_97/n1127 , \mult_97/n1126 , \mult_97/n1125 , \mult_97/n1124 ,
         \mult_97/n1123 , \mult_97/n1122 , \mult_97/n1121 , \mult_97/n1120 ,
         \mult_97/n1119 , \mult_97/n1118 , \mult_97/n1117 , \mult_97/n1116 ,
         \mult_97/n1115 , \mult_97/n1114 , \mult_97/n1113 , \mult_97/n1112 ,
         \mult_97/n1111 , \mult_97/n1110 , \mult_97/n1109 , \mult_97/n1108 ,
         \mult_97/n1107 , \mult_97/n1106 , \mult_97/n1105 , \mult_97/n1104 ,
         \mult_97/n1103 , \mult_97/n1102 , \mult_97/n1101 , \mult_97/n1100 ,
         \mult_97/n1099 , \mult_97/n1098 , \mult_97/n1097 , \mult_97/n1096 ,
         \mult_97/n1095 , \mult_97/n1094 , \mult_97/n1093 , \mult_97/n1092 ,
         \mult_97/n1091 , \mult_97/n1090 , \mult_97/n1089 , \mult_97/n1088 ,
         \mult_97/n1087 , \mult_97/n1086 , \mult_97/n1085 , \mult_97/n1084 ,
         \mult_97/n1083 , \mult_97/n1082 , \mult_97/n1081 , \mult_97/n1080 ,
         \mult_97/n1079 , \mult_97/n1078 , \mult_97/n1077 , \mult_97/n1076 ,
         \mult_97/n1075 , \mult_97/n1074 , \mult_97/n1073 , \mult_97/n1072 ,
         \mult_97/n1071 , \mult_97/n1070 , \mult_97/n1069 , \mult_97/n1068 ,
         \mult_97/n1067 , \mult_97/n1066 , \mult_97/n1065 , \mult_97/n1064 ,
         \mult_97/n1063 , \mult_97/n1062 , \mult_97/n1061 , \mult_97/n1060 ,
         \mult_97/n1059 , \mult_97/n1058 , \mult_97/n1057 , \mult_97/n1056 ,
         \mult_97/n1055 , \mult_97/n1054 , \mult_97/n1053 , \mult_97/n1052 ,
         \mult_97/n1051 , \mult_97/n1050 , \mult_97/n1049 , \mult_97/n1048 ,
         \mult_97/n1047 , \mult_97/n1046 , \mult_97/n1045 , \mult_97/n1044 ,
         \mult_97/n1043 , \mult_97/n1042 , \mult_97/n1041 , \mult_97/n1040 ,
         \mult_97/n1039 , \mult_97/n1038 , \mult_97/n1037 , \mult_97/n1036 ,
         \mult_97/n1035 , \mult_97/n1034 , \mult_97/n1033 , \mult_97/n1032 ,
         \mult_97/n1031 , \mult_97/n1030 , \mult_97/n1029 , \mult_97/n1028 ,
         \mult_97/n1027 , \mult_97/n1026 , \mult_97/n1025 , \mult_97/n1024 ,
         \mult_97/n1023 , \mult_97/n1022 , \mult_97/n1021 , \mult_97/n1020 ,
         \mult_97/n1019 , \mult_97/n1018 , \mult_97/n1017 , \mult_97/n1016 ,
         \mult_97/n1015 , \mult_97/n1014 , \mult_97/n1013 , \mult_97/n1012 ,
         \mult_97/n1011 , \mult_97/n1010 , \mult_97/n1009 , \mult_97/n1008 ,
         \mult_97/n1007 , \mult_97/n1006 , \mult_97/n1005 , \mult_97/n1004 ,
         \mult_97/n1003 , \mult_97/n1002 , \mult_97/n1001 , \mult_97/n1000 ,
         \mult_97/n999 , \mult_97/n998 , \mult_97/n997 , \mult_97/n996 ,
         \mult_97/n995 , \mult_97/n994 , \mult_97/n993 , \mult_97/n992 ,
         \mult_97/n991 , \mult_97/n990 , \mult_97/n989 , \mult_97/n988 ,
         \mult_97/n987 , \mult_97/n986 , \mult_97/n985 , \mult_97/n984 ,
         \mult_97/n983 , \mult_97/n982 , \mult_97/n981 , \mult_97/n980 ,
         \mult_97/n979 , \mult_97/n978 , \mult_97/n977 , \mult_97/n976 ,
         \mult_97/n975 , \mult_97/n974 , \mult_97/n973 , \mult_97/n972 ,
         \mult_97/n971 , \mult_97/n970 , \mult_97/n969 , \mult_97/n968 ,
         \mult_97/n967 , \mult_97/n966 , \mult_97/n965 , \mult_97/n964 ,
         \mult_97/n963 , \mult_97/n962 , \mult_97/n961 , \mult_97/n960 ,
         \mult_97/n959 , \mult_97/n958 , \mult_97/n957 , \mult_97/n956 ,
         \mult_97/n955 , \mult_97/n954 , \mult_97/n953 , \mult_97/n952 ,
         \mult_97/n951 , \mult_97/n950 , \mult_97/n949 , \mult_97/n948 ,
         \mult_97/n947 , \mult_97/n946 , \mult_97/n945 , \mult_97/n944 ,
         \mult_97/n943 , \mult_97/n942 , \mult_97/n941 , \mult_97/n940 ,
         \mult_97/n939 , \mult_97/n938 , \mult_97/n937 , \mult_97/n936 ,
         \mult_97/n935 , \mult_97/n934 , \mult_97/n933 , \mult_97/n932 ,
         \mult_97/n931 , \mult_97/n930 , \mult_97/n929 , \mult_97/n928 ,
         \mult_97/n927 , \mult_97/n926 , \mult_97/n925 , \mult_97/n924 ,
         \mult_97/n923 , \mult_97/n922 , \mult_97/n921 , \mult_97/n911 ,
         \mult_97/n905 , \mult_97/n904 , \mult_97/n903 , \mult_97/n901 ,
         \mult_97/n897 , \mult_97/n893 , \mult_97/n887 , \mult_97/n885 ,
         \mult_97/n883 , \mult_97/n881 , \mult_97/n880 , \mult_97/n878 ,
         \mult_97/n876 , \mult_97/n874 , \mult_97/n872 , \mult_97/n871 ,
         \mult_97/n868 , \mult_97/n862 , \mult_97/n861 , \mult_97/n859 ,
         \mult_97/n858 , \mult_97/n856 , \mult_97/n854 , \mult_97/n853 ,
         \mult_97/n852 , \mult_97/n851 , \mult_97/n850 , \mult_97/n848 ,
         \mult_97/n846 , \mult_97/n845 , \mult_97/n844 , \mult_97/n843 ,
         \mult_97/n842 , \mult_97/n841 , \mult_97/n840 , \mult_97/n838 ,
         \mult_97/n837 , \mult_97/n836 , \mult_97/n835 , \mult_97/n834 ,
         \mult_97/n833 , \mult_97/n832 , \mult_97/n831 , \mult_97/n830 ,
         \mult_97/n829 , \mult_97/n828 , \mult_97/n827 , \mult_97/n826 ,
         \mult_97/n825 , \mult_97/n822 , \mult_97/n821 , \mult_97/n820 ,
         \mult_97/n818 , \mult_97/n815 , \mult_97/n809 , \mult_97/n808 ,
         \mult_97/n807 , \mult_97/n806 , \mult_97/n804 , \mult_97/n803 ,
         \mult_97/n800 , \mult_97/n799 , \mult_97/n798 , \mult_97/n796 ,
         \mult_97/n793 , \mult_97/n792 , \mult_97/n791 , \mult_97/n789 ,
         \mult_97/n788 , \mult_97/n787 , \mult_97/n786 , \mult_97/n781 ,
         \mult_97/n780 , \mult_97/n778 , \mult_97/n777 , \mult_97/n774 ,
         \mult_97/n773 , \mult_97/n771 , \mult_97/n770 , \mult_97/n769 ,
         \mult_97/n768 , \mult_97/n767 , \mult_97/n766 , \mult_97/n765 ,
         \mult_97/n764 , \mult_97/n760 , \mult_97/n759 , \mult_97/n758 ,
         \mult_97/n757 , \mult_97/n756 , \mult_97/n755 , \mult_97/n754 ,
         \mult_97/n752 , \mult_97/n751 , \mult_97/n750 , \mult_97/n749 ,
         \mult_97/n748 , \mult_97/n747 , \mult_97/n746 , \mult_97/n745 ,
         \mult_97/n740 , \mult_97/n739 , \mult_97/n737 , \mult_97/n733 ,
         \mult_97/n732 , \mult_97/n731 , \mult_97/n730 , \mult_97/n728 ,
         \mult_97/n725 , \mult_97/n723 , \mult_97/n721 , \mult_97/n720 ,
         \mult_97/n719 , \mult_97/n718 , \mult_97/n717 , \mult_97/n716 ,
         \mult_97/n715 , \mult_97/n714 , \mult_97/n710 , \mult_97/n709 ,
         \mult_97/n708 , \mult_97/n707 , \mult_97/n706 , \mult_97/n705 ,
         \mult_97/n704 , \mult_97/n702 , \mult_97/n701 , \mult_97/n700 ,
         \mult_97/n699 , \mult_97/n698 , \mult_97/n697 , \mult_97/n696 ,
         \mult_97/n695 , \mult_97/n694 , \mult_97/n693 , \mult_97/n691 ,
         \mult_97/n690 , \mult_97/n689 , \mult_97/n688 , \mult_97/n687 ,
         \mult_97/n686 , \mult_97/n685 , \mult_97/n684 , \mult_97/n683 ,
         \mult_97/n679 , \mult_97/n678 , \mult_97/n677 , \mult_97/n676 ,
         \mult_97/n675 , \mult_97/n674 , \mult_97/n673 , \mult_97/n672 ,
         \mult_97/n671 , \mult_97/n670 , \mult_97/n666 , \mult_97/n665 ,
         \mult_97/n664 , \mult_97/n663 , \mult_97/n662 , \mult_97/n661 ,
         \mult_97/n660 , \mult_97/n659 , \mult_97/n658 , \mult_97/n654 ,
         \mult_97/n653 , \mult_97/n652 , \mult_97/n651 , \mult_97/n650 ,
         \mult_97/n649 , \mult_97/n648 , \mult_97/n647 , \mult_97/n646 ,
         \mult_97/n645 , \mult_97/n644 , \mult_97/n643 , \mult_97/n642 ,
         \mult_97/n640 , \mult_97/n637 , \mult_97/n635 , \mult_97/n634 ,
         \mult_97/n632 , \mult_97/n630 , \mult_97/n628 , \mult_97/n627 ,
         \mult_97/n626 , \mult_97/n625 , \mult_97/n624 , \mult_97/n623 ,
         \mult_97/n620 , \mult_97/n618 , \mult_97/n617 , \mult_97/n615 ,
         \mult_97/n613 , \mult_97/n611 , \mult_97/n610 , \mult_97/n609 ,
         \mult_97/n608 , \mult_97/n607 , \mult_97/n606 , \mult_97/n605 ,
         \mult_97/n604 , \mult_97/n600 , \mult_97/n599 , \mult_97/n598 ,
         \mult_97/n597 , \mult_97/n596 , \mult_97/n595 , \mult_97/n594 ,
         \mult_97/n593 , \mult_97/n592 , \mult_97/n588 , \mult_97/n587 ,
         \mult_97/n586 , \mult_97/n585 , \mult_97/n584 , \mult_97/n583 ,
         \mult_97/n582 , \mult_97/n581 , \mult_97/n580 , \mult_97/n579 ,
         \mult_97/n578 , \mult_97/n577 , \mult_97/n576 , \mult_97/n575 ,
         \mult_97/n572 , \mult_97/n570 , \mult_97/n569 , \mult_97/n567 ,
         \mult_97/n566 , \mult_97/n565 , \mult_97/n563 , \mult_97/n562 ,
         \mult_97/n561 , \mult_97/n560 , \mult_97/n559 , \mult_97/n558 ,
         \mult_97/n557 , \mult_97/n556 , \mult_97/n554 , \mult_97/n553 ,
         \mult_97/n552 , \mult_97/n551 , \mult_97/n549 , \mult_97/n548 ,
         \mult_97/n547 , \mult_97/n545 , \mult_97/n544 , \mult_97/n543 ,
         \mult_97/n542 , \mult_97/n541 , \mult_97/n540 , \mult_97/n538 ,
         \mult_97/n536 , \mult_97/n535 , \mult_97/n531 , \mult_97/n530 ,
         \mult_97/n529 , \mult_97/n528 , \mult_97/n526 , \mult_97/n524 ,
         \mult_97/n522 , \mult_97/n521 , \mult_97/n520 , \mult_97/n519 ,
         \mult_97/n517 , \mult_97/n511 , \mult_97/n510 , \mult_97/n508 ,
         \mult_97/n506 , \mult_97/n505 , \mult_97/n504 , \mult_97/n503 ,
         \mult_97/n502 , \mult_97/n492 , \mult_97/n485 , \mult_97/n478 ,
         \mult_97/n466 , \mult_97/n461 , \mult_97/n448 , \mult_97/n374 ,
         \mult_97/n371 , \mult_97/n368 , \mult_97/n362 , \mult_97/n353 , n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n55, n56, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n96,
         n97, n98, n99, n101, n102, n103, n104, n105, n106, n107, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n156, n157, n158, n159, n160, n161, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n559, n561, n563, n565, n567, n569, n571,
         n573, n575, n577;
  assign \A_extended[32]  = A[31];
  assign \B_extended[32]  = B[31];

  DFFPOSX1 clk_r_REG15_S2 ( .D(n632), .CLK(CLK), .Q(PRODUCT[63]) );
  DFFPOSX1 clk_r_REG16_S2 ( .D(n633), .CLK(CLK), .Q(PRODUCT[62]) );
  DFFPOSX1 clk_r_REG17_S2 ( .D(n634), .CLK(CLK), .Q(PRODUCT[61]) );
  DFFPOSX1 clk_r_REG18_S2 ( .D(n635), .CLK(CLK), .Q(PRODUCT[60]) );
  DFFPOSX1 clk_r_REG8_S2 ( .D(n642), .CLK(CLK), .Q(PRODUCT[53]) );
  DFFPOSX1 clk_r_REG10_S2 ( .D(n34), .CLK(CLK), .Q(PRODUCT[52]) );
  DFFPOSX1 clk_r_REG9_S2 ( .D(n644), .CLK(CLK), .Q(PRODUCT[51]) );
  DFFPOSX1 clk_r_REG4_S2 ( .D(n647), .CLK(CLK), .Q(PRODUCT[48]) );
  DFFPOSX1 clk_r_REG3_S2 ( .D(n648), .CLK(CLK), .Q(PRODUCT[47]) );
  DFFPOSX1 clk_r_REG2_S2 ( .D(n649), .CLK(CLK), .Q(PRODUCT[46]) );
  DFFPOSX1 clk_r_REG197_S1 ( .D(n686), .CLK(CLK), .Q(n577) );
  DFFPOSX1 clk_r_REG200_S1 ( .D(n687), .CLK(CLK), .Q(n575) );
  DFFPOSX1 clk_r_REG202_S1 ( .D(n688), .CLK(CLK), .Q(n573) );
  DFFPOSX1 clk_r_REG204_S1 ( .D(n689), .CLK(CLK), .Q(n571) );
  DFFPOSX1 clk_r_REG206_S1 ( .D(n690), .CLK(CLK), .Q(n569) );
  DFFPOSX1 clk_r_REG208_S1 ( .D(n691), .CLK(CLK), .Q(n567) );
  DFFPOSX1 \mult_97/clk_r_REG87_S1  ( .D(\mult_97/n1348 ), .CLK(CLK), .Q(n520)
         );
  DFFPOSX1 \mult_97/clk_r_REG86_S1  ( .D(\mult_97/n1347 ), .CLK(CLK), .Q(n519)
         );
  DFFPOSX1 \mult_97/clk_r_REG74_S1  ( .D(\mult_97/n1346 ), .CLK(CLK), .Q(n518)
         );
  DFFPOSX1 \mult_97/clk_r_REG73_S1  ( .D(\mult_97/n1345 ), .CLK(CLK), .Q(n517)
         );
  DFFPOSX1 \mult_97/clk_r_REG91_S1  ( .D(\mult_97/n1320 ), .CLK(CLK), .Q(n516)
         );
  DFFPOSX1 \mult_97/clk_r_REG90_S1  ( .D(\mult_97/n1319 ), .CLK(CLK), .Q(n515)
         );
  DFFPOSX1 \mult_97/clk_r_REG71_S1  ( .D(\mult_97/n1318 ), .CLK(CLK), .Q(n514)
         );
  DFFPOSX1 \mult_97/clk_r_REG66_S1  ( .D(\mult_97/n1317 ), .CLK(CLK), .Q(n513)
         );
  DFFPOSX1 \mult_97/clk_r_REG95_S1  ( .D(\mult_97/n1292 ), .CLK(CLK), .Q(n512)
         );
  DFFPOSX1 \mult_97/clk_r_REG94_S1  ( .D(\mult_97/n1291 ), .CLK(CLK), .Q(n511)
         );
  DFFPOSX1 \mult_97/clk_r_REG85_S1  ( .D(\mult_97/n1290 ), .CLK(CLK), .Q(n510)
         );
  DFFPOSX1 \mult_97/clk_r_REG84_S1  ( .D(\mult_97/n1289 ), .CLK(CLK), .Q(n509)
         );
  DFFPOSX1 \mult_97/clk_r_REG101_S1  ( .D(\mult_97/n1266 ), .CLK(CLK), .Q(n508) );
  DFFPOSX1 \mult_97/clk_r_REG89_S1  ( .D(\mult_97/n1264 ), .CLK(CLK), .Q(n507)
         );
  DFFPOSX1 \mult_97/clk_r_REG93_S1  ( .D(\mult_97/n1238 ), .CLK(CLK), .Q(n506)
         );
  DFFPOSX1 \mult_97/clk_r_REG104_S1  ( .D(\mult_97/n1214 ), .CLK(CLK), .Q(n505) );
  DFFPOSX1 \mult_97/clk_r_REG31_S1  ( .D(\mult_97/n1190 ), .CLK(CLK), .Q(n504)
         );
  DFFPOSX1 \mult_97/clk_r_REG30_S1  ( .D(\mult_97/n1189 ), .CLK(CLK), .Q(n503)
         );
  DFFPOSX1 \mult_97/clk_r_REG28_S1  ( .D(\mult_97/n1166 ), .CLK(CLK), .Q(n502)
         );
  DFFPOSX1 \mult_97/clk_r_REG27_S1  ( .D(\mult_97/n1165 ), .CLK(CLK), .Q(n501)
         );
  DFFPOSX1 \mult_97/clk_r_REG35_S1  ( .D(\mult_97/n1146 ), .CLK(CLK), .Q(n500)
         );
  DFFPOSX1 \mult_97/clk_r_REG25_S1  ( .D(\mult_97/n1144 ), .CLK(CLK), .Q(n499)
         );
  DFFPOSX1 \mult_97/clk_r_REG24_S1  ( .D(\mult_97/n1143 ), .CLK(CLK), .Q(n498)
         );
  DFFPOSX1 \mult_97/clk_r_REG125_S1  ( .D(\mult_97/n1126 ), .CLK(CLK), .Q(n497) );
  DFFPOSX1 \mult_97/clk_r_REG22_S1  ( .D(\mult_97/n1124 ), .CLK(CLK), .Q(n496)
         );
  DFFPOSX1 \mult_97/clk_r_REG0_S1  ( .D(\mult_97/n1123 ), .CLK(CLK), .Q(n495)
         );
  DFFPOSX1 \mult_97/clk_r_REG124_S1  ( .D(\mult_97/n1106 ), .CLK(CLK), .Q(n494) );
  DFFPOSX1 \mult_97/clk_r_REG34_S1  ( .D(\mult_97/n1104 ), .CLK(CLK), .Q(n493)
         );
  DFFPOSX1 \mult_97/clk_r_REG33_S1  ( .D(\mult_97/n1103 ), .CLK(CLK), .Q(n492)
         );
  DFFPOSX1 \mult_97/clk_r_REG63_S1  ( .D(\mult_97/n1088 ), .CLK(CLK), .Q(n491)
         );
  DFFPOSX1 \mult_97/clk_r_REG65_S1  ( .D(\mult_97/n1086 ), .CLK(CLK), .Q(n490)
         );
  DFFPOSX1 \mult_97/clk_r_REG64_S1  ( .D(\mult_97/n1085 ), .CLK(CLK), .Q(n489)
         );
  DFFPOSX1 \mult_97/clk_r_REG62_S1  ( .D(\mult_97/n1070 ), .CLK(CLK), .Q(n488)
         );
  DFFPOSX1 \mult_97/clk_r_REG61_S1  ( .D(\mult_97/n1068 ), .CLK(CLK), .Q(n487)
         );
  DFFPOSX1 \mult_97/clk_r_REG60_S1  ( .D(\mult_97/n1067 ), .CLK(CLK), .Q(n486)
         );
  DFFPOSX1 \mult_97/clk_r_REG126_S1  ( .D(\mult_97/n1054 ), .CLK(CLK), .Q(n485) );
  DFFPOSX1 \mult_97/clk_r_REG59_S1  ( .D(\mult_97/n1052 ), .CLK(CLK), .Q(n484)
         );
  DFFPOSX1 \mult_97/clk_r_REG58_S1  ( .D(\mult_97/n1051 ), .CLK(CLK), .Q(n483)
         );
  DFFPOSX1 \mult_97/clk_r_REG113_S1  ( .D(\mult_97/n1038 ), .CLK(CLK), .Q(n482) );
  DFFPOSX1 \mult_97/clk_r_REG57_S1  ( .D(\mult_97/n1036 ), .CLK(CLK), .Q(n481)
         );
  DFFPOSX1 \mult_97/clk_r_REG110_S1  ( .D(\mult_97/n1006 ), .CLK(CLK), .Q(n480) );
  DFFPOSX1 \mult_97/clk_r_REG196_S1  ( .D(\mult_97/n822 ), .CLK(CLK), .Q(n474)
         );
  DFFPOSX1 \mult_97/clk_r_REG193_S1  ( .D(\mult_97/n820 ), .CLK(CLK), .Q(n473)
         );
  DFFPOSX1 \mult_97/clk_r_REG190_S1  ( .D(\mult_97/n815 ), .CLK(CLK), .Q(n472)
         );
  DFFPOSX1 \mult_97/clk_r_REG187_S1  ( .D(\mult_97/n807 ), .CLK(CLK), .Q(n471)
         );
  DFFPOSX1 \mult_97/clk_r_REG185_S1  ( .D(\mult_97/n806 ), .CLK(CLK), .Q(n470)
         );
  DFFPOSX1 \mult_97/clk_r_REG184_S1  ( .D(\mult_97/n804 ), .CLK(CLK), .Q(n469)
         );
  DFFPOSX1 \mult_97/clk_r_REG182_S1  ( .D(\mult_97/n803 ), .CLK(CLK), .Q(n468)
         );
  DFFPOSX1 \mult_97/clk_r_REG181_S1  ( .D(\mult_97/n798 ), .CLK(CLK), .Q(n467)
         );
  DFFPOSX1 \mult_97/clk_r_REG178_S1  ( .D(\mult_97/n793 ), .CLK(CLK), .Q(n466)
         );
  DFFPOSX1 \mult_97/clk_r_REG176_S1  ( .D(\mult_97/n792 ), .CLK(CLK), .Q(n465)
         );
  DFFPOSX1 \mult_97/clk_r_REG175_S1  ( .D(\mult_97/n781 ), .CLK(CLK), .Q(n464)
         );
  DFFPOSX1 \mult_97/clk_r_REG173_S1  ( .D(\mult_97/n780 ), .CLK(CLK), .Q(n463)
         );
  DFFPOSX1 \mult_97/clk_r_REG172_S1  ( .D(\mult_97/n778 ), .CLK(CLK), .Q(n462)
         );
  DFFPOSX1 \mult_97/clk_r_REG170_S1  ( .D(\mult_97/n777 ), .CLK(CLK), .Q(n461)
         );
  DFFPOSX1 \mult_97/clk_r_REG109_S1  ( .D(\mult_97/n567 ), .CLK(CLK), .Q(n460)
         );
  DFFPOSX1 \mult_97/clk_r_REG108_S1  ( .D(\mult_97/n566 ), .CLK(CLK), .Q(n459)
         );
  DFFPOSX1 \mult_97/clk_r_REG107_S1  ( .D(\mult_97/n557 ), .CLK(CLK), .Q(n458)
         );
  DFFPOSX1 \mult_97/clk_r_REG106_S1  ( .D(\mult_97/n556 ), .CLK(CLK), .Q(n457)
         );
  DFFPOSX1 \mult_97/clk_r_REG55_S1  ( .D(\mult_97/n554 ), .CLK(CLK), .Q(n456)
         );
  DFFPOSX1 \mult_97/clk_r_REG54_S1  ( .D(\mult_97/n553 ), .CLK(CLK), .Q(n455)
         );
  DFFPOSX1 \mult_97/clk_r_REG41_S1  ( .D(\mult_97/n549 ), .CLK(CLK), .Q(n454)
         );
  DFFPOSX1 \mult_97/clk_r_REG40_S1  ( .D(\mult_97/n548 ), .CLK(CLK), .Q(n453)
         );
  DFFPOSX1 \mult_97/clk_r_REG39_S1  ( .D(\mult_97/n540 ), .CLK(CLK), .Q(n452)
         );
  DFFPOSX1 \mult_97/clk_r_REG37_S1  ( .D(\mult_97/n531 ), .CLK(CLK), .Q(n451)
         );
  DFFPOSX1 \mult_97/clk_r_REG36_S1  ( .D(\mult_97/n530 ), .CLK(CLK), .Q(n450)
         );
  DFFPOSX1 \mult_97/clk_r_REG43_S1  ( .D(\mult_97/n526 ), .CLK(CLK), .Q(n449)
         );
  DFFPOSX1 \mult_97/clk_r_REG47_S1  ( .D(\mult_97/n517 ), .CLK(CLK), .Q(n448)
         );
  DFFPOSX1 \mult_97/clk_r_REG45_S1  ( .D(\mult_97/n510 ), .CLK(CLK), .Q(n447)
         );
  DFFPOSX1 \mult_97/clk_r_REG169_S1  ( .D(\mult_97/n1707 ), .CLK(CLK), .Q(n445) );
  DFFPOSX1 \mult_97/clk_r_REG164_S1  ( .D(\mult_97/n1690 ), .CLK(CLK), .Q(n444) );
  DFFPOSX1 \mult_97/clk_r_REG163_S1  ( .D(\mult_97/n1689 ), .CLK(CLK), .Q(n443) );
  DFFPOSX1 \mult_97/clk_r_REG151_S1  ( .D(\mult_97/n1633 ), .CLK(CLK), .Q(n442) );
  DFFPOSX1 \mult_97/clk_r_REG149_S1  ( .D(\mult_97/n1614 ), .CLK(CLK), .Q(n441) );
  DFFPOSX1 \mult_97/clk_r_REG155_S1  ( .D(\mult_97/n1612 ), .CLK(CLK), .Q(n440) );
  DFFPOSX1 \mult_97/clk_r_REG154_S1  ( .D(\mult_97/n1611 ), .CLK(CLK), .Q(n439) );
  DFFPOSX1 \mult_97/clk_r_REG148_S1  ( .D(\mult_97/n1592 ), .CLK(CLK), .Q(n438) );
  DFFPOSX1 \mult_97/clk_r_REG146_S1  ( .D(\mult_97/n1590 ), .CLK(CLK), .Q(n437) );
  DFFPOSX1 \mult_97/clk_r_REG145_S1  ( .D(\mult_97/n1589 ), .CLK(CLK), .Q(n436) );
  DFFPOSX1 \mult_97/clk_r_REG144_S1  ( .D(\mult_97/n1568 ), .CLK(CLK), .Q(n435) );
  DFFPOSX1 \mult_97/clk_r_REG142_S1  ( .D(\mult_97/n1566 ), .CLK(CLK), .Q(n434) );
  DFFPOSX1 \mult_97/clk_r_REG141_S1  ( .D(\mult_97/n1565 ), .CLK(CLK), .Q(n433) );
  DFFPOSX1 \mult_97/clk_r_REG137_S1  ( .D(\mult_97/n1544 ), .CLK(CLK), .Q(n432) );
  DFFPOSX1 \mult_97/clk_r_REG140_S1  ( .D(\mult_97/n1542 ), .CLK(CLK), .Q(n431) );
  DFFPOSX1 \mult_97/clk_r_REG139_S1  ( .D(\mult_97/n1541 ), .CLK(CLK), .Q(n430) );
  DFFPOSX1 \mult_97/clk_r_REG132_S1  ( .D(\mult_97/n1518 ), .CLK(CLK), .Q(n429) );
  DFFPOSX1 \mult_97/clk_r_REG136_S1  ( .D(\mult_97/n1516 ), .CLK(CLK), .Q(n428) );
  DFFPOSX1 \mult_97/clk_r_REG135_S1  ( .D(\mult_97/n1515 ), .CLK(CLK), .Q(n427) );
  DFFPOSX1 \mult_97/clk_r_REG134_S1  ( .D(\mult_97/n1492 ), .CLK(CLK), .Q(n426) );
  DFFPOSX1 \mult_97/clk_r_REG130_S1  ( .D(\mult_97/n1490 ), .CLK(CLK), .Q(n425) );
  DFFPOSX1 \mult_97/clk_r_REG129_S1  ( .D(\mult_97/n1489 ), .CLK(CLK), .Q(n424) );
  DFFPOSX1 \mult_97/clk_r_REG120_S1  ( .D(\mult_97/n1464 ), .CLK(CLK), .Q(n423) );
  DFFPOSX1 \mult_97/clk_r_REG128_S1  ( .D(\mult_97/n1462 ), .CLK(CLK), .Q(n422) );
  DFFPOSX1 \mult_97/clk_r_REG127_S1  ( .D(\mult_97/n1461 ), .CLK(CLK), .Q(n421) );
  DFFPOSX1 \mult_97/clk_r_REG123_S1  ( .D(\mult_97/n1436 ), .CLK(CLK), .Q(n420) );
  DFFPOSX1 \mult_97/clk_r_REG117_S1  ( .D(\mult_97/n1434 ), .CLK(CLK), .Q(n419) );
  DFFPOSX1 \mult_97/clk_r_REG116_S1  ( .D(\mult_97/n1433 ), .CLK(CLK), .Q(n418) );
  DFFPOSX1 \mult_97/clk_r_REG115_S1  ( .D(\mult_97/n1406 ), .CLK(CLK), .Q(n417) );
  DFFPOSX1 \mult_97/clk_r_REG114_S1  ( .D(\mult_97/n1405 ), .CLK(CLK), .Q(n416) );
  DFFPOSX1 \mult_97/clk_r_REG79_S1  ( .D(\mult_97/n1380 ), .CLK(CLK), .Q(n415)
         );
  DFFPOSX1 \mult_97/clk_r_REG77_S1  ( .D(\mult_97/n1378 ), .CLK(CLK), .Q(n414)
         );
  DFFPOSX1 \mult_97/clk_r_REG76_S1  ( .D(\mult_97/n1377 ), .CLK(CLK), .Q(n413)
         );
  DFFPOSX1 \mult_97/clk_r_REG81_S1  ( .D(\mult_97/n1376 ), .CLK(CLK), .Q(n412)
         );
  DFFPOSX1 \mult_97/clk_r_REG80_S1  ( .D(\mult_97/n1375 ), .CLK(CLK), .Q(n411)
         );
  DFFPOSX1 \mult_97/clk_r_REG44_S1  ( .D(n526), .CLK(CLK), .Q(n409) );
  DFFPOSX1 \mult_97/clk_r_REG46_S1  ( .D(n527), .CLK(CLK), .Q(n408) );
  DFFPOSX1 \mult_97/clk_r_REG42_S1  ( .D(n525), .CLK(CLK), .Q(n407) );
  DFFPOSX1 \mult_97/clk_r_REG38_S1  ( .D(n524), .CLK(CLK), .Q(n406) );
  DFFPOSX1 \mult_97/clk_r_REG179_S1  ( .D(n523), .CLK(CLK), .Q(n405) );
  DFFPOSX1 \mult_97/clk_r_REG188_S1  ( .D(n522), .CLK(CLK), .Q(n404) );
  DFFPOSX1 \mult_97/clk_r_REG191_S1  ( .D(n521), .CLK(CLK), .Q(n403) );
  XOR2X1 \mult_97/U2375  ( .A(A[2]), .B(n304), .Y(\mult_97/n2953 ) );
  XNOR2X1 \mult_97/U2373  ( .A(A[4]), .B(n305), .Y(\mult_97/n353 ) );
  XOR2X1 \mult_97/U2372  ( .A(n302), .B(A[4]), .Y(\mult_97/n2952 ) );
  XOR2X1 \mult_97/U2369  ( .A(A[6]), .B(n299), .Y(\mult_97/n2951 ) );
  XOR2X1 \mult_97/U2366  ( .A(A[8]), .B(n296), .Y(\mult_97/n2950 ) );
  XNOR2X1 \mult_97/U2364  ( .A(A[10]), .B(n297), .Y(\mult_97/n362 ) );
  XOR2X1 \mult_97/U2363  ( .A(n294), .B(A[10]), .Y(\mult_97/n2949 ) );
  XOR2X1 \mult_97/U2360  ( .A(A[12]), .B(n291), .Y(\mult_97/n2948 ) );
  XNOR2X1 \mult_97/U2358  ( .A(A[14]), .B(n292), .Y(\mult_97/n368 ) );
  XOR2X1 \mult_97/U2357  ( .A(A[14]), .B(n289), .Y(\mult_97/n2947 ) );
  XNOR2X1 \mult_97/U2355  ( .A(A[16]), .B(A[15]), .Y(\mult_97/n371 ) );
  XOR2X1 \mult_97/U2354  ( .A(n286), .B(A[16]), .Y(\mult_97/n2946 ) );
  XNOR2X1 \mult_97/U2352  ( .A(n287), .B(A[18]), .Y(\mult_97/n374 ) );
  XOR2X1 \mult_97/U2351  ( .A(A[18]), .B(n283), .Y(\mult_97/n2945 ) );
  XOR2X1 \mult_97/U2348  ( .A(A[20]), .B(n281), .Y(\mult_97/n2944 ) );
  XOR2X1 \mult_97/U2345  ( .A(n279), .B(A[22]), .Y(\mult_97/n2943 ) );
  XOR2X1 \mult_97/U2342  ( .A(A[24]), .B(n276), .Y(\mult_97/n2942 ) );
  XOR2X1 \mult_97/U2339  ( .A(A[26]), .B(n274), .Y(\mult_97/n2941 ) );
  XOR2X1 \mult_97/U2336  ( .A(n272), .B(A[28]), .Y(\mult_97/n2940 ) );
  XOR2X1 \mult_97/U2333  ( .A(\A_extended[32] ), .B(A[30]), .Y(\mult_97/n2939 ) );
  XNOR2X1 \mult_97/U2269  ( .A(n251), .B(n308), .Y(\mult_97/n2905 ) );
  XNOR2X1 \mult_97/U2268  ( .A(n400), .B(n308), .Y(\mult_97/n2904 ) );
  XNOR2X1 \mult_97/U2267  ( .A(n398), .B(n308), .Y(\mult_97/n2903 ) );
  XNOR2X1 \mult_97/U2266  ( .A(n396), .B(n308), .Y(\mult_97/n2902 ) );
  XNOR2X1 \mult_97/U2265  ( .A(n394), .B(n308), .Y(\mult_97/n2901 ) );
  XNOR2X1 \mult_97/U2264  ( .A(n392), .B(n308), .Y(\mult_97/n2900 ) );
  XNOR2X1 \mult_97/U2263  ( .A(n390), .B(n308), .Y(\mult_97/n2899 ) );
  XNOR2X1 \mult_97/U2262  ( .A(n388), .B(n308), .Y(\mult_97/n2898 ) );
  XNOR2X1 \mult_97/U2261  ( .A(n386), .B(n307), .Y(\mult_97/n2897 ) );
  XNOR2X1 \mult_97/U2260  ( .A(n384), .B(n308), .Y(\mult_97/n2896 ) );
  XNOR2X1 \mult_97/U2259  ( .A(n382), .B(n308), .Y(\mult_97/n2895 ) );
  XNOR2X1 \mult_97/U2258  ( .A(n380), .B(n307), .Y(\mult_97/n2894 ) );
  XNOR2X1 \mult_97/U2257  ( .A(n378), .B(n307), .Y(\mult_97/n2893 ) );
  XNOR2X1 \mult_97/U2256  ( .A(n376), .B(n307), .Y(\mult_97/n2892 ) );
  XNOR2X1 \mult_97/U2255  ( .A(n374), .B(n307), .Y(\mult_97/n2891 ) );
  XNOR2X1 \mult_97/U2254  ( .A(n372), .B(n307), .Y(\mult_97/n2890 ) );
  XNOR2X1 \mult_97/U2253  ( .A(n370), .B(n307), .Y(\mult_97/n2889 ) );
  XNOR2X1 \mult_97/U2252  ( .A(n368), .B(n307), .Y(\mult_97/n2888 ) );
  XNOR2X1 \mult_97/U2251  ( .A(n366), .B(n307), .Y(\mult_97/n2887 ) );
  XNOR2X1 \mult_97/U2250  ( .A(n364), .B(n307), .Y(\mult_97/n2886 ) );
  XNOR2X1 \mult_97/U2249  ( .A(n362), .B(n307), .Y(\mult_97/n2885 ) );
  XNOR2X1 \mult_97/U2248  ( .A(n360), .B(n307), .Y(\mult_97/n2884 ) );
  XNOR2X1 \mult_97/U2247  ( .A(n358), .B(n307), .Y(\mult_97/n2883 ) );
  XNOR2X1 \mult_97/U2246  ( .A(n356), .B(n307), .Y(\mult_97/n2882 ) );
  XNOR2X1 \mult_97/U2245  ( .A(n354), .B(n307), .Y(\mult_97/n2881 ) );
  XNOR2X1 \mult_97/U2244  ( .A(n352), .B(n307), .Y(\mult_97/n2880 ) );
  XNOR2X1 \mult_97/U2243  ( .A(n350), .B(n307), .Y(\mult_97/n2879 ) );
  XNOR2X1 \mult_97/U2242  ( .A(n348), .B(n307), .Y(\mult_97/n2878 ) );
  XNOR2X1 \mult_97/U2241  ( .A(n346), .B(n307), .Y(\mult_97/n2877 ) );
  XNOR2X1 \mult_97/U2240  ( .A(n344), .B(n307), .Y(\mult_97/n2876 ) );
  XNOR2X1 \mult_97/U2239  ( .A(n342), .B(n307), .Y(\mult_97/n2875 ) );
  XNOR2X1 \mult_97/U2238  ( .A(n340), .B(n308), .Y(\mult_97/n2874 ) );
  OAI22X1 \mult_97/U2237  ( .A(n309), .B(\mult_97/n2904 ), .C(n246), .D(
        \mult_97/n2905 ), .Y(\mult_97/n2378 ) );
  OAI22X1 \mult_97/U2236  ( .A(n246), .B(\mult_97/n2904 ), .C(n309), .D(
        \mult_97/n2903 ), .Y(\mult_97/n2377 ) );
  OAI22X1 \mult_97/U2235  ( .A(n246), .B(\mult_97/n2903 ), .C(n309), .D(
        \mult_97/n2902 ), .Y(\mult_97/n2376 ) );
  OAI22X1 \mult_97/U2234  ( .A(n246), .B(\mult_97/n2902 ), .C(n309), .D(
        \mult_97/n2901 ), .Y(\mult_97/n2375 ) );
  OAI22X1 \mult_97/U2233  ( .A(n246), .B(\mult_97/n2901 ), .C(n309), .D(
        \mult_97/n2900 ), .Y(\mult_97/n2374 ) );
  OAI22X1 \mult_97/U2232  ( .A(n246), .B(\mult_97/n2900 ), .C(n309), .D(
        \mult_97/n2899 ), .Y(\mult_97/n2373 ) );
  OAI22X1 \mult_97/U2231  ( .A(n309), .B(\mult_97/n2898 ), .C(n246), .D(
        \mult_97/n2899 ), .Y(\mult_97/n2372 ) );
  OAI22X1 \mult_97/U2230  ( .A(n246), .B(\mult_97/n2898 ), .C(n309), .D(
        \mult_97/n2897 ), .Y(\mult_97/n2371 ) );
  OAI22X1 \mult_97/U2229  ( .A(n246), .B(\mult_97/n2897 ), .C(n309), .D(
        \mult_97/n2896 ), .Y(\mult_97/n2370 ) );
  OAI22X1 \mult_97/U2228  ( .A(n246), .B(\mult_97/n2896 ), .C(n309), .D(
        \mult_97/n2895 ), .Y(\mult_97/n2369 ) );
  OAI22X1 \mult_97/U2227  ( .A(n246), .B(\mult_97/n2895 ), .C(n309), .D(
        \mult_97/n2894 ), .Y(\mult_97/n2368 ) );
  OAI22X1 \mult_97/U2226  ( .A(n246), .B(\mult_97/n2894 ), .C(n309), .D(
        \mult_97/n2893 ), .Y(\mult_97/n2367 ) );
  OAI22X1 \mult_97/U2225  ( .A(n246), .B(\mult_97/n2893 ), .C(n309), .D(
        \mult_97/n2892 ), .Y(\mult_97/n2366 ) );
  OAI22X1 \mult_97/U2224  ( .A(n246), .B(\mult_97/n2892 ), .C(n309), .D(
        \mult_97/n2891 ), .Y(\mult_97/n2365 ) );
  OAI22X1 \mult_97/U2223  ( .A(n246), .B(\mult_97/n2891 ), .C(n309), .D(
        \mult_97/n2890 ), .Y(\mult_97/n2364 ) );
  OAI22X1 \mult_97/U2222  ( .A(n246), .B(\mult_97/n2890 ), .C(n309), .D(
        \mult_97/n2889 ), .Y(\mult_97/n2363 ) );
  OAI22X1 \mult_97/U2221  ( .A(n246), .B(\mult_97/n2889 ), .C(n309), .D(
        \mult_97/n2888 ), .Y(\mult_97/n2362 ) );
  OAI22X1 \mult_97/U2220  ( .A(n246), .B(\mult_97/n2888 ), .C(n309), .D(
        \mult_97/n2887 ), .Y(\mult_97/n2361 ) );
  OAI22X1 \mult_97/U2219  ( .A(n246), .B(\mult_97/n2887 ), .C(n309), .D(
        \mult_97/n2886 ), .Y(\mult_97/n2360 ) );
  OAI22X1 \mult_97/U2218  ( .A(n246), .B(\mult_97/n2886 ), .C(n309), .D(
        \mult_97/n2885 ), .Y(\mult_97/n2359 ) );
  OAI22X1 \mult_97/U2217  ( .A(n246), .B(\mult_97/n2885 ), .C(n309), .D(
        \mult_97/n2884 ), .Y(\mult_97/n2358 ) );
  OAI22X1 \mult_97/U2216  ( .A(n246), .B(\mult_97/n2884 ), .C(n309), .D(
        \mult_97/n2883 ), .Y(\mult_97/n2357 ) );
  OAI22X1 \mult_97/U2215  ( .A(n246), .B(\mult_97/n2883 ), .C(n309), .D(
        \mult_97/n2882 ), .Y(\mult_97/n2356 ) );
  OAI22X1 \mult_97/U2214  ( .A(n246), .B(\mult_97/n2882 ), .C(n309), .D(
        \mult_97/n2881 ), .Y(\mult_97/n2355 ) );
  OAI22X1 \mult_97/U2213  ( .A(n246), .B(\mult_97/n2881 ), .C(n309), .D(
        \mult_97/n2880 ), .Y(\mult_97/n2354 ) );
  OAI22X1 \mult_97/U2212  ( .A(n246), .B(\mult_97/n2880 ), .C(n309), .D(
        \mult_97/n2879 ), .Y(\mult_97/n2353 ) );
  OAI22X1 \mult_97/U2211  ( .A(n246), .B(\mult_97/n2879 ), .C(n309), .D(
        \mult_97/n2878 ), .Y(\mult_97/n2352 ) );
  OAI22X1 \mult_97/U2210  ( .A(n246), .B(\mult_97/n2878 ), .C(n309), .D(
        \mult_97/n2877 ), .Y(\mult_97/n2351 ) );
  OAI22X1 \mult_97/U2209  ( .A(n246), .B(\mult_97/n2877 ), .C(n309), .D(
        \mult_97/n2876 ), .Y(\mult_97/n2350 ) );
  OAI22X1 \mult_97/U2208  ( .A(n309), .B(\mult_97/n2875 ), .C(n246), .D(
        \mult_97/n2876 ), .Y(\mult_97/n2349 ) );
  OAI22X1 \mult_97/U2207  ( .A(n246), .B(\mult_97/n2875 ), .C(n309), .D(
        \mult_97/n2874 ), .Y(\mult_97/n2348 ) );
  OAI22X1 \mult_97/U2206  ( .A(n306), .B(n246), .C(n309), .D(\mult_97/n2906 ), 
        .Y(\mult_97/n1866 ) );
  XNOR2X1 \mult_97/U2205  ( .A(n251), .B(n305), .Y(\mult_97/n2872 ) );
  XNOR2X1 \mult_97/U2204  ( .A(n400), .B(n305), .Y(\mult_97/n2871 ) );
  XNOR2X1 \mult_97/U2203  ( .A(n398), .B(n305), .Y(\mult_97/n2870 ) );
  XNOR2X1 \mult_97/U2202  ( .A(n396), .B(n305), .Y(\mult_97/n2869 ) );
  XNOR2X1 \mult_97/U2201  ( .A(n394), .B(n305), .Y(\mult_97/n2868 ) );
  XNOR2X1 \mult_97/U2200  ( .A(n392), .B(n305), .Y(\mult_97/n2867 ) );
  XNOR2X1 \mult_97/U2199  ( .A(n390), .B(n305), .Y(\mult_97/n2866 ) );
  XNOR2X1 \mult_97/U2198  ( .A(n388), .B(n305), .Y(\mult_97/n2865 ) );
  XNOR2X1 \mult_97/U2197  ( .A(n386), .B(n304), .Y(\mult_97/n2864 ) );
  XNOR2X1 \mult_97/U2196  ( .A(n384), .B(n305), .Y(\mult_97/n2863 ) );
  XNOR2X1 \mult_97/U2195  ( .A(n382), .B(n305), .Y(\mult_97/n2862 ) );
  XNOR2X1 \mult_97/U2194  ( .A(n380), .B(n304), .Y(\mult_97/n2861 ) );
  XNOR2X1 \mult_97/U2193  ( .A(n378), .B(n304), .Y(\mult_97/n2860 ) );
  XNOR2X1 \mult_97/U2192  ( .A(n376), .B(n304), .Y(\mult_97/n2859 ) );
  XNOR2X1 \mult_97/U2191  ( .A(n374), .B(n304), .Y(\mult_97/n2858 ) );
  XNOR2X1 \mult_97/U2190  ( .A(n372), .B(n304), .Y(\mult_97/n2857 ) );
  XNOR2X1 \mult_97/U2189  ( .A(n370), .B(n304), .Y(\mult_97/n2856 ) );
  XNOR2X1 \mult_97/U2188  ( .A(n368), .B(n304), .Y(\mult_97/n2855 ) );
  XNOR2X1 \mult_97/U2187  ( .A(n366), .B(n304), .Y(\mult_97/n2854 ) );
  XNOR2X1 \mult_97/U2186  ( .A(B[19]), .B(n304), .Y(\mult_97/n2853 ) );
  XNOR2X1 \mult_97/U2185  ( .A(n362), .B(n304), .Y(\mult_97/n2852 ) );
  XNOR2X1 \mult_97/U2184  ( .A(n360), .B(n304), .Y(\mult_97/n2851 ) );
  XNOR2X1 \mult_97/U2183  ( .A(n358), .B(n304), .Y(\mult_97/n2850 ) );
  XNOR2X1 \mult_97/U2182  ( .A(n356), .B(n304), .Y(\mult_97/n2849 ) );
  XNOR2X1 \mult_97/U2181  ( .A(n354), .B(n304), .Y(\mult_97/n2848 ) );
  XNOR2X1 \mult_97/U2180  ( .A(n352), .B(n304), .Y(\mult_97/n2847 ) );
  XNOR2X1 \mult_97/U2179  ( .A(n350), .B(n304), .Y(\mult_97/n2846 ) );
  XNOR2X1 \mult_97/U2178  ( .A(n348), .B(n304), .Y(\mult_97/n2845 ) );
  XNOR2X1 \mult_97/U2177  ( .A(n346), .B(n304), .Y(\mult_97/n2844 ) );
  XNOR2X1 \mult_97/U2176  ( .A(n344), .B(n304), .Y(\mult_97/n2843 ) );
  XNOR2X1 \mult_97/U2175  ( .A(n342), .B(n304), .Y(\mult_97/n2842 ) );
  XNOR2X1 \mult_97/U2174  ( .A(n340), .B(n305), .Y(\mult_97/n2841 ) );
  OAI22X1 \mult_97/U2173  ( .A(\mult_97/n2871 ), .B(n311), .C(\mult_97/n2872 ), 
        .D(n244), .Y(\mult_97/n2345 ) );
  OAI22X1 \mult_97/U2172  ( .A(\mult_97/n2870 ), .B(n311), .C(\mult_97/n2871 ), 
        .D(n244), .Y(\mult_97/n2344 ) );
  OAI22X1 \mult_97/U2171  ( .A(\mult_97/n2869 ), .B(n311), .C(\mult_97/n2870 ), 
        .D(n244), .Y(\mult_97/n2343 ) );
  OAI22X1 \mult_97/U2170  ( .A(\mult_97/n2868 ), .B(n311), .C(\mult_97/n2869 ), 
        .D(n244), .Y(\mult_97/n2342 ) );
  OAI22X1 \mult_97/U2169  ( .A(\mult_97/n2867 ), .B(n311), .C(\mult_97/n2868 ), 
        .D(n244), .Y(\mult_97/n2341 ) );
  OAI22X1 \mult_97/U2168  ( .A(\mult_97/n2866 ), .B(n311), .C(\mult_97/n2867 ), 
        .D(n244), .Y(\mult_97/n2340 ) );
  OAI22X1 \mult_97/U2167  ( .A(\mult_97/n2865 ), .B(n311), .C(\mult_97/n2866 ), 
        .D(n244), .Y(\mult_97/n2339 ) );
  OAI22X1 \mult_97/U2166  ( .A(\mult_97/n2864 ), .B(n311), .C(\mult_97/n2865 ), 
        .D(n244), .Y(\mult_97/n2338 ) );
  OAI22X1 \mult_97/U2165  ( .A(\mult_97/n2863 ), .B(n311), .C(\mult_97/n2864 ), 
        .D(n244), .Y(\mult_97/n2337 ) );
  OAI22X1 \mult_97/U2164  ( .A(\mult_97/n2862 ), .B(n311), .C(\mult_97/n2863 ), 
        .D(n244), .Y(\mult_97/n2336 ) );
  OAI22X1 \mult_97/U2163  ( .A(\mult_97/n2861 ), .B(n311), .C(\mult_97/n2862 ), 
        .D(n244), .Y(\mult_97/n2335 ) );
  OAI22X1 \mult_97/U2162  ( .A(\mult_97/n2860 ), .B(n311), .C(\mult_97/n2861 ), 
        .D(n244), .Y(\mult_97/n2334 ) );
  OAI22X1 \mult_97/U2161  ( .A(\mult_97/n2859 ), .B(n311), .C(\mult_97/n2860 ), 
        .D(n244), .Y(\mult_97/n2333 ) );
  OAI22X1 \mult_97/U2160  ( .A(\mult_97/n2858 ), .B(n311), .C(\mult_97/n2859 ), 
        .D(n244), .Y(\mult_97/n2332 ) );
  OAI22X1 \mult_97/U2159  ( .A(\mult_97/n2857 ), .B(n310), .C(\mult_97/n2858 ), 
        .D(n244), .Y(\mult_97/n2331 ) );
  OAI22X1 \mult_97/U2158  ( .A(\mult_97/n2856 ), .B(n310), .C(\mult_97/n2857 ), 
        .D(n244), .Y(\mult_97/n2330 ) );
  OAI22X1 \mult_97/U2157  ( .A(\mult_97/n2855 ), .B(n310), .C(\mult_97/n2856 ), 
        .D(n244), .Y(\mult_97/n2329 ) );
  OAI22X1 \mult_97/U2156  ( .A(\mult_97/n2854 ), .B(n310), .C(\mult_97/n2855 ), 
        .D(n244), .Y(\mult_97/n2328 ) );
  OAI22X1 \mult_97/U2155  ( .A(\mult_97/n2853 ), .B(n310), .C(\mult_97/n2854 ), 
        .D(n244), .Y(\mult_97/n2327 ) );
  OAI22X1 \mult_97/U2154  ( .A(\mult_97/n2852 ), .B(n310), .C(\mult_97/n2853 ), 
        .D(n244), .Y(\mult_97/n2326 ) );
  OAI22X1 \mult_97/U2153  ( .A(\mult_97/n2851 ), .B(n310), .C(\mult_97/n2852 ), 
        .D(n244), .Y(\mult_97/n2325 ) );
  OAI22X1 \mult_97/U2152  ( .A(\mult_97/n2850 ), .B(n311), .C(\mult_97/n2851 ), 
        .D(n244), .Y(\mult_97/n2324 ) );
  OAI22X1 \mult_97/U2151  ( .A(\mult_97/n2849 ), .B(n311), .C(\mult_97/n2850 ), 
        .D(n244), .Y(\mult_97/n2323 ) );
  OAI22X1 \mult_97/U2150  ( .A(\mult_97/n2848 ), .B(n311), .C(\mult_97/n2849 ), 
        .D(n244), .Y(\mult_97/n2322 ) );
  OAI22X1 \mult_97/U2149  ( .A(\mult_97/n2847 ), .B(n311), .C(\mult_97/n2848 ), 
        .D(n244), .Y(\mult_97/n2321 ) );
  OAI22X1 \mult_97/U2148  ( .A(\mult_97/n2846 ), .B(n311), .C(\mult_97/n2847 ), 
        .D(n244), .Y(\mult_97/n2320 ) );
  OAI22X1 \mult_97/U2147  ( .A(\mult_97/n2845 ), .B(n311), .C(\mult_97/n2846 ), 
        .D(n244), .Y(\mult_97/n2319 ) );
  OAI22X1 \mult_97/U2146  ( .A(\mult_97/n2844 ), .B(n311), .C(\mult_97/n2845 ), 
        .D(n244), .Y(\mult_97/n2318 ) );
  OAI22X1 \mult_97/U2145  ( .A(\mult_97/n2843 ), .B(n311), .C(\mult_97/n2844 ), 
        .D(n244), .Y(\mult_97/n2317 ) );
  OAI22X1 \mult_97/U2144  ( .A(\mult_97/n2842 ), .B(n311), .C(\mult_97/n2843 ), 
        .D(n244), .Y(\mult_97/n2316 ) );
  OAI22X1 \mult_97/U2143  ( .A(\mult_97/n2841 ), .B(n311), .C(\mult_97/n2842 ), 
        .D(n244), .Y(\mult_97/n2315 ) );
  OAI22X1 \mult_97/U2142  ( .A(n310), .B(\mult_97/n2873 ), .C(n303), .D(n244), 
        .Y(\mult_97/n1865 ) );
  XNOR2X1 \mult_97/U2141  ( .A(n302), .B(n251), .Y(\mult_97/n2839 ) );
  XNOR2X1 \mult_97/U2140  ( .A(n302), .B(n400), .Y(\mult_97/n2838 ) );
  XNOR2X1 \mult_97/U2139  ( .A(n302), .B(n398), .Y(\mult_97/n2837 ) );
  XNOR2X1 \mult_97/U2138  ( .A(n302), .B(n396), .Y(\mult_97/n2836 ) );
  XNOR2X1 \mult_97/U2137  ( .A(n302), .B(n394), .Y(\mult_97/n2835 ) );
  XNOR2X1 \mult_97/U2136  ( .A(n302), .B(n392), .Y(\mult_97/n2834 ) );
  XNOR2X1 \mult_97/U2135  ( .A(n302), .B(n390), .Y(\mult_97/n2833 ) );
  XNOR2X1 \mult_97/U2134  ( .A(n302), .B(n388), .Y(\mult_97/n2832 ) );
  XNOR2X1 \mult_97/U2133  ( .A(n302), .B(n386), .Y(\mult_97/n2831 ) );
  XNOR2X1 \mult_97/U2132  ( .A(n302), .B(n384), .Y(\mult_97/n2830 ) );
  XNOR2X1 \mult_97/U2131  ( .A(n302), .B(n382), .Y(\mult_97/n2829 ) );
  XNOR2X1 \mult_97/U2130  ( .A(n302), .B(n380), .Y(\mult_97/n2828 ) );
  XNOR2X1 \mult_97/U2129  ( .A(n302), .B(n378), .Y(\mult_97/n2827 ) );
  XNOR2X1 \mult_97/U2128  ( .A(n302), .B(n376), .Y(\mult_97/n2826 ) );
  XNOR2X1 \mult_97/U2127  ( .A(n302), .B(n374), .Y(\mult_97/n2825 ) );
  XNOR2X1 \mult_97/U2126  ( .A(n302), .B(n372), .Y(\mult_97/n2824 ) );
  XNOR2X1 \mult_97/U2125  ( .A(n302), .B(n370), .Y(\mult_97/n2823 ) );
  XNOR2X1 \mult_97/U2124  ( .A(n302), .B(n368), .Y(\mult_97/n2822 ) );
  XNOR2X1 \mult_97/U2123  ( .A(n302), .B(n366), .Y(\mult_97/n2821 ) );
  XNOR2X1 \mult_97/U2122  ( .A(n302), .B(n364), .Y(\mult_97/n2820 ) );
  XNOR2X1 \mult_97/U2121  ( .A(n302), .B(n362), .Y(\mult_97/n2819 ) );
  XNOR2X1 \mult_97/U2120  ( .A(n302), .B(n360), .Y(\mult_97/n2818 ) );
  XNOR2X1 \mult_97/U2119  ( .A(n302), .B(n358), .Y(\mult_97/n2817 ) );
  XNOR2X1 \mult_97/U2118  ( .A(n302), .B(n356), .Y(\mult_97/n2816 ) );
  XNOR2X1 \mult_97/U2117  ( .A(n302), .B(n354), .Y(\mult_97/n2815 ) );
  XNOR2X1 \mult_97/U2116  ( .A(n302), .B(n352), .Y(\mult_97/n2814 ) );
  XNOR2X1 \mult_97/U2115  ( .A(n302), .B(n350), .Y(\mult_97/n2813 ) );
  XNOR2X1 \mult_97/U2114  ( .A(n302), .B(n348), .Y(\mult_97/n2812 ) );
  XNOR2X1 \mult_97/U2113  ( .A(n302), .B(n346), .Y(\mult_97/n2811 ) );
  XNOR2X1 \mult_97/U2112  ( .A(n302), .B(n344), .Y(\mult_97/n2810 ) );
  XNOR2X1 \mult_97/U2111  ( .A(n302), .B(n342), .Y(\mult_97/n2809 ) );
  XNOR2X1 \mult_97/U2110  ( .A(n302), .B(n340), .Y(\mult_97/n2808 ) );
  OAI22X1 \mult_97/U2109  ( .A(n313), .B(\mult_97/n2838 ), .C(\mult_97/n2839 ), 
        .D(n332), .Y(\mult_97/n2312 ) );
  OAI22X1 \mult_97/U2108  ( .A(n313), .B(\mult_97/n2837 ), .C(\mult_97/n2838 ), 
        .D(n332), .Y(\mult_97/n2311 ) );
  OAI22X1 \mult_97/U2107  ( .A(n313), .B(\mult_97/n2836 ), .C(\mult_97/n2837 ), 
        .D(n332), .Y(\mult_97/n2310 ) );
  OAI22X1 \mult_97/U2106  ( .A(n313), .B(\mult_97/n2835 ), .C(\mult_97/n2836 ), 
        .D(n332), .Y(\mult_97/n2309 ) );
  OAI22X1 \mult_97/U2105  ( .A(n313), .B(\mult_97/n2834 ), .C(\mult_97/n2835 ), 
        .D(n332), .Y(\mult_97/n2308 ) );
  OAI22X1 \mult_97/U2104  ( .A(n313), .B(\mult_97/n2833 ), .C(\mult_97/n2834 ), 
        .D(n332), .Y(\mult_97/n2307 ) );
  OAI22X1 \mult_97/U2103  ( .A(n313), .B(\mult_97/n2832 ), .C(\mult_97/n2833 ), 
        .D(n332), .Y(\mult_97/n2306 ) );
  OAI22X1 \mult_97/U2102  ( .A(n313), .B(\mult_97/n2831 ), .C(\mult_97/n2832 ), 
        .D(n332), .Y(\mult_97/n2305 ) );
  OAI22X1 \mult_97/U2101  ( .A(n313), .B(\mult_97/n2830 ), .C(\mult_97/n2831 ), 
        .D(n332), .Y(\mult_97/n2304 ) );
  OAI22X1 \mult_97/U2100  ( .A(n313), .B(\mult_97/n2829 ), .C(\mult_97/n2830 ), 
        .D(n332), .Y(\mult_97/n2303 ) );
  OAI22X1 \mult_97/U2099  ( .A(n313), .B(\mult_97/n2828 ), .C(\mult_97/n2829 ), 
        .D(n332), .Y(\mult_97/n2302 ) );
  OAI22X1 \mult_97/U2098  ( .A(n313), .B(\mult_97/n2827 ), .C(\mult_97/n2828 ), 
        .D(n332), .Y(\mult_97/n2301 ) );
  OAI22X1 \mult_97/U2097  ( .A(n313), .B(\mult_97/n2826 ), .C(\mult_97/n2827 ), 
        .D(n332), .Y(\mult_97/n2300 ) );
  OAI22X1 \mult_97/U2096  ( .A(\mult_97/n353 ), .B(\mult_97/n2825 ), .C(
        \mult_97/n2826 ), .D(n332), .Y(\mult_97/n2299 ) );
  OAI22X1 \mult_97/U2095  ( .A(n313), .B(\mult_97/n2824 ), .C(\mult_97/n2825 ), 
        .D(n332), .Y(\mult_97/n2298 ) );
  OAI22X1 \mult_97/U2094  ( .A(\mult_97/n353 ), .B(\mult_97/n2823 ), .C(
        \mult_97/n2824 ), .D(n332), .Y(\mult_97/n2297 ) );
  OAI22X1 \mult_97/U2093  ( .A(\mult_97/n353 ), .B(\mult_97/n2822 ), .C(
        \mult_97/n2823 ), .D(n332), .Y(\mult_97/n2296 ) );
  OAI22X1 \mult_97/U2092  ( .A(\mult_97/n353 ), .B(\mult_97/n2821 ), .C(
        \mult_97/n2822 ), .D(n332), .Y(\mult_97/n2295 ) );
  OAI22X1 \mult_97/U2091  ( .A(\mult_97/n353 ), .B(\mult_97/n2820 ), .C(
        \mult_97/n2821 ), .D(n332), .Y(\mult_97/n2294 ) );
  OAI22X1 \mult_97/U2090  ( .A(\mult_97/n353 ), .B(\mult_97/n2819 ), .C(
        \mult_97/n2820 ), .D(n332), .Y(\mult_97/n2293 ) );
  OAI22X1 \mult_97/U2089  ( .A(n313), .B(\mult_97/n2818 ), .C(\mult_97/n2819 ), 
        .D(n332), .Y(\mult_97/n2292 ) );
  OAI22X1 \mult_97/U2088  ( .A(n313), .B(\mult_97/n2817 ), .C(\mult_97/n2818 ), 
        .D(n332), .Y(\mult_97/n2291 ) );
  OAI22X1 \mult_97/U2087  ( .A(n313), .B(\mult_97/n2816 ), .C(\mult_97/n2817 ), 
        .D(n332), .Y(\mult_97/n2290 ) );
  OAI22X1 \mult_97/U2086  ( .A(n313), .B(\mult_97/n2815 ), .C(\mult_97/n2816 ), 
        .D(n332), .Y(\mult_97/n2289 ) );
  OAI22X1 \mult_97/U2085  ( .A(n313), .B(\mult_97/n2814 ), .C(\mult_97/n2815 ), 
        .D(n332), .Y(\mult_97/n2288 ) );
  OAI22X1 \mult_97/U2084  ( .A(n313), .B(\mult_97/n2813 ), .C(\mult_97/n2814 ), 
        .D(n332), .Y(\mult_97/n2287 ) );
  OAI22X1 \mult_97/U2083  ( .A(n313), .B(\mult_97/n2812 ), .C(\mult_97/n2813 ), 
        .D(n332), .Y(\mult_97/n2286 ) );
  OAI22X1 \mult_97/U2082  ( .A(n313), .B(\mult_97/n2811 ), .C(\mult_97/n2812 ), 
        .D(n332), .Y(\mult_97/n2285 ) );
  OAI22X1 \mult_97/U2081  ( .A(n313), .B(\mult_97/n2810 ), .C(\mult_97/n2811 ), 
        .D(n332), .Y(\mult_97/n2284 ) );
  OAI22X1 \mult_97/U2080  ( .A(n313), .B(\mult_97/n2809 ), .C(\mult_97/n2810 ), 
        .D(n332), .Y(\mult_97/n2283 ) );
  OAI22X1 \mult_97/U2079  ( .A(n313), .B(\mult_97/n2808 ), .C(\mult_97/n2809 ), 
        .D(n332), .Y(\mult_97/n2282 ) );
  OAI22X1 \mult_97/U2078  ( .A(n313), .B(\mult_97/n2840 ), .C(n301), .D(n332), 
        .Y(\mult_97/n1864 ) );
  XNOR2X1 \mult_97/U2077  ( .A(n251), .B(n300), .Y(\mult_97/n2806 ) );
  XNOR2X1 \mult_97/U2076  ( .A(n400), .B(n300), .Y(\mult_97/n2805 ) );
  XNOR2X1 \mult_97/U2075  ( .A(n398), .B(n300), .Y(\mult_97/n2804 ) );
  XNOR2X1 \mult_97/U2074  ( .A(n396), .B(n300), .Y(\mult_97/n2803 ) );
  XNOR2X1 \mult_97/U2073  ( .A(n394), .B(n300), .Y(\mult_97/n2802 ) );
  XNOR2X1 \mult_97/U2072  ( .A(n392), .B(n300), .Y(\mult_97/n2801 ) );
  XNOR2X1 \mult_97/U2071  ( .A(n390), .B(n300), .Y(\mult_97/n2800 ) );
  XNOR2X1 \mult_97/U2070  ( .A(n388), .B(n300), .Y(\mult_97/n2799 ) );
  XNOR2X1 \mult_97/U2069  ( .A(n386), .B(n299), .Y(\mult_97/n2798 ) );
  XNOR2X1 \mult_97/U2068  ( .A(n384), .B(n300), .Y(\mult_97/n2797 ) );
  XNOR2X1 \mult_97/U2067  ( .A(n382), .B(n300), .Y(\mult_97/n2796 ) );
  XNOR2X1 \mult_97/U2066  ( .A(n380), .B(n299), .Y(\mult_97/n2795 ) );
  XNOR2X1 \mult_97/U2065  ( .A(n378), .B(n299), .Y(\mult_97/n2794 ) );
  XNOR2X1 \mult_97/U2064  ( .A(n376), .B(n299), .Y(\mult_97/n2793 ) );
  XNOR2X1 \mult_97/U2063  ( .A(B[14]), .B(n299), .Y(\mult_97/n2792 ) );
  XNOR2X1 \mult_97/U2062  ( .A(n372), .B(n299), .Y(\mult_97/n2791 ) );
  XNOR2X1 \mult_97/U2061  ( .A(n370), .B(n299), .Y(\mult_97/n2790 ) );
  XNOR2X1 \mult_97/U2060  ( .A(n368), .B(n299), .Y(\mult_97/n2789 ) );
  XNOR2X1 \mult_97/U2059  ( .A(n366), .B(n299), .Y(\mult_97/n2788 ) );
  XNOR2X1 \mult_97/U2058  ( .A(n364), .B(n299), .Y(\mult_97/n2787 ) );
  XNOR2X1 \mult_97/U2057  ( .A(n362), .B(n299), .Y(\mult_97/n2786 ) );
  XNOR2X1 \mult_97/U2056  ( .A(n360), .B(n299), .Y(\mult_97/n2785 ) );
  XNOR2X1 \mult_97/U2055  ( .A(n358), .B(n299), .Y(\mult_97/n2784 ) );
  XNOR2X1 \mult_97/U2054  ( .A(n356), .B(n299), .Y(\mult_97/n2783 ) );
  XNOR2X1 \mult_97/U2053  ( .A(n354), .B(n299), .Y(\mult_97/n2782 ) );
  XNOR2X1 \mult_97/U2052  ( .A(n352), .B(n299), .Y(\mult_97/n2781 ) );
  XNOR2X1 \mult_97/U2051  ( .A(n350), .B(n299), .Y(\mult_97/n2780 ) );
  XNOR2X1 \mult_97/U2050  ( .A(n348), .B(n299), .Y(\mult_97/n2779 ) );
  XNOR2X1 \mult_97/U2049  ( .A(n346), .B(n299), .Y(\mult_97/n2778 ) );
  XNOR2X1 \mult_97/U2048  ( .A(n344), .B(n299), .Y(\mult_97/n2777 ) );
  XNOR2X1 \mult_97/U2047  ( .A(n342), .B(n299), .Y(\mult_97/n2776 ) );
  XNOR2X1 \mult_97/U2046  ( .A(n340), .B(n300), .Y(\mult_97/n2775 ) );
  OAI22X1 \mult_97/U2045  ( .A(\mult_97/n2805 ), .B(n314), .C(\mult_97/n2806 ), 
        .D(n245), .Y(\mult_97/n2279 ) );
  OAI22X1 \mult_97/U2044  ( .A(\mult_97/n2804 ), .B(n314), .C(\mult_97/n2805 ), 
        .D(n245), .Y(\mult_97/n2278 ) );
  OAI22X1 \mult_97/U2043  ( .A(\mult_97/n2803 ), .B(n314), .C(\mult_97/n2804 ), 
        .D(n245), .Y(\mult_97/n2277 ) );
  OAI22X1 \mult_97/U2042  ( .A(\mult_97/n2802 ), .B(n314), .C(\mult_97/n2803 ), 
        .D(n245), .Y(\mult_97/n2276 ) );
  OAI22X1 \mult_97/U2041  ( .A(\mult_97/n2801 ), .B(n314), .C(\mult_97/n2802 ), 
        .D(n245), .Y(\mult_97/n2275 ) );
  OAI22X1 \mult_97/U2040  ( .A(\mult_97/n2800 ), .B(n314), .C(\mult_97/n2801 ), 
        .D(n245), .Y(\mult_97/n2274 ) );
  OAI22X1 \mult_97/U2039  ( .A(\mult_97/n2799 ), .B(n314), .C(\mult_97/n2800 ), 
        .D(n245), .Y(\mult_97/n2273 ) );
  OAI22X1 \mult_97/U2038  ( .A(\mult_97/n2798 ), .B(n314), .C(\mult_97/n2799 ), 
        .D(n245), .Y(\mult_97/n2272 ) );
  OAI22X1 \mult_97/U2037  ( .A(\mult_97/n2797 ), .B(n314), .C(\mult_97/n2798 ), 
        .D(n245), .Y(\mult_97/n2271 ) );
  OAI22X1 \mult_97/U2036  ( .A(\mult_97/n2796 ), .B(n314), .C(\mult_97/n2797 ), 
        .D(n245), .Y(\mult_97/n2270 ) );
  OAI22X1 \mult_97/U2035  ( .A(\mult_97/n2795 ), .B(n314), .C(\mult_97/n2796 ), 
        .D(n245), .Y(\mult_97/n2269 ) );
  OAI22X1 \mult_97/U2034  ( .A(\mult_97/n2794 ), .B(n314), .C(\mult_97/n2795 ), 
        .D(n245), .Y(\mult_97/n2268 ) );
  OAI22X1 \mult_97/U2033  ( .A(\mult_97/n2793 ), .B(n314), .C(\mult_97/n2794 ), 
        .D(n245), .Y(\mult_97/n2267 ) );
  OAI22X1 \mult_97/U2032  ( .A(\mult_97/n2792 ), .B(n314), .C(\mult_97/n2793 ), 
        .D(n245), .Y(\mult_97/n2266 ) );
  OAI22X1 \mult_97/U2031  ( .A(\mult_97/n2791 ), .B(n314), .C(\mult_97/n2792 ), 
        .D(n245), .Y(\mult_97/n2265 ) );
  OAI22X1 \mult_97/U2030  ( .A(\mult_97/n2790 ), .B(n314), .C(\mult_97/n2791 ), 
        .D(n245), .Y(\mult_97/n2264 ) );
  OAI22X1 \mult_97/U2029  ( .A(\mult_97/n2789 ), .B(n314), .C(\mult_97/n2790 ), 
        .D(n245), .Y(\mult_97/n2263 ) );
  OAI22X1 \mult_97/U2028  ( .A(\mult_97/n2788 ), .B(n314), .C(\mult_97/n2789 ), 
        .D(n245), .Y(\mult_97/n2262 ) );
  OAI22X1 \mult_97/U2027  ( .A(\mult_97/n2787 ), .B(n314), .C(\mult_97/n2788 ), 
        .D(n245), .Y(\mult_97/n2261 ) );
  OAI22X1 \mult_97/U2026  ( .A(\mult_97/n2786 ), .B(n314), .C(\mult_97/n2787 ), 
        .D(n245), .Y(\mult_97/n2260 ) );
  OAI22X1 \mult_97/U2025  ( .A(\mult_97/n2785 ), .B(n314), .C(\mult_97/n2786 ), 
        .D(n245), .Y(\mult_97/n2259 ) );
  OAI22X1 \mult_97/U2024  ( .A(\mult_97/n2784 ), .B(n314), .C(\mult_97/n2785 ), 
        .D(n245), .Y(\mult_97/n2258 ) );
  OAI22X1 \mult_97/U2023  ( .A(\mult_97/n2783 ), .B(n314), .C(\mult_97/n2784 ), 
        .D(n245), .Y(\mult_97/n2257 ) );
  OAI22X1 \mult_97/U2022  ( .A(\mult_97/n2782 ), .B(n314), .C(\mult_97/n2783 ), 
        .D(n245), .Y(\mult_97/n2256 ) );
  OAI22X1 \mult_97/U2021  ( .A(\mult_97/n2781 ), .B(n314), .C(\mult_97/n2782 ), 
        .D(n245), .Y(\mult_97/n2255 ) );
  OAI22X1 \mult_97/U2020  ( .A(\mult_97/n2780 ), .B(n314), .C(\mult_97/n2781 ), 
        .D(n245), .Y(\mult_97/n2254 ) );
  OAI22X1 \mult_97/U2019  ( .A(\mult_97/n2779 ), .B(n314), .C(\mult_97/n2780 ), 
        .D(n245), .Y(\mult_97/n1369 ) );
  OAI22X1 \mult_97/U2018  ( .A(\mult_97/n2778 ), .B(n314), .C(\mult_97/n2779 ), 
        .D(n245), .Y(\mult_97/n2253 ) );
  OAI22X1 \mult_97/U2017  ( .A(\mult_97/n2777 ), .B(n314), .C(\mult_97/n2778 ), 
        .D(n245), .Y(\mult_97/n2252 ) );
  OAI22X1 \mult_97/U2016  ( .A(\mult_97/n2776 ), .B(n314), .C(\mult_97/n2777 ), 
        .D(n245), .Y(\mult_97/n2251 ) );
  OAI22X1 \mult_97/U2015  ( .A(\mult_97/n2775 ), .B(n314), .C(\mult_97/n2776 ), 
        .D(n245), .Y(\mult_97/n1257 ) );
  OAI22X1 \mult_97/U2014  ( .A(n314), .B(\mult_97/n2807 ), .C(n298), .D(n245), 
        .Y(\mult_97/n1863 ) );
  XNOR2X1 \mult_97/U2013  ( .A(n251), .B(n297), .Y(\mult_97/n2773 ) );
  XNOR2X1 \mult_97/U2012  ( .A(B[1]), .B(n297), .Y(\mult_97/n2772 ) );
  XNOR2X1 \mult_97/U2011  ( .A(B[2]), .B(n297), .Y(\mult_97/n2771 ) );
  XNOR2X1 \mult_97/U2010  ( .A(B[3]), .B(n297), .Y(\mult_97/n2770 ) );
  XNOR2X1 \mult_97/U2009  ( .A(n394), .B(n297), .Y(\mult_97/n2769 ) );
  XNOR2X1 \mult_97/U2008  ( .A(n392), .B(n297), .Y(\mult_97/n2768 ) );
  XNOR2X1 \mult_97/U2007  ( .A(n390), .B(n297), .Y(\mult_97/n2767 ) );
  XNOR2X1 \mult_97/U2006  ( .A(n388), .B(n297), .Y(\mult_97/n2766 ) );
  XNOR2X1 \mult_97/U2005  ( .A(n386), .B(n296), .Y(\mult_97/n2765 ) );
  XNOR2X1 \mult_97/U2004  ( .A(n384), .B(n297), .Y(\mult_97/n2764 ) );
  XNOR2X1 \mult_97/U2003  ( .A(n382), .B(n297), .Y(\mult_97/n2763 ) );
  XNOR2X1 \mult_97/U2002  ( .A(n380), .B(n296), .Y(\mult_97/n2762 ) );
  XNOR2X1 \mult_97/U2001  ( .A(B[12]), .B(n296), .Y(\mult_97/n2761 ) );
  XNOR2X1 \mult_97/U2000  ( .A(B[13]), .B(n296), .Y(\mult_97/n2760 ) );
  XNOR2X1 \mult_97/U1999  ( .A(n374), .B(n296), .Y(\mult_97/n2759 ) );
  XNOR2X1 \mult_97/U1998  ( .A(n372), .B(n296), .Y(\mult_97/n2758 ) );
  XNOR2X1 \mult_97/U1997  ( .A(n370), .B(n296), .Y(\mult_97/n2757 ) );
  XNOR2X1 \mult_97/U1996  ( .A(n368), .B(n296), .Y(\mult_97/n2756 ) );
  XNOR2X1 \mult_97/U1995  ( .A(n366), .B(n296), .Y(\mult_97/n2755 ) );
  XNOR2X1 \mult_97/U1994  ( .A(n364), .B(n296), .Y(\mult_97/n2754 ) );
  XNOR2X1 \mult_97/U1993  ( .A(n362), .B(n296), .Y(\mult_97/n2753 ) );
  XNOR2X1 \mult_97/U1992  ( .A(n360), .B(n296), .Y(\mult_97/n2752 ) );
  XNOR2X1 \mult_97/U1991  ( .A(n358), .B(n296), .Y(\mult_97/n2751 ) );
  XNOR2X1 \mult_97/U1990  ( .A(n356), .B(n296), .Y(\mult_97/n2750 ) );
  XNOR2X1 \mult_97/U1989  ( .A(n354), .B(n296), .Y(\mult_97/n2749 ) );
  XNOR2X1 \mult_97/U1988  ( .A(n352), .B(n296), .Y(\mult_97/n2748 ) );
  XNOR2X1 \mult_97/U1987  ( .A(n350), .B(n296), .Y(\mult_97/n2747 ) );
  XNOR2X1 \mult_97/U1986  ( .A(n348), .B(n296), .Y(\mult_97/n2746 ) );
  XNOR2X1 \mult_97/U1985  ( .A(n346), .B(n296), .Y(\mult_97/n2745 ) );
  XNOR2X1 \mult_97/U1984  ( .A(n344), .B(n296), .Y(\mult_97/n2744 ) );
  XNOR2X1 \mult_97/U1983  ( .A(n342), .B(n296), .Y(\mult_97/n2743 ) );
  XNOR2X1 \mult_97/U1982  ( .A(n340), .B(n297), .Y(\mult_97/n2742 ) );
  OAI22X1 \mult_97/U1981  ( .A(\mult_97/n2772 ), .B(n316), .C(\mult_97/n2773 ), 
        .D(n333), .Y(\mult_97/n2248 ) );
  OAI22X1 \mult_97/U1980  ( .A(\mult_97/n2771 ), .B(n316), .C(\mult_97/n2772 ), 
        .D(n333), .Y(\mult_97/n2247 ) );
  OAI22X1 \mult_97/U1979  ( .A(\mult_97/n2770 ), .B(n316), .C(\mult_97/n2771 ), 
        .D(n333), .Y(\mult_97/n2246 ) );
  OAI22X1 \mult_97/U1978  ( .A(\mult_97/n2769 ), .B(n316), .C(\mult_97/n2770 ), 
        .D(n333), .Y(\mult_97/n2245 ) );
  OAI22X1 \mult_97/U1977  ( .A(\mult_97/n2768 ), .B(n316), .C(\mult_97/n2769 ), 
        .D(n333), .Y(\mult_97/n2244 ) );
  OAI22X1 \mult_97/U1976  ( .A(\mult_97/n2767 ), .B(n316), .C(\mult_97/n2768 ), 
        .D(n333), .Y(\mult_97/n2243 ) );
  OAI22X1 \mult_97/U1975  ( .A(\mult_97/n2766 ), .B(n316), .C(\mult_97/n2767 ), 
        .D(n333), .Y(\mult_97/n2242 ) );
  OAI22X1 \mult_97/U1974  ( .A(\mult_97/n2765 ), .B(n316), .C(\mult_97/n2766 ), 
        .D(n333), .Y(\mult_97/n2241 ) );
  OAI22X1 \mult_97/U1973  ( .A(\mult_97/n2764 ), .B(n316), .C(\mult_97/n2765 ), 
        .D(n333), .Y(\mult_97/n2240 ) );
  OAI22X1 \mult_97/U1972  ( .A(\mult_97/n2763 ), .B(n316), .C(\mult_97/n2764 ), 
        .D(n333), .Y(\mult_97/n2239 ) );
  OAI22X1 \mult_97/U1971  ( .A(\mult_97/n2762 ), .B(n316), .C(\mult_97/n2763 ), 
        .D(n333), .Y(\mult_97/n2238 ) );
  OAI22X1 \mult_97/U1970  ( .A(\mult_97/n2761 ), .B(n316), .C(\mult_97/n2762 ), 
        .D(n333), .Y(\mult_97/n2237 ) );
  OAI22X1 \mult_97/U1969  ( .A(\mult_97/n2760 ), .B(n316), .C(\mult_97/n2761 ), 
        .D(n333), .Y(\mult_97/n2236 ) );
  OAI22X1 \mult_97/U1968  ( .A(\mult_97/n2759 ), .B(n316), .C(\mult_97/n2760 ), 
        .D(n333), .Y(\mult_97/n2235 ) );
  OAI22X1 \mult_97/U1967  ( .A(\mult_97/n2758 ), .B(n315), .C(\mult_97/n2759 ), 
        .D(n333), .Y(\mult_97/n2234 ) );
  OAI22X1 \mult_97/U1966  ( .A(\mult_97/n2757 ), .B(n315), .C(\mult_97/n2758 ), 
        .D(n333), .Y(\mult_97/n2233 ) );
  OAI22X1 \mult_97/U1965  ( .A(\mult_97/n2756 ), .B(n315), .C(\mult_97/n2757 ), 
        .D(n333), .Y(\mult_97/n2232 ) );
  OAI22X1 \mult_97/U1964  ( .A(\mult_97/n2755 ), .B(n315), .C(\mult_97/n2756 ), 
        .D(n333), .Y(\mult_97/n2231 ) );
  OAI22X1 \mult_97/U1963  ( .A(\mult_97/n2754 ), .B(n315), .C(\mult_97/n2755 ), 
        .D(n333), .Y(\mult_97/n2230 ) );
  OAI22X1 \mult_97/U1962  ( .A(\mult_97/n2753 ), .B(n315), .C(\mult_97/n2754 ), 
        .D(n333), .Y(\mult_97/n2229 ) );
  OAI22X1 \mult_97/U1961  ( .A(\mult_97/n2752 ), .B(n315), .C(\mult_97/n2753 ), 
        .D(n333), .Y(\mult_97/n2228 ) );
  OAI22X1 \mult_97/U1960  ( .A(\mult_97/n2751 ), .B(n316), .C(\mult_97/n2752 ), 
        .D(n333), .Y(\mult_97/n2227 ) );
  OAI22X1 \mult_97/U1959  ( .A(\mult_97/n2750 ), .B(n316), .C(\mult_97/n2751 ), 
        .D(n333), .Y(\mult_97/n2226 ) );
  OAI22X1 \mult_97/U1958  ( .A(\mult_97/n2749 ), .B(n316), .C(\mult_97/n2750 ), 
        .D(n333), .Y(\mult_97/n2225 ) );
  OAI22X1 \mult_97/U1957  ( .A(\mult_97/n2748 ), .B(n316), .C(\mult_97/n2749 ), 
        .D(n333), .Y(\mult_97/n2224 ) );
  OAI22X1 \mult_97/U1956  ( .A(\mult_97/n2747 ), .B(n316), .C(\mult_97/n2748 ), 
        .D(n333), .Y(\mult_97/n2223 ) );
  OAI22X1 \mult_97/U1955  ( .A(\mult_97/n2746 ), .B(n316), .C(\mult_97/n2747 ), 
        .D(n333), .Y(\mult_97/n2222 ) );
  OAI22X1 \mult_97/U1954  ( .A(\mult_97/n2745 ), .B(n316), .C(\mult_97/n2746 ), 
        .D(n333), .Y(\mult_97/n2221 ) );
  OAI22X1 \mult_97/U1953  ( .A(\mult_97/n2744 ), .B(n316), .C(\mult_97/n2745 ), 
        .D(n333), .Y(\mult_97/n2220 ) );
  OAI22X1 \mult_97/U1952  ( .A(\mult_97/n2743 ), .B(n316), .C(\mult_97/n2744 ), 
        .D(n333), .Y(\mult_97/n2219 ) );
  OAI22X1 \mult_97/U1951  ( .A(\mult_97/n2742 ), .B(n316), .C(\mult_97/n2743 ), 
        .D(n333), .Y(\mult_97/n2218 ) );
  OAI22X1 \mult_97/U1950  ( .A(n315), .B(\mult_97/n2774 ), .C(n295), .D(n333), 
        .Y(\mult_97/n1862 ) );
  XNOR2X1 \mult_97/U1949  ( .A(n294), .B(n251), .Y(\mult_97/n2740 ) );
  XNOR2X1 \mult_97/U1948  ( .A(n294), .B(n400), .Y(\mult_97/n2739 ) );
  XNOR2X1 \mult_97/U1947  ( .A(n294), .B(n398), .Y(\mult_97/n2738 ) );
  XNOR2X1 \mult_97/U1946  ( .A(n294), .B(n396), .Y(\mult_97/n2737 ) );
  XNOR2X1 \mult_97/U1945  ( .A(n294), .B(n394), .Y(\mult_97/n2736 ) );
  XNOR2X1 \mult_97/U1944  ( .A(n294), .B(n392), .Y(\mult_97/n2735 ) );
  XNOR2X1 \mult_97/U1943  ( .A(n294), .B(n390), .Y(\mult_97/n2734 ) );
  XNOR2X1 \mult_97/U1942  ( .A(n294), .B(n388), .Y(\mult_97/n2733 ) );
  XNOR2X1 \mult_97/U1941  ( .A(n294), .B(n386), .Y(\mult_97/n2732 ) );
  XNOR2X1 \mult_97/U1940  ( .A(n294), .B(n384), .Y(\mult_97/n2731 ) );
  XNOR2X1 \mult_97/U1939  ( .A(n294), .B(n382), .Y(\mult_97/n2730 ) );
  XNOR2X1 \mult_97/U1938  ( .A(n294), .B(n380), .Y(\mult_97/n2729 ) );
  XNOR2X1 \mult_97/U1937  ( .A(n294), .B(n378), .Y(\mult_97/n2728 ) );
  XNOR2X1 \mult_97/U1936  ( .A(n294), .B(n376), .Y(\mult_97/n2727 ) );
  XNOR2X1 \mult_97/U1935  ( .A(n294), .B(n374), .Y(\mult_97/n2726 ) );
  XNOR2X1 \mult_97/U1934  ( .A(n294), .B(n372), .Y(\mult_97/n2725 ) );
  XNOR2X1 \mult_97/U1933  ( .A(n294), .B(n370), .Y(\mult_97/n2724 ) );
  XNOR2X1 \mult_97/U1932  ( .A(n294), .B(n368), .Y(\mult_97/n2723 ) );
  XNOR2X1 \mult_97/U1931  ( .A(n294), .B(n366), .Y(\mult_97/n2722 ) );
  XNOR2X1 \mult_97/U1930  ( .A(n294), .B(n364), .Y(\mult_97/n2721 ) );
  XNOR2X1 \mult_97/U1929  ( .A(n294), .B(n362), .Y(\mult_97/n2720 ) );
  XNOR2X1 \mult_97/U1928  ( .A(n294), .B(n360), .Y(\mult_97/n2719 ) );
  XNOR2X1 \mult_97/U1927  ( .A(n294), .B(n358), .Y(\mult_97/n2718 ) );
  XNOR2X1 \mult_97/U1926  ( .A(n294), .B(n356), .Y(\mult_97/n2717 ) );
  XNOR2X1 \mult_97/U1925  ( .A(n294), .B(n354), .Y(\mult_97/n2716 ) );
  XNOR2X1 \mult_97/U1924  ( .A(n294), .B(n352), .Y(\mult_97/n2715 ) );
  XNOR2X1 \mult_97/U1923  ( .A(n294), .B(n350), .Y(\mult_97/n2714 ) );
  XNOR2X1 \mult_97/U1922  ( .A(n294), .B(n348), .Y(\mult_97/n2713 ) );
  XNOR2X1 \mult_97/U1921  ( .A(n294), .B(n346), .Y(\mult_97/n2712 ) );
  XNOR2X1 \mult_97/U1920  ( .A(n294), .B(n344), .Y(\mult_97/n2711 ) );
  XNOR2X1 \mult_97/U1919  ( .A(n294), .B(n342), .Y(\mult_97/n2710 ) );
  XNOR2X1 \mult_97/U1918  ( .A(n294), .B(n340), .Y(\mult_97/n2709 ) );
  OAI22X1 \mult_97/U1917  ( .A(n318), .B(\mult_97/n2739 ), .C(\mult_97/n2740 ), 
        .D(n243), .Y(\mult_97/n2215 ) );
  OAI22X1 \mult_97/U1916  ( .A(n318), .B(\mult_97/n2738 ), .C(\mult_97/n2739 ), 
        .D(n243), .Y(\mult_97/n2214 ) );
  OAI22X1 \mult_97/U1915  ( .A(n318), .B(\mult_97/n2737 ), .C(\mult_97/n2738 ), 
        .D(n243), .Y(\mult_97/n2213 ) );
  OAI22X1 \mult_97/U1914  ( .A(n318), .B(\mult_97/n2736 ), .C(\mult_97/n2737 ), 
        .D(n243), .Y(\mult_97/n2212 ) );
  OAI22X1 \mult_97/U1913  ( .A(n318), .B(\mult_97/n2735 ), .C(\mult_97/n2736 ), 
        .D(n243), .Y(\mult_97/n2211 ) );
  OAI22X1 \mult_97/U1912  ( .A(n318), .B(\mult_97/n2734 ), .C(\mult_97/n2735 ), 
        .D(n243), .Y(\mult_97/n2210 ) );
  OAI22X1 \mult_97/U1911  ( .A(n318), .B(\mult_97/n2733 ), .C(\mult_97/n2734 ), 
        .D(n243), .Y(\mult_97/n2209 ) );
  OAI22X1 \mult_97/U1910  ( .A(n318), .B(\mult_97/n2732 ), .C(\mult_97/n2733 ), 
        .D(n243), .Y(\mult_97/n2208 ) );
  OAI22X1 \mult_97/U1909  ( .A(n318), .B(\mult_97/n2731 ), .C(\mult_97/n2732 ), 
        .D(n243), .Y(\mult_97/n2207 ) );
  OAI22X1 \mult_97/U1908  ( .A(n318), .B(\mult_97/n2730 ), .C(\mult_97/n2731 ), 
        .D(n243), .Y(\mult_97/n2206 ) );
  OAI22X1 \mult_97/U1907  ( .A(n318), .B(\mult_97/n2729 ), .C(\mult_97/n2730 ), 
        .D(n243), .Y(\mult_97/n2205 ) );
  OAI22X1 \mult_97/U1906  ( .A(n318), .B(\mult_97/n2728 ), .C(\mult_97/n2729 ), 
        .D(n243), .Y(\mult_97/n2204 ) );
  OAI22X1 \mult_97/U1905  ( .A(n318), .B(\mult_97/n2727 ), .C(\mult_97/n2728 ), 
        .D(n243), .Y(\mult_97/n2203 ) );
  OAI22X1 \mult_97/U1904  ( .A(\mult_97/n362 ), .B(\mult_97/n2726 ), .C(
        \mult_97/n2727 ), .D(n243), .Y(\mult_97/n2202 ) );
  OAI22X1 \mult_97/U1903  ( .A(n318), .B(\mult_97/n2725 ), .C(\mult_97/n2726 ), 
        .D(n243), .Y(\mult_97/n2201 ) );
  OAI22X1 \mult_97/U1902  ( .A(\mult_97/n362 ), .B(\mult_97/n2724 ), .C(
        \mult_97/n2725 ), .D(n243), .Y(\mult_97/n2200 ) );
  OAI22X1 \mult_97/U1901  ( .A(n318), .B(\mult_97/n2723 ), .C(\mult_97/n2724 ), 
        .D(n243), .Y(\mult_97/n2199 ) );
  OAI22X1 \mult_97/U1900  ( .A(\mult_97/n362 ), .B(\mult_97/n2722 ), .C(
        \mult_97/n2723 ), .D(n243), .Y(\mult_97/n2198 ) );
  OAI22X1 \mult_97/U1899  ( .A(\mult_97/n362 ), .B(\mult_97/n2721 ), .C(
        \mult_97/n2722 ), .D(n243), .Y(\mult_97/n2197 ) );
  OAI22X1 \mult_97/U1898  ( .A(\mult_97/n362 ), .B(\mult_97/n2720 ), .C(
        \mult_97/n2721 ), .D(n243), .Y(\mult_97/n2196 ) );
  OAI22X1 \mult_97/U1897  ( .A(\mult_97/n362 ), .B(\mult_97/n2719 ), .C(
        \mult_97/n2720 ), .D(n243), .Y(\mult_97/n2195 ) );
  OAI22X1 \mult_97/U1896  ( .A(n318), .B(\mult_97/n2718 ), .C(\mult_97/n2719 ), 
        .D(n243), .Y(\mult_97/n2194 ) );
  OAI22X1 \mult_97/U1895  ( .A(n318), .B(\mult_97/n2717 ), .C(\mult_97/n2718 ), 
        .D(n243), .Y(\mult_97/n2193 ) );
  OAI22X1 \mult_97/U1894  ( .A(n318), .B(\mult_97/n2716 ), .C(\mult_97/n2717 ), 
        .D(n243), .Y(\mult_97/n2192 ) );
  OAI22X1 \mult_97/U1893  ( .A(n318), .B(\mult_97/n2715 ), .C(\mult_97/n2716 ), 
        .D(n243), .Y(\mult_97/n2191 ) );
  OAI22X1 \mult_97/U1892  ( .A(n318), .B(\mult_97/n2714 ), .C(\mult_97/n2715 ), 
        .D(n243), .Y(\mult_97/n2190 ) );
  OAI22X1 \mult_97/U1891  ( .A(n318), .B(\mult_97/n2713 ), .C(\mult_97/n2714 ), 
        .D(n243), .Y(\mult_97/n2189 ) );
  OAI22X1 \mult_97/U1890  ( .A(n318), .B(\mult_97/n2712 ), .C(\mult_97/n2713 ), 
        .D(n243), .Y(\mult_97/n2188 ) );
  OAI22X1 \mult_97/U1889  ( .A(n318), .B(\mult_97/n2711 ), .C(\mult_97/n2712 ), 
        .D(n243), .Y(\mult_97/n2187 ) );
  OAI22X1 \mult_97/U1888  ( .A(n318), .B(\mult_97/n2710 ), .C(\mult_97/n2711 ), 
        .D(n243), .Y(\mult_97/n2186 ) );
  OAI22X1 \mult_97/U1887  ( .A(n318), .B(\mult_97/n2709 ), .C(\mult_97/n2710 ), 
        .D(n243), .Y(\mult_97/n2185 ) );
  OAI22X1 \mult_97/U1886  ( .A(n318), .B(\mult_97/n2741 ), .C(n293), .D(n243), 
        .Y(\mult_97/n1861 ) );
  XNOR2X1 \mult_97/U1885  ( .A(n251), .B(n292), .Y(\mult_97/n2707 ) );
  XNOR2X1 \mult_97/U1884  ( .A(n400), .B(n292), .Y(\mult_97/n2706 ) );
  XNOR2X1 \mult_97/U1883  ( .A(n398), .B(n292), .Y(\mult_97/n2705 ) );
  XNOR2X1 \mult_97/U1882  ( .A(n396), .B(n292), .Y(\mult_97/n2704 ) );
  XNOR2X1 \mult_97/U1881  ( .A(n394), .B(n292), .Y(\mult_97/n2703 ) );
  XNOR2X1 \mult_97/U1880  ( .A(n392), .B(n292), .Y(\mult_97/n2702 ) );
  XNOR2X1 \mult_97/U1879  ( .A(n390), .B(n292), .Y(\mult_97/n2701 ) );
  XNOR2X1 \mult_97/U1878  ( .A(n388), .B(n292), .Y(\mult_97/n2700 ) );
  XNOR2X1 \mult_97/U1877  ( .A(B[8]), .B(n291), .Y(\mult_97/n2699 ) );
  XNOR2X1 \mult_97/U1876  ( .A(n384), .B(n292), .Y(\mult_97/n2698 ) );
  XNOR2X1 \mult_97/U1875  ( .A(n382), .B(n292), .Y(\mult_97/n2697 ) );
  XNOR2X1 \mult_97/U1874  ( .A(n380), .B(n291), .Y(\mult_97/n2696 ) );
  XNOR2X1 \mult_97/U1873  ( .A(n378), .B(n291), .Y(\mult_97/n2695 ) );
  XNOR2X1 \mult_97/U1872  ( .A(n376), .B(n291), .Y(\mult_97/n2694 ) );
  XNOR2X1 \mult_97/U1871  ( .A(n374), .B(n291), .Y(\mult_97/n2693 ) );
  XNOR2X1 \mult_97/U1870  ( .A(n372), .B(n291), .Y(\mult_97/n2692 ) );
  XNOR2X1 \mult_97/U1869  ( .A(n370), .B(n291), .Y(\mult_97/n2691 ) );
  XNOR2X1 \mult_97/U1868  ( .A(n368), .B(n291), .Y(\mult_97/n2690 ) );
  XNOR2X1 \mult_97/U1867  ( .A(n366), .B(n291), .Y(\mult_97/n2689 ) );
  XNOR2X1 \mult_97/U1866  ( .A(n364), .B(n291), .Y(\mult_97/n2688 ) );
  XNOR2X1 \mult_97/U1865  ( .A(n362), .B(n291), .Y(\mult_97/n2687 ) );
  XNOR2X1 \mult_97/U1864  ( .A(n360), .B(n291), .Y(\mult_97/n2686 ) );
  XNOR2X1 \mult_97/U1863  ( .A(n358), .B(n291), .Y(\mult_97/n2685 ) );
  XNOR2X1 \mult_97/U1862  ( .A(n356), .B(n291), .Y(\mult_97/n2684 ) );
  XNOR2X1 \mult_97/U1861  ( .A(n354), .B(n291), .Y(\mult_97/n2683 ) );
  XNOR2X1 \mult_97/U1860  ( .A(n352), .B(n291), .Y(\mult_97/n2682 ) );
  XNOR2X1 \mult_97/U1859  ( .A(n350), .B(n291), .Y(\mult_97/n2681 ) );
  XNOR2X1 \mult_97/U1858  ( .A(n348), .B(n291), .Y(\mult_97/n2680 ) );
  XNOR2X1 \mult_97/U1857  ( .A(n346), .B(n291), .Y(\mult_97/n2679 ) );
  XNOR2X1 \mult_97/U1856  ( .A(n344), .B(n291), .Y(\mult_97/n2678 ) );
  XNOR2X1 \mult_97/U1855  ( .A(n342), .B(n291), .Y(\mult_97/n2677 ) );
  XNOR2X1 \mult_97/U1854  ( .A(n340), .B(n292), .Y(\mult_97/n2676 ) );
  OAI22X1 \mult_97/U1853  ( .A(\mult_97/n2706 ), .B(n319), .C(\mult_97/n2707 ), 
        .D(n249), .Y(\mult_97/n2182 ) );
  OAI22X1 \mult_97/U1852  ( .A(\mult_97/n2705 ), .B(n319), .C(\mult_97/n2706 ), 
        .D(n249), .Y(\mult_97/n2181 ) );
  OAI22X1 \mult_97/U1851  ( .A(\mult_97/n2704 ), .B(n319), .C(\mult_97/n2705 ), 
        .D(n249), .Y(\mult_97/n2180 ) );
  OAI22X1 \mult_97/U1850  ( .A(\mult_97/n2703 ), .B(n319), .C(\mult_97/n2704 ), 
        .D(n249), .Y(\mult_97/n2179 ) );
  OAI22X1 \mult_97/U1849  ( .A(\mult_97/n2702 ), .B(n319), .C(\mult_97/n2703 ), 
        .D(n249), .Y(\mult_97/n2178 ) );
  OAI22X1 \mult_97/U1848  ( .A(\mult_97/n2701 ), .B(n319), .C(\mult_97/n2702 ), 
        .D(n249), .Y(\mult_97/n2177 ) );
  OAI22X1 \mult_97/U1847  ( .A(\mult_97/n2700 ), .B(n319), .C(\mult_97/n2701 ), 
        .D(n249), .Y(\mult_97/n2176 ) );
  OAI22X1 \mult_97/U1846  ( .A(\mult_97/n2699 ), .B(n319), .C(\mult_97/n2700 ), 
        .D(n249), .Y(\mult_97/n2175 ) );
  OAI22X1 \mult_97/U1845  ( .A(\mult_97/n2698 ), .B(n319), .C(\mult_97/n2699 ), 
        .D(n249), .Y(\mult_97/n2174 ) );
  OAI22X1 \mult_97/U1844  ( .A(\mult_97/n2697 ), .B(n319), .C(\mult_97/n2698 ), 
        .D(n249), .Y(\mult_97/n2173 ) );
  OAI22X1 \mult_97/U1843  ( .A(\mult_97/n2696 ), .B(n319), .C(\mult_97/n2697 ), 
        .D(n249), .Y(\mult_97/n2172 ) );
  OAI22X1 \mult_97/U1842  ( .A(\mult_97/n2695 ), .B(n319), .C(\mult_97/n2696 ), 
        .D(n249), .Y(\mult_97/n2171 ) );
  OAI22X1 \mult_97/U1841  ( .A(\mult_97/n2694 ), .B(n319), .C(\mult_97/n2695 ), 
        .D(n249), .Y(\mult_97/n2170 ) );
  OAI22X1 \mult_97/U1840  ( .A(\mult_97/n2693 ), .B(n319), .C(\mult_97/n2694 ), 
        .D(n249), .Y(\mult_97/n2169 ) );
  OAI22X1 \mult_97/U1839  ( .A(\mult_97/n2692 ), .B(n319), .C(\mult_97/n2693 ), 
        .D(n249), .Y(\mult_97/n2168 ) );
  OAI22X1 \mult_97/U1838  ( .A(\mult_97/n2691 ), .B(n319), .C(\mult_97/n2692 ), 
        .D(n249), .Y(\mult_97/n2167 ) );
  OAI22X1 \mult_97/U1837  ( .A(\mult_97/n2690 ), .B(n319), .C(\mult_97/n2691 ), 
        .D(n249), .Y(\mult_97/n2166 ) );
  OAI22X1 \mult_97/U1836  ( .A(\mult_97/n2689 ), .B(n319), .C(\mult_97/n2690 ), 
        .D(n249), .Y(\mult_97/n2165 ) );
  OAI22X1 \mult_97/U1835  ( .A(\mult_97/n2688 ), .B(n319), .C(\mult_97/n2689 ), 
        .D(n249), .Y(\mult_97/n2164 ) );
  OAI22X1 \mult_97/U1834  ( .A(\mult_97/n2687 ), .B(n319), .C(\mult_97/n2688 ), 
        .D(n249), .Y(\mult_97/n2163 ) );
  OAI22X1 \mult_97/U1833  ( .A(\mult_97/n2686 ), .B(n319), .C(\mult_97/n2687 ), 
        .D(n249), .Y(\mult_97/n2162 ) );
  OAI22X1 \mult_97/U1832  ( .A(\mult_97/n2685 ), .B(n319), .C(\mult_97/n2686 ), 
        .D(n249), .Y(\mult_97/n2161 ) );
  OAI22X1 \mult_97/U1831  ( .A(\mult_97/n2684 ), .B(n319), .C(\mult_97/n2685 ), 
        .D(n249), .Y(\mult_97/n1311 ) );
  OAI22X1 \mult_97/U1830  ( .A(\mult_97/n2683 ), .B(n319), .C(\mult_97/n2684 ), 
        .D(n249), .Y(\mult_97/n2160 ) );
  OAI22X1 \mult_97/U1829  ( .A(\mult_97/n2682 ), .B(n319), .C(\mult_97/n2683 ), 
        .D(n249), .Y(\mult_97/n2159 ) );
  OAI22X1 \mult_97/U1828  ( .A(\mult_97/n2681 ), .B(n319), .C(\mult_97/n2682 ), 
        .D(n249), .Y(\mult_97/n2158 ) );
  OAI22X1 \mult_97/U1827  ( .A(\mult_97/n2680 ), .B(n319), .C(\mult_97/n2681 ), 
        .D(n249), .Y(\mult_97/n2157 ) );
  OAI22X1 \mult_97/U1826  ( .A(\mult_97/n2679 ), .B(n319), .C(\mult_97/n2680 ), 
        .D(n249), .Y(\mult_97/n2156 ) );
  OAI22X1 \mult_97/U1825  ( .A(\mult_97/n2678 ), .B(n319), .C(\mult_97/n2679 ), 
        .D(n249), .Y(\mult_97/n2155 ) );
  OAI22X1 \mult_97/U1824  ( .A(\mult_97/n2677 ), .B(n319), .C(\mult_97/n2678 ), 
        .D(n249), .Y(\mult_97/n2154 ) );
  OAI22X1 \mult_97/U1823  ( .A(\mult_97/n2676 ), .B(n319), .C(\mult_97/n2677 ), 
        .D(n249), .Y(\mult_97/n1119 ) );
  OAI22X1 \mult_97/U1822  ( .A(n319), .B(\mult_97/n2708 ), .C(n290), .D(n249), 
        .Y(\mult_97/n1860 ) );
  XNOR2X1 \mult_97/U1821  ( .A(n251), .B(A[15]), .Y(\mult_97/n2674 ) );
  XNOR2X1 \mult_97/U1820  ( .A(n400), .B(n289), .Y(\mult_97/n2673 ) );
  XNOR2X1 \mult_97/U1819  ( .A(n398), .B(n289), .Y(\mult_97/n2672 ) );
  XNOR2X1 \mult_97/U1818  ( .A(n396), .B(n289), .Y(\mult_97/n2671 ) );
  XNOR2X1 \mult_97/U1817  ( .A(n394), .B(n289), .Y(\mult_97/n2670 ) );
  XNOR2X1 \mult_97/U1816  ( .A(n392), .B(n289), .Y(\mult_97/n2669 ) );
  XNOR2X1 \mult_97/U1815  ( .A(B[6]), .B(n289), .Y(\mult_97/n2668 ) );
  XNOR2X1 \mult_97/U1814  ( .A(n388), .B(n289), .Y(\mult_97/n2667 ) );
  XNOR2X1 \mult_97/U1813  ( .A(n386), .B(n289), .Y(\mult_97/n2666 ) );
  XNOR2X1 \mult_97/U1812  ( .A(n384), .B(n289), .Y(\mult_97/n2665 ) );
  XNOR2X1 \mult_97/U1811  ( .A(n382), .B(n289), .Y(\mult_97/n2664 ) );
  XNOR2X1 \mult_97/U1810  ( .A(n380), .B(n289), .Y(\mult_97/n2663 ) );
  XNOR2X1 \mult_97/U1809  ( .A(n378), .B(n289), .Y(\mult_97/n2662 ) );
  XNOR2X1 \mult_97/U1808  ( .A(n376), .B(n289), .Y(\mult_97/n2661 ) );
  XNOR2X1 \mult_97/U1807  ( .A(n374), .B(n289), .Y(\mult_97/n2660 ) );
  XNOR2X1 \mult_97/U1806  ( .A(n372), .B(n289), .Y(\mult_97/n2659 ) );
  XNOR2X1 \mult_97/U1805  ( .A(n370), .B(n289), .Y(\mult_97/n2658 ) );
  XNOR2X1 \mult_97/U1804  ( .A(n368), .B(n289), .Y(\mult_97/n2657 ) );
  XNOR2X1 \mult_97/U1803  ( .A(n366), .B(n289), .Y(\mult_97/n2656 ) );
  XNOR2X1 \mult_97/U1802  ( .A(n364), .B(n289), .Y(\mult_97/n2655 ) );
  XNOR2X1 \mult_97/U1801  ( .A(B[20]), .B(n289), .Y(\mult_97/n2654 ) );
  XNOR2X1 \mult_97/U1800  ( .A(B[21]), .B(n289), .Y(\mult_97/n2653 ) );
  XNOR2X1 \mult_97/U1799  ( .A(n358), .B(n289), .Y(\mult_97/n2652 ) );
  XNOR2X1 \mult_97/U1798  ( .A(n356), .B(n289), .Y(\mult_97/n2651 ) );
  XNOR2X1 \mult_97/U1797  ( .A(n354), .B(n289), .Y(\mult_97/n2650 ) );
  XNOR2X1 \mult_97/U1796  ( .A(n352), .B(n289), .Y(\mult_97/n2649 ) );
  XNOR2X1 \mult_97/U1795  ( .A(n350), .B(n289), .Y(\mult_97/n2648 ) );
  XNOR2X1 \mult_97/U1794  ( .A(n348), .B(n289), .Y(\mult_97/n2647 ) );
  XNOR2X1 \mult_97/U1793  ( .A(n346), .B(n289), .Y(\mult_97/n2646 ) );
  XNOR2X1 \mult_97/U1792  ( .A(n344), .B(n289), .Y(\mult_97/n2645 ) );
  XNOR2X1 \mult_97/U1791  ( .A(n342), .B(n289), .Y(\mult_97/n2644 ) );
  XNOR2X1 \mult_97/U1790  ( .A(n340), .B(A[15]), .Y(\mult_97/n2643 ) );
  OAI22X1 \mult_97/U1789  ( .A(\mult_97/n2673 ), .B(n321), .C(\mult_97/n2674 ), 
        .D(n334), .Y(\mult_97/n2151 ) );
  OAI22X1 \mult_97/U1788  ( .A(\mult_97/n2672 ), .B(n321), .C(\mult_97/n2673 ), 
        .D(n334), .Y(\mult_97/n2150 ) );
  OAI22X1 \mult_97/U1787  ( .A(\mult_97/n2671 ), .B(n321), .C(\mult_97/n2672 ), 
        .D(n334), .Y(\mult_97/n2149 ) );
  OAI22X1 \mult_97/U1786  ( .A(\mult_97/n2670 ), .B(n321), .C(\mult_97/n2671 ), 
        .D(n334), .Y(\mult_97/n2148 ) );
  OAI22X1 \mult_97/U1785  ( .A(\mult_97/n2669 ), .B(n321), .C(\mult_97/n2670 ), 
        .D(n334), .Y(\mult_97/n2147 ) );
  OAI22X1 \mult_97/U1784  ( .A(\mult_97/n2668 ), .B(n321), .C(\mult_97/n2669 ), 
        .D(n334), .Y(\mult_97/n2146 ) );
  OAI22X1 \mult_97/U1783  ( .A(\mult_97/n2667 ), .B(n321), .C(\mult_97/n2668 ), 
        .D(n334), .Y(\mult_97/n2145 ) );
  OAI22X1 \mult_97/U1782  ( .A(\mult_97/n2666 ), .B(n321), .C(\mult_97/n2667 ), 
        .D(n334), .Y(\mult_97/n2144 ) );
  OAI22X1 \mult_97/U1781  ( .A(\mult_97/n2665 ), .B(n321), .C(\mult_97/n2666 ), 
        .D(n334), .Y(\mult_97/n2143 ) );
  OAI22X1 \mult_97/U1780  ( .A(\mult_97/n2664 ), .B(n321), .C(\mult_97/n2665 ), 
        .D(n334), .Y(\mult_97/n2142 ) );
  OAI22X1 \mult_97/U1779  ( .A(\mult_97/n2663 ), .B(n321), .C(\mult_97/n2664 ), 
        .D(n334), .Y(\mult_97/n2141 ) );
  OAI22X1 \mult_97/U1778  ( .A(\mult_97/n2662 ), .B(n321), .C(\mult_97/n2663 ), 
        .D(n334), .Y(\mult_97/n2140 ) );
  OAI22X1 \mult_97/U1777  ( .A(\mult_97/n2661 ), .B(n321), .C(\mult_97/n2662 ), 
        .D(n334), .Y(\mult_97/n2139 ) );
  OAI22X1 \mult_97/U1776  ( .A(\mult_97/n2660 ), .B(n321), .C(\mult_97/n2661 ), 
        .D(n334), .Y(\mult_97/n2138 ) );
  OAI22X1 \mult_97/U1775  ( .A(\mult_97/n2659 ), .B(\mult_97/n368 ), .C(
        \mult_97/n2660 ), .D(n334), .Y(\mult_97/n2137 ) );
  OAI22X1 \mult_97/U1774  ( .A(\mult_97/n2658 ), .B(n321), .C(\mult_97/n2659 ), 
        .D(n334), .Y(\mult_97/n2136 ) );
  OAI22X1 \mult_97/U1773  ( .A(\mult_97/n2657 ), .B(\mult_97/n368 ), .C(
        \mult_97/n2658 ), .D(n334), .Y(\mult_97/n2135 ) );
  OAI22X1 \mult_97/U1772  ( .A(\mult_97/n2656 ), .B(\mult_97/n368 ), .C(
        \mult_97/n2657 ), .D(n334), .Y(\mult_97/n2134 ) );
  OAI22X1 \mult_97/U1771  ( .A(\mult_97/n2655 ), .B(\mult_97/n368 ), .C(
        \mult_97/n2656 ), .D(n334), .Y(\mult_97/n2133 ) );
  OAI22X1 \mult_97/U1770  ( .A(\mult_97/n2654 ), .B(\mult_97/n368 ), .C(
        \mult_97/n2655 ), .D(n334), .Y(\mult_97/n2132 ) );
  OAI22X1 \mult_97/U1769  ( .A(\mult_97/n2653 ), .B(\mult_97/n368 ), .C(
        \mult_97/n2654 ), .D(n334), .Y(\mult_97/n2131 ) );
  OAI22X1 \mult_97/U1768  ( .A(\mult_97/n2652 ), .B(n321), .C(\mult_97/n2653 ), 
        .D(n334), .Y(\mult_97/n2130 ) );
  OAI22X1 \mult_97/U1767  ( .A(\mult_97/n2651 ), .B(n321), .C(\mult_97/n2652 ), 
        .D(n334), .Y(\mult_97/n2129 ) );
  OAI22X1 \mult_97/U1766  ( .A(\mult_97/n2650 ), .B(n321), .C(\mult_97/n2651 ), 
        .D(n334), .Y(\mult_97/n2128 ) );
  OAI22X1 \mult_97/U1765  ( .A(\mult_97/n2649 ), .B(n321), .C(\mult_97/n2650 ), 
        .D(n334), .Y(\mult_97/n2127 ) );
  OAI22X1 \mult_97/U1764  ( .A(\mult_97/n2648 ), .B(n321), .C(\mult_97/n2649 ), 
        .D(n334), .Y(\mult_97/n2126 ) );
  OAI22X1 \mult_97/U1763  ( .A(\mult_97/n2647 ), .B(n321), .C(\mult_97/n2648 ), 
        .D(n334), .Y(\mult_97/n2125 ) );
  OAI22X1 \mult_97/U1762  ( .A(\mult_97/n2646 ), .B(n321), .C(\mult_97/n2647 ), 
        .D(n334), .Y(\mult_97/n2124 ) );
  OAI22X1 \mult_97/U1761  ( .A(\mult_97/n2645 ), .B(n321), .C(\mult_97/n2646 ), 
        .D(n334), .Y(\mult_97/n2123 ) );
  OAI22X1 \mult_97/U1760  ( .A(\mult_97/n2644 ), .B(n321), .C(\mult_97/n2645 ), 
        .D(n334), .Y(\mult_97/n2122 ) );
  OAI22X1 \mult_97/U1759  ( .A(\mult_97/n2643 ), .B(n321), .C(\mult_97/n2644 ), 
        .D(n334), .Y(\mult_97/n2121 ) );
  OAI22X1 \mult_97/U1758  ( .A(\mult_97/n368 ), .B(\mult_97/n2675 ), .C(n288), 
        .D(n334), .Y(\mult_97/n1859 ) );
  XNOR2X1 \mult_97/U1757  ( .A(n287), .B(n251), .Y(\mult_97/n2641 ) );
  XNOR2X1 \mult_97/U1756  ( .A(n287), .B(n400), .Y(\mult_97/n2640 ) );
  XNOR2X1 \mult_97/U1755  ( .A(n287), .B(n398), .Y(\mult_97/n2639 ) );
  XNOR2X1 \mult_97/U1754  ( .A(n287), .B(n396), .Y(\mult_97/n2638 ) );
  XNOR2X1 \mult_97/U1753  ( .A(n287), .B(n394), .Y(\mult_97/n2637 ) );
  XNOR2X1 \mult_97/U1752  ( .A(n287), .B(n392), .Y(\mult_97/n2636 ) );
  XNOR2X1 \mult_97/U1751  ( .A(n287), .B(n390), .Y(\mult_97/n2635 ) );
  XNOR2X1 \mult_97/U1750  ( .A(n287), .B(n388), .Y(\mult_97/n2634 ) );
  XNOR2X1 \mult_97/U1749  ( .A(n286), .B(n386), .Y(\mult_97/n2633 ) );
  XNOR2X1 \mult_97/U1748  ( .A(n287), .B(n384), .Y(\mult_97/n2632 ) );
  XNOR2X1 \mult_97/U1747  ( .A(n287), .B(n382), .Y(\mult_97/n2631 ) );
  XNOR2X1 \mult_97/U1746  ( .A(n286), .B(n380), .Y(\mult_97/n2630 ) );
  XNOR2X1 \mult_97/U1745  ( .A(n286), .B(n378), .Y(\mult_97/n2629 ) );
  XNOR2X1 \mult_97/U1744  ( .A(n286), .B(n376), .Y(\mult_97/n2628 ) );
  XNOR2X1 \mult_97/U1743  ( .A(n286), .B(n374), .Y(\mult_97/n2627 ) );
  XNOR2X1 \mult_97/U1742  ( .A(n286), .B(n372), .Y(\mult_97/n2626 ) );
  XNOR2X1 \mult_97/U1741  ( .A(n286), .B(n370), .Y(\mult_97/n2625 ) );
  XNOR2X1 \mult_97/U1740  ( .A(n286), .B(n368), .Y(\mult_97/n2624 ) );
  XNOR2X1 \mult_97/U1739  ( .A(n286), .B(n366), .Y(\mult_97/n2623 ) );
  XNOR2X1 \mult_97/U1738  ( .A(n286), .B(n364), .Y(\mult_97/n2622 ) );
  XNOR2X1 \mult_97/U1737  ( .A(n286), .B(n362), .Y(\mult_97/n2621 ) );
  XNOR2X1 \mult_97/U1736  ( .A(n286), .B(n360), .Y(\mult_97/n2620 ) );
  XNOR2X1 \mult_97/U1735  ( .A(n286), .B(n358), .Y(\mult_97/n2619 ) );
  XNOR2X1 \mult_97/U1734  ( .A(n286), .B(n356), .Y(\mult_97/n2618 ) );
  XNOR2X1 \mult_97/U1733  ( .A(n286), .B(n354), .Y(\mult_97/n2617 ) );
  XNOR2X1 \mult_97/U1732  ( .A(n286), .B(n352), .Y(\mult_97/n2616 ) );
  XNOR2X1 \mult_97/U1731  ( .A(n286), .B(n350), .Y(\mult_97/n2615 ) );
  XNOR2X1 \mult_97/U1730  ( .A(n286), .B(n348), .Y(\mult_97/n2614 ) );
  XNOR2X1 \mult_97/U1729  ( .A(n286), .B(n346), .Y(\mult_97/n2613 ) );
  XNOR2X1 \mult_97/U1728  ( .A(n286), .B(n344), .Y(\mult_97/n2612 ) );
  XNOR2X1 \mult_97/U1727  ( .A(n286), .B(n342), .Y(\mult_97/n2611 ) );
  XNOR2X1 \mult_97/U1726  ( .A(n287), .B(n340), .Y(\mult_97/n2610 ) );
  OAI22X1 \mult_97/U1725  ( .A(n323), .B(\mult_97/n2640 ), .C(\mult_97/n2641 ), 
        .D(n335), .Y(\mult_97/n2118 ) );
  OAI22X1 \mult_97/U1724  ( .A(n323), .B(\mult_97/n2639 ), .C(\mult_97/n2640 ), 
        .D(n335), .Y(\mult_97/n2117 ) );
  OAI22X1 \mult_97/U1723  ( .A(n323), .B(\mult_97/n2638 ), .C(\mult_97/n2639 ), 
        .D(n335), .Y(\mult_97/n2116 ) );
  OAI22X1 \mult_97/U1722  ( .A(n323), .B(\mult_97/n2637 ), .C(\mult_97/n2638 ), 
        .D(n335), .Y(\mult_97/n2115 ) );
  OAI22X1 \mult_97/U1721  ( .A(n323), .B(\mult_97/n2636 ), .C(\mult_97/n2637 ), 
        .D(n335), .Y(\mult_97/n2114 ) );
  OAI22X1 \mult_97/U1720  ( .A(n323), .B(\mult_97/n2635 ), .C(\mult_97/n2636 ), 
        .D(n335), .Y(\mult_97/n2113 ) );
  OAI22X1 \mult_97/U1719  ( .A(n323), .B(\mult_97/n2634 ), .C(\mult_97/n2635 ), 
        .D(n335), .Y(\mult_97/n2112 ) );
  OAI22X1 \mult_97/U1718  ( .A(n323), .B(\mult_97/n2633 ), .C(\mult_97/n2634 ), 
        .D(n335), .Y(\mult_97/n2111 ) );
  OAI22X1 \mult_97/U1717  ( .A(n323), .B(\mult_97/n2632 ), .C(\mult_97/n2633 ), 
        .D(n335), .Y(\mult_97/n2110 ) );
  OAI22X1 \mult_97/U1716  ( .A(n323), .B(\mult_97/n2631 ), .C(\mult_97/n2632 ), 
        .D(n335), .Y(\mult_97/n2109 ) );
  OAI22X1 \mult_97/U1715  ( .A(n323), .B(\mult_97/n2630 ), .C(\mult_97/n2631 ), 
        .D(n335), .Y(\mult_97/n2108 ) );
  OAI22X1 \mult_97/U1714  ( .A(n323), .B(\mult_97/n2629 ), .C(\mult_97/n2630 ), 
        .D(n335), .Y(\mult_97/n2107 ) );
  OAI22X1 \mult_97/U1713  ( .A(n323), .B(\mult_97/n2628 ), .C(\mult_97/n2629 ), 
        .D(n335), .Y(\mult_97/n2106 ) );
  OAI22X1 \mult_97/U1712  ( .A(\mult_97/n371 ), .B(\mult_97/n2627 ), .C(
        \mult_97/n2628 ), .D(n335), .Y(\mult_97/n2105 ) );
  OAI22X1 \mult_97/U1711  ( .A(n323), .B(\mult_97/n2626 ), .C(\mult_97/n2627 ), 
        .D(n335), .Y(\mult_97/n2104 ) );
  OAI22X1 \mult_97/U1710  ( .A(\mult_97/n371 ), .B(\mult_97/n2625 ), .C(
        \mult_97/n2626 ), .D(n335), .Y(\mult_97/n2103 ) );
  OAI22X1 \mult_97/U1709  ( .A(\mult_97/n371 ), .B(\mult_97/n2624 ), .C(
        \mult_97/n2625 ), .D(n335), .Y(\mult_97/n2102 ) );
  OAI22X1 \mult_97/U1708  ( .A(\mult_97/n371 ), .B(\mult_97/n2623 ), .C(
        \mult_97/n2624 ), .D(n335), .Y(\mult_97/n2101 ) );
  OAI22X1 \mult_97/U1707  ( .A(\mult_97/n371 ), .B(\mult_97/n2622 ), .C(
        \mult_97/n2623 ), .D(n335), .Y(\mult_97/n2100 ) );
  OAI22X1 \mult_97/U1706  ( .A(\mult_97/n371 ), .B(\mult_97/n2621 ), .C(
        \mult_97/n2622 ), .D(n335), .Y(\mult_97/n2099 ) );
  OAI22X1 \mult_97/U1705  ( .A(\mult_97/n371 ), .B(\mult_97/n2620 ), .C(
        \mult_97/n2621 ), .D(n335), .Y(\mult_97/n2098 ) );
  OAI22X1 \mult_97/U1704  ( .A(n323), .B(\mult_97/n2619 ), .C(\mult_97/n2620 ), 
        .D(n335), .Y(\mult_97/n2097 ) );
  OAI22X1 \mult_97/U1703  ( .A(n323), .B(\mult_97/n2618 ), .C(\mult_97/n2619 ), 
        .D(n335), .Y(\mult_97/n2096 ) );
  OAI22X1 \mult_97/U1702  ( .A(n323), .B(\mult_97/n2617 ), .C(\mult_97/n2618 ), 
        .D(n335), .Y(\mult_97/n2095 ) );
  OAI22X1 \mult_97/U1701  ( .A(n323), .B(\mult_97/n2616 ), .C(\mult_97/n2617 ), 
        .D(n335), .Y(\mult_97/n2094 ) );
  OAI22X1 \mult_97/U1700  ( .A(n323), .B(\mult_97/n2615 ), .C(\mult_97/n2616 ), 
        .D(n335), .Y(\mult_97/n2093 ) );
  OAI22X1 \mult_97/U1699  ( .A(n323), .B(\mult_97/n2614 ), .C(\mult_97/n2615 ), 
        .D(n335), .Y(\mult_97/n2092 ) );
  OAI22X1 \mult_97/U1698  ( .A(n323), .B(\mult_97/n2613 ), .C(\mult_97/n2614 ), 
        .D(n335), .Y(\mult_97/n2091 ) );
  OAI22X1 \mult_97/U1697  ( .A(n323), .B(\mult_97/n2612 ), .C(\mult_97/n2613 ), 
        .D(n335), .Y(\mult_97/n2090 ) );
  OAI22X1 \mult_97/U1696  ( .A(n323), .B(\mult_97/n2611 ), .C(\mult_97/n2612 ), 
        .D(n335), .Y(\mult_97/n2089 ) );
  OAI22X1 \mult_97/U1695  ( .A(n323), .B(\mult_97/n2610 ), .C(\mult_97/n2611 ), 
        .D(n335), .Y(\mult_97/n2088 ) );
  OAI22X1 \mult_97/U1694  ( .A(n323), .B(\mult_97/n2642 ), .C(n285), .D(n335), 
        .Y(\mult_97/n1858 ) );
  XNOR2X1 \mult_97/U1693  ( .A(n251), .B(n284), .Y(\mult_97/n2608 ) );
  XNOR2X1 \mult_97/U1692  ( .A(n400), .B(n284), .Y(\mult_97/n2607 ) );
  XNOR2X1 \mult_97/U1691  ( .A(n398), .B(n284), .Y(\mult_97/n2606 ) );
  XNOR2X1 \mult_97/U1690  ( .A(n396), .B(n284), .Y(\mult_97/n2605 ) );
  XNOR2X1 \mult_97/U1689  ( .A(B[4]), .B(n284), .Y(\mult_97/n2604 ) );
  XNOR2X1 \mult_97/U1688  ( .A(n392), .B(n284), .Y(\mult_97/n2603 ) );
  XNOR2X1 \mult_97/U1687  ( .A(n390), .B(n284), .Y(\mult_97/n2602 ) );
  XNOR2X1 \mult_97/U1686  ( .A(n388), .B(n284), .Y(\mult_97/n2601 ) );
  XNOR2X1 \mult_97/U1685  ( .A(n386), .B(n283), .Y(\mult_97/n2600 ) );
  XNOR2X1 \mult_97/U1684  ( .A(n384), .B(n284), .Y(\mult_97/n2599 ) );
  XNOR2X1 \mult_97/U1683  ( .A(n382), .B(n284), .Y(\mult_97/n2598 ) );
  XNOR2X1 \mult_97/U1682  ( .A(n380), .B(n283), .Y(\mult_97/n2597 ) );
  XNOR2X1 \mult_97/U1681  ( .A(n378), .B(n283), .Y(\mult_97/n2596 ) );
  XNOR2X1 \mult_97/U1680  ( .A(n376), .B(n283), .Y(\mult_97/n2595 ) );
  XNOR2X1 \mult_97/U1679  ( .A(n374), .B(n283), .Y(\mult_97/n2594 ) );
  XNOR2X1 \mult_97/U1678  ( .A(n372), .B(n283), .Y(\mult_97/n2593 ) );
  XNOR2X1 \mult_97/U1677  ( .A(n370), .B(n283), .Y(\mult_97/n2592 ) );
  XNOR2X1 \mult_97/U1676  ( .A(n368), .B(n283), .Y(\mult_97/n2591 ) );
  XNOR2X1 \mult_97/U1675  ( .A(n366), .B(n283), .Y(\mult_97/n2590 ) );
  XNOR2X1 \mult_97/U1674  ( .A(n364), .B(n283), .Y(\mult_97/n2589 ) );
  XNOR2X1 \mult_97/U1673  ( .A(n362), .B(n283), .Y(\mult_97/n2588 ) );
  XNOR2X1 \mult_97/U1672  ( .A(n360), .B(n283), .Y(\mult_97/n2587 ) );
  XNOR2X1 \mult_97/U1671  ( .A(n358), .B(n283), .Y(\mult_97/n2586 ) );
  XNOR2X1 \mult_97/U1670  ( .A(n356), .B(n283), .Y(\mult_97/n2585 ) );
  XNOR2X1 \mult_97/U1669  ( .A(n354), .B(n283), .Y(\mult_97/n2584 ) );
  XNOR2X1 \mult_97/U1668  ( .A(n352), .B(n283), .Y(\mult_97/n2583 ) );
  XNOR2X1 \mult_97/U1667  ( .A(B[26]), .B(n283), .Y(\mult_97/n2582 ) );
  XNOR2X1 \mult_97/U1666  ( .A(n348), .B(n283), .Y(\mult_97/n2581 ) );
  XNOR2X1 \mult_97/U1665  ( .A(n346), .B(n283), .Y(\mult_97/n2580 ) );
  XNOR2X1 \mult_97/U1664  ( .A(n344), .B(n283), .Y(\mult_97/n2579 ) );
  XNOR2X1 \mult_97/U1663  ( .A(n342), .B(n283), .Y(\mult_97/n2578 ) );
  XNOR2X1 \mult_97/U1662  ( .A(n340), .B(n284), .Y(\mult_97/n2577 ) );
  OAI22X1 \mult_97/U1661  ( .A(\mult_97/n2607 ), .B(n325), .C(\mult_97/n2608 ), 
        .D(n336), .Y(\mult_97/n2085 ) );
  OAI22X1 \mult_97/U1660  ( .A(\mult_97/n2606 ), .B(n325), .C(\mult_97/n2607 ), 
        .D(n336), .Y(\mult_97/n2084 ) );
  OAI22X1 \mult_97/U1659  ( .A(\mult_97/n2605 ), .B(n325), .C(\mult_97/n2606 ), 
        .D(n336), .Y(\mult_97/n2083 ) );
  OAI22X1 \mult_97/U1658  ( .A(\mult_97/n2604 ), .B(n325), .C(\mult_97/n2605 ), 
        .D(n336), .Y(\mult_97/n2082 ) );
  OAI22X1 \mult_97/U1657  ( .A(\mult_97/n2603 ), .B(n325), .C(\mult_97/n2604 ), 
        .D(n336), .Y(\mult_97/n2081 ) );
  OAI22X1 \mult_97/U1656  ( .A(\mult_97/n2602 ), .B(n325), .C(\mult_97/n2603 ), 
        .D(n336), .Y(\mult_97/n2080 ) );
  OAI22X1 \mult_97/U1655  ( .A(\mult_97/n2601 ), .B(n325), .C(\mult_97/n2602 ), 
        .D(n336), .Y(\mult_97/n2079 ) );
  OAI22X1 \mult_97/U1654  ( .A(\mult_97/n2600 ), .B(n325), .C(\mult_97/n2601 ), 
        .D(n336), .Y(\mult_97/n2078 ) );
  OAI22X1 \mult_97/U1653  ( .A(\mult_97/n2599 ), .B(n325), .C(\mult_97/n2600 ), 
        .D(n336), .Y(\mult_97/n2077 ) );
  OAI22X1 \mult_97/U1652  ( .A(\mult_97/n2598 ), .B(n325), .C(\mult_97/n2599 ), 
        .D(n336), .Y(\mult_97/n2076 ) );
  OAI22X1 \mult_97/U1651  ( .A(\mult_97/n2597 ), .B(n325), .C(\mult_97/n2598 ), 
        .D(n336), .Y(\mult_97/n2075 ) );
  OAI22X1 \mult_97/U1650  ( .A(\mult_97/n2596 ), .B(n325), .C(\mult_97/n2597 ), 
        .D(n336), .Y(\mult_97/n2074 ) );
  OAI22X1 \mult_97/U1649  ( .A(\mult_97/n2595 ), .B(n325), .C(\mult_97/n2596 ), 
        .D(n336), .Y(\mult_97/n2073 ) );
  OAI22X1 \mult_97/U1648  ( .A(\mult_97/n2594 ), .B(n325), .C(\mult_97/n2595 ), 
        .D(n336), .Y(\mult_97/n2072 ) );
  OAI22X1 \mult_97/U1647  ( .A(\mult_97/n2593 ), .B(\mult_97/n374 ), .C(
        \mult_97/n2594 ), .D(n336), .Y(\mult_97/n2071 ) );
  OAI22X1 \mult_97/U1646  ( .A(\mult_97/n2592 ), .B(\mult_97/n374 ), .C(
        \mult_97/n2593 ), .D(n336), .Y(\mult_97/n2070 ) );
  OAI22X1 \mult_97/U1645  ( .A(\mult_97/n2591 ), .B(\mult_97/n374 ), .C(
        \mult_97/n2592 ), .D(n336), .Y(\mult_97/n2069 ) );
  OAI22X1 \mult_97/U1644  ( .A(\mult_97/n2590 ), .B(\mult_97/n374 ), .C(
        \mult_97/n2591 ), .D(n336), .Y(\mult_97/n2068 ) );
  OAI22X1 \mult_97/U1643  ( .A(\mult_97/n2589 ), .B(\mult_97/n374 ), .C(
        \mult_97/n2590 ), .D(n336), .Y(\mult_97/n2067 ) );
  OAI22X1 \mult_97/U1642  ( .A(\mult_97/n2588 ), .B(\mult_97/n374 ), .C(
        \mult_97/n2589 ), .D(n336), .Y(\mult_97/n2066 ) );
  OAI22X1 \mult_97/U1641  ( .A(\mult_97/n2587 ), .B(n325), .C(\mult_97/n2588 ), 
        .D(n336), .Y(\mult_97/n1207 ) );
  OAI22X1 \mult_97/U1640  ( .A(\mult_97/n2586 ), .B(n325), .C(\mult_97/n2587 ), 
        .D(n336), .Y(\mult_97/n2065 ) );
  OAI22X1 \mult_97/U1639  ( .A(\mult_97/n2585 ), .B(n325), .C(\mult_97/n2586 ), 
        .D(n336), .Y(\mult_97/n2064 ) );
  OAI22X1 \mult_97/U1638  ( .A(\mult_97/n2584 ), .B(n325), .C(\mult_97/n2585 ), 
        .D(n336), .Y(\mult_97/n2063 ) );
  OAI22X1 \mult_97/U1637  ( .A(\mult_97/n2583 ), .B(n325), .C(\mult_97/n2584 ), 
        .D(n336), .Y(\mult_97/n2062 ) );
  OAI22X1 \mult_97/U1636  ( .A(\mult_97/n2582 ), .B(n325), .C(\mult_97/n2583 ), 
        .D(n336), .Y(\mult_97/n2061 ) );
  OAI22X1 \mult_97/U1635  ( .A(\mult_97/n2581 ), .B(n325), .C(\mult_97/n2582 ), 
        .D(n336), .Y(\mult_97/n2060 ) );
  OAI22X1 \mult_97/U1634  ( .A(\mult_97/n2580 ), .B(n325), .C(\mult_97/n2581 ), 
        .D(n336), .Y(\mult_97/n2059 ) );
  OAI22X1 \mult_97/U1633  ( .A(\mult_97/n2579 ), .B(n325), .C(\mult_97/n2580 ), 
        .D(n336), .Y(\mult_97/n2058 ) );
  OAI22X1 \mult_97/U1632  ( .A(\mult_97/n2578 ), .B(n325), .C(\mult_97/n2579 ), 
        .D(n336), .Y(\mult_97/n2057 ) );
  OAI22X1 \mult_97/U1631  ( .A(\mult_97/n2577 ), .B(n325), .C(\mult_97/n2578 ), 
        .D(n336), .Y(\mult_97/n1017 ) );
  OAI22X1 \mult_97/U1630  ( .A(\mult_97/n374 ), .B(\mult_97/n2609 ), .C(n282), 
        .D(n336), .Y(\mult_97/n1857 ) );
  XNOR2X1 \mult_97/U1629  ( .A(n251), .B(A[21]), .Y(\mult_97/n2575 ) );
  XNOR2X1 \mult_97/U1628  ( .A(n400), .B(n281), .Y(\mult_97/n2574 ) );
  XNOR2X1 \mult_97/U1627  ( .A(n398), .B(n281), .Y(\mult_97/n2573 ) );
  XNOR2X1 \mult_97/U1626  ( .A(n396), .B(n281), .Y(\mult_97/n2572 ) );
  XNOR2X1 \mult_97/U1625  ( .A(n394), .B(n281), .Y(\mult_97/n2571 ) );
  XNOR2X1 \mult_97/U1624  ( .A(n392), .B(n281), .Y(\mult_97/n2570 ) );
  XNOR2X1 \mult_97/U1623  ( .A(n390), .B(n281), .Y(\mult_97/n2569 ) );
  XNOR2X1 \mult_97/U1622  ( .A(n388), .B(n281), .Y(\mult_97/n2568 ) );
  XNOR2X1 \mult_97/U1621  ( .A(n386), .B(n281), .Y(\mult_97/n2567 ) );
  XNOR2X1 \mult_97/U1620  ( .A(n384), .B(n281), .Y(\mult_97/n2566 ) );
  XNOR2X1 \mult_97/U1619  ( .A(n382), .B(A[21]), .Y(\mult_97/n2565 ) );
  XNOR2X1 \mult_97/U1618  ( .A(n380), .B(n281), .Y(\mult_97/n2564 ) );
  XNOR2X1 \mult_97/U1617  ( .A(n378), .B(n281), .Y(\mult_97/n2563 ) );
  XNOR2X1 \mult_97/U1616  ( .A(n376), .B(n281), .Y(\mult_97/n2562 ) );
  XNOR2X1 \mult_97/U1615  ( .A(n374), .B(n281), .Y(\mult_97/n2561 ) );
  XNOR2X1 \mult_97/U1614  ( .A(n372), .B(n281), .Y(\mult_97/n2560 ) );
  XNOR2X1 \mult_97/U1613  ( .A(n370), .B(n281), .Y(\mult_97/n2559 ) );
  XNOR2X1 \mult_97/U1612  ( .A(B[17]), .B(n281), .Y(\mult_97/n2558 ) );
  XNOR2X1 \mult_97/U1611  ( .A(n366), .B(n281), .Y(\mult_97/n2557 ) );
  XNOR2X1 \mult_97/U1610  ( .A(n364), .B(n281), .Y(\mult_97/n2556 ) );
  XNOR2X1 \mult_97/U1609  ( .A(n362), .B(n281), .Y(\mult_97/n2555 ) );
  XNOR2X1 \mult_97/U1608  ( .A(n360), .B(n281), .Y(\mult_97/n2554 ) );
  XNOR2X1 \mult_97/U1607  ( .A(n358), .B(n281), .Y(\mult_97/n2553 ) );
  XNOR2X1 \mult_97/U1606  ( .A(B[23]), .B(n281), .Y(\mult_97/n2552 ) );
  XNOR2X1 \mult_97/U1605  ( .A(B[24]), .B(n281), .Y(\mult_97/n2551 ) );
  XNOR2X1 \mult_97/U1604  ( .A(n352), .B(n281), .Y(\mult_97/n2550 ) );
  XNOR2X1 \mult_97/U1603  ( .A(n350), .B(n281), .Y(\mult_97/n2549 ) );
  XNOR2X1 \mult_97/U1602  ( .A(n348), .B(n281), .Y(\mult_97/n2548 ) );
  XNOR2X1 \mult_97/U1601  ( .A(n346), .B(n281), .Y(\mult_97/n2547 ) );
  XNOR2X1 \mult_97/U1600  ( .A(n344), .B(n281), .Y(\mult_97/n2546 ) );
  XNOR2X1 \mult_97/U1599  ( .A(n342), .B(n281), .Y(\mult_97/n2545 ) );
  XNOR2X1 \mult_97/U1598  ( .A(n340), .B(n281), .Y(\mult_97/n2544 ) );
  OAI22X1 \mult_97/U1597  ( .A(\mult_97/n2574 ), .B(n326), .C(\mult_97/n2575 ), 
        .D(n337), .Y(\mult_97/n2054 ) );
  OAI22X1 \mult_97/U1596  ( .A(\mult_97/n2573 ), .B(n326), .C(\mult_97/n2574 ), 
        .D(n337), .Y(\mult_97/n2053 ) );
  OAI22X1 \mult_97/U1595  ( .A(\mult_97/n2572 ), .B(n326), .C(\mult_97/n2573 ), 
        .D(n337), .Y(\mult_97/n2052 ) );
  OAI22X1 \mult_97/U1594  ( .A(\mult_97/n2571 ), .B(n326), .C(\mult_97/n2572 ), 
        .D(n337), .Y(\mult_97/n2051 ) );
  OAI22X1 \mult_97/U1593  ( .A(\mult_97/n2570 ), .B(n326), .C(\mult_97/n2571 ), 
        .D(n337), .Y(\mult_97/n2050 ) );
  OAI22X1 \mult_97/U1592  ( .A(\mult_97/n2569 ), .B(n326), .C(\mult_97/n2570 ), 
        .D(n337), .Y(\mult_97/n2049 ) );
  OAI22X1 \mult_97/U1591  ( .A(\mult_97/n2568 ), .B(n326), .C(\mult_97/n2569 ), 
        .D(n337), .Y(\mult_97/n2048 ) );
  OAI22X1 \mult_97/U1590  ( .A(\mult_97/n2567 ), .B(n326), .C(\mult_97/n2568 ), 
        .D(n337), .Y(\mult_97/n2047 ) );
  OAI22X1 \mult_97/U1589  ( .A(\mult_97/n2566 ), .B(n326), .C(\mult_97/n2567 ), 
        .D(n337), .Y(\mult_97/n2046 ) );
  OAI22X1 \mult_97/U1588  ( .A(\mult_97/n2565 ), .B(n326), .C(\mult_97/n2566 ), 
        .D(n337), .Y(\mult_97/n2045 ) );
  OAI22X1 \mult_97/U1587  ( .A(\mult_97/n2564 ), .B(n326), .C(\mult_97/n2565 ), 
        .D(n337), .Y(\mult_97/n2044 ) );
  OAI22X1 \mult_97/U1586  ( .A(\mult_97/n2563 ), .B(n326), .C(\mult_97/n2564 ), 
        .D(n337), .Y(\mult_97/n2043 ) );
  OAI22X1 \mult_97/U1585  ( .A(\mult_97/n2562 ), .B(n326), .C(\mult_97/n2563 ), 
        .D(n337), .Y(\mult_97/n2042 ) );
  OAI22X1 \mult_97/U1584  ( .A(\mult_97/n2561 ), .B(n326), .C(\mult_97/n2562 ), 
        .D(n337), .Y(\mult_97/n2041 ) );
  OAI22X1 \mult_97/U1583  ( .A(\mult_97/n2560 ), .B(n326), .C(\mult_97/n2561 ), 
        .D(n337), .Y(\mult_97/n2040 ) );
  OAI22X1 \mult_97/U1582  ( .A(\mult_97/n2559 ), .B(n326), .C(\mult_97/n2560 ), 
        .D(n337), .Y(\mult_97/n2039 ) );
  OAI22X1 \mult_97/U1581  ( .A(\mult_97/n2558 ), .B(n326), .C(\mult_97/n2559 ), 
        .D(n337), .Y(\mult_97/n2038 ) );
  OAI22X1 \mult_97/U1580  ( .A(\mult_97/n2557 ), .B(n326), .C(\mult_97/n2558 ), 
        .D(n337), .Y(\mult_97/n2037 ) );
  OAI22X1 \mult_97/U1579  ( .A(\mult_97/n2556 ), .B(n326), .C(\mult_97/n2557 ), 
        .D(n337), .Y(\mult_97/n2036 ) );
  OAI22X1 \mult_97/U1578  ( .A(\mult_97/n2555 ), .B(n326), .C(\mult_97/n2556 ), 
        .D(n337), .Y(\mult_97/n2035 ) );
  OAI22X1 \mult_97/U1577  ( .A(\mult_97/n2554 ), .B(n326), .C(\mult_97/n2555 ), 
        .D(n337), .Y(\mult_97/n2034 ) );
  OAI22X1 \mult_97/U1576  ( .A(\mult_97/n2553 ), .B(n326), .C(\mult_97/n2554 ), 
        .D(n337), .Y(\mult_97/n2033 ) );
  OAI22X1 \mult_97/U1575  ( .A(\mult_97/n2552 ), .B(n326), .C(\mult_97/n2553 ), 
        .D(n337), .Y(\mult_97/n2032 ) );
  OAI22X1 \mult_97/U1574  ( .A(\mult_97/n2551 ), .B(n326), .C(\mult_97/n2552 ), 
        .D(n337), .Y(\mult_97/n2031 ) );
  OAI22X1 \mult_97/U1573  ( .A(\mult_97/n2550 ), .B(n326), .C(\mult_97/n2551 ), 
        .D(n337), .Y(\mult_97/n2030 ) );
  OAI22X1 \mult_97/U1572  ( .A(\mult_97/n2549 ), .B(n326), .C(\mult_97/n2550 ), 
        .D(n337), .Y(\mult_97/n2029 ) );
  OAI22X1 \mult_97/U1571  ( .A(\mult_97/n2548 ), .B(n326), .C(\mult_97/n2549 ), 
        .D(n337), .Y(\mult_97/n2028 ) );
  OAI22X1 \mult_97/U1570  ( .A(\mult_97/n2547 ), .B(n326), .C(\mult_97/n2548 ), 
        .D(n337), .Y(\mult_97/n2027 ) );
  OAI22X1 \mult_97/U1569  ( .A(\mult_97/n2546 ), .B(n326), .C(\mult_97/n2547 ), 
        .D(n337), .Y(\mult_97/n2026 ) );
  OAI22X1 \mult_97/U1568  ( .A(\mult_97/n2545 ), .B(n326), .C(\mult_97/n2546 ), 
        .D(n337), .Y(\mult_97/n2025 ) );
  OAI22X1 \mult_97/U1567  ( .A(\mult_97/n2544 ), .B(n326), .C(\mult_97/n2545 ), 
        .D(n337), .Y(\mult_97/n2024 ) );
  OAI22X1 \mult_97/U1566  ( .A(n326), .B(\mult_97/n2576 ), .C(n280), .D(n337), 
        .Y(\mult_97/n1856 ) );
  XNOR2X1 \mult_97/U1565  ( .A(n279), .B(n251), .Y(\mult_97/n2542 ) );
  XNOR2X1 \mult_97/U1564  ( .A(n279), .B(n400), .Y(\mult_97/n2541 ) );
  XNOR2X1 \mult_97/U1563  ( .A(n279), .B(n398), .Y(\mult_97/n2540 ) );
  XNOR2X1 \mult_97/U1562  ( .A(n279), .B(n396), .Y(\mult_97/n2539 ) );
  XNOR2X1 \mult_97/U1561  ( .A(n279), .B(n394), .Y(\mult_97/n2538 ) );
  XNOR2X1 \mult_97/U1560  ( .A(n279), .B(n392), .Y(\mult_97/n2537 ) );
  XNOR2X1 \mult_97/U1559  ( .A(n279), .B(n390), .Y(\mult_97/n2536 ) );
  XNOR2X1 \mult_97/U1558  ( .A(n279), .B(n388), .Y(\mult_97/n2535 ) );
  XNOR2X1 \mult_97/U1557  ( .A(n279), .B(n386), .Y(\mult_97/n2534 ) );
  XNOR2X1 \mult_97/U1556  ( .A(n279), .B(n384), .Y(\mult_97/n2533 ) );
  XNOR2X1 \mult_97/U1555  ( .A(n279), .B(n382), .Y(\mult_97/n2532 ) );
  XNOR2X1 \mult_97/U1554  ( .A(n279), .B(n380), .Y(\mult_97/n2531 ) );
  XNOR2X1 \mult_97/U1553  ( .A(n279), .B(n378), .Y(\mult_97/n2530 ) );
  XNOR2X1 \mult_97/U1552  ( .A(n279), .B(n376), .Y(\mult_97/n2529 ) );
  XNOR2X1 \mult_97/U1551  ( .A(n279), .B(n374), .Y(\mult_97/n2528 ) );
  XNOR2X1 \mult_97/U1550  ( .A(n279), .B(n372), .Y(\mult_97/n2527 ) );
  XNOR2X1 \mult_97/U1549  ( .A(n279), .B(n370), .Y(\mult_97/n2526 ) );
  XNOR2X1 \mult_97/U1548  ( .A(n279), .B(n368), .Y(\mult_97/n2525 ) );
  XNOR2X1 \mult_97/U1547  ( .A(n279), .B(n366), .Y(\mult_97/n2524 ) );
  XNOR2X1 \mult_97/U1546  ( .A(n279), .B(n364), .Y(\mult_97/n2523 ) );
  XNOR2X1 \mult_97/U1545  ( .A(n279), .B(n362), .Y(\mult_97/n2522 ) );
  XNOR2X1 \mult_97/U1544  ( .A(n279), .B(n360), .Y(\mult_97/n2521 ) );
  XNOR2X1 \mult_97/U1543  ( .A(n279), .B(n358), .Y(\mult_97/n2520 ) );
  XNOR2X1 \mult_97/U1542  ( .A(n279), .B(n356), .Y(\mult_97/n2519 ) );
  XNOR2X1 \mult_97/U1541  ( .A(n279), .B(n354), .Y(\mult_97/n2518 ) );
  XNOR2X1 \mult_97/U1540  ( .A(n279), .B(n352), .Y(\mult_97/n2517 ) );
  XNOR2X1 \mult_97/U1539  ( .A(n279), .B(n350), .Y(\mult_97/n2516 ) );
  XNOR2X1 \mult_97/U1538  ( .A(n279), .B(n348), .Y(\mult_97/n2515 ) );
  XNOR2X1 \mult_97/U1537  ( .A(n279), .B(n346), .Y(\mult_97/n2514 ) );
  XNOR2X1 \mult_97/U1536  ( .A(n279), .B(n344), .Y(\mult_97/n2513 ) );
  XNOR2X1 \mult_97/U1535  ( .A(n279), .B(n342), .Y(\mult_97/n2512 ) );
  XNOR2X1 \mult_97/U1534  ( .A(n279), .B(n340), .Y(\mult_97/n2511 ) );
  OAI22X1 \mult_97/U1533  ( .A(n327), .B(\mult_97/n2541 ), .C(\mult_97/n2542 ), 
        .D(n247), .Y(\mult_97/n2021 ) );
  OAI22X1 \mult_97/U1532  ( .A(n327), .B(\mult_97/n2540 ), .C(\mult_97/n2541 ), 
        .D(n247), .Y(\mult_97/n2020 ) );
  OAI22X1 \mult_97/U1531  ( .A(n327), .B(\mult_97/n2539 ), .C(\mult_97/n2540 ), 
        .D(n247), .Y(\mult_97/n2019 ) );
  OAI22X1 \mult_97/U1530  ( .A(n327), .B(\mult_97/n2538 ), .C(\mult_97/n2539 ), 
        .D(n247), .Y(\mult_97/n2018 ) );
  OAI22X1 \mult_97/U1529  ( .A(n327), .B(\mult_97/n2537 ), .C(\mult_97/n2538 ), 
        .D(n247), .Y(\mult_97/n2017 ) );
  OAI22X1 \mult_97/U1528  ( .A(n327), .B(\mult_97/n2536 ), .C(\mult_97/n2537 ), 
        .D(n247), .Y(\mult_97/n2016 ) );
  OAI22X1 \mult_97/U1527  ( .A(n327), .B(\mult_97/n2535 ), .C(\mult_97/n2536 ), 
        .D(n247), .Y(\mult_97/n2015 ) );
  OAI22X1 \mult_97/U1526  ( .A(n327), .B(\mult_97/n2534 ), .C(\mult_97/n2535 ), 
        .D(n247), .Y(\mult_97/n2014 ) );
  OAI22X1 \mult_97/U1525  ( .A(n327), .B(\mult_97/n2533 ), .C(\mult_97/n2534 ), 
        .D(n247), .Y(\mult_97/n2013 ) );
  OAI22X1 \mult_97/U1524  ( .A(n327), .B(\mult_97/n2532 ), .C(\mult_97/n2533 ), 
        .D(n247), .Y(\mult_97/n2012 ) );
  OAI22X1 \mult_97/U1523  ( .A(n327), .B(\mult_97/n2531 ), .C(\mult_97/n2532 ), 
        .D(n247), .Y(\mult_97/n2011 ) );
  OAI22X1 \mult_97/U1522  ( .A(n327), .B(\mult_97/n2530 ), .C(\mult_97/n2531 ), 
        .D(n247), .Y(\mult_97/n2010 ) );
  OAI22X1 \mult_97/U1521  ( .A(n327), .B(\mult_97/n2529 ), .C(\mult_97/n2530 ), 
        .D(n247), .Y(\mult_97/n2009 ) );
  OAI22X1 \mult_97/U1520  ( .A(n327), .B(\mult_97/n2528 ), .C(\mult_97/n2529 ), 
        .D(n247), .Y(\mult_97/n2008 ) );
  OAI22X1 \mult_97/U1519  ( .A(n327), .B(\mult_97/n2527 ), .C(\mult_97/n2528 ), 
        .D(n247), .Y(\mult_97/n2007 ) );
  OAI22X1 \mult_97/U1518  ( .A(n327), .B(\mult_97/n2526 ), .C(\mult_97/n2527 ), 
        .D(n247), .Y(\mult_97/n2006 ) );
  OAI22X1 \mult_97/U1517  ( .A(n327), .B(\mult_97/n2525 ), .C(\mult_97/n2526 ), 
        .D(n247), .Y(\mult_97/n2005 ) );
  OAI22X1 \mult_97/U1516  ( .A(n327), .B(\mult_97/n2524 ), .C(\mult_97/n2525 ), 
        .D(n247), .Y(\mult_97/n2004 ) );
  OAI22X1 \mult_97/U1515  ( .A(n327), .B(\mult_97/n2523 ), .C(\mult_97/n2524 ), 
        .D(n247), .Y(\mult_97/n2003 ) );
  OAI22X1 \mult_97/U1514  ( .A(n327), .B(\mult_97/n2522 ), .C(\mult_97/n2523 ), 
        .D(n247), .Y(\mult_97/n2002 ) );
  OAI22X1 \mult_97/U1513  ( .A(n327), .B(\mult_97/n2521 ), .C(\mult_97/n2522 ), 
        .D(n247), .Y(\mult_97/n2001 ) );
  OAI22X1 \mult_97/U1512  ( .A(n327), .B(\mult_97/n2520 ), .C(\mult_97/n2521 ), 
        .D(n247), .Y(\mult_97/n2000 ) );
  OAI22X1 \mult_97/U1511  ( .A(n327), .B(\mult_97/n2519 ), .C(\mult_97/n2520 ), 
        .D(n247), .Y(\mult_97/n1999 ) );
  OAI22X1 \mult_97/U1510  ( .A(n327), .B(\mult_97/n2518 ), .C(\mult_97/n2519 ), 
        .D(n247), .Y(\mult_97/n1998 ) );
  OAI22X1 \mult_97/U1509  ( .A(n327), .B(\mult_97/n2517 ), .C(\mult_97/n2518 ), 
        .D(n247), .Y(\mult_97/n1997 ) );
  OAI22X1 \mult_97/U1508  ( .A(n327), .B(\mult_97/n2516 ), .C(\mult_97/n2517 ), 
        .D(n247), .Y(\mult_97/n1996 ) );
  OAI22X1 \mult_97/U1507  ( .A(n327), .B(\mult_97/n2515 ), .C(\mult_97/n2516 ), 
        .D(n247), .Y(\mult_97/n1995 ) );
  OAI22X1 \mult_97/U1506  ( .A(n327), .B(\mult_97/n2514 ), .C(\mult_97/n2515 ), 
        .D(n247), .Y(\mult_97/n1994 ) );
  OAI22X1 \mult_97/U1505  ( .A(n327), .B(\mult_97/n2513 ), .C(\mult_97/n2514 ), 
        .D(n247), .Y(\mult_97/n1993 ) );
  OAI22X1 \mult_97/U1504  ( .A(n327), .B(\mult_97/n2512 ), .C(\mult_97/n2513 ), 
        .D(n247), .Y(\mult_97/n1992 ) );
  OAI22X1 \mult_97/U1503  ( .A(n327), .B(\mult_97/n2511 ), .C(\mult_97/n2512 ), 
        .D(n247), .Y(\mult_97/n1991 ) );
  OAI22X1 \mult_97/U1502  ( .A(n327), .B(\mult_97/n2543 ), .C(n278), .D(n247), 
        .Y(\mult_97/n1855 ) );
  XNOR2X1 \mult_97/U1501  ( .A(n251), .B(n277), .Y(\mult_97/n2509 ) );
  XNOR2X1 \mult_97/U1500  ( .A(n400), .B(n277), .Y(\mult_97/n2508 ) );
  XNOR2X1 \mult_97/U1499  ( .A(n398), .B(n277), .Y(\mult_97/n2507 ) );
  XNOR2X1 \mult_97/U1498  ( .A(n396), .B(n277), .Y(\mult_97/n2506 ) );
  XNOR2X1 \mult_97/U1497  ( .A(n394), .B(n277), .Y(\mult_97/n2505 ) );
  XNOR2X1 \mult_97/U1496  ( .A(n392), .B(n277), .Y(\mult_97/n2504 ) );
  XNOR2X1 \mult_97/U1495  ( .A(n390), .B(n277), .Y(\mult_97/n2503 ) );
  XNOR2X1 \mult_97/U1494  ( .A(B[7]), .B(n277), .Y(\mult_97/n2502 ) );
  XNOR2X1 \mult_97/U1493  ( .A(n386), .B(n276), .Y(\mult_97/n2501 ) );
  XNOR2X1 \mult_97/U1492  ( .A(n384), .B(n277), .Y(\mult_97/n2500 ) );
  XNOR2X1 \mult_97/U1491  ( .A(n382), .B(n277), .Y(\mult_97/n2499 ) );
  XNOR2X1 \mult_97/U1490  ( .A(n380), .B(n276), .Y(\mult_97/n2498 ) );
  XNOR2X1 \mult_97/U1489  ( .A(n378), .B(n276), .Y(\mult_97/n2497 ) );
  XNOR2X1 \mult_97/U1488  ( .A(n376), .B(n276), .Y(\mult_97/n2496 ) );
  XNOR2X1 \mult_97/U1487  ( .A(n374), .B(n276), .Y(\mult_97/n2495 ) );
  XNOR2X1 \mult_97/U1486  ( .A(n372), .B(n276), .Y(\mult_97/n2494 ) );
  XNOR2X1 \mult_97/U1485  ( .A(n370), .B(n276), .Y(\mult_97/n2493 ) );
  XNOR2X1 \mult_97/U1484  ( .A(n368), .B(n276), .Y(\mult_97/n2492 ) );
  XNOR2X1 \mult_97/U1483  ( .A(n366), .B(n276), .Y(\mult_97/n2491 ) );
  XNOR2X1 \mult_97/U1482  ( .A(n364), .B(n276), .Y(\mult_97/n2490 ) );
  XNOR2X1 \mult_97/U1481  ( .A(n362), .B(n276), .Y(\mult_97/n2489 ) );
  XNOR2X1 \mult_97/U1480  ( .A(n360), .B(n276), .Y(\mult_97/n2488 ) );
  XNOR2X1 \mult_97/U1479  ( .A(n358), .B(n276), .Y(\mult_97/n2487 ) );
  XNOR2X1 \mult_97/U1478  ( .A(n356), .B(n276), .Y(\mult_97/n2486 ) );
  XNOR2X1 \mult_97/U1477  ( .A(n354), .B(n276), .Y(\mult_97/n2485 ) );
  XNOR2X1 \mult_97/U1476  ( .A(n352), .B(n276), .Y(\mult_97/n2484 ) );
  XNOR2X1 \mult_97/U1475  ( .A(n350), .B(n276), .Y(\mult_97/n2483 ) );
  XNOR2X1 \mult_97/U1474  ( .A(n348), .B(n276), .Y(\mult_97/n2482 ) );
  XNOR2X1 \mult_97/U1473  ( .A(n346), .B(n276), .Y(\mult_97/n2481 ) );
  XNOR2X1 \mult_97/U1472  ( .A(n344), .B(n276), .Y(\mult_97/n2480 ) );
  XNOR2X1 \mult_97/U1471  ( .A(n342), .B(n276), .Y(\mult_97/n2479 ) );
  XNOR2X1 \mult_97/U1470  ( .A(n340), .B(n277), .Y(\mult_97/n2478 ) );
  OAI22X1 \mult_97/U1469  ( .A(\mult_97/n2508 ), .B(n328), .C(\mult_97/n2509 ), 
        .D(n250), .Y(\mult_97/n1988 ) );
  OAI22X1 \mult_97/U1468  ( .A(\mult_97/n2507 ), .B(n328), .C(\mult_97/n2508 ), 
        .D(n250), .Y(\mult_97/n1987 ) );
  OAI22X1 \mult_97/U1467  ( .A(\mult_97/n2506 ), .B(n328), .C(\mult_97/n2507 ), 
        .D(n250), .Y(\mult_97/n1986 ) );
  OAI22X1 \mult_97/U1466  ( .A(\mult_97/n2505 ), .B(n328), .C(\mult_97/n2506 ), 
        .D(n250), .Y(\mult_97/n1985 ) );
  OAI22X1 \mult_97/U1465  ( .A(\mult_97/n2504 ), .B(n328), .C(\mult_97/n2505 ), 
        .D(n250), .Y(\mult_97/n1984 ) );
  OAI22X1 \mult_97/U1464  ( .A(\mult_97/n2503 ), .B(n328), .C(\mult_97/n2504 ), 
        .D(n250), .Y(\mult_97/n1983 ) );
  OAI22X1 \mult_97/U1463  ( .A(\mult_97/n2502 ), .B(n328), .C(\mult_97/n2503 ), 
        .D(n250), .Y(\mult_97/n1982 ) );
  OAI22X1 \mult_97/U1462  ( .A(\mult_97/n2501 ), .B(n328), .C(\mult_97/n2502 ), 
        .D(n250), .Y(\mult_97/n1981 ) );
  OAI22X1 \mult_97/U1461  ( .A(\mult_97/n2500 ), .B(n328), .C(\mult_97/n2501 ), 
        .D(n250), .Y(\mult_97/n1980 ) );
  OAI22X1 \mult_97/U1460  ( .A(\mult_97/n2499 ), .B(n328), .C(\mult_97/n2500 ), 
        .D(n250), .Y(\mult_97/n1979 ) );
  OAI22X1 \mult_97/U1459  ( .A(\mult_97/n2498 ), .B(n328), .C(\mult_97/n2499 ), 
        .D(n250), .Y(\mult_97/n1978 ) );
  OAI22X1 \mult_97/U1458  ( .A(\mult_97/n2497 ), .B(n328), .C(\mult_97/n2498 ), 
        .D(n250), .Y(\mult_97/n1977 ) );
  OAI22X1 \mult_97/U1457  ( .A(\mult_97/n2496 ), .B(n328), .C(\mult_97/n2497 ), 
        .D(n250), .Y(\mult_97/n1976 ) );
  OAI22X1 \mult_97/U1456  ( .A(\mult_97/n2495 ), .B(n328), .C(\mult_97/n2496 ), 
        .D(n250), .Y(\mult_97/n1975 ) );
  OAI22X1 \mult_97/U1455  ( .A(\mult_97/n2494 ), .B(n328), .C(\mult_97/n2495 ), 
        .D(n250), .Y(\mult_97/n1974 ) );
  OAI22X1 \mult_97/U1454  ( .A(\mult_97/n2493 ), .B(n328), .C(\mult_97/n2494 ), 
        .D(n250), .Y(\mult_97/n1973 ) );
  OAI22X1 \mult_97/U1453  ( .A(\mult_97/n2492 ), .B(n328), .C(\mult_97/n2493 ), 
        .D(n250), .Y(\mult_97/n1161 ) );
  OAI22X1 \mult_97/U1452  ( .A(\mult_97/n2491 ), .B(n328), .C(\mult_97/n2492 ), 
        .D(n250), .Y(\mult_97/n1972 ) );
  OAI22X1 \mult_97/U1451  ( .A(\mult_97/n2490 ), .B(n328), .C(\mult_97/n2491 ), 
        .D(n250), .Y(\mult_97/n1971 ) );
  OAI22X1 \mult_97/U1450  ( .A(\mult_97/n2489 ), .B(n328), .C(\mult_97/n2490 ), 
        .D(n250), .Y(\mult_97/n1970 ) );
  OAI22X1 \mult_97/U1449  ( .A(\mult_97/n2488 ), .B(n328), .C(\mult_97/n2489 ), 
        .D(n250), .Y(\mult_97/n1081 ) );
  OAI22X1 \mult_97/U1448  ( .A(\mult_97/n2487 ), .B(n328), .C(\mult_97/n2488 ), 
        .D(n250), .Y(\mult_97/n1969 ) );
  OAI22X1 \mult_97/U1447  ( .A(\mult_97/n2486 ), .B(n328), .C(\mult_97/n2487 ), 
        .D(n250), .Y(\mult_97/n1047 ) );
  OAI22X1 \mult_97/U1446  ( .A(\mult_97/n2485 ), .B(n328), .C(\mult_97/n2486 ), 
        .D(n250), .Y(\mult_97/n1968 ) );
  OAI22X1 \mult_97/U1445  ( .A(\mult_97/n2484 ), .B(n328), .C(\mult_97/n2485 ), 
        .D(n250), .Y(\mult_97/n1967 ) );
  OAI22X1 \mult_97/U1444  ( .A(\mult_97/n2483 ), .B(n328), .C(\mult_97/n2484 ), 
        .D(n250), .Y(\mult_97/n1966 ) );
  OAI22X1 \mult_97/U1443  ( .A(\mult_97/n2482 ), .B(n328), .C(\mult_97/n2483 ), 
        .D(n250), .Y(\mult_97/n991 ) );
  OAI22X1 \mult_97/U1442  ( .A(\mult_97/n2481 ), .B(n328), .C(\mult_97/n2482 ), 
        .D(n250), .Y(\mult_97/n1965 ) );
  OAI22X1 \mult_97/U1441  ( .A(\mult_97/n2480 ), .B(n328), .C(\mult_97/n2481 ), 
        .D(n250), .Y(\mult_97/n969 ) );
  OAI22X1 \mult_97/U1440  ( .A(\mult_97/n2479 ), .B(n328), .C(\mult_97/n2480 ), 
        .D(n250), .Y(\mult_97/n1964 ) );
  OAI22X1 \mult_97/U1439  ( .A(\mult_97/n2478 ), .B(n328), .C(\mult_97/n2479 ), 
        .D(n250), .Y(\mult_97/n951 ) );
  OAI22X1 \mult_97/U1438  ( .A(n328), .B(\mult_97/n2510 ), .C(n275), .D(n250), 
        .Y(\mult_97/n1854 ) );
  XNOR2X1 \mult_97/U1437  ( .A(n251), .B(n274), .Y(\mult_97/n2476 ) );
  XNOR2X1 \mult_97/U1436  ( .A(n400), .B(n274), .Y(\mult_97/n2475 ) );
  XNOR2X1 \mult_97/U1435  ( .A(n398), .B(n274), .Y(\mult_97/n2474 ) );
  XNOR2X1 \mult_97/U1434  ( .A(n396), .B(n274), .Y(\mult_97/n2473 ) );
  XNOR2X1 \mult_97/U1433  ( .A(n394), .B(n274), .Y(\mult_97/n2472 ) );
  XNOR2X1 \mult_97/U1432  ( .A(n392), .B(n274), .Y(\mult_97/n2471 ) );
  XNOR2X1 \mult_97/U1431  ( .A(n390), .B(n274), .Y(\mult_97/n2470 ) );
  XNOR2X1 \mult_97/U1430  ( .A(n388), .B(n274), .Y(\mult_97/n2469 ) );
  XNOR2X1 \mult_97/U1429  ( .A(n386), .B(n274), .Y(\mult_97/n2468 ) );
  XNOR2X1 \mult_97/U1428  ( .A(B[9]), .B(A[27]), .Y(\mult_97/n2467 ) );
  XNOR2X1 \mult_97/U1427  ( .A(B[10]), .B(n274), .Y(\mult_97/n2466 ) );
  XNOR2X1 \mult_97/U1426  ( .A(n380), .B(n274), .Y(\mult_97/n2465 ) );
  XNOR2X1 \mult_97/U1425  ( .A(n378), .B(n274), .Y(\mult_97/n2464 ) );
  XNOR2X1 \mult_97/U1424  ( .A(n376), .B(n274), .Y(\mult_97/n2463 ) );
  XNOR2X1 \mult_97/U1423  ( .A(n374), .B(n274), .Y(\mult_97/n2462 ) );
  XNOR2X1 \mult_97/U1422  ( .A(n372), .B(n274), .Y(\mult_97/n2461 ) );
  XNOR2X1 \mult_97/U1421  ( .A(n370), .B(n274), .Y(\mult_97/n2460 ) );
  XNOR2X1 \mult_97/U1420  ( .A(n368), .B(n274), .Y(\mult_97/n2459 ) );
  XNOR2X1 \mult_97/U1419  ( .A(B[18]), .B(n274), .Y(\mult_97/n2458 ) );
  XNOR2X1 \mult_97/U1418  ( .A(n364), .B(n274), .Y(\mult_97/n2457 ) );
  XNOR2X1 \mult_97/U1417  ( .A(n362), .B(n274), .Y(\mult_97/n2456 ) );
  XNOR2X1 \mult_97/U1416  ( .A(n360), .B(n274), .Y(\mult_97/n2455 ) );
  XNOR2X1 \mult_97/U1415  ( .A(n358), .B(n274), .Y(\mult_97/n2454 ) );
  XNOR2X1 \mult_97/U1414  ( .A(n356), .B(n274), .Y(\mult_97/n2453 ) );
  XNOR2X1 \mult_97/U1413  ( .A(n354), .B(n274), .Y(\mult_97/n2452 ) );
  XNOR2X1 \mult_97/U1412  ( .A(n352), .B(n274), .Y(\mult_97/n2451 ) );
  XNOR2X1 \mult_97/U1411  ( .A(n350), .B(n274), .Y(\mult_97/n2450 ) );
  XNOR2X1 \mult_97/U1410  ( .A(n348), .B(n274), .Y(\mult_97/n2449 ) );
  XNOR2X1 \mult_97/U1409  ( .A(n346), .B(n274), .Y(\mult_97/n2448 ) );
  XNOR2X1 \mult_97/U1408  ( .A(n344), .B(n274), .Y(\mult_97/n2447 ) );
  XNOR2X1 \mult_97/U1407  ( .A(n342), .B(n274), .Y(\mult_97/n2446 ) );
  XNOR2X1 \mult_97/U1406  ( .A(n340), .B(A[27]), .Y(\mult_97/n2445 ) );
  OAI22X1 \mult_97/U1405  ( .A(\mult_97/n2475 ), .B(n329), .C(\mult_97/n2476 ), 
        .D(n338), .Y(\mult_97/n1961 ) );
  OAI22X1 \mult_97/U1404  ( .A(\mult_97/n2474 ), .B(n329), .C(\mult_97/n2475 ), 
        .D(n338), .Y(\mult_97/n1960 ) );
  OAI22X1 \mult_97/U1403  ( .A(\mult_97/n2473 ), .B(n329), .C(\mult_97/n2474 ), 
        .D(n338), .Y(\mult_97/n1959 ) );
  OAI22X1 \mult_97/U1402  ( .A(\mult_97/n2472 ), .B(n329), .C(\mult_97/n2473 ), 
        .D(n338), .Y(\mult_97/n1958 ) );
  OAI22X1 \mult_97/U1401  ( .A(\mult_97/n2471 ), .B(n329), .C(\mult_97/n2472 ), 
        .D(n338), .Y(\mult_97/n1957 ) );
  OAI22X1 \mult_97/U1400  ( .A(\mult_97/n2470 ), .B(n329), .C(\mult_97/n2471 ), 
        .D(n338), .Y(\mult_97/n1956 ) );
  OAI22X1 \mult_97/U1399  ( .A(\mult_97/n2469 ), .B(n329), .C(\mult_97/n2470 ), 
        .D(n338), .Y(\mult_97/n1955 ) );
  OAI22X1 \mult_97/U1398  ( .A(\mult_97/n2468 ), .B(n329), .C(\mult_97/n2469 ), 
        .D(n338), .Y(\mult_97/n1954 ) );
  OAI22X1 \mult_97/U1397  ( .A(\mult_97/n2467 ), .B(n329), .C(\mult_97/n2468 ), 
        .D(n338), .Y(\mult_97/n1953 ) );
  OAI22X1 \mult_97/U1396  ( .A(\mult_97/n2466 ), .B(n329), .C(\mult_97/n2467 ), 
        .D(n338), .Y(\mult_97/n1952 ) );
  OAI22X1 \mult_97/U1395  ( .A(\mult_97/n2465 ), .B(n329), .C(\mult_97/n2466 ), 
        .D(n338), .Y(\mult_97/n1951 ) );
  OAI22X1 \mult_97/U1394  ( .A(\mult_97/n2464 ), .B(n329), .C(\mult_97/n2465 ), 
        .D(n338), .Y(\mult_97/n1950 ) );
  OAI22X1 \mult_97/U1393  ( .A(\mult_97/n2463 ), .B(n329), .C(\mult_97/n2464 ), 
        .D(n338), .Y(\mult_97/n1949 ) );
  OAI22X1 \mult_97/U1392  ( .A(\mult_97/n2462 ), .B(n329), .C(\mult_97/n2463 ), 
        .D(n338), .Y(\mult_97/n1948 ) );
  OAI22X1 \mult_97/U1391  ( .A(\mult_97/n2461 ), .B(n329), .C(\mult_97/n2462 ), 
        .D(n338), .Y(\mult_97/n1947 ) );
  OAI22X1 \mult_97/U1390  ( .A(\mult_97/n2460 ), .B(n329), .C(\mult_97/n2461 ), 
        .D(n338), .Y(\mult_97/n1946 ) );
  OAI22X1 \mult_97/U1389  ( .A(\mult_97/n2459 ), .B(n329), .C(\mult_97/n2460 ), 
        .D(n338), .Y(\mult_97/n1945 ) );
  OAI22X1 \mult_97/U1388  ( .A(\mult_97/n2458 ), .B(n329), .C(\mult_97/n2459 ), 
        .D(n338), .Y(\mult_97/n1944 ) );
  OAI22X1 \mult_97/U1387  ( .A(\mult_97/n2457 ), .B(n329), .C(\mult_97/n2458 ), 
        .D(n338), .Y(\mult_97/n1943 ) );
  OAI22X1 \mult_97/U1386  ( .A(\mult_97/n2456 ), .B(n329), .C(\mult_97/n2457 ), 
        .D(n338), .Y(\mult_97/n1942 ) );
  OAI22X1 \mult_97/U1385  ( .A(\mult_97/n2455 ), .B(n329), .C(\mult_97/n2456 ), 
        .D(n338), .Y(\mult_97/n1941 ) );
  OAI22X1 \mult_97/U1384  ( .A(\mult_97/n2454 ), .B(n329), .C(\mult_97/n2455 ), 
        .D(n338), .Y(\mult_97/n1940 ) );
  OAI22X1 \mult_97/U1383  ( .A(\mult_97/n2453 ), .B(n329), .C(\mult_97/n2454 ), 
        .D(n338), .Y(\mult_97/n1939 ) );
  OAI22X1 \mult_97/U1382  ( .A(\mult_97/n2452 ), .B(n329), .C(\mult_97/n2453 ), 
        .D(n338), .Y(\mult_97/n1938 ) );
  OAI22X1 \mult_97/U1381  ( .A(\mult_97/n2451 ), .B(n329), .C(\mult_97/n2452 ), 
        .D(n338), .Y(\mult_97/n1937 ) );
  OAI22X1 \mult_97/U1380  ( .A(\mult_97/n2450 ), .B(n329), .C(\mult_97/n2451 ), 
        .D(n338), .Y(\mult_97/n1936 ) );
  OAI22X1 \mult_97/U1379  ( .A(\mult_97/n2449 ), .B(n329), .C(\mult_97/n2450 ), 
        .D(n338), .Y(\mult_97/n1935 ) );
  OAI22X1 \mult_97/U1378  ( .A(\mult_97/n2448 ), .B(n329), .C(\mult_97/n2449 ), 
        .D(n338), .Y(\mult_97/n1934 ) );
  OAI22X1 \mult_97/U1377  ( .A(\mult_97/n2447 ), .B(n329), .C(\mult_97/n2448 ), 
        .D(n338), .Y(\mult_97/n1933 ) );
  OAI22X1 \mult_97/U1376  ( .A(\mult_97/n2446 ), .B(n329), .C(\mult_97/n2447 ), 
        .D(n338), .Y(\mult_97/n1932 ) );
  OAI22X1 \mult_97/U1375  ( .A(\mult_97/n2445 ), .B(n329), .C(\mult_97/n2446 ), 
        .D(n338), .Y(\mult_97/n1931 ) );
  OAI22X1 \mult_97/U1374  ( .A(n329), .B(\mult_97/n2477 ), .C(n273), .D(n338), 
        .Y(\mult_97/n1853 ) );
  XNOR2X1 \mult_97/U1373  ( .A(n272), .B(n251), .Y(\mult_97/n2443 ) );
  XNOR2X1 \mult_97/U1372  ( .A(n272), .B(n400), .Y(\mult_97/n2442 ) );
  XNOR2X1 \mult_97/U1371  ( .A(n272), .B(n398), .Y(\mult_97/n2441 ) );
  XNOR2X1 \mult_97/U1370  ( .A(n272), .B(n396), .Y(\mult_97/n2440 ) );
  XNOR2X1 \mult_97/U1369  ( .A(n272), .B(n394), .Y(\mult_97/n2439 ) );
  XNOR2X1 \mult_97/U1368  ( .A(n272), .B(n392), .Y(\mult_97/n2438 ) );
  XNOR2X1 \mult_97/U1367  ( .A(n272), .B(n390), .Y(\mult_97/n2437 ) );
  XNOR2X1 \mult_97/U1366  ( .A(n272), .B(n388), .Y(\mult_97/n2436 ) );
  XNOR2X1 \mult_97/U1365  ( .A(n272), .B(n386), .Y(\mult_97/n2435 ) );
  XNOR2X1 \mult_97/U1364  ( .A(n272), .B(n384), .Y(\mult_97/n2434 ) );
  XNOR2X1 \mult_97/U1363  ( .A(n272), .B(n382), .Y(\mult_97/n2433 ) );
  XNOR2X1 \mult_97/U1362  ( .A(n272), .B(n380), .Y(\mult_97/n2432 ) );
  XNOR2X1 \mult_97/U1361  ( .A(n272), .B(n378), .Y(\mult_97/n2431 ) );
  XNOR2X1 \mult_97/U1360  ( .A(n272), .B(n376), .Y(\mult_97/n2430 ) );
  XNOR2X1 \mult_97/U1359  ( .A(n272), .B(n374), .Y(\mult_97/n2429 ) );
  XNOR2X1 \mult_97/U1358  ( .A(n272), .B(n372), .Y(\mult_97/n2428 ) );
  XNOR2X1 \mult_97/U1357  ( .A(n272), .B(n370), .Y(\mult_97/n2427 ) );
  XNOR2X1 \mult_97/U1356  ( .A(n272), .B(n368), .Y(\mult_97/n2426 ) );
  XNOR2X1 \mult_97/U1355  ( .A(n272), .B(n366), .Y(\mult_97/n2425 ) );
  XNOR2X1 \mult_97/U1354  ( .A(n272), .B(n364), .Y(\mult_97/n2424 ) );
  XNOR2X1 \mult_97/U1353  ( .A(n272), .B(n362), .Y(\mult_97/n2423 ) );
  XNOR2X1 \mult_97/U1352  ( .A(n272), .B(n360), .Y(\mult_97/n2422 ) );
  XNOR2X1 \mult_97/U1351  ( .A(n272), .B(n358), .Y(\mult_97/n2421 ) );
  XNOR2X1 \mult_97/U1350  ( .A(n272), .B(n356), .Y(\mult_97/n2420 ) );
  XNOR2X1 \mult_97/U1349  ( .A(n272), .B(n354), .Y(\mult_97/n2419 ) );
  XNOR2X1 \mult_97/U1348  ( .A(n272), .B(n352), .Y(\mult_97/n2418 ) );
  XNOR2X1 \mult_97/U1347  ( .A(n272), .B(n350), .Y(\mult_97/n2417 ) );
  XNOR2X1 \mult_97/U1346  ( .A(n272), .B(n348), .Y(\mult_97/n2416 ) );
  XNOR2X1 \mult_97/U1345  ( .A(n272), .B(n346), .Y(\mult_97/n2415 ) );
  XNOR2X1 \mult_97/U1344  ( .A(n272), .B(n344), .Y(\mult_97/n2414 ) );
  XNOR2X1 \mult_97/U1343  ( .A(n272), .B(n342), .Y(\mult_97/n2413 ) );
  XNOR2X1 \mult_97/U1342  ( .A(n272), .B(n340), .Y(\mult_97/n2412 ) );
  OAI22X1 \mult_97/U1341  ( .A(n330), .B(\mult_97/n2442 ), .C(\mult_97/n2443 ), 
        .D(n248), .Y(\mult_97/n1928 ) );
  OAI22X1 \mult_97/U1340  ( .A(n330), .B(\mult_97/n2441 ), .C(\mult_97/n2442 ), 
        .D(n248), .Y(\mult_97/n1927 ) );
  OAI22X1 \mult_97/U1339  ( .A(n330), .B(\mult_97/n2440 ), .C(\mult_97/n2441 ), 
        .D(n248), .Y(\mult_97/n1926 ) );
  OAI22X1 \mult_97/U1338  ( .A(n330), .B(\mult_97/n2439 ), .C(\mult_97/n2440 ), 
        .D(n248), .Y(\mult_97/n1925 ) );
  OAI22X1 \mult_97/U1337  ( .A(n330), .B(\mult_97/n2438 ), .C(\mult_97/n2439 ), 
        .D(n248), .Y(\mult_97/n1924 ) );
  OAI22X1 \mult_97/U1336  ( .A(n330), .B(\mult_97/n2437 ), .C(\mult_97/n2438 ), 
        .D(n248), .Y(\mult_97/n1923 ) );
  OAI22X1 \mult_97/U1335  ( .A(n330), .B(\mult_97/n2436 ), .C(\mult_97/n2437 ), 
        .D(n248), .Y(\mult_97/n1922 ) );
  OAI22X1 \mult_97/U1334  ( .A(n330), .B(\mult_97/n2435 ), .C(\mult_97/n2436 ), 
        .D(n248), .Y(\mult_97/n1921 ) );
  OAI22X1 \mult_97/U1333  ( .A(n330), .B(\mult_97/n2434 ), .C(\mult_97/n2435 ), 
        .D(n248), .Y(\mult_97/n1920 ) );
  OAI22X1 \mult_97/U1332  ( .A(n330), .B(\mult_97/n2433 ), .C(\mult_97/n2434 ), 
        .D(n248), .Y(\mult_97/n1919 ) );
  OAI22X1 \mult_97/U1331  ( .A(n330), .B(\mult_97/n2432 ), .C(\mult_97/n2433 ), 
        .D(n248), .Y(\mult_97/n1918 ) );
  OAI22X1 \mult_97/U1330  ( .A(n330), .B(\mult_97/n2431 ), .C(\mult_97/n2432 ), 
        .D(n248), .Y(\mult_97/n1917 ) );
  OAI22X1 \mult_97/U1329  ( .A(n330), .B(\mult_97/n2430 ), .C(\mult_97/n2431 ), 
        .D(n248), .Y(\mult_97/n1916 ) );
  OAI22X1 \mult_97/U1328  ( .A(n330), .B(\mult_97/n2429 ), .C(\mult_97/n2430 ), 
        .D(n248), .Y(\mult_97/n1915 ) );
  OAI22X1 \mult_97/U1327  ( .A(n330), .B(\mult_97/n2428 ), .C(\mult_97/n2429 ), 
        .D(n248), .Y(\mult_97/n1914 ) );
  OAI22X1 \mult_97/U1326  ( .A(n330), .B(\mult_97/n2427 ), .C(\mult_97/n2428 ), 
        .D(n248), .Y(\mult_97/n1913 ) );
  OAI22X1 \mult_97/U1325  ( .A(n330), .B(\mult_97/n2426 ), .C(\mult_97/n2427 ), 
        .D(n248), .Y(\mult_97/n1912 ) );
  OAI22X1 \mult_97/U1324  ( .A(n330), .B(\mult_97/n2425 ), .C(\mult_97/n2426 ), 
        .D(n248), .Y(\mult_97/n1911 ) );
  OAI22X1 \mult_97/U1323  ( .A(n330), .B(\mult_97/n2424 ), .C(\mult_97/n2425 ), 
        .D(n248), .Y(\mult_97/n1910 ) );
  OAI22X1 \mult_97/U1322  ( .A(n330), .B(\mult_97/n2423 ), .C(\mult_97/n2424 ), 
        .D(n248), .Y(\mult_97/n1909 ) );
  OAI22X1 \mult_97/U1321  ( .A(n330), .B(\mult_97/n2422 ), .C(\mult_97/n2423 ), 
        .D(n248), .Y(\mult_97/n1908 ) );
  OAI22X1 \mult_97/U1320  ( .A(n330), .B(\mult_97/n2421 ), .C(\mult_97/n2422 ), 
        .D(n248), .Y(\mult_97/n1907 ) );
  OAI22X1 \mult_97/U1319  ( .A(n330), .B(\mult_97/n2420 ), .C(\mult_97/n2421 ), 
        .D(n248), .Y(\mult_97/n1906 ) );
  OAI22X1 \mult_97/U1318  ( .A(n330), .B(\mult_97/n2419 ), .C(\mult_97/n2420 ), 
        .D(n248), .Y(\mult_97/n1905 ) );
  OAI22X1 \mult_97/U1317  ( .A(n330), .B(\mult_97/n2418 ), .C(\mult_97/n2419 ), 
        .D(n248), .Y(\mult_97/n1904 ) );
  OAI22X1 \mult_97/U1316  ( .A(n330), .B(\mult_97/n2417 ), .C(\mult_97/n2418 ), 
        .D(n248), .Y(\mult_97/n1903 ) );
  OAI22X1 \mult_97/U1315  ( .A(n330), .B(\mult_97/n2416 ), .C(\mult_97/n2417 ), 
        .D(n248), .Y(\mult_97/n1902 ) );
  OAI22X1 \mult_97/U1314  ( .A(n330), .B(\mult_97/n2415 ), .C(\mult_97/n2416 ), 
        .D(n248), .Y(\mult_97/n1901 ) );
  OAI22X1 \mult_97/U1313  ( .A(n330), .B(\mult_97/n2414 ), .C(\mult_97/n2415 ), 
        .D(n248), .Y(\mult_97/n937 ) );
  OAI22X1 \mult_97/U1312  ( .A(n330), .B(\mult_97/n2413 ), .C(\mult_97/n2414 ), 
        .D(n248), .Y(\mult_97/n1900 ) );
  OAI22X1 \mult_97/U1311  ( .A(n330), .B(\mult_97/n2412 ), .C(\mult_97/n2413 ), 
        .D(n248), .Y(\mult_97/n927 ) );
  OAI22X1 \mult_97/U1310  ( .A(n330), .B(\mult_97/n2444 ), .C(n271), .D(n248), 
        .Y(\mult_97/n1852 ) );
  XNOR2X1 \mult_97/U1309  ( .A(n270), .B(n251), .Y(\mult_97/n2410 ) );
  XNOR2X1 \mult_97/U1308  ( .A(n270), .B(n400), .Y(\mult_97/n2409 ) );
  XNOR2X1 \mult_97/U1307  ( .A(n270), .B(n398), .Y(\mult_97/n2408 ) );
  XNOR2X1 \mult_97/U1306  ( .A(n270), .B(n396), .Y(\mult_97/n2407 ) );
  XNOR2X1 \mult_97/U1305  ( .A(n270), .B(n394), .Y(\mult_97/n2406 ) );
  XNOR2X1 \mult_97/U1304  ( .A(n270), .B(n392), .Y(\mult_97/n2405 ) );
  XNOR2X1 \mult_97/U1303  ( .A(n270), .B(n390), .Y(\mult_97/n2404 ) );
  XNOR2X1 \mult_97/U1302  ( .A(n270), .B(n388), .Y(\mult_97/n2403 ) );
  XNOR2X1 \mult_97/U1301  ( .A(n270), .B(n386), .Y(\mult_97/n2402 ) );
  XNOR2X1 \mult_97/U1300  ( .A(n270), .B(n384), .Y(\mult_97/n2401 ) );
  XNOR2X1 \mult_97/U1299  ( .A(n270), .B(n382), .Y(\mult_97/n2400 ) );
  XNOR2X1 \mult_97/U1298  ( .A(n270), .B(n380), .Y(\mult_97/n2399 ) );
  XNOR2X1 \mult_97/U1297  ( .A(n269), .B(n378), .Y(\mult_97/n2398 ) );
  XNOR2X1 \mult_97/U1296  ( .A(n269), .B(n376), .Y(\mult_97/n2397 ) );
  XNOR2X1 \mult_97/U1295  ( .A(n269), .B(n374), .Y(\mult_97/n2396 ) );
  XNOR2X1 \mult_97/U1294  ( .A(n269), .B(n372), .Y(\mult_97/n2395 ) );
  XNOR2X1 \mult_97/U1293  ( .A(n269), .B(n370), .Y(\mult_97/n2394 ) );
  XNOR2X1 \mult_97/U1292  ( .A(n269), .B(n368), .Y(\mult_97/n2393 ) );
  XNOR2X1 \mult_97/U1291  ( .A(n269), .B(n366), .Y(\mult_97/n2392 ) );
  XNOR2X1 \mult_97/U1290  ( .A(n269), .B(n364), .Y(\mult_97/n2391 ) );
  XNOR2X1 \mult_97/U1289  ( .A(n269), .B(n362), .Y(\mult_97/n2390 ) );
  XNOR2X1 \mult_97/U1288  ( .A(n269), .B(n360), .Y(\mult_97/n2389 ) );
  XNOR2X1 \mult_97/U1287  ( .A(n269), .B(n358), .Y(\mult_97/n2388 ) );
  XNOR2X1 \mult_97/U1286  ( .A(n269), .B(n356), .Y(\mult_97/n2387 ) );
  XNOR2X1 \mult_97/U1285  ( .A(n270), .B(n354), .Y(\mult_97/n2386 ) );
  XNOR2X1 \mult_97/U1284  ( .A(n270), .B(n352), .Y(\mult_97/n2385 ) );
  XNOR2X1 \mult_97/U1283  ( .A(n270), .B(n350), .Y(\mult_97/n2384 ) );
  XNOR2X1 \mult_97/U1282  ( .A(n270), .B(n348), .Y(\mult_97/n2383 ) );
  XNOR2X1 \mult_97/U1281  ( .A(n270), .B(n346), .Y(\mult_97/n2382 ) );
  XNOR2X1 \mult_97/U1280  ( .A(n270), .B(n344), .Y(\mult_97/n2381 ) );
  XNOR2X1 \mult_97/U1279  ( .A(n270), .B(n342), .Y(\mult_97/n2380 ) );
  XNOR2X1 \mult_97/U1278  ( .A(n270), .B(n340), .Y(\mult_97/n2379 ) );
  OAI22X1 \mult_97/U1277  ( .A(\mult_97/n2409 ), .B(n331), .C(\mult_97/n2410 ), 
        .D(n339), .Y(\mult_97/n1897 ) );
  OAI22X1 \mult_97/U1276  ( .A(\mult_97/n2408 ), .B(n331), .C(\mult_97/n2409 ), 
        .D(n339), .Y(\mult_97/n1896 ) );
  OAI22X1 \mult_97/U1275  ( .A(\mult_97/n2407 ), .B(n331), .C(\mult_97/n2408 ), 
        .D(n339), .Y(\mult_97/n1895 ) );
  OAI22X1 \mult_97/U1274  ( .A(\mult_97/n2406 ), .B(n331), .C(\mult_97/n2407 ), 
        .D(n339), .Y(\mult_97/n1894 ) );
  OAI22X1 \mult_97/U1273  ( .A(\mult_97/n2405 ), .B(n331), .C(\mult_97/n2406 ), 
        .D(n339), .Y(\mult_97/n1893 ) );
  OAI22X1 \mult_97/U1272  ( .A(\mult_97/n2404 ), .B(n331), .C(\mult_97/n2405 ), 
        .D(n339), .Y(\mult_97/n1892 ) );
  OAI22X1 \mult_97/U1271  ( .A(\mult_97/n2403 ), .B(n331), .C(\mult_97/n2404 ), 
        .D(n339), .Y(\mult_97/n1891 ) );
  OAI22X1 \mult_97/U1270  ( .A(\mult_97/n2402 ), .B(n331), .C(\mult_97/n2403 ), 
        .D(n339), .Y(\mult_97/n1890 ) );
  OAI22X1 \mult_97/U1269  ( .A(\mult_97/n2401 ), .B(n331), .C(\mult_97/n2402 ), 
        .D(n339), .Y(\mult_97/n1889 ) );
  OAI22X1 \mult_97/U1268  ( .A(\mult_97/n2400 ), .B(n331), .C(\mult_97/n2401 ), 
        .D(n339), .Y(\mult_97/n1888 ) );
  OAI22X1 \mult_97/U1267  ( .A(\mult_97/n2399 ), .B(n331), .C(\mult_97/n2400 ), 
        .D(n339), .Y(\mult_97/n1887 ) );
  OAI22X1 \mult_97/U1266  ( .A(\mult_97/n2398 ), .B(n331), .C(\mult_97/n2399 ), 
        .D(n339), .Y(\mult_97/n1886 ) );
  OAI22X1 \mult_97/U1265  ( .A(\mult_97/n2397 ), .B(n331), .C(\mult_97/n2398 ), 
        .D(n339), .Y(\mult_97/n1885 ) );
  OAI22X1 \mult_97/U1264  ( .A(\mult_97/n2396 ), .B(n331), .C(\mult_97/n2397 ), 
        .D(n339), .Y(\mult_97/n1884 ) );
  OAI22X1 \mult_97/U1263  ( .A(\mult_97/n2395 ), .B(n331), .C(\mult_97/n2396 ), 
        .D(n339), .Y(\mult_97/n1883 ) );
  OAI22X1 \mult_97/U1262  ( .A(\mult_97/n2394 ), .B(n331), .C(\mult_97/n2395 ), 
        .D(n339), .Y(\mult_97/n1882 ) );
  OAI22X1 \mult_97/U1261  ( .A(\mult_97/n2393 ), .B(n331), .C(\mult_97/n2394 ), 
        .D(n339), .Y(\mult_97/n1881 ) );
  OAI22X1 \mult_97/U1260  ( .A(\mult_97/n2392 ), .B(n331), .C(\mult_97/n2393 ), 
        .D(n339), .Y(\mult_97/n1880 ) );
  OAI22X1 \mult_97/U1259  ( .A(\mult_97/n2391 ), .B(n331), .C(\mult_97/n2392 ), 
        .D(n339), .Y(\mult_97/n1879 ) );
  OAI22X1 \mult_97/U1258  ( .A(\mult_97/n2390 ), .B(n331), .C(\mult_97/n2391 ), 
        .D(n339), .Y(\mult_97/n1878 ) );
  OAI22X1 \mult_97/U1257  ( .A(\mult_97/n2389 ), .B(n331), .C(\mult_97/n2390 ), 
        .D(n339), .Y(\mult_97/n1877 ) );
  OAI22X1 \mult_97/U1256  ( .A(\mult_97/n2388 ), .B(n331), .C(\mult_97/n2389 ), 
        .D(n339), .Y(\mult_97/n1876 ) );
  OAI22X1 \mult_97/U1255  ( .A(\mult_97/n2387 ), .B(n331), .C(\mult_97/n2388 ), 
        .D(n339), .Y(\mult_97/n1875 ) );
  OAI22X1 \mult_97/U1254  ( .A(\mult_97/n2386 ), .B(n331), .C(\mult_97/n2387 ), 
        .D(n339), .Y(\mult_97/n1874 ) );
  OAI22X1 \mult_97/U1253  ( .A(\mult_97/n2385 ), .B(n331), .C(\mult_97/n2386 ), 
        .D(n339), .Y(\mult_97/n1873 ) );
  OAI22X1 \mult_97/U1252  ( .A(\mult_97/n2384 ), .B(n331), .C(\mult_97/n2385 ), 
        .D(n339), .Y(\mult_97/n1872 ) );
  OAI22X1 \mult_97/U1251  ( .A(\mult_97/n2383 ), .B(n331), .C(\mult_97/n2384 ), 
        .D(n339), .Y(\mult_97/n1871 ) );
  OAI22X1 \mult_97/U1250  ( .A(\mult_97/n2382 ), .B(n331), .C(\mult_97/n2383 ), 
        .D(n339), .Y(\mult_97/n1870 ) );
  OAI22X1 \mult_97/U1249  ( .A(\mult_97/n2381 ), .B(n331), .C(\mult_97/n2382 ), 
        .D(n339), .Y(\mult_97/n1869 ) );
  OAI22X1 \mult_97/U1248  ( .A(\mult_97/n2380 ), .B(n331), .C(\mult_97/n2381 ), 
        .D(n339), .Y(\mult_97/n1868 ) );
  OAI22X1 \mult_97/U1247  ( .A(n331), .B(\mult_97/n2379 ), .C(\mult_97/n2380 ), 
        .D(n339), .Y(\mult_97/n921 ) );
  OAI22X1 \mult_97/U1246  ( .A(n331), .B(\mult_97/n2411 ), .C(n268), .D(n339), 
        .Y(\mult_97/n1851 ) );
  HAX1 \mult_97/U1245  ( .A(\mult_97/n2376 ), .B(\mult_97/n2345 ), .YC(
        \mult_97/n1849 ), .YS(\mult_97/n1850 ) );
  FAX1 \mult_97/U1244  ( .A(\mult_97/n2375 ), .B(\mult_97/n2313 ), .C(
        \mult_97/n2344 ), .YC(\mult_97/n1847 ), .YS(\mult_97/n1848 ) );
  HAX1 \mult_97/U1243  ( .A(\mult_97/n2374 ), .B(\mult_97/n1864 ), .YC(
        \mult_97/n1845 ), .YS(\mult_97/n1846 ) );
  FAX1 \mult_97/U1242  ( .A(\mult_97/n2312 ), .B(\mult_97/n2343 ), .C(
        \mult_97/n1846 ), .YC(\mult_97/n1843 ), .YS(\mult_97/n1844 ) );
  FAX1 \mult_97/U1241  ( .A(\mult_97/n2373 ), .B(\mult_97/n2311 ), .C(
        \mult_97/n2342 ), .YC(\mult_97/n1841 ), .YS(\mult_97/n1842 ) );
  FAX1 \mult_97/U1240  ( .A(\mult_97/n2280 ), .B(\mult_97/n1845 ), .C(
        \mult_97/n1842 ), .YC(\mult_97/n1839 ), .YS(\mult_97/n1840 ) );
  HAX1 \mult_97/U1239  ( .A(\mult_97/n2372 ), .B(\mult_97/n1863 ), .YC(
        \mult_97/n1837 ), .YS(\mult_97/n1838 ) );
  FAX1 \mult_97/U1238  ( .A(\mult_97/n2279 ), .B(\mult_97/n2310 ), .C(
        \mult_97/n2341 ), .YC(\mult_97/n1835 ), .YS(\mult_97/n1836 ) );
  FAX1 \mult_97/U1237  ( .A(\mult_97/n1838 ), .B(\mult_97/n1841 ), .C(
        \mult_97/n1836 ), .YC(\mult_97/n1833 ), .YS(\mult_97/n1834 ) );
  FAX1 \mult_97/U1236  ( .A(\mult_97/n2371 ), .B(\mult_97/n2278 ), .C(
        \mult_97/n2309 ), .YC(\mult_97/n1831 ), .YS(\mult_97/n1832 ) );
  FAX1 \mult_97/U1235  ( .A(\mult_97/n2340 ), .B(\mult_97/n2249 ), .C(
        \mult_97/n1837 ), .YC(\mult_97/n1829 ), .YS(\mult_97/n1830 ) );
  FAX1 \mult_97/U1234  ( .A(\mult_97/n1835 ), .B(\mult_97/n1832 ), .C(
        \mult_97/n1830 ), .YC(\mult_97/n1827 ), .YS(\mult_97/n1828 ) );
  HAX1 \mult_97/U1233  ( .A(\mult_97/n2370 ), .B(\mult_97/n2277 ), .YC(
        \mult_97/n1825 ), .YS(\mult_97/n1826 ) );
  FAX1 \mult_97/U1232  ( .A(\mult_97/n2308 ), .B(\mult_97/n2339 ), .C(
        \mult_97/n1862 ), .YC(\mult_97/n1823 ), .YS(\mult_97/n1824 ) );
  FAX1 \mult_97/U1231  ( .A(\mult_97/n2248 ), .B(\mult_97/n1826 ), .C(
        \mult_97/n1831 ), .YC(\mult_97/n1821 ), .YS(\mult_97/n1822 ) );
  FAX1 \mult_97/U1230  ( .A(\mult_97/n1824 ), .B(\mult_97/n1829 ), .C(
        \mult_97/n1822 ), .YC(\mult_97/n1819 ), .YS(\mult_97/n1820 ) );
  FAX1 \mult_97/U1229  ( .A(\mult_97/n2369 ), .B(\mult_97/n2216 ), .C(
        \mult_97/n2276 ), .YC(\mult_97/n1817 ), .YS(\mult_97/n1818 ) );
  FAX1 \mult_97/U1228  ( .A(\mult_97/n2307 ), .B(\mult_97/n2338 ), .C(
        \mult_97/n2247 ), .YC(\mult_97/n1815 ), .YS(\mult_97/n1816 ) );
  FAX1 \mult_97/U1227  ( .A(\mult_97/n1825 ), .B(\mult_97/n1823 ), .C(
        \mult_97/n1818 ), .YC(\mult_97/n1813 ), .YS(\mult_97/n1814 ) );
  FAX1 \mult_97/U1226  ( .A(\mult_97/n1816 ), .B(\mult_97/n1821 ), .C(
        \mult_97/n1814 ), .YC(\mult_97/n1811 ), .YS(\mult_97/n1812 ) );
  HAX1 \mult_97/U1225  ( .A(\mult_97/n2368 ), .B(\mult_97/n2275 ), .YC(
        \mult_97/n1809 ), .YS(\mult_97/n1810 ) );
  FAX1 \mult_97/U1224  ( .A(\mult_97/n1861 ), .B(\mult_97/n2215 ), .C(
        \mult_97/n2337 ), .YC(\mult_97/n1807 ), .YS(\mult_97/n1808 ) );
  FAX1 \mult_97/U1223  ( .A(\mult_97/n2306 ), .B(\mult_97/n2246 ), .C(
        \mult_97/n1810 ), .YC(\mult_97/n1805 ), .YS(\mult_97/n1806 ) );
  FAX1 \mult_97/U1222  ( .A(\mult_97/n1817 ), .B(\mult_97/n1815 ), .C(
        \mult_97/n1808 ), .YC(\mult_97/n1803 ), .YS(\mult_97/n1804 ) );
  FAX1 \mult_97/U1221  ( .A(\mult_97/n1806 ), .B(\mult_97/n1813 ), .C(
        \mult_97/n1804 ), .YC(\mult_97/n1801 ), .YS(\mult_97/n1802 ) );
  FAX1 \mult_97/U1220  ( .A(\mult_97/n2367 ), .B(\mult_97/n2274 ), .C(
        \mult_97/n2305 ), .YC(\mult_97/n1799 ), .YS(\mult_97/n1800 ) );
  FAX1 \mult_97/U1219  ( .A(\mult_97/n2214 ), .B(\mult_97/n2336 ), .C(
        \mult_97/n2245 ), .YC(\mult_97/n1797 ), .YS(\mult_97/n1798 ) );
  FAX1 \mult_97/U1218  ( .A(\mult_97/n2183 ), .B(\mult_97/n1809 ), .C(
        \mult_97/n1807 ), .YC(\mult_97/n1795 ), .YS(\mult_97/n1796 ) );
  FAX1 \mult_97/U1217  ( .A(\mult_97/n1800 ), .B(\mult_97/n1798 ), .C(
        \mult_97/n1805 ), .YC(\mult_97/n1793 ), .YS(\mult_97/n1794 ) );
  FAX1 \mult_97/U1216  ( .A(\mult_97/n1803 ), .B(\mult_97/n1796 ), .C(
        \mult_97/n1794 ), .YC(\mult_97/n1791 ), .YS(\mult_97/n1792 ) );
  HAX1 \mult_97/U1215  ( .A(\mult_97/n2366 ), .B(\mult_97/n1860 ), .YC(
        \mult_97/n1789 ), .YS(\mult_97/n1790 ) );
  FAX1 \mult_97/U1214  ( .A(\mult_97/n2273 ), .B(\mult_97/n2213 ), .C(
        \mult_97/n2335 ), .YC(\mult_97/n1787 ), .YS(\mult_97/n1788 ) );
  FAX1 \mult_97/U1213  ( .A(\mult_97/n2182 ), .B(\mult_97/n2304 ), .C(
        \mult_97/n2244 ), .YC(\mult_97/n1785 ), .YS(\mult_97/n1786 ) );
  FAX1 \mult_97/U1212  ( .A(\mult_97/n1790 ), .B(\mult_97/n1799 ), .C(
        \mult_97/n1797 ), .YC(\mult_97/n1783 ), .YS(\mult_97/n1784 ) );
  FAX1 \mult_97/U1211  ( .A(\mult_97/n1786 ), .B(\mult_97/n1788 ), .C(
        \mult_97/n1795 ), .YC(\mult_97/n1781 ), .YS(\mult_97/n1782 ) );
  FAX1 \mult_97/U1210  ( .A(\mult_97/n1784 ), .B(\mult_97/n1793 ), .C(
        \mult_97/n1782 ), .YC(\mult_97/n1779 ), .YS(\mult_97/n1780 ) );
  FAX1 \mult_97/U1209  ( .A(\mult_97/n2365 ), .B(\mult_97/n2272 ), .C(
        \mult_97/n2181 ), .YC(\mult_97/n1777 ), .YS(\mult_97/n1778 ) );
  FAX1 \mult_97/U1208  ( .A(\mult_97/n2303 ), .B(\mult_97/n2212 ), .C(
        \mult_97/n2243 ), .YC(\mult_97/n1775 ), .YS(\mult_97/n1776 ) );
  FAX1 \mult_97/U1207  ( .A(\mult_97/n2334 ), .B(\mult_97/n2152 ), .C(
        \mult_97/n1789 ), .YC(\mult_97/n1773 ), .YS(\mult_97/n1774 ) );
  FAX1 \mult_97/U1206  ( .A(\mult_97/n1787 ), .B(\mult_97/n1785 ), .C(
        \mult_97/n1778 ), .YC(\mult_97/n1771 ), .YS(\mult_97/n1772 ) );
  FAX1 \mult_97/U1205  ( .A(\mult_97/n1776 ), .B(\mult_97/n1774 ), .C(
        \mult_97/n1783 ), .YC(\mult_97/n1769 ), .YS(\mult_97/n1770 ) );
  FAX1 \mult_97/U1204  ( .A(\mult_97/n1772 ), .B(\mult_97/n1781 ), .C(
        \mult_97/n1770 ), .YC(\mult_97/n1767 ), .YS(\mult_97/n1768 ) );
  HAX1 \mult_97/U1203  ( .A(\mult_97/n2364 ), .B(\mult_97/n2271 ), .YC(
        \mult_97/n1765 ), .YS(\mult_97/n1766 ) );
  FAX1 \mult_97/U1202  ( .A(\mult_97/n2180 ), .B(\mult_97/n2302 ), .C(
        \mult_97/n1859 ), .YC(\mult_97/n1763 ), .YS(\mult_97/n1764 ) );
  FAX1 \mult_97/U1201  ( .A(\mult_97/n2211 ), .B(\mult_97/n2333 ), .C(
        \mult_97/n2151 ), .YC(\mult_97/n1761 ), .YS(\mult_97/n1762 ) );
  FAX1 \mult_97/U1200  ( .A(\mult_97/n2242 ), .B(\mult_97/n1766 ), .C(
        \mult_97/n1777 ), .YC(\mult_97/n1759 ), .YS(\mult_97/n1760 ) );
  FAX1 \mult_97/U1199  ( .A(\mult_97/n1775 ), .B(\mult_97/n1764 ), .C(
        \mult_97/n1762 ), .YC(\mult_97/n1757 ), .YS(\mult_97/n1758 ) );
  FAX1 \mult_97/U1198  ( .A(\mult_97/n1773 ), .B(\mult_97/n1771 ), .C(
        \mult_97/n1760 ), .YC(\mult_97/n1755 ), .YS(\mult_97/n1756 ) );
  FAX1 \mult_97/U1197  ( .A(\mult_97/n1758 ), .B(\mult_97/n1769 ), .C(
        \mult_97/n1756 ), .YC(\mult_97/n1753 ), .YS(\mult_97/n1754 ) );
  FAX1 \mult_97/U1196  ( .A(\mult_97/n2363 ), .B(\mult_97/n2119 ), .C(
        \mult_97/n2270 ), .YC(\mult_97/n1751 ), .YS(\mult_97/n1752 ) );
  FAX1 \mult_97/U1195  ( .A(\mult_97/n2179 ), .B(\mult_97/n2210 ), .C(
        \mult_97/n2150 ), .YC(\mult_97/n1749 ), .YS(\mult_97/n1750 ) );
  FAX1 \mult_97/U1194  ( .A(\mult_97/n2301 ), .B(\mult_97/n2332 ), .C(
        \mult_97/n2241 ), .YC(\mult_97/n1747 ), .YS(\mult_97/n1748 ) );
  FAX1 \mult_97/U1193  ( .A(\mult_97/n1765 ), .B(\mult_97/n1763 ), .C(
        \mult_97/n1761 ), .YC(\mult_97/n1745 ), .YS(\mult_97/n1746 ) );
  FAX1 \mult_97/U1192  ( .A(\mult_97/n1752 ), .B(\mult_97/n1750 ), .C(
        \mult_97/n1748 ), .YC(\mult_97/n1743 ), .YS(\mult_97/n1744 ) );
  FAX1 \mult_97/U1191  ( .A(\mult_97/n1759 ), .B(\mult_97/n1757 ), .C(
        \mult_97/n1746 ), .YC(\mult_97/n1741 ), .YS(\mult_97/n1742 ) );
  FAX1 \mult_97/U1190  ( .A(\mult_97/n1744 ), .B(\mult_97/n1755 ), .C(
        \mult_97/n1742 ), .YC(\mult_97/n1739 ), .YS(\mult_97/n1740 ) );
  HAX1 \mult_97/U1189  ( .A(\mult_97/n2362 ), .B(\mult_97/n2269 ), .YC(
        \mult_97/n1737 ), .YS(\mult_97/n1738 ) );
  FAX1 \mult_97/U1188  ( .A(\mult_97/n2178 ), .B(\mult_97/n1858 ), .C(
        \mult_97/n2331 ), .YC(\mult_97/n1735 ), .YS(\mult_97/n1736 ) );
  FAX1 \mult_97/U1187  ( .A(\mult_97/n2118 ), .B(\mult_97/n2209 ), .C(
        \mult_97/n2149 ), .YC(\mult_97/n1733 ), .YS(\mult_97/n1734 ) );
  FAX1 \mult_97/U1186  ( .A(\mult_97/n2300 ), .B(\mult_97/n2240 ), .C(
        \mult_97/n1738 ), .YC(\mult_97/n1731 ), .YS(\mult_97/n1732 ) );
  FAX1 \mult_97/U1185  ( .A(\mult_97/n1751 ), .B(\mult_97/n1749 ), .C(
        \mult_97/n1747 ), .YC(\mult_97/n1729 ), .YS(\mult_97/n1730 ) );
  FAX1 \mult_97/U1184  ( .A(\mult_97/n1736 ), .B(\mult_97/n1734 ), .C(
        \mult_97/n1732 ), .YC(\mult_97/n1727 ), .YS(\mult_97/n1728 ) );
  FAX1 \mult_97/U1183  ( .A(\mult_97/n1745 ), .B(\mult_97/n1743 ), .C(
        \mult_97/n1730 ), .YC(\mult_97/n1725 ), .YS(\mult_97/n1726 ) );
  FAX1 \mult_97/U1182  ( .A(\mult_97/n1728 ), .B(\mult_97/n1741 ), .C(
        \mult_97/n1726 ), .YC(\mult_97/n1723 ), .YS(\mult_97/n1724 ) );
  FAX1 \mult_97/U1181  ( .A(\mult_97/n2361 ), .B(\mult_97/n2268 ), .C(
        \mult_97/n2177 ), .YC(\mult_97/n1721 ), .YS(\mult_97/n1722 ) );
  FAX1 \mult_97/U1180  ( .A(\mult_97/n2208 ), .B(\mult_97/n2117 ), .C(
        \mult_97/n2148 ), .YC(\mult_97/n1719 ), .YS(\mult_97/n1720 ) );
  FAX1 \mult_97/U1179  ( .A(\mult_97/n2299 ), .B(\mult_97/n2330 ), .C(
        \mult_97/n2239 ), .YC(\mult_97/n1717 ), .YS(\mult_97/n1718 ) );
  FAX1 \mult_97/U1178  ( .A(\mult_97/n2086 ), .B(\mult_97/n1737 ), .C(
        \mult_97/n1735 ), .YC(\mult_97/n1715 ), .YS(\mult_97/n1716 ) );
  FAX1 \mult_97/U1177  ( .A(\mult_97/n1733 ), .B(\mult_97/n1722 ), .C(
        \mult_97/n1720 ), .YC(\mult_97/n1713 ), .YS(\mult_97/n1714 ) );
  FAX1 \mult_97/U1176  ( .A(\mult_97/n1718 ), .B(\mult_97/n1731 ), .C(
        \mult_97/n1729 ), .YC(\mult_97/n1711 ), .YS(\mult_97/n1712 ) );
  FAX1 \mult_97/U1175  ( .A(\mult_97/n1716 ), .B(\mult_97/n1714 ), .C(
        \mult_97/n1727 ), .YC(\mult_97/n1709 ), .YS(\mult_97/n1710 ) );
  FAX1 \mult_97/U1174  ( .A(\mult_97/n1712 ), .B(\mult_97/n1725 ), .C(
        \mult_97/n1710 ), .YC(\mult_97/n1707 ), .YS(\mult_97/n1708 ) );
  HAX1 \mult_97/U1173  ( .A(\mult_97/n2360 ), .B(\mult_97/n1857 ), .YC(
        \mult_97/n1705 ), .YS(\mult_97/n1706 ) );
  FAX1 \mult_97/U1172  ( .A(\mult_97/n2085 ), .B(\mult_97/n2298 ), .C(
        \mult_97/n2238 ), .YC(\mult_97/n1703 ), .YS(\mult_97/n1704 ) );
  FAX1 \mult_97/U1171  ( .A(\mult_97/n2267 ), .B(\mult_97/n2116 ), .C(
        \mult_97/n2147 ), .YC(\mult_97/n1701 ), .YS(\mult_97/n1702 ) );
  FAX1 \mult_97/U1170  ( .A(\mult_97/n2176 ), .B(\mult_97/n2207 ), .C(
        \mult_97/n2329 ), .YC(\mult_97/n1699 ), .YS(\mult_97/n1700 ) );
  FAX1 \mult_97/U1169  ( .A(\mult_97/n1706 ), .B(\mult_97/n1721 ), .C(
        \mult_97/n1719 ), .YC(\mult_97/n1697 ), .YS(\mult_97/n1698 ) );
  FAX1 \mult_97/U1168  ( .A(\mult_97/n1717 ), .B(\mult_97/n1700 ), .C(
        \mult_97/n1702 ), .YC(\mult_97/n1695 ), .YS(\mult_97/n1696 ) );
  FAX1 \mult_97/U1167  ( .A(\mult_97/n1704 ), .B(\mult_97/n1715 ), .C(
        \mult_97/n1713 ), .YC(\mult_97/n1693 ), .YS(\mult_97/n1694 ) );
  FAX1 \mult_97/U1166  ( .A(\mult_97/n1698 ), .B(\mult_97/n1696 ), .C(
        \mult_97/n1711 ), .YC(\mult_97/n1691 ), .YS(\mult_97/n1692 ) );
  FAX1 \mult_97/U1165  ( .A(\mult_97/n1694 ), .B(\mult_97/n1709 ), .C(
        \mult_97/n1692 ), .YC(\mult_97/n1689 ), .YS(\mult_97/n1690 ) );
  FAX1 \mult_97/U1164  ( .A(\mult_97/n2359 ), .B(\mult_97/n2084 ), .C(
        \mult_97/n2175 ), .YC(\mult_97/n1687 ), .YS(\mult_97/n1688 ) );
  FAX1 \mult_97/U1163  ( .A(\mult_97/n2266 ), .B(\mult_97/n2115 ), .C(
        \mult_97/n2146 ), .YC(\mult_97/n1685 ), .YS(\mult_97/n1686 ) );
  FAX1 \mult_97/U1162  ( .A(\mult_97/n2206 ), .B(\mult_97/n2297 ), .C(
        \mult_97/n2237 ), .YC(\mult_97/n1683 ), .YS(\mult_97/n1684 ) );
  FAX1 \mult_97/U1161  ( .A(\mult_97/n2328 ), .B(\mult_97/n2055 ), .C(
        \mult_97/n1705 ), .YC(\mult_97/n1681 ), .YS(\mult_97/n1682 ) );
  FAX1 \mult_97/U1160  ( .A(\mult_97/n1703 ), .B(\mult_97/n1699 ), .C(
        \mult_97/n1701 ), .YC(\mult_97/n1679 ), .YS(\mult_97/n1680 ) );
  FAX1 \mult_97/U1159  ( .A(\mult_97/n1688 ), .B(\mult_97/n1686 ), .C(
        \mult_97/n1684 ), .YC(\mult_97/n1677 ), .YS(\mult_97/n1678 ) );
  FAX1 \mult_97/U1158  ( .A(\mult_97/n1682 ), .B(\mult_97/n1697 ), .C(
        \mult_97/n1695 ), .YC(\mult_97/n1675 ), .YS(\mult_97/n1676 ) );
  FAX1 \mult_97/U1157  ( .A(\mult_97/n1680 ), .B(\mult_97/n1678 ), .C(
        \mult_97/n1693 ), .YC(\mult_97/n1673 ), .YS(\mult_97/n1674 ) );
  FAX1 \mult_97/U1156  ( .A(\mult_97/n1676 ), .B(\mult_97/n1691 ), .C(
        \mult_97/n1674 ), .YC(n242), .YS(n241) );
  HAX1 \mult_97/U1155  ( .A(\mult_97/n2358 ), .B(\mult_97/n2083 ), .YC(
        \mult_97/n1669 ), .YS(\mult_97/n1670 ) );
  FAX1 \mult_97/U1154  ( .A(\mult_97/n2174 ), .B(\mult_97/n2114 ), .C(
        \mult_97/n2327 ), .YC(\mult_97/n1667 ), .YS(\mult_97/n1668 ) );
  FAX1 \mult_97/U1153  ( .A(\mult_97/n2265 ), .B(\mult_97/n2205 ), .C(
        \mult_97/n1856 ), .YC(\mult_97/n1665 ), .YS(\mult_97/n1666 ) );
  FAX1 \mult_97/U1152  ( .A(\mult_97/n2296 ), .B(\mult_97/n2236 ), .C(
        \mult_97/n2054 ), .YC(\mult_97/n1663 ), .YS(\mult_97/n1664 ) );
  FAX1 \mult_97/U1151  ( .A(\mult_97/n2145 ), .B(\mult_97/n1670 ), .C(
        \mult_97/n1687 ), .YC(\mult_97/n1661 ), .YS(\mult_97/n1662 ) );
  FAX1 \mult_97/U1150  ( .A(\mult_97/n1685 ), .B(\mult_97/n1683 ), .C(
        \mult_97/n1666 ), .YC(\mult_97/n1659 ), .YS(\mult_97/n1660 ) );
  FAX1 \mult_97/U1149  ( .A(\mult_97/n1668 ), .B(\mult_97/n1664 ), .C(
        \mult_97/n1681 ), .YC(\mult_97/n1657 ), .YS(\mult_97/n1658 ) );
  FAX1 \mult_97/U1148  ( .A(\mult_97/n1679 ), .B(\mult_97/n1662 ), .C(
        \mult_97/n1677 ), .YC(\mult_97/n1655 ), .YS(\mult_97/n1656 ) );
  FAX1 \mult_97/U1147  ( .A(\mult_97/n1660 ), .B(\mult_97/n1658 ), .C(
        \mult_97/n1675 ), .YC(\mult_97/n1653 ), .YS(\mult_97/n1654 ) );
  FAX1 \mult_97/U1146  ( .A(\mult_97/n1656 ), .B(\mult_97/n1673 ), .C(
        \mult_97/n1654 ), .YC(n240), .YS(n239) );
  FAX1 \mult_97/U1145  ( .A(\mult_97/n2357 ), .B(\mult_97/n2022 ), .C(
        \mult_97/n2082 ), .YC(\mult_97/n1649 ), .YS(\mult_97/n1650 ) );
  FAX1 \mult_97/U1144  ( .A(\mult_97/n2173 ), .B(\mult_97/n2113 ), .C(
        \mult_97/n2053 ), .YC(\mult_97/n1647 ), .YS(\mult_97/n1648 ) );
  FAX1 \mult_97/U1143  ( .A(\mult_97/n2264 ), .B(\mult_97/n2295 ), .C(
        \mult_97/n2144 ), .YC(\mult_97/n1645 ), .YS(\mult_97/n1646 ) );
  FAX1 \mult_97/U1142  ( .A(\mult_97/n2204 ), .B(\mult_97/n2326 ), .C(
        \mult_97/n2235 ), .YC(\mult_97/n1643 ), .YS(\mult_97/n1644 ) );
  FAX1 \mult_97/U1141  ( .A(\mult_97/n1669 ), .B(\mult_97/n1667 ), .C(
        \mult_97/n1665 ), .YC(\mult_97/n1641 ), .YS(\mult_97/n1642 ) );
  FAX1 \mult_97/U1140  ( .A(\mult_97/n1663 ), .B(\mult_97/n1650 ), .C(
        \mult_97/n1646 ), .YC(\mult_97/n1639 ), .YS(\mult_97/n1640 ) );
  FAX1 \mult_97/U1139  ( .A(\mult_97/n1648 ), .B(\mult_97/n1644 ), .C(
        \mult_97/n1661 ), .YC(\mult_97/n1637 ), .YS(\mult_97/n1638 ) );
  FAX1 \mult_97/U1138  ( .A(\mult_97/n1659 ), .B(\mult_97/n1642 ), .C(
        \mult_97/n1657 ), .YC(\mult_97/n1635 ), .YS(\mult_97/n1636 ) );
  FAX1 \mult_97/U1137  ( .A(\mult_97/n1640 ), .B(\mult_97/n1638 ), .C(
        \mult_97/n1655 ), .YC(\mult_97/n1633 ), .YS(\mult_97/n1634 ) );
  FAX1 \mult_97/U1136  ( .A(\mult_97/n1636 ), .B(\mult_97/n1653 ), .C(
        \mult_97/n1634 ), .YC(n238), .YS(n237) );
  HAX1 \mult_97/U1135  ( .A(\mult_97/n2356 ), .B(\mult_97/n2081 ), .YC(
        \mult_97/n1629 ), .YS(\mult_97/n1630 ) );
  FAX1 \mult_97/U1134  ( .A(\mult_97/n2172 ), .B(\mult_97/n1855 ), .C(
        \mult_97/n2234 ), .YC(\mult_97/n1627 ), .YS(\mult_97/n1628 ) );
  FAX1 \mult_97/U1133  ( .A(\mult_97/n2263 ), .B(\mult_97/n2021 ), .C(
        \mult_97/n2325 ), .YC(\mult_97/n1625 ), .YS(\mult_97/n1626 ) );
  FAX1 \mult_97/U1132  ( .A(\mult_97/n2294 ), .B(\mult_97/n2112 ), .C(
        \mult_97/n2052 ), .YC(\mult_97/n1623 ), .YS(\mult_97/n1624 ) );
  FAX1 \mult_97/U1131  ( .A(\mult_97/n2203 ), .B(\mult_97/n2143 ), .C(
        \mult_97/n1630 ), .YC(\mult_97/n1621 ), .YS(\mult_97/n1622 ) );
  FAX1 \mult_97/U1130  ( .A(\mult_97/n1649 ), .B(\mult_97/n1647 ), .C(
        \mult_97/n1645 ), .YC(\mult_97/n1619 ), .YS(\mult_97/n1620 ) );
  FAX1 \mult_97/U1129  ( .A(\mult_97/n1643 ), .B(\mult_97/n1628 ), .C(
        \mult_97/n1626 ), .YC(\mult_97/n1617 ), .YS(\mult_97/n1618 ) );
  FAX1 \mult_97/U1128  ( .A(\mult_97/n1624 ), .B(\mult_97/n1622 ), .C(
        \mult_97/n1641 ), .YC(\mult_97/n1615 ), .YS(\mult_97/n1616 ) );
  FAX1 \mult_97/U1127  ( .A(\mult_97/n1639 ), .B(\mult_97/n1620 ), .C(
        \mult_97/n1618 ), .YC(\mult_97/n1613 ), .YS(\mult_97/n1614 ) );
  FAX1 \mult_97/U1126  ( .A(\mult_97/n1637 ), .B(\mult_97/n1616 ), .C(
        \mult_97/n1635 ), .YC(\mult_97/n1611 ), .YS(\mult_97/n1612 ) );
  FAX1 \mult_97/U1125  ( .A(n441), .B(n442), .C(n440), .YC(\mult_97/n1609 ), 
        .YS(\mult_97/n1610 ) );
  FAX1 \mult_97/U1124  ( .A(\mult_97/n2355 ), .B(\mult_97/n2171 ), .C(
        \mult_97/n2262 ), .YC(\mult_97/n1607 ), .YS(\mult_97/n1608 ) );
  FAX1 \mult_97/U1123  ( .A(\mult_97/n2080 ), .B(\mult_97/n2020 ), .C(
        \mult_97/n2051 ), .YC(\mult_97/n1605 ), .YS(\mult_97/n1606 ) );
  FAX1 \mult_97/U1122  ( .A(\mult_97/n2293 ), .B(\mult_97/n2202 ), .C(
        \mult_97/n2233 ), .YC(\mult_97/n1603 ), .YS(\mult_97/n1604 ) );
  FAX1 \mult_97/U1121  ( .A(\mult_97/n2111 ), .B(\mult_97/n2324 ), .C(
        \mult_97/n2142 ), .YC(\mult_97/n1601 ), .YS(\mult_97/n1602 ) );
  FAX1 \mult_97/U1120  ( .A(\mult_97/n1989 ), .B(\mult_97/n1629 ), .C(
        \mult_97/n1627 ), .YC(\mult_97/n1599 ), .YS(\mult_97/n1600 ) );
  FAX1 \mult_97/U1119  ( .A(\mult_97/n1625 ), .B(\mult_97/n1623 ), .C(
        \mult_97/n1608 ), .YC(\mult_97/n1597 ), .YS(\mult_97/n1598 ) );
  FAX1 \mult_97/U1118  ( .A(\mult_97/n1606 ), .B(\mult_97/n1604 ), .C(
        \mult_97/n1602 ), .YC(\mult_97/n1595 ), .YS(\mult_97/n1596 ) );
  FAX1 \mult_97/U1117  ( .A(\mult_97/n1621 ), .B(\mult_97/n1619 ), .C(
        \mult_97/n1600 ), .YC(\mult_97/n1593 ), .YS(\mult_97/n1594 ) );
  FAX1 \mult_97/U1116  ( .A(\mult_97/n1617 ), .B(\mult_97/n1598 ), .C(
        \mult_97/n1596 ), .YC(\mult_97/n1591 ), .YS(\mult_97/n1592 ) );
  FAX1 \mult_97/U1115  ( .A(\mult_97/n1615 ), .B(\mult_97/n1594 ), .C(
        \mult_97/n1613 ), .YC(\mult_97/n1589 ), .YS(\mult_97/n1590 ) );
  FAX1 \mult_97/U1114  ( .A(n438), .B(n439), .C(n437), .YC(\mult_97/n1587 ), 
        .YS(\mult_97/n1588 ) );
  HAX1 \mult_97/U1113  ( .A(\mult_97/n2354 ), .B(\mult_97/n1854 ), .YC(
        \mult_97/n1585 ), .YS(\mult_97/n1586 ) );
  FAX1 \mult_97/U1112  ( .A(\mult_97/n2170 ), .B(\mult_97/n2110 ), .C(
        \mult_97/n2323 ), .YC(\mult_97/n1583 ), .YS(\mult_97/n1584 ) );
  FAX1 \mult_97/U1111  ( .A(\mult_97/n2079 ), .B(\mult_97/n2019 ), .C(
        \mult_97/n2141 ), .YC(\mult_97/n1581 ), .YS(\mult_97/n1582 ) );
  FAX1 \mult_97/U1110  ( .A(\mult_97/n1988 ), .B(\mult_97/n2201 ), .C(
        \mult_97/n2050 ), .YC(\mult_97/n1579 ), .YS(\mult_97/n1580 ) );
  FAX1 \mult_97/U1109  ( .A(\mult_97/n2261 ), .B(\mult_97/n2292 ), .C(
        \mult_97/n2232 ), .YC(\mult_97/n1577 ), .YS(\mult_97/n1578 ) );
  FAX1 \mult_97/U1108  ( .A(\mult_97/n1586 ), .B(\mult_97/n1607 ), .C(
        \mult_97/n1605 ), .YC(\mult_97/n1575 ), .YS(\mult_97/n1576 ) );
  FAX1 \mult_97/U1107  ( .A(\mult_97/n1603 ), .B(\mult_97/n1601 ), .C(
        \mult_97/n1578 ), .YC(\mult_97/n1573 ), .YS(\mult_97/n1574 ) );
  FAX1 \mult_97/U1106  ( .A(\mult_97/n1580 ), .B(\mult_97/n1584 ), .C(
        \mult_97/n1582 ), .YC(\mult_97/n1571 ), .YS(\mult_97/n1572 ) );
  FAX1 \mult_97/U1105  ( .A(\mult_97/n1599 ), .B(\mult_97/n1597 ), .C(
        \mult_97/n1576 ), .YC(\mult_97/n1569 ), .YS(\mult_97/n1570 ) );
  FAX1 \mult_97/U1104  ( .A(\mult_97/n1595 ), .B(\mult_97/n1574 ), .C(
        \mult_97/n1572 ), .YC(\mult_97/n1567 ), .YS(\mult_97/n1568 ) );
  FAX1 \mult_97/U1103  ( .A(\mult_97/n1593 ), .B(\mult_97/n1591 ), .C(
        \mult_97/n1570 ), .YC(\mult_97/n1565 ), .YS(\mult_97/n1566 ) );
  FAX1 \mult_97/U1102  ( .A(n435), .B(n436), .C(n434), .YC(\mult_97/n1563 ), 
        .YS(\mult_97/n1564 ) );
  FAX1 \mult_97/U1101  ( .A(\mult_97/n2353 ), .B(\mult_97/n2169 ), .C(
        \mult_97/n1987 ), .YC(\mult_97/n1561 ), .YS(\mult_97/n1562 ) );
  FAX1 \mult_97/U1100  ( .A(\mult_97/n2260 ), .B(\mult_97/n2018 ), .C(
        \mult_97/n2049 ), .YC(\mult_97/n1559 ), .YS(\mult_97/n1560 ) );
  FAX1 \mult_97/U1099  ( .A(\mult_97/n2078 ), .B(\mult_97/n2109 ), .C(
        \mult_97/n2140 ), .YC(\mult_97/n1557 ), .YS(\mult_97/n1558 ) );
  FAX1 \mult_97/U1098  ( .A(\mult_97/n2291 ), .B(\mult_97/n2200 ), .C(
        \mult_97/n2231 ), .YC(\mult_97/n1555 ), .YS(\mult_97/n1556 ) );
  FAX1 \mult_97/U1097  ( .A(\mult_97/n2322 ), .B(\mult_97/n1962 ), .C(
        \mult_97/n1585 ), .YC(\mult_97/n1553 ), .YS(\mult_97/n1554 ) );
  FAX1 \mult_97/U1096  ( .A(\mult_97/n1583 ), .B(\mult_97/n1577 ), .C(
        \mult_97/n1579 ), .YC(\mult_97/n1551 ), .YS(\mult_97/n1552 ) );
  FAX1 \mult_97/U1095  ( .A(\mult_97/n1581 ), .B(\mult_97/n1562 ), .C(
        \mult_97/n1560 ), .YC(\mult_97/n1549 ), .YS(\mult_97/n1550 ) );
  FAX1 \mult_97/U1094  ( .A(\mult_97/n1558 ), .B(\mult_97/n1556 ), .C(
        \mult_97/n1554 ), .YC(\mult_97/n1547 ), .YS(\mult_97/n1548 ) );
  FAX1 \mult_97/U1093  ( .A(\mult_97/n1575 ), .B(\mult_97/n1573 ), .C(
        \mult_97/n1571 ), .YC(\mult_97/n1545 ), .YS(\mult_97/n1546 ) );
  FAX1 \mult_97/U1092  ( .A(\mult_97/n1552 ), .B(\mult_97/n1550 ), .C(
        \mult_97/n1548 ), .YC(\mult_97/n1543 ), .YS(\mult_97/n1544 ) );
  FAX1 \mult_97/U1091  ( .A(\mult_97/n1569 ), .B(\mult_97/n1567 ), .C(
        \mult_97/n1546 ), .YC(\mult_97/n1541 ), .YS(\mult_97/n1542 ) );
  FAX1 \mult_97/U1090  ( .A(n432), .B(n433), .C(n431), .YC(\mult_97/n1539 ), 
        .YS(\mult_97/n1540 ) );
  HAX1 \mult_97/U1089  ( .A(\mult_97/n2352 ), .B(\mult_97/n2077 ), .YC(
        \mult_97/n1537 ), .YS(\mult_97/n1538 ) );
  FAX1 \mult_97/U1088  ( .A(\mult_97/n2259 ), .B(\mult_97/n2199 ), .C(
        \mult_97/n2321 ), .YC(\mult_97/n1535 ), .YS(\mult_97/n1536 ) );
  FAX1 \mult_97/U1087  ( .A(\mult_97/n2168 ), .B(\mult_97/n2108 ), .C(
        \mult_97/n1961 ), .YC(\mult_97/n1533 ), .YS(\mult_97/n1534 ) );
  FAX1 \mult_97/U1086  ( .A(\mult_97/n1986 ), .B(\mult_97/n2017 ), .C(
        \mult_97/n1853 ), .YC(\mult_97/n1531 ), .YS(\mult_97/n1532 ) );
  FAX1 \mult_97/U1085  ( .A(\mult_97/n2290 ), .B(\mult_97/n2230 ), .C(
        \mult_97/n2048 ), .YC(\mult_97/n1529 ), .YS(\mult_97/n1530 ) );
  FAX1 \mult_97/U1084  ( .A(\mult_97/n2139 ), .B(\mult_97/n1538 ), .C(
        \mult_97/n1561 ), .YC(\mult_97/n1527 ), .YS(\mult_97/n1528 ) );
  FAX1 \mult_97/U1083  ( .A(\mult_97/n1557 ), .B(\mult_97/n1559 ), .C(
        \mult_97/n1555 ), .YC(\mult_97/n1525 ), .YS(\mult_97/n1526 ) );
  FAX1 \mult_97/U1082  ( .A(\mult_97/n1534 ), .B(\mult_97/n1532 ), .C(
        \mult_97/n1530 ), .YC(\mult_97/n1523 ), .YS(\mult_97/n1524 ) );
  FAX1 \mult_97/U1081  ( .A(\mult_97/n1536 ), .B(\mult_97/n1553 ), .C(
        \mult_97/n1551 ), .YC(\mult_97/n1521 ), .YS(\mult_97/n1522 ) );
  FAX1 \mult_97/U1080  ( .A(\mult_97/n1528 ), .B(\mult_97/n1549 ), .C(
        \mult_97/n1526 ), .YC(\mult_97/n1519 ), .YS(\mult_97/n1520 ) );
  FAX1 \mult_97/U1079  ( .A(\mult_97/n1524 ), .B(\mult_97/n1547 ), .C(
        \mult_97/n1545 ), .YC(\mult_97/n1517 ), .YS(\mult_97/n1518 ) );
  FAX1 \mult_97/U1078  ( .A(\mult_97/n1522 ), .B(\mult_97/n1520 ), .C(
        \mult_97/n1543 ), .YC(\mult_97/n1515 ), .YS(\mult_97/n1516 ) );
  FAX1 \mult_97/U1077  ( .A(n429), .B(n430), .C(n428), .YC(\mult_97/n1513 ), 
        .YS(\mult_97/n1514 ) );
  FAX1 \mult_97/U1076  ( .A(\mult_97/n2351 ), .B(\mult_97/n1929 ), .C(
        \mult_97/n2167 ), .YC(\mult_97/n1511 ), .YS(\mult_97/n1512 ) );
  FAX1 \mult_97/U1075  ( .A(\mult_97/n2258 ), .B(\mult_97/n2016 ), .C(
        \mult_97/n1960 ), .YC(\mult_97/n1509 ), .YS(\mult_97/n1510 ) );
  FAX1 \mult_97/U1074  ( .A(\mult_97/n2076 ), .B(\mult_97/n2198 ), .C(
        \mult_97/n2229 ), .YC(\mult_97/n1507 ), .YS(\mult_97/n1508 ) );
  FAX1 \mult_97/U1073  ( .A(\mult_97/n1985 ), .B(\mult_97/n2107 ), .C(
        \mult_97/n2047 ), .YC(\mult_97/n1505 ), .YS(\mult_97/n1506 ) );
  FAX1 \mult_97/U1072  ( .A(\mult_97/n2289 ), .B(\mult_97/n2320 ), .C(
        \mult_97/n2138 ), .YC(\mult_97/n1503 ), .YS(\mult_97/n1504 ) );
  FAX1 \mult_97/U1071  ( .A(\mult_97/n1537 ), .B(\mult_97/n1535 ), .C(
        \mult_97/n1533 ), .YC(\mult_97/n1501 ), .YS(\mult_97/n1502 ) );
  FAX1 \mult_97/U1070  ( .A(\mult_97/n1531 ), .B(\mult_97/n1529 ), .C(
        \mult_97/n1512 ), .YC(\mult_97/n1499 ), .YS(\mult_97/n1500 ) );
  FAX1 \mult_97/U1069  ( .A(\mult_97/n1508 ), .B(\mult_97/n1506 ), .C(
        \mult_97/n1504 ), .YC(\mult_97/n1497 ), .YS(\mult_97/n1498 ) );
  FAX1 \mult_97/U1068  ( .A(\mult_97/n1510 ), .B(\mult_97/n1527 ), .C(
        \mult_97/n1525 ), .YC(\mult_97/n1495 ), .YS(\mult_97/n1496 ) );
  FAX1 \mult_97/U1067  ( .A(\mult_97/n1502 ), .B(\mult_97/n1523 ), .C(
        \mult_97/n1500 ), .YC(\mult_97/n1493 ), .YS(\mult_97/n1494 ) );
  FAX1 \mult_97/U1066  ( .A(\mult_97/n1498 ), .B(\mult_97/n1521 ), .C(
        \mult_97/n1496 ), .YC(\mult_97/n1491 ), .YS(\mult_97/n1492 ) );
  FAX1 \mult_97/U1065  ( .A(\mult_97/n1519 ), .B(\mult_97/n1494 ), .C(
        \mult_97/n1517 ), .YC(\mult_97/n1489 ), .YS(\mult_97/n1490 ) );
  FAX1 \mult_97/U1064  ( .A(n426), .B(n427), .C(n425), .YC(\mult_97/n1487 ), 
        .YS(\mult_97/n1488 ) );
  HAX1 \mult_97/U1063  ( .A(\mult_97/n2350 ), .B(\mult_97/n2166 ), .YC(
        \mult_97/n1485 ), .YS(\mult_97/n1486 ) );
  FAX1 \mult_97/U1062  ( .A(\mult_97/n2257 ), .B(\mult_97/n1928 ), .C(
        \mult_97/n2319 ), .YC(\mult_97/n1483 ), .YS(\mult_97/n1484 ) );
  FAX1 \mult_97/U1061  ( .A(\mult_97/n1984 ), .B(\mult_97/n2288 ), .C(
        \mult_97/n2137 ), .YC(\mult_97/n1481 ), .YS(\mult_97/n1482 ) );
  FAX1 \mult_97/U1060  ( .A(\mult_97/n2075 ), .B(\mult_97/n1852 ), .C(
        \mult_97/n1959 ), .YC(\mult_97/n1479 ), .YS(\mult_97/n1480 ) );
  FAX1 \mult_97/U1059  ( .A(\mult_97/n2106 ), .B(\mult_97/n2015 ), .C(
        \mult_97/n2046 ), .YC(\mult_97/n1477 ), .YS(\mult_97/n1478 ) );
  FAX1 \mult_97/U1058  ( .A(\mult_97/n2197 ), .B(\mult_97/n2228 ), .C(
        \mult_97/n1486 ), .YC(\mult_97/n1475 ), .YS(\mult_97/n1476 ) );
  FAX1 \mult_97/U1057  ( .A(\mult_97/n1511 ), .B(\mult_97/n1505 ), .C(
        \mult_97/n1507 ), .YC(\mult_97/n1473 ), .YS(\mult_97/n1474 ) );
  FAX1 \mult_97/U1056  ( .A(\mult_97/n1509 ), .B(\mult_97/n1503 ), .C(
        \mult_97/n1482 ), .YC(\mult_97/n1471 ), .YS(\mult_97/n1472 ) );
  FAX1 \mult_97/U1055  ( .A(\mult_97/n1480 ), .B(\mult_97/n1484 ), .C(
        \mult_97/n1478 ), .YC(\mult_97/n1469 ), .YS(\mult_97/n1470 ) );
  FAX1 \mult_97/U1054  ( .A(\mult_97/n1476 ), .B(\mult_97/n1501 ), .C(
        \mult_97/n1499 ), .YC(\mult_97/n1467 ), .YS(\mult_97/n1468 ) );
  FAX1 \mult_97/U1053  ( .A(\mult_97/n1474 ), .B(\mult_97/n1497 ), .C(
        \mult_97/n1472 ), .YC(\mult_97/n1465 ), .YS(\mult_97/n1466 ) );
  FAX1 \mult_97/U1052  ( .A(\mult_97/n1470 ), .B(\mult_97/n1495 ), .C(
        \mult_97/n1468 ), .YC(\mult_97/n1463 ), .YS(\mult_97/n1464 ) );
  FAX1 \mult_97/U1051  ( .A(\mult_97/n1493 ), .B(\mult_97/n1466 ), .C(
        \mult_97/n1491 ), .YC(\mult_97/n1461 ), .YS(\mult_97/n1462 ) );
  FAX1 \mult_97/U1050  ( .A(n423), .B(n424), .C(n422), .YC(\mult_97/n1459 ), 
        .YS(\mult_97/n1460 ) );
  FAX1 \mult_97/U1049  ( .A(\mult_97/n2349 ), .B(\mult_97/n2256 ), .C(
        \mult_97/n2165 ), .YC(\mult_97/n1457 ), .YS(\mult_97/n1458 ) );
  FAX1 \mult_97/U1048  ( .A(\mult_97/n2074 ), .B(\mult_97/n2014 ), .C(
        \mult_97/n2136 ), .YC(\mult_97/n1455 ), .YS(\mult_97/n1456 ) );
  FAX1 \mult_97/U1047  ( .A(\mult_97/n1983 ), .B(\mult_97/n2196 ), .C(
        \mult_97/n2045 ), .YC(\mult_97/n1453 ), .YS(\mult_97/n1454 ) );
  FAX1 \mult_97/U1046  ( .A(\mult_97/n2287 ), .B(\mult_97/n1927 ), .C(
        \mult_97/n1958 ), .YC(\mult_97/n1451 ), .YS(\mult_97/n1452 ) );
  FAX1 \mult_97/U1045  ( .A(\mult_97/n2105 ), .B(\mult_97/n2318 ), .C(
        \mult_97/n2227 ), .YC(\mult_97/n1449 ), .YS(\mult_97/n1450 ) );
  FAX1 \mult_97/U1044  ( .A(\mult_97/n1898 ), .B(\mult_97/n1485 ), .C(
        \mult_97/n1483 ), .YC(\mult_97/n1447 ), .YS(\mult_97/n1448 ) );
  FAX1 \mult_97/U1043  ( .A(\mult_97/n1481 ), .B(\mult_97/n1479 ), .C(
        \mult_97/n1477 ), .YC(\mult_97/n1445 ), .YS(\mult_97/n1446 ) );
  FAX1 \mult_97/U1042  ( .A(\mult_97/n1458 ), .B(\mult_97/n1456 ), .C(
        \mult_97/n1450 ), .YC(\mult_97/n1443 ), .YS(\mult_97/n1444 ) );
  FAX1 \mult_97/U1041  ( .A(\mult_97/n1454 ), .B(\mult_97/n1452 ), .C(
        \mult_97/n1475 ), .YC(\mult_97/n1441 ), .YS(\mult_97/n1442 ) );
  FAX1 \mult_97/U1040  ( .A(\mult_97/n1473 ), .B(\mult_97/n1471 ), .C(
        \mult_97/n1448 ), .YC(\mult_97/n1439 ), .YS(\mult_97/n1440 ) );
  FAX1 \mult_97/U1039  ( .A(\mult_97/n1469 ), .B(\mult_97/n1446 ), .C(
        \mult_97/n1444 ), .YC(\mult_97/n1437 ), .YS(\mult_97/n1438 ) );
  FAX1 \mult_97/U1038  ( .A(\mult_97/n1442 ), .B(\mult_97/n1467 ), .C(
        \mult_97/n1465 ), .YC(\mult_97/n1435 ), .YS(\mult_97/n1436 ) );
  FAX1 \mult_97/U1037  ( .A(\mult_97/n1440 ), .B(\mult_97/n1438 ), .C(
        \mult_97/n1463 ), .YC(\mult_97/n1433 ), .YS(\mult_97/n1434 ) );
  FAX1 \mult_97/U1036  ( .A(n420), .B(n421), .C(n419), .YC(\mult_97/n1431 ), 
        .YS(\mult_97/n1432 ) );
  HAX1 \mult_97/U1035  ( .A(\mult_97/n2348 ), .B(\mult_97/n2164 ), .YC(
        \mult_97/n1429 ), .YS(\mult_97/n1430 ) );
  FAX1 \mult_97/U1034  ( .A(\mult_97/n2073 ), .B(\mult_97/n2013 ), .C(
        \mult_97/n2317 ), .YC(\mult_97/n1427 ), .YS(\mult_97/n1428 ) );
  FAX1 \mult_97/U1033  ( .A(\mult_97/n2255 ), .B(\mult_97/n2286 ), .C(
        \mult_97/n2226 ), .YC(\mult_97/n1425 ), .YS(\mult_97/n1426 ) );
  FAX1 \mult_97/U1032  ( .A(\mult_97/n1982 ), .B(\mult_97/n2104 ), .C(
        \mult_97/n2044 ), .YC(\mult_97/n1423 ), .YS(\mult_97/n1424 ) );
  FAX1 \mult_97/U1031  ( .A(\mult_97/n2195 ), .B(\mult_97/n1926 ), .C(
        \mult_97/n1957 ), .YC(\mult_97/n1421 ), .YS(\mult_97/n1422 ) );
  FAX1 \mult_97/U1030  ( .A(\mult_97/n1897 ), .B(\mult_97/n1851 ), .C(
        \mult_97/n2135 ), .YC(\mult_97/n1419 ), .YS(\mult_97/n1420 ) );
  FAX1 \mult_97/U1029  ( .A(\mult_97/n1430 ), .B(\mult_97/n1457 ), .C(
        \mult_97/n1455 ), .YC(\mult_97/n1417 ), .YS(\mult_97/n1418 ) );
  FAX1 \mult_97/U1028  ( .A(\mult_97/n1453 ), .B(\mult_97/n1451 ), .C(
        \mult_97/n1449 ), .YC(\mult_97/n1415 ), .YS(\mult_97/n1416 ) );
  FAX1 \mult_97/U1027  ( .A(\mult_97/n1426 ), .B(\mult_97/n1422 ), .C(
        \mult_97/n1420 ), .YC(\mult_97/n1413 ), .YS(\mult_97/n1414 ) );
  FAX1 \mult_97/U1026  ( .A(\mult_97/n1424 ), .B(\mult_97/n1428 ), .C(
        \mult_97/n1447 ), .YC(\mult_97/n1411 ), .YS(\mult_97/n1412 ) );
  FAX1 \mult_97/U1025  ( .A(\mult_97/n1445 ), .B(\mult_97/n1418 ), .C(
        \mult_97/n1443 ), .YC(\mult_97/n1409 ), .YS(\mult_97/n1410 ) );
  FAX1 \mult_97/U1024  ( .A(\mult_97/n1416 ), .B(\mult_97/n1441 ), .C(
        \mult_97/n1414 ), .YC(\mult_97/n1407 ), .YS(\mult_97/n1408 ) );
  FAX1 \mult_97/U1023  ( .A(\mult_97/n1412 ), .B(\mult_97/n1439 ), .C(
        \mult_97/n1437 ), .YC(\mult_97/n1405 ), .YS(\mult_97/n1406 ) );
  FAX1 \mult_97/U1022  ( .A(\mult_97/n1410 ), .B(\mult_97/n1408 ), .C(
        \mult_97/n1435 ), .YC(n236), .YS(n235) );
  FAX1 \mult_97/U1021  ( .A(n417), .B(n418), .C(\mult_97/n1404 ), .YC(
        \mult_97/n1401 ), .YS(\mult_97/n1402 ) );
  OR2X2 \mult_97/U1020  ( .A(\mult_97/n2163 ), .B(\mult_97/n1981 ), .Y(
        \mult_97/n1399 ) );
  XNOR2X1 \mult_97/U1019  ( .A(\mult_97/n2163 ), .B(\mult_97/n1981 ), .Y(
        \mult_97/n1400 ) );
  FAX1 \mult_97/U1018  ( .A(\mult_97/n2254 ), .B(\mult_97/n1925 ), .C(
        \mult_97/n2347 ), .YC(\mult_97/n1397 ), .YS(\mult_97/n1398 ) );
  FAX1 \mult_97/U1017  ( .A(\mult_97/n2072 ), .B(\mult_97/n2194 ), .C(
        \mult_97/n2134 ), .YC(\mult_97/n1395 ), .YS(\mult_97/n1396 ) );
  FAX1 \mult_97/U1016  ( .A(\mult_97/n2012 ), .B(\mult_97/n2103 ), .C(
        \mult_97/n2043 ), .YC(\mult_97/n1393 ), .YS(\mult_97/n1394 ) );
  FAX1 \mult_97/U1015  ( .A(\mult_97/n2285 ), .B(\mult_97/n1896 ), .C(
        \mult_97/n1956 ), .YC(\mult_97/n1391 ), .YS(\mult_97/n1392 ) );
  FAX1 \mult_97/U1014  ( .A(\mult_97/n2316 ), .B(\mult_97/n2225 ), .C(
        \mult_97/n1429 ), .YC(\mult_97/n1389 ), .YS(\mult_97/n1390 ) );
  FAX1 \mult_97/U1013  ( .A(\mult_97/n1427 ), .B(\mult_97/n1421 ), .C(
        \mult_97/n1400 ), .YC(\mult_97/n1387 ), .YS(\mult_97/n1388 ) );
  FAX1 \mult_97/U1012  ( .A(\mult_97/n1425 ), .B(\mult_97/n1423 ), .C(
        \mult_97/n1419 ), .YC(\mult_97/n1385 ), .YS(\mult_97/n1386 ) );
  FAX1 \mult_97/U1011  ( .A(\mult_97/n1396 ), .B(\mult_97/n1394 ), .C(
        \mult_97/n1392 ), .YC(\mult_97/n1383 ), .YS(\mult_97/n1384 ) );
  FAX1 \mult_97/U1010  ( .A(\mult_97/n1398 ), .B(\mult_97/n1390 ), .C(
        \mult_97/n1417 ), .YC(\mult_97/n1381 ), .YS(\mult_97/n1382 ) );
  FAX1 \mult_97/U1009  ( .A(\mult_97/n1415 ), .B(\mult_97/n1413 ), .C(
        \mult_97/n1388 ), .YC(\mult_97/n1379 ), .YS(\mult_97/n1380 ) );
  FAX1 \mult_97/U1008  ( .A(\mult_97/n1386 ), .B(\mult_97/n1384 ), .C(
        \mult_97/n1411 ), .YC(\mult_97/n1377 ), .YS(\mult_97/n1378 ) );
  FAX1 \mult_97/U1007  ( .A(\mult_97/n1382 ), .B(\mult_97/n1409 ), .C(
        \mult_97/n1407 ), .YC(\mult_97/n1375 ), .YS(\mult_97/n1376 ) );
  FAX1 \mult_97/U1006  ( .A(n415), .B(n414), .C(n416), .YC(\mult_97/n1373 ), 
        .YS(\mult_97/n1374 ) );
  FAX1 \mult_97/U1005  ( .A(n412), .B(\mult_97/n1403 ), .C(\mult_97/n1374 ), 
        .YC(\mult_97/n1371 ), .YS(\mult_97/n1372 ) );
  FAX1 \mult_97/U1003  ( .A(\mult_97/n2071 ), .B(\mult_97/n2193 ), .C(
        \mult_97/n1955 ), .YC(\mult_97/n1367 ), .YS(\mult_97/n1368 ) );
  FAX1 \mult_97/U1002  ( .A(\mult_97/n1980 ), .B(\mult_97/n2011 ), .C(
        \mult_97/n2315 ), .YC(\mult_97/n1365 ), .YS(\mult_97/n1366 ) );
  FAX1 \mult_97/U1001  ( .A(\mult_97/n2162 ), .B(\mult_97/n1924 ), .C(
        \mult_97/n2224 ), .YC(\mult_97/n1363 ), .YS(\mult_97/n1364 ) );
  FAX1 \mult_97/U1000  ( .A(\mult_97/n2284 ), .B(\mult_97/n2102 ), .C(
        \mult_97/n2133 ), .YC(\mult_97/n1361 ), .YS(\mult_97/n1362 ) );
  FAX1 \mult_97/U999  ( .A(\mult_97/n1895 ), .B(\mult_97/n2042 ), .C(
        \mult_97/n1370 ), .YC(\mult_97/n1359 ), .YS(\mult_97/n1360 ) );
  FAX1 \mult_97/U998  ( .A(\mult_97/n1399 ), .B(\mult_97/n1397 ), .C(
        \mult_97/n1395 ), .YC(\mult_97/n1357 ), .YS(\mult_97/n1358 ) );
  FAX1 \mult_97/U997  ( .A(\mult_97/n1393 ), .B(\mult_97/n1391 ), .C(
        \mult_97/n1366 ), .YC(\mult_97/n1355 ), .YS(\mult_97/n1356 ) );
  FAX1 \mult_97/U996  ( .A(\mult_97/n1368 ), .B(\mult_97/n1362 ), .C(
        \mult_97/n1360 ), .YC(\mult_97/n1353 ), .YS(\mult_97/n1354 ) );
  FAX1 \mult_97/U995  ( .A(\mult_97/n1364 ), .B(\mult_97/n1389 ), .C(
        \mult_97/n1387 ), .YC(\mult_97/n1351 ), .YS(\mult_97/n1352 ) );
  FAX1 \mult_97/U994  ( .A(\mult_97/n1385 ), .B(\mult_97/n1358 ), .C(
        \mult_97/n1383 ), .YC(\mult_97/n1349 ), .YS(\mult_97/n1350 ) );
  FAX1 \mult_97/U993  ( .A(\mult_97/n1356 ), .B(\mult_97/n1354 ), .C(
        \mult_97/n1381 ), .YC(\mult_97/n1347 ), .YS(\mult_97/n1348 ) );
  FAX1 \mult_97/U992  ( .A(\mult_97/n1352 ), .B(\mult_97/n1379 ), .C(
        \mult_97/n1350 ), .YC(\mult_97/n1345 ), .YS(\mult_97/n1346 ) );
  FAX1 \mult_97/U991  ( .A(n413), .B(n520), .C(n411), .YC(\mult_97/n1343 ), 
        .YS(\mult_97/n1344 ) );
  FAX1 \mult_97/U990  ( .A(n518), .B(\mult_97/n1373 ), .C(\mult_97/n1344 ), 
        .YC(\mult_97/n1341 ), .YS(\mult_97/n1342 ) );
  FAX1 \mult_97/U989  ( .A(\mult_97/n1369 ), .B(\mult_97/n2192 ), .C(
        \mult_97/n1954 ), .YC(\mult_97/n1339 ), .YS(\mult_97/n1340 ) );
  FAX1 \mult_97/U988  ( .A(\mult_97/n1979 ), .B(\mult_97/n2101 ), .C(
        \mult_97/n2041 ), .YC(\mult_97/n1337 ), .YS(\mult_97/n1338 ) );
  FAX1 \mult_97/U987  ( .A(\mult_97/n2253 ), .B(\mult_97/n2010 ), .C(
        \mult_97/n2132 ), .YC(\mult_97/n1335 ), .YS(\mult_97/n1336 ) );
  FAX1 \mult_97/U986  ( .A(\mult_97/n2070 ), .B(\mult_97/n2283 ), .C(
        \mult_97/n2223 ), .YC(\mult_97/n1333 ), .YS(\mult_97/n1334 ) );
  FAX1 \mult_97/U985  ( .A(\mult_97/n2161 ), .B(\mult_97/n1923 ), .C(
        \mult_97/n1894 ), .YC(\mult_97/n1331 ), .YS(\mult_97/n1332 ) );
  FAX1 \mult_97/U984  ( .A(\mult_97/n2314 ), .B(\mult_97/n1367 ), .C(
        \mult_97/n1365 ), .YC(\mult_97/n1329 ), .YS(\mult_97/n1330 ) );
  FAX1 \mult_97/U983  ( .A(\mult_97/n1363 ), .B(\mult_97/n1361 ), .C(
        \mult_97/n1359 ), .YC(\mult_97/n1327 ), .YS(\mult_97/n1328 ) );
  FAX1 \mult_97/U982  ( .A(\mult_97/n1332 ), .B(\mult_97/n1340 ), .C(
        \mult_97/n1338 ), .YC(\mult_97/n1325 ), .YS(\mult_97/n1326 ) );
  FAX1 \mult_97/U981  ( .A(\mult_97/n1336 ), .B(\mult_97/n1334 ), .C(
        \mult_97/n1357 ), .YC(\mult_97/n1323 ), .YS(\mult_97/n1324 ) );
  FAX1 \mult_97/U980  ( .A(\mult_97/n1355 ), .B(\mult_97/n1330 ), .C(
        \mult_97/n1353 ), .YC(\mult_97/n1321 ), .YS(\mult_97/n1322 ) );
  FAX1 \mult_97/U979  ( .A(\mult_97/n1328 ), .B(\mult_97/n1326 ), .C(
        \mult_97/n1351 ), .YC(\mult_97/n1319 ), .YS(\mult_97/n1320 ) );
  FAX1 \mult_97/U978  ( .A(\mult_97/n1324 ), .B(\mult_97/n1349 ), .C(
        \mult_97/n1322 ), .YC(\mult_97/n1317 ), .YS(\mult_97/n1318 ) );
  FAX1 \mult_97/U977  ( .A(n519), .B(n516), .C(n517), .YC(\mult_97/n1315 ), 
        .YS(\mult_97/n1316 ) );
  FAX1 \mult_97/U976  ( .A(n514), .B(\mult_97/n1343 ), .C(\mult_97/n1316 ), 
        .YC(\mult_97/n1313 ), .YS(\mult_97/n1314 ) );
  FAX1 \mult_97/U974  ( .A(\mult_97/n2069 ), .B(\mult_97/n2009 ), .C(
        \mult_97/n2131 ), .YC(\mult_97/n1309 ), .YS(\mult_97/n1310 ) );
  FAX1 \mult_97/U973  ( .A(\mult_97/n1978 ), .B(\mult_97/n2100 ), .C(
        \mult_97/n2222 ), .YC(\mult_97/n1307 ), .YS(\mult_97/n1308 ) );
  FAX1 \mult_97/U972  ( .A(\mult_97/n2252 ), .B(\mult_97/n1922 ), .C(
        \mult_97/n2040 ), .YC(\mult_97/n1305 ), .YS(\mult_97/n1306 ) );
  FAX1 \mult_97/U971  ( .A(\mult_97/n2282 ), .B(\mult_97/n2191 ), .C(
        \mult_97/n1953 ), .YC(\mult_97/n1303 ), .YS(\mult_97/n1304 ) );
  FAX1 \mult_97/U970  ( .A(\mult_97/n1893 ), .B(\mult_97/n1312 ), .C(
        \mult_97/n1339 ), .YC(\mult_97/n1301 ), .YS(\mult_97/n1302 ) );
  FAX1 \mult_97/U969  ( .A(\mult_97/n1333 ), .B(\mult_97/n1337 ), .C(
        \mult_97/n1331 ), .YC(\mult_97/n1299 ), .YS(\mult_97/n1300 ) );
  FAX1 \mult_97/U968  ( .A(\mult_97/n1335 ), .B(\mult_97/n1308 ), .C(
        \mult_97/n1310 ), .YC(\mult_97/n1297 ), .YS(\mult_97/n1298 ) );
  FAX1 \mult_97/U967  ( .A(\mult_97/n1306 ), .B(\mult_97/n1304 ), .C(
        \mult_97/n1329 ), .YC(\mult_97/n1295 ), .YS(\mult_97/n1296 ) );
  FAX1 \mult_97/U966  ( .A(\mult_97/n1327 ), .B(\mult_97/n1302 ), .C(
        \mult_97/n1325 ), .YC(\mult_97/n1293 ), .YS(\mult_97/n1294 ) );
  FAX1 \mult_97/U965  ( .A(\mult_97/n1300 ), .B(\mult_97/n1298 ), .C(
        \mult_97/n1323 ), .YC(\mult_97/n1291 ), .YS(\mult_97/n1292 ) );
  FAX1 \mult_97/U964  ( .A(\mult_97/n1296 ), .B(\mult_97/n1321 ), .C(
        \mult_97/n1294 ), .YC(\mult_97/n1289 ), .YS(\mult_97/n1290 ) );
  FAX1 \mult_97/U963  ( .A(n515), .B(n512), .C(n513), .YC(\mult_97/n1287 ), 
        .YS(\mult_97/n1288 ) );
  FAX1 \mult_97/U962  ( .A(n510), .B(\mult_97/n1315 ), .C(\mult_97/n1288 ), 
        .YC(\mult_97/n1285 ), .YS(\mult_97/n1286 ) );
  FAX1 \mult_97/U961  ( .A(\mult_97/n1311 ), .B(\mult_97/n2099 ), .C(
        \mult_97/n2130 ), .YC(\mult_97/n1283 ), .YS(\mult_97/n1284 ) );
  FAX1 \mult_97/U960  ( .A(\mult_97/n2068 ), .B(\mult_97/n1921 ), .C(
        \mult_97/n1952 ), .YC(\mult_97/n1281 ), .YS(\mult_97/n1282 ) );
  FAX1 \mult_97/U959  ( .A(\mult_97/n1977 ), .B(\mult_97/n2190 ), .C(
        \mult_97/n2039 ), .YC(\mult_97/n1279 ), .YS(\mult_97/n1280 ) );
  FAX1 \mult_97/U958  ( .A(\mult_97/n2251 ), .B(\mult_97/n2008 ), .C(
        \mult_97/n2221 ), .YC(\mult_97/n1277 ), .YS(\mult_97/n1278 ) );
  FAX1 \mult_97/U957  ( .A(\mult_97/n2160 ), .B(\mult_97/n1892 ), .C(
        \mult_97/n2281 ), .YC(\mult_97/n1275 ), .YS(\mult_97/n1276 ) );
  FAX1 \mult_97/U956  ( .A(\mult_97/n1305 ), .B(\mult_97/n1309 ), .C(
        \mult_97/n1303 ), .YC(\mult_97/n1273 ), .YS(\mult_97/n1274 ) );
  FAX1 \mult_97/U955  ( .A(\mult_97/n1307 ), .B(\mult_97/n1278 ), .C(
        \mult_97/n1280 ), .YC(\mult_97/n1271 ), .YS(\mult_97/n1272 ) );
  FAX1 \mult_97/U954  ( .A(\mult_97/n1282 ), .B(\mult_97/n1284 ), .C(
        \mult_97/n1276 ), .YC(\mult_97/n1269 ), .YS(\mult_97/n1270 ) );
  FAX1 \mult_97/U953  ( .A(\mult_97/n1301 ), .B(\mult_97/n1299 ), .C(
        \mult_97/n1297 ), .YC(\mult_97/n1267 ), .YS(\mult_97/n1268 ) );
  FAX1 \mult_97/U952  ( .A(\mult_97/n1274 ), .B(\mult_97/n1272 ), .C(
        \mult_97/n1270 ), .YC(\mult_97/n1265 ), .YS(\mult_97/n1266 ) );
  FAX1 \mult_97/U951  ( .A(\mult_97/n1295 ), .B(\mult_97/n1293 ), .C(
        \mult_97/n1268 ), .YC(\mult_97/n1263 ), .YS(\mult_97/n1264 ) );
  FAX1 \mult_97/U950  ( .A(n511), .B(n508), .C(n509), .YC(\mult_97/n1261 ), 
        .YS(\mult_97/n1262 ) );
  FAX1 \mult_97/U949  ( .A(n507), .B(\mult_97/n1287 ), .C(\mult_97/n1262 ), 
        .YC(\mult_97/n1259 ), .YS(\mult_97/n1260 ) );
  FAX1 \mult_97/U947  ( .A(\mult_97/n2159 ), .B(\mult_97/n1920 ), .C(
        \mult_97/n2220 ), .YC(\mult_97/n1255 ), .YS(\mult_97/n1256 ) );
  FAX1 \mult_97/U946  ( .A(\mult_97/n1976 ), .B(\mult_97/n2098 ), .C(
        \mult_97/n1951 ), .YC(\mult_97/n1253 ), .YS(\mult_97/n1254 ) );
  FAX1 \mult_97/U945  ( .A(\mult_97/n2067 ), .B(\mult_97/n2007 ), .C(
        \mult_97/n2038 ), .YC(\mult_97/n1251 ), .YS(\mult_97/n1252 ) );
  FAX1 \mult_97/U944  ( .A(\mult_97/n2189 ), .B(\mult_97/n1891 ), .C(
        \mult_97/n2129 ), .YC(\mult_97/n1249 ), .YS(\mult_97/n1250 ) );
  FAX1 \mult_97/U943  ( .A(\mult_97/n1258 ), .B(\mult_97/n1283 ), .C(
        \mult_97/n1281 ), .YC(\mult_97/n1247 ), .YS(\mult_97/n1248 ) );
  FAX1 \mult_97/U942  ( .A(\mult_97/n1279 ), .B(\mult_97/n1277 ), .C(
        \mult_97/n1252 ), .YC(\mult_97/n1245 ), .YS(\mult_97/n1246 ) );
  FAX1 \mult_97/U941  ( .A(\mult_97/n1254 ), .B(\mult_97/n1256 ), .C(
        \mult_97/n1275 ), .YC(\mult_97/n1243 ), .YS(\mult_97/n1244 ) );
  FAX1 \mult_97/U940  ( .A(\mult_97/n1250 ), .B(\mult_97/n1273 ), .C(
        \mult_97/n1271 ), .YC(\mult_97/n1241 ), .YS(\mult_97/n1242 ) );
  FAX1 \mult_97/U939  ( .A(\mult_97/n1248 ), .B(\mult_97/n1246 ), .C(
        \mult_97/n1269 ), .YC(\mult_97/n1239 ), .YS(\mult_97/n1240 ) );
  FAX1 \mult_97/U938  ( .A(\mult_97/n1244 ), .B(\mult_97/n1267 ), .C(
        \mult_97/n1242 ), .YC(\mult_97/n1237 ), .YS(\mult_97/n1238 ) );
  FAX1 \mult_97/U937  ( .A(\mult_97/n1265 ), .B(\mult_97/n1240 ), .C(
        \mult_97/n1263 ), .YC(n234), .YS(n233) );
  FAX1 \mult_97/U936  ( .A(n506), .B(\mult_97/n1261 ), .C(\mult_97/n1236 ), 
        .YC(\mult_97/n1233 ), .YS(\mult_97/n1234 ) );
  FAX1 \mult_97/U935  ( .A(\mult_97/n1257 ), .B(\mult_97/n1919 ), .C(
        \mult_97/n2219 ), .YC(\mult_97/n1231 ), .YS(\mult_97/n1232 ) );
  FAX1 \mult_97/U934  ( .A(\mult_97/n2066 ), .B(\mult_97/n2006 ), .C(
        \mult_97/n1950 ), .YC(\mult_97/n1229 ), .YS(\mult_97/n1230 ) );
  FAX1 \mult_97/U933  ( .A(\mult_97/n2158 ), .B(\mult_97/n2188 ), .C(
        \mult_97/n2037 ), .YC(\mult_97/n1227 ), .YS(\mult_97/n1228 ) );
  FAX1 \mult_97/U932  ( .A(\mult_97/n1975 ), .B(\mult_97/n2097 ), .C(
        \mult_97/n2128 ), .YC(\mult_97/n1225 ), .YS(\mult_97/n1226 ) );
  FAX1 \mult_97/U931  ( .A(\mult_97/n1890 ), .B(\mult_97/n2250 ), .C(
        \mult_97/n1255 ), .YC(\mult_97/n1223 ), .YS(\mult_97/n1224 ) );
  FAX1 \mult_97/U930  ( .A(\mult_97/n1253 ), .B(\mult_97/n1251 ), .C(
        \mult_97/n1249 ), .YC(\mult_97/n1221 ), .YS(\mult_97/n1222 ) );
  FAX1 \mult_97/U929  ( .A(\mult_97/n1226 ), .B(\mult_97/n1232 ), .C(
        \mult_97/n1230 ), .YC(\mult_97/n1219 ), .YS(\mult_97/n1220 ) );
  FAX1 \mult_97/U928  ( .A(\mult_97/n1228 ), .B(\mult_97/n1247 ), .C(
        \mult_97/n1245 ), .YC(\mult_97/n1217 ), .YS(\mult_97/n1218 ) );
  FAX1 \mult_97/U927  ( .A(\mult_97/n1224 ), .B(\mult_97/n1243 ), .C(
        \mult_97/n1222 ), .YC(\mult_97/n1215 ), .YS(\mult_97/n1216 ) );
  FAX1 \mult_97/U926  ( .A(\mult_97/n1220 ), .B(\mult_97/n1241 ), .C(
        \mult_97/n1218 ), .YC(\mult_97/n1213 ), .YS(\mult_97/n1214 ) );
  FAX1 \mult_97/U925  ( .A(\mult_97/n1239 ), .B(\mult_97/n1216 ), .C(
        \mult_97/n1237 ), .YC(n232), .YS(n231) );
  FAX1 \mult_97/U924  ( .A(n505), .B(\mult_97/n1235 ), .C(\mult_97/n1212 ), 
        .YC(\mult_97/n1209 ), .YS(\mult_97/n1210 ) );
  FAX1 \mult_97/U922  ( .A(\mult_97/n2157 ), .B(\mult_97/n1918 ), .C(
        \mult_97/n2036 ), .YC(\mult_97/n1205 ), .YS(\mult_97/n1206 ) );
  FAX1 \mult_97/U921  ( .A(\mult_97/n1974 ), .B(\mult_97/n2096 ), .C(
        \mult_97/n2218 ), .YC(\mult_97/n1203 ), .YS(\mult_97/n1204 ) );
  FAX1 \mult_97/U920  ( .A(\mult_97/n2187 ), .B(\mult_97/n2005 ), .C(
        \mult_97/n1949 ), .YC(\mult_97/n1201 ), .YS(\mult_97/n1202 ) );
  FAX1 \mult_97/U919  ( .A(\mult_97/n1889 ), .B(\mult_97/n2127 ), .C(
        \mult_97/n1208 ), .YC(\mult_97/n1199 ), .YS(\mult_97/n1200 ) );
  FAX1 \mult_97/U918  ( .A(\mult_97/n1231 ), .B(\mult_97/n1225 ), .C(
        \mult_97/n1227 ), .YC(\mult_97/n1197 ), .YS(\mult_97/n1198 ) );
  FAX1 \mult_97/U917  ( .A(\mult_97/n1229 ), .B(\mult_97/n1206 ), .C(
        \mult_97/n1204 ), .YC(\mult_97/n1195 ), .YS(\mult_97/n1196 ) );
  FAX1 \mult_97/U916  ( .A(\mult_97/n1202 ), .B(\mult_97/n1200 ), .C(
        \mult_97/n1223 ), .YC(\mult_97/n1193 ), .YS(\mult_97/n1194 ) );
  FAX1 \mult_97/U915  ( .A(\mult_97/n1221 ), .B(\mult_97/n1219 ), .C(
        \mult_97/n1198 ), .YC(\mult_97/n1191 ), .YS(\mult_97/n1192 ) );
  FAX1 \mult_97/U914  ( .A(\mult_97/n1196 ), .B(\mult_97/n1194 ), .C(
        \mult_97/n1217 ), .YC(\mult_97/n1189 ), .YS(\mult_97/n1190 ) );
  FAX1 \mult_97/U913  ( .A(\mult_97/n1215 ), .B(\mult_97/n1192 ), .C(
        \mult_97/n1213 ), .YC(n230), .YS(n229) );
  FAX1 \mult_97/U912  ( .A(n504), .B(\mult_97/n1211 ), .C(\mult_97/n1188 ), 
        .YC(\mult_97/n1185 ), .YS(\mult_97/n1186 ) );
  FAX1 \mult_97/U911  ( .A(\mult_97/n1207 ), .B(\mult_97/n2004 ), .C(
        \mult_97/n2126 ), .YC(\mult_97/n1183 ), .YS(\mult_97/n1184 ) );
  FAX1 \mult_97/U910  ( .A(\mult_97/n2065 ), .B(\mult_97/n1917 ), .C(
        \mult_97/n1948 ), .YC(\mult_97/n1181 ), .YS(\mult_97/n1182 ) );
  FAX1 \mult_97/U909  ( .A(\mult_97/n1973 ), .B(\mult_97/n2095 ), .C(
        \mult_97/n2035 ), .YC(\mult_97/n1179 ), .YS(\mult_97/n1180 ) );
  FAX1 \mult_97/U908  ( .A(\mult_97/n2156 ), .B(\mult_97/n2186 ), .C(
        \mult_97/n1888 ), .YC(\mult_97/n1177 ), .YS(\mult_97/n1178 ) );
  FAX1 \mult_97/U907  ( .A(\mult_97/n2217 ), .B(\mult_97/n1205 ), .C(
        \mult_97/n1203 ), .YC(\mult_97/n1175 ), .YS(\mult_97/n1176 ) );
  FAX1 \mult_97/U906  ( .A(\mult_97/n1201 ), .B(\mult_97/n1199 ), .C(
        \mult_97/n1178 ), .YC(\mult_97/n1173 ), .YS(\mult_97/n1174 ) );
  FAX1 \mult_97/U905  ( .A(\mult_97/n1180 ), .B(\mult_97/n1184 ), .C(
        \mult_97/n1182 ), .YC(\mult_97/n1171 ), .YS(\mult_97/n1172 ) );
  FAX1 \mult_97/U904  ( .A(\mult_97/n1197 ), .B(\mult_97/n1195 ), .C(
        \mult_97/n1176 ), .YC(\mult_97/n1169 ), .YS(\mult_97/n1170 ) );
  FAX1 \mult_97/U903  ( .A(\mult_97/n1174 ), .B(\mult_97/n1172 ), .C(
        \mult_97/n1193 ), .YC(\mult_97/n1167 ), .YS(\mult_97/n1168 ) );
  FAX1 \mult_97/U902  ( .A(\mult_97/n1191 ), .B(\mult_97/n1170 ), .C(
        \mult_97/n1168 ), .YC(\mult_97/n1165 ), .YS(\mult_97/n1166 ) );
  FAX1 \mult_97/U901  ( .A(n503), .B(n502), .C(\mult_97/n1187 ), .YC(
        \mult_97/n1163 ), .YS(\mult_97/n1164 ) );
  FAX1 \mult_97/U899  ( .A(\mult_97/n2064 ), .B(\mult_97/n2185 ), .C(
        \mult_97/n2034 ), .YC(\mult_97/n1159 ), .YS(\mult_97/n1160 ) );
  FAX1 \mult_97/U898  ( .A(\mult_97/n2155 ), .B(\mult_97/n1916 ), .C(
        \mult_97/n2125 ), .YC(\mult_97/n1157 ), .YS(\mult_97/n1158 ) );
  FAX1 \mult_97/U897  ( .A(\mult_97/n2094 ), .B(\mult_97/n2003 ), .C(
        \mult_97/n1947 ), .YC(\mult_97/n1155 ), .YS(\mult_97/n1156 ) );
  FAX1 \mult_97/U896  ( .A(\mult_97/n1887 ), .B(\mult_97/n1162 ), .C(
        \mult_97/n1183 ), .YC(\mult_97/n1153 ), .YS(\mult_97/n1154 ) );
  FAX1 \mult_97/U895  ( .A(\mult_97/n1181 ), .B(\mult_97/n1177 ), .C(
        \mult_97/n1179 ), .YC(\mult_97/n1151 ), .YS(\mult_97/n1152 ) );
  FAX1 \mult_97/U894  ( .A(\mult_97/n1160 ), .B(\mult_97/n1158 ), .C(
        \mult_97/n1156 ), .YC(\mult_97/n1149 ), .YS(\mult_97/n1150 ) );
  FAX1 \mult_97/U893  ( .A(\mult_97/n1175 ), .B(\mult_97/n1154 ), .C(
        \mult_97/n1173 ), .YC(\mult_97/n1147 ), .YS(\mult_97/n1148 ) );
  FAX1 \mult_97/U892  ( .A(\mult_97/n1171 ), .B(\mult_97/n1152 ), .C(
        \mult_97/n1150 ), .YC(\mult_97/n1145 ), .YS(\mult_97/n1146 ) );
  FAX1 \mult_97/U891  ( .A(\mult_97/n1169 ), .B(\mult_97/n1148 ), .C(
        \mult_97/n1167 ), .YC(\mult_97/n1143 ), .YS(\mult_97/n1144 ) );
  FAX1 \mult_97/U890  ( .A(n500), .B(n501), .C(n499), .YC(\mult_97/n1141 ), 
        .YS(\mult_97/n1142 ) );
  FAX1 \mult_97/U889  ( .A(\mult_97/n1161 ), .B(\mult_97/n2002 ), .C(
        \mult_97/n2033 ), .YC(\mult_97/n1139 ), .YS(\mult_97/n1140 ) );
  FAX1 \mult_97/U888  ( .A(\mult_97/n2063 ), .B(\mult_97/n1915 ), .C(
        \mult_97/n2124 ), .YC(\mult_97/n1137 ), .YS(\mult_97/n1138 ) );
  FAX1 \mult_97/U887  ( .A(\mult_97/n2154 ), .B(\mult_97/n2093 ), .C(
        \mult_97/n1946 ), .YC(\mult_97/n1135 ), .YS(\mult_97/n1136 ) );
  FAX1 \mult_97/U886  ( .A(\mult_97/n1972 ), .B(\mult_97/n1886 ), .C(
        \mult_97/n2184 ), .YC(\mult_97/n1133 ), .YS(\mult_97/n1134 ) );
  FAX1 \mult_97/U885  ( .A(\mult_97/n1159 ), .B(\mult_97/n1157 ), .C(
        \mult_97/n1155 ), .YC(\mult_97/n1131 ), .YS(\mult_97/n1132 ) );
  FAX1 \mult_97/U884  ( .A(\mult_97/n1136 ), .B(\mult_97/n1140 ), .C(
        \mult_97/n1138 ), .YC(\mult_97/n1129 ), .YS(\mult_97/n1130 ) );
  FAX1 \mult_97/U883  ( .A(\mult_97/n1134 ), .B(\mult_97/n1153 ), .C(
        \mult_97/n1151 ), .YC(\mult_97/n1127 ), .YS(\mult_97/n1128 ) );
  FAX1 \mult_97/U882  ( .A(\mult_97/n1149 ), .B(\mult_97/n1132 ), .C(
        \mult_97/n1130 ), .YC(\mult_97/n1125 ), .YS(\mult_97/n1126 ) );
  FAX1 \mult_97/U881  ( .A(\mult_97/n1147 ), .B(\mult_97/n1128 ), .C(
        \mult_97/n1145 ), .YC(\mult_97/n1123 ), .YS(\mult_97/n1124 ) );
  FAX1 \mult_97/U880  ( .A(n497), .B(n498), .C(n496), .YC(\mult_97/n1121 ), 
        .YS(\mult_97/n1122 ) );
  FAX1 \mult_97/U878  ( .A(\mult_97/n1971 ), .B(\mult_97/n1914 ), .C(
        \mult_97/n2123 ), .YC(\mult_97/n1117 ), .YS(\mult_97/n1118 ) );
  FAX1 \mult_97/U877  ( .A(\mult_97/n2062 ), .B(\mult_97/n2001 ), .C(
        \mult_97/n1945 ), .YC(\mult_97/n1115 ), .YS(\mult_97/n1116 ) );
  FAX1 \mult_97/U876  ( .A(\mult_97/n2092 ), .B(\mult_97/n1885 ), .C(
        \mult_97/n2032 ), .YC(\mult_97/n1113 ), .YS(\mult_97/n1114 ) );
  FAX1 \mult_97/U875  ( .A(\mult_97/n1120 ), .B(\mult_97/n1139 ), .C(
        \mult_97/n1137 ), .YC(\mult_97/n1111 ), .YS(\mult_97/n1112 ) );
  FAX1 \mult_97/U874  ( .A(\mult_97/n1135 ), .B(\mult_97/n1116 ), .C(
        \mult_97/n1118 ), .YC(\mult_97/n1109 ), .YS(\mult_97/n1110 ) );
  FAX1 \mult_97/U873  ( .A(\mult_97/n1114 ), .B(\mult_97/n1133 ), .C(
        \mult_97/n1131 ), .YC(\mult_97/n1107 ), .YS(\mult_97/n1108 ) );
  FAX1 \mult_97/U872  ( .A(\mult_97/n1112 ), .B(\mult_97/n1129 ), .C(
        \mult_97/n1110 ), .YC(\mult_97/n1105 ), .YS(\mult_97/n1106 ) );
  FAX1 \mult_97/U871  ( .A(\mult_97/n1127 ), .B(\mult_97/n1108 ), .C(
        \mult_97/n1125 ), .YC(\mult_97/n1103 ), .YS(\mult_97/n1104 ) );
  FAX1 \mult_97/U870  ( .A(n494), .B(n495), .C(n493), .YC(\mult_97/n1101 ), 
        .YS(\mult_97/n1102 ) );
  FAX1 \mult_97/U869  ( .A(\mult_97/n1119 ), .B(\mult_97/n2000 ), .C(
        \mult_97/n1944 ), .YC(\mult_97/n1099 ), .YS(\mult_97/n1100 ) );
  FAX1 \mult_97/U868  ( .A(\mult_97/n2061 ), .B(\mult_97/n1913 ), .C(
        \mult_97/n2122 ), .YC(\mult_97/n1097 ), .YS(\mult_97/n1098 ) );
  FAX1 \mult_97/U867  ( .A(\mult_97/n1970 ), .B(\mult_97/n2091 ), .C(
        \mult_97/n2031 ), .YC(\mult_97/n1095 ), .YS(\mult_97/n1096 ) );
  FAX1 \mult_97/U866  ( .A(\mult_97/n1884 ), .B(\mult_97/n2153 ), .C(
        \mult_97/n1117 ), .YC(\mult_97/n1093 ), .YS(\mult_97/n1094 ) );
  FAX1 \mult_97/U865  ( .A(\mult_97/n1115 ), .B(\mult_97/n1113 ), .C(
        \mult_97/n1096 ), .YC(\mult_97/n1091 ), .YS(\mult_97/n1092 ) );
  FAX1 \mult_97/U864  ( .A(\mult_97/n1098 ), .B(\mult_97/n1100 ), .C(
        \mult_97/n1111 ), .YC(\mult_97/n1089 ), .YS(\mult_97/n1090 ) );
  FAX1 \mult_97/U863  ( .A(\mult_97/n1094 ), .B(\mult_97/n1109 ), .C(
        \mult_97/n1092 ), .YC(\mult_97/n1087 ), .YS(\mult_97/n1088 ) );
  FAX1 \mult_97/U862  ( .A(\mult_97/n1107 ), .B(\mult_97/n1090 ), .C(
        \mult_97/n1105 ), .YC(\mult_97/n1085 ), .YS(\mult_97/n1086 ) );
  FAX1 \mult_97/U861  ( .A(n491), .B(n492), .C(n490), .YC(\mult_97/n1083 ), 
        .YS(\mult_97/n1084 ) );
  FAX1 \mult_97/U859  ( .A(\mult_97/n2060 ), .B(\mult_97/n1912 ), .C(
        \mult_97/n2030 ), .YC(\mult_97/n1079 ), .YS(\mult_97/n1080 ) );
  FAX1 \mult_97/U858  ( .A(\mult_97/n2090 ), .B(\mult_97/n1999 ), .C(
        \mult_97/n1943 ), .YC(\mult_97/n1077 ), .YS(\mult_97/n1078 ) );
  FAX1 \mult_97/U857  ( .A(\mult_97/n1883 ), .B(\mult_97/n2121 ), .C(
        \mult_97/n1082 ), .YC(\mult_97/n1075 ), .YS(\mult_97/n1076 ) );
  FAX1 \mult_97/U856  ( .A(\mult_97/n1099 ), .B(\mult_97/n1095 ), .C(
        \mult_97/n1097 ), .YC(\mult_97/n1073 ), .YS(\mult_97/n1074 ) );
  FAX1 \mult_97/U855  ( .A(\mult_97/n1080 ), .B(\mult_97/n1078 ), .C(
        \mult_97/n1076 ), .YC(\mult_97/n1071 ), .YS(\mult_97/n1072 ) );
  FAX1 \mult_97/U854  ( .A(\mult_97/n1093 ), .B(\mult_97/n1091 ), .C(
        \mult_97/n1074 ), .YC(\mult_97/n1069 ), .YS(\mult_97/n1070 ) );
  FAX1 \mult_97/U853  ( .A(\mult_97/n1072 ), .B(\mult_97/n1089 ), .C(
        \mult_97/n1087 ), .YC(\mult_97/n1067 ), .YS(\mult_97/n1068 ) );
  FAX1 \mult_97/U852  ( .A(n488), .B(n489), .C(n487), .YC(\mult_97/n1065 ), 
        .YS(\mult_97/n1066 ) );
  FAX1 \mult_97/U851  ( .A(\mult_97/n1081 ), .B(\mult_97/n1911 ), .C(
        \mult_97/n1942 ), .YC(\mult_97/n1063 ), .YS(\mult_97/n1064 ) );
  FAX1 \mult_97/U850  ( .A(\mult_97/n2059 ), .B(\mult_97/n2089 ), .C(
        \mult_97/n2029 ), .YC(\mult_97/n1061 ), .YS(\mult_97/n1062 ) );
  FAX1 \mult_97/U849  ( .A(\mult_97/n1969 ), .B(\mult_97/n1998 ), .C(
        \mult_97/n1882 ), .YC(\mult_97/n1059 ), .YS(\mult_97/n1060 ) );
  FAX1 \mult_97/U848  ( .A(\mult_97/n2120 ), .B(\mult_97/n1079 ), .C(
        \mult_97/n1077 ), .YC(\mult_97/n1057 ), .YS(\mult_97/n1058 ) );
  FAX1 \mult_97/U847  ( .A(\mult_97/n1075 ), .B(\mult_97/n1060 ), .C(
        \mult_97/n1064 ), .YC(\mult_97/n1055 ), .YS(\mult_97/n1056 ) );
  FAX1 \mult_97/U846  ( .A(\mult_97/n1062 ), .B(\mult_97/n1073 ), .C(
        \mult_97/n1058 ), .YC(\mult_97/n1053 ), .YS(\mult_97/n1054 ) );
  FAX1 \mult_97/U845  ( .A(\mult_97/n1071 ), .B(\mult_97/n1056 ), .C(
        \mult_97/n1069 ), .YC(\mult_97/n1051 ), .YS(\mult_97/n1052 ) );
  FAX1 \mult_97/U844  ( .A(n485), .B(n486), .C(n484), .YC(\mult_97/n1049 ), 
        .YS(\mult_97/n1050 ) );
  FAX1 \mult_97/U842  ( .A(\mult_97/n2058 ), .B(\mult_97/n2088 ), .C(
        \mult_97/n2028 ), .YC(\mult_97/n1045 ), .YS(\mult_97/n1046 ) );
  FAX1 \mult_97/U841  ( .A(\mult_97/n1997 ), .B(\mult_97/n1910 ), .C(
        \mult_97/n1941 ), .YC(\mult_97/n1043 ), .YS(\mult_97/n1044 ) );
  FAX1 \mult_97/U840  ( .A(\mult_97/n1881 ), .B(\mult_97/n1048 ), .C(
        \mult_97/n1063 ), .YC(\mult_97/n1041 ), .YS(\mult_97/n1042 ) );
  FAX1 \mult_97/U839  ( .A(\mult_97/n1061 ), .B(\mult_97/n1059 ), .C(
        \mult_97/n1046 ), .YC(\mult_97/n1039 ), .YS(\mult_97/n1040 ) );
  FAX1 \mult_97/U838  ( .A(\mult_97/n1044 ), .B(\mult_97/n1057 ), .C(
        \mult_97/n1042 ), .YC(\mult_97/n1037 ), .YS(\mult_97/n1038 ) );
  FAX1 \mult_97/U837  ( .A(\mult_97/n1055 ), .B(\mult_97/n1040 ), .C(
        \mult_97/n1053 ), .YC(\mult_97/n1035 ), .YS(\mult_97/n1036 ) );
  FAX1 \mult_97/U836  ( .A(n482), .B(n483), .C(n481), .YC(\mult_97/n1033 ), 
        .YS(\mult_97/n1034 ) );
  FAX1 \mult_97/U835  ( .A(\mult_97/n1047 ), .B(\mult_97/n1996 ), .C(
        \mult_97/n2027 ), .YC(\mult_97/n1031 ), .YS(\mult_97/n1032 ) );
  FAX1 \mult_97/U834  ( .A(\mult_97/n2057 ), .B(\mult_97/n1909 ), .C(
        \mult_97/n1940 ), .YC(\mult_97/n1029 ), .YS(\mult_97/n1030 ) );
  FAX1 \mult_97/U833  ( .A(\mult_97/n1968 ), .B(\mult_97/n1880 ), .C(
        \mult_97/n2087 ), .YC(\mult_97/n1027 ), .YS(\mult_97/n1028 ) );
  FAX1 \mult_97/U832  ( .A(\mult_97/n1045 ), .B(\mult_97/n1043 ), .C(
        \mult_97/n1030 ), .YC(\mult_97/n1025 ), .YS(\mult_97/n1026 ) );
  FAX1 \mult_97/U831  ( .A(\mult_97/n1032 ), .B(\mult_97/n1028 ), .C(
        \mult_97/n1041 ), .YC(\mult_97/n1023 ), .YS(\mult_97/n1024 ) );
  FAX1 \mult_97/U830  ( .A(\mult_97/n1039 ), .B(\mult_97/n1026 ), .C(
        \mult_97/n1024 ), .YC(\mult_97/n1021 ), .YS(\mult_97/n1022 ) );
  FAX1 \mult_97/U829  ( .A(\mult_97/n1037 ), .B(\mult_97/n1035 ), .C(
        \mult_97/n1022 ), .YC(n228), .YS(n227) );
  FAX1 \mult_97/U827  ( .A(\mult_97/n1967 ), .B(\mult_97/n1908 ), .C(
        \mult_97/n2026 ), .YC(\mult_97/n1015 ), .YS(\mult_97/n1016 ) );
  FAX1 \mult_97/U826  ( .A(\mult_97/n1995 ), .B(\mult_97/n1879 ), .C(
        \mult_97/n1939 ), .YC(\mult_97/n1013 ), .YS(\mult_97/n1014 ) );
  FAX1 \mult_97/U825  ( .A(\mult_97/n1018 ), .B(\mult_97/n1031 ), .C(
        \mult_97/n1029 ), .YC(\mult_97/n1011 ), .YS(\mult_97/n1012 ) );
  FAX1 \mult_97/U824  ( .A(\mult_97/n1016 ), .B(\mult_97/n1014 ), .C(
        \mult_97/n1027 ), .YC(\mult_97/n1009 ), .YS(\mult_97/n1010 ) );
  FAX1 \mult_97/U823  ( .A(\mult_97/n1025 ), .B(\mult_97/n1012 ), .C(
        \mult_97/n1010 ), .YC(\mult_97/n1007 ), .YS(\mult_97/n1008 ) );
  FAX1 \mult_97/U822  ( .A(\mult_97/n1023 ), .B(\mult_97/n1008 ), .C(
        \mult_97/n1021 ), .YC(\mult_97/n1005 ), .YS(\mult_97/n1006 ) );
  FAX1 \mult_97/U821  ( .A(\mult_97/n1017 ), .B(\mult_97/n1994 ), .C(
        \mult_97/n1938 ), .YC(\mult_97/n1003 ), .YS(\mult_97/n1004 ) );
  FAX1 \mult_97/U820  ( .A(\mult_97/n1966 ), .B(\mult_97/n1907 ), .C(
        \mult_97/n2025 ), .YC(\mult_97/n1001 ), .YS(\mult_97/n1002 ) );
  FAX1 \mult_97/U819  ( .A(\mult_97/n1878 ), .B(\mult_97/n2056 ), .C(
        \mult_97/n1015 ), .YC(\mult_97/n999 ), .YS(\mult_97/n1000 ) );
  FAX1 \mult_97/U818  ( .A(\mult_97/n1013 ), .B(\mult_97/n1002 ), .C(
        \mult_97/n1004 ), .YC(\mult_97/n997 ), .YS(\mult_97/n998 ) );
  FAX1 \mult_97/U817  ( .A(\mult_97/n1011 ), .B(\mult_97/n1000 ), .C(
        \mult_97/n1009 ), .YC(\mult_97/n995 ), .YS(\mult_97/n996 ) );
  FAX1 \mult_97/U816  ( .A(\mult_97/n998 ), .B(\mult_97/n1007 ), .C(
        \mult_97/n996 ), .YC(\mult_97/n993 ), .YS(\mult_97/n994 ) );
  FAX1 \mult_97/U814  ( .A(\mult_97/n1993 ), .B(\mult_97/n1906 ), .C(
        \mult_97/n2024 ), .YC(\mult_97/n989 ), .YS(\mult_97/n990 ) );
  FAX1 \mult_97/U813  ( .A(\mult_97/n1877 ), .B(\mult_97/n1937 ), .C(
        \mult_97/n992 ), .YC(\mult_97/n987 ), .YS(\mult_97/n988 ) );
  FAX1 \mult_97/U812  ( .A(\mult_97/n1003 ), .B(\mult_97/n1001 ), .C(
        \mult_97/n990 ), .YC(\mult_97/n985 ), .YS(\mult_97/n986 ) );
  FAX1 \mult_97/U811  ( .A(\mult_97/n988 ), .B(\mult_97/n999 ), .C(
        \mult_97/n997 ), .YC(\mult_97/n983 ), .YS(\mult_97/n984 ) );
  FAX1 \mult_97/U810  ( .A(\mult_97/n986 ), .B(\mult_97/n995 ), .C(
        \mult_97/n984 ), .YC(\mult_97/n981 ), .YS(\mult_97/n982 ) );
  FAX1 \mult_97/U809  ( .A(\mult_97/n991 ), .B(\mult_97/n1992 ), .C(
        \mult_97/n1936 ), .YC(\mult_97/n979 ), .YS(\mult_97/n980 ) );
  FAX1 \mult_97/U808  ( .A(\mult_97/n1965 ), .B(\mult_97/n1905 ), .C(
        \mult_97/n1876 ), .YC(\mult_97/n977 ), .YS(\mult_97/n978 ) );
  FAX1 \mult_97/U807  ( .A(\mult_97/n2023 ), .B(\mult_97/n989 ), .C(
        \mult_97/n987 ), .YC(\mult_97/n975 ), .YS(\mult_97/n976 ) );
  FAX1 \mult_97/U806  ( .A(\mult_97/n978 ), .B(\mult_97/n980 ), .C(
        \mult_97/n985 ), .YC(\mult_97/n973 ), .YS(\mult_97/n974 ) );
  FAX1 \mult_97/U805  ( .A(\mult_97/n976 ), .B(\mult_97/n983 ), .C(
        \mult_97/n974 ), .YC(\mult_97/n971 ), .YS(\mult_97/n972 ) );
  FAX1 \mult_97/U803  ( .A(\mult_97/n1904 ), .B(\mult_97/n1991 ), .C(
        \mult_97/n1935 ), .YC(\mult_97/n967 ), .YS(\mult_97/n968 ) );
  FAX1 \mult_97/U802  ( .A(\mult_97/n1875 ), .B(\mult_97/n970 ), .C(
        \mult_97/n979 ), .YC(\mult_97/n965 ), .YS(\mult_97/n966 ) );
  FAX1 \mult_97/U801  ( .A(\mult_97/n977 ), .B(\mult_97/n968 ), .C(
        \mult_97/n975 ), .YC(\mult_97/n963 ), .YS(\mult_97/n964 ) );
  FAX1 \mult_97/U800  ( .A(\mult_97/n966 ), .B(\mult_97/n973 ), .C(
        \mult_97/n964 ), .YC(\mult_97/n961 ), .YS(\mult_97/n962 ) );
  FAX1 \mult_97/U799  ( .A(\mult_97/n969 ), .B(\mult_97/n1903 ), .C(
        \mult_97/n1934 ), .YC(\mult_97/n959 ), .YS(\mult_97/n960 ) );
  FAX1 \mult_97/U798  ( .A(\mult_97/n1964 ), .B(\mult_97/n1874 ), .C(
        \mult_97/n1990 ), .YC(\mult_97/n957 ), .YS(\mult_97/n958 ) );
  FAX1 \mult_97/U797  ( .A(\mult_97/n967 ), .B(\mult_97/n960 ), .C(
        \mult_97/n958 ), .YC(\mult_97/n955 ), .YS(\mult_97/n956 ) );
  FAX1 \mult_97/U796  ( .A(\mult_97/n965 ), .B(\mult_97/n956 ), .C(
        \mult_97/n963 ), .YC(\mult_97/n953 ), .YS(\mult_97/n954 ) );
  FAX1 \mult_97/U794  ( .A(\mult_97/n1902 ), .B(\mult_97/n1873 ), .C(
        \mult_97/n1933 ), .YC(\mult_97/n949 ), .YS(\mult_97/n950 ) );
  FAX1 \mult_97/U793  ( .A(\mult_97/n952 ), .B(\mult_97/n959 ), .C(
        \mult_97/n950 ), .YC(\mult_97/n947 ), .YS(\mult_97/n948 ) );
  FAX1 \mult_97/U792  ( .A(\mult_97/n957 ), .B(\mult_97/n948 ), .C(
        \mult_97/n955 ), .YC(\mult_97/n945 ), .YS(\mult_97/n946 ) );
  FAX1 \mult_97/U791  ( .A(\mult_97/n951 ), .B(\mult_97/n1901 ), .C(
        \mult_97/n1932 ), .YC(\mult_97/n943 ), .YS(\mult_97/n944 ) );
  FAX1 \mult_97/U790  ( .A(\mult_97/n1872 ), .B(\mult_97/n1963 ), .C(
        \mult_97/n949 ), .YC(\mult_97/n941 ), .YS(\mult_97/n942 ) );
  FAX1 \mult_97/U789  ( .A(\mult_97/n944 ), .B(\mult_97/n947 ), .C(
        \mult_97/n942 ), .YC(\mult_97/n939 ), .YS(\mult_97/n940 ) );
  FAX1 \mult_97/U787  ( .A(\mult_97/n1871 ), .B(\mult_97/n1931 ), .C(
        \mult_97/n938 ), .YC(\mult_97/n935 ), .YS(\mult_97/n936 ) );
  FAX1 \mult_97/U786  ( .A(\mult_97/n943 ), .B(\mult_97/n936 ), .C(
        \mult_97/n941 ), .YC(\mult_97/n933 ), .YS(\mult_97/n934 ) );
  FAX1 \mult_97/U785  ( .A(\mult_97/n937 ), .B(\mult_97/n1900 ), .C(
        \mult_97/n1870 ), .YC(\mult_97/n931 ), .YS(\mult_97/n932 ) );
  FAX1 \mult_97/U784  ( .A(\mult_97/n1930 ), .B(\mult_97/n935 ), .C(
        \mult_97/n932 ), .YC(\mult_97/n929 ), .YS(\mult_97/n930 ) );
  FAX1 \mult_97/U782  ( .A(\mult_97/n1869 ), .B(\mult_97/n928 ), .C(
        \mult_97/n931 ), .YC(\mult_97/n925 ), .YS(\mult_97/n926 ) );
  FAX1 \mult_97/U781  ( .A(\mult_97/n927 ), .B(\mult_97/n1868 ), .C(
        \mult_97/n1899 ), .YC(\mult_97/n923 ), .YS(\mult_97/n924 ) );
  NAND2X1 \mult_97/U779  ( .A(\mult_97/n2378 ), .B(\mult_97/n1866 ), .Y(
        \mult_97/n861 ) );
  NAND2X1 \mult_97/U773  ( .A(\mult_97/n2377 ), .B(\mult_97/n2346 ), .Y(
        \mult_97/n858 ) );
  AOI21X1 \mult_97/U767  ( .A(\mult_97/n859 ), .B(n529), .C(\mult_97/n856 ), 
        .Y(\mult_97/n854 ) );
  NAND2X1 \mult_97/U765  ( .A(\mult_97/n1865 ), .B(\mult_97/n1850 ), .Y(
        \mult_97/n853 ) );
  NOR2X1 \mult_97/U764  ( .A(\mult_97/n1865 ), .B(\mult_97/n1850 ), .Y(
        \mult_97/n852 ) );
  OAI21X1 \mult_97/U761  ( .A(\mult_97/n852 ), .B(\mult_97/n854 ), .C(
        \mult_97/n853 ), .Y(\mult_97/n851 ) );
  NAND2X1 \mult_97/U759  ( .A(\mult_97/n1849 ), .B(\mult_97/n1848 ), .Y(
        \mult_97/n850 ) );
  AOI21X1 \mult_97/U753  ( .A(n528), .B(\mult_97/n851 ), .C(\mult_97/n848 ), 
        .Y(\mult_97/n846 ) );
  NAND2X1 \mult_97/U751  ( .A(\mult_97/n1847 ), .B(\mult_97/n1844 ), .Y(
        \mult_97/n845 ) );
  NOR2X1 \mult_97/U750  ( .A(\mult_97/n1847 ), .B(\mult_97/n1844 ), .Y(
        \mult_97/n844 ) );
  OAI21X1 \mult_97/U747  ( .A(\mult_97/n844 ), .B(\mult_97/n846 ), .C(
        \mult_97/n845 ), .Y(\mult_97/n843 ) );
  NAND2X1 \mult_97/U744  ( .A(\mult_97/n1843 ), .B(\mult_97/n1840 ), .Y(
        \mult_97/n841 ) );
  NOR2X1 \mult_97/U743  ( .A(\mult_97/n1843 ), .B(\mult_97/n1840 ), .Y(
        \mult_97/n840 ) );
  NAND2X1 \mult_97/U738  ( .A(\mult_97/n1839 ), .B(\mult_97/n1834 ), .Y(
        \mult_97/n838 ) );
  NOR2X1 \mult_97/U737  ( .A(\mult_97/n1839 ), .B(\mult_97/n1834 ), .Y(
        \mult_97/n837 ) );
  OAI21X1 \mult_97/U734  ( .A(\mult_97/n841 ), .B(\mult_97/n837 ), .C(
        \mult_97/n838 ), .Y(\mult_97/n836 ) );
  NOR2X1 \mult_97/U733  ( .A(\mult_97/n840 ), .B(\mult_97/n837 ), .Y(
        \mult_97/n835 ) );
  AOI21X1 \mult_97/U732  ( .A(\mult_97/n843 ), .B(\mult_97/n835 ), .C(
        \mult_97/n836 ), .Y(\mult_97/n834 ) );
  NAND2X1 \mult_97/U730  ( .A(\mult_97/n1833 ), .B(\mult_97/n1828 ), .Y(
        \mult_97/n833 ) );
  NOR2X1 \mult_97/U729  ( .A(\mult_97/n1833 ), .B(\mult_97/n1828 ), .Y(
        \mult_97/n832 ) );
  OAI21X1 \mult_97/U726  ( .A(\mult_97/n832 ), .B(\mult_97/n834 ), .C(
        \mult_97/n833 ), .Y(\mult_97/n831 ) );
  NAND2X1 \mult_97/U723  ( .A(\mult_97/n1827 ), .B(\mult_97/n1820 ), .Y(
        \mult_97/n829 ) );
  NOR2X1 \mult_97/U722  ( .A(\mult_97/n1827 ), .B(\mult_97/n1820 ), .Y(
        \mult_97/n828 ) );
  OAI21X1 \mult_97/U719  ( .A(\mult_97/n828 ), .B(\mult_97/n830 ), .C(
        \mult_97/n829 ), .Y(\mult_97/n827 ) );
  NAND2X1 \mult_97/U717  ( .A(\mult_97/n1819 ), .B(\mult_97/n1812 ), .Y(
        \mult_97/n826 ) );
  NOR2X1 \mult_97/U716  ( .A(\mult_97/n1819 ), .B(\mult_97/n1812 ), .Y(
        \mult_97/n825 ) );
  NAND2X1 \mult_97/U714  ( .A(\mult_97/n826 ), .B(\mult_97/n911 ), .Y(
        \mult_97/n492 ) );
  XNOR2X1 \mult_97/U709  ( .A(\mult_97/n827 ), .B(\mult_97/n492 ), .Y(n226) );
  NAND2X1 \mult_97/U708  ( .A(\mult_97/n1811 ), .B(\mult_97/n1802 ), .Y(
        \mult_97/n820 ) );
  NAND2X1 \mult_97/U700  ( .A(\mult_97/n1801 ), .B(\mult_97/n1792 ), .Y(
        \mult_97/n815 ) );
  NAND2X1 \mult_97/U689  ( .A(\mult_97/n1791 ), .B(\mult_97/n1780 ), .Y(
        \mult_97/n807 ) );
  NOR2X1 \mult_97/U688  ( .A(\mult_97/n1791 ), .B(\mult_97/n1780 ), .Y(
        \mult_97/n806 ) );
  NAND2X1 \mult_97/U683  ( .A(\mult_97/n1779 ), .B(\mult_97/n1768 ), .Y(
        \mult_97/n804 ) );
  NOR2X1 \mult_97/U682  ( .A(\mult_97/n1779 ), .B(\mult_97/n1768 ), .Y(
        \mult_97/n803 ) );
  NAND2X1 \mult_97/U674  ( .A(\mult_97/n1767 ), .B(\mult_97/n1754 ), .Y(
        \mult_97/n798 ) );
  NAND2X1 \mult_97/U666  ( .A(\mult_97/n1753 ), .B(\mult_97/n1740 ), .Y(
        \mult_97/n793 ) );
  NOR2X1 \mult_97/U665  ( .A(\mult_97/n1753 ), .B(\mult_97/n1740 ), .Y(
        \mult_97/n792 ) );
  AOI21X1 \mult_97/U660  ( .A(\mult_97/n796 ), .B(\mult_97/n905 ), .C(
        \mult_97/n791 ), .Y(\mult_97/n789 ) );
  NAND2X1 \mult_97/U659  ( .A(n405), .B(\mult_97/n905 ), .Y(\mult_97/n788 ) );
  OAI21X1 \mult_97/U658  ( .A(\mult_97/n788 ), .B(\mult_97/n800 ), .C(
        \mult_97/n789 ), .Y(\mult_97/n787 ) );
  NAND2X1 \mult_97/U655  ( .A(\mult_97/n1739 ), .B(\mult_97/n1724 ), .Y(
        \mult_97/n781 ) );
  NOR2X1 \mult_97/U654  ( .A(\mult_97/n1739 ), .B(\mult_97/n1724 ), .Y(
        \mult_97/n780 ) );
  NAND2X1 \mult_97/U652  ( .A(n464), .B(\mult_97/n904 ), .Y(\mult_97/n485 ) );
  XOR2X1 \mult_97/U646  ( .A(\mult_97/n786 ), .B(\mult_97/n485 ), .Y(n678) );
  NAND2X1 \mult_97/U645  ( .A(\mult_97/n1723 ), .B(\mult_97/n1708 ), .Y(
        \mult_97/n778 ) );
  NOR2X1 \mult_97/U644  ( .A(\mult_97/n1723 ), .B(\mult_97/n1708 ), .Y(
        \mult_97/n777 ) );
  NAND2X1 \mult_97/U638  ( .A(\mult_97/n904 ), .B(\mult_97/n903 ), .Y(
        \mult_97/n773 ) );
  NAND2X1 \mult_97/U635  ( .A(n445), .B(n444), .Y(\mult_97/n771 ) );
  NOR2X1 \mult_97/U634  ( .A(n445), .B(n444), .Y(\mult_97/n770 ) );
  OAI21X1 \mult_97/U631  ( .A(\mult_97/n770 ), .B(\mult_97/n774 ), .C(
        \mult_97/n771 ), .Y(\mult_97/n769 ) );
  NOR2X1 \mult_97/U630  ( .A(\mult_97/n770 ), .B(\mult_97/n773 ), .Y(
        \mult_97/n768 ) );
  AOI21X1 \mult_97/U629  ( .A(\mult_97/n787 ), .B(\mult_97/n768 ), .C(
        \mult_97/n769 ), .Y(\mult_97/n767 ) );
  NAND2X1 \mult_97/U626  ( .A(n443), .B(\mult_97/n1672 ), .Y(\mult_97/n765 )
         );
  NOR2X1 \mult_97/U625  ( .A(n443), .B(\mult_97/n1672 ), .Y(\mult_97/n764 ) );
  NAND2X1 \mult_97/U618  ( .A(\mult_97/n1671 ), .B(\mult_97/n1652 ), .Y(
        \mult_97/n760 ) );
  NOR2X1 \mult_97/U617  ( .A(\mult_97/n1671 ), .B(\mult_97/n1652 ), .Y(
        \mult_97/n759 ) );
  OAI21X1 \mult_97/U614  ( .A(\mult_97/n765 ), .B(\mult_97/n759 ), .C(
        \mult_97/n760 ), .Y(\mult_97/n758 ) );
  NOR2X1 \mult_97/U613  ( .A(\mult_97/n764 ), .B(\mult_97/n759 ), .Y(
        \mult_97/n757 ) );
  AOI21X1 \mult_97/U612  ( .A(\mult_97/n757 ), .B(\mult_97/n766 ), .C(
        \mult_97/n758 ), .Y(\mult_97/n756 ) );
  NAND2X1 \mult_97/U610  ( .A(\mult_97/n1651 ), .B(\mult_97/n1632 ), .Y(
        \mult_97/n755 ) );
  NOR2X1 \mult_97/U609  ( .A(\mult_97/n1651 ), .B(\mult_97/n1632 ), .Y(
        \mult_97/n754 ) );
  NAND2X1 \mult_97/U604  ( .A(\mult_97/n1631 ), .B(\mult_97/n1610 ), .Y(
        \mult_97/n752 ) );
  NOR2X1 \mult_97/U603  ( .A(\mult_97/n1631 ), .B(\mult_97/n1610 ), .Y(
        \mult_97/n751 ) );
  OAI21X1 \mult_97/U600  ( .A(\mult_97/n755 ), .B(\mult_97/n751 ), .C(
        \mult_97/n752 ), .Y(\mult_97/n750 ) );
  NOR2X1 \mult_97/U599  ( .A(\mult_97/n754 ), .B(\mult_97/n751 ), .Y(
        \mult_97/n749 ) );
  AOI21X1 \mult_97/U598  ( .A(\mult_97/n758 ), .B(\mult_97/n749 ), .C(
        \mult_97/n750 ), .Y(\mult_97/n748 ) );
  NAND2X1 \mult_97/U597  ( .A(\mult_97/n757 ), .B(\mult_97/n749 ), .Y(
        \mult_97/n747 ) );
  OAI21X1 \mult_97/U596  ( .A(\mult_97/n767 ), .B(\mult_97/n747 ), .C(
        \mult_97/n748 ), .Y(\mult_97/n746 ) );
  NAND2X1 \mult_97/U593  ( .A(\mult_97/n1609 ), .B(\mult_97/n1588 ), .Y(
        \mult_97/n740 ) );
  NOR2X1 \mult_97/U592  ( .A(\mult_97/n1609 ), .B(\mult_97/n1588 ), .Y(
        \mult_97/n739 ) );
  NAND2X1 \mult_97/U590  ( .A(\mult_97/n740 ), .B(\mult_97/n897 ), .Y(
        \mult_97/n478 ) );
  XOR2X1 \mult_97/U584  ( .A(\mult_97/n745 ), .B(\mult_97/n478 ), .Y(n671) );
  NAND2X1 \mult_97/U583  ( .A(\mult_97/n1587 ), .B(\mult_97/n1564 ), .Y(
        \mult_97/n737 ) );
  NAND2X1 \mult_97/U576  ( .A(\mult_97/n897 ), .B(n533), .Y(\mult_97/n732 ) );
  OAI21X1 \mult_97/U575  ( .A(\mult_97/n732 ), .B(\mult_97/n745 ), .C(
        \mult_97/n733 ), .Y(\mult_97/n731 ) );
  NAND2X1 \mult_97/U573  ( .A(\mult_97/n1563 ), .B(\mult_97/n1540 ), .Y(
        \mult_97/n730 ) );
  NAND2X1 \mult_97/U565  ( .A(\mult_97/n1539 ), .B(\mult_97/n1514 ), .Y(
        \mult_97/n725 ) );
  AOI21X1 \mult_97/U559  ( .A(\mult_97/n728 ), .B(n556), .C(\mult_97/n723 ), 
        .Y(\mult_97/n721 ) );
  NAND2X1 \mult_97/U558  ( .A(n531), .B(n556), .Y(\mult_97/n720 ) );
  OAI21X1 \mult_97/U557  ( .A(\mult_97/n733 ), .B(\mult_97/n720 ), .C(
        \mult_97/n721 ), .Y(\mult_97/n719 ) );
  NOR2X1 \mult_97/U556  ( .A(\mult_97/n732 ), .B(\mult_97/n720 ), .Y(
        \mult_97/n718 ) );
  AOI21X1 \mult_97/U555  ( .A(\mult_97/n718 ), .B(\mult_97/n746 ), .C(
        \mult_97/n719 ), .Y(\mult_97/n717 ) );
  NAND2X1 \mult_97/U552  ( .A(\mult_97/n1513 ), .B(\mult_97/n1488 ), .Y(
        \mult_97/n715 ) );
  NOR2X1 \mult_97/U551  ( .A(\mult_97/n1513 ), .B(\mult_97/n1488 ), .Y(
        \mult_97/n714 ) );
  NAND2X1 \mult_97/U544  ( .A(\mult_97/n1487 ), .B(\mult_97/n1460 ), .Y(
        \mult_97/n710 ) );
  NOR2X1 \mult_97/U543  ( .A(\mult_97/n1487 ), .B(\mult_97/n1460 ), .Y(
        \mult_97/n709 ) );
  OAI21X1 \mult_97/U540  ( .A(\mult_97/n715 ), .B(\mult_97/n709 ), .C(
        \mult_97/n710 ), .Y(\mult_97/n708 ) );
  NOR2X1 \mult_97/U539  ( .A(\mult_97/n714 ), .B(\mult_97/n709 ), .Y(
        \mult_97/n707 ) );
  AOI21X1 \mult_97/U538  ( .A(\mult_97/n707 ), .B(\mult_97/n716 ), .C(
        \mult_97/n708 ), .Y(\mult_97/n706 ) );
  NAND2X1 \mult_97/U536  ( .A(\mult_97/n1459 ), .B(\mult_97/n1432 ), .Y(
        \mult_97/n705 ) );
  NOR2X1 \mult_97/U535  ( .A(\mult_97/n1459 ), .B(\mult_97/n1432 ), .Y(
        \mult_97/n704 ) );
  NAND2X1 \mult_97/U530  ( .A(\mult_97/n1431 ), .B(\mult_97/n1402 ), .Y(
        \mult_97/n702 ) );
  NOR2X1 \mult_97/U529  ( .A(\mult_97/n1431 ), .B(\mult_97/n1402 ), .Y(
        \mult_97/n701 ) );
  OAI21X1 \mult_97/U526  ( .A(\mult_97/n705 ), .B(\mult_97/n701 ), .C(
        \mult_97/n702 ), .Y(\mult_97/n700 ) );
  NOR2X1 \mult_97/U525  ( .A(\mult_97/n704 ), .B(\mult_97/n701 ), .Y(
        \mult_97/n699 ) );
  AOI21X1 \mult_97/U524  ( .A(\mult_97/n708 ), .B(\mult_97/n699 ), .C(
        \mult_97/n700 ), .Y(\mult_97/n698 ) );
  NAND2X1 \mult_97/U523  ( .A(\mult_97/n707 ), .B(\mult_97/n699 ), .Y(
        \mult_97/n697 ) );
  OAI21X1 \mult_97/U522  ( .A(\mult_97/n697 ), .B(\mult_97/n717 ), .C(
        \mult_97/n698 ), .Y(\mult_97/n696 ) );
  NAND2X1 \mult_97/U519  ( .A(\mult_97/n1401 ), .B(\mult_97/n1372 ), .Y(
        \mult_97/n694 ) );
  NOR2X1 \mult_97/U518  ( .A(\mult_97/n1401 ), .B(\mult_97/n1372 ), .Y(
        \mult_97/n693 ) );
  NAND2X1 \mult_97/U513  ( .A(\mult_97/n1371 ), .B(\mult_97/n1342 ), .Y(
        \mult_97/n691 ) );
  NOR2X1 \mult_97/U512  ( .A(\mult_97/n1371 ), .B(\mult_97/n1342 ), .Y(
        \mult_97/n690 ) );
  OAI21X1 \mult_97/U509  ( .A(\mult_97/n694 ), .B(\mult_97/n690 ), .C(
        \mult_97/n691 ), .Y(\mult_97/n689 ) );
  NOR2X1 \mult_97/U508  ( .A(\mult_97/n693 ), .B(\mult_97/n690 ), .Y(
        \mult_97/n688 ) );
  OAI21X1 \mult_97/U505  ( .A(\mult_97/n686 ), .B(\mult_97/n695 ), .C(
        \mult_97/n687 ), .Y(\mult_97/n685 ) );
  NAND2X1 \mult_97/U503  ( .A(\mult_97/n1341 ), .B(\mult_97/n1314 ), .Y(
        \mult_97/n684 ) );
  NOR2X1 \mult_97/U502  ( .A(\mult_97/n1341 ), .B(\mult_97/n1314 ), .Y(
        \mult_97/n683 ) );
  NAND2X1 \mult_97/U495  ( .A(\mult_97/n1313 ), .B(\mult_97/n1286 ), .Y(
        \mult_97/n679 ) );
  NOR2X1 \mult_97/U494  ( .A(\mult_97/n1313 ), .B(\mult_97/n1286 ), .Y(
        \mult_97/n678 ) );
  OAI21X1 \mult_97/U491  ( .A(\mult_97/n684 ), .B(\mult_97/n678 ), .C(
        \mult_97/n679 ), .Y(\mult_97/n677 ) );
  NOR2X1 \mult_97/U490  ( .A(\mult_97/n678 ), .B(\mult_97/n683 ), .Y(
        \mult_97/n676 ) );
  AOI21X1 \mult_97/U489  ( .A(\mult_97/n689 ), .B(\mult_97/n676 ), .C(
        \mult_97/n677 ), .Y(\mult_97/n675 ) );
  NAND2X1 \mult_97/U488  ( .A(\mult_97/n688 ), .B(\mult_97/n676 ), .Y(
        \mult_97/n674 ) );
  OAI21X1 \mult_97/U487  ( .A(\mult_97/n674 ), .B(\mult_97/n695 ), .C(
        \mult_97/n675 ), .Y(\mult_97/n673 ) );
  NAND2X1 \mult_97/U484  ( .A(\mult_97/n1285 ), .B(\mult_97/n1260 ), .Y(
        \mult_97/n671 ) );
  NOR2X1 \mult_97/U483  ( .A(\mult_97/n1285 ), .B(\mult_97/n1260 ), .Y(
        \mult_97/n670 ) );
  NAND2X1 \mult_97/U481  ( .A(\mult_97/n671 ), .B(\mult_97/n885 ), .Y(
        \mult_97/n466 ) );
  XOR2X1 \mult_97/U477  ( .A(\mult_97/n672 ), .B(\mult_97/n466 ), .Y(n659) );
  NAND2X1 \mult_97/U476  ( .A(\mult_97/n1259 ), .B(\mult_97/n1234 ), .Y(
        \mult_97/n666 ) );
  NOR2X1 \mult_97/U475  ( .A(\mult_97/n1259 ), .B(\mult_97/n1234 ), .Y(
        \mult_97/n665 ) );
  OAI21X1 \mult_97/U472  ( .A(\mult_97/n671 ), .B(\mult_97/n665 ), .C(
        \mult_97/n666 ), .Y(\mult_97/n664 ) );
  NOR2X1 \mult_97/U471  ( .A(\mult_97/n665 ), .B(\mult_97/n670 ), .Y(
        \mult_97/n663 ) );
  OAI21X1 \mult_97/U468  ( .A(\mult_97/n661 ), .B(\mult_97/n672 ), .C(
        \mult_97/n662 ), .Y(\mult_97/n660 ) );
  NAND2X1 \mult_97/U466  ( .A(\mult_97/n1233 ), .B(\mult_97/n1210 ), .Y(
        \mult_97/n659 ) );
  NOR2X1 \mult_97/U465  ( .A(\mult_97/n1233 ), .B(\mult_97/n1210 ), .Y(
        \mult_97/n658 ) );
  NAND2X1 \mult_97/U458  ( .A(\mult_97/n1209 ), .B(\mult_97/n1186 ), .Y(
        \mult_97/n654 ) );
  NOR2X1 \mult_97/U457  ( .A(\mult_97/n1209 ), .B(\mult_97/n1186 ), .Y(
        \mult_97/n653 ) );
  OAI21X1 \mult_97/U454  ( .A(\mult_97/n659 ), .B(\mult_97/n653 ), .C(
        \mult_97/n654 ), .Y(\mult_97/n652 ) );
  NOR2X1 \mult_97/U453  ( .A(\mult_97/n653 ), .B(\mult_97/n658 ), .Y(
        \mult_97/n651 ) );
  AOI21X1 \mult_97/U452  ( .A(\mult_97/n664 ), .B(\mult_97/n651 ), .C(
        \mult_97/n652 ), .Y(\mult_97/n650 ) );
  NAND2X1 \mult_97/U451  ( .A(\mult_97/n651 ), .B(\mult_97/n663 ), .Y(
        \mult_97/n649 ) );
  OAI21X1 \mult_97/U450  ( .A(\mult_97/n649 ), .B(\mult_97/n675 ), .C(
        \mult_97/n650 ), .Y(\mult_97/n648 ) );
  NOR2X1 \mult_97/U449  ( .A(\mult_97/n649 ), .B(\mult_97/n674 ), .Y(
        \mult_97/n647 ) );
  AOI21X1 \mult_97/U448  ( .A(\mult_97/n696 ), .B(\mult_97/n647 ), .C(
        \mult_97/n648 ), .Y(\mult_97/n646 ) );
  NAND2X1 \mult_97/U445  ( .A(\mult_97/n1185 ), .B(\mult_97/n1164 ), .Y(
        \mult_97/n644 ) );
  NOR2X1 \mult_97/U444  ( .A(\mult_97/n1185 ), .B(\mult_97/n1164 ), .Y(
        \mult_97/n643 ) );
  AOI21X1 \mult_97/U439  ( .A(\mult_97/n881 ), .B(\mult_97/n645 ), .C(
        \mult_97/n642 ), .Y(\mult_97/n640 ) );
  NAND2X1 \mult_97/U437  ( .A(\mult_97/n1142 ), .B(\mult_97/n1163 ), .Y(
        \mult_97/n635 ) );
  NOR2X1 \mult_97/U436  ( .A(\mult_97/n1142 ), .B(\mult_97/n1163 ), .Y(
        \mult_97/n634 ) );
  NAND2X1 \mult_97/U434  ( .A(\mult_97/n635 ), .B(\mult_97/n880 ), .Y(
        \mult_97/n461 ) );
  XOR2X1 \mult_97/U428  ( .A(\mult_97/n640 ), .B(\mult_97/n461 ), .Y(n654) );
  NAND2X1 \mult_97/U427  ( .A(\mult_97/n1122 ), .B(\mult_97/n1141 ), .Y(
        \mult_97/n632 ) );
  AOI21X1 \mult_97/U421  ( .A(n530), .B(\mult_97/n637 ), .C(\mult_97/n630 ), 
        .Y(\mult_97/n628 ) );
  NAND2X1 \mult_97/U420  ( .A(n530), .B(\mult_97/n880 ), .Y(\mult_97/n627 ) );
  OAI21X1 \mult_97/U419  ( .A(\mult_97/n644 ), .B(\mult_97/n627 ), .C(
        \mult_97/n628 ), .Y(\mult_97/n626 ) );
  NOR2X1 \mult_97/U418  ( .A(\mult_97/n643 ), .B(\mult_97/n627 ), .Y(
        \mult_97/n625 ) );
  AOI21X1 \mult_97/U417  ( .A(\mult_97/n625 ), .B(\mult_97/n645 ), .C(
        \mult_97/n626 ), .Y(\mult_97/n624 ) );
  NAND2X1 \mult_97/U414  ( .A(\mult_97/n1121 ), .B(\mult_97/n1102 ), .Y(
        \mult_97/n618 ) );
  NOR2X1 \mult_97/U413  ( .A(\mult_97/n1121 ), .B(\mult_97/n1102 ), .Y(
        \mult_97/n617 ) );
  NAND2X1 \mult_97/U404  ( .A(\mult_97/n1101 ), .B(\mult_97/n1084 ), .Y(
        \mult_97/n615 ) );
  AOI21X1 \mult_97/U398  ( .A(\mult_97/n620 ), .B(n532), .C(\mult_97/n613 ), 
        .Y(\mult_97/n611 ) );
  NAND2X1 \mult_97/U397  ( .A(n532), .B(\mult_97/n878 ), .Y(\mult_97/n610 ) );
  AOI21X1 \mult_97/U394  ( .A(\mult_97/n608 ), .B(\mult_97/n623 ), .C(
        \mult_97/n609 ), .Y(\mult_97/n607 ) );
  NAND2X1 \mult_97/U391  ( .A(\mult_97/n1083 ), .B(\mult_97/n1066 ), .Y(
        \mult_97/n605 ) );
  NOR2X1 \mult_97/U390  ( .A(\mult_97/n1083 ), .B(\mult_97/n1066 ), .Y(
        \mult_97/n604 ) );
  NAND2X1 \mult_97/U383  ( .A(\mult_97/n1065 ), .B(\mult_97/n1050 ), .Y(
        \mult_97/n600 ) );
  NOR2X1 \mult_97/U382  ( .A(\mult_97/n1065 ), .B(\mult_97/n1050 ), .Y(
        \mult_97/n599 ) );
  OAI21X1 \mult_97/U379  ( .A(\mult_97/n605 ), .B(\mult_97/n599 ), .C(
        \mult_97/n600 ), .Y(\mult_97/n598 ) );
  NOR2X1 \mult_97/U378  ( .A(\mult_97/n599 ), .B(\mult_97/n604 ), .Y(
        \mult_97/n597 ) );
  OAI21X1 \mult_97/U375  ( .A(\mult_97/n595 ), .B(\mult_97/n607 ), .C(
        \mult_97/n596 ), .Y(\mult_97/n594 ) );
  NAND2X1 \mult_97/U373  ( .A(\mult_97/n1049 ), .B(\mult_97/n1034 ), .Y(
        \mult_97/n593 ) );
  NOR2X1 \mult_97/U372  ( .A(\mult_97/n1049 ), .B(\mult_97/n1034 ), .Y(
        \mult_97/n592 ) );
  NAND2X1 \mult_97/U365  ( .A(\mult_97/n1033 ), .B(\mult_97/n1020 ), .Y(
        \mult_97/n588 ) );
  NOR2X1 \mult_97/U364  ( .A(\mult_97/n1033 ), .B(\mult_97/n1020 ), .Y(
        \mult_97/n587 ) );
  OAI21X1 \mult_97/U361  ( .A(\mult_97/n593 ), .B(\mult_97/n587 ), .C(
        \mult_97/n588 ), .Y(\mult_97/n586 ) );
  NOR2X1 \mult_97/U360  ( .A(\mult_97/n587 ), .B(\mult_97/n592 ), .Y(
        \mult_97/n585 ) );
  AOI21X1 \mult_97/U359  ( .A(\mult_97/n585 ), .B(\mult_97/n598 ), .C(
        \mult_97/n586 ), .Y(\mult_97/n584 ) );
  NAND2X1 \mult_97/U358  ( .A(\mult_97/n585 ), .B(\mult_97/n597 ), .Y(
        \mult_97/n583 ) );
  OAI21X1 \mult_97/U357  ( .A(\mult_97/n611 ), .B(\mult_97/n583 ), .C(
        \mult_97/n584 ), .Y(\mult_97/n582 ) );
  NOR2X1 \mult_97/U356  ( .A(\mult_97/n610 ), .B(\mult_97/n583 ), .Y(
        \mult_97/n581 ) );
  AOI21X1 \mult_97/U355  ( .A(\mult_97/n626 ), .B(\mult_97/n581 ), .C(
        \mult_97/n582 ), .Y(\mult_97/n580 ) );
  NAND2X1 \mult_97/U354  ( .A(\mult_97/n625 ), .B(\mult_97/n581 ), .Y(
        \mult_97/n579 ) );
  AOI21X1 \mult_97/U351  ( .A(\mult_97/n577 ), .B(\mult_97/n645 ), .C(
        \mult_97/n578 ), .Y(\mult_97/n576 ) );
  NAND2X1 \mult_97/U348  ( .A(n480), .B(\mult_97/n1019 ), .Y(\mult_97/n570 )
         );
  NOR2X1 \mult_97/U347  ( .A(n480), .B(\mult_97/n1019 ), .Y(\mult_97/n569 ) );
  NAND2X1 \mult_97/U338  ( .A(\mult_97/n994 ), .B(\mult_97/n1005 ), .Y(
        \mult_97/n567 ) );
  NOR2X1 \mult_97/U337  ( .A(\mult_97/n994 ), .B(\mult_97/n1005 ), .Y(
        \mult_97/n566 ) );
  AOI21X1 \mult_97/U332  ( .A(\mult_97/n871 ), .B(\mult_97/n572 ), .C(
        \mult_97/n565 ), .Y(\mult_97/n563 ) );
  NAND2X1 \mult_97/U331  ( .A(\mult_97/n871 ), .B(\mult_97/n872 ), .Y(
        \mult_97/n562 ) );
  AOI21X1 \mult_97/U328  ( .A(\mult_97/n560 ), .B(\mult_97/n575 ), .C(
        \mult_97/n561 ), .Y(\mult_97/n559 ) );
  NAND2X1 \mult_97/U325  ( .A(\mult_97/n993 ), .B(\mult_97/n982 ), .Y(
        \mult_97/n557 ) );
  NOR2X1 \mult_97/U324  ( .A(\mult_97/n993 ), .B(\mult_97/n982 ), .Y(
        \mult_97/n556 ) );
  NAND2X1 \mult_97/U319  ( .A(\mult_97/n981 ), .B(\mult_97/n972 ), .Y(
        \mult_97/n554 ) );
  NOR2X1 \mult_97/U318  ( .A(\mult_97/n981 ), .B(\mult_97/n972 ), .Y(
        \mult_97/n553 ) );
  OAI21X1 \mult_97/U309  ( .A(n458), .B(n455), .C(n456), .Y(\mult_97/n552 ) );
  NOR2X1 \mult_97/U308  ( .A(n455), .B(n457), .Y(\mult_97/n551 ) );
  NAND2X1 \mult_97/U305  ( .A(\mult_97/n971 ), .B(\mult_97/n962 ), .Y(
        \mult_97/n549 ) );
  NOR2X1 \mult_97/U304  ( .A(\mult_97/n971 ), .B(\mult_97/n962 ), .Y(
        \mult_97/n548 ) );
  AOI21X1 \mult_97/U299  ( .A(\mult_97/n868 ), .B(\mult_97/n552 ), .C(
        \mult_97/n547 ), .Y(\mult_97/n545 ) );
  NAND2X1 \mult_97/U298  ( .A(\mult_97/n868 ), .B(\mult_97/n551 ), .Y(
        \mult_97/n544 ) );
  OAI21X1 \mult_97/U297  ( .A(\mult_97/n563 ), .B(\mult_97/n544 ), .C(
        \mult_97/n545 ), .Y(\mult_97/n543 ) );
  NOR2X1 \mult_97/U296  ( .A(\mult_97/n544 ), .B(\mult_97/n562 ), .Y(
        \mult_97/n542 ) );
  AOI21X1 \mult_97/U295  ( .A(\mult_97/n542 ), .B(\mult_97/n575 ), .C(
        \mult_97/n543 ), .Y(\mult_97/n541 ) );
  NAND2X1 \mult_97/U293  ( .A(\mult_97/n961 ), .B(\mult_97/n954 ), .Y(
        \mult_97/n540 ) );
  NAND2X1 \mult_97/U290  ( .A(n452), .B(n406), .Y(\mult_97/n448 ) );
  AOI21X1 \mult_97/U287  ( .A(n406), .B(\mult_97/n543 ), .C(\mult_97/n538 ), 
        .Y(\mult_97/n536 ) );
  NAND2X1 \mult_97/U286  ( .A(n406), .B(\mult_97/n542 ), .Y(\mult_97/n535 ) );
  XOR2X1 \mult_97/U282  ( .A(\mult_97/n541 ), .B(\mult_97/n448 ), .Y(n641) );
  NAND2X1 \mult_97/U281  ( .A(\mult_97/n946 ), .B(\mult_97/n953 ), .Y(
        \mult_97/n531 ) );
  NOR2X1 \mult_97/U280  ( .A(\mult_97/n946 ), .B(\mult_97/n953 ), .Y(
        \mult_97/n530 ) );
  OAI21X1 \mult_97/U277  ( .A(n450), .B(\mult_97/n536 ), .C(n451), .Y(
        \mult_97/n529 ) );
  NOR2X1 \mult_97/U276  ( .A(n450), .B(\mult_97/n535 ), .Y(\mult_97/n528 ) );
  NAND2X1 \mult_97/U273  ( .A(\mult_97/n940 ), .B(\mult_97/n945 ), .Y(
        \mult_97/n526 ) );
  AOI21X1 \mult_97/U267  ( .A(n407), .B(\mult_97/n529 ), .C(\mult_97/n524 ), 
        .Y(\mult_97/n522 ) );
  NAND2X1 \mult_97/U266  ( .A(n407), .B(\mult_97/n528 ), .Y(\mult_97/n521 ) );
  OAI21X1 \mult_97/U265  ( .A(\mult_97/n521 ), .B(\mult_97/n580 ), .C(
        \mult_97/n522 ), .Y(\mult_97/n520 ) );
  NOR2X1 \mult_97/U264  ( .A(\mult_97/n521 ), .B(\mult_97/n579 ), .Y(
        \mult_97/n519 ) );
  NAND2X1 \mult_97/U261  ( .A(\mult_97/n934 ), .B(\mult_97/n939 ), .Y(
        \mult_97/n517 ) );
  NAND2X1 \mult_97/U251  ( .A(\mult_97/n930 ), .B(\mult_97/n933 ), .Y(
        \mult_97/n510 ) );
  AOI21X1 \mult_97/U245  ( .A(n409), .B(\mult_97/n511 ), .C(\mult_97/n508 ), 
        .Y(\mult_97/n506 ) );
  FAX1 \mult_97/U242  ( .A(n478), .B(n479), .C(\mult_97/n862 ), .YC(
        \mult_97/n505 ), .YS(n636) );
  FAX1 \mult_97/U241  ( .A(n476), .B(n477), .C(\mult_97/n505 ), .YC(
        \mult_97/n504 ), .YS(n635) );
  FAX1 \mult_97/U240  ( .A(\mult_97/n922 ), .B(n475), .C(\mult_97/n504 ), .YC(
        \mult_97/n503 ), .YS(n634) );
  FAX1 \mult_97/U239  ( .A(n446), .B(n410), .C(\mult_97/n503 ), .YC(
        \mult_97/n502 ), .YS(n633) );
  DFFPOSX1 clk_r_REG217_S2 ( .D(n32), .CLK(CLK), .Q(PRODUCT[0]) );
  DFFPOSX1 clk_r_REG215_S2 ( .D(n30), .CLK(CLK), .Q(PRODUCT[1]) );
  DFFPOSX1 clk_r_REG213_S2 ( .D(n28), .CLK(CLK), .Q(PRODUCT[2]) );
  DFFPOSX1 clk_r_REG211_S2 ( .D(n26), .CLK(CLK), .Q(PRODUCT[3]) );
  DFFPOSX1 clk_r_REG209_S2 ( .D(n24), .CLK(CLK), .Q(PRODUCT[4]) );
  DFFPOSX1 clk_r_REG207_S2 ( .D(n22), .CLK(CLK), .Q(PRODUCT[5]) );
  DFFPOSX1 clk_r_REG205_S2 ( .D(n20), .CLK(CLK), .Q(PRODUCT[6]) );
  DFFPOSX1 clk_r_REG203_S2 ( .D(n18), .CLK(CLK), .Q(PRODUCT[7]) );
  DFFPOSX1 clk_r_REG201_S2 ( .D(n16), .CLK(CLK), .Q(PRODUCT[8]) );
  DFFPOSX1 clk_r_REG198_S2 ( .D(n14), .CLK(CLK), .Q(PRODUCT[9]) );
  DFFPOSX1 clk_r_REG195_S2 ( .D(n12), .CLK(CLK), .Q(PRODUCT[10]) );
  DFFPOSX1 clk_r_REG192_S2 ( .D(n684), .CLK(CLK), .Q(PRODUCT[11]) );
  DFFPOSX1 clk_r_REG189_S2 ( .D(n683), .CLK(CLK), .Q(PRODUCT[12]) );
  DFFPOSX1 clk_r_REG186_S2 ( .D(n682), .CLK(CLK), .Q(PRODUCT[13]) );
  DFFPOSX1 clk_r_REG180_S2 ( .D(n680), .CLK(CLK), .Q(PRODUCT[15]) );
  DFFPOSX1 clk_r_REG183_S2 ( .D(n11), .CLK(CLK), .Q(PRODUCT[14]) );
  DFFPOSX1 clk_r_REG177_S2 ( .D(n679), .CLK(CLK), .Q(PRODUCT[16]) );
  DFFPOSX1 clk_r_REG216_S1 ( .D(n695), .CLK(CLK), .Q(n559) );
  DFFPOSX1 clk_r_REG174_S2 ( .D(n678), .CLK(CLK), .Q(PRODUCT[17]) );
  DFFPOSX1 clk_r_REG161_S2 ( .D(n675), .CLK(CLK), .Q(PRODUCT[20]) );
  DFFPOSX1 clk_r_REG171_S2 ( .D(n10), .CLK(CLK), .Q(PRODUCT[18]) );
  DFFPOSX1 clk_r_REG165_S2 ( .D(n676), .CLK(CLK), .Q(PRODUCT[19]) );
  DFFPOSX1 clk_r_REG159_S2 ( .D(n674), .CLK(CLK), .Q(PRODUCT[21]) );
  DFFPOSX1 clk_r_REG153_S2 ( .D(n673), .CLK(CLK), .Q(PRODUCT[22]) );
  DFFPOSX1 clk_r_REG147_S2 ( .D(n671), .CLK(CLK), .Q(PRODUCT[24]) );
  DFFPOSX1 clk_r_REG131_S2 ( .D(n667), .CLK(CLK), .Q(PRODUCT[28]) );
  DFFPOSX1 clk_r_REG150_S2 ( .D(n672), .CLK(CLK), .Q(PRODUCT[23]) );
  DFFPOSX1 clk_r_REG143_S2 ( .D(n670), .CLK(CLK), .Q(PRODUCT[25]) );
  DFFPOSX1 clk_r_REG138_S2 ( .D(n669), .CLK(CLK), .Q(PRODUCT[26]) );
  DFFPOSX1 \mult_97/clk_r_REG53_S1  ( .D(\mult_97/n921 ), .CLK(CLK), .Q(n446)
         );
  DFFPOSX1 clk_r_REG121_S2 ( .D(n666), .CLK(CLK), .Q(PRODUCT[29]) );
  DFFPOSX1 clk_r_REG118_S2 ( .D(n665), .CLK(CLK), .Q(PRODUCT[30]) );
  DFFPOSX1 clk_r_REG133_S2 ( .D(n668), .CLK(CLK), .Q(PRODUCT[27]) );
  DFFPOSX1 \mult_97/clk_r_REG105_S1  ( .D(\mult_97/n1867 ), .CLK(CLK), .Q(n410) );
  DFFPOSX1 clk_r_REG78_S2 ( .D(n663), .CLK(CLK), .Q(PRODUCT[32]) );
  DFFPOSX1 clk_r_REG83_S2 ( .D(n664), .CLK(CLK), .Q(PRODUCT[31]) );
  DFFPOSX1 clk_r_REG75_S2 ( .D(n662), .CLK(CLK), .Q(PRODUCT[33]) );
  DFFPOSX1 clk_r_REG29_S2 ( .D(n655), .CLK(CLK), .Q(PRODUCT[40]) );
  DFFPOSX1 clk_r_REG14_S2 ( .D(n9), .CLK(CLK), .Q(PRODUCT[58]) );
  DFFPOSX1 clk_r_REG72_S2 ( .D(n661), .CLK(CLK), .Q(PRODUCT[34]) );
  DFFPOSX1 clk_r_REG214_S1 ( .D(n694), .CLK(CLK), .Q(n561) );
  DFFPOSX1 clk_r_REG69_S2 ( .D(n659), .CLK(CLK), .Q(PRODUCT[36]) );
  DFFPOSX1 clk_r_REG67_S2 ( .D(n658), .CLK(CLK), .Q(PRODUCT[37]) );
  DFFPOSX1 \mult_97/clk_r_REG51_S1  ( .D(\mult_97/n923 ), .CLK(CLK), .Q(n475)
         );
  DFFPOSX1 clk_r_REG70_S2 ( .D(n660), .CLK(CLK), .Q(PRODUCT[35]) );
  DFFPOSX1 clk_r_REG13_S2 ( .D(n638), .CLK(CLK), .Q(PRODUCT[57]) );
  DFFPOSX1 clk_r_REG212_S1 ( .D(n693), .CLK(CLK), .Q(n563) );
  DFFPOSX1 clk_r_REG26_S2 ( .D(n654), .CLK(CLK), .Q(PRODUCT[41]) );
  DFFPOSX1 \mult_97/clk_r_REG52_S1  ( .D(\mult_97/n924 ), .CLK(CLK), .Q(n476)
         );
  DFFPOSX1 clk_r_REG21_S2 ( .D(n652), .CLK(CLK), .Q(PRODUCT[43]) );
  DFFPOSX1 clk_r_REG12_S2 ( .D(n8), .CLK(CLK), .Q(PRODUCT[50]) );
  DFFPOSX1 clk_r_REG20_S2 ( .D(n651), .CLK(CLK), .Q(PRODUCT[44]) );
  DFFPOSX1 clk_r_REG68_S2 ( .D(n657), .CLK(CLK), .Q(PRODUCT[38]) );
  DFFPOSX1 clk_r_REG23_S2 ( .D(n653), .CLK(CLK), .Q(PRODUCT[42]) );
  DFFPOSX1 clk_r_REG11_S2 ( .D(n646), .CLK(CLK), .Q(PRODUCT[49]) );
  DFFPOSX1 \mult_97/clk_r_REG49_S1  ( .D(\mult_97/n925 ), .CLK(CLK), .Q(n477)
         );
  DFFPOSX1 clk_r_REG19_S2 ( .D(n636), .CLK(CLK), .Q(PRODUCT[59]) );
  DFFPOSX1 clk_r_REG32_S2 ( .D(n656), .CLK(CLK), .Q(PRODUCT[39]) );
  DFFPOSX1 clk_r_REG6_S2 ( .D(n7), .CLK(CLK), .Q(PRODUCT[55]) );
  DFFPOSX1 clk_r_REG5_S2 ( .D(n639), .CLK(CLK), .Q(PRODUCT[56]) );
  DFFPOSX1 clk_r_REG7_S2 ( .D(n641), .CLK(CLK), .Q(PRODUCT[54]) );
  DFFPOSX1 \mult_97/clk_r_REG50_S1  ( .D(\mult_97/n926 ), .CLK(CLK), .Q(n478)
         );
  DFFPOSX1 clk_r_REG210_S1 ( .D(n692), .CLK(CLK), .Q(n565) );
  DFFPOSX1 clk_r_REG1_S2 ( .D(n650), .CLK(CLK), .Q(PRODUCT[45]) );
  DFFPOSX1 \mult_97/clk_r_REG48_S1  ( .D(\mult_97/n929 ), .CLK(CLK), .Q(n479)
         );
  DFFPOSX1 R_0 ( .D(n242), .CLK(CLK), .Q(\mult_97/n1671 ) );
  DFFPOSX1 R_1 ( .D(n241), .CLK(CLK), .Q(\mult_97/n1672 ) );
  DFFPOSX1 R_2 ( .D(n240), .CLK(CLK), .Q(\mult_97/n1651 ) );
  DFFPOSX1 R_3 ( .D(n239), .CLK(CLK), .Q(\mult_97/n1652 ) );
  DFFPOSX1 R_4 ( .D(n238), .CLK(CLK), .Q(\mult_97/n1631 ) );
  DFFPOSX1 R_5 ( .D(n237), .CLK(CLK), .Q(\mult_97/n1632 ) );
  DFFPOSX1 R_22 ( .D(n236), .CLK(CLK), .Q(\mult_97/n1403 ) );
  DFFPOSX1 R_23 ( .D(n235), .CLK(CLK), .Q(\mult_97/n1404 ) );
  DFFPOSX1 R_34 ( .D(n234), .CLK(CLK), .Q(\mult_97/n1235 ) );
  DFFPOSX1 R_35 ( .D(n233), .CLK(CLK), .Q(\mult_97/n1236 ) );
  DFFPOSX1 R_36 ( .D(n232), .CLK(CLK), .Q(\mult_97/n1211 ) );
  DFFPOSX1 R_37 ( .D(n231), .CLK(CLK), .Q(\mult_97/n1212 ) );
  DFFPOSX1 R_38 ( .D(n230), .CLK(CLK), .Q(\mult_97/n1187 ) );
  DFFPOSX1 R_39 ( .D(n229), .CLK(CLK), .Q(\mult_97/n1188 ) );
  DFFPOSX1 R_54 ( .D(n228), .CLK(CLK), .Q(\mult_97/n1019 ) );
  DFFPOSX1 R_55 ( .D(n227), .CLK(CLK), .Q(\mult_97/n1020 ) );
  DFFPOSX1 R_56 ( .D(n226), .CLK(CLK), .Q(n685) );
  OAI21X1 U1 ( .A(\mult_97/n825 ), .B(\mult_97/n828 ), .C(1'b1), .Y(n109) );
  OAI21X1 U2 ( .A(n470), .B(n468), .C(1'b1), .Y(n38) );
  OAI21X1 U3 ( .A(1'b0), .B(\mult_97/n868 ), .C(n454), .Y(n222) );
  OAI21X1 U4 ( .A(1'b0), .B(n404), .C(n472), .Y(n163) );
  OAI21X1 U5 ( .A(1'b0), .B(\mult_97/n905 ), .C(n466), .Y(n156) );
  OAI21X1 U6 ( .A(1'b0), .B(n556), .C(\mult_97/n725 ), .Y(n101) );
  OAI21X1 U7 ( .A(1'b0), .B(n408), .C(n448), .Y(n96) );
  OAI21X1 U8 ( .A(1'b0), .B(\mult_97/n519 ), .C(n408), .Y(n59) );
  OAI21X1 U9 ( .A(1'b0), .B(n404), .C(n403), .Y(n55) );
  OAI21X1 U10 ( .A(1'b0), .B(n407), .C(n449), .Y(n44) );
  BUFX2 U11 ( .A(n640), .Y(n7) );
  BUFX2 U12 ( .A(n645), .Y(n8) );
  BUFX2 U13 ( .A(n637), .Y(n9) );
  BUFX2 U14 ( .A(n677), .Y(n10) );
  BUFX2 U15 ( .A(n681), .Y(n11) );
  BUFX4 U16 ( .A(n685), .Y(n13) );
  BUFX2 U17 ( .A(n13), .Y(n12) );
  BUFX4 U18 ( .A(n577), .Y(n15) );
  BUFX2 U19 ( .A(n15), .Y(n14) );
  BUFX4 U20 ( .A(n575), .Y(n17) );
  BUFX2 U21 ( .A(n17), .Y(n16) );
  BUFX4 U22 ( .A(n573), .Y(n19) );
  BUFX2 U23 ( .A(n19), .Y(n18) );
  BUFX4 U24 ( .A(n571), .Y(n21) );
  BUFX2 U25 ( .A(n21), .Y(n20) );
  BUFX4 U26 ( .A(n569), .Y(n23) );
  BUFX2 U27 ( .A(n23), .Y(n22) );
  BUFX4 U28 ( .A(n567), .Y(n25) );
  BUFX2 U29 ( .A(n25), .Y(n24) );
  BUFX4 U30 ( .A(n565), .Y(n27) );
  BUFX2 U31 ( .A(n27), .Y(n26) );
  BUFX4 U32 ( .A(n563), .Y(n29) );
  BUFX2 U33 ( .A(n29), .Y(n28) );
  BUFX4 U34 ( .A(n561), .Y(n31) );
  BUFX2 U35 ( .A(n31), .Y(n30) );
  BUFX4 U36 ( .A(n559), .Y(n33) );
  BUFX2 U37 ( .A(n33), .Y(n32) );
  BUFX2 U38 ( .A(n643), .Y(n34) );
  INVX2 U39 ( .A(A[17]), .Y(n285) );
  INVX2 U40 ( .A(n551), .Y(n315) );
  INVX2 U41 ( .A(n552), .Y(n310) );
  INVX4 U42 ( .A(n535), .Y(n250) );
  INVX4 U43 ( .A(n317), .Y(n318) );
  INVX4 U44 ( .A(n548), .Y(n327) );
  INVX4 U45 ( .A(n322), .Y(n323) );
  INVX4 U46 ( .A(n537), .Y(n249) );
  INVX4 U47 ( .A(n545), .Y(n330) );
  INVX1 U48 ( .A(n533), .Y(n35) );
  OAI21X1 U49 ( .A(\mult_97/n740 ), .B(n35), .C(\mult_97/n737 ), .Y(n36) );
  INVX1 U50 ( .A(n36), .Y(\mult_97/n733 ) );
  OAI21X1 U52 ( .A(n468), .B(n471), .C(n469), .Y(n39) );
  AOI21X1 U53 ( .A(\mult_97/n809 ), .B(n38), .C(n39), .Y(\mult_97/n800 ) );
  NAND2X1 U54 ( .A(\mult_97/n876 ), .B(\mult_97/n605 ), .Y(n40) );
  NAND2X1 U55 ( .A(\mult_97/n606 ), .B(n40), .Y(n41) );
  OAI21X1 U56 ( .A(\mult_97/n606 ), .B(n40), .C(n41), .Y(n650) );
  AOI21X1 U57 ( .A(\mult_97/n528 ), .B(\mult_97/n575 ), .C(\mult_97/n529 ), 
        .Y(n42) );
  XOR2X1 U59 ( .A(n42), .B(n44), .Y(n639) );
  OAI21X1 U60 ( .A(\mult_97/n634 ), .B(\mult_97/n640 ), .C(\mult_97/n635 ), 
        .Y(n45) );
  NAND2X1 U61 ( .A(\mult_97/n632 ), .B(n530), .Y(n46) );
  NAND2X1 U62 ( .A(n45), .B(n46), .Y(n47) );
  OAI21X1 U63 ( .A(n45), .B(n46), .C(n47), .Y(n653) );
  INVX1 U64 ( .A(\mult_97/n685 ), .Y(n48) );
  INVX1 U65 ( .A(\mult_97/n887 ), .Y(n49) );
  OAI21X1 U66 ( .A(n48), .B(n49), .C(\mult_97/n684 ), .Y(n50) );
  INVX1 U67 ( .A(\mult_97/n678 ), .Y(n51) );
  NAND2X1 U68 ( .A(n51), .B(\mult_97/n679 ), .Y(n52) );
  NAND2X1 U69 ( .A(n50), .B(n52), .Y(n53) );
  OAI21X1 U70 ( .A(n50), .B(n52), .C(n53), .Y(n660) );
  INVX1 U72 ( .A(n472), .Y(n56) );
  AOI21X1 U73 ( .A(n404), .B(\mult_97/n818 ), .C(n56), .Y(n57) );
  OAI21X1 U74 ( .A(n474), .B(n55), .C(n57), .Y(\mult_97/n809 ) );
  INVX1 U76 ( .A(n448), .Y(n60) );
  AOI21X1 U77 ( .A(n408), .B(\mult_97/n520 ), .C(n60), .Y(n61) );
  OAI21X1 U78 ( .A(\mult_97/n646 ), .B(n59), .C(n61), .Y(\mult_97/n511 ) );
  INVX1 U79 ( .A(n450), .Y(n62) );
  INVX1 U80 ( .A(\mult_97/n575 ), .Y(n63) );
  OAI21X1 U81 ( .A(\mult_97/n535 ), .B(n63), .C(\mult_97/n536 ), .Y(n64) );
  NAND2X1 U82 ( .A(n62), .B(n451), .Y(n65) );
  NAND2X1 U83 ( .A(n64), .B(n65), .Y(n66) );
  OAI21X1 U84 ( .A(n64), .B(n65), .C(n66), .Y(n640) );
  OAI21X1 U85 ( .A(\mult_97/n617 ), .B(\mult_97/n624 ), .C(\mult_97/n618 ), 
        .Y(n67) );
  NAND2X1 U86 ( .A(\mult_97/n615 ), .B(n532), .Y(n68) );
  NAND2X1 U87 ( .A(n67), .B(n68), .Y(n69) );
  OAI21X1 U88 ( .A(n67), .B(n68), .C(n69), .Y(n651) );
  INVX1 U89 ( .A(\mult_97/n673 ), .Y(n70) );
  INVX1 U90 ( .A(\mult_97/n885 ), .Y(n71) );
  OAI21X1 U91 ( .A(n70), .B(n71), .C(\mult_97/n671 ), .Y(n72) );
  INVX1 U92 ( .A(\mult_97/n665 ), .Y(n73) );
  NAND2X1 U93 ( .A(n73), .B(\mult_97/n666 ), .Y(n74) );
  NAND2X1 U94 ( .A(n72), .B(n74), .Y(n75) );
  OAI21X1 U95 ( .A(n72), .B(n74), .C(n75), .Y(n658) );
  OAI21X1 U96 ( .A(\mult_97/n706 ), .B(\mult_97/n704 ), .C(\mult_97/n705 ), 
        .Y(n76) );
  INVX1 U97 ( .A(\mult_97/n701 ), .Y(n77) );
  NAND2X1 U98 ( .A(n77), .B(\mult_97/n702 ), .Y(n78) );
  NAND2X1 U99 ( .A(n76), .B(n78), .Y(n79) );
  OAI21X1 U100 ( .A(n76), .B(n78), .C(n79), .Y(n664) );
  OAI21X1 U101 ( .A(\mult_97/n756 ), .B(\mult_97/n754 ), .C(\mult_97/n755 ), 
        .Y(n80) );
  INVX1 U102 ( .A(\mult_97/n751 ), .Y(n81) );
  NAND2X1 U103 ( .A(n81), .B(\mult_97/n752 ), .Y(n82) );
  NAND2X1 U104 ( .A(n80), .B(n82), .Y(n83) );
  OAI21X1 U105 ( .A(n80), .B(n82), .C(n83), .Y(n672) );
  INVX1 U106 ( .A(\mult_97/n903 ), .Y(n84) );
  OAI21X1 U107 ( .A(n464), .B(n84), .C(n462), .Y(n85) );
  INVX1 U108 ( .A(n85), .Y(\mult_97/n774 ) );
  INVX1 U109 ( .A(\mult_97/n660 ), .Y(n86) );
  INVX1 U110 ( .A(\mult_97/n883 ), .Y(n87) );
  OAI21X1 U111 ( .A(n86), .B(n87), .C(\mult_97/n659 ), .Y(n88) );
  INVX1 U112 ( .A(\mult_97/n653 ), .Y(n89) );
  NAND2X1 U113 ( .A(n89), .B(\mult_97/n654 ), .Y(n90) );
  NAND2X1 U114 ( .A(n88), .B(n90), .Y(n91) );
  OAI21X1 U115 ( .A(n88), .B(n90), .C(n91), .Y(n656) );
  NAND2X1 U116 ( .A(\mult_97/n872 ), .B(\mult_97/n570 ), .Y(n92) );
  NAND2X1 U117 ( .A(\mult_97/n575 ), .B(n92), .Y(n93) );
  OAI21X1 U118 ( .A(\mult_97/n575 ), .B(n92), .C(n93), .Y(n646) );
  AOI21X1 U119 ( .A(\mult_97/n519 ), .B(\mult_97/n645 ), .C(\mult_97/n520 ), 
        .Y(n94) );
  XOR2X1 U121 ( .A(n94), .B(n96), .Y(n638) );
  NAND2X1 U122 ( .A(\mult_97/n887 ), .B(\mult_97/n684 ), .Y(n97) );
  NAND2X1 U123 ( .A(\mult_97/n685 ), .B(n97), .Y(n98) );
  OAI21X1 U124 ( .A(\mult_97/n685 ), .B(n97), .C(n98), .Y(n661) );
  AOI21X1 U125 ( .A(n531), .B(\mult_97/n731 ), .C(\mult_97/n728 ), .Y(n99) );
  XOR2X1 U127 ( .A(n99), .B(n101), .Y(n668) );
  INVX1 U128 ( .A(\mult_97/n705 ), .Y(n102) );
  NOR2X1 U129 ( .A(n102), .B(\mult_97/n704 ), .Y(n103) );
  NAND2X1 U130 ( .A(\mult_97/n706 ), .B(n103), .Y(n104) );
  OAI21X1 U131 ( .A(n103), .B(\mult_97/n706 ), .C(n104), .Y(n665) );
  INVX1 U132 ( .A(\mult_97/n755 ), .Y(n105) );
  NOR2X1 U133 ( .A(n105), .B(\mult_97/n754 ), .Y(n106) );
  NAND2X1 U134 ( .A(\mult_97/n756 ), .B(n106), .Y(n107) );
  OAI21X1 U135 ( .A(n106), .B(\mult_97/n756 ), .C(n107), .Y(n673) );
  OAI21X1 U137 ( .A(\mult_97/n825 ), .B(\mult_97/n829 ), .C(\mult_97/n826 ), 
        .Y(n110) );
  AOI21X1 U138 ( .A(\mult_97/n831 ), .B(n109), .C(n110), .Y(\mult_97/n822 ) );
  INVX1 U139 ( .A(\mult_97/n841 ), .Y(n111) );
  NOR2X1 U140 ( .A(n111), .B(\mult_97/n840 ), .Y(n112) );
  NAND2X1 U141 ( .A(\mult_97/n842 ), .B(n112), .Y(n113) );
  OAI21X1 U142 ( .A(n112), .B(\mult_97/n842 ), .C(n113), .Y(n689) );
  INVX1 U143 ( .A(\mult_97/n606 ), .Y(n114) );
  INVX1 U144 ( .A(\mult_97/n876 ), .Y(n115) );
  OAI21X1 U145 ( .A(n114), .B(n115), .C(\mult_97/n605 ), .Y(n116) );
  INVX1 U146 ( .A(\mult_97/n599 ), .Y(n117) );
  NAND2X1 U147 ( .A(n117), .B(\mult_97/n600 ), .Y(n118) );
  NAND2X1 U148 ( .A(n116), .B(n118), .Y(n119) );
  OAI21X1 U149 ( .A(n116), .B(n118), .C(n119), .Y(n649) );
  INVX1 U150 ( .A(n457), .Y(n120) );
  NAND2X1 U151 ( .A(n120), .B(n458), .Y(n121) );
  NAND2X1 U152 ( .A(\mult_97/n558 ), .B(n121), .Y(n122) );
  OAI21X1 U153 ( .A(\mult_97/n558 ), .B(n121), .C(n122), .Y(n644) );
  OAI21X1 U154 ( .A(A[0]), .B(n307), .C(n309), .Y(n123) );
  AOI21X1 U155 ( .A(A[0]), .B(n307), .C(n123), .Y(n553) );
  INVX1 U156 ( .A(\mult_97/n853 ), .Y(n124) );
  NOR2X1 U157 ( .A(n124), .B(\mult_97/n852 ), .Y(n125) );
  NAND2X1 U158 ( .A(\mult_97/n854 ), .B(n125), .Y(n126) );
  OAI21X1 U159 ( .A(n125), .B(\mult_97/n854 ), .C(n126), .Y(n692) );
  NAND2X1 U160 ( .A(\mult_97/n878 ), .B(\mult_97/n618 ), .Y(n127) );
  NAND2X1 U161 ( .A(\mult_97/n623 ), .B(n127), .Y(n128) );
  OAI21X1 U162 ( .A(\mult_97/n623 ), .B(n127), .C(n128), .Y(n652) );
  OAI21X1 U163 ( .A(\mult_97/n2378 ), .B(\mult_97/n1866 ), .C(\mult_97/n861 ), 
        .Y(n129) );
  INVX1 U164 ( .A(n129), .Y(n694) );
  NAND2X1 U165 ( .A(\mult_97/n881 ), .B(\mult_97/n644 ), .Y(n130) );
  NAND2X1 U166 ( .A(\mult_97/n645 ), .B(n130), .Y(n131) );
  OAI21X1 U167 ( .A(\mult_97/n645 ), .B(n130), .C(n131), .Y(n655) );
  OAI21X1 U168 ( .A(\mult_97/n695 ), .B(\mult_97/n693 ), .C(\mult_97/n694 ), 
        .Y(n132) );
  INVX1 U169 ( .A(\mult_97/n690 ), .Y(n133) );
  NAND2X1 U170 ( .A(n133), .B(\mult_97/n691 ), .Y(n134) );
  NAND2X1 U171 ( .A(n132), .B(n134), .Y(n135) );
  OAI21X1 U172 ( .A(n132), .B(n134), .C(n135), .Y(n662) );
  INVX1 U173 ( .A(\mult_97/n716 ), .Y(n136) );
  INVX1 U174 ( .A(\mult_97/n893 ), .Y(n137) );
  OAI21X1 U175 ( .A(n136), .B(n137), .C(\mult_97/n715 ), .Y(n138) );
  INVX1 U176 ( .A(\mult_97/n709 ), .Y(n139) );
  NAND2X1 U177 ( .A(n139), .B(\mult_97/n710 ), .Y(n140) );
  NAND2X1 U178 ( .A(n138), .B(n140), .Y(n141) );
  OAI21X1 U179 ( .A(n138), .B(n140), .C(n141), .Y(n666) );
  NAND2X1 U180 ( .A(n531), .B(\mult_97/n730 ), .Y(n142) );
  NAND2X1 U181 ( .A(\mult_97/n731 ), .B(n142), .Y(n143) );
  OAI21X1 U182 ( .A(\mult_97/n731 ), .B(n142), .C(n143), .Y(n669) );
  INVX1 U183 ( .A(\mult_97/n766 ), .Y(n144) );
  INVX1 U184 ( .A(\mult_97/n901 ), .Y(n145) );
  OAI21X1 U185 ( .A(n144), .B(n145), .C(\mult_97/n765 ), .Y(n146) );
  INVX1 U186 ( .A(\mult_97/n759 ), .Y(n147) );
  NAND2X1 U187 ( .A(n147), .B(\mult_97/n760 ), .Y(n148) );
  NAND2X1 U188 ( .A(n146), .B(n148), .Y(n149) );
  OAI21X1 U189 ( .A(n146), .B(n148), .C(n149), .Y(n674) );
  OAI21X1 U190 ( .A(\mult_97/n786 ), .B(\mult_97/n773 ), .C(\mult_97/n774 ), 
        .Y(n150) );
  INVX1 U191 ( .A(\mult_97/n770 ), .Y(n151) );
  NAND2X1 U192 ( .A(n151), .B(\mult_97/n771 ), .Y(n152) );
  NAND2X1 U193 ( .A(n150), .B(n152), .Y(n153) );
  OAI21X1 U194 ( .A(n150), .B(n152), .C(n153), .Y(n676) );
  AOI21X1 U195 ( .A(n405), .B(\mult_97/n799 ), .C(\mult_97/n796 ), .Y(n154) );
  XOR2X1 U197 ( .A(n154), .B(n156), .Y(n679) );
  OAI21X1 U198 ( .A(\mult_97/n808 ), .B(n470), .C(n471), .Y(n157) );
  INVX1 U199 ( .A(n468), .Y(n158) );
  NAND2X1 U200 ( .A(n158), .B(n469), .Y(n159) );
  NAND2X1 U201 ( .A(n157), .B(n159), .Y(n160) );
  OAI21X1 U202 ( .A(n157), .B(n159), .C(n160), .Y(n681) );
  AOI21X1 U203 ( .A(n403), .B(\mult_97/n821 ), .C(\mult_97/n818 ), .Y(n161) );
  XOR2X1 U205 ( .A(n161), .B(n163), .Y(n683) );
  INVX1 U206 ( .A(\mult_97/n845 ), .Y(n164) );
  NOR2X1 U207 ( .A(n164), .B(\mult_97/n844 ), .Y(n165) );
  NAND2X1 U208 ( .A(\mult_97/n846 ), .B(n165), .Y(n166) );
  OAI21X1 U209 ( .A(n165), .B(\mult_97/n846 ), .C(n166), .Y(n690) );
  INVX1 U210 ( .A(\mult_97/n833 ), .Y(n167) );
  NOR2X1 U211 ( .A(n167), .B(\mult_97/n832 ), .Y(n168) );
  NAND2X1 U212 ( .A(\mult_97/n834 ), .B(n168), .Y(n169) );
  OAI21X1 U213 ( .A(n168), .B(\mult_97/n834 ), .C(n169), .Y(n687) );
  NAND2X1 U214 ( .A(\mult_97/n874 ), .B(\mult_97/n593 ), .Y(n170) );
  NAND2X1 U215 ( .A(\mult_97/n594 ), .B(n170), .Y(n171) );
  OAI21X1 U216 ( .A(\mult_97/n594 ), .B(n170), .C(n171), .Y(n648) );
  OAI21X1 U217 ( .A(\mult_97/n559 ), .B(n457), .C(n458), .Y(n172) );
  INVX1 U218 ( .A(n455), .Y(n173) );
  NAND2X1 U219 ( .A(n173), .B(n456), .Y(n174) );
  NAND2X1 U220 ( .A(n172), .B(n174), .Y(n175) );
  OAI21X1 U221 ( .A(n172), .B(n174), .C(n175), .Y(n643) );
  NAND2X1 U222 ( .A(\mult_97/n883 ), .B(\mult_97/n659 ), .Y(n176) );
  NAND2X1 U223 ( .A(\mult_97/n660 ), .B(n176), .Y(n177) );
  OAI21X1 U224 ( .A(\mult_97/n660 ), .B(n176), .C(n177), .Y(n657) );
  OAI21X1 U225 ( .A(\mult_97/n569 ), .B(\mult_97/n576 ), .C(\mult_97/n570 ), 
        .Y(n178) );
  NAND2X1 U226 ( .A(n460), .B(\mult_97/n871 ), .Y(n179) );
  NAND2X1 U227 ( .A(n178), .B(n179), .Y(n180) );
  OAI21X1 U228 ( .A(n178), .B(n179), .C(n180), .Y(n645) );
  NAND2X1 U229 ( .A(\mult_97/n858 ), .B(n529), .Y(n181) );
  NAND2X1 U230 ( .A(\mult_97/n859 ), .B(n181), .Y(n182) );
  OAI21X1 U231 ( .A(\mult_97/n859 ), .B(n181), .C(n182), .Y(n693) );
  NAND2X1 U232 ( .A(n409), .B(n447), .Y(n183) );
  NAND2X1 U233 ( .A(\mult_97/n511 ), .B(n183), .Y(n184) );
  OAI21X1 U234 ( .A(\mult_97/n511 ), .B(n183), .C(n184), .Y(n637) );
  INVX1 U235 ( .A(\mult_97/n694 ), .Y(n185) );
  NOR2X1 U236 ( .A(n185), .B(\mult_97/n693 ), .Y(n186) );
  NAND2X1 U237 ( .A(\mult_97/n695 ), .B(n186), .Y(n187) );
  OAI21X1 U238 ( .A(n186), .B(\mult_97/n695 ), .C(n187), .Y(n663) );
  OAI21X1 U239 ( .A(\mult_97/n739 ), .B(\mult_97/n745 ), .C(\mult_97/n740 ), 
        .Y(n188) );
  NAND2X1 U240 ( .A(\mult_97/n737 ), .B(n533), .Y(n189) );
  NAND2X1 U241 ( .A(n188), .B(n189), .Y(n190) );
  OAI21X1 U242 ( .A(n188), .B(n189), .C(n190), .Y(n670) );
  NAND2X1 U243 ( .A(\mult_97/n893 ), .B(\mult_97/n715 ), .Y(n191) );
  NAND2X1 U244 ( .A(\mult_97/n716 ), .B(n191), .Y(n192) );
  OAI21X1 U245 ( .A(\mult_97/n716 ), .B(n191), .C(n192), .Y(n667) );
  OAI21X1 U246 ( .A(n463), .B(\mult_97/n786 ), .C(n464), .Y(n193) );
  NAND2X1 U247 ( .A(n462), .B(\mult_97/n903 ), .Y(n194) );
  NAND2X1 U248 ( .A(n193), .B(n194), .Y(n195) );
  OAI21X1 U249 ( .A(n193), .B(n194), .C(n195), .Y(n677) );
  NAND2X1 U250 ( .A(\mult_97/n901 ), .B(\mult_97/n765 ), .Y(n196) );
  NAND2X1 U251 ( .A(\mult_97/n766 ), .B(n196), .Y(n197) );
  OAI21X1 U252 ( .A(\mult_97/n766 ), .B(n196), .C(n197), .Y(n675) );
  NAND2X1 U253 ( .A(n405), .B(n467), .Y(n198) );
  NAND2X1 U254 ( .A(\mult_97/n799 ), .B(n198), .Y(n199) );
  OAI21X1 U255 ( .A(\mult_97/n799 ), .B(n198), .C(n199), .Y(n680) );
  INVX1 U256 ( .A(n471), .Y(n200) );
  NOR2X1 U257 ( .A(n200), .B(n470), .Y(n201) );
  NAND2X1 U258 ( .A(\mult_97/n808 ), .B(n201), .Y(n202) );
  OAI21X1 U259 ( .A(n201), .B(\mult_97/n808 ), .C(n202), .Y(n682) );
  NAND2X1 U260 ( .A(n403), .B(n473), .Y(n203) );
  NAND2X1 U261 ( .A(\mult_97/n821 ), .B(n203), .Y(n204) );
  OAI21X1 U262 ( .A(\mult_97/n821 ), .B(n203), .C(n204), .Y(n684) );
  NAND2X1 U263 ( .A(\mult_97/n850 ), .B(n528), .Y(n205) );
  NAND2X1 U264 ( .A(\mult_97/n851 ), .B(n205), .Y(n206) );
  OAI21X1 U265 ( .A(\mult_97/n851 ), .B(n205), .C(n206), .Y(n691) );
  INVX1 U266 ( .A(\mult_97/n837 ), .Y(n207) );
  OAI21X1 U267 ( .A(\mult_97/n840 ), .B(\mult_97/n842 ), .C(\mult_97/n841 ), 
        .Y(n208) );
  NAND2X1 U268 ( .A(n207), .B(\mult_97/n838 ), .Y(n209) );
  NAND2X1 U269 ( .A(n208), .B(n209), .Y(n210) );
  OAI21X1 U270 ( .A(n208), .B(n209), .C(n210), .Y(n688) );
  INVX1 U271 ( .A(\mult_97/n829 ), .Y(n211) );
  NOR2X1 U272 ( .A(n211), .B(\mult_97/n828 ), .Y(n212) );
  NAND2X1 U273 ( .A(\mult_97/n830 ), .B(n212), .Y(n213) );
  OAI21X1 U274 ( .A(n212), .B(\mult_97/n830 ), .C(n213), .Y(n686) );
  INVX1 U275 ( .A(\mult_97/n587 ), .Y(n214) );
  INVX1 U276 ( .A(\mult_97/n594 ), .Y(n215) );
  INVX1 U277 ( .A(\mult_97/n874 ), .Y(n216) );
  OAI21X1 U278 ( .A(n215), .B(n216), .C(\mult_97/n593 ), .Y(n217) );
  NAND2X1 U279 ( .A(n214), .B(\mult_97/n588 ), .Y(n218) );
  NAND2X1 U280 ( .A(n217), .B(n218), .Y(n219) );
  OAI21X1 U281 ( .A(n217), .B(n218), .C(n219), .Y(n647) );
  AOI21X1 U282 ( .A(\mult_97/n551 ), .B(\mult_97/n558 ), .C(\mult_97/n552 ), 
        .Y(n220) );
  XOR2X1 U284 ( .A(n220), .B(n222), .Y(n642) );
  INVX4 U285 ( .A(A[15]), .Y(n288) );
  INVX8 U286 ( .A(n288), .Y(n289) );
  INVX8 U287 ( .A(n224), .Y(n335) );
  INVX8 U288 ( .A(n225), .Y(n334) );
  AND2X2 U289 ( .A(\mult_97/n362 ), .B(\mult_97/n2949 ), .Y(n223) );
  INVX8 U290 ( .A(n540), .Y(n338) );
  INVX8 U291 ( .A(n541), .Y(n337) );
  INVX8 U292 ( .A(n536), .Y(n336) );
  INVX8 U293 ( .A(n557), .Y(n332) );
  INVX8 U294 ( .A(n542), .Y(n333) );
  AND2X2 U295 ( .A(\mult_97/n371 ), .B(\mult_97/n2946 ), .Y(n224) );
  AND2X2 U296 ( .A(\mult_97/n368 ), .B(\mult_97/n2947 ), .Y(n225) );
  OR2X1 U297 ( .A(\mult_97/n1767 ), .B(\mult_97/n1754 ), .Y(n523) );
  OR2X1 U298 ( .A(\mult_97/n961 ), .B(\mult_97/n954 ), .Y(n524) );
  OR2X1 U299 ( .A(\mult_97/n1801 ), .B(\mult_97/n1792 ), .Y(n522) );
  OR2X1 U300 ( .A(\mult_97/n1811 ), .B(\mult_97/n1802 ), .Y(n521) );
  OR2X1 U301 ( .A(\mult_97/n940 ), .B(\mult_97/n945 ), .Y(n525) );
  OR2X1 U302 ( .A(\mult_97/n930 ), .B(\mult_97/n933 ), .Y(n526) );
  OR2X1 U303 ( .A(\mult_97/n934 ), .B(\mult_97/n939 ), .Y(n527) );
  INVX1 U304 ( .A(\mult_97/n850 ), .Y(\mult_97/n848 ) );
  INVX2 U305 ( .A(\mult_97/n717 ), .Y(\mult_97/n716 ) );
  INVX1 U306 ( .A(\mult_97/n858 ), .Y(\mult_97/n856 ) );
  INVX2 U307 ( .A(\mult_97/n746 ), .Y(\mult_97/n745 ) );
  INVX1 U308 ( .A(n252), .Y(\mult_97/n1867 ) );
  INVX8 U309 ( .A(n223), .Y(n243) );
  INVX8 U310 ( .A(n543), .Y(n244) );
  INVX4 U311 ( .A(n320), .Y(n321) );
  INVX4 U312 ( .A(n324), .Y(n325) );
  INVX1 U313 ( .A(\mult_97/n610 ), .Y(\mult_97/n608 ) );
  INVX1 U314 ( .A(\mult_97/n611 ), .Y(\mult_97/n609 ) );
  INVX4 U315 ( .A(n312), .Y(n313) );
  INVX1 U316 ( .A(\mult_97/n644 ), .Y(\mult_97/n642 ) );
  INVX8 U317 ( .A(n554), .Y(n245) );
  INVX8 U318 ( .A(n553), .Y(n246) );
  INVX1 U319 ( .A(\mult_97/n635 ), .Y(\mult_97/n637 ) );
  INVX1 U320 ( .A(\mult_97/n598 ), .Y(\mult_97/n596 ) );
  INVX8 U321 ( .A(n539), .Y(n247) );
  INVX8 U322 ( .A(n538), .Y(n248) );
  INVX1 U323 ( .A(\mult_97/n2874 ), .Y(n267) );
  INVX1 U324 ( .A(\mult_97/n632 ), .Y(\mult_97/n630 ) );
  INVX1 U325 ( .A(\mult_97/n618 ), .Y(\mult_97/n620 ) );
  INVX1 U326 ( .A(\mult_97/n615 ), .Y(\mult_97/n613 ) );
  INVX1 U327 ( .A(\mult_97/n725 ), .Y(\mult_97/n723 ) );
  INVX1 U328 ( .A(\mult_97/n730 ), .Y(\mult_97/n728 ) );
  INVX1 U329 ( .A(\mult_97/n570 ), .Y(\mult_97/n572 ) );
  INVX1 U330 ( .A(\mult_97/n604 ), .Y(\mult_97/n876 ) );
  INVX1 U331 ( .A(\mult_97/n714 ), .Y(\mult_97/n893 ) );
  INVX1 U332 ( .A(\mult_97/n764 ), .Y(\mult_97/n901 ) );
  INVX4 U333 ( .A(n544), .Y(n331) );
  INVX2 U334 ( .A(n453), .Y(\mult_97/n868 ) );
  INVX2 U335 ( .A(n459), .Y(\mult_97/n871 ) );
  INVX2 U336 ( .A(n446), .Y(\mult_97/n922 ) );
  INVX2 U337 ( .A(n473), .Y(\mult_97/n818 ) );
  INVX2 U338 ( .A(n467), .Y(\mult_97/n796 ) );
  INVX2 U339 ( .A(n465), .Y(\mult_97/n905 ) );
  INVX2 U340 ( .A(n463), .Y(\mult_97/n904 ) );
  INVX4 U341 ( .A(n402), .Y(n251) );
  INVX2 U342 ( .A(A[9]), .Y(n295) );
  INVX2 U343 ( .A(A[7]), .Y(n298) );
  INVX2 U344 ( .A(A[5]), .Y(n301) );
  INVX2 U345 ( .A(n474), .Y(\mult_97/n821 ) );
  INVX2 U346 ( .A(\A_extended[32] ), .Y(n268) );
  INVX2 U347 ( .A(n461), .Y(\mult_97/n903 ) );
  AOI21X1 U348 ( .A(n331), .B(n339), .C(\mult_97/n2379 ), .Y(n252) );
  NOR2X1 U349 ( .A(n402), .B(n331), .Y(\mult_97/n1898 ) );
  AOI21X1 U350 ( .A(n330), .B(n248), .C(\mult_97/n2412 ), .Y(n253) );
  NOR2X1 U351 ( .A(n402), .B(n330), .Y(\mult_97/n1929 ) );
  AOI21X1 U352 ( .A(n329), .B(n338), .C(\mult_97/n2445 ), .Y(n254) );
  NOR2X1 U353 ( .A(n402), .B(n329), .Y(\mult_97/n1962 ) );
  AOI21X1 U354 ( .A(n328), .B(n250), .C(\mult_97/n2478 ), .Y(n255) );
  NOR2X1 U355 ( .A(n402), .B(n328), .Y(\mult_97/n1989 ) );
  AOI21X1 U356 ( .A(n327), .B(n247), .C(\mult_97/n2511 ), .Y(n256) );
  NOR2X1 U357 ( .A(n402), .B(n327), .Y(\mult_97/n2022 ) );
  AOI21X1 U358 ( .A(n326), .B(n337), .C(\mult_97/n2544 ), .Y(n257) );
  NOR2X1 U359 ( .A(n402), .B(n326), .Y(\mult_97/n2055 ) );
  AOI21X1 U360 ( .A(\mult_97/n374 ), .B(n336), .C(\mult_97/n2577 ), .Y(n258)
         );
  NOR2X1 U361 ( .A(n402), .B(\mult_97/n374 ), .Y(\mult_97/n2086 ) );
  AOI21X1 U362 ( .A(n323), .B(n335), .C(\mult_97/n2610 ), .Y(n259) );
  NOR2X1 U363 ( .A(n402), .B(n323), .Y(\mult_97/n2119 ) );
  AOI21X1 U364 ( .A(\mult_97/n368 ), .B(n334), .C(\mult_97/n2643 ), .Y(n260)
         );
  NOR2X1 U365 ( .A(n402), .B(\mult_97/n368 ), .Y(\mult_97/n2152 ) );
  AOI21X1 U366 ( .A(n319), .B(n249), .C(\mult_97/n2676 ), .Y(n261) );
  NOR2X1 U367 ( .A(n402), .B(n319), .Y(\mult_97/n2183 ) );
  AOI21X1 U368 ( .A(n318), .B(n243), .C(\mult_97/n2709 ), .Y(n262) );
  NOR2X1 U369 ( .A(n402), .B(\mult_97/n362 ), .Y(\mult_97/n2216 ) );
  AOI21X1 U370 ( .A(n315), .B(n333), .C(\mult_97/n2742 ), .Y(n263) );
  NOR2X1 U371 ( .A(n402), .B(n315), .Y(\mult_97/n2249 ) );
  AOI21X1 U372 ( .A(n314), .B(n245), .C(\mult_97/n2775 ), .Y(n264) );
  NOR2X1 U373 ( .A(n402), .B(n314), .Y(\mult_97/n2280 ) );
  AOI21X1 U374 ( .A(n313), .B(n332), .C(\mult_97/n2808 ), .Y(n265) );
  NOR2X1 U375 ( .A(n402), .B(\mult_97/n353 ), .Y(\mult_97/n2313 ) );
  AOI21X1 U376 ( .A(n310), .B(n244), .C(\mult_97/n2841 ), .Y(n266) );
  NOR2X1 U377 ( .A(n402), .B(n310), .Y(\mult_97/n2346 ) );
  OAI21X1 U378 ( .A(A[0]), .B(n553), .C(n267), .Y(\mult_97/n2347 ) );
  NAND2X1 U379 ( .A(n270), .B(n402), .Y(\mult_97/n2411 ) );
  NAND2X1 U380 ( .A(n272), .B(n402), .Y(\mult_97/n2444 ) );
  NAND2X1 U381 ( .A(n274), .B(n402), .Y(\mult_97/n2477 ) );
  NAND2X1 U382 ( .A(n276), .B(n402), .Y(\mult_97/n2510 ) );
  NAND2X1 U383 ( .A(n279), .B(n402), .Y(\mult_97/n2543 ) );
  NAND2X1 U384 ( .A(n281), .B(n402), .Y(\mult_97/n2576 ) );
  NAND2X1 U385 ( .A(n283), .B(n402), .Y(\mult_97/n2609 ) );
  NAND2X1 U386 ( .A(n286), .B(n402), .Y(\mult_97/n2642 ) );
  NAND2X1 U387 ( .A(n289), .B(n402), .Y(\mult_97/n2675 ) );
  NAND2X1 U388 ( .A(n291), .B(n402), .Y(\mult_97/n2708 ) );
  NAND2X1 U389 ( .A(n294), .B(n402), .Y(\mult_97/n2741 ) );
  NAND2X1 U390 ( .A(n296), .B(n402), .Y(\mult_97/n2774 ) );
  NAND2X1 U391 ( .A(n299), .B(n402), .Y(\mult_97/n2807 ) );
  NAND2X1 U392 ( .A(n302), .B(n402), .Y(\mult_97/n2840 ) );
  NAND2X1 U393 ( .A(n304), .B(n402), .Y(\mult_97/n2873 ) );
  NAND2X1 U394 ( .A(n307), .B(n402), .Y(\mult_97/n2906 ) );
  INVX2 U395 ( .A(\mult_97/n576 ), .Y(\mult_97/n575 ) );
  INVX2 U396 ( .A(\mult_97/n646 ), .Y(\mult_97/n645 ) );
  INVX2 U397 ( .A(\mult_97/n767 ), .Y(\mult_97/n766 ) );
  INVX2 U398 ( .A(\mult_97/n787 ), .Y(\mult_97/n786 ) );
  NOR2X1 U399 ( .A(n402), .B(n309), .Y(n695) );
  INVX8 U400 ( .A(n273), .Y(n274) );
  INVX8 U401 ( .A(n275), .Y(n277) );
  INVX8 U402 ( .A(n280), .Y(n281) );
  INVX8 U403 ( .A(n282), .Y(n284) );
  INVX8 U404 ( .A(n285), .Y(n287) );
  INVX8 U405 ( .A(n290), .Y(n292) );
  INVX8 U406 ( .A(n295), .Y(n297) );
  INVX8 U407 ( .A(n298), .Y(n300) );
  INVX8 U408 ( .A(n303), .Y(n305) );
  INVX8 U409 ( .A(n306), .Y(n307) );
  INVX8 U410 ( .A(n306), .Y(n308) );
  INVX1 U411 ( .A(\mult_97/n502 ), .Y(n632) );
  OR2X2 U412 ( .A(\mult_97/n1849 ), .B(\mult_97/n1848 ), .Y(n528) );
  OR2X2 U413 ( .A(\mult_97/n2377 ), .B(\mult_97/n2346 ), .Y(n529) );
  OR2X2 U414 ( .A(\mult_97/n1122 ), .B(\mult_97/n1141 ), .Y(n530) );
  OR2X2 U415 ( .A(\mult_97/n1563 ), .B(\mult_97/n1540 ), .Y(n531) );
  OR2X2 U416 ( .A(\mult_97/n1101 ), .B(\mult_97/n1084 ), .Y(n532) );
  OR2X2 U417 ( .A(\mult_97/n1587 ), .B(\mult_97/n1564 ), .Y(n533) );
  INVX2 U418 ( .A(\mult_97/n371 ), .Y(n322) );
  INVX2 U419 ( .A(\mult_97/n362 ), .Y(n317) );
  INVX2 U420 ( .A(\mult_97/n374 ), .Y(n324) );
  AND2X2 U421 ( .A(\mult_97/n2939 ), .B(n331), .Y(n534) );
  AND2X2 U422 ( .A(\mult_97/n2942 ), .B(n328), .Y(n535) );
  AND2X2 U423 ( .A(\mult_97/n2945 ), .B(\mult_97/n374 ), .Y(n536) );
  AND2X2 U424 ( .A(\mult_97/n2948 ), .B(n319), .Y(n537) );
  AND2X2 U425 ( .A(n330), .B(\mult_97/n2940 ), .Y(n538) );
  AND2X2 U426 ( .A(n327), .B(\mult_97/n2943 ), .Y(n539) );
  AND2X2 U427 ( .A(n329), .B(\mult_97/n2941 ), .Y(n540) );
  AND2X2 U428 ( .A(n326), .B(\mult_97/n2944 ), .Y(n541) );
  AND2X2 U429 ( .A(n315), .B(\mult_97/n2950 ), .Y(n542) );
  AND2X2 U430 ( .A(n310), .B(\mult_97/n2953 ), .Y(n543) );
  XOR2X1 U431 ( .A(A[29]), .B(A[30]), .Y(n544) );
  XOR2X1 U432 ( .A(A[28]), .B(A[27]), .Y(n545) );
  XOR2X1 U433 ( .A(A[26]), .B(n277), .Y(n546) );
  XOR2X1 U434 ( .A(A[23]), .B(A[24]), .Y(n547) );
  XOR2X1 U435 ( .A(A[22]), .B(A[21]), .Y(n548) );
  XOR2X1 U436 ( .A(A[20]), .B(n284), .Y(n549) );
  XOR2X1 U437 ( .A(A[11]), .B(A[12]), .Y(n550) );
  XOR2X1 U438 ( .A(A[8]), .B(n300), .Y(n551) );
  XOR2X1 U439 ( .A(A[2]), .B(n308), .Y(n552) );
  AND2X2 U440 ( .A(\mult_97/n2951 ), .B(n314), .Y(n554) );
  XOR2X1 U441 ( .A(A[5]), .B(A[6]), .Y(n555) );
  OR2X2 U442 ( .A(\mult_97/n1539 ), .B(\mult_97/n1514 ), .Y(n556) );
  INVX2 U443 ( .A(\mult_97/n353 ), .Y(n312) );
  INVX2 U444 ( .A(\mult_97/n368 ), .Y(n320) );
  AND2X2 U445 ( .A(\mult_97/n353 ), .B(\mult_97/n2952 ), .Y(n557) );
  INVX8 U446 ( .A(n275), .Y(n276) );
  INVX8 U447 ( .A(n271), .Y(n272) );
  INVX1 U448 ( .A(\mult_97/n825 ), .Y(\mult_97/n911 ) );
  INVX1 U449 ( .A(n466), .Y(\mult_97/n791 ) );
  INVX1 U450 ( .A(n460), .Y(\mult_97/n565 ) );
  INVX1 U451 ( .A(n454), .Y(\mult_97/n547 ) );
  INVX1 U452 ( .A(n452), .Y(\mult_97/n538 ) );
  INVX1 U453 ( .A(n449), .Y(\mult_97/n524 ) );
  INVX1 U454 ( .A(n447), .Y(\mult_97/n508 ) );
  INVX1 U455 ( .A(\mult_97/n562 ), .Y(\mult_97/n560 ) );
  INVX1 U456 ( .A(\mult_97/n579 ), .Y(\mult_97/n577 ) );
  INVX1 U457 ( .A(\mult_97/n580 ), .Y(\mult_97/n578 ) );
  INVX1 U458 ( .A(\mult_97/n563 ), .Y(\mult_97/n561 ) );
  INVX1 U459 ( .A(\mult_97/n663 ), .Y(\mult_97/n661 ) );
  INVX1 U460 ( .A(\mult_97/n688 ), .Y(\mult_97/n686 ) );
  INVX4 U461 ( .A(A[1]), .Y(n306) );
  INVX4 U462 ( .A(A[13]), .Y(n290) );
  INVX8 U463 ( .A(n550), .Y(n319) );
  INVX4 U464 ( .A(A[25]), .Y(n275) );
  INVX8 U465 ( .A(n547), .Y(n328) );
  INVX8 U466 ( .A(n549), .Y(n326) );
  INVX8 U467 ( .A(n293), .Y(n294) );
  INVX8 U468 ( .A(n555), .Y(n314) );
  INVX2 U469 ( .A(A[23]), .Y(n278) );
  INVX8 U470 ( .A(n278), .Y(n279) );
  INVX2 U471 ( .A(A[27]), .Y(n273) );
  INVX8 U472 ( .A(n546), .Y(n329) );
  INVX4 U473 ( .A(A[3]), .Y(n303) );
  INVX8 U474 ( .A(n301), .Y(n302) );
  INVX2 U475 ( .A(n263), .Y(\mult_97/n2217 ) );
  INVX2 U476 ( .A(\mult_97/n1207 ), .Y(\mult_97/n1208 ) );
  INVX2 U477 ( .A(n264), .Y(\mult_97/n2250 ) );
  INVX2 U478 ( .A(\mult_97/n861 ), .Y(\mult_97/n859 ) );
  INVX2 U479 ( .A(\mult_97/n831 ), .Y(\mult_97/n830 ) );
  INVX2 U480 ( .A(\mult_97/n1017 ), .Y(\mult_97/n1018 ) );
  INVX2 U481 ( .A(n259), .Y(\mult_97/n2087 ) );
  INVX2 U482 ( .A(n258), .Y(\mult_97/n2056 ) );
  INVX2 U483 ( .A(\mult_97/n1047 ), .Y(\mult_97/n1048 ) );
  INVX2 U484 ( .A(\mult_97/n1161 ), .Y(\mult_97/n1162 ) );
  INVX2 U485 ( .A(n266), .Y(\mult_97/n2314 ) );
  INVX2 U486 ( .A(n257), .Y(\mult_97/n2023 ) );
  INVX2 U487 ( .A(\mult_97/n969 ), .Y(\mult_97/n970 ) );
  INVX2 U488 ( .A(n256), .Y(\mult_97/n1990 ) );
  INVX2 U489 ( .A(n265), .Y(\mult_97/n2281 ) );
  INVX2 U490 ( .A(n262), .Y(\mult_97/n2184 ) );
  INVX2 U491 ( .A(\mult_97/n1119 ), .Y(\mult_97/n1120 ) );
  INVX2 U492 ( .A(\mult_97/n1257 ), .Y(\mult_97/n1258 ) );
  INVX2 U493 ( .A(n261), .Y(\mult_97/n2153 ) );
  INVX2 U494 ( .A(n260), .Y(\mult_97/n2120 ) );
  INVX2 U495 ( .A(\mult_97/n843 ), .Y(\mult_97/n842 ) );
  INVX2 U496 ( .A(n255), .Y(\mult_97/n1963 ) );
  INVX2 U497 ( .A(\mult_97/n634 ), .Y(\mult_97/n880 ) );
  INVX2 U498 ( .A(\mult_97/n617 ), .Y(\mult_97/n878 ) );
  INVX2 U499 ( .A(\mult_97/n739 ), .Y(\mult_97/n897 ) );
  INVX2 U500 ( .A(\mult_97/n506 ), .Y(\mult_97/n862 ) );
  INVX2 U501 ( .A(n254), .Y(\mult_97/n1930 ) );
  INVX2 U502 ( .A(\mult_97/n927 ), .Y(\mult_97/n928 ) );
  INVX2 U503 ( .A(\mult_97/n559 ), .Y(\mult_97/n558 ) );
  INVX2 U504 ( .A(\mult_97/n624 ), .Y(\mult_97/n623 ) );
  INVX2 U505 ( .A(\mult_97/n607 ), .Y(\mult_97/n606 ) );
  INVX2 U506 ( .A(n253), .Y(\mult_97/n1899 ) );
  INVX2 U507 ( .A(\mult_97/n673 ), .Y(\mult_97/n672 ) );
  INVX2 U508 ( .A(\mult_97/n991 ), .Y(\mult_97/n992 ) );
  INVX2 U509 ( .A(\mult_97/n1369 ), .Y(\mult_97/n1370 ) );
  INVX2 U510 ( .A(\mult_97/n1311 ), .Y(\mult_97/n1312 ) );
  INVX2 U511 ( .A(\mult_97/n1081 ), .Y(\mult_97/n1082 ) );
  INVX2 U512 ( .A(\mult_97/n951 ), .Y(\mult_97/n952 ) );
  INVX2 U513 ( .A(\mult_97/n569 ), .Y(\mult_97/n872 ) );
  INVX1 U514 ( .A(\mult_97/n658 ), .Y(\mult_97/n883 ) );
  INVX4 U515 ( .A(A[0]), .Y(n309) );
  INVX1 U516 ( .A(B[3]), .Y(n397) );
  INVX1 U517 ( .A(B[12]), .Y(n379) );
  INVX1 U518 ( .A(B[8]), .Y(n387) );
  INVX1 U519 ( .A(B[7]), .Y(n389) );
  INVX1 U520 ( .A(B[10]), .Y(n383) );
  INVX1 U521 ( .A(B[9]), .Y(n385) );
  INVX1 U522 ( .A(B[17]), .Y(n369) );
  INVX1 U523 ( .A(B[20]), .Y(n363) );
  INVX1 U524 ( .A(B[6]), .Y(n391) );
  INVX1 U525 ( .A(B[2]), .Y(n399) );
  INVX1 U526 ( .A(B[1]), .Y(n401) );
  INVX1 U527 ( .A(B[24]), .Y(n355) );
  INVX1 U528 ( .A(B[23]), .Y(n357) );
  INVX1 U529 ( .A(B[26]), .Y(n351) );
  INVX1 U530 ( .A(B[25]), .Y(n353) );
  INVX1 U531 ( .A(B[14]), .Y(n375) );
  INVX1 U532 ( .A(B[13]), .Y(n377) );
  INVX2 U533 ( .A(\mult_97/n937 ), .Y(\mult_97/n938 ) );
  INVX1 U534 ( .A(B[27]), .Y(n349) );
  INVX1 U535 ( .A(B[28]), .Y(n347) );
  INVX1 U536 ( .A(B[16]), .Y(n371) );
  INVX1 U537 ( .A(B[15]), .Y(n373) );
  INVX1 U538 ( .A(B[4]), .Y(n395) );
  INVX1 U539 ( .A(B[11]), .Y(n381) );
  INVX1 U540 ( .A(B[18]), .Y(n367) );
  INVX1 U541 ( .A(B[19]), .Y(n365) );
  INVX1 U542 ( .A(B[22]), .Y(n359) );
  INVX1 U543 ( .A(B[21]), .Y(n361) );
  INVX1 U544 ( .A(B[5]), .Y(n393) );
  INVX1 U545 ( .A(B[29]), .Y(n345) );
  INVX1 U546 ( .A(B[30]), .Y(n343) );
  INVX1 U547 ( .A(\B_extended[32] ), .Y(n341) );
  INVX2 U548 ( .A(B[0]), .Y(n402) );
  INVX4 U549 ( .A(n285), .Y(n286) );
  INVX2 U550 ( .A(n268), .Y(n269) );
  INVX2 U551 ( .A(n349), .Y(n348) );
  INVX2 U552 ( .A(n347), .Y(n346) );
  INVX2 U553 ( .A(n371), .Y(n370) );
  INVX2 U554 ( .A(n373), .Y(n372) );
  INVX2 U555 ( .A(n379), .Y(n378) );
  INVX2 U556 ( .A(n381), .Y(n380) );
  INVX2 U557 ( .A(n387), .Y(n386) );
  INVX4 U558 ( .A(n282), .Y(n283) );
  INVX2 U559 ( .A(n359), .Y(n358) );
  INVX2 U560 ( .A(n393), .Y(n392) );
  INVX2 U561 ( .A(n355), .Y(n354) );
  INVX2 U562 ( .A(n353), .Y(n352) );
  INVX2 U563 ( .A(n377), .Y(n376) );
  INVX2 U564 ( .A(n345), .Y(n344) );
  INVX2 U565 ( .A(n343), .Y(n342) );
  INVX2 U566 ( .A(n341), .Y(n340) );
  INVX2 U567 ( .A(n395), .Y(n394) );
  INVX2 U568 ( .A(n397), .Y(n396) );
  INVX2 U569 ( .A(A[21]), .Y(n280) );
  INVX2 U570 ( .A(A[19]), .Y(n282) );
  INVX2 U571 ( .A(n389), .Y(n388) );
  INVX2 U572 ( .A(n383), .Y(n382) );
  INVX2 U573 ( .A(n385), .Y(n384) );
  INVX2 U574 ( .A(n367), .Y(n366) );
  INVX2 U575 ( .A(n369), .Y(n368) );
  INVX2 U576 ( .A(n363), .Y(n362) );
  INVX4 U577 ( .A(n295), .Y(n296) );
  INVX2 U578 ( .A(n365), .Y(n364) );
  INVX2 U579 ( .A(n361), .Y(n360) );
  INVX2 U580 ( .A(n391), .Y(n390) );
  INVX2 U581 ( .A(n399), .Y(n398) );
  INVX2 U582 ( .A(n401), .Y(n400) );
  INVX2 U583 ( .A(n357), .Y(n356) );
  INVX2 U584 ( .A(n351), .Y(n350) );
  INVX4 U585 ( .A(n303), .Y(n304) );
  INVX2 U586 ( .A(n552), .Y(n311) );
  INVX2 U587 ( .A(n375), .Y(n374) );
  INVX2 U588 ( .A(n551), .Y(n316) );
  INVX2 U589 ( .A(\mult_97/n592 ), .Y(\mult_97/n874 ) );
  INVX2 U590 ( .A(\mult_97/n800 ), .Y(\mult_97/n799 ) );
  INVX2 U591 ( .A(\mult_97/n809 ), .Y(\mult_97/n808 ) );
  INVX2 U592 ( .A(n268), .Y(n270) );
  INVX4 U593 ( .A(n534), .Y(n339) );
  INVX8 U594 ( .A(n290), .Y(n291) );
  INVX2 U595 ( .A(A[11]), .Y(n293) );
  INVX8 U596 ( .A(n298), .Y(n299) );
  INVX2 U597 ( .A(A[29]), .Y(n271) );
  INVX1 U598 ( .A(\mult_97/n597 ), .Y(\mult_97/n595 ) );
  INVX2 U599 ( .A(\mult_97/n696 ), .Y(\mult_97/n695 ) );
  INVX1 U600 ( .A(\mult_97/n664 ), .Y(\mult_97/n662 ) );
  INVX1 U601 ( .A(\mult_97/n643 ), .Y(\mult_97/n881 ) );
  INVX1 U602 ( .A(\mult_97/n683 ), .Y(\mult_97/n887 ) );
  INVX1 U603 ( .A(\mult_97/n689 ), .Y(\mult_97/n687 ) );
  INVX1 U604 ( .A(\mult_97/n670 ), .Y(\mult_97/n885 ) );
endmodule


module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push_2, _pushout_d, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90,
         N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103,
         N104, N105, N106, N107, N108, N109, N110, N111, N113, N114, N115,
         N116, N117, N118, N119, N120, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N143, push_0, push_1, \C2/DATA3_1 , n66, n74, n76,
         n281, n283, n285, n287, n289, n291, n293, n295, n297, n299, n301,
         n303, n305, n307, n309, n311, n313, n315, n317, n319, n321, n323,
         n325, n327, n329, n331, n333, n335, n337, n339, n341, n343, n346,
         n349, n352, n355, n358, n361, n364, n367, n370, n373, n376, n379,
         n382, n385, n388, n391, n394, n397, n400, n403, n406, n409, n412,
         n415, n418, n421, n424, n427, n430, n433, n436, n439, n441, n443,
         n445, n447, n449, n451, n453, n455, n457, n459, n461, n463, n465,
         n467, n469, n471, n473, n475, n477, n479, n481, n483, n485, n487,
         n489, n491, n493, n495, n497, n499, n501, n503, n505, n507, n509,
         n511, n512, n513, n514, n515, n516, n517, n524, n527, n530, n533,
         n536, n539, n542, n544, n546, n548, n550, n552, n554, n556, n558,
         n560, n562, n564, n566, n568, n570, n572, n574, n576, n578, n580,
         n582, n584, n586, n588, n590, n592, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n629, n630, n631, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, \C2/Z_63 , \C2/Z_62 , \C2/Z_61 ,
         \C2/Z_60 , \C2/Z_59 , \C2/Z_58 , \C2/Z_57 , \C2/Z_56 , \C2/Z_55 ,
         \C2/Z_54 , \C2/Z_53 , \C2/Z_52 , \C2/Z_51 , \C2/Z_50 , \C2/Z_49 ,
         \C2/Z_48 , \C2/Z_47 , \C2/Z_46 , \C2/Z_45 , \C2/Z_44 , \C2/Z_43 ,
         \C2/Z_42 , \C2/Z_41 , \C2/Z_40 , \C2/Z_39 , \C2/Z_38 , \C2/Z_37 ,
         \C2/Z_36 , \C2/Z_35 , \C2/Z_34 , \C2/Z_33 , \C2/Z_32 , \C2/Z_31 ,
         \C2/Z_30 , \C2/Z_29 , \C2/Z_28 , \C2/Z_27 , \C2/Z_26 , \C2/Z_25 ,
         \C2/Z_24 , \C2/Z_23 , \C2/Z_22 , \C2/Z_21 , \C2/Z_20 , \C2/Z_19 ,
         \C2/Z_18 , \C2/Z_17 , \C2/Z_16 , \C2/Z_15 , \C2/Z_14 , \C2/Z_13 ,
         \C2/Z_12 , \C2/Z_11 , \C2/Z_10 , \C2/Z_9 , \C2/Z_8 , \C2/Z_7 ,
         \C2/Z_6 , \C2/Z_5 , \C2/Z_4 , \C2/Z_3 , \C2/Z_2 , \C2/Z_1 ,
         \ashr_28_1/SH[5] , \ashr_28_1/n969 , \ashr_28_1/n968 ,
         \ashr_28_1/n967 , \ashr_28_1/n966 , \ashr_28_1/n965 ,
         \ashr_28_1/n964 , \ashr_28_1/n963 , \ashr_28_1/n962 ,
         \ashr_28_1/n961 , \ashr_28_1/n960 , \ashr_28_1/n959 ,
         \ashr_28_1/n958 , \ashr_28_1/n957 , \ashr_28_1/n956 ,
         \ashr_28_1/n955 , \ashr_28_1/n954 , \ashr_28_1/n953 ,
         \ashr_28_1/n952 , \ashr_28_1/n951 , \ashr_28_1/n950 ,
         \ashr_28_1/n949 , \ashr_28_1/n948 , \ashr_28_1/n947 ,
         \ashr_28_1/n946 , \ashr_28_1/n945 , \ashr_28_1/n944 ,
         \ashr_28_1/n943 , \ashr_28_1/n942 , \ashr_28_1/n941 ,
         \ashr_28_1/n940 , \ashr_28_1/n939 , \ashr_28_1/n938 ,
         \ashr_28_1/n937 , \ashr_28_1/n936 , \ashr_28_1/n935 ,
         \ashr_28_1/n934 , \ashr_28_1/n933 , \ashr_28_1/n932 ,
         \ashr_28_1/n931 , \ashr_28_1/n930 , \ashr_28_1/n929 ,
         \ashr_28_1/n928 , \ashr_28_1/n927 , \ashr_28_1/n926 ,
         \ashr_28_1/n925 , \ashr_28_1/n924 , \ashr_28_1/n923 ,
         \ashr_28_1/n922 , \ashr_28_1/n921 , \ashr_28_1/n920 ,
         \ashr_28_1/n919 , \ashr_28_1/n918 , \ashr_28_1/n917 ,
         \ashr_28_1/n916 , \ashr_28_1/n915 , \ashr_28_1/n914 ,
         \ashr_28_1/n913 , \ashr_28_1/n912 , \ashr_28_1/n911 ,
         \ashr_28_1/n910 , \ashr_28_1/n909 , \ashr_28_1/n908 ,
         \ashr_28_1/n907 , \ashr_28_1/n906 , \ashr_28_1/n905 ,
         \ashr_28_1/n904 , \ashr_28_1/n903 , \ashr_28_1/n902 ,
         \ashr_28_1/n901 , \ashr_28_1/n900 , \ashr_28_1/n899 ,
         \ashr_28_1/n898 , \ashr_28_1/n897 , \ashr_28_1/n896 ,
         \ashr_28_1/n895 , \ashr_28_1/n894 , \ashr_28_1/n893 ,
         \ashr_28_1/n892 , \ashr_28_1/n891 , \ashr_28_1/n890 ,
         \ashr_28_1/n889 , \ashr_28_1/n888 , \ashr_28_1/n887 ,
         \ashr_28_1/n886 , \ashr_28_1/n885 , \ashr_28_1/n884 ,
         \ashr_28_1/n883 , \ashr_28_1/n882 , \ashr_28_1/n881 ,
         \ashr_28_1/n880 , \ashr_28_1/n879 , \ashr_28_1/n878 ,
         \ashr_28_1/n877 , \ashr_28_1/n876 , \ashr_28_1/n875 ,
         \ashr_28_1/n874 , \ashr_28_1/n873 , \ashr_28_1/n872 ,
         \ashr_28_1/n871 , \ashr_28_1/n870 , \ashr_28_1/n869 ,
         \ashr_28_1/n868 , \ashr_28_1/n867 , \ashr_28_1/n866 ,
         \ashr_28_1/n865 , \ashr_28_1/n864 , \ashr_28_1/n863 ,
         \ashr_28_1/n862 , \ashr_28_1/n861 , \ashr_28_1/n860 ,
         \ashr_28_1/n859 , \ashr_28_1/n858 , \ashr_28_1/n857 ,
         \ashr_28_1/n856 , \ashr_28_1/n855 , \ashr_28_1/n854 ,
         \ashr_28_1/n853 , \ashr_28_1/n852 , \ashr_28_1/n851 ,
         \ashr_28_1/n850 , \ashr_28_1/n849 , \ashr_28_1/n848 ,
         \ashr_28_1/n847 , \ashr_28_1/n846 , \ashr_28_1/n845 ,
         \ashr_28_1/n844 , \ashr_28_1/n843 , \ashr_28_1/n842 ,
         \ashr_28_1/n841 , \ashr_28_1/n840 , \ashr_28_1/n839 ,
         \ashr_28_1/n838 , \ashr_28_1/n837 , \ashr_28_1/n836 ,
         \ashr_28_1/n835 , \ashr_28_1/n834 , \ashr_28_1/n833 ,
         \ashr_28_1/n832 , \ashr_28_1/n831 , \ashr_28_1/n830 ,
         \ashr_28_1/n829 , \ashr_28_1/n828 , \ashr_28_1/n827 ,
         \ashr_28_1/n826 , \ashr_28_1/n825 , \ashr_28_1/n824 ,
         \ashr_28_1/n823 , \ashr_28_1/n822 , \ashr_28_1/n821 ,
         \ashr_28_1/n820 , \ashr_28_1/n819 , \ashr_28_1/n818 ,
         \ashr_28_1/n817 , \ashr_28_1/n816 , \ashr_28_1/n815 ,
         \ashr_28_1/n814 , \ashr_28_1/n813 , \ashr_28_1/n812 ,
         \ashr_28_1/n811 , \ashr_28_1/n810 , \ashr_28_1/n809 ,
         \ashr_28_1/n808 , \ashr_28_1/n807 , \ashr_28_1/n806 ,
         \ashr_28_1/n805 , \ashr_28_1/n804 , \ashr_28_1/n803 ,
         \ashr_28_1/n802 , \ashr_28_1/n801 , \ashr_28_1/n800 ,
         \ashr_28_1/n799 , \ashr_28_1/n798 , \ashr_28_1/n797 ,
         \ashr_28_1/n796 , \ashr_28_1/n795 , \ashr_28_1/n794 ,
         \ashr_28_1/n793 , \ashr_28_1/n792 , \ashr_28_1/n791 ,
         \ashr_28_1/n790 , \ashr_28_1/n789 , \ashr_28_1/n788 ,
         \ashr_28_1/n787 , \ashr_28_1/n786 , \ashr_28_1/n785 ,
         \ashr_28_1/n784 , \ashr_28_1/n783 , \ashr_28_1/n782 ,
         \ashr_28_1/n781 , \ashr_28_1/n780 , \ashr_28_1/n779 ,
         \ashr_28_1/n778 , \ashr_28_1/n777 , \ashr_28_1/n776 ,
         \ashr_28_1/n775 , \ashr_28_1/n774 , \ashr_28_1/n773 ,
         \ashr_28_1/n772 , \ashr_28_1/n771 , \ashr_28_1/n770 ,
         \ashr_28_1/n769 , \ashr_28_1/n768 , \ashr_28_1/n767 ,
         \ashr_28_1/n766 , \ashr_28_1/n765 , \ashr_28_1/n764 ,
         \ashr_28_1/n763 , \ashr_28_1/n762 , \ashr_28_1/n761 ,
         \ashr_28_1/n760 , \ashr_28_1/n759 , \ashr_28_1/n758 ,
         \ashr_28_1/n757 , \ashr_28_1/n756 , \ashr_28_1/n755 ,
         \ashr_28_1/n754 , \ashr_28_1/n753 , \ashr_28_1/n752 ,
         \ashr_28_1/n751 , \ashr_28_1/n750 , \ashr_28_1/n749 ,
         \ashr_28_1/n748 , \ashr_28_1/n747 , \ashr_28_1/n746 ,
         \ashr_28_1/n745 , \ashr_28_1/n744 , \ashr_28_1/n743 ,
         \ashr_28_1/n742 , \ashr_28_1/n741 , \ashr_28_1/n740 ,
         \ashr_28_1/n739 , \ashr_28_1/n738 , \ashr_28_1/n737 ,
         \ashr_28_1/n736 , \ashr_28_1/n735 , \ashr_28_1/n734 ,
         \ashr_28_1/n733 , \ashr_28_1/n732 , \ashr_28_1/n731 ,
         \ashr_28_1/n730 , \ashr_28_1/n729 , \ashr_28_1/n728 ,
         \ashr_28_1/n727 , \ashr_28_1/n726 , \ashr_28_1/n725 ,
         \ashr_28_1/n724 , \ashr_28_1/n723 , \ashr_28_1/n722 ,
         \ashr_28_1/n721 , \ashr_28_1/n720 , \ashr_28_1/n719 ,
         \ashr_28_1/n718 , \ashr_28_1/n717 , \ashr_28_1/n716 ,
         \ashr_28_1/n715 , \ashr_28_1/n714 , \ashr_28_1/n713 ,
         \ashr_28_1/n712 , \ashr_28_1/n711 , \ashr_28_1/n710 ,
         \ashr_28_1/n709 , \ashr_28_1/n708 , \ashr_28_1/n707 ,
         \ashr_28_1/n706 , \ashr_28_1/n705 , \ashr_28_1/n704 ,
         \ashr_28_1/n703 , \ashr_28_1/n702 , \ashr_28_1/n701 ,
         \ashr_28_1/n700 , \ashr_28_1/n699 , \ashr_28_1/n698 ,
         \ashr_28_1/n697 , \ashr_28_1/n696 , \ashr_28_1/n695 ,
         \ashr_28_1/n694 , \ashr_28_1/n693 , \ashr_28_1/n692 ,
         \ashr_28_1/n691 , \ashr_28_1/n690 , \ashr_28_1/n689 ,
         \ashr_28_1/n688 , \ashr_28_1/n687 , \ashr_28_1/n686 ,
         \ashr_28_1/n685 , \ashr_28_1/n684 , \ashr_28_1/n683 ,
         \ashr_28_1/n682 , \ashr_28_1/n681 , \ashr_28_1/n680 ,
         \ashr_28_1/n679 , \ashr_28_1/n678 , \ashr_28_1/n677 ,
         \ashr_28_1/n676 , \ashr_28_1/n675 , \ashr_28_1/n674 ,
         \ashr_28_1/n673 , \ashr_28_1/n672 , \ashr_28_1/n671 ,
         \ashr_28_1/n670 , \ashr_28_1/n669 , \ashr_28_1/n668 ,
         \ashr_28_1/n667 , \ashr_28_1/n666 , \ashr_28_1/n665 ,
         \ashr_28_1/n664 , \ashr_28_1/n663 , \ashr_28_1/n662 ,
         \ashr_28_1/n661 , \ashr_28_1/n660 , \ashr_28_1/n659 ,
         \ashr_28_1/n658 , \ashr_28_1/n657 , \ashr_28_1/n656 ,
         \ashr_28_1/n655 , \ashr_28_1/n654 , \ashr_28_1/n653 ,
         \ashr_28_1/n652 , \ashr_28_1/n651 , \ashr_28_1/n650 ,
         \ashr_28_1/n649 , \ashr_28_1/n648 , \ashr_28_1/n647 ,
         \ashr_28_1/n646 , \ashr_28_1/n645 , \ashr_28_1/n644 ,
         \ashr_28_1/n643 , \ashr_28_1/n642 , \ashr_28_1/n641 ,
         \ashr_28_1/n640 , \ashr_28_1/n639 , \ashr_28_1/n638 ,
         \ashr_28_1/n637 , \ashr_28_1/n636 , \ashr_28_1/n635 ,
         \ashr_28_1/n634 , \ashr_28_1/n633 , \ashr_28_1/n632 ,
         \ashr_28_1/n631 , \ashr_28_1/n630 , \ashr_28_1/n629 ,
         \ashr_28_1/n628 , \ashr_28_1/n627 , \ashr_28_1/n626 ,
         \ashr_28_1/n625 , \ashr_28_1/n624 , \ashr_28_1/n623 ,
         \ashr_28_1/n622 , \ashr_28_1/n621 , \ashr_28_1/n620 ,
         \ashr_28_1/n619 , \ashr_28_1/n618 , \ashr_28_1/n617 ,
         \ashr_28_1/n616 , \ashr_28_1/n615 , \ashr_28_1/n614 ,
         \ashr_28_1/n613 , \ashr_28_1/n612 , \ashr_28_1/n611 ,
         \ashr_28_1/n610 , \ashr_28_1/n609 , \ashr_28_1/n608 ,
         \ashr_28_1/n607 , \ashr_28_1/n606 , \ashr_28_1/n605 ,
         \ashr_28_1/n604 , \ashr_28_1/n603 , \ashr_28_1/n602 ,
         \ashr_28_1/n601 , \ashr_28_1/n600 , \ashr_28_1/n599 ,
         \ashr_28_1/n598 , \ashr_28_1/n597 , \ashr_28_1/n596 ,
         \ashr_28_1/n595 , \ashr_28_1/n594 , \ashr_28_1/n593 ,
         \ashr_28_1/n592 , \ashr_28_1/n591 , \ashr_28_1/n590 ,
         \ashr_28_1/n589 , \ashr_28_1/n588 , \ashr_28_1/n587 ,
         \ashr_28_1/n586 , \ashr_28_1/n585 , \ashr_28_1/n584 ,
         \ashr_28_1/n583 , \ashr_28_1/n582 , \ashr_28_1/n581 ,
         \ashr_28_1/n580 , \DP_OP_19_294_9081/n716 , \DP_OP_19_294_9081/n715 ,
         \DP_OP_19_294_9081/n714 , \DP_OP_19_294_9081/n713 ,
         \DP_OP_19_294_9081/n712 , \DP_OP_19_294_9081/n711 ,
         \DP_OP_19_294_9081/n710 , \DP_OP_19_294_9081/n709 ,
         \DP_OP_19_294_9081/n708 , \DP_OP_19_294_9081/n707 ,
         \DP_OP_19_294_9081/n706 , \DP_OP_19_294_9081/n705 ,
         \DP_OP_19_294_9081/n704 , \DP_OP_19_294_9081/n703 ,
         \DP_OP_19_294_9081/n702 , \DP_OP_19_294_9081/n701 ,
         \DP_OP_19_294_9081/n700 , \DP_OP_19_294_9081/n699 ,
         \DP_OP_19_294_9081/n698 , \DP_OP_19_294_9081/n697 ,
         \DP_OP_19_294_9081/n696 , \DP_OP_19_294_9081/n695 ,
         \DP_OP_19_294_9081/n694 , \DP_OP_19_294_9081/n693 ,
         \DP_OP_19_294_9081/n692 , \DP_OP_19_294_9081/n691 ,
         \DP_OP_19_294_9081/n690 , \DP_OP_19_294_9081/n689 ,
         \DP_OP_19_294_9081/n688 , \DP_OP_19_294_9081/n687 ,
         \DP_OP_19_294_9081/n686 , \DP_OP_19_294_9081/n685 ,
         \DP_OP_19_294_9081/n684 , \DP_OP_19_294_9081/n683 ,
         \DP_OP_19_294_9081/n682 , \DP_OP_19_294_9081/n681 ,
         \DP_OP_19_294_9081/n680 , \DP_OP_19_294_9081/n679 ,
         \DP_OP_19_294_9081/n678 , \DP_OP_19_294_9081/n677 ,
         \DP_OP_19_294_9081/n676 , \DP_OP_19_294_9081/n675 ,
         \DP_OP_19_294_9081/n674 , \DP_OP_19_294_9081/n673 ,
         \DP_OP_19_294_9081/n672 , \DP_OP_19_294_9081/n671 ,
         \DP_OP_19_294_9081/n670 , \DP_OP_19_294_9081/n669 ,
         \DP_OP_19_294_9081/n668 , \DP_OP_19_294_9081/n667 ,
         \DP_OP_19_294_9081/n666 , \DP_OP_19_294_9081/n665 ,
         \DP_OP_19_294_9081/n664 , \DP_OP_19_294_9081/n663 ,
         \DP_OP_19_294_9081/n662 , \DP_OP_19_294_9081/n661 ,
         \DP_OP_19_294_9081/n660 , \DP_OP_19_294_9081/n659 ,
         \DP_OP_19_294_9081/n658 , \DP_OP_19_294_9081/n657 ,
         \DP_OP_19_294_9081/n656 , \DP_OP_19_294_9081/n655 ,
         \DP_OP_19_294_9081/n654 , \DP_OP_19_294_9081/n653 ,
         \DP_OP_19_294_9081/n589 , \DP_OP_19_294_9081/n519 ,
         \DP_OP_19_294_9081/n518 , \DP_OP_19_294_9081/n517 ,
         \DP_OP_19_294_9081/n516 , \DP_OP_19_294_9081/n515 ,
         \DP_OP_19_294_9081/n514 , \DP_OP_19_294_9081/n513 ,
         \DP_OP_19_294_9081/n512 , \DP_OP_19_294_9081/n511 ,
         \DP_OP_19_294_9081/n510 , \DP_OP_19_294_9081/n509 ,
         \DP_OP_19_294_9081/n508 , \DP_OP_19_294_9081/n507 ,
         \DP_OP_19_294_9081/n506 , \DP_OP_19_294_9081/n505 ,
         \DP_OP_19_294_9081/n504 , \DP_OP_19_294_9081/n503 ,
         \DP_OP_19_294_9081/n502 , \DP_OP_19_294_9081/n501 ,
         \DP_OP_19_294_9081/n500 , \DP_OP_19_294_9081/n499 ,
         \DP_OP_19_294_9081/n498 , \DP_OP_19_294_9081/n497 ,
         \DP_OP_19_294_9081/n496 , \DP_OP_19_294_9081/n495 ,
         \DP_OP_19_294_9081/n494 , \DP_OP_19_294_9081/n493 ,
         \DP_OP_19_294_9081/n492 , \DP_OP_19_294_9081/n491 ,
         \DP_OP_19_294_9081/n490 , \DP_OP_19_294_9081/n489 ,
         \DP_OP_19_294_9081/n488 , \DP_OP_19_294_9081/n487 ,
         \DP_OP_19_294_9081/n486 , \DP_OP_19_294_9081/n485 ,
         \DP_OP_19_294_9081/n484 , \DP_OP_19_294_9081/n483 ,
         \DP_OP_19_294_9081/n482 , \DP_OP_19_294_9081/n481 ,
         \DP_OP_19_294_9081/n479 , \DP_OP_19_294_9081/n478 ,
         \DP_OP_19_294_9081/n477 , \DP_OP_19_294_9081/n476 ,
         \DP_OP_19_294_9081/n475 , \DP_OP_19_294_9081/n474 ,
         \DP_OP_19_294_9081/n473 , \DP_OP_19_294_9081/n472 ,
         \DP_OP_19_294_9081/n471 , \DP_OP_19_294_9081/n470 ,
         \DP_OP_19_294_9081/n469 , \DP_OP_19_294_9081/n468 ,
         \DP_OP_19_294_9081/n467 , \DP_OP_19_294_9081/n466 ,
         \DP_OP_19_294_9081/n465 , \DP_OP_19_294_9081/n464 ,
         \DP_OP_19_294_9081/n463 , \DP_OP_19_294_9081/n462 ,
         \DP_OP_19_294_9081/n461 , \DP_OP_19_294_9081/n458 ,
         \DP_OP_19_294_9081/n457 , \DP_OP_19_294_9081/n455 ,
         \DP_OP_19_294_9081/n454 , \DP_OP_19_294_9081/n453 ,
         \DP_OP_19_294_9081/n452 , \DP_OP_19_294_9081/n451 ,
         \DP_OP_19_294_9081/n450 , \DP_OP_19_294_9081/n449 ,
         \DP_OP_19_294_9081/n448 , \DP_OP_19_294_9081/n447 ,
         \DP_OP_19_294_9081/n444 , \DP_OP_19_294_9081/n443 ,
         \DP_OP_19_294_9081/n442 , \DP_OP_19_294_9081/n441 ,
         \DP_OP_19_294_9081/n440 , \DP_OP_19_294_9081/n438 ,
         \DP_OP_19_294_9081/n437 , \DP_OP_19_294_9081/n436 ,
         \DP_OP_19_294_9081/n435 , \DP_OP_19_294_9081/n434 ,
         \DP_OP_19_294_9081/n433 , \DP_OP_19_294_9081/n432 ,
         \DP_OP_19_294_9081/n431 , \DP_OP_19_294_9081/n430 ,
         \DP_OP_19_294_9081/n429 , \DP_OP_19_294_9081/n428 ,
         \DP_OP_19_294_9081/n427 , \DP_OP_19_294_9081/n426 ,
         \DP_OP_19_294_9081/n425 , \DP_OP_19_294_9081/n424 ,
         \DP_OP_19_294_9081/n423 , \DP_OP_19_294_9081/n422 ,
         \DP_OP_19_294_9081/n421 , \DP_OP_19_294_9081/n420 ,
         \DP_OP_19_294_9081/n419 , \DP_OP_19_294_9081/n418 ,
         \DP_OP_19_294_9081/n417 , \DP_OP_19_294_9081/n416 ,
         \DP_OP_19_294_9081/n415 , \DP_OP_19_294_9081/n414 ,
         \DP_OP_19_294_9081/n413 , \DP_OP_19_294_9081/n412 ,
         \DP_OP_19_294_9081/n411 , \DP_OP_19_294_9081/n410 ,
         \DP_OP_19_294_9081/n409 , \DP_OP_19_294_9081/n407 ,
         \DP_OP_19_294_9081/n406 , \DP_OP_19_294_9081/n405 ,
         \DP_OP_19_294_9081/n404 , \DP_OP_19_294_9081/n403 ,
         \DP_OP_19_294_9081/n402 , \DP_OP_19_294_9081/n401 ,
         \DP_OP_19_294_9081/n400 , \DP_OP_19_294_9081/n399 ,
         \DP_OP_19_294_9081/n398 , \DP_OP_19_294_9081/n397 ,
         \DP_OP_19_294_9081/n396 , \DP_OP_19_294_9081/n395 ,
         \DP_OP_19_294_9081/n394 , \DP_OP_19_294_9081/n393 ,
         \DP_OP_19_294_9081/n392 , \DP_OP_19_294_9081/n391 ,
         \DP_OP_19_294_9081/n390 , \DP_OP_19_294_9081/n389 ,
         \DP_OP_19_294_9081/n388 , \DP_OP_19_294_9081/n387 ,
         \DP_OP_19_294_9081/n386 , \DP_OP_19_294_9081/n385 ,
         \DP_OP_19_294_9081/n384 , \DP_OP_19_294_9081/n383 ,
         \DP_OP_19_294_9081/n382 , \DP_OP_19_294_9081/n378 ,
         \DP_OP_19_294_9081/n377 , \DP_OP_19_294_9081/n376 ,
         \DP_OP_19_294_9081/n375 , \DP_OP_19_294_9081/n373 ,
         \DP_OP_19_294_9081/n372 , \DP_OP_19_294_9081/n371 ,
         \DP_OP_19_294_9081/n370 , \DP_OP_19_294_9081/n369 ,
         \DP_OP_19_294_9081/n368 , \DP_OP_19_294_9081/n367 ,
         \DP_OP_19_294_9081/n366 , \DP_OP_19_294_9081/n365 ,
         \DP_OP_19_294_9081/n364 , \DP_OP_19_294_9081/n363 ,
         \DP_OP_19_294_9081/n362 , \DP_OP_19_294_9081/n361 ,
         \DP_OP_19_294_9081/n360 , \DP_OP_19_294_9081/n359 ,
         \DP_OP_19_294_9081/n358 , \DP_OP_19_294_9081/n357 ,
         \DP_OP_19_294_9081/n356 , \DP_OP_19_294_9081/n355 ,
         \DP_OP_19_294_9081/n354 , \DP_OP_19_294_9081/n353 ,
         \DP_OP_19_294_9081/n352 , \DP_OP_19_294_9081/n351 ,
         \DP_OP_19_294_9081/n350 , \DP_OP_19_294_9081/n349 ,
         \DP_OP_19_294_9081/n348 , \DP_OP_19_294_9081/n347 ,
         \DP_OP_19_294_9081/n346 , \DP_OP_19_294_9081/n345 ,
         \DP_OP_19_294_9081/n344 , \DP_OP_19_294_9081/n343 ,
         \DP_OP_19_294_9081/n342 , \DP_OP_19_294_9081/n341 ,
         \DP_OP_19_294_9081/n340 , \DP_OP_19_294_9081/n339 ,
         \DP_OP_19_294_9081/n338 , \DP_OP_19_294_9081/n337 ,
         \DP_OP_19_294_9081/n336 , \DP_OP_19_294_9081/n335 ,
         \DP_OP_19_294_9081/n334 , \DP_OP_19_294_9081/n333 ,
         \DP_OP_19_294_9081/n332 , \DP_OP_19_294_9081/n331 ,
         \DP_OP_19_294_9081/n330 , \DP_OP_19_294_9081/n329 ,
         \DP_OP_19_294_9081/n328 , \DP_OP_19_294_9081/n327 ,
         \DP_OP_19_294_9081/n326 , \DP_OP_19_294_9081/n325 ,
         \DP_OP_19_294_9081/n324 , \DP_OP_19_294_9081/n323 ,
         \DP_OP_19_294_9081/n322 , \DP_OP_19_294_9081/n321 ,
         \DP_OP_19_294_9081/n320 , \DP_OP_19_294_9081/n319 ,
         \DP_OP_19_294_9081/n318 , \DP_OP_19_294_9081/n317 ,
         \DP_OP_19_294_9081/n316 , \DP_OP_19_294_9081/n315 ,
         \DP_OP_19_294_9081/n314 , \DP_OP_19_294_9081/n313 ,
         \DP_OP_19_294_9081/n312 , \DP_OP_19_294_9081/n311 ,
         \DP_OP_19_294_9081/n310 , \DP_OP_19_294_9081/n309 ,
         \DP_OP_19_294_9081/n308 , \DP_OP_19_294_9081/n307 ,
         \DP_OP_19_294_9081/n306 , \DP_OP_19_294_9081/n305 ,
         \DP_OP_19_294_9081/n304 , \DP_OP_19_294_9081/n303 ,
         \DP_OP_19_294_9081/n302 , \DP_OP_19_294_9081/n301 ,
         \DP_OP_19_294_9081/n300 , \DP_OP_19_294_9081/n299 ,
         \DP_OP_19_294_9081/n298 , \DP_OP_19_294_9081/n297 ,
         \DP_OP_19_294_9081/n296 , \DP_OP_19_294_9081/n295 ,
         \DP_OP_19_294_9081/n294 , \DP_OP_19_294_9081/n293 ,
         \DP_OP_19_294_9081/n292 , \DP_OP_19_294_9081/n291 ,
         \DP_OP_19_294_9081/n290 , \DP_OP_19_294_9081/n288 ,
         \DP_OP_19_294_9081/n287 , \DP_OP_19_294_9081/n286 ,
         \DP_OP_19_294_9081/n285 , \DP_OP_19_294_9081/n284 ,
         \DP_OP_19_294_9081/n283 , \DP_OP_19_294_9081/n282 ,
         \DP_OP_19_294_9081/n281 , \DP_OP_19_294_9081/n280 ,
         \DP_OP_19_294_9081/n279 , \DP_OP_19_294_9081/n278 ,
         \DP_OP_19_294_9081/n277 , \DP_OP_19_294_9081/n276 ,
         \DP_OP_19_294_9081/n275 , \DP_OP_19_294_9081/n274 ,
         \DP_OP_19_294_9081/n273 , \DP_OP_19_294_9081/n268 ,
         \DP_OP_19_294_9081/n267 , \DP_OP_19_294_9081/n266 ,
         \DP_OP_19_294_9081/n265 , \DP_OP_19_294_9081/n264 ,
         \DP_OP_19_294_9081/n263 , \DP_OP_19_294_9081/n262 ,
         \DP_OP_19_294_9081/n261 , \DP_OP_19_294_9081/n260 ,
         \DP_OP_19_294_9081/n259 , \DP_OP_19_294_9081/n258 ,
         \DP_OP_19_294_9081/n257 , \DP_OP_19_294_9081/n256 ,
         \DP_OP_19_294_9081/n255 , \DP_OP_19_294_9081/n254 ,
         \DP_OP_19_294_9081/n253 , \DP_OP_19_294_9081/n252 ,
         \DP_OP_19_294_9081/n251 , \DP_OP_19_294_9081/n250 ,
         \DP_OP_19_294_9081/n249 , \DP_OP_19_294_9081/n248 ,
         \DP_OP_19_294_9081/n247 , \DP_OP_19_294_9081/n246 ,
         \DP_OP_19_294_9081/n245 , \DP_OP_19_294_9081/n244 ,
         \DP_OP_19_294_9081/n243 , \DP_OP_19_294_9081/n240 ,
         \DP_OP_19_294_9081/n239 , \DP_OP_19_294_9081/n238 ,
         \DP_OP_19_294_9081/n237 , \DP_OP_19_294_9081/n236 ,
         \DP_OP_19_294_9081/n235 , \DP_OP_19_294_9081/n234 ,
         \DP_OP_19_294_9081/n233 , \DP_OP_19_294_9081/n232 ,
         \DP_OP_19_294_9081/n231 , \DP_OP_19_294_9081/n230 ,
         \DP_OP_19_294_9081/n229 , \DP_OP_19_294_9081/n228 ,
         \DP_OP_19_294_9081/n227 , \DP_OP_19_294_9081/n226 ,
         \DP_OP_19_294_9081/n225 , \DP_OP_19_294_9081/n224 ,
         \DP_OP_19_294_9081/n223 , \DP_OP_19_294_9081/n222 ,
         \DP_OP_19_294_9081/n221 , \DP_OP_19_294_9081/n220 ,
         \DP_OP_19_294_9081/n219 , \DP_OP_19_294_9081/n218 ,
         \DP_OP_19_294_9081/n217 , \DP_OP_19_294_9081/n216 ,
         \DP_OP_19_294_9081/n215 , \DP_OP_19_294_9081/n214 ,
         \DP_OP_19_294_9081/n213 , \DP_OP_19_294_9081/n212 ,
         \DP_OP_19_294_9081/n211 , \DP_OP_19_294_9081/n210 ,
         \DP_OP_19_294_9081/n209 , \DP_OP_19_294_9081/n208 ,
         \DP_OP_19_294_9081/n207 , \DP_OP_19_294_9081/n206 ,
         \DP_OP_19_294_9081/n205 , \DP_OP_19_294_9081/n204 ,
         \DP_OP_19_294_9081/n203 , \DP_OP_19_294_9081/n202 ,
         \DP_OP_19_294_9081/n201 , \DP_OP_19_294_9081/n200 ,
         \DP_OP_19_294_9081/n199 , \DP_OP_19_294_9081/n198 ,
         \DP_OP_19_294_9081/n197 , \DP_OP_19_294_9081/n196 ,
         \DP_OP_19_294_9081/n195 , \DP_OP_19_294_9081/n194 ,
         \DP_OP_19_294_9081/n193 , \DP_OP_19_294_9081/n192 ,
         \DP_OP_19_294_9081/n191 , \DP_OP_19_294_9081/n190 ,
         \DP_OP_19_294_9081/n189 , \DP_OP_19_294_9081/n188 ,
         \DP_OP_19_294_9081/n187 , \DP_OP_19_294_9081/n186 ,
         \DP_OP_19_294_9081/n185 , \DP_OP_19_294_9081/n182 ,
         \DP_OP_19_294_9081/n181 , \DP_OP_19_294_9081/n180 ,
         \DP_OP_19_294_9081/n179 , \DP_OP_19_294_9081/n178 ,
         \DP_OP_19_294_9081/n177 , \DP_OP_19_294_9081/n176 ,
         \DP_OP_19_294_9081/n175 , \DP_OP_19_294_9081/n174 ,
         \DP_OP_19_294_9081/n173 , \DP_OP_19_294_9081/n172 ,
         \DP_OP_19_294_9081/n171 , \DP_OP_19_294_9081/n170 ,
         \DP_OP_19_294_9081/n169 , \DP_OP_19_294_9081/n168 ,
         \DP_OP_19_294_9081/n167 , \DP_OP_19_294_9081/n166 ,
         \DP_OP_19_294_9081/n165 , \DP_OP_19_294_9081/n164 ,
         \DP_OP_19_294_9081/n163 , \DP_OP_19_294_9081/n162 ,
         \DP_OP_19_294_9081/n161 , \DP_OP_19_294_9081/n158 ,
         \DP_OP_19_294_9081/n157 , \DP_OP_19_294_9081/n156 ,
         \DP_OP_19_294_9081/n155 , \DP_OP_19_294_9081/n154 ,
         \DP_OP_19_294_9081/n153 , \DP_OP_19_294_9081/n152 ,
         \DP_OP_19_294_9081/n151 , \DP_OP_19_294_9081/n150 ,
         \DP_OP_19_294_9081/n149 , \DP_OP_19_294_9081/n148 ,
         \DP_OP_19_294_9081/n147 , \DP_OP_19_294_9081/n146 ,
         \DP_OP_19_294_9081/n143 , \DP_OP_19_294_9081/n142 ,
         \DP_OP_19_294_9081/n141 , \DP_OP_19_294_9081/n140 ,
         \DP_OP_19_294_9081/n139 , \DP_OP_19_294_9081/n138 ,
         \DP_OP_19_294_9081/n137 , \DP_OP_19_294_9081/n136 ,
         \DP_OP_19_294_9081/n135 , \DP_OP_19_294_9081/n134 ,
         \DP_OP_19_294_9081/n133 , \DP_OP_19_294_9081/n132 ,
         \DP_OP_19_294_9081/n131 , \DP_OP_19_294_9081/n130 ,
         \DP_OP_19_294_9081/n129 , \DP_OP_19_294_9081/n128 ,
         \DP_OP_19_294_9081/n127 , \DP_OP_19_294_9081/n126 ,
         \DP_OP_19_294_9081/n125 , \DP_OP_19_294_9081/n124 ,
         \DP_OP_19_294_9081/n123 , \DP_OP_19_294_9081/n122 ,
         \DP_OP_19_294_9081/n121 , \DP_OP_19_294_9081/n120 ,
         \DP_OP_19_294_9081/n119 , \DP_OP_19_294_9081/n118 ,
         \DP_OP_19_294_9081/n117 , \DP_OP_19_294_9081/n116 ,
         \DP_OP_19_294_9081/n113 , \DP_OP_19_294_9081/n112 ,
         \DP_OP_19_294_9081/n111 , \DP_OP_19_294_9081/n110 ,
         \DP_OP_19_294_9081/n109 , \DP_OP_19_294_9081/n108 ,
         \DP_OP_19_294_9081/n107 , \DP_OP_19_294_9081/n106 ,
         \DP_OP_19_294_9081/n105 , \DP_OP_19_294_9081/n104 ,
         \DP_OP_19_294_9081/n103 , \DP_OP_19_294_9081/n102 ,
         \DP_OP_19_294_9081/n101 , \DP_OP_19_294_9081/n100 ,
         \DP_OP_19_294_9081/n99 , \DP_OP_19_294_9081/n98 ,
         \DP_OP_19_294_9081/n97 , \DP_OP_19_294_9081/n96 ,
         \DP_OP_19_294_9081/n95 , \DP_OP_19_294_9081/n94 ,
         \DP_OP_19_294_9081/n93 , \DP_OP_19_294_9081/n92 ,
         \DP_OP_19_294_9081/n89 , \DP_OP_19_294_9081/n88 ,
         \DP_OP_19_294_9081/n87 , \DP_OP_19_294_9081/n86 ,
         \DP_OP_19_294_9081/n85 , \DP_OP_19_294_9081/n84 ,
         \DP_OP_19_294_9081/n82 , \DP_OP_19_294_9081/n80 ,
         \DP_OP_19_294_9081/n79 , \DP_OP_19_294_9081/n78 ,
         \DP_OP_19_294_9081/n77 , \DP_OP_19_294_9081/n76 ,
         \DP_OP_19_294_9081/n75 , \DP_OP_19_294_9081/n74 ,
         \DP_OP_19_294_9081/n73 , \DP_OP_19_294_9081/n72 ,
         \DP_OP_19_294_9081/n71 , \DP_OP_19_294_9081/n70 ,
         \DP_OP_19_294_9081/n69 , \DP_OP_19_294_9081/n67 ,
         \DP_OP_19_294_9081/n64 , \DP_OP_19_294_9081/n63 ,
         \DP_OP_19_294_9081/n62 , \DP_OP_19_294_9081/n61 ,
         \DP_OP_19_294_9081/n60 , \DP_OP_19_294_9081/n59 ,
         \DP_OP_19_294_9081/n58 , \DP_OP_19_294_9081/n57 ,
         \DP_OP_19_294_9081/n56 , \DP_OP_19_294_9081/n55 ,
         \DP_OP_19_294_9081/n54 , \DP_OP_19_294_9081/n53 ,
         \DP_OP_19_294_9081/n52 , \DP_OP_19_294_9081/n51 ,
         \DP_OP_19_294_9081/n50 , \DP_OP_19_294_9081/n49 ,
         \DP_OP_19_294_9081/n48 , \DP_OP_19_294_9081/n47 ,
         \DP_OP_19_294_9081/n46 , \DP_OP_19_294_9081/n45 ,
         \DP_OP_19_294_9081/n44 , \DP_OP_19_294_9081/n43 ,
         \DP_OP_19_294_9081/n42 , \DP_OP_19_294_9081/n41 ,
         \DP_OP_19_294_9081/n40 , \DP_OP_19_294_9081/n39 ,
         \DP_OP_19_294_9081/n38 , \DP_OP_19_294_9081/n37 ,
         \DP_OP_19_294_9081/n36 , \DP_OP_19_294_9081/n34 ,
         \DP_OP_19_294_9081/n33 , \DP_OP_19_294_9081/n32 ,
         \DP_OP_19_294_9081/n30 , \DP_OP_19_294_9081/n26 ,
         \DP_OP_19_294_9081/n24 , \DP_OP_19_294_9081/n22 ,
         \DP_OP_19_294_9081/n21 , \DP_OP_19_294_9081/n20 ,
         \DP_OP_19_294_9081/n18 , \DP_OP_19_294_9081/n17 ,
         \DP_OP_19_294_9081/n16 , \DP_OP_19_294_9081/n15 ,
         \DP_OP_19_294_9081/n14 , \DP_OP_19_294_9081/n13 ,
         \DP_OP_19_294_9081/n12 , \DP_OP_19_294_9081/n11 ,
         \DP_OP_19_294_9081/n10 , \DP_OP_19_294_9081/n9 ,
         \DP_OP_19_294_9081/n8 , \DP_OP_19_294_9081/n7 ,
         \DP_OP_19_294_9081/n6 , \DP_OP_19_294_9081/n5 ,
         \DP_OP_19_294_9081/n4 , \DP_OP_19_294_9081/n3 ,
         \DP_OP_19_294_9081/n2 , \DP_OP_19_294_9081/n1 , n672, n674, n675,
         n677, n678, n680, n681, n682, n684, n685, n686, n687, n688, n689,
         n690, n692, n693, n694, n695, n696, n697, n699, n700, n701, n702,
         n703, n704, n706, n708, n709, n710, n711, n712, n714, n715, n716,
         n717, n718, n720, n721, n723, n724, n726, n727, n729, n730, n732,
         n733, n735, n736, n738, n739, n741, n743, n745, n747, n748, n750,
         n751, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n788, n790, n792, n793, n795, n796, n798, n799, n801,
         n802, n804, n805, n807, n808, n810, n811, n813, n814, n816, n817,
         n819, n820, n822, n823, n825, n826, n828, n829, n831, n832, n834,
         n835, n837, n838, n840, n841, n843, n844, n846, n847, n849, n850,
         n852, n853, n855, n856, n858, n859, n861, n862, n864, n865, n867,
         n868, n870, n871, n873, n874, n876, n877, n879, n880, n882, n883,
         n885, n886, n888, n889, n891, n892, n894, n895, n897, n898, n900,
         n901, n903, n904, n906, n907, n909, n910, n912, n913, n915, n916,
         n918, n919, n921, n922, n924, n925, n927, n928, n930, n931, n933,
         n934, n936, n937, n939, n940, n942, n943, n945, n946, n948, n949,
         n951, n952, n954, n955, n957, n958, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] mulout;
  wire   [63:0] acc;
  wire   [6:0] h2;
  wire   [1:0] cmd0;
  wire   [6:0] h1;
  wire   [1:0] cmd_1;

  sfilt_DW02_mult_3_stage_0 pipe ( .A(q0), .B(h0), .TC(1'b1), .CLK(clk), 
        .PRODUCT(mulout) );
  DFFSR \cmd0_reg[1]  ( .D(cmd[1]), .CLK(clk), .R(n630), .S(1'b1), .Q(cmd0[1])
         );
  DFFSR \cmd0_reg[0]  ( .D(cmd[0]), .CLK(clk), .R(n1181), .S(1'b1), .Q(cmd0[0]) );
  DFFSR \h0_reg[31]  ( .D(n592), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[31]) );
  DFFSR \h0_reg[30]  ( .D(n590), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[30]) );
  DFFSR \h0_reg[29]  ( .D(n588), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[29]) );
  DFFSR \h0_reg[28]  ( .D(n586), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[28]) );
  DFFSR \h0_reg[27]  ( .D(n584), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[27]) );
  DFFSR \h0_reg[26]  ( .D(n582), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[26]) );
  DFFSR \h0_reg[25]  ( .D(n580), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[25]) );
  DFFSR \h0_reg[24]  ( .D(n578), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[24]) );
  DFFSR \h0_reg[23]  ( .D(n576), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[23]) );
  DFFSR \h0_reg[22]  ( .D(n574), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[22]) );
  DFFSR \h0_reg[21]  ( .D(n572), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[21]) );
  DFFSR \h0_reg[20]  ( .D(n570), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[20]) );
  DFFSR \h0_reg[19]  ( .D(n568), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[19]) );
  DFFSR \h0_reg[18]  ( .D(n566), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[18]) );
  DFFSR \h0_reg[17]  ( .D(n564), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[17]) );
  DFFSR \h0_reg[16]  ( .D(n562), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[16]) );
  DFFSR \h0_reg[15]  ( .D(n560), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[15]) );
  DFFSR \h0_reg[14]  ( .D(n558), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[14]) );
  DFFSR \h0_reg[13]  ( .D(n556), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[13]) );
  DFFSR \h0_reg[12]  ( .D(n554), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[12]) );
  DFFSR \h0_reg[11]  ( .D(n552), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[11]) );
  DFFSR \h0_reg[10]  ( .D(n550), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[10]) );
  DFFSR \h0_reg[9]  ( .D(n548), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[9]) );
  DFFSR \h0_reg[8]  ( .D(n546), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[8]) );
  DFFSR \h0_reg[7]  ( .D(n544), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[7]) );
  DFFSR \h0_reg[6]  ( .D(n542), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[6]) );
  DFFSR \h1_reg[6]  ( .D(h0[6]), .CLK(clk), .R(n630), .S(1'b1), .Q(h1[6]) );
  DFFSR \h0_reg[5]  ( .D(n539), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[5]) );
  DFFSR \h1_reg[5]  ( .D(h0[5]), .CLK(clk), .R(n630), .S(1'b1), .Q(h1[5]) );
  DFFSR \h0_reg[4]  ( .D(n536), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[4]) );
  DFFSR \h1_reg[4]  ( .D(h0[4]), .CLK(clk), .R(n1181), .S(1'b1), .Q(h1[4]) );
  DFFSR \h0_reg[3]  ( .D(n533), .CLK(clk), .R(n1181), .S(1'b1), .Q(h0[3]) );
  DFFSR \h1_reg[3]  ( .D(h0[3]), .CLK(clk), .R(n630), .S(1'b1), .Q(h1[3]) );
  DFFSR \h0_reg[2]  ( .D(n530), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[2]) );
  DFFSR \h1_reg[2]  ( .D(h0[2]), .CLK(clk), .R(n630), .S(1'b1), .Q(h1[2]) );
  DFFSR \h0_reg[1]  ( .D(n527), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[1]) );
  DFFSR \h1_reg[1]  ( .D(h0[1]), .CLK(clk), .R(n630), .S(1'b1), .Q(h1[1]) );
  DFFSR \h0_reg[0]  ( .D(n524), .CLK(clk), .R(n630), .S(1'b1), .Q(h0[0]) );
  DFFSR \h1_reg[0]  ( .D(h0[0]), .CLK(clk), .R(n630), .S(1'b1), .Q(h1[0]) );
  DFFSR \cmd_1_reg[1]  ( .D(n1087), .CLK(clk), .R(n630), .S(1'b1), .Q(cmd_1[1]) );
  DFFSR \cmd_1_reg[0]  ( .D(n1086), .CLK(clk), .R(n630), .S(1'b1), .Q(cmd_1[0]) );
  DFFSR push_0_reg ( .D(n1169), .CLK(clk), .R(n630), .S(1'b1), .Q(push_0) );
  DFFSR push_1_reg ( .D(n1085), .CLK(clk), .R(n630), .S(1'b1), .Q(push_1) );
  DFFPOSX1 \h2_reg[6]  ( .D(n1063), .CLK(clk), .Q(h2[6]) );
  DFFPOSX1 \h2_reg[5]  ( .D(n516), .CLK(clk), .Q(h2[5]) );
  DFFPOSX1 \h2_reg[4]  ( .D(n515), .CLK(clk), .Q(h2[4]) );
  DFFPOSX1 \h2_reg[3]  ( .D(n514), .CLK(clk), .Q(h2[3]) );
  DFFPOSX1 \h2_reg[2]  ( .D(n1062), .CLK(clk), .Q(h2[2]) );
  DFFPOSX1 \h2_reg[1]  ( .D(n1061), .CLK(clk), .Q(h2[1]) );
  DFFPOSX1 \h2_reg[0]  ( .D(n511), .CLK(clk), .Q(h2[0]) );
  DFFSR push_2_reg ( .D(n1084), .CLK(clk), .R(n1181), .S(1'b1), .Q(push_2) );
  DFFSR \q0_reg[31]  ( .D(n509), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[31]) );
  DFFSR \q0_reg[30]  ( .D(n507), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[30]) );
  DFFSR \q0_reg[29]  ( .D(n505), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[29]) );
  DFFSR \q0_reg[28]  ( .D(n503), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[28]) );
  DFFSR \q0_reg[27]  ( .D(n501), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[27]) );
  DFFSR \q0_reg[26]  ( .D(n499), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[26]) );
  DFFSR \q0_reg[25]  ( .D(n497), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[25]) );
  DFFSR \q0_reg[24]  ( .D(n495), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[24]) );
  DFFSR \q0_reg[23]  ( .D(n493), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[23]) );
  DFFSR \q0_reg[22]  ( .D(n491), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[22]) );
  DFFSR \q0_reg[21]  ( .D(n489), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[21]) );
  DFFSR \q0_reg[20]  ( .D(n487), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[20]) );
  DFFSR \q0_reg[19]  ( .D(n485), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[19]) );
  DFFSR \q0_reg[18]  ( .D(n483), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[18]) );
  DFFSR \q0_reg[17]  ( .D(n481), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[17]) );
  DFFSR \q0_reg[16]  ( .D(n479), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[16]) );
  DFFSR \q0_reg[15]  ( .D(n477), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[15]) );
  DFFSR \q0_reg[14]  ( .D(n475), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[14]) );
  DFFSR \q0_reg[13]  ( .D(n473), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[13]) );
  DFFSR \q0_reg[12]  ( .D(n471), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[12]) );
  DFFSR \q0_reg[11]  ( .D(n469), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[11]) );
  DFFSR \q0_reg[10]  ( .D(n467), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[10]) );
  DFFSR \q0_reg[9]  ( .D(n465), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[9]) );
  DFFSR \q0_reg[8]  ( .D(n463), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[8]) );
  DFFSR \q0_reg[7]  ( .D(n461), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[7]) );
  DFFSR \q0_reg[6]  ( .D(n459), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[6]) );
  DFFSR \q0_reg[5]  ( .D(n457), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[5]) );
  DFFSR \q0_reg[4]  ( .D(n455), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[4]) );
  DFFSR \q0_reg[3]  ( .D(n453), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[3]) );
  DFFSR \q0_reg[2]  ( .D(n451), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[2]) );
  DFFSR \q0_reg[1]  ( .D(n449), .CLK(clk), .R(n1181), .S(1'b1), .Q(q0[1]) );
  DFFSR \q0_reg[0]  ( .D(n447), .CLK(clk), .R(n630), .S(1'b1), .Q(q0[0]) );
  DFFSR \cmd_2_reg[1]  ( .D(n443), .CLK(clk), .R(1'b1), .S(n630), .Q(n445) );
  DFFSR \cmd_2_reg[0]  ( .D(n441), .CLK(clk), .R(1'b1), .S(n630), .Q(n629) );
  DFFSR _pushout_reg ( .D(_pushout_d), .CLK(clk), .R(n1181), .S(1'b1), .Q(
        pushout) );
  DFFSR \acc_reg[0]  ( .D(n439), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[0]) );
  DFFSR \dout_reg[0]  ( .D(n626), .CLK(clk), .R(n630), .S(1'b1), .Q(z[0]) );
  DFFSR \acc_reg[1]  ( .D(n436), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[1]) );
  DFFSR \dout_reg[1]  ( .D(n625), .CLK(clk), .R(n630), .S(1'b1), .Q(z[1]) );
  DFFSR \acc_reg[2]  ( .D(n433), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[2]) );
  DFFSR \dout_reg[2]  ( .D(n624), .CLK(clk), .R(n630), .S(1'b1), .Q(z[2]) );
  DFFSR \acc_reg[3]  ( .D(n430), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[3]) );
  DFFSR \dout_reg[3]  ( .D(n623), .CLK(clk), .R(n630), .S(1'b1), .Q(z[3]) );
  DFFSR \acc_reg[4]  ( .D(n1060), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[4]) );
  DFFSR \dout_reg[4]  ( .D(n622), .CLK(clk), .R(n630), .S(1'b1), .Q(z[4]) );
  DFFSR \acc_reg[5]  ( .D(n1059), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[5]) );
  DFFSR \dout_reg[5]  ( .D(n621), .CLK(clk), .R(n630), .S(1'b1), .Q(z[5]) );
  DFFSR \acc_reg[6]  ( .D(n1058), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[6]) );
  DFFSR \dout_reg[6]  ( .D(n620), .CLK(clk), .R(n630), .S(1'b1), .Q(z[6]) );
  DFFSR \acc_reg[7]  ( .D(n1057), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[7]) );
  DFFSR \dout_reg[7]  ( .D(n619), .CLK(clk), .R(n630), .S(1'b1), .Q(z[7]) );
  DFFSR \acc_reg[8]  ( .D(n1056), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[8]) );
  DFFSR \dout_reg[8]  ( .D(n618), .CLK(clk), .R(n630), .S(1'b1), .Q(z[8]) );
  DFFSR \acc_reg[9]  ( .D(n1055), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[9])
         );
  DFFSR \dout_reg[9]  ( .D(n617), .CLK(clk), .R(n630), .S(1'b1), .Q(z[9]) );
  DFFSR \acc_reg[10]  ( .D(n1054), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[10])
         );
  DFFSR \dout_reg[10]  ( .D(n616), .CLK(clk), .R(n630), .S(1'b1), .Q(z[10]) );
  DFFSR \acc_reg[11]  ( .D(n1053), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[11])
         );
  DFFSR \dout_reg[11]  ( .D(n615), .CLK(clk), .R(n630), .S(1'b1), .Q(z[11]) );
  DFFSR \acc_reg[12]  ( .D(n1052), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[12])
         );
  DFFSR \dout_reg[12]  ( .D(n614), .CLK(clk), .R(n630), .S(1'b1), .Q(z[12]) );
  DFFSR \acc_reg[13]  ( .D(n1051), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[13])
         );
  DFFSR \dout_reg[13]  ( .D(n613), .CLK(clk), .R(n630), .S(1'b1), .Q(z[13]) );
  DFFSR \acc_reg[14]  ( .D(n1050), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[14])
         );
  DFFSR \dout_reg[14]  ( .D(n612), .CLK(clk), .R(n630), .S(1'b1), .Q(z[14]) );
  DFFSR \acc_reg[15]  ( .D(n1049), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[15])
         );
  DFFSR \dout_reg[15]  ( .D(n611), .CLK(clk), .R(n630), .S(1'b1), .Q(z[15]) );
  DFFSR \acc_reg[16]  ( .D(n1048), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[16])
         );
  DFFSR \dout_reg[16]  ( .D(n610), .CLK(clk), .R(n630), .S(1'b1), .Q(z[16]) );
  DFFSR \acc_reg[17]  ( .D(n1047), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[17])
         );
  DFFSR \dout_reg[17]  ( .D(n609), .CLK(clk), .R(n630), .S(1'b1), .Q(z[17]) );
  DFFSR \acc_reg[18]  ( .D(n1046), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[18])
         );
  DFFSR \dout_reg[18]  ( .D(n608), .CLK(clk), .R(n630), .S(1'b1), .Q(z[18]) );
  DFFSR \acc_reg[19]  ( .D(n1083), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[19])
         );
  DFFSR \dout_reg[19]  ( .D(n607), .CLK(clk), .R(n630), .S(1'b1), .Q(z[19]) );
  DFFSR \acc_reg[20]  ( .D(n1045), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[20])
         );
  DFFSR \dout_reg[20]  ( .D(n606), .CLK(clk), .R(n630), .S(1'b1), .Q(z[20]) );
  DFFSR \acc_reg[21]  ( .D(n1044), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[21])
         );
  DFFSR \dout_reg[21]  ( .D(n605), .CLK(clk), .R(n630), .S(1'b1), .Q(z[21]) );
  DFFSR \acc_reg[22]  ( .D(n1043), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[22])
         );
  DFFSR \dout_reg[22]  ( .D(n604), .CLK(clk), .R(n630), .S(1'b1), .Q(z[22]) );
  DFFSR \acc_reg[23]  ( .D(n1042), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[23])
         );
  DFFSR \dout_reg[23]  ( .D(n603), .CLK(clk), .R(n630), .S(1'b1), .Q(z[23]) );
  DFFSR \acc_reg[24]  ( .D(n1041), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[24])
         );
  DFFSR \dout_reg[24]  ( .D(n602), .CLK(clk), .R(n630), .S(1'b1), .Q(z[24]) );
  DFFSR \acc_reg[25]  ( .D(n1040), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[25])
         );
  DFFSR \dout_reg[25]  ( .D(n601), .CLK(clk), .R(n630), .S(1'b1), .Q(z[25]) );
  DFFSR \acc_reg[26]  ( .D(n1039), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[26])
         );
  DFFSR \dout_reg[26]  ( .D(n600), .CLK(clk), .R(n630), .S(1'b1), .Q(z[26]) );
  DFFSR \acc_reg[27]  ( .D(n1038), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[27])
         );
  DFFSR \dout_reg[27]  ( .D(n599), .CLK(clk), .R(n630), .S(1'b1), .Q(z[27]) );
  DFFSR \acc_reg[28]  ( .D(n1037), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[28])
         );
  DFFSR \dout_reg[28]  ( .D(n598), .CLK(clk), .R(n630), .S(1'b1), .Q(z[28]) );
  DFFSR \acc_reg[29]  ( .D(n1036), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[29])
         );
  DFFSR \dout_reg[29]  ( .D(n597), .CLK(clk), .R(n630), .S(1'b1), .Q(z[29]) );
  DFFSR \acc_reg[30]  ( .D(n1035), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[30])
         );
  DFFSR \dout_reg[30]  ( .D(n596), .CLK(clk), .R(n630), .S(1'b1), .Q(z[30]) );
  DFFSR \acc_reg[31]  ( .D(n1034), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[31])
         );
  DFFSR \dout_reg[31]  ( .D(n595), .CLK(clk), .R(n630), .S(1'b1), .Q(z[31]) );
  DFFSR \acc_reg[32]  ( .D(n1082), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[32])
         );
  DFFSR \acc_reg[33]  ( .D(n341), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[33])
         );
  DFFSR \acc_reg[34]  ( .D(n1081), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[34])
         );
  DFFSR \acc_reg[35]  ( .D(n337), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[35])
         );
  DFFSR \acc_reg[36]  ( .D(n1080), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[36])
         );
  DFFSR \acc_reg[37]  ( .D(n333), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[37])
         );
  DFFSR \acc_reg[38]  ( .D(n1079), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[38])
         );
  DFFSR \acc_reg[39]  ( .D(n329), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[39])
         );
  DFFSR \acc_reg[40]  ( .D(n327), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[40])
         );
  DFFSR \acc_reg[41]  ( .D(n325), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[41])
         );
  DFFSR \acc_reg[42]  ( .D(n1078), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[42])
         );
  DFFSR \acc_reg[43]  ( .D(n321), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[43])
         );
  DFFSR \acc_reg[44]  ( .D(n1077), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[44])
         );
  DFFSR \acc_reg[45]  ( .D(n317), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[45])
         );
  DFFSR \acc_reg[46]  ( .D(n1076), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[46])
         );
  DFFSR \acc_reg[47]  ( .D(n313), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[47])
         );
  DFFSR \acc_reg[48]  ( .D(n1075), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[48])
         );
  DFFSR \acc_reg[49]  ( .D(n309), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[49])
         );
  DFFSR \acc_reg[50]  ( .D(n1074), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[50])
         );
  DFFSR \acc_reg[51]  ( .D(n305), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[51])
         );
  DFFSR \acc_reg[52]  ( .D(n1073), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[52])
         );
  DFFSR \acc_reg[53]  ( .D(n301), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[53])
         );
  DFFSR \acc_reg[54]  ( .D(n1072), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[54])
         );
  DFFSR \acc_reg[55]  ( .D(n297), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[55])
         );
  DFFSR \acc_reg[56]  ( .D(n1071), .CLK(clk), .R(n1181), .S(1'b1), .Q(acc[56])
         );
  DFFSR \acc_reg[57]  ( .D(n293), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[57])
         );
  DFFSR \acc_reg[58]  ( .D(n1070), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[58])
         );
  DFFSR \acc_reg[59]  ( .D(n289), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[59])
         );
  DFFSR \acc_reg[60]  ( .D(n1069), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[60])
         );
  DFFSR \acc_reg[61]  ( .D(n285), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[61])
         );
  DFFSR \acc_reg[62]  ( .D(n1068), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[62])
         );
  DFFSR \acc_reg[63]  ( .D(n281), .CLK(clk), .R(n630), .S(1'b1), .Q(acc[63])
         );
  OAI21X1 U103 ( .A(n1147), .B(n630), .C(n66), .Y(n517) );
  OAI21X1 U115 ( .A(n630), .B(n1157), .C(n74), .Y(n513) );
  OAI21X1 U118 ( .A(n630), .B(n1161), .C(n76), .Y(n512) );
  INVX1 U516 ( .A(cmd_1[0]), .Y(n441) );
  INVX1 U518 ( .A(cmd_1[1]), .Y(n443) );
  AOI22X1 U632 ( .A(n1378), .B(acc[0]), .C(z[0]), .D(n1180), .Y(n631) );
  AOI22X1 U633 ( .A(n1378), .B(acc[1]), .C(z[1]), .D(n1180), .Y(n633) );
  AOI22X1 U634 ( .A(n1378), .B(acc[2]), .C(z[2]), .D(n1180), .Y(n634) );
  AOI22X1 U635 ( .A(n1378), .B(acc[3]), .C(z[3]), .D(n1180), .Y(n635) );
  AOI22X1 U636 ( .A(n1378), .B(acc[4]), .C(z[4]), .D(n1180), .Y(n636) );
  AOI22X1 U637 ( .A(n1378), .B(acc[5]), .C(z[5]), .D(n1180), .Y(n637) );
  AOI22X1 U638 ( .A(n1378), .B(acc[6]), .C(z[6]), .D(n1180), .Y(n638) );
  AOI22X1 U639 ( .A(n1378), .B(acc[7]), .C(z[7]), .D(n1180), .Y(n639) );
  AOI22X1 U640 ( .A(n1378), .B(acc[8]), .C(z[8]), .D(n1180), .Y(n640) );
  AOI22X1 U641 ( .A(n1378), .B(acc[9]), .C(z[9]), .D(n1180), .Y(n641) );
  AOI22X1 U642 ( .A(n1378), .B(acc[10]), .C(z[10]), .D(n1180), .Y(n642) );
  AOI22X1 U643 ( .A(n1378), .B(acc[11]), .C(z[11]), .D(n1180), .Y(n643) );
  AOI22X1 U644 ( .A(n1378), .B(acc[12]), .C(z[12]), .D(n1180), .Y(n644) );
  AOI22X1 U645 ( .A(n1378), .B(acc[13]), .C(z[13]), .D(n1180), .Y(n645) );
  AOI22X1 U646 ( .A(n1378), .B(acc[14]), .C(z[14]), .D(n1180), .Y(n646) );
  AOI22X1 U647 ( .A(n1378), .B(acc[15]), .C(z[15]), .D(n1180), .Y(n647) );
  AOI22X1 U648 ( .A(n1378), .B(acc[16]), .C(z[16]), .D(n1180), .Y(n648) );
  AOI22X1 U649 ( .A(n1378), .B(acc[17]), .C(z[17]), .D(n1180), .Y(n649) );
  AOI22X1 U650 ( .A(n1378), .B(acc[18]), .C(z[18]), .D(n1180), .Y(n650) );
  AOI22X1 U651 ( .A(n1378), .B(acc[19]), .C(z[19]), .D(n1180), .Y(n651) );
  AOI22X1 U652 ( .A(n1378), .B(acc[20]), .C(z[20]), .D(n1180), .Y(n652) );
  AOI22X1 U653 ( .A(n1378), .B(acc[21]), .C(z[21]), .D(n1180), .Y(n653) );
  AOI22X1 U654 ( .A(n1378), .B(acc[22]), .C(z[22]), .D(n1180), .Y(n654) );
  AOI22X1 U655 ( .A(n1378), .B(acc[23]), .C(z[23]), .D(n1180), .Y(n655) );
  AOI22X1 U656 ( .A(n1378), .B(acc[24]), .C(z[24]), .D(n1180), .Y(n656) );
  AOI22X1 U657 ( .A(n1378), .B(acc[25]), .C(z[25]), .D(n1180), .Y(n657) );
  AOI22X1 U658 ( .A(n1378), .B(acc[26]), .C(z[26]), .D(n1180), .Y(n658) );
  AOI22X1 U659 ( .A(n1378), .B(acc[27]), .C(z[27]), .D(n1180), .Y(n659) );
  AOI22X1 U660 ( .A(n1378), .B(acc[28]), .C(z[28]), .D(n1180), .Y(n660) );
  AOI22X1 U661 ( .A(n1378), .B(acc[29]), .C(z[29]), .D(n1180), .Y(n661) );
  AOI22X1 U662 ( .A(n1378), .B(acc[30]), .C(z[30]), .D(n1180), .Y(n662) );
  AOI22X1 U663 ( .A(n1378), .B(acc[31]), .C(z[31]), .D(n1180), .Y(n663) );
  NAND2X1 \ashr_28_1/U440  ( .A(n1153), .B(acc[31]), .Y(\ashr_28_1/n905 ) );
  MUX2X1 \ashr_28_1/U439  ( .B(acc[0]), .A(acc[32]), .S(n1152), .Y(
        \ashr_28_1/n906 ) );
  MUX2X1 \ashr_28_1/U438  ( .B(acc[1]), .A(acc[33]), .S(n1153), .Y(
        \ashr_28_1/n907 ) );
  MUX2X1 \ashr_28_1/U437  ( .B(acc[2]), .A(acc[34]), .S(n1152), .Y(
        \ashr_28_1/n908 ) );
  MUX2X1 \ashr_28_1/U436  ( .B(acc[3]), .A(acc[35]), .S(n1153), .Y(
        \ashr_28_1/n909 ) );
  MUX2X1 \ashr_28_1/U435  ( .B(acc[4]), .A(acc[36]), .S(n1153), .Y(
        \ashr_28_1/n910 ) );
  MUX2X1 \ashr_28_1/U434  ( .B(acc[5]), .A(acc[37]), .S(n1152), .Y(
        \ashr_28_1/n911 ) );
  MUX2X1 \ashr_28_1/U433  ( .B(acc[6]), .A(acc[38]), .S(n1152), .Y(
        \ashr_28_1/n912 ) );
  MUX2X1 \ashr_28_1/U432  ( .B(acc[7]), .A(acc[39]), .S(n1153), .Y(
        \ashr_28_1/n913 ) );
  MUX2X1 \ashr_28_1/U431  ( .B(acc[8]), .A(acc[40]), .S(n1152), .Y(
        \ashr_28_1/n914 ) );
  MUX2X1 \ashr_28_1/U430  ( .B(acc[9]), .A(acc[41]), .S(n1152), .Y(
        \ashr_28_1/n915 ) );
  MUX2X1 \ashr_28_1/U429  ( .B(acc[10]), .A(acc[42]), .S(n1152), .Y(
        \ashr_28_1/n916 ) );
  MUX2X1 \ashr_28_1/U428  ( .B(acc[11]), .A(acc[43]), .S(n1152), .Y(
        \ashr_28_1/n917 ) );
  MUX2X1 \ashr_28_1/U427  ( .B(acc[12]), .A(acc[44]), .S(n1152), .Y(
        \ashr_28_1/n918 ) );
  MUX2X1 \ashr_28_1/U426  ( .B(acc[13]), .A(acc[45]), .S(n1152), .Y(
        \ashr_28_1/n919 ) );
  MUX2X1 \ashr_28_1/U425  ( .B(acc[14]), .A(acc[46]), .S(n1152), .Y(
        \ashr_28_1/n920 ) );
  MUX2X1 \ashr_28_1/U424  ( .B(acc[15]), .A(acc[47]), .S(n1152), .Y(
        \ashr_28_1/n921 ) );
  MUX2X1 \ashr_28_1/U423  ( .B(acc[16]), .A(acc[48]), .S(n1152), .Y(
        \ashr_28_1/n922 ) );
  MUX2X1 \ashr_28_1/U422  ( .B(acc[17]), .A(acc[49]), .S(n1152), .Y(
        \ashr_28_1/n923 ) );
  MUX2X1 \ashr_28_1/U421  ( .B(acc[18]), .A(acc[50]), .S(n1152), .Y(
        \ashr_28_1/n924 ) );
  MUX2X1 \ashr_28_1/U420  ( .B(acc[19]), .A(acc[51]), .S(n1152), .Y(
        \ashr_28_1/n925 ) );
  MUX2X1 \ashr_28_1/U419  ( .B(acc[20]), .A(acc[52]), .S(n1153), .Y(
        \ashr_28_1/n926 ) );
  MUX2X1 \ashr_28_1/U418  ( .B(acc[21]), .A(acc[53]), .S(n1153), .Y(
        \ashr_28_1/n927 ) );
  MUX2X1 \ashr_28_1/U417  ( .B(acc[22]), .A(acc[54]), .S(n1153), .Y(
        \ashr_28_1/n928 ) );
  MUX2X1 \ashr_28_1/U416  ( .B(acc[23]), .A(acc[55]), .S(n1153), .Y(
        \ashr_28_1/n929 ) );
  MUX2X1 \ashr_28_1/U415  ( .B(acc[24]), .A(acc[56]), .S(n1153), .Y(
        \ashr_28_1/n930 ) );
  MUX2X1 \ashr_28_1/U414  ( .B(acc[25]), .A(acc[57]), .S(n1153), .Y(
        \ashr_28_1/n931 ) );
  MUX2X1 \ashr_28_1/U413  ( .B(acc[26]), .A(acc[58]), .S(n1153), .Y(
        \ashr_28_1/n932 ) );
  MUX2X1 \ashr_28_1/U412  ( .B(acc[27]), .A(acc[59]), .S(n1153), .Y(
        \ashr_28_1/n933 ) );
  MUX2X1 \ashr_28_1/U411  ( .B(acc[28]), .A(acc[60]), .S(n1153), .Y(
        \ashr_28_1/n934 ) );
  MUX2X1 \ashr_28_1/U410  ( .B(acc[29]), .A(acc[61]), .S(n1153), .Y(
        \ashr_28_1/n935 ) );
  MUX2X1 \ashr_28_1/U409  ( .B(acc[30]), .A(acc[62]), .S(n1153), .Y(
        \ashr_28_1/n936 ) );
  MUX2X1 \ashr_28_1/U408  ( .B(acc[31]), .A(acc[63]), .S(n1153), .Y(
        \ashr_28_1/n937 ) );
  MUX2X1 \ashr_28_1/U407  ( .B(\ashr_28_1/n905 ), .A(\ashr_28_1/n969 ), .S(
        n1148), .Y(\ashr_28_1/n840 ) );
  NOR2X1 \ashr_28_1/U406  ( .A(n1149), .B(\ashr_28_1/n906 ), .Y(
        \ashr_28_1/n841 ) );
  NOR2X1 \ashr_28_1/U405  ( .A(n1148), .B(\ashr_28_1/n907 ), .Y(
        \ashr_28_1/n842 ) );
  NOR2X1 \ashr_28_1/U404  ( .A(n1148), .B(\ashr_28_1/n908 ), .Y(
        \ashr_28_1/n843 ) );
  NOR2X1 \ashr_28_1/U403  ( .A(n1149), .B(\ashr_28_1/n909 ), .Y(
        \ashr_28_1/n844 ) );
  NOR2X1 \ashr_28_1/U402  ( .A(n1149), .B(\ashr_28_1/n910 ), .Y(
        \ashr_28_1/n845 ) );
  NOR2X1 \ashr_28_1/U401  ( .A(n1148), .B(\ashr_28_1/n911 ), .Y(
        \ashr_28_1/n846 ) );
  NOR2X1 \ashr_28_1/U400  ( .A(n1148), .B(\ashr_28_1/n912 ), .Y(
        \ashr_28_1/n847 ) );
  NOR2X1 \ashr_28_1/U399  ( .A(n1149), .B(\ashr_28_1/n913 ), .Y(
        \ashr_28_1/n848 ) );
  NOR2X1 \ashr_28_1/U398  ( .A(n1148), .B(\ashr_28_1/n914 ), .Y(
        \ashr_28_1/n849 ) );
  NOR2X1 \ashr_28_1/U397  ( .A(n1149), .B(\ashr_28_1/n915 ), .Y(
        \ashr_28_1/n850 ) );
  NOR2X1 \ashr_28_1/U396  ( .A(n1149), .B(\ashr_28_1/n916 ), .Y(
        \ashr_28_1/n851 ) );
  NOR2X1 \ashr_28_1/U395  ( .A(n1149), .B(\ashr_28_1/n917 ), .Y(
        \ashr_28_1/n852 ) );
  NOR2X1 \ashr_28_1/U394  ( .A(n1148), .B(\ashr_28_1/n918 ), .Y(
        \ashr_28_1/n853 ) );
  NOR2X1 \ashr_28_1/U393  ( .A(n1149), .B(\ashr_28_1/n919 ), .Y(
        \ashr_28_1/n854 ) );
  NOR2X1 \ashr_28_1/U392  ( .A(n1149), .B(\ashr_28_1/n920 ), .Y(
        \ashr_28_1/n855 ) );
  NOR2X1 \ashr_28_1/U391  ( .A(n1149), .B(\ashr_28_1/n921 ), .Y(
        \ashr_28_1/n856 ) );
  NOR2X1 \ashr_28_1/U390  ( .A(n1149), .B(\ashr_28_1/n922 ), .Y(
        \ashr_28_1/n857 ) );
  NOR2X1 \ashr_28_1/U389  ( .A(n1149), .B(\ashr_28_1/n923 ), .Y(
        \ashr_28_1/n858 ) );
  NOR2X1 \ashr_28_1/U388  ( .A(n1149), .B(\ashr_28_1/n924 ), .Y(
        \ashr_28_1/n859 ) );
  NOR2X1 \ashr_28_1/U387  ( .A(n1149), .B(\ashr_28_1/n925 ), .Y(
        \ashr_28_1/n860 ) );
  NOR2X1 \ashr_28_1/U386  ( .A(n1149), .B(\ashr_28_1/n926 ), .Y(
        \ashr_28_1/n861 ) );
  NOR2X1 \ashr_28_1/U385  ( .A(n1149), .B(\ashr_28_1/n927 ), .Y(
        \ashr_28_1/n862 ) );
  NOR2X1 \ashr_28_1/U384  ( .A(n1149), .B(\ashr_28_1/n928 ), .Y(
        \ashr_28_1/n863 ) );
  NOR2X1 \ashr_28_1/U383  ( .A(n1149), .B(\ashr_28_1/n929 ), .Y(
        \ashr_28_1/n864 ) );
  NOR2X1 \ashr_28_1/U382  ( .A(n1149), .B(\ashr_28_1/n930 ), .Y(
        \ashr_28_1/n865 ) );
  NOR2X1 \ashr_28_1/U381  ( .A(n1149), .B(\ashr_28_1/n931 ), .Y(
        \ashr_28_1/n866 ) );
  NOR2X1 \ashr_28_1/U380  ( .A(n1149), .B(\ashr_28_1/n932 ), .Y(
        \ashr_28_1/n867 ) );
  NOR2X1 \ashr_28_1/U379  ( .A(n1149), .B(\ashr_28_1/n933 ), .Y(
        \ashr_28_1/n868 ) );
  NOR2X1 \ashr_28_1/U378  ( .A(n1149), .B(\ashr_28_1/n934 ), .Y(
        \ashr_28_1/n869 ) );
  NOR2X1 \ashr_28_1/U377  ( .A(n1149), .B(\ashr_28_1/n935 ), .Y(
        \ashr_28_1/n870 ) );
  NOR2X1 \ashr_28_1/U376  ( .A(n1149), .B(\ashr_28_1/n936 ), .Y(
        \ashr_28_1/n871 ) );
  NOR2X1 \ashr_28_1/U375  ( .A(n1149), .B(\ashr_28_1/n937 ), .Y(
        \ashr_28_1/n872 ) );
  NOR2X1 \ashr_28_1/U374  ( .A(n1149), .B(\ashr_28_1/n938 ), .Y(
        \ashr_28_1/n873 ) );
  NOR2X1 \ashr_28_1/U373  ( .A(n1149), .B(\ashr_28_1/n939 ), .Y(
        \ashr_28_1/n874 ) );
  NOR2X1 \ashr_28_1/U372  ( .A(n1149), .B(\ashr_28_1/n940 ), .Y(
        \ashr_28_1/n875 ) );
  NOR2X1 \ashr_28_1/U371  ( .A(n1149), .B(\ashr_28_1/n941 ), .Y(
        \ashr_28_1/n876 ) );
  NOR2X1 \ashr_28_1/U370  ( .A(n1149), .B(\ashr_28_1/n942 ), .Y(
        \ashr_28_1/n877 ) );
  NOR2X1 \ashr_28_1/U369  ( .A(n1149), .B(\ashr_28_1/n943 ), .Y(
        \ashr_28_1/n878 ) );
  NOR2X1 \ashr_28_1/U368  ( .A(n1149), .B(\ashr_28_1/n944 ), .Y(
        \ashr_28_1/n879 ) );
  NOR2X1 \ashr_28_1/U367  ( .A(n1149), .B(\ashr_28_1/n945 ), .Y(
        \ashr_28_1/n880 ) );
  NOR2X1 \ashr_28_1/U366  ( .A(n1149), .B(\ashr_28_1/n946 ), .Y(
        \ashr_28_1/n881 ) );
  NOR2X1 \ashr_28_1/U365  ( .A(n1149), .B(\ashr_28_1/n947 ), .Y(
        \ashr_28_1/n882 ) );
  NOR2X1 \ashr_28_1/U364  ( .A(n1149), .B(\ashr_28_1/n948 ), .Y(
        \ashr_28_1/n883 ) );
  NOR2X1 \ashr_28_1/U363  ( .A(n1149), .B(\ashr_28_1/n949 ), .Y(
        \ashr_28_1/n884 ) );
  NOR2X1 \ashr_28_1/U362  ( .A(n1149), .B(\ashr_28_1/n950 ), .Y(
        \ashr_28_1/n885 ) );
  NOR2X1 \ashr_28_1/U361  ( .A(n1149), .B(\ashr_28_1/n951 ), .Y(
        \ashr_28_1/n886 ) );
  NOR2X1 \ashr_28_1/U360  ( .A(n1149), .B(\ashr_28_1/n952 ), .Y(
        \ashr_28_1/n887 ) );
  NOR2X1 \ashr_28_1/U359  ( .A(n1149), .B(\ashr_28_1/n953 ), .Y(
        \ashr_28_1/n888 ) );
  NOR2X1 \ashr_28_1/U358  ( .A(n1149), .B(\ashr_28_1/n954 ), .Y(
        \ashr_28_1/n889 ) );
  NOR2X1 \ashr_28_1/U357  ( .A(n1149), .B(\ashr_28_1/n955 ), .Y(
        \ashr_28_1/n890 ) );
  NOR2X1 \ashr_28_1/U356  ( .A(n1148), .B(\ashr_28_1/n956 ), .Y(
        \ashr_28_1/n891 ) );
  NOR2X1 \ashr_28_1/U355  ( .A(n1148), .B(\ashr_28_1/n957 ), .Y(
        \ashr_28_1/n892 ) );
  NOR2X1 \ashr_28_1/U354  ( .A(n1148), .B(\ashr_28_1/n958 ), .Y(
        \ashr_28_1/n893 ) );
  NOR2X1 \ashr_28_1/U353  ( .A(n1148), .B(\ashr_28_1/n959 ), .Y(
        \ashr_28_1/n894 ) );
  NOR2X1 \ashr_28_1/U352  ( .A(n1148), .B(\ashr_28_1/n960 ), .Y(
        \ashr_28_1/n895 ) );
  NOR2X1 \ashr_28_1/U351  ( .A(n1148), .B(\ashr_28_1/n961 ), .Y(
        \ashr_28_1/n896 ) );
  NOR2X1 \ashr_28_1/U350  ( .A(n1148), .B(\ashr_28_1/n962 ), .Y(
        \ashr_28_1/n897 ) );
  NOR2X1 \ashr_28_1/U349  ( .A(n1148), .B(\ashr_28_1/n963 ), .Y(
        \ashr_28_1/n898 ) );
  NOR2X1 \ashr_28_1/U348  ( .A(n1148), .B(\ashr_28_1/n964 ), .Y(
        \ashr_28_1/n899 ) );
  NOR2X1 \ashr_28_1/U347  ( .A(n1148), .B(\ashr_28_1/n965 ), .Y(
        \ashr_28_1/n900 ) );
  NOR2X1 \ashr_28_1/U346  ( .A(n1148), .B(\ashr_28_1/n966 ), .Y(
        \ashr_28_1/n901 ) );
  NOR2X1 \ashr_28_1/U345  ( .A(n1148), .B(\ashr_28_1/n967 ), .Y(
        \ashr_28_1/n902 ) );
  NOR2X1 \ashr_28_1/U344  ( .A(n1148), .B(\ashr_28_1/n968 ), .Y(
        \ashr_28_1/n903 ) );
  NOR2X1 \ashr_28_1/U343  ( .A(n1148), .B(\ashr_28_1/n969 ), .Y(
        \ashr_28_1/n904 ) );
  MUX2X1 \ashr_28_1/U342  ( .B(\ashr_28_1/n840 ), .A(\ashr_28_1/n856 ), .S(
        n1065), .Y(\ashr_28_1/n775 ) );
  MUX2X1 \ashr_28_1/U341  ( .B(\ashr_28_1/n841 ), .A(\ashr_28_1/n857 ), .S(
        n1065), .Y(\ashr_28_1/n776 ) );
  MUX2X1 \ashr_28_1/U340  ( .B(\ashr_28_1/n842 ), .A(\ashr_28_1/n858 ), .S(
        n1065), .Y(\ashr_28_1/n777 ) );
  MUX2X1 \ashr_28_1/U339  ( .B(\ashr_28_1/n843 ), .A(\ashr_28_1/n859 ), .S(
        n1065), .Y(\ashr_28_1/n778 ) );
  MUX2X1 \ashr_28_1/U338  ( .B(\ashr_28_1/n844 ), .A(\ashr_28_1/n860 ), .S(
        n1065), .Y(\ashr_28_1/n779 ) );
  MUX2X1 \ashr_28_1/U337  ( .B(\ashr_28_1/n845 ), .A(\ashr_28_1/n861 ), .S(
        n1065), .Y(\ashr_28_1/n780 ) );
  MUX2X1 \ashr_28_1/U336  ( .B(\ashr_28_1/n846 ), .A(\ashr_28_1/n862 ), .S(
        n1065), .Y(\ashr_28_1/n781 ) );
  MUX2X1 \ashr_28_1/U335  ( .B(\ashr_28_1/n847 ), .A(\ashr_28_1/n863 ), .S(
        n1065), .Y(\ashr_28_1/n782 ) );
  MUX2X1 \ashr_28_1/U333  ( .B(\ashr_28_1/n849 ), .A(\ashr_28_1/n865 ), .S(
        n1065), .Y(\ashr_28_1/n784 ) );
  MUX2X1 \ashr_28_1/U332  ( .B(\ashr_28_1/n850 ), .A(\ashr_28_1/n866 ), .S(
        n1065), .Y(\ashr_28_1/n785 ) );
  MUX2X1 \ashr_28_1/U331  ( .B(\ashr_28_1/n851 ), .A(\ashr_28_1/n867 ), .S(
        n1065), .Y(\ashr_28_1/n786 ) );
  MUX2X1 \ashr_28_1/U330  ( .B(\ashr_28_1/n852 ), .A(\ashr_28_1/n868 ), .S(
        n1065), .Y(\ashr_28_1/n787 ) );
  MUX2X1 \ashr_28_1/U329  ( .B(\ashr_28_1/n853 ), .A(\ashr_28_1/n869 ), .S(
        n1065), .Y(\ashr_28_1/n788 ) );
  MUX2X1 \ashr_28_1/U328  ( .B(\ashr_28_1/n854 ), .A(\ashr_28_1/n870 ), .S(
        n1065), .Y(\ashr_28_1/n789 ) );
  MUX2X1 \ashr_28_1/U326  ( .B(\ashr_28_1/n856 ), .A(\ashr_28_1/n872 ), .S(
        n1065), .Y(\ashr_28_1/n791 ) );
  MUX2X1 \ashr_28_1/U325  ( .B(\ashr_28_1/n857 ), .A(\ashr_28_1/n873 ), .S(
        n1065), .Y(\ashr_28_1/n792 ) );
  MUX2X1 \ashr_28_1/U324  ( .B(\ashr_28_1/n858 ), .A(\ashr_28_1/n874 ), .S(
        n1065), .Y(\ashr_28_1/n793 ) );
  MUX2X1 \ashr_28_1/U322  ( .B(\ashr_28_1/n860 ), .A(\ashr_28_1/n876 ), .S(
        n1065), .Y(\ashr_28_1/n795 ) );
  MUX2X1 \ashr_28_1/U320  ( .B(\ashr_28_1/n862 ), .A(\ashr_28_1/n878 ), .S(
        n1065), .Y(\ashr_28_1/n797 ) );
  MUX2X1 \ashr_28_1/U318  ( .B(\ashr_28_1/n864 ), .A(\ashr_28_1/n880 ), .S(
        n1065), .Y(\ashr_28_1/n799 ) );
  MUX2X1 \ashr_28_1/U317  ( .B(\ashr_28_1/n865 ), .A(\ashr_28_1/n881 ), .S(
        n1067), .Y(\ashr_28_1/n800 ) );
  MUX2X1 \ashr_28_1/U316  ( .B(\ashr_28_1/n866 ), .A(\ashr_28_1/n882 ), .S(
        n1067), .Y(\ashr_28_1/n801 ) );
  MUX2X1 \ashr_28_1/U315  ( .B(\ashr_28_1/n867 ), .A(\ashr_28_1/n883 ), .S(
        n1067), .Y(\ashr_28_1/n802 ) );
  MUX2X1 \ashr_28_1/U314  ( .B(\ashr_28_1/n868 ), .A(\ashr_28_1/n884 ), .S(
        n1067), .Y(\ashr_28_1/n803 ) );
  MUX2X1 \ashr_28_1/U313  ( .B(\ashr_28_1/n869 ), .A(\ashr_28_1/n885 ), .S(
        n1067), .Y(\ashr_28_1/n804 ) );
  MUX2X1 \ashr_28_1/U312  ( .B(\ashr_28_1/n870 ), .A(\ashr_28_1/n886 ), .S(
        n1067), .Y(\ashr_28_1/n805 ) );
  MUX2X1 \ashr_28_1/U311  ( .B(\ashr_28_1/n871 ), .A(\ashr_28_1/n887 ), .S(
        n1067), .Y(\ashr_28_1/n806 ) );
  MUX2X1 \ashr_28_1/U310  ( .B(\ashr_28_1/n872 ), .A(\ashr_28_1/n888 ), .S(
        n1067), .Y(\ashr_28_1/n807 ) );
  MUX2X1 \ashr_28_1/U309  ( .B(\ashr_28_1/n873 ), .A(\ashr_28_1/n889 ), .S(
        n1067), .Y(\ashr_28_1/n808 ) );
  MUX2X1 \ashr_28_1/U308  ( .B(\ashr_28_1/n874 ), .A(\ashr_28_1/n890 ), .S(
        n1067), .Y(\ashr_28_1/n809 ) );
  MUX2X1 \ashr_28_1/U307  ( .B(\ashr_28_1/n875 ), .A(\ashr_28_1/n891 ), .S(
        n1067), .Y(\ashr_28_1/n810 ) );
  MUX2X1 \ashr_28_1/U306  ( .B(\ashr_28_1/n876 ), .A(\ashr_28_1/n892 ), .S(
        n1067), .Y(\ashr_28_1/n811 ) );
  MUX2X1 \ashr_28_1/U305  ( .B(\ashr_28_1/n877 ), .A(\ashr_28_1/n893 ), .S(
        n1067), .Y(\ashr_28_1/n812 ) );
  MUX2X1 \ashr_28_1/U304  ( .B(\ashr_28_1/n878 ), .A(\ashr_28_1/n894 ), .S(
        n1067), .Y(\ashr_28_1/n813 ) );
  MUX2X1 \ashr_28_1/U303  ( .B(\ashr_28_1/n879 ), .A(\ashr_28_1/n895 ), .S(
        n1067), .Y(\ashr_28_1/n814 ) );
  MUX2X1 \ashr_28_1/U302  ( .B(\ashr_28_1/n880 ), .A(\ashr_28_1/n896 ), .S(
        n1067), .Y(\ashr_28_1/n815 ) );
  MUX2X1 \ashr_28_1/U301  ( .B(\ashr_28_1/n881 ), .A(\ashr_28_1/n897 ), .S(
        n1067), .Y(\ashr_28_1/n816 ) );
  MUX2X1 \ashr_28_1/U300  ( .B(\ashr_28_1/n882 ), .A(\ashr_28_1/n898 ), .S(
        n1067), .Y(\ashr_28_1/n817 ) );
  MUX2X1 \ashr_28_1/U299  ( .B(\ashr_28_1/n883 ), .A(\ashr_28_1/n899 ), .S(
        n1067), .Y(\ashr_28_1/n818 ) );
  MUX2X1 \ashr_28_1/U298  ( .B(\ashr_28_1/n884 ), .A(\ashr_28_1/n900 ), .S(
        n1067), .Y(\ashr_28_1/n819 ) );
  MUX2X1 \ashr_28_1/U297  ( .B(\ashr_28_1/n885 ), .A(\ashr_28_1/n901 ), .S(
        n1067), .Y(\ashr_28_1/n820 ) );
  MUX2X1 \ashr_28_1/U296  ( .B(\ashr_28_1/n886 ), .A(\ashr_28_1/n902 ), .S(
        n1067), .Y(\ashr_28_1/n821 ) );
  MUX2X1 \ashr_28_1/U295  ( .B(\ashr_28_1/n887 ), .A(\ashr_28_1/n903 ), .S(
        n1067), .Y(\ashr_28_1/n822 ) );
  MUX2X1 \ashr_28_1/U294  ( .B(\ashr_28_1/n888 ), .A(\ashr_28_1/n904 ), .S(
        n1067), .Y(\ashr_28_1/n823 ) );
  MUX2X1 \ashr_28_1/U293  ( .B(\ashr_28_1/n775 ), .A(\ashr_28_1/n783 ), .S(
        n1156), .Y(\ashr_28_1/n710 ) );
  MUX2X1 \ashr_28_1/U292  ( .B(\ashr_28_1/n776 ), .A(\ashr_28_1/n784 ), .S(
        n1156), .Y(\ashr_28_1/n711 ) );
  MUX2X1 \ashr_28_1/U291  ( .B(\ashr_28_1/n777 ), .A(\ashr_28_1/n785 ), .S(
        n1156), .Y(\ashr_28_1/n712 ) );
  MUX2X1 \ashr_28_1/U290  ( .B(\ashr_28_1/n778 ), .A(\ashr_28_1/n786 ), .S(
        n1156), .Y(\ashr_28_1/n713 ) );
  MUX2X1 \ashr_28_1/U289  ( .B(\ashr_28_1/n779 ), .A(\ashr_28_1/n787 ), .S(
        n1156), .Y(\ashr_28_1/n714 ) );
  MUX2X1 \ashr_28_1/U288  ( .B(\ashr_28_1/n780 ), .A(\ashr_28_1/n788 ), .S(
        n1156), .Y(\ashr_28_1/n715 ) );
  MUX2X1 \ashr_28_1/U287  ( .B(\ashr_28_1/n781 ), .A(\ashr_28_1/n789 ), .S(
        n1156), .Y(\ashr_28_1/n716 ) );
  MUX2X1 \ashr_28_1/U285  ( .B(\ashr_28_1/n783 ), .A(\ashr_28_1/n791 ), .S(
        n1156), .Y(\ashr_28_1/n718 ) );
  MUX2X1 \ashr_28_1/U284  ( .B(\ashr_28_1/n784 ), .A(\ashr_28_1/n792 ), .S(
        n1156), .Y(\ashr_28_1/n719 ) );
  MUX2X1 \ashr_28_1/U283  ( .B(\ashr_28_1/n785 ), .A(\ashr_28_1/n793 ), .S(
        n1156), .Y(\ashr_28_1/n720 ) );
  MUX2X1 \ashr_28_1/U282  ( .B(\ashr_28_1/n786 ), .A(\ashr_28_1/n794 ), .S(
        n1156), .Y(\ashr_28_1/n721 ) );
  MUX2X1 \ashr_28_1/U281  ( .B(\ashr_28_1/n787 ), .A(\ashr_28_1/n795 ), .S(
        n1155), .Y(\ashr_28_1/n722 ) );
  MUX2X1 \ashr_28_1/U280  ( .B(\ashr_28_1/n788 ), .A(\ashr_28_1/n796 ), .S(
        n1155), .Y(\ashr_28_1/n723 ) );
  MUX2X1 \ashr_28_1/U279  ( .B(\ashr_28_1/n789 ), .A(\ashr_28_1/n797 ), .S(
        n1155), .Y(\ashr_28_1/n724 ) );
  MUX2X1 \ashr_28_1/U278  ( .B(\ashr_28_1/n790 ), .A(\ashr_28_1/n798 ), .S(
        n1155), .Y(\ashr_28_1/n725 ) );
  MUX2X1 \ashr_28_1/U277  ( .B(\ashr_28_1/n791 ), .A(\ashr_28_1/n799 ), .S(
        n1155), .Y(\ashr_28_1/n726 ) );
  MUX2X1 \ashr_28_1/U276  ( .B(\ashr_28_1/n792 ), .A(\ashr_28_1/n800 ), .S(
        n1155), .Y(\ashr_28_1/n727 ) );
  MUX2X1 \ashr_28_1/U275  ( .B(\ashr_28_1/n793 ), .A(\ashr_28_1/n801 ), .S(
        n1155), .Y(\ashr_28_1/n728 ) );
  MUX2X1 \ashr_28_1/U274  ( .B(\ashr_28_1/n794 ), .A(\ashr_28_1/n802 ), .S(
        n1155), .Y(\ashr_28_1/n729 ) );
  MUX2X1 \ashr_28_1/U273  ( .B(\ashr_28_1/n795 ), .A(\ashr_28_1/n803 ), .S(
        n1155), .Y(\ashr_28_1/n730 ) );
  MUX2X1 \ashr_28_1/U272  ( .B(\ashr_28_1/n796 ), .A(\ashr_28_1/n804 ), .S(
        n1155), .Y(\ashr_28_1/n731 ) );
  MUX2X1 \ashr_28_1/U271  ( .B(\ashr_28_1/n797 ), .A(\ashr_28_1/n805 ), .S(
        n1155), .Y(\ashr_28_1/n732 ) );
  MUX2X1 \ashr_28_1/U270  ( .B(\ashr_28_1/n798 ), .A(\ashr_28_1/n806 ), .S(
        n1155), .Y(\ashr_28_1/n733 ) );
  MUX2X1 \ashr_28_1/U269  ( .B(\ashr_28_1/n799 ), .A(\ashr_28_1/n807 ), .S(
        n1155), .Y(\ashr_28_1/n734 ) );
  MUX2X1 \ashr_28_1/U268  ( .B(\ashr_28_1/n800 ), .A(\ashr_28_1/n808 ), .S(
        n1155), .Y(\ashr_28_1/n735 ) );
  MUX2X1 \ashr_28_1/U267  ( .B(\ashr_28_1/n801 ), .A(\ashr_28_1/n809 ), .S(
        n1155), .Y(\ashr_28_1/n736 ) );
  MUX2X1 \ashr_28_1/U266  ( .B(\ashr_28_1/n802 ), .A(\ashr_28_1/n810 ), .S(
        n1155), .Y(\ashr_28_1/n737 ) );
  MUX2X1 \ashr_28_1/U265  ( .B(\ashr_28_1/n803 ), .A(\ashr_28_1/n811 ), .S(
        n1155), .Y(\ashr_28_1/n738 ) );
  MUX2X1 \ashr_28_1/U264  ( .B(\ashr_28_1/n804 ), .A(\ashr_28_1/n812 ), .S(
        n1155), .Y(\ashr_28_1/n739 ) );
  MUX2X1 \ashr_28_1/U263  ( .B(\ashr_28_1/n805 ), .A(\ashr_28_1/n813 ), .S(
        n1155), .Y(\ashr_28_1/n740 ) );
  MUX2X1 \ashr_28_1/U262  ( .B(\ashr_28_1/n806 ), .A(\ashr_28_1/n814 ), .S(
        n1155), .Y(\ashr_28_1/n741 ) );
  MUX2X1 \ashr_28_1/U261  ( .B(\ashr_28_1/n807 ), .A(\ashr_28_1/n815 ), .S(
        n1155), .Y(\ashr_28_1/n742 ) );
  MUX2X1 \ashr_28_1/U260  ( .B(\ashr_28_1/n808 ), .A(\ashr_28_1/n816 ), .S(
        n1155), .Y(\ashr_28_1/n743 ) );
  MUX2X1 \ashr_28_1/U259  ( .B(\ashr_28_1/n809 ), .A(\ashr_28_1/n817 ), .S(
        n1155), .Y(\ashr_28_1/n744 ) );
  MUX2X1 \ashr_28_1/U258  ( .B(\ashr_28_1/n810 ), .A(\ashr_28_1/n818 ), .S(
        n1155), .Y(\ashr_28_1/n745 ) );
  MUX2X1 \ashr_28_1/U257  ( .B(\ashr_28_1/n811 ), .A(\ashr_28_1/n819 ), .S(
        n1155), .Y(\ashr_28_1/n746 ) );
  MUX2X1 \ashr_28_1/U256  ( .B(\ashr_28_1/n812 ), .A(\ashr_28_1/n820 ), .S(
        n1155), .Y(\ashr_28_1/n747 ) );
  MUX2X1 \ashr_28_1/U255  ( .B(\ashr_28_1/n813 ), .A(\ashr_28_1/n821 ), .S(
        n1155), .Y(\ashr_28_1/n748 ) );
  MUX2X1 \ashr_28_1/U254  ( .B(\ashr_28_1/n814 ), .A(\ashr_28_1/n822 ), .S(
        n1155), .Y(\ashr_28_1/n749 ) );
  MUX2X1 \ashr_28_1/U253  ( .B(\ashr_28_1/n815 ), .A(\ashr_28_1/n823 ), .S(
        n1155), .Y(\ashr_28_1/n750 ) );
  MUX2X1 \ashr_28_1/U252  ( .B(\ashr_28_1/n816 ), .A(\ashr_28_1/n824 ), .S(
        n1155), .Y(\ashr_28_1/n751 ) );
  MUX2X1 \ashr_28_1/U251  ( .B(\ashr_28_1/n817 ), .A(\ashr_28_1/n825 ), .S(
        n1155), .Y(\ashr_28_1/n752 ) );
  MUX2X1 \ashr_28_1/U250  ( .B(\ashr_28_1/n818 ), .A(\ashr_28_1/n826 ), .S(
        n1155), .Y(\ashr_28_1/n753 ) );
  MUX2X1 \ashr_28_1/U249  ( .B(\ashr_28_1/n819 ), .A(\ashr_28_1/n827 ), .S(
        n1155), .Y(\ashr_28_1/n754 ) );
  MUX2X1 \ashr_28_1/U248  ( .B(\ashr_28_1/n820 ), .A(\ashr_28_1/n828 ), .S(
        n1155), .Y(\ashr_28_1/n755 ) );
  MUX2X1 \ashr_28_1/U247  ( .B(\ashr_28_1/n821 ), .A(\ashr_28_1/n829 ), .S(
        n1155), .Y(\ashr_28_1/n756 ) );
  MUX2X1 \ashr_28_1/U246  ( .B(\ashr_28_1/n822 ), .A(\ashr_28_1/n830 ), .S(
        n1155), .Y(\ashr_28_1/n757 ) );
  MUX2X1 \ashr_28_1/U245  ( .B(\ashr_28_1/n823 ), .A(\ashr_28_1/n831 ), .S(
        n1156), .Y(\ashr_28_1/n758 ) );
  MUX2X1 \ashr_28_1/U244  ( .B(\ashr_28_1/n824 ), .A(\ashr_28_1/n832 ), .S(
        n1155), .Y(\ashr_28_1/n759 ) );
  MUX2X1 \ashr_28_1/U243  ( .B(\ashr_28_1/n825 ), .A(\ashr_28_1/n833 ), .S(
        n1156), .Y(\ashr_28_1/n760 ) );
  MUX2X1 \ashr_28_1/U242  ( .B(\ashr_28_1/n826 ), .A(\ashr_28_1/n834 ), .S(
        n1155), .Y(\ashr_28_1/n761 ) );
  MUX2X1 \ashr_28_1/U241  ( .B(\ashr_28_1/n827 ), .A(\ashr_28_1/n835 ), .S(
        n1156), .Y(\ashr_28_1/n762 ) );
  MUX2X1 \ashr_28_1/U240  ( .B(\ashr_28_1/n828 ), .A(\ashr_28_1/n836 ), .S(
        n1155), .Y(\ashr_28_1/n763 ) );
  MUX2X1 \ashr_28_1/U239  ( .B(\ashr_28_1/n829 ), .A(\ashr_28_1/n837 ), .S(
        n1156), .Y(\ashr_28_1/n764 ) );
  MUX2X1 \ashr_28_1/U238  ( .B(\ashr_28_1/n830 ), .A(\ashr_28_1/n838 ), .S(
        n1155), .Y(\ashr_28_1/n765 ) );
  MUX2X1 \ashr_28_1/U237  ( .B(\ashr_28_1/n831 ), .A(\ashr_28_1/n839 ), .S(
        n1155), .Y(\ashr_28_1/n766 ) );
  NOR2X1 \ashr_28_1/U236  ( .A(n1156), .B(\ashr_28_1/n832 ), .Y(
        \ashr_28_1/n767 ) );
  NOR2X1 \ashr_28_1/U235  ( .A(n1155), .B(\ashr_28_1/n833 ), .Y(
        \ashr_28_1/n768 ) );
  NOR2X1 \ashr_28_1/U234  ( .A(n1156), .B(\ashr_28_1/n834 ), .Y(
        \ashr_28_1/n769 ) );
  NOR2X1 \ashr_28_1/U233  ( .A(n1155), .B(\ashr_28_1/n835 ), .Y(
        \ashr_28_1/n770 ) );
  NOR2X1 \ashr_28_1/U232  ( .A(n1155), .B(\ashr_28_1/n836 ), .Y(
        \ashr_28_1/n771 ) );
  NOR2X1 \ashr_28_1/U231  ( .A(n1156), .B(\ashr_28_1/n837 ), .Y(
        \ashr_28_1/n772 ) );
  NOR2X1 \ashr_28_1/U230  ( .A(n1155), .B(\ashr_28_1/n838 ), .Y(
        \ashr_28_1/n773 ) );
  NOR2X1 \ashr_28_1/U229  ( .A(n1155), .B(\ashr_28_1/n839 ), .Y(
        \ashr_28_1/n774 ) );
  MUX2X1 \ashr_28_1/U228  ( .B(\ashr_28_1/n710 ), .A(\ashr_28_1/n714 ), .S(
        n1160), .Y(\ashr_28_1/n645 ) );
  MUX2X1 \ashr_28_1/U227  ( .B(\ashr_28_1/n711 ), .A(\ashr_28_1/n715 ), .S(
        n1158), .Y(\ashr_28_1/n646 ) );
  MUX2X1 \ashr_28_1/U226  ( .B(\ashr_28_1/n712 ), .A(\ashr_28_1/n716 ), .S(
        n1158), .Y(\ashr_28_1/n647 ) );
  MUX2X1 \ashr_28_1/U225  ( .B(\ashr_28_1/n713 ), .A(\ashr_28_1/n717 ), .S(
        n1158), .Y(\ashr_28_1/n648 ) );
  MUX2X1 \ashr_28_1/U224  ( .B(\ashr_28_1/n714 ), .A(\ashr_28_1/n718 ), .S(
        n1158), .Y(\ashr_28_1/n649 ) );
  MUX2X1 \ashr_28_1/U223  ( .B(\ashr_28_1/n715 ), .A(\ashr_28_1/n719 ), .S(
        n1158), .Y(\ashr_28_1/n650 ) );
  MUX2X1 \ashr_28_1/U222  ( .B(\ashr_28_1/n716 ), .A(\ashr_28_1/n720 ), .S(
        n1158), .Y(\ashr_28_1/n651 ) );
  MUX2X1 \ashr_28_1/U221  ( .B(\ashr_28_1/n717 ), .A(\ashr_28_1/n721 ), .S(
        n1158), .Y(\ashr_28_1/n652 ) );
  MUX2X1 \ashr_28_1/U220  ( .B(\ashr_28_1/n718 ), .A(\ashr_28_1/n722 ), .S(
        n1158), .Y(\ashr_28_1/n653 ) );
  MUX2X1 \ashr_28_1/U219  ( .B(\ashr_28_1/n719 ), .A(\ashr_28_1/n723 ), .S(
        n1158), .Y(\ashr_28_1/n654 ) );
  MUX2X1 \ashr_28_1/U218  ( .B(\ashr_28_1/n720 ), .A(\ashr_28_1/n724 ), .S(
        n1158), .Y(\ashr_28_1/n655 ) );
  MUX2X1 \ashr_28_1/U217  ( .B(\ashr_28_1/n721 ), .A(\ashr_28_1/n725 ), .S(
        n1158), .Y(\ashr_28_1/n656 ) );
  MUX2X1 \ashr_28_1/U216  ( .B(\ashr_28_1/n722 ), .A(\ashr_28_1/n726 ), .S(
        n1158), .Y(\ashr_28_1/n657 ) );
  MUX2X1 \ashr_28_1/U215  ( .B(\ashr_28_1/n723 ), .A(\ashr_28_1/n727 ), .S(
        n1159), .Y(\ashr_28_1/n658 ) );
  MUX2X1 \ashr_28_1/U214  ( .B(\ashr_28_1/n724 ), .A(\ashr_28_1/n728 ), .S(
        n1159), .Y(\ashr_28_1/n659 ) );
  MUX2X1 \ashr_28_1/U213  ( .B(\ashr_28_1/n725 ), .A(\ashr_28_1/n729 ), .S(
        n1160), .Y(\ashr_28_1/n660 ) );
  MUX2X1 \ashr_28_1/U212  ( .B(\ashr_28_1/n726 ), .A(\ashr_28_1/n730 ), .S(
        n1160), .Y(\ashr_28_1/n661 ) );
  MUX2X1 \ashr_28_1/U211  ( .B(\ashr_28_1/n727 ), .A(\ashr_28_1/n731 ), .S(
        n1160), .Y(\ashr_28_1/n662 ) );
  MUX2X1 \ashr_28_1/U210  ( .B(\ashr_28_1/n728 ), .A(\ashr_28_1/n732 ), .S(
        n1159), .Y(\ashr_28_1/n663 ) );
  MUX2X1 \ashr_28_1/U209  ( .B(\ashr_28_1/n729 ), .A(\ashr_28_1/n733 ), .S(
        n1159), .Y(\ashr_28_1/n664 ) );
  MUX2X1 \ashr_28_1/U208  ( .B(\ashr_28_1/n730 ), .A(\ashr_28_1/n734 ), .S(
        n1159), .Y(\ashr_28_1/n665 ) );
  MUX2X1 \ashr_28_1/U207  ( .B(\ashr_28_1/n731 ), .A(\ashr_28_1/n735 ), .S(
        n1160), .Y(\ashr_28_1/n666 ) );
  MUX2X1 \ashr_28_1/U206  ( .B(\ashr_28_1/n732 ), .A(\ashr_28_1/n736 ), .S(
        n1160), .Y(\ashr_28_1/n667 ) );
  MUX2X1 \ashr_28_1/U205  ( .B(\ashr_28_1/n733 ), .A(\ashr_28_1/n737 ), .S(
        n1159), .Y(\ashr_28_1/n668 ) );
  MUX2X1 \ashr_28_1/U204  ( .B(\ashr_28_1/n734 ), .A(\ashr_28_1/n738 ), .S(
        n1159), .Y(\ashr_28_1/n669 ) );
  MUX2X1 \ashr_28_1/U203  ( .B(\ashr_28_1/n735 ), .A(\ashr_28_1/n739 ), .S(
        n1159), .Y(\ashr_28_1/n670 ) );
  MUX2X1 \ashr_28_1/U202  ( .B(\ashr_28_1/n736 ), .A(\ashr_28_1/n740 ), .S(
        n1159), .Y(\ashr_28_1/n671 ) );
  MUX2X1 \ashr_28_1/U201  ( .B(\ashr_28_1/n737 ), .A(\ashr_28_1/n741 ), .S(
        n1159), .Y(\ashr_28_1/n672 ) );
  MUX2X1 \ashr_28_1/U200  ( .B(\ashr_28_1/n738 ), .A(\ashr_28_1/n742 ), .S(
        n1159), .Y(\ashr_28_1/n673 ) );
  MUX2X1 \ashr_28_1/U109  ( .B(\ashr_28_1/n739 ), .A(\ashr_28_1/n743 ), .S(
        n1159), .Y(\ashr_28_1/n674 ) );
  MUX2X1 \ashr_28_1/U108  ( .B(\ashr_28_1/n740 ), .A(\ashr_28_1/n744 ), .S(
        n1159), .Y(\ashr_28_1/n675 ) );
  MUX2X1 \ashr_28_1/U107  ( .B(\ashr_28_1/n741 ), .A(\ashr_28_1/n745 ), .S(
        n1159), .Y(\ashr_28_1/n676 ) );
  MUX2X1 \ashr_28_1/U106  ( .B(\ashr_28_1/n742 ), .A(\ashr_28_1/n746 ), .S(
        n1159), .Y(\ashr_28_1/n677 ) );
  MUX2X1 \ashr_28_1/U105  ( .B(\ashr_28_1/n743 ), .A(\ashr_28_1/n747 ), .S(
        n1159), .Y(\ashr_28_1/n678 ) );
  MUX2X1 \ashr_28_1/U104  ( .B(\ashr_28_1/n744 ), .A(\ashr_28_1/n748 ), .S(
        n1159), .Y(\ashr_28_1/n679 ) );
  MUX2X1 \ashr_28_1/U103  ( .B(\ashr_28_1/n745 ), .A(\ashr_28_1/n749 ), .S(
        n1159), .Y(\ashr_28_1/n680 ) );
  MUX2X1 \ashr_28_1/U102  ( .B(\ashr_28_1/n746 ), .A(\ashr_28_1/n750 ), .S(
        n1159), .Y(\ashr_28_1/n681 ) );
  MUX2X1 \ashr_28_1/U101  ( .B(\ashr_28_1/n747 ), .A(\ashr_28_1/n751 ), .S(
        n1160), .Y(\ashr_28_1/n682 ) );
  MUX2X1 \ashr_28_1/U100  ( .B(\ashr_28_1/n748 ), .A(\ashr_28_1/n752 ), .S(
        n1160), .Y(\ashr_28_1/n683 ) );
  MUX2X1 \ashr_28_1/U99  ( .B(\ashr_28_1/n749 ), .A(\ashr_28_1/n753 ), .S(
        n1160), .Y(\ashr_28_1/n684 ) );
  MUX2X1 \ashr_28_1/U98  ( .B(\ashr_28_1/n750 ), .A(\ashr_28_1/n754 ), .S(
        n1160), .Y(\ashr_28_1/n685 ) );
  MUX2X1 \ashr_28_1/U97  ( .B(\ashr_28_1/n751 ), .A(\ashr_28_1/n755 ), .S(
        n1160), .Y(\ashr_28_1/n686 ) );
  MUX2X1 \ashr_28_1/U96  ( .B(\ashr_28_1/n752 ), .A(\ashr_28_1/n756 ), .S(
        n1160), .Y(\ashr_28_1/n687 ) );
  MUX2X1 \ashr_28_1/U95  ( .B(\ashr_28_1/n753 ), .A(\ashr_28_1/n757 ), .S(
        n1160), .Y(\ashr_28_1/n688 ) );
  MUX2X1 \ashr_28_1/U94  ( .B(\ashr_28_1/n754 ), .A(\ashr_28_1/n758 ), .S(
        n1160), .Y(\ashr_28_1/n689 ) );
  MUX2X1 \ashr_28_1/U93  ( .B(\ashr_28_1/n755 ), .A(\ashr_28_1/n759 ), .S(
        n1160), .Y(\ashr_28_1/n690 ) );
  MUX2X1 \ashr_28_1/U92  ( .B(\ashr_28_1/n756 ), .A(\ashr_28_1/n760 ), .S(
        n1160), .Y(\ashr_28_1/n691 ) );
  MUX2X1 \ashr_28_1/U91  ( .B(\ashr_28_1/n757 ), .A(\ashr_28_1/n761 ), .S(
        n1160), .Y(\ashr_28_1/n692 ) );
  MUX2X1 \ashr_28_1/U90  ( .B(\ashr_28_1/n758 ), .A(\ashr_28_1/n762 ), .S(
        n1160), .Y(\ashr_28_1/n693 ) );
  MUX2X1 \ashr_28_1/U89  ( .B(\ashr_28_1/n759 ), .A(\ashr_28_1/n763 ), .S(
        n1160), .Y(\ashr_28_1/n694 ) );
  MUX2X1 \ashr_28_1/U88  ( .B(\ashr_28_1/n760 ), .A(\ashr_28_1/n764 ), .S(
        n1158), .Y(\ashr_28_1/n695 ) );
  MUX2X1 \ashr_28_1/U87  ( .B(\ashr_28_1/n761 ), .A(\ashr_28_1/n765 ), .S(
        n1159), .Y(\ashr_28_1/n696 ) );
  MUX2X1 \ashr_28_1/U86  ( .B(\ashr_28_1/n762 ), .A(\ashr_28_1/n766 ), .S(
        n1158), .Y(\ashr_28_1/n697 ) );
  MUX2X1 \ashr_28_1/U85  ( .B(\ashr_28_1/n763 ), .A(\ashr_28_1/n767 ), .S(
        n1160), .Y(\ashr_28_1/n698 ) );
  MUX2X1 \ashr_28_1/U84  ( .B(\ashr_28_1/n764 ), .A(\ashr_28_1/n768 ), .S(
        n1159), .Y(\ashr_28_1/n699 ) );
  MUX2X1 \ashr_28_1/U83  ( .B(\ashr_28_1/n765 ), .A(\ashr_28_1/n769 ), .S(
        n1158), .Y(\ashr_28_1/n700 ) );
  MUX2X1 \ashr_28_1/U82  ( .B(\ashr_28_1/n766 ), .A(\ashr_28_1/n770 ), .S(
        n1158), .Y(\ashr_28_1/n701 ) );
  MUX2X1 \ashr_28_1/U81  ( .B(\ashr_28_1/n767 ), .A(\ashr_28_1/n771 ), .S(
        n1160), .Y(\ashr_28_1/n702 ) );
  MUX2X1 \ashr_28_1/U80  ( .B(\ashr_28_1/n768 ), .A(\ashr_28_1/n772 ), .S(
        n1158), .Y(\ashr_28_1/n703 ) );
  MUX2X1 \ashr_28_1/U79  ( .B(\ashr_28_1/n769 ), .A(\ashr_28_1/n773 ), .S(
        n1159), .Y(\ashr_28_1/n704 ) );
  MUX2X1 \ashr_28_1/U78  ( .B(\ashr_28_1/n770 ), .A(\ashr_28_1/n774 ), .S(
        n1160), .Y(\ashr_28_1/n705 ) );
  MUX2X1 \ashr_28_1/U77  ( .B(\ashr_28_1/n645 ), .A(\ashr_28_1/n646 ), .S(
        n1166), .Y(\ashr_28_1/n580 ) );
  MUX2X1 \ashr_28_1/U76  ( .B(\ashr_28_1/n646 ), .A(\ashr_28_1/n647 ), .S(
        n1166), .Y(\ashr_28_1/n581 ) );
  MUX2X1 \ashr_28_1/U75  ( .B(\ashr_28_1/n647 ), .A(\ashr_28_1/n648 ), .S(
        n1166), .Y(\ashr_28_1/n582 ) );
  MUX2X1 \ashr_28_1/U73  ( .B(\ashr_28_1/n649 ), .A(\ashr_28_1/n650 ), .S(
        n1166), .Y(\ashr_28_1/n584 ) );
  MUX2X1 \ashr_28_1/U72  ( .B(\ashr_28_1/n650 ), .A(\ashr_28_1/n651 ), .S(
        n1166), .Y(\ashr_28_1/n585 ) );
  MUX2X1 \ashr_28_1/U71  ( .B(\ashr_28_1/n651 ), .A(\ashr_28_1/n652 ), .S(
        n1166), .Y(\ashr_28_1/n586 ) );
  MUX2X1 \ashr_28_1/U70  ( .B(\ashr_28_1/n652 ), .A(\ashr_28_1/n653 ), .S(
        n1166), .Y(\ashr_28_1/n587 ) );
  MUX2X1 \ashr_28_1/U69  ( .B(\ashr_28_1/n653 ), .A(\ashr_28_1/n654 ), .S(
        n1166), .Y(\ashr_28_1/n588 ) );
  MUX2X1 \ashr_28_1/U68  ( .B(\ashr_28_1/n654 ), .A(\ashr_28_1/n655 ), .S(
        n1166), .Y(\ashr_28_1/n589 ) );
  MUX2X1 \ashr_28_1/U67  ( .B(\ashr_28_1/n655 ), .A(\ashr_28_1/n656 ), .S(
        n1166), .Y(\ashr_28_1/n590 ) );
  MUX2X1 \ashr_28_1/U66  ( .B(\ashr_28_1/n656 ), .A(\ashr_28_1/n657 ), .S(
        n1166), .Y(\ashr_28_1/n591 ) );
  MUX2X1 \ashr_28_1/U65  ( .B(\ashr_28_1/n657 ), .A(\ashr_28_1/n658 ), .S(
        n1166), .Y(\ashr_28_1/n592 ) );
  MUX2X1 \ashr_28_1/U64  ( .B(\ashr_28_1/n658 ), .A(\ashr_28_1/n659 ), .S(
        n1166), .Y(\ashr_28_1/n593 ) );
  MUX2X1 \ashr_28_1/U63  ( .B(\ashr_28_1/n659 ), .A(\ashr_28_1/n660 ), .S(
        n1166), .Y(\ashr_28_1/n594 ) );
  MUX2X1 \ashr_28_1/U62  ( .B(\ashr_28_1/n660 ), .A(\ashr_28_1/n661 ), .S(
        n1166), .Y(\ashr_28_1/n595 ) );
  MUX2X1 \ashr_28_1/U61  ( .B(\ashr_28_1/n661 ), .A(\ashr_28_1/n662 ), .S(
        n1166), .Y(\ashr_28_1/n596 ) );
  MUX2X1 \ashr_28_1/U60  ( .B(\ashr_28_1/n662 ), .A(\ashr_28_1/n663 ), .S(
        n1166), .Y(\ashr_28_1/n597 ) );
  MUX2X1 \ashr_28_1/U59  ( .B(\ashr_28_1/n663 ), .A(\ashr_28_1/n664 ), .S(
        n1166), .Y(\ashr_28_1/n598 ) );
  MUX2X1 \ashr_28_1/U58  ( .B(\ashr_28_1/n664 ), .A(\ashr_28_1/n665 ), .S(
        n1166), .Y(\ashr_28_1/n599 ) );
  MUX2X1 \ashr_28_1/U57  ( .B(\ashr_28_1/n665 ), .A(\ashr_28_1/n666 ), .S(
        n1166), .Y(\ashr_28_1/n600 ) );
  MUX2X1 \ashr_28_1/U56  ( .B(\ashr_28_1/n666 ), .A(\ashr_28_1/n667 ), .S(
        n1166), .Y(\ashr_28_1/n601 ) );
  MUX2X1 \ashr_28_1/U55  ( .B(\ashr_28_1/n667 ), .A(\ashr_28_1/n668 ), .S(
        n1166), .Y(\ashr_28_1/n602 ) );
  MUX2X1 \ashr_28_1/U54  ( .B(\ashr_28_1/n668 ), .A(\ashr_28_1/n669 ), .S(
        n1166), .Y(\ashr_28_1/n603 ) );
  MUX2X1 \ashr_28_1/U53  ( .B(\ashr_28_1/n669 ), .A(\ashr_28_1/n670 ), .S(
        n1165), .Y(\ashr_28_1/n604 ) );
  MUX2X1 \ashr_28_1/U52  ( .B(\ashr_28_1/n670 ), .A(\ashr_28_1/n671 ), .S(
        n1165), .Y(\ashr_28_1/n605 ) );
  MUX2X1 \ashr_28_1/U51  ( .B(\ashr_28_1/n671 ), .A(\ashr_28_1/n672 ), .S(
        n1165), .Y(\ashr_28_1/n606 ) );
  MUX2X1 \ashr_28_1/U50  ( .B(\ashr_28_1/n672 ), .A(\ashr_28_1/n673 ), .S(
        n1165), .Y(\ashr_28_1/n607 ) );
  MUX2X1 \ashr_28_1/U49  ( .B(\ashr_28_1/n673 ), .A(\ashr_28_1/n674 ), .S(
        n1165), .Y(\ashr_28_1/n608 ) );
  MUX2X1 \ashr_28_1/U48  ( .B(\ashr_28_1/n674 ), .A(\ashr_28_1/n675 ), .S(
        n1165), .Y(\ashr_28_1/n609 ) );
  MUX2X1 \ashr_28_1/U47  ( .B(\ashr_28_1/n675 ), .A(\ashr_28_1/n676 ), .S(
        n1165), .Y(\ashr_28_1/n610 ) );
  MUX2X1 \ashr_28_1/U46  ( .B(\ashr_28_1/n676 ), .A(\ashr_28_1/n677 ), .S(
        n1165), .Y(\ashr_28_1/n611 ) );
  MUX2X1 \ashr_28_1/U45  ( .B(\ashr_28_1/n677 ), .A(\ashr_28_1/n678 ), .S(
        n1165), .Y(\ashr_28_1/n612 ) );
  MUX2X1 \ashr_28_1/U44  ( .B(\ashr_28_1/n678 ), .A(\ashr_28_1/n679 ), .S(
        n1165), .Y(\ashr_28_1/n613 ) );
  MUX2X1 \ashr_28_1/U43  ( .B(\ashr_28_1/n679 ), .A(\ashr_28_1/n680 ), .S(
        n1165), .Y(\ashr_28_1/n614 ) );
  MUX2X1 \ashr_28_1/U42  ( .B(\ashr_28_1/n680 ), .A(\ashr_28_1/n681 ), .S(
        n1165), .Y(\ashr_28_1/n615 ) );
  MUX2X1 \ashr_28_1/U41  ( .B(\ashr_28_1/n681 ), .A(\ashr_28_1/n682 ), .S(
        n1165), .Y(\ashr_28_1/n616 ) );
  MUX2X1 \ashr_28_1/U40  ( .B(\ashr_28_1/n682 ), .A(\ashr_28_1/n683 ), .S(
        n1165), .Y(\ashr_28_1/n617 ) );
  MUX2X1 \ashr_28_1/U39  ( .B(\ashr_28_1/n683 ), .A(\ashr_28_1/n684 ), .S(
        n1165), .Y(\ashr_28_1/n618 ) );
  MUX2X1 \ashr_28_1/U38  ( .B(\ashr_28_1/n684 ), .A(\ashr_28_1/n685 ), .S(
        n1165), .Y(\ashr_28_1/n619 ) );
  MUX2X1 \ashr_28_1/U37  ( .B(\ashr_28_1/n685 ), .A(\ashr_28_1/n686 ), .S(
        n1165), .Y(\ashr_28_1/n620 ) );
  MUX2X1 \ashr_28_1/U36  ( .B(\ashr_28_1/n686 ), .A(\ashr_28_1/n687 ), .S(
        n1165), .Y(\ashr_28_1/n621 ) );
  MUX2X1 \ashr_28_1/U35  ( .B(\ashr_28_1/n687 ), .A(\ashr_28_1/n688 ), .S(
        n1165), .Y(\ashr_28_1/n622 ) );
  MUX2X1 \ashr_28_1/U34  ( .B(\ashr_28_1/n688 ), .A(\ashr_28_1/n689 ), .S(
        n1165), .Y(\ashr_28_1/n623 ) );
  MUX2X1 \ashr_28_1/U33  ( .B(\ashr_28_1/n689 ), .A(\ashr_28_1/n690 ), .S(
        n1165), .Y(\ashr_28_1/n624 ) );
  MUX2X1 \ashr_28_1/U32  ( .B(\ashr_28_1/n690 ), .A(\ashr_28_1/n691 ), .S(
        n1165), .Y(\ashr_28_1/n625 ) );
  MUX2X1 \ashr_28_1/U31  ( .B(\ashr_28_1/n691 ), .A(\ashr_28_1/n692 ), .S(
        n1165), .Y(\ashr_28_1/n626 ) );
  MUX2X1 \ashr_28_1/U30  ( .B(\ashr_28_1/n692 ), .A(\ashr_28_1/n693 ), .S(
        n1165), .Y(\ashr_28_1/n627 ) );
  MUX2X1 \ashr_28_1/U29  ( .B(\ashr_28_1/n693 ), .A(\ashr_28_1/n694 ), .S(
        n1166), .Y(\ashr_28_1/n628 ) );
  MUX2X1 \ashr_28_1/U28  ( .B(\ashr_28_1/n694 ), .A(\ashr_28_1/n695 ), .S(
        n1166), .Y(\ashr_28_1/n629 ) );
  MUX2X1 \ashr_28_1/U27  ( .B(\ashr_28_1/n695 ), .A(\ashr_28_1/n696 ), .S(
        n1165), .Y(\ashr_28_1/n630 ) );
  MUX2X1 \ashr_28_1/U26  ( .B(\ashr_28_1/n696 ), .A(\ashr_28_1/n697 ), .S(
        n1166), .Y(\ashr_28_1/n631 ) );
  MUX2X1 \ashr_28_1/U25  ( .B(\ashr_28_1/n697 ), .A(\ashr_28_1/n698 ), .S(
        n1166), .Y(\ashr_28_1/n632 ) );
  MUX2X1 \ashr_28_1/U24  ( .B(\ashr_28_1/n698 ), .A(\ashr_28_1/n699 ), .S(
        n1166), .Y(\ashr_28_1/n633 ) );
  MUX2X1 \ashr_28_1/U23  ( .B(\ashr_28_1/n699 ), .A(\ashr_28_1/n700 ), .S(
        n1165), .Y(\ashr_28_1/n634 ) );
  MUX2X1 \ashr_28_1/U22  ( .B(\ashr_28_1/n700 ), .A(\ashr_28_1/n701 ), .S(
        n1166), .Y(\ashr_28_1/n635 ) );
  MUX2X1 \ashr_28_1/U20  ( .B(\ashr_28_1/n701 ), .A(\ashr_28_1/n702 ), .S(
        h2[0]), .Y(\ashr_28_1/n636 ) );
  MUX2X1 \ashr_28_1/U10  ( .B(\ashr_28_1/n702 ), .A(\ashr_28_1/n703 ), .S(
        h2[0]), .Y(\ashr_28_1/n637 ) );
  MUX2X1 \ashr_28_1/U9  ( .B(\ashr_28_1/n703 ), .A(\ashr_28_1/n704 ), .S(n1166), .Y(\ashr_28_1/n638 ) );
  MUX2X1 \ashr_28_1/U8  ( .B(\ashr_28_1/n704 ), .A(\ashr_28_1/n705 ), .S(h2[0]), .Y(\ashr_28_1/n639 ) );
  MUX2X1 \ashr_28_1/U7  ( .B(\ashr_28_1/n705 ), .A(\ashr_28_1/n706 ), .S(n1165), .Y(\ashr_28_1/n640 ) );
  MUX2X1 \ashr_28_1/U6  ( .B(\ashr_28_1/n706 ), .A(\ashr_28_1/n707 ), .S(n1166), .Y(\ashr_28_1/n641 ) );
  MUX2X1 \ashr_28_1/U5  ( .B(\ashr_28_1/n707 ), .A(\ashr_28_1/n708 ), .S(n1165), .Y(\ashr_28_1/n642 ) );
  MUX2X1 \ashr_28_1/U4  ( .B(\ashr_28_1/n708 ), .A(\ashr_28_1/n709 ), .S(h2[0]), .Y(\ashr_28_1/n643 ) );
  NOR2X1 \ashr_28_1/U3  ( .A(n1165), .B(\ashr_28_1/n709 ), .Y(\ashr_28_1/n644 ) );
  NAND2X1 \DP_OP_19_294_9081/U584  ( .A(\DP_OP_19_294_9081/n653 ), .B(
        \DP_OP_19_294_9081/n589 ), .Y(\DP_OP_19_294_9081/n457 ) );
  NAND2X1 \DP_OP_19_294_9081/U579  ( .A(\C2/Z_1 ), .B(\DP_OP_19_294_9081/n654 ), .Y(\DP_OP_19_294_9081/n455 ) );
  NOR2X1 \DP_OP_19_294_9081/U578  ( .A(\C2/Z_1 ), .B(\DP_OP_19_294_9081/n654 ), 
        .Y(\DP_OP_19_294_9081/n454 ) );
  NAND2X1 \DP_OP_19_294_9081/U576  ( .A(\DP_OP_19_294_9081/n455 ), .B(
        \DP_OP_19_294_9081/n519 ), .Y(\DP_OP_19_294_9081/n67 ) );
  OAI21X1 \DP_OP_19_294_9081/U575  ( .A(\DP_OP_19_294_9081/n457 ), .B(
        \DP_OP_19_294_9081/n454 ), .C(\DP_OP_19_294_9081/n455 ), .Y(
        \DP_OP_19_294_9081/n453 ) );
  XOR2X1 \DP_OP_19_294_9081/U573  ( .A(\DP_OP_19_294_9081/n457 ), .B(
        \DP_OP_19_294_9081/n67 ), .Y(\C2/DATA3_1 ) );
  NAND2X1 \DP_OP_19_294_9081/U572  ( .A(\C2/Z_2 ), .B(\DP_OP_19_294_9081/n655 ), .Y(\DP_OP_19_294_9081/n451 ) );
  NOR2X1 \DP_OP_19_294_9081/U571  ( .A(\C2/Z_2 ), .B(\DP_OP_19_294_9081/n655 ), 
        .Y(\DP_OP_19_294_9081/n450 ) );
  OAI21X1 \DP_OP_19_294_9081/U568  ( .A(\DP_OP_19_294_9081/n450 ), .B(
        \DP_OP_19_294_9081/n452 ), .C(\DP_OP_19_294_9081/n451 ), .Y(
        \DP_OP_19_294_9081/n449 ) );
  NAND2X1 \DP_OP_19_294_9081/U566  ( .A(\C2/Z_3 ), .B(\DP_OP_19_294_9081/n656 ), .Y(\DP_OP_19_294_9081/n448 ) );
  NOR2X1 \DP_OP_19_294_9081/U565  ( .A(\C2/Z_3 ), .B(\DP_OP_19_294_9081/n656 ), 
        .Y(\DP_OP_19_294_9081/n447 ) );
  NAND2X1 \DP_OP_19_294_9081/U557  ( .A(\C2/Z_4 ), .B(\DP_OP_19_294_9081/n657 ), .Y(\DP_OP_19_294_9081/n442 ) );
  NOR2X1 \DP_OP_19_294_9081/U556  ( .A(\C2/Z_4 ), .B(\DP_OP_19_294_9081/n657 ), 
        .Y(\DP_OP_19_294_9081/n441 ) );
  NAND2X1 \DP_OP_19_294_9081/U554  ( .A(\DP_OP_19_294_9081/n442 ), .B(
        \DP_OP_19_294_9081/n516 ), .Y(\DP_OP_19_294_9081/n64 ) );
  AOI21X1 \DP_OP_19_294_9081/U551  ( .A(\DP_OP_19_294_9081/n516 ), .B(
        \DP_OP_19_294_9081/n443 ), .C(\DP_OP_19_294_9081/n440 ), .Y(
        \DP_OP_19_294_9081/n438 ) );
  NAND2X1 \DP_OP_19_294_9081/U549  ( .A(\C2/Z_5 ), .B(\DP_OP_19_294_9081/n658 ), .Y(\DP_OP_19_294_9081/n437 ) );
  NOR2X1 \DP_OP_19_294_9081/U548  ( .A(\C2/Z_5 ), .B(\DP_OP_19_294_9081/n658 ), 
        .Y(\DP_OP_19_294_9081/n436 ) );
  NAND2X1 \DP_OP_19_294_9081/U546  ( .A(\DP_OP_19_294_9081/n437 ), .B(
        \DP_OP_19_294_9081/n515 ), .Y(\DP_OP_19_294_9081/n63 ) );
  OAI21X1 \DP_OP_19_294_9081/U545  ( .A(\DP_OP_19_294_9081/n442 ), .B(
        \DP_OP_19_294_9081/n436 ), .C(\DP_OP_19_294_9081/n437 ), .Y(
        \DP_OP_19_294_9081/n435 ) );
  NOR2X1 \DP_OP_19_294_9081/U544  ( .A(\DP_OP_19_294_9081/n436 ), .B(
        \DP_OP_19_294_9081/n441 ), .Y(\DP_OP_19_294_9081/n434 ) );
  AOI21X1 \DP_OP_19_294_9081/U543  ( .A(\DP_OP_19_294_9081/n434 ), .B(
        \DP_OP_19_294_9081/n443 ), .C(\DP_OP_19_294_9081/n435 ), .Y(
        \DP_OP_19_294_9081/n433 ) );
  NAND2X1 \DP_OP_19_294_9081/U541  ( .A(\C2/Z_6 ), .B(\DP_OP_19_294_9081/n659 ), .Y(\DP_OP_19_294_9081/n432 ) );
  NOR2X1 \DP_OP_19_294_9081/U540  ( .A(\C2/Z_6 ), .B(\DP_OP_19_294_9081/n659 ), 
        .Y(\DP_OP_19_294_9081/n431 ) );
  NAND2X1 \DP_OP_19_294_9081/U538  ( .A(\DP_OP_19_294_9081/n432 ), .B(
        \DP_OP_19_294_9081/n514 ), .Y(\DP_OP_19_294_9081/n62 ) );
  OAI21X1 \DP_OP_19_294_9081/U537  ( .A(\DP_OP_19_294_9081/n431 ), .B(
        \DP_OP_19_294_9081/n433 ), .C(\DP_OP_19_294_9081/n432 ), .Y(
        \DP_OP_19_294_9081/n430 ) );
  NAND2X1 \DP_OP_19_294_9081/U535  ( .A(\C2/Z_7 ), .B(\DP_OP_19_294_9081/n660 ), .Y(\DP_OP_19_294_9081/n429 ) );
  NOR2X1 \DP_OP_19_294_9081/U534  ( .A(\C2/Z_7 ), .B(\DP_OP_19_294_9081/n660 ), 
        .Y(\DP_OP_19_294_9081/n428 ) );
  NAND2X1 \DP_OP_19_294_9081/U532  ( .A(\DP_OP_19_294_9081/n429 ), .B(
        \DP_OP_19_294_9081/n513 ), .Y(\DP_OP_19_294_9081/n61 ) );
  OAI21X1 \DP_OP_19_294_9081/U531  ( .A(\DP_OP_19_294_9081/n432 ), .B(
        \DP_OP_19_294_9081/n428 ), .C(\DP_OP_19_294_9081/n429 ), .Y(
        \DP_OP_19_294_9081/n427 ) );
  NOR2X1 \DP_OP_19_294_9081/U530  ( .A(\DP_OP_19_294_9081/n428 ), .B(
        \DP_OP_19_294_9081/n431 ), .Y(\DP_OP_19_294_9081/n426 ) );
  AOI21X1 \DP_OP_19_294_9081/U529  ( .A(\DP_OP_19_294_9081/n435 ), .B(
        \DP_OP_19_294_9081/n426 ), .C(\DP_OP_19_294_9081/n427 ), .Y(
        \DP_OP_19_294_9081/n425 ) );
  NAND2X1 \DP_OP_19_294_9081/U528  ( .A(\DP_OP_19_294_9081/n434 ), .B(
        \DP_OP_19_294_9081/n426 ), .Y(\DP_OP_19_294_9081/n424 ) );
  OAI21X1 \DP_OP_19_294_9081/U527  ( .A(\DP_OP_19_294_9081/n424 ), .B(
        \DP_OP_19_294_9081/n444 ), .C(\DP_OP_19_294_9081/n425 ), .Y(
        \DP_OP_19_294_9081/n423 ) );
  NAND2X1 \DP_OP_19_294_9081/U524  ( .A(\C2/Z_8 ), .B(\DP_OP_19_294_9081/n661 ), .Y(\DP_OP_19_294_9081/n421 ) );
  NOR2X1 \DP_OP_19_294_9081/U523  ( .A(\C2/Z_8 ), .B(\DP_OP_19_294_9081/n661 ), 
        .Y(\DP_OP_19_294_9081/n420 ) );
  NAND2X1 \DP_OP_19_294_9081/U521  ( .A(\DP_OP_19_294_9081/n421 ), .B(
        \DP_OP_19_294_9081/n512 ), .Y(\DP_OP_19_294_9081/n60 ) );
  OAI21X1 \DP_OP_19_294_9081/U520  ( .A(\DP_OP_19_294_9081/n420 ), .B(
        \DP_OP_19_294_9081/n422 ), .C(\DP_OP_19_294_9081/n421 ), .Y(
        \DP_OP_19_294_9081/n419 ) );
  NAND2X1 \DP_OP_19_294_9081/U518  ( .A(\C2/Z_9 ), .B(\DP_OP_19_294_9081/n662 ), .Y(\DP_OP_19_294_9081/n418 ) );
  NOR2X1 \DP_OP_19_294_9081/U517  ( .A(\C2/Z_9 ), .B(\DP_OP_19_294_9081/n662 ), 
        .Y(\DP_OP_19_294_9081/n417 ) );
  NAND2X1 \DP_OP_19_294_9081/U515  ( .A(\DP_OP_19_294_9081/n418 ), .B(
        \DP_OP_19_294_9081/n511 ), .Y(\DP_OP_19_294_9081/n59 ) );
  OAI21X1 \DP_OP_19_294_9081/U514  ( .A(\DP_OP_19_294_9081/n421 ), .B(
        \DP_OP_19_294_9081/n417 ), .C(\DP_OP_19_294_9081/n418 ), .Y(
        \DP_OP_19_294_9081/n416 ) );
  NOR2X1 \DP_OP_19_294_9081/U513  ( .A(\DP_OP_19_294_9081/n417 ), .B(
        \DP_OP_19_294_9081/n420 ), .Y(\DP_OP_19_294_9081/n415 ) );
  OAI21X1 \DP_OP_19_294_9081/U510  ( .A(\DP_OP_19_294_9081/n413 ), .B(
        \DP_OP_19_294_9081/n422 ), .C(\DP_OP_19_294_9081/n414 ), .Y(
        \DP_OP_19_294_9081/n412 ) );
  NAND2X1 \DP_OP_19_294_9081/U508  ( .A(\C2/Z_10 ), .B(
        \DP_OP_19_294_9081/n663 ), .Y(\DP_OP_19_294_9081/n411 ) );
  NOR2X1 \DP_OP_19_294_9081/U507  ( .A(\C2/Z_10 ), .B(\DP_OP_19_294_9081/n663 ), .Y(\DP_OP_19_294_9081/n410 ) );
  NAND2X1 \DP_OP_19_294_9081/U505  ( .A(\DP_OP_19_294_9081/n411 ), .B(
        \DP_OP_19_294_9081/n510 ), .Y(\DP_OP_19_294_9081/n58 ) );
  AOI21X1 \DP_OP_19_294_9081/U502  ( .A(\DP_OP_19_294_9081/n510 ), .B(
        \DP_OP_19_294_9081/n412 ), .C(\DP_OP_19_294_9081/n409 ), .Y(
        \DP_OP_19_294_9081/n407 ) );
  NAND2X1 \DP_OP_19_294_9081/U500  ( .A(\C2/Z_11 ), .B(
        \DP_OP_19_294_9081/n664 ), .Y(\DP_OP_19_294_9081/n406 ) );
  NOR2X1 \DP_OP_19_294_9081/U499  ( .A(\C2/Z_11 ), .B(\DP_OP_19_294_9081/n664 ), .Y(\DP_OP_19_294_9081/n405 ) );
  NAND2X1 \DP_OP_19_294_9081/U497  ( .A(\DP_OP_19_294_9081/n406 ), .B(
        \DP_OP_19_294_9081/n509 ), .Y(\DP_OP_19_294_9081/n57 ) );
  OAI21X1 \DP_OP_19_294_9081/U496  ( .A(\DP_OP_19_294_9081/n411 ), .B(
        \DP_OP_19_294_9081/n405 ), .C(\DP_OP_19_294_9081/n406 ), .Y(
        \DP_OP_19_294_9081/n404 ) );
  NOR2X1 \DP_OP_19_294_9081/U495  ( .A(\DP_OP_19_294_9081/n405 ), .B(
        \DP_OP_19_294_9081/n410 ), .Y(\DP_OP_19_294_9081/n403 ) );
  AOI21X1 \DP_OP_19_294_9081/U494  ( .A(\DP_OP_19_294_9081/n416 ), .B(
        \DP_OP_19_294_9081/n403 ), .C(\DP_OP_19_294_9081/n404 ), .Y(
        \DP_OP_19_294_9081/n402 ) );
  NAND2X1 \DP_OP_19_294_9081/U493  ( .A(\DP_OP_19_294_9081/n403 ), .B(
        \DP_OP_19_294_9081/n415 ), .Y(\DP_OP_19_294_9081/n401 ) );
  OAI21X1 \DP_OP_19_294_9081/U492  ( .A(\DP_OP_19_294_9081/n401 ), .B(
        \DP_OP_19_294_9081/n422 ), .C(\DP_OP_19_294_9081/n402 ), .Y(
        \DP_OP_19_294_9081/n400 ) );
  NAND2X1 \DP_OP_19_294_9081/U489  ( .A(\C2/Z_12 ), .B(
        \DP_OP_19_294_9081/n665 ), .Y(\DP_OP_19_294_9081/n398 ) );
  NOR2X1 \DP_OP_19_294_9081/U488  ( .A(\C2/Z_12 ), .B(\DP_OP_19_294_9081/n665 ), .Y(\DP_OP_19_294_9081/n397 ) );
  NAND2X1 \DP_OP_19_294_9081/U486  ( .A(\DP_OP_19_294_9081/n398 ), .B(
        \DP_OP_19_294_9081/n508 ), .Y(\DP_OP_19_294_9081/n56 ) );
  OAI21X1 \DP_OP_19_294_9081/U485  ( .A(\DP_OP_19_294_9081/n397 ), .B(
        \DP_OP_19_294_9081/n399 ), .C(\DP_OP_19_294_9081/n398 ), .Y(
        \DP_OP_19_294_9081/n396 ) );
  NAND2X1 \DP_OP_19_294_9081/U483  ( .A(\C2/Z_13 ), .B(
        \DP_OP_19_294_9081/n666 ), .Y(\DP_OP_19_294_9081/n395 ) );
  NOR2X1 \DP_OP_19_294_9081/U482  ( .A(\C2/Z_13 ), .B(\DP_OP_19_294_9081/n666 ), .Y(\DP_OP_19_294_9081/n394 ) );
  NAND2X1 \DP_OP_19_294_9081/U480  ( .A(\DP_OP_19_294_9081/n395 ), .B(
        \DP_OP_19_294_9081/n507 ), .Y(\DP_OP_19_294_9081/n55 ) );
  OAI21X1 \DP_OP_19_294_9081/U479  ( .A(\DP_OP_19_294_9081/n398 ), .B(
        \DP_OP_19_294_9081/n394 ), .C(\DP_OP_19_294_9081/n395 ), .Y(
        \DP_OP_19_294_9081/n393 ) );
  NOR2X1 \DP_OP_19_294_9081/U478  ( .A(\DP_OP_19_294_9081/n394 ), .B(
        \DP_OP_19_294_9081/n397 ), .Y(\DP_OP_19_294_9081/n392 ) );
  AOI21X1 \DP_OP_19_294_9081/U477  ( .A(\DP_OP_19_294_9081/n392 ), .B(
        \DP_OP_19_294_9081/n400 ), .C(\DP_OP_19_294_9081/n393 ), .Y(
        \DP_OP_19_294_9081/n391 ) );
  NAND2X1 \DP_OP_19_294_9081/U475  ( .A(\C2/Z_14 ), .B(
        \DP_OP_19_294_9081/n667 ), .Y(\DP_OP_19_294_9081/n390 ) );
  NOR2X1 \DP_OP_19_294_9081/U474  ( .A(\C2/Z_14 ), .B(\DP_OP_19_294_9081/n667 ), .Y(\DP_OP_19_294_9081/n389 ) );
  NAND2X1 \DP_OP_19_294_9081/U472  ( .A(\DP_OP_19_294_9081/n390 ), .B(
        \DP_OP_19_294_9081/n506 ), .Y(\DP_OP_19_294_9081/n54 ) );
  OAI21X1 \DP_OP_19_294_9081/U471  ( .A(\DP_OP_19_294_9081/n389 ), .B(
        \DP_OP_19_294_9081/n391 ), .C(\DP_OP_19_294_9081/n390 ), .Y(
        \DP_OP_19_294_9081/n388 ) );
  NAND2X1 \DP_OP_19_294_9081/U469  ( .A(\C2/Z_15 ), .B(
        \DP_OP_19_294_9081/n668 ), .Y(\DP_OP_19_294_9081/n387 ) );
  NOR2X1 \DP_OP_19_294_9081/U468  ( .A(\C2/Z_15 ), .B(\DP_OP_19_294_9081/n668 ), .Y(\DP_OP_19_294_9081/n386 ) );
  NAND2X1 \DP_OP_19_294_9081/U466  ( .A(\DP_OP_19_294_9081/n387 ), .B(
        \DP_OP_19_294_9081/n505 ), .Y(\DP_OP_19_294_9081/n53 ) );
  OAI21X1 \DP_OP_19_294_9081/U465  ( .A(\DP_OP_19_294_9081/n390 ), .B(
        \DP_OP_19_294_9081/n386 ), .C(\DP_OP_19_294_9081/n387 ), .Y(
        \DP_OP_19_294_9081/n385 ) );
  NOR2X1 \DP_OP_19_294_9081/U464  ( .A(\DP_OP_19_294_9081/n389 ), .B(
        \DP_OP_19_294_9081/n386 ), .Y(\DP_OP_19_294_9081/n384 ) );
  AOI21X1 \DP_OP_19_294_9081/U463  ( .A(\DP_OP_19_294_9081/n393 ), .B(
        \DP_OP_19_294_9081/n384 ), .C(\DP_OP_19_294_9081/n385 ), .Y(
        \DP_OP_19_294_9081/n383 ) );
  NAND2X1 \DP_OP_19_294_9081/U462  ( .A(\DP_OP_19_294_9081/n384 ), .B(
        \DP_OP_19_294_9081/n392 ), .Y(\DP_OP_19_294_9081/n382 ) );
  NAND2X1 \DP_OP_19_294_9081/U456  ( .A(\C2/Z_16 ), .B(
        \DP_OP_19_294_9081/n669 ), .Y(\DP_OP_19_294_9081/n377 ) );
  NOR2X1 \DP_OP_19_294_9081/U455  ( .A(\C2/Z_16 ), .B(\DP_OP_19_294_9081/n669 ), .Y(\DP_OP_19_294_9081/n376 ) );
  NAND2X1 \DP_OP_19_294_9081/U453  ( .A(\DP_OP_19_294_9081/n377 ), .B(
        \DP_OP_19_294_9081/n504 ), .Y(\DP_OP_19_294_9081/n52 ) );
  AOI21X1 \DP_OP_19_294_9081/U450  ( .A(\DP_OP_19_294_9081/n504 ), .B(
        \DP_OP_19_294_9081/n378 ), .C(\DP_OP_19_294_9081/n375 ), .Y(
        \DP_OP_19_294_9081/n373 ) );
  NAND2X1 \DP_OP_19_294_9081/U448  ( .A(\C2/Z_17 ), .B(
        \DP_OP_19_294_9081/n670 ), .Y(\DP_OP_19_294_9081/n372 ) );
  NOR2X1 \DP_OP_19_294_9081/U447  ( .A(\C2/Z_17 ), .B(\DP_OP_19_294_9081/n670 ), .Y(\DP_OP_19_294_9081/n371 ) );
  NAND2X1 \DP_OP_19_294_9081/U445  ( .A(\DP_OP_19_294_9081/n372 ), .B(
        \DP_OP_19_294_9081/n503 ), .Y(\DP_OP_19_294_9081/n51 ) );
  OAI21X1 \DP_OP_19_294_9081/U444  ( .A(\DP_OP_19_294_9081/n377 ), .B(
        \DP_OP_19_294_9081/n371 ), .C(\DP_OP_19_294_9081/n372 ), .Y(
        \DP_OP_19_294_9081/n370 ) );
  NOR2X1 \DP_OP_19_294_9081/U443  ( .A(\DP_OP_19_294_9081/n371 ), .B(
        \DP_OP_19_294_9081/n376 ), .Y(\DP_OP_19_294_9081/n369 ) );
  AOI21X1 \DP_OP_19_294_9081/U442  ( .A(\DP_OP_19_294_9081/n369 ), .B(
        \DP_OP_19_294_9081/n378 ), .C(\DP_OP_19_294_9081/n370 ), .Y(
        \DP_OP_19_294_9081/n368 ) );
  NAND2X1 \DP_OP_19_294_9081/U440  ( .A(\C2/Z_18 ), .B(
        \DP_OP_19_294_9081/n671 ), .Y(\DP_OP_19_294_9081/n367 ) );
  NOR2X1 \DP_OP_19_294_9081/U439  ( .A(\C2/Z_18 ), .B(\DP_OP_19_294_9081/n671 ), .Y(\DP_OP_19_294_9081/n366 ) );
  NAND2X1 \DP_OP_19_294_9081/U437  ( .A(\DP_OP_19_294_9081/n367 ), .B(
        \DP_OP_19_294_9081/n502 ), .Y(\DP_OP_19_294_9081/n50 ) );
  OAI21X1 \DP_OP_19_294_9081/U436  ( .A(\DP_OP_19_294_9081/n366 ), .B(
        \DP_OP_19_294_9081/n368 ), .C(\DP_OP_19_294_9081/n367 ), .Y(
        \DP_OP_19_294_9081/n365 ) );
  NAND2X1 \DP_OP_19_294_9081/U434  ( .A(\C2/Z_19 ), .B(
        \DP_OP_19_294_9081/n672 ), .Y(\DP_OP_19_294_9081/n364 ) );
  NOR2X1 \DP_OP_19_294_9081/U433  ( .A(\C2/Z_19 ), .B(\DP_OP_19_294_9081/n672 ), .Y(\DP_OP_19_294_9081/n363 ) );
  NAND2X1 \DP_OP_19_294_9081/U431  ( .A(\DP_OP_19_294_9081/n364 ), .B(
        \DP_OP_19_294_9081/n501 ), .Y(\DP_OP_19_294_9081/n49 ) );
  OAI21X1 \DP_OP_19_294_9081/U430  ( .A(\DP_OP_19_294_9081/n367 ), .B(
        \DP_OP_19_294_9081/n363 ), .C(\DP_OP_19_294_9081/n364 ), .Y(
        \DP_OP_19_294_9081/n362 ) );
  NOR2X1 \DP_OP_19_294_9081/U429  ( .A(\DP_OP_19_294_9081/n363 ), .B(
        \DP_OP_19_294_9081/n366 ), .Y(\DP_OP_19_294_9081/n361 ) );
  AOI21X1 \DP_OP_19_294_9081/U428  ( .A(\DP_OP_19_294_9081/n370 ), .B(
        \DP_OP_19_294_9081/n361 ), .C(\DP_OP_19_294_9081/n362 ), .Y(
        \DP_OP_19_294_9081/n360 ) );
  NAND2X1 \DP_OP_19_294_9081/U427  ( .A(\DP_OP_19_294_9081/n361 ), .B(
        \DP_OP_19_294_9081/n369 ), .Y(\DP_OP_19_294_9081/n359 ) );
  OAI21X1 \DP_OP_19_294_9081/U426  ( .A(\DP_OP_19_294_9081/n359 ), .B(
        \DP_OP_19_294_9081/n1 ), .C(\DP_OP_19_294_9081/n360 ), .Y(
        \DP_OP_19_294_9081/n358 ) );
  NAND2X1 \DP_OP_19_294_9081/U423  ( .A(\C2/Z_20 ), .B(
        \DP_OP_19_294_9081/n673 ), .Y(\DP_OP_19_294_9081/n356 ) );
  NOR2X1 \DP_OP_19_294_9081/U422  ( .A(\C2/Z_20 ), .B(\DP_OP_19_294_9081/n673 ), .Y(\DP_OP_19_294_9081/n355 ) );
  NAND2X1 \DP_OP_19_294_9081/U420  ( .A(\DP_OP_19_294_9081/n356 ), .B(
        \DP_OP_19_294_9081/n500 ), .Y(\DP_OP_19_294_9081/n48 ) );
  OAI21X1 \DP_OP_19_294_9081/U419  ( .A(\DP_OP_19_294_9081/n355 ), .B(
        \DP_OP_19_294_9081/n357 ), .C(\DP_OP_19_294_9081/n356 ), .Y(
        \DP_OP_19_294_9081/n354 ) );
  NAND2X1 \DP_OP_19_294_9081/U417  ( .A(\C2/Z_21 ), .B(
        \DP_OP_19_294_9081/n674 ), .Y(\DP_OP_19_294_9081/n353 ) );
  NOR2X1 \DP_OP_19_294_9081/U416  ( .A(\C2/Z_21 ), .B(\DP_OP_19_294_9081/n674 ), .Y(\DP_OP_19_294_9081/n352 ) );
  NAND2X1 \DP_OP_19_294_9081/U414  ( .A(\DP_OP_19_294_9081/n353 ), .B(
        \DP_OP_19_294_9081/n499 ), .Y(\DP_OP_19_294_9081/n47 ) );
  OAI21X1 \DP_OP_19_294_9081/U413  ( .A(\DP_OP_19_294_9081/n356 ), .B(
        \DP_OP_19_294_9081/n352 ), .C(\DP_OP_19_294_9081/n353 ), .Y(
        \DP_OP_19_294_9081/n351 ) );
  NOR2X1 \DP_OP_19_294_9081/U412  ( .A(\DP_OP_19_294_9081/n352 ), .B(
        \DP_OP_19_294_9081/n355 ), .Y(\DP_OP_19_294_9081/n350 ) );
  AOI21X1 \DP_OP_19_294_9081/U411  ( .A(\DP_OP_19_294_9081/n350 ), .B(
        \DP_OP_19_294_9081/n358 ), .C(\DP_OP_19_294_9081/n351 ), .Y(
        \DP_OP_19_294_9081/n349 ) );
  NAND2X1 \DP_OP_19_294_9081/U409  ( .A(\C2/Z_22 ), .B(
        \DP_OP_19_294_9081/n675 ), .Y(\DP_OP_19_294_9081/n348 ) );
  NOR2X1 \DP_OP_19_294_9081/U408  ( .A(\C2/Z_22 ), .B(\DP_OP_19_294_9081/n675 ), .Y(\DP_OP_19_294_9081/n347 ) );
  NAND2X1 \DP_OP_19_294_9081/U406  ( .A(\DP_OP_19_294_9081/n348 ), .B(
        \DP_OP_19_294_9081/n498 ), .Y(\DP_OP_19_294_9081/n46 ) );
  OAI21X1 \DP_OP_19_294_9081/U405  ( .A(\DP_OP_19_294_9081/n347 ), .B(
        \DP_OP_19_294_9081/n349 ), .C(\DP_OP_19_294_9081/n348 ), .Y(
        \DP_OP_19_294_9081/n346 ) );
  NAND2X1 \DP_OP_19_294_9081/U403  ( .A(\C2/Z_23 ), .B(
        \DP_OP_19_294_9081/n676 ), .Y(\DP_OP_19_294_9081/n345 ) );
  NOR2X1 \DP_OP_19_294_9081/U402  ( .A(\C2/Z_23 ), .B(\DP_OP_19_294_9081/n676 ), .Y(\DP_OP_19_294_9081/n344 ) );
  NAND2X1 \DP_OP_19_294_9081/U400  ( .A(\DP_OP_19_294_9081/n345 ), .B(
        \DP_OP_19_294_9081/n497 ), .Y(\DP_OP_19_294_9081/n45 ) );
  OAI21X1 \DP_OP_19_294_9081/U399  ( .A(\DP_OP_19_294_9081/n348 ), .B(
        \DP_OP_19_294_9081/n344 ), .C(\DP_OP_19_294_9081/n345 ), .Y(
        \DP_OP_19_294_9081/n343 ) );
  NOR2X1 \DP_OP_19_294_9081/U398  ( .A(\DP_OP_19_294_9081/n344 ), .B(
        \DP_OP_19_294_9081/n347 ), .Y(\DP_OP_19_294_9081/n342 ) );
  AOI21X1 \DP_OP_19_294_9081/U397  ( .A(\DP_OP_19_294_9081/n351 ), .B(
        \DP_OP_19_294_9081/n342 ), .C(\DP_OP_19_294_9081/n343 ), .Y(
        \DP_OP_19_294_9081/n341 ) );
  NAND2X1 \DP_OP_19_294_9081/U396  ( .A(\DP_OP_19_294_9081/n342 ), .B(
        \DP_OP_19_294_9081/n350 ), .Y(\DP_OP_19_294_9081/n340 ) );
  OAI21X1 \DP_OP_19_294_9081/U395  ( .A(\DP_OP_19_294_9081/n340 ), .B(
        \DP_OP_19_294_9081/n360 ), .C(\DP_OP_19_294_9081/n341 ), .Y(
        \DP_OP_19_294_9081/n339 ) );
  NOR2X1 \DP_OP_19_294_9081/U394  ( .A(\DP_OP_19_294_9081/n340 ), .B(
        \DP_OP_19_294_9081/n359 ), .Y(\DP_OP_19_294_9081/n338 ) );
  OAI21X1 \DP_OP_19_294_9081/U391  ( .A(\DP_OP_19_294_9081/n336 ), .B(
        \DP_OP_19_294_9081/n1 ), .C(\DP_OP_19_294_9081/n337 ), .Y(
        \DP_OP_19_294_9081/n335 ) );
  NAND2X1 \DP_OP_19_294_9081/U388  ( .A(\C2/Z_24 ), .B(
        \DP_OP_19_294_9081/n677 ), .Y(\DP_OP_19_294_9081/n333 ) );
  NOR2X1 \DP_OP_19_294_9081/U387  ( .A(\C2/Z_24 ), .B(\DP_OP_19_294_9081/n677 ), .Y(\DP_OP_19_294_9081/n332 ) );
  NAND2X1 \DP_OP_19_294_9081/U385  ( .A(\DP_OP_19_294_9081/n333 ), .B(
        \DP_OP_19_294_9081/n496 ), .Y(\DP_OP_19_294_9081/n44 ) );
  OAI21X1 \DP_OP_19_294_9081/U384  ( .A(\DP_OP_19_294_9081/n332 ), .B(
        \DP_OP_19_294_9081/n334 ), .C(\DP_OP_19_294_9081/n333 ), .Y(
        \DP_OP_19_294_9081/n331 ) );
  NAND2X1 \DP_OP_19_294_9081/U382  ( .A(\C2/Z_25 ), .B(
        \DP_OP_19_294_9081/n678 ), .Y(\DP_OP_19_294_9081/n330 ) );
  NOR2X1 \DP_OP_19_294_9081/U381  ( .A(\C2/Z_25 ), .B(\DP_OP_19_294_9081/n678 ), .Y(\DP_OP_19_294_9081/n329 ) );
  NAND2X1 \DP_OP_19_294_9081/U379  ( .A(\DP_OP_19_294_9081/n330 ), .B(
        \DP_OP_19_294_9081/n495 ), .Y(\DP_OP_19_294_9081/n43 ) );
  OAI21X1 \DP_OP_19_294_9081/U378  ( .A(\DP_OP_19_294_9081/n333 ), .B(
        \DP_OP_19_294_9081/n329 ), .C(\DP_OP_19_294_9081/n330 ), .Y(
        \DP_OP_19_294_9081/n328 ) );
  NOR2X1 \DP_OP_19_294_9081/U377  ( .A(\DP_OP_19_294_9081/n329 ), .B(
        \DP_OP_19_294_9081/n332 ), .Y(\DP_OP_19_294_9081/n327 ) );
  AOI21X1 \DP_OP_19_294_9081/U376  ( .A(\DP_OP_19_294_9081/n327 ), .B(
        \DP_OP_19_294_9081/n335 ), .C(\DP_OP_19_294_9081/n328 ), .Y(
        \DP_OP_19_294_9081/n326 ) );
  NAND2X1 \DP_OP_19_294_9081/U374  ( .A(\C2/Z_26 ), .B(
        \DP_OP_19_294_9081/n679 ), .Y(\DP_OP_19_294_9081/n325 ) );
  NOR2X1 \DP_OP_19_294_9081/U373  ( .A(\C2/Z_26 ), .B(\DP_OP_19_294_9081/n679 ), .Y(\DP_OP_19_294_9081/n324 ) );
  NAND2X1 \DP_OP_19_294_9081/U371  ( .A(\DP_OP_19_294_9081/n325 ), .B(
        \DP_OP_19_294_9081/n494 ), .Y(\DP_OP_19_294_9081/n42 ) );
  OAI21X1 \DP_OP_19_294_9081/U370  ( .A(\DP_OP_19_294_9081/n324 ), .B(
        \DP_OP_19_294_9081/n326 ), .C(\DP_OP_19_294_9081/n325 ), .Y(
        \DP_OP_19_294_9081/n323 ) );
  NAND2X1 \DP_OP_19_294_9081/U368  ( .A(\C2/Z_27 ), .B(
        \DP_OP_19_294_9081/n680 ), .Y(\DP_OP_19_294_9081/n322 ) );
  NOR2X1 \DP_OP_19_294_9081/U367  ( .A(\C2/Z_27 ), .B(\DP_OP_19_294_9081/n680 ), .Y(\DP_OP_19_294_9081/n321 ) );
  NAND2X1 \DP_OP_19_294_9081/U365  ( .A(\DP_OP_19_294_9081/n322 ), .B(
        \DP_OP_19_294_9081/n493 ), .Y(\DP_OP_19_294_9081/n41 ) );
  OAI21X1 \DP_OP_19_294_9081/U364  ( .A(\DP_OP_19_294_9081/n325 ), .B(
        \DP_OP_19_294_9081/n321 ), .C(\DP_OP_19_294_9081/n322 ), .Y(
        \DP_OP_19_294_9081/n320 ) );
  NOR2X1 \DP_OP_19_294_9081/U363  ( .A(\DP_OP_19_294_9081/n321 ), .B(
        \DP_OP_19_294_9081/n324 ), .Y(\DP_OP_19_294_9081/n319 ) );
  AOI21X1 \DP_OP_19_294_9081/U362  ( .A(\DP_OP_19_294_9081/n328 ), .B(
        \DP_OP_19_294_9081/n319 ), .C(\DP_OP_19_294_9081/n320 ), .Y(
        \DP_OP_19_294_9081/n318 ) );
  NAND2X1 \DP_OP_19_294_9081/U361  ( .A(\DP_OP_19_294_9081/n319 ), .B(
        \DP_OP_19_294_9081/n327 ), .Y(\DP_OP_19_294_9081/n317 ) );
  AOI21X1 \DP_OP_19_294_9081/U358  ( .A(\DP_OP_19_294_9081/n315 ), .B(
        \DP_OP_19_294_9081/n339 ), .C(\DP_OP_19_294_9081/n316 ), .Y(
        \DP_OP_19_294_9081/n314 ) );
  NAND2X1 \DP_OP_19_294_9081/U357  ( .A(\DP_OP_19_294_9081/n315 ), .B(
        \DP_OP_19_294_9081/n338 ), .Y(\DP_OP_19_294_9081/n313 ) );
  OAI21X1 \DP_OP_19_294_9081/U356  ( .A(\DP_OP_19_294_9081/n313 ), .B(
        \DP_OP_19_294_9081/n1 ), .C(\DP_OP_19_294_9081/n314 ), .Y(
        \DP_OP_19_294_9081/n312 ) );
  NAND2X1 \DP_OP_19_294_9081/U353  ( .A(\C2/Z_28 ), .B(
        \DP_OP_19_294_9081/n681 ), .Y(\DP_OP_19_294_9081/n310 ) );
  NOR2X1 \DP_OP_19_294_9081/U352  ( .A(\C2/Z_28 ), .B(\DP_OP_19_294_9081/n681 ), .Y(\DP_OP_19_294_9081/n309 ) );
  NAND2X1 \DP_OP_19_294_9081/U350  ( .A(\DP_OP_19_294_9081/n310 ), .B(
        \DP_OP_19_294_9081/n492 ), .Y(\DP_OP_19_294_9081/n40 ) );
  OAI21X1 \DP_OP_19_294_9081/U349  ( .A(\DP_OP_19_294_9081/n309 ), .B(
        \DP_OP_19_294_9081/n311 ), .C(\DP_OP_19_294_9081/n310 ), .Y(
        \DP_OP_19_294_9081/n308 ) );
  NAND2X1 \DP_OP_19_294_9081/U347  ( .A(\C2/Z_29 ), .B(
        \DP_OP_19_294_9081/n682 ), .Y(\DP_OP_19_294_9081/n307 ) );
  NOR2X1 \DP_OP_19_294_9081/U346  ( .A(\C2/Z_29 ), .B(\DP_OP_19_294_9081/n682 ), .Y(\DP_OP_19_294_9081/n306 ) );
  NAND2X1 \DP_OP_19_294_9081/U344  ( .A(\DP_OP_19_294_9081/n307 ), .B(
        \DP_OP_19_294_9081/n491 ), .Y(\DP_OP_19_294_9081/n39 ) );
  OAI21X1 \DP_OP_19_294_9081/U343  ( .A(\DP_OP_19_294_9081/n310 ), .B(
        \DP_OP_19_294_9081/n306 ), .C(\DP_OP_19_294_9081/n307 ), .Y(
        \DP_OP_19_294_9081/n305 ) );
  NOR2X1 \DP_OP_19_294_9081/U342  ( .A(\DP_OP_19_294_9081/n306 ), .B(
        \DP_OP_19_294_9081/n309 ), .Y(\DP_OP_19_294_9081/n304 ) );
  AOI21X1 \DP_OP_19_294_9081/U341  ( .A(\DP_OP_19_294_9081/n304 ), .B(
        \DP_OP_19_294_9081/n312 ), .C(\DP_OP_19_294_9081/n305 ), .Y(
        \DP_OP_19_294_9081/n303 ) );
  NAND2X1 \DP_OP_19_294_9081/U339  ( .A(\C2/Z_30 ), .B(
        \DP_OP_19_294_9081/n683 ), .Y(\DP_OP_19_294_9081/n302 ) );
  NOR2X1 \DP_OP_19_294_9081/U338  ( .A(\C2/Z_30 ), .B(\DP_OP_19_294_9081/n683 ), .Y(\DP_OP_19_294_9081/n301 ) );
  NAND2X1 \DP_OP_19_294_9081/U336  ( .A(\DP_OP_19_294_9081/n302 ), .B(
        \DP_OP_19_294_9081/n490 ), .Y(\DP_OP_19_294_9081/n38 ) );
  OAI21X1 \DP_OP_19_294_9081/U335  ( .A(\DP_OP_19_294_9081/n301 ), .B(
        \DP_OP_19_294_9081/n303 ), .C(\DP_OP_19_294_9081/n302 ), .Y(
        \DP_OP_19_294_9081/n300 ) );
  NAND2X1 \DP_OP_19_294_9081/U333  ( .A(\C2/Z_31 ), .B(
        \DP_OP_19_294_9081/n684 ), .Y(\DP_OP_19_294_9081/n299 ) );
  NOR2X1 \DP_OP_19_294_9081/U332  ( .A(\C2/Z_31 ), .B(\DP_OP_19_294_9081/n684 ), .Y(\DP_OP_19_294_9081/n298 ) );
  NAND2X1 \DP_OP_19_294_9081/U330  ( .A(\DP_OP_19_294_9081/n299 ), .B(
        \DP_OP_19_294_9081/n489 ), .Y(\DP_OP_19_294_9081/n37 ) );
  OAI21X1 \DP_OP_19_294_9081/U329  ( .A(\DP_OP_19_294_9081/n302 ), .B(
        \DP_OP_19_294_9081/n298 ), .C(\DP_OP_19_294_9081/n299 ), .Y(
        \DP_OP_19_294_9081/n297 ) );
  NOR2X1 \DP_OP_19_294_9081/U328  ( .A(\DP_OP_19_294_9081/n298 ), .B(
        \DP_OP_19_294_9081/n301 ), .Y(\DP_OP_19_294_9081/n296 ) );
  AOI21X1 \DP_OP_19_294_9081/U327  ( .A(\DP_OP_19_294_9081/n305 ), .B(
        \DP_OP_19_294_9081/n296 ), .C(\DP_OP_19_294_9081/n297 ), .Y(
        \DP_OP_19_294_9081/n295 ) );
  NAND2X1 \DP_OP_19_294_9081/U326  ( .A(\DP_OP_19_294_9081/n296 ), .B(
        \DP_OP_19_294_9081/n304 ), .Y(\DP_OP_19_294_9081/n294 ) );
  OAI21X1 \DP_OP_19_294_9081/U325  ( .A(\DP_OP_19_294_9081/n294 ), .B(
        \DP_OP_19_294_9081/n318 ), .C(\DP_OP_19_294_9081/n295 ), .Y(
        \DP_OP_19_294_9081/n293 ) );
  NOR2X1 \DP_OP_19_294_9081/U324  ( .A(\DP_OP_19_294_9081/n294 ), .B(
        \DP_OP_19_294_9081/n317 ), .Y(\DP_OP_19_294_9081/n292 ) );
  AOI21X1 \DP_OP_19_294_9081/U323  ( .A(\DP_OP_19_294_9081/n339 ), .B(
        \DP_OP_19_294_9081/n292 ), .C(\DP_OP_19_294_9081/n293 ), .Y(
        \DP_OP_19_294_9081/n291 ) );
  NAND2X1 \DP_OP_19_294_9081/U322  ( .A(\DP_OP_19_294_9081/n292 ), .B(
        \DP_OP_19_294_9081/n338 ), .Y(\DP_OP_19_294_9081/n290 ) );
  OAI21X1 \DP_OP_19_294_9081/U321  ( .A(\DP_OP_19_294_9081/n290 ), .B(
        \DP_OP_19_294_9081/n1 ), .C(\DP_OP_19_294_9081/n291 ), .Y(
        \DP_OP_19_294_9081/n2 ) );
  NAND2X1 \DP_OP_19_294_9081/U318  ( .A(\C2/Z_32 ), .B(
        \DP_OP_19_294_9081/n685 ), .Y(\DP_OP_19_294_9081/n287 ) );
  NOR2X1 \DP_OP_19_294_9081/U317  ( .A(\C2/Z_32 ), .B(\DP_OP_19_294_9081/n685 ), .Y(\DP_OP_19_294_9081/n286 ) );
  NAND2X1 \DP_OP_19_294_9081/U315  ( .A(\DP_OP_19_294_9081/n287 ), .B(
        \DP_OP_19_294_9081/n488 ), .Y(\DP_OP_19_294_9081/n36 ) );
  OAI21X1 \DP_OP_19_294_9081/U314  ( .A(\DP_OP_19_294_9081/n286 ), .B(
        \DP_OP_19_294_9081/n288 ), .C(\DP_OP_19_294_9081/n287 ), .Y(
        \DP_OP_19_294_9081/n285 ) );
  NAND2X1 \DP_OP_19_294_9081/U312  ( .A(\C2/Z_33 ), .B(
        \DP_OP_19_294_9081/n686 ), .Y(\DP_OP_19_294_9081/n284 ) );
  NOR2X1 \DP_OP_19_294_9081/U311  ( .A(\C2/Z_33 ), .B(\DP_OP_19_294_9081/n686 ), .Y(\DP_OP_19_294_9081/n283 ) );
  OAI21X1 \DP_OP_19_294_9081/U308  ( .A(\DP_OP_19_294_9081/n287 ), .B(
        \DP_OP_19_294_9081/n283 ), .C(\DP_OP_19_294_9081/n284 ), .Y(
        \DP_OP_19_294_9081/n282 ) );
  NOR2X1 \DP_OP_19_294_9081/U307  ( .A(\DP_OP_19_294_9081/n286 ), .B(
        \DP_OP_19_294_9081/n283 ), .Y(\DP_OP_19_294_9081/n281 ) );
  AOI21X1 \DP_OP_19_294_9081/U306  ( .A(\DP_OP_19_294_9081/n281 ), .B(n1064), 
        .C(\DP_OP_19_294_9081/n282 ), .Y(\DP_OP_19_294_9081/n280 ) );
  NAND2X1 \DP_OP_19_294_9081/U304  ( .A(\C2/Z_34 ), .B(
        \DP_OP_19_294_9081/n687 ), .Y(\DP_OP_19_294_9081/n279 ) );
  NOR2X1 \DP_OP_19_294_9081/U303  ( .A(\C2/Z_34 ), .B(\DP_OP_19_294_9081/n687 ), .Y(\DP_OP_19_294_9081/n278 ) );
  NAND2X1 \DP_OP_19_294_9081/U301  ( .A(\DP_OP_19_294_9081/n279 ), .B(
        \DP_OP_19_294_9081/n486 ), .Y(\DP_OP_19_294_9081/n34 ) );
  OAI21X1 \DP_OP_19_294_9081/U300  ( .A(\DP_OP_19_294_9081/n280 ), .B(
        \DP_OP_19_294_9081/n278 ), .C(\DP_OP_19_294_9081/n279 ), .Y(
        \DP_OP_19_294_9081/n277 ) );
  NAND2X1 \DP_OP_19_294_9081/U298  ( .A(\C2/Z_35 ), .B(
        \DP_OP_19_294_9081/n688 ), .Y(\DP_OP_19_294_9081/n276 ) );
  NOR2X1 \DP_OP_19_294_9081/U297  ( .A(\C2/Z_35 ), .B(\DP_OP_19_294_9081/n688 ), .Y(\DP_OP_19_294_9081/n275 ) );
  NAND2X1 \DP_OP_19_294_9081/U295  ( .A(\DP_OP_19_294_9081/n276 ), .B(
        \DP_OP_19_294_9081/n485 ), .Y(\DP_OP_19_294_9081/n33 ) );
  OAI21X1 \DP_OP_19_294_9081/U294  ( .A(\DP_OP_19_294_9081/n279 ), .B(
        \DP_OP_19_294_9081/n275 ), .C(\DP_OP_19_294_9081/n276 ), .Y(
        \DP_OP_19_294_9081/n274 ) );
  NOR2X1 \DP_OP_19_294_9081/U293  ( .A(\DP_OP_19_294_9081/n278 ), .B(
        \DP_OP_19_294_9081/n275 ), .Y(\DP_OP_19_294_9081/n273 ) );
  AOI21X1 \DP_OP_19_294_9081/U292  ( .A(\DP_OP_19_294_9081/n282 ), .B(
        \DP_OP_19_294_9081/n273 ), .C(\DP_OP_19_294_9081/n274 ), .Y(
        \DP_OP_19_294_9081/n268 ) );
  NAND2X1 \DP_OP_19_294_9081/U291  ( .A(\DP_OP_19_294_9081/n273 ), .B(
        \DP_OP_19_294_9081/n281 ), .Y(\DP_OP_19_294_9081/n267 ) );
  AOI21X1 \DP_OP_19_294_9081/U284  ( .A(\DP_OP_19_294_9081/n265 ), .B(n1064), 
        .C(\DP_OP_19_294_9081/n266 ), .Y(\DP_OP_19_294_9081/n264 ) );
  NAND2X1 \DP_OP_19_294_9081/U282  ( .A(\C2/Z_36 ), .B(
        \DP_OP_19_294_9081/n689 ), .Y(\DP_OP_19_294_9081/n263 ) );
  NOR2X1 \DP_OP_19_294_9081/U281  ( .A(\C2/Z_36 ), .B(\DP_OP_19_294_9081/n689 ), .Y(\DP_OP_19_294_9081/n262 ) );
  NAND2X1 \DP_OP_19_294_9081/U279  ( .A(\DP_OP_19_294_9081/n263 ), .B(
        \DP_OP_19_294_9081/n484 ), .Y(\DP_OP_19_294_9081/n32 ) );
  OAI21X1 \DP_OP_19_294_9081/U278  ( .A(\DP_OP_19_294_9081/n262 ), .B(
        \DP_OP_19_294_9081/n264 ), .C(\DP_OP_19_294_9081/n263 ), .Y(
        \DP_OP_19_294_9081/n261 ) );
  NAND2X1 \DP_OP_19_294_9081/U276  ( .A(\C2/Z_37 ), .B(
        \DP_OP_19_294_9081/n690 ), .Y(\DP_OP_19_294_9081/n260 ) );
  NOR2X1 \DP_OP_19_294_9081/U275  ( .A(\C2/Z_37 ), .B(\DP_OP_19_294_9081/n690 ), .Y(\DP_OP_19_294_9081/n259 ) );
  OAI21X1 \DP_OP_19_294_9081/U272  ( .A(\DP_OP_19_294_9081/n263 ), .B(
        \DP_OP_19_294_9081/n259 ), .C(\DP_OP_19_294_9081/n260 ), .Y(
        \DP_OP_19_294_9081/n258 ) );
  NOR2X1 \DP_OP_19_294_9081/U271  ( .A(\DP_OP_19_294_9081/n262 ), .B(
        \DP_OP_19_294_9081/n259 ), .Y(\DP_OP_19_294_9081/n257 ) );
  OAI21X1 \DP_OP_19_294_9081/U268  ( .A(\DP_OP_19_294_9081/n255 ), .B(
        \DP_OP_19_294_9081/n268 ), .C(\DP_OP_19_294_9081/n256 ), .Y(
        \DP_OP_19_294_9081/n254 ) );
  NOR2X1 \DP_OP_19_294_9081/U267  ( .A(\DP_OP_19_294_9081/n255 ), .B(
        \DP_OP_19_294_9081/n267 ), .Y(\DP_OP_19_294_9081/n253 ) );
  AOI21X1 \DP_OP_19_294_9081/U266  ( .A(\DP_OP_19_294_9081/n253 ), .B(n1064), 
        .C(\DP_OP_19_294_9081/n254 ), .Y(\DP_OP_19_294_9081/n252 ) );
  NAND2X1 \DP_OP_19_294_9081/U264  ( .A(\C2/Z_38 ), .B(
        \DP_OP_19_294_9081/n691 ), .Y(\DP_OP_19_294_9081/n251 ) );
  NOR2X1 \DP_OP_19_294_9081/U263  ( .A(\C2/Z_38 ), .B(\DP_OP_19_294_9081/n691 ), .Y(\DP_OP_19_294_9081/n250 ) );
  NAND2X1 \DP_OP_19_294_9081/U261  ( .A(\DP_OP_19_294_9081/n251 ), .B(
        \DP_OP_19_294_9081/n482 ), .Y(\DP_OP_19_294_9081/n30 ) );
  OAI21X1 \DP_OP_19_294_9081/U260  ( .A(\DP_OP_19_294_9081/n250 ), .B(
        \DP_OP_19_294_9081/n252 ), .C(\DP_OP_19_294_9081/n251 ), .Y(
        \DP_OP_19_294_9081/n249 ) );
  NAND2X1 \DP_OP_19_294_9081/U258  ( .A(\C2/Z_39 ), .B(
        \DP_OP_19_294_9081/n692 ), .Y(\DP_OP_19_294_9081/n248 ) );
  NOR2X1 \DP_OP_19_294_9081/U257  ( .A(\C2/Z_39 ), .B(\DP_OP_19_294_9081/n692 ), .Y(\DP_OP_19_294_9081/n247 ) );
  OAI21X1 \DP_OP_19_294_9081/U254  ( .A(\DP_OP_19_294_9081/n251 ), .B(
        \DP_OP_19_294_9081/n247 ), .C(\DP_OP_19_294_9081/n248 ), .Y(
        \DP_OP_19_294_9081/n246 ) );
  NOR2X1 \DP_OP_19_294_9081/U253  ( .A(\DP_OP_19_294_9081/n250 ), .B(
        \DP_OP_19_294_9081/n247 ), .Y(\DP_OP_19_294_9081/n245 ) );
  AOI21X1 \DP_OP_19_294_9081/U252  ( .A(\DP_OP_19_294_9081/n258 ), .B(
        \DP_OP_19_294_9081/n245 ), .C(\DP_OP_19_294_9081/n246 ), .Y(
        \DP_OP_19_294_9081/n244 ) );
  NAND2X1 \DP_OP_19_294_9081/U251  ( .A(\DP_OP_19_294_9081/n245 ), .B(
        \DP_OP_19_294_9081/n257 ), .Y(\DP_OP_19_294_9081/n243 ) );
  OAI21X1 \DP_OP_19_294_9081/U250  ( .A(\DP_OP_19_294_9081/n243 ), .B(
        \DP_OP_19_294_9081/n268 ), .C(\DP_OP_19_294_9081/n244 ), .Y(
        \DP_OP_19_294_9081/n238 ) );
  NOR2X1 \DP_OP_19_294_9081/U249  ( .A(\DP_OP_19_294_9081/n267 ), .B(
        \DP_OP_19_294_9081/n243 ), .Y(\DP_OP_19_294_9081/n237 ) );
  AOI21X1 \DP_OP_19_294_9081/U244  ( .A(\DP_OP_19_294_9081/n237 ), .B(n1064), 
        .C(\DP_OP_19_294_9081/n238 ), .Y(\DP_OP_19_294_9081/n236 ) );
  NAND2X1 \DP_OP_19_294_9081/U242  ( .A(\C2/Z_40 ), .B(
        \DP_OP_19_294_9081/n693 ), .Y(\DP_OP_19_294_9081/n235 ) );
  NOR2X1 \DP_OP_19_294_9081/U241  ( .A(\C2/Z_40 ), .B(\DP_OP_19_294_9081/n693 ), .Y(\DP_OP_19_294_9081/n234 ) );
  OAI21X1 \DP_OP_19_294_9081/U238  ( .A(\DP_OP_19_294_9081/n234 ), .B(
        \DP_OP_19_294_9081/n236 ), .C(\DP_OP_19_294_9081/n235 ), .Y(
        \DP_OP_19_294_9081/n233 ) );
  NAND2X1 \DP_OP_19_294_9081/U236  ( .A(\C2/Z_41 ), .B(
        \DP_OP_19_294_9081/n694 ), .Y(\DP_OP_19_294_9081/n232 ) );
  NOR2X1 \DP_OP_19_294_9081/U235  ( .A(\C2/Z_41 ), .B(\DP_OP_19_294_9081/n694 ), .Y(\DP_OP_19_294_9081/n231 ) );
  OAI21X1 \DP_OP_19_294_9081/U232  ( .A(\DP_OP_19_294_9081/n235 ), .B(
        \DP_OP_19_294_9081/n231 ), .C(\DP_OP_19_294_9081/n232 ), .Y(
        \DP_OP_19_294_9081/n230 ) );
  NOR2X1 \DP_OP_19_294_9081/U231  ( .A(\DP_OP_19_294_9081/n234 ), .B(
        \DP_OP_19_294_9081/n231 ), .Y(\DP_OP_19_294_9081/n229 ) );
  OAI21X1 \DP_OP_19_294_9081/U228  ( .A(\DP_OP_19_294_9081/n227 ), .B(
        \DP_OP_19_294_9081/n240 ), .C(\DP_OP_19_294_9081/n228 ), .Y(
        \DP_OP_19_294_9081/n226 ) );
  NOR2X1 \DP_OP_19_294_9081/U227  ( .A(\DP_OP_19_294_9081/n227 ), .B(
        \DP_OP_19_294_9081/n239 ), .Y(\DP_OP_19_294_9081/n225 ) );
  AOI21X1 \DP_OP_19_294_9081/U226  ( .A(\DP_OP_19_294_9081/n225 ), .B(n1064), 
        .C(\DP_OP_19_294_9081/n226 ), .Y(\DP_OP_19_294_9081/n224 ) );
  NAND2X1 \DP_OP_19_294_9081/U224  ( .A(\C2/Z_42 ), .B(
        \DP_OP_19_294_9081/n695 ), .Y(\DP_OP_19_294_9081/n223 ) );
  NOR2X1 \DP_OP_19_294_9081/U223  ( .A(\C2/Z_42 ), .B(\DP_OP_19_294_9081/n695 ), .Y(\DP_OP_19_294_9081/n222 ) );
  NAND2X1 \DP_OP_19_294_9081/U221  ( .A(\DP_OP_19_294_9081/n223 ), .B(
        \DP_OP_19_294_9081/n478 ), .Y(\DP_OP_19_294_9081/n26 ) );
  OAI21X1 \DP_OP_19_294_9081/U220  ( .A(\DP_OP_19_294_9081/n222 ), .B(
        \DP_OP_19_294_9081/n224 ), .C(\DP_OP_19_294_9081/n223 ), .Y(
        \DP_OP_19_294_9081/n221 ) );
  NAND2X1 \DP_OP_19_294_9081/U218  ( .A(\C2/Z_43 ), .B(
        \DP_OP_19_294_9081/n696 ), .Y(\DP_OP_19_294_9081/n220 ) );
  NOR2X1 \DP_OP_19_294_9081/U217  ( .A(\C2/Z_43 ), .B(\DP_OP_19_294_9081/n696 ), .Y(\DP_OP_19_294_9081/n219 ) );
  OAI21X1 \DP_OP_19_294_9081/U214  ( .A(\DP_OP_19_294_9081/n223 ), .B(
        \DP_OP_19_294_9081/n219 ), .C(\DP_OP_19_294_9081/n220 ), .Y(
        \DP_OP_19_294_9081/n218 ) );
  NOR2X1 \DP_OP_19_294_9081/U213  ( .A(\DP_OP_19_294_9081/n222 ), .B(
        \DP_OP_19_294_9081/n219 ), .Y(\DP_OP_19_294_9081/n217 ) );
  AOI21X1 \DP_OP_19_294_9081/U212  ( .A(\DP_OP_19_294_9081/n230 ), .B(
        \DP_OP_19_294_9081/n217 ), .C(\DP_OP_19_294_9081/n218 ), .Y(
        \DP_OP_19_294_9081/n216 ) );
  NAND2X1 \DP_OP_19_294_9081/U211  ( .A(\DP_OP_19_294_9081/n217 ), .B(
        \DP_OP_19_294_9081/n229 ), .Y(\DP_OP_19_294_9081/n215 ) );
  AOI21X1 \DP_OP_19_294_9081/U208  ( .A(\DP_OP_19_294_9081/n213 ), .B(
        \DP_OP_19_294_9081/n238 ), .C(\DP_OP_19_294_9081/n214 ), .Y(
        \DP_OP_19_294_9081/n212 ) );
  NAND2X1 \DP_OP_19_294_9081/U207  ( .A(\DP_OP_19_294_9081/n213 ), .B(
        \DP_OP_19_294_9081/n237 ), .Y(\DP_OP_19_294_9081/n211 ) );
  AOI21X1 \DP_OP_19_294_9081/U204  ( .A(\DP_OP_19_294_9081/n209 ), .B(n1064), 
        .C(\DP_OP_19_294_9081/n210 ), .Y(\DP_OP_19_294_9081/n208 ) );
  NAND2X1 \DP_OP_19_294_9081/U202  ( .A(\C2/Z_44 ), .B(
        \DP_OP_19_294_9081/n697 ), .Y(\DP_OP_19_294_9081/n207 ) );
  NOR2X1 \DP_OP_19_294_9081/U201  ( .A(\C2/Z_44 ), .B(\DP_OP_19_294_9081/n697 ), .Y(\DP_OP_19_294_9081/n206 ) );
  NAND2X1 \DP_OP_19_294_9081/U199  ( .A(\DP_OP_19_294_9081/n207 ), .B(
        \DP_OP_19_294_9081/n476 ), .Y(\DP_OP_19_294_9081/n24 ) );
  OAI21X1 \DP_OP_19_294_9081/U198  ( .A(\DP_OP_19_294_9081/n206 ), .B(
        \DP_OP_19_294_9081/n208 ), .C(\DP_OP_19_294_9081/n207 ), .Y(
        \DP_OP_19_294_9081/n205 ) );
  NAND2X1 \DP_OP_19_294_9081/U196  ( .A(\C2/Z_45 ), .B(
        \DP_OP_19_294_9081/n698 ), .Y(\DP_OP_19_294_9081/n204 ) );
  NOR2X1 \DP_OP_19_294_9081/U195  ( .A(\C2/Z_45 ), .B(\DP_OP_19_294_9081/n698 ), .Y(\DP_OP_19_294_9081/n203 ) );
  OAI21X1 \DP_OP_19_294_9081/U192  ( .A(\DP_OP_19_294_9081/n207 ), .B(
        \DP_OP_19_294_9081/n203 ), .C(\DP_OP_19_294_9081/n204 ), .Y(
        \DP_OP_19_294_9081/n202 ) );
  NOR2X1 \DP_OP_19_294_9081/U191  ( .A(\DP_OP_19_294_9081/n206 ), .B(
        \DP_OP_19_294_9081/n203 ), .Y(\DP_OP_19_294_9081/n201 ) );
  OAI21X1 \DP_OP_19_294_9081/U188  ( .A(\DP_OP_19_294_9081/n199 ), .B(
        \DP_OP_19_294_9081/n212 ), .C(\DP_OP_19_294_9081/n200 ), .Y(
        \DP_OP_19_294_9081/n198 ) );
  NOR2X1 \DP_OP_19_294_9081/U187  ( .A(\DP_OP_19_294_9081/n199 ), .B(
        \DP_OP_19_294_9081/n211 ), .Y(\DP_OP_19_294_9081/n197 ) );
  AOI21X1 \DP_OP_19_294_9081/U186  ( .A(n1064), .B(\DP_OP_19_294_9081/n197 ), 
        .C(\DP_OP_19_294_9081/n198 ), .Y(\DP_OP_19_294_9081/n196 ) );
  NAND2X1 \DP_OP_19_294_9081/U184  ( .A(\C2/Z_46 ), .B(
        \DP_OP_19_294_9081/n699 ), .Y(\DP_OP_19_294_9081/n195 ) );
  NOR2X1 \DP_OP_19_294_9081/U183  ( .A(\C2/Z_46 ), .B(\DP_OP_19_294_9081/n699 ), .Y(\DP_OP_19_294_9081/n194 ) );
  NAND2X1 \DP_OP_19_294_9081/U181  ( .A(\DP_OP_19_294_9081/n195 ), .B(
        \DP_OP_19_294_9081/n474 ), .Y(\DP_OP_19_294_9081/n22 ) );
  OAI21X1 \DP_OP_19_294_9081/U180  ( .A(\DP_OP_19_294_9081/n194 ), .B(
        \DP_OP_19_294_9081/n196 ), .C(\DP_OP_19_294_9081/n195 ), .Y(
        \DP_OP_19_294_9081/n193 ) );
  NAND2X1 \DP_OP_19_294_9081/U178  ( .A(\C2/Z_47 ), .B(
        \DP_OP_19_294_9081/n700 ), .Y(\DP_OP_19_294_9081/n192 ) );
  NOR2X1 \DP_OP_19_294_9081/U177  ( .A(\C2/Z_47 ), .B(\DP_OP_19_294_9081/n700 ), .Y(\DP_OP_19_294_9081/n191 ) );
  NAND2X1 \DP_OP_19_294_9081/U175  ( .A(\DP_OP_19_294_9081/n192 ), .B(
        \DP_OP_19_294_9081/n473 ), .Y(\DP_OP_19_294_9081/n21 ) );
  OAI21X1 \DP_OP_19_294_9081/U174  ( .A(\DP_OP_19_294_9081/n195 ), .B(
        \DP_OP_19_294_9081/n191 ), .C(\DP_OP_19_294_9081/n192 ), .Y(
        \DP_OP_19_294_9081/n190 ) );
  NOR2X1 \DP_OP_19_294_9081/U173  ( .A(\DP_OP_19_294_9081/n194 ), .B(
        \DP_OP_19_294_9081/n191 ), .Y(\DP_OP_19_294_9081/n189 ) );
  AOI21X1 \DP_OP_19_294_9081/U172  ( .A(\DP_OP_19_294_9081/n202 ), .B(
        \DP_OP_19_294_9081/n189 ), .C(\DP_OP_19_294_9081/n190 ), .Y(
        \DP_OP_19_294_9081/n188 ) );
  NAND2X1 \DP_OP_19_294_9081/U171  ( .A(\DP_OP_19_294_9081/n189 ), .B(
        \DP_OP_19_294_9081/n201 ), .Y(\DP_OP_19_294_9081/n187 ) );
  OAI21X1 \DP_OP_19_294_9081/U170  ( .A(\DP_OP_19_294_9081/n187 ), .B(
        \DP_OP_19_294_9081/n216 ), .C(\DP_OP_19_294_9081/n188 ), .Y(
        \DP_OP_19_294_9081/n186 ) );
  NOR2X1 \DP_OP_19_294_9081/U169  ( .A(\DP_OP_19_294_9081/n215 ), .B(
        \DP_OP_19_294_9081/n187 ), .Y(\DP_OP_19_294_9081/n185 ) );
  AOI21X1 \DP_OP_19_294_9081/U168  ( .A(\DP_OP_19_294_9081/n238 ), .B(
        \DP_OP_19_294_9081/n185 ), .C(\DP_OP_19_294_9081/n186 ), .Y(
        \DP_OP_19_294_9081/n3 ) );
  NAND2X1 \DP_OP_19_294_9081/U167  ( .A(\DP_OP_19_294_9081/n237 ), .B(
        \DP_OP_19_294_9081/n185 ), .Y(\DP_OP_19_294_9081/n4 ) );
  AOI21X1 \DP_OP_19_294_9081/U164  ( .A(\DP_OP_19_294_9081/n181 ), .B(n1064), 
        .C(\DP_OP_19_294_9081/n182 ), .Y(\DP_OP_19_294_9081/n180 ) );
  NAND2X1 \DP_OP_19_294_9081/U162  ( .A(\C2/Z_48 ), .B(
        \DP_OP_19_294_9081/n701 ), .Y(\DP_OP_19_294_9081/n179 ) );
  NOR2X1 \DP_OP_19_294_9081/U161  ( .A(\C2/Z_48 ), .B(\DP_OP_19_294_9081/n701 ), .Y(\DP_OP_19_294_9081/n178 ) );
  NAND2X1 \DP_OP_19_294_9081/U159  ( .A(\DP_OP_19_294_9081/n179 ), .B(
        \DP_OP_19_294_9081/n472 ), .Y(\DP_OP_19_294_9081/n20 ) );
  OAI21X1 \DP_OP_19_294_9081/U158  ( .A(\DP_OP_19_294_9081/n178 ), .B(
        \DP_OP_19_294_9081/n180 ), .C(\DP_OP_19_294_9081/n179 ), .Y(
        \DP_OP_19_294_9081/n177 ) );
  NAND2X1 \DP_OP_19_294_9081/U156  ( .A(\C2/Z_49 ), .B(
        \DP_OP_19_294_9081/n702 ), .Y(\DP_OP_19_294_9081/n176 ) );
  NOR2X1 \DP_OP_19_294_9081/U155  ( .A(\C2/Z_49 ), .B(\DP_OP_19_294_9081/n702 ), .Y(\DP_OP_19_294_9081/n175 ) );
  OAI21X1 \DP_OP_19_294_9081/U152  ( .A(\DP_OP_19_294_9081/n179 ), .B(
        \DP_OP_19_294_9081/n175 ), .C(\DP_OP_19_294_9081/n176 ), .Y(
        \DP_OP_19_294_9081/n174 ) );
  NOR2X1 \DP_OP_19_294_9081/U151  ( .A(\DP_OP_19_294_9081/n178 ), .B(
        \DP_OP_19_294_9081/n175 ), .Y(\DP_OP_19_294_9081/n173 ) );
  OAI21X1 \DP_OP_19_294_9081/U148  ( .A(\DP_OP_19_294_9081/n171 ), .B(
        \DP_OP_19_294_9081/n3 ), .C(\DP_OP_19_294_9081/n172 ), .Y(
        \DP_OP_19_294_9081/n170 ) );
  NOR2X1 \DP_OP_19_294_9081/U147  ( .A(\DP_OP_19_294_9081/n171 ), .B(
        \DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n169 ) );
  AOI21X1 \DP_OP_19_294_9081/U146  ( .A(n1064), .B(\DP_OP_19_294_9081/n169 ), 
        .C(\DP_OP_19_294_9081/n170 ), .Y(\DP_OP_19_294_9081/n168 ) );
  NAND2X1 \DP_OP_19_294_9081/U144  ( .A(\C2/Z_50 ), .B(
        \DP_OP_19_294_9081/n703 ), .Y(\DP_OP_19_294_9081/n167 ) );
  NOR2X1 \DP_OP_19_294_9081/U143  ( .A(\C2/Z_50 ), .B(\DP_OP_19_294_9081/n703 ), .Y(\DP_OP_19_294_9081/n166 ) );
  NAND2X1 \DP_OP_19_294_9081/U141  ( .A(\DP_OP_19_294_9081/n167 ), .B(
        \DP_OP_19_294_9081/n470 ), .Y(\DP_OP_19_294_9081/n18 ) );
  OAI21X1 \DP_OP_19_294_9081/U140  ( .A(\DP_OP_19_294_9081/n166 ), .B(
        \DP_OP_19_294_9081/n168 ), .C(\DP_OP_19_294_9081/n167 ), .Y(
        \DP_OP_19_294_9081/n165 ) );
  NAND2X1 \DP_OP_19_294_9081/U138  ( .A(\C2/Z_51 ), .B(
        \DP_OP_19_294_9081/n704 ), .Y(\DP_OP_19_294_9081/n164 ) );
  NOR2X1 \DP_OP_19_294_9081/U137  ( .A(\C2/Z_51 ), .B(\DP_OP_19_294_9081/n704 ), .Y(\DP_OP_19_294_9081/n163 ) );
  NAND2X1 \DP_OP_19_294_9081/U135  ( .A(\DP_OP_19_294_9081/n164 ), .B(
        \DP_OP_19_294_9081/n469 ), .Y(\DP_OP_19_294_9081/n17 ) );
  OAI21X1 \DP_OP_19_294_9081/U134  ( .A(\DP_OP_19_294_9081/n167 ), .B(
        \DP_OP_19_294_9081/n163 ), .C(\DP_OP_19_294_9081/n164 ), .Y(
        \DP_OP_19_294_9081/n162 ) );
  NOR2X1 \DP_OP_19_294_9081/U133  ( .A(\DP_OP_19_294_9081/n166 ), .B(
        \DP_OP_19_294_9081/n163 ), .Y(\DP_OP_19_294_9081/n161 ) );
  AOI21X1 \DP_OP_19_294_9081/U132  ( .A(\DP_OP_19_294_9081/n174 ), .B(
        \DP_OP_19_294_9081/n161 ), .C(\DP_OP_19_294_9081/n162 ), .Y(
        \DP_OP_19_294_9081/n156 ) );
  NAND2X1 \DP_OP_19_294_9081/U131  ( .A(\DP_OP_19_294_9081/n161 ), .B(
        \DP_OP_19_294_9081/n173 ), .Y(\DP_OP_19_294_9081/n155 ) );
  OAI21X1 \DP_OP_19_294_9081/U126  ( .A(\DP_OP_19_294_9081/n155 ), .B(
        \DP_OP_19_294_9081/n3 ), .C(\DP_OP_19_294_9081/n156 ), .Y(
        \DP_OP_19_294_9081/n154 ) );
  NOR2X1 \DP_OP_19_294_9081/U125  ( .A(\DP_OP_19_294_9081/n155 ), .B(
        \DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n153 ) );
  AOI21X1 \DP_OP_19_294_9081/U124  ( .A(n1064), .B(\DP_OP_19_294_9081/n153 ), 
        .C(\DP_OP_19_294_9081/n154 ), .Y(\DP_OP_19_294_9081/n152 ) );
  NAND2X1 \DP_OP_19_294_9081/U122  ( .A(\C2/Z_52 ), .B(
        \DP_OP_19_294_9081/n705 ), .Y(\DP_OP_19_294_9081/n151 ) );
  NOR2X1 \DP_OP_19_294_9081/U121  ( .A(\C2/Z_52 ), .B(\DP_OP_19_294_9081/n705 ), .Y(\DP_OP_19_294_9081/n150 ) );
  NAND2X1 \DP_OP_19_294_9081/U119  ( .A(\DP_OP_19_294_9081/n151 ), .B(
        \DP_OP_19_294_9081/n468 ), .Y(\DP_OP_19_294_9081/n16 ) );
  OAI21X1 \DP_OP_19_294_9081/U118  ( .A(\DP_OP_19_294_9081/n150 ), .B(
        \DP_OP_19_294_9081/n152 ), .C(\DP_OP_19_294_9081/n151 ), .Y(
        \DP_OP_19_294_9081/n149 ) );
  NAND2X1 \DP_OP_19_294_9081/U116  ( .A(\C2/Z_53 ), .B(
        \DP_OP_19_294_9081/n706 ), .Y(\DP_OP_19_294_9081/n148 ) );
  NOR2X1 \DP_OP_19_294_9081/U115  ( .A(\C2/Z_53 ), .B(\DP_OP_19_294_9081/n706 ), .Y(\DP_OP_19_294_9081/n147 ) );
  NAND2X1 \DP_OP_19_294_9081/U113  ( .A(\DP_OP_19_294_9081/n148 ), .B(
        \DP_OP_19_294_9081/n467 ), .Y(\DP_OP_19_294_9081/n15 ) );
  OAI21X1 \DP_OP_19_294_9081/U112  ( .A(\DP_OP_19_294_9081/n151 ), .B(
        \DP_OP_19_294_9081/n147 ), .C(\DP_OP_19_294_9081/n148 ), .Y(
        \DP_OP_19_294_9081/n146 ) );
  NOR2X1 \DP_OP_19_294_9081/U111  ( .A(\DP_OP_19_294_9081/n150 ), .B(
        \DP_OP_19_294_9081/n147 ), .Y(\DP_OP_19_294_9081/n143 ) );
  AOI21X1 \DP_OP_19_294_9081/U108  ( .A(\DP_OP_19_294_9081/n143 ), .B(
        \DP_OP_19_294_9081/n158 ), .C(\DP_OP_19_294_9081/n146 ), .Y(
        \DP_OP_19_294_9081/n142 ) );
  NAND2X1 \DP_OP_19_294_9081/U107  ( .A(\DP_OP_19_294_9081/n143 ), .B(
        \DP_OP_19_294_9081/n157 ), .Y(\DP_OP_19_294_9081/n141 ) );
  OAI21X1 \DP_OP_19_294_9081/U106  ( .A(\DP_OP_19_294_9081/n141 ), .B(
        \DP_OP_19_294_9081/n3 ), .C(\DP_OP_19_294_9081/n142 ), .Y(
        \DP_OP_19_294_9081/n140 ) );
  NOR2X1 \DP_OP_19_294_9081/U105  ( .A(\DP_OP_19_294_9081/n141 ), .B(
        \DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n139 ) );
  AOI21X1 \DP_OP_19_294_9081/U104  ( .A(n1064), .B(\DP_OP_19_294_9081/n139 ), 
        .C(\DP_OP_19_294_9081/n140 ), .Y(\DP_OP_19_294_9081/n138 ) );
  NAND2X1 \DP_OP_19_294_9081/U102  ( .A(\C2/Z_54 ), .B(
        \DP_OP_19_294_9081/n707 ), .Y(\DP_OP_19_294_9081/n137 ) );
  NOR2X1 \DP_OP_19_294_9081/U101  ( .A(\C2/Z_54 ), .B(\DP_OP_19_294_9081/n707 ), .Y(\DP_OP_19_294_9081/n136 ) );
  NAND2X1 \DP_OP_19_294_9081/U99  ( .A(\DP_OP_19_294_9081/n137 ), .B(
        \DP_OP_19_294_9081/n466 ), .Y(\DP_OP_19_294_9081/n14 ) );
  OAI21X1 \DP_OP_19_294_9081/U98  ( .A(\DP_OP_19_294_9081/n136 ), .B(
        \DP_OP_19_294_9081/n138 ), .C(\DP_OP_19_294_9081/n137 ), .Y(
        \DP_OP_19_294_9081/n135 ) );
  NAND2X1 \DP_OP_19_294_9081/U96  ( .A(\C2/Z_55 ), .B(\DP_OP_19_294_9081/n708 ), .Y(\DP_OP_19_294_9081/n134 ) );
  NOR2X1 \DP_OP_19_294_9081/U95  ( .A(\C2/Z_55 ), .B(\DP_OP_19_294_9081/n708 ), 
        .Y(\DP_OP_19_294_9081/n133 ) );
  NAND2X1 \DP_OP_19_294_9081/U93  ( .A(\DP_OP_19_294_9081/n134 ), .B(
        \DP_OP_19_294_9081/n465 ), .Y(\DP_OP_19_294_9081/n13 ) );
  OAI21X1 \DP_OP_19_294_9081/U92  ( .A(\DP_OP_19_294_9081/n137 ), .B(
        \DP_OP_19_294_9081/n133 ), .C(\DP_OP_19_294_9081/n134 ), .Y(
        \DP_OP_19_294_9081/n132 ) );
  NOR2X1 \DP_OP_19_294_9081/U91  ( .A(\DP_OP_19_294_9081/n136 ), .B(
        \DP_OP_19_294_9081/n133 ), .Y(\DP_OP_19_294_9081/n131 ) );
  AOI21X1 \DP_OP_19_294_9081/U90  ( .A(\DP_OP_19_294_9081/n146 ), .B(
        \DP_OP_19_294_9081/n131 ), .C(\DP_OP_19_294_9081/n132 ), .Y(
        \DP_OP_19_294_9081/n130 ) );
  NAND2X1 \DP_OP_19_294_9081/U89  ( .A(\DP_OP_19_294_9081/n131 ), .B(
        \DP_OP_19_294_9081/n143 ), .Y(\DP_OP_19_294_9081/n129 ) );
  OAI21X1 \DP_OP_19_294_9081/U88  ( .A(\DP_OP_19_294_9081/n129 ), .B(
        \DP_OP_19_294_9081/n156 ), .C(\DP_OP_19_294_9081/n130 ), .Y(
        \DP_OP_19_294_9081/n128 ) );
  NOR2X1 \DP_OP_19_294_9081/U87  ( .A(\DP_OP_19_294_9081/n155 ), .B(
        \DP_OP_19_294_9081/n129 ), .Y(\DP_OP_19_294_9081/n127 ) );
  OAI21X1 \DP_OP_19_294_9081/U84  ( .A(\DP_OP_19_294_9081/n125 ), .B(
        \DP_OP_19_294_9081/n3 ), .C(\DP_OP_19_294_9081/n126 ), .Y(
        \DP_OP_19_294_9081/n124 ) );
  NOR2X1 \DP_OP_19_294_9081/U83  ( .A(\DP_OP_19_294_9081/n125 ), .B(
        \DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n123 ) );
  AOI21X1 \DP_OP_19_294_9081/U82  ( .A(n1064), .B(\DP_OP_19_294_9081/n123 ), 
        .C(\DP_OP_19_294_9081/n124 ), .Y(\DP_OP_19_294_9081/n122 ) );
  NAND2X1 \DP_OP_19_294_9081/U80  ( .A(\C2/Z_56 ), .B(\DP_OP_19_294_9081/n709 ), .Y(\DP_OP_19_294_9081/n121 ) );
  NOR2X1 \DP_OP_19_294_9081/U79  ( .A(\C2/Z_56 ), .B(\DP_OP_19_294_9081/n709 ), 
        .Y(\DP_OP_19_294_9081/n120 ) );
  NAND2X1 \DP_OP_19_294_9081/U77  ( .A(\DP_OP_19_294_9081/n121 ), .B(
        \DP_OP_19_294_9081/n464 ), .Y(\DP_OP_19_294_9081/n12 ) );
  OAI21X1 \DP_OP_19_294_9081/U76  ( .A(\DP_OP_19_294_9081/n120 ), .B(
        \DP_OP_19_294_9081/n122 ), .C(\DP_OP_19_294_9081/n121 ), .Y(
        \DP_OP_19_294_9081/n119 ) );
  NAND2X1 \DP_OP_19_294_9081/U74  ( .A(\C2/Z_57 ), .B(\DP_OP_19_294_9081/n710 ), .Y(\DP_OP_19_294_9081/n118 ) );
  NOR2X1 \DP_OP_19_294_9081/U73  ( .A(\C2/Z_57 ), .B(\DP_OP_19_294_9081/n710 ), 
        .Y(\DP_OP_19_294_9081/n117 ) );
  NAND2X1 \DP_OP_19_294_9081/U71  ( .A(\DP_OP_19_294_9081/n118 ), .B(
        \DP_OP_19_294_9081/n463 ), .Y(\DP_OP_19_294_9081/n11 ) );
  OAI21X1 \DP_OP_19_294_9081/U70  ( .A(\DP_OP_19_294_9081/n121 ), .B(
        \DP_OP_19_294_9081/n117 ), .C(\DP_OP_19_294_9081/n118 ), .Y(
        \DP_OP_19_294_9081/n116 ) );
  NOR2X1 \DP_OP_19_294_9081/U69  ( .A(\DP_OP_19_294_9081/n120 ), .B(
        \DP_OP_19_294_9081/n117 ), .Y(\DP_OP_19_294_9081/n113 ) );
  AOI21X1 \DP_OP_19_294_9081/U66  ( .A(\DP_OP_19_294_9081/n113 ), .B(
        \DP_OP_19_294_9081/n128 ), .C(\DP_OP_19_294_9081/n116 ), .Y(
        \DP_OP_19_294_9081/n112 ) );
  NAND2X1 \DP_OP_19_294_9081/U65  ( .A(\DP_OP_19_294_9081/n113 ), .B(
        \DP_OP_19_294_9081/n127 ), .Y(\DP_OP_19_294_9081/n111 ) );
  OAI21X1 \DP_OP_19_294_9081/U64  ( .A(\DP_OP_19_294_9081/n3 ), .B(
        \DP_OP_19_294_9081/n111 ), .C(\DP_OP_19_294_9081/n112 ), .Y(
        \DP_OP_19_294_9081/n110 ) );
  NOR2X1 \DP_OP_19_294_9081/U63  ( .A(\DP_OP_19_294_9081/n111 ), .B(
        \DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n109 ) );
  AOI21X1 \DP_OP_19_294_9081/U62  ( .A(n1064), .B(\DP_OP_19_294_9081/n109 ), 
        .C(\DP_OP_19_294_9081/n110 ), .Y(\DP_OP_19_294_9081/n108 ) );
  NAND2X1 \DP_OP_19_294_9081/U60  ( .A(\C2/Z_58 ), .B(\DP_OP_19_294_9081/n711 ), .Y(\DP_OP_19_294_9081/n107 ) );
  NOR2X1 \DP_OP_19_294_9081/U59  ( .A(\C2/Z_58 ), .B(\DP_OP_19_294_9081/n711 ), 
        .Y(\DP_OP_19_294_9081/n106 ) );
  NAND2X1 \DP_OP_19_294_9081/U57  ( .A(\DP_OP_19_294_9081/n107 ), .B(
        \DP_OP_19_294_9081/n462 ), .Y(\DP_OP_19_294_9081/n10 ) );
  OAI21X1 \DP_OP_19_294_9081/U56  ( .A(\DP_OP_19_294_9081/n106 ), .B(
        \DP_OP_19_294_9081/n108 ), .C(\DP_OP_19_294_9081/n107 ), .Y(
        \DP_OP_19_294_9081/n105 ) );
  NAND2X1 \DP_OP_19_294_9081/U54  ( .A(\C2/Z_59 ), .B(\DP_OP_19_294_9081/n712 ), .Y(\DP_OP_19_294_9081/n104 ) );
  NOR2X1 \DP_OP_19_294_9081/U53  ( .A(\C2/Z_59 ), .B(\DP_OP_19_294_9081/n712 ), 
        .Y(\DP_OP_19_294_9081/n103 ) );
  NAND2X1 \DP_OP_19_294_9081/U51  ( .A(\DP_OP_19_294_9081/n104 ), .B(
        \DP_OP_19_294_9081/n461 ), .Y(\DP_OP_19_294_9081/n9 ) );
  OAI21X1 \DP_OP_19_294_9081/U50  ( .A(\DP_OP_19_294_9081/n107 ), .B(
        \DP_OP_19_294_9081/n103 ), .C(\DP_OP_19_294_9081/n104 ), .Y(
        \DP_OP_19_294_9081/n102 ) );
  NOR2X1 \DP_OP_19_294_9081/U49  ( .A(\DP_OP_19_294_9081/n106 ), .B(
        \DP_OP_19_294_9081/n103 ), .Y(\DP_OP_19_294_9081/n101 ) );
  AOI21X1 \DP_OP_19_294_9081/U48  ( .A(\DP_OP_19_294_9081/n116 ), .B(
        \DP_OP_19_294_9081/n101 ), .C(\DP_OP_19_294_9081/n102 ), .Y(
        \DP_OP_19_294_9081/n100 ) );
  NAND2X1 \DP_OP_19_294_9081/U47  ( .A(\DP_OP_19_294_9081/n101 ), .B(
        \DP_OP_19_294_9081/n113 ), .Y(\DP_OP_19_294_9081/n99 ) );
  AOI21X1 \DP_OP_19_294_9081/U44  ( .A(\DP_OP_19_294_9081/n97 ), .B(
        \DP_OP_19_294_9081/n128 ), .C(\DP_OP_19_294_9081/n98 ), .Y(
        \DP_OP_19_294_9081/n96 ) );
  NAND2X1 \DP_OP_19_294_9081/U43  ( .A(\DP_OP_19_294_9081/n97 ), .B(
        \DP_OP_19_294_9081/n127 ), .Y(\DP_OP_19_294_9081/n95 ) );
  OAI21X1 \DP_OP_19_294_9081/U42  ( .A(\DP_OP_19_294_9081/n95 ), .B(
        \DP_OP_19_294_9081/n3 ), .C(\DP_OP_19_294_9081/n96 ), .Y(
        \DP_OP_19_294_9081/n94 ) );
  NOR2X1 \DP_OP_19_294_9081/U41  ( .A(\DP_OP_19_294_9081/n95 ), .B(
        \DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n93 ) );
  AOI21X1 \DP_OP_19_294_9081/U40  ( .A(n1064), .B(\DP_OP_19_294_9081/n93 ), 
        .C(\DP_OP_19_294_9081/n94 ), .Y(\DP_OP_19_294_9081/n92 ) );
  NAND2X1 \DP_OP_19_294_9081/U38  ( .A(\C2/Z_60 ), .B(\DP_OP_19_294_9081/n713 ), .Y(\DP_OP_19_294_9081/n87 ) );
  NOR2X1 \DP_OP_19_294_9081/U37  ( .A(\C2/Z_60 ), .B(\DP_OP_19_294_9081/n713 ), 
        .Y(\DP_OP_19_294_9081/n86 ) );
  NAND2X1 \DP_OP_19_294_9081/U35  ( .A(\DP_OP_19_294_9081/n87 ), .B(
        \DP_OP_19_294_9081/n88 ), .Y(\DP_OP_19_294_9081/n8 ) );
  OAI21X1 \DP_OP_19_294_9081/U30  ( .A(\DP_OP_19_294_9081/n86 ), .B(
        \DP_OP_19_294_9081/n92 ), .C(\DP_OP_19_294_9081/n87 ), .Y(
        \DP_OP_19_294_9081/n85 ) );
  NAND2X1 \DP_OP_19_294_9081/U28  ( .A(\C2/Z_61 ), .B(\DP_OP_19_294_9081/n714 ), .Y(\DP_OP_19_294_9081/n84 ) );
  NAND2X1 \DP_OP_19_294_9081/U25  ( .A(\DP_OP_19_294_9081/n84 ), .B(n1089), 
        .Y(\DP_OP_19_294_9081/n7 ) );
  AOI21X1 \DP_OP_19_294_9081/U22  ( .A(\DP_OP_19_294_9081/n89 ), .B(n1089), 
        .C(\DP_OP_19_294_9081/n82 ), .Y(\DP_OP_19_294_9081/n80 ) );
  NAND2X1 \DP_OP_19_294_9081/U21  ( .A(n1089), .B(\DP_OP_19_294_9081/n88 ), 
        .Y(\DP_OP_19_294_9081/n79 ) );
  OAI21X1 \DP_OP_19_294_9081/U20  ( .A(\DP_OP_19_294_9081/n79 ), .B(
        \DP_OP_19_294_9081/n100 ), .C(\DP_OP_19_294_9081/n80 ), .Y(
        \DP_OP_19_294_9081/n78 ) );
  NOR2X1 \DP_OP_19_294_9081/U19  ( .A(\DP_OP_19_294_9081/n79 ), .B(
        \DP_OP_19_294_9081/n99 ), .Y(\DP_OP_19_294_9081/n77 ) );
  AOI21X1 \DP_OP_19_294_9081/U18  ( .A(\DP_OP_19_294_9081/n77 ), .B(
        \DP_OP_19_294_9081/n128 ), .C(\DP_OP_19_294_9081/n78 ), .Y(
        \DP_OP_19_294_9081/n76 ) );
  NAND2X1 \DP_OP_19_294_9081/U17  ( .A(\DP_OP_19_294_9081/n77 ), .B(
        \DP_OP_19_294_9081/n127 ), .Y(\DP_OP_19_294_9081/n75 ) );
  OAI21X1 \DP_OP_19_294_9081/U16  ( .A(\DP_OP_19_294_9081/n75 ), .B(
        \DP_OP_19_294_9081/n3 ), .C(\DP_OP_19_294_9081/n76 ), .Y(
        \DP_OP_19_294_9081/n74 ) );
  NOR2X1 \DP_OP_19_294_9081/U15  ( .A(\DP_OP_19_294_9081/n75 ), .B(
        \DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n73 ) );
  AOI21X1 \DP_OP_19_294_9081/U14  ( .A(n1064), .B(\DP_OP_19_294_9081/n73 ), 
        .C(\DP_OP_19_294_9081/n74 ), .Y(\DP_OP_19_294_9081/n72 ) );
  NAND2X1 \DP_OP_19_294_9081/U12  ( .A(\C2/Z_62 ), .B(\DP_OP_19_294_9081/n715 ), .Y(\DP_OP_19_294_9081/n71 ) );
  NOR2X1 \DP_OP_19_294_9081/U11  ( .A(\C2/Z_62 ), .B(\DP_OP_19_294_9081/n715 ), 
        .Y(\DP_OP_19_294_9081/n70 ) );
  NAND2X1 \DP_OP_19_294_9081/U9  ( .A(\DP_OP_19_294_9081/n71 ), .B(
        \DP_OP_19_294_9081/n458 ), .Y(\DP_OP_19_294_9081/n6 ) );
  OAI21X1 \DP_OP_19_294_9081/U8  ( .A(\DP_OP_19_294_9081/n70 ), .B(
        \DP_OP_19_294_9081/n72 ), .C(\DP_OP_19_294_9081/n71 ), .Y(
        \DP_OP_19_294_9081/n69 ) );
  XOR2X1 \DP_OP_19_294_9081/U6  ( .A(\DP_OP_19_294_9081/n716 ), .B(\C2/Z_63 ), 
        .Y(\DP_OP_19_294_9081/n5 ) );
  INVX1 U627 ( .A(n634), .Y(n624) );
  INVX1 U598 ( .A(n663), .Y(n595) );
  INVX1 U616 ( .A(n645), .Y(n613) );
  INVX1 U615 ( .A(n646), .Y(n612) );
  INVX1 U628 ( .A(n633), .Y(n625) );
  INVX1 U611 ( .A(n650), .Y(n608) );
  INVX1 U607 ( .A(n654), .Y(n604) );
  INVX1 U624 ( .A(n637), .Y(n621) );
  INVX1 U626 ( .A(n635), .Y(n623) );
  INVX1 U629 ( .A(n631), .Y(n626) );
  INVX1 U609 ( .A(n652), .Y(n606) );
  INVX1 U612 ( .A(n649), .Y(n609) );
  INVX1 U625 ( .A(n636), .Y(n622) );
  INVX1 U608 ( .A(n653), .Y(n605) );
  INVX1 U614 ( .A(n647), .Y(n611) );
  INVX1 U610 ( .A(n651), .Y(n607) );
  INVX1 U613 ( .A(n648), .Y(n610) );
  INVX1 U603 ( .A(n658), .Y(n600) );
  INVX1 U619 ( .A(n642), .Y(n616) );
  INVX1 U621 ( .A(n640), .Y(n618) );
  INVX1 U600 ( .A(n661), .Y(n597) );
  INVX1 U605 ( .A(n656), .Y(n602) );
  INVX1 U622 ( .A(n639), .Y(n619) );
  INVX1 U618 ( .A(n643), .Y(n615) );
  INVX1 U604 ( .A(n657), .Y(n601) );
  INVX1 U601 ( .A(n660), .Y(n598) );
  INVX1 U599 ( .A(n662), .Y(n596) );
  INVX1 U620 ( .A(n641), .Y(n617) );
  INVX1 U623 ( .A(n638), .Y(n620) );
  INVX1 U602 ( .A(n659), .Y(n599) );
  INVX1 U606 ( .A(n655), .Y(n603) );
  INVX1 U617 ( .A(n644), .Y(n614) );
  OAI21X1 U673 ( .A(n1179), .B(n788), .C(1'b1), .Y(_pushout_d) );
  OAI21X1 U674 ( .A(\DP_OP_19_294_9081/n382 ), .B(\DP_OP_19_294_9081/n401 ), 
        .C(1'b1), .Y(n708) );
  OAI21X1 U675 ( .A(n1179), .B(n445), .C(1'b1), .Y(n706) );
  OAI21X1 U676 ( .A(\DP_OP_19_294_9081/n447 ), .B(\DP_OP_19_294_9081/n450 ), 
        .C(1'b1), .Y(n680) );
  OAI21X1 U677 ( .A(1'b0), .B(h[31]), .C(n1171), .Y(n960) );
  OAI21X1 U678 ( .A(1'b0), .B(h[30]), .C(n1171), .Y(n957) );
  OAI21X1 U679 ( .A(1'b0), .B(h[29]), .C(n1171), .Y(n954) );
  OAI21X1 U680 ( .A(1'b0), .B(h[28]), .C(n1169), .Y(n951) );
  OAI21X1 U681 ( .A(1'b0), .B(h[27]), .C(n1171), .Y(n948) );
  OAI21X1 U682 ( .A(1'b0), .B(h[26]), .C(n1171), .Y(n945) );
  OAI21X1 U683 ( .A(1'b0), .B(h[25]), .C(n1170), .Y(n942) );
  OAI21X1 U684 ( .A(1'b0), .B(n1169), .C(h[24]), .Y(n939) );
  OAI21X1 U685 ( .A(1'b0), .B(h[23]), .C(n1170), .Y(n936) );
  OAI21X1 U686 ( .A(1'b0), .B(n1171), .C(h[22]), .Y(n933) );
  OAI21X1 U687 ( .A(1'b0), .B(h[21]), .C(n1171), .Y(n930) );
  OAI21X1 U688 ( .A(1'b0), .B(n1169), .C(h[20]), .Y(n927) );
  OAI21X1 U689 ( .A(1'b0), .B(h[19]), .C(n1169), .Y(n924) );
  OAI21X1 U690 ( .A(1'b0), .B(n1170), .C(h[18]), .Y(n921) );
  OAI21X1 U691 ( .A(1'b0), .B(n1171), .C(h[17]), .Y(n918) );
  OAI21X1 U692 ( .A(1'b0), .B(h[16]), .C(n1170), .Y(n915) );
  OAI21X1 U693 ( .A(1'b0), .B(h[15]), .C(n1171), .Y(n912) );
  OAI21X1 U694 ( .A(1'b0), .B(n1170), .C(h[14]), .Y(n909) );
  OAI21X1 U695 ( .A(1'b0), .B(h[13]), .C(n1170), .Y(n906) );
  OAI21X1 U696 ( .A(1'b0), .B(h[12]), .C(n1170), .Y(n903) );
  OAI21X1 U697 ( .A(1'b0), .B(n1170), .C(h[11]), .Y(n900) );
  OAI21X1 U698 ( .A(1'b0), .B(h[10]), .C(n1169), .Y(n897) );
  OAI21X1 U699 ( .A(1'b0), .B(h[9]), .C(n1171), .Y(n894) );
  OAI21X1 U700 ( .A(1'b0), .B(h[8]), .C(n1169), .Y(n891) );
  OAI21X1 U701 ( .A(1'b0), .B(h[7]), .C(n1169), .Y(n888) );
  OAI21X1 U702 ( .A(1'b0), .B(n1171), .C(h[6]), .Y(n885) );
  OAI21X1 U703 ( .A(1'b0), .B(h[5]), .C(n1169), .Y(n882) );
  OAI21X1 U704 ( .A(1'b0), .B(h[4]), .C(n1170), .Y(n879) );
  OAI21X1 U705 ( .A(1'b0), .B(h[3]), .C(n1169), .Y(n876) );
  OAI21X1 U706 ( .A(1'b0), .B(h[2]), .C(n1170), .Y(n873) );
  OAI21X1 U707 ( .A(1'b0), .B(h[1]), .C(n1171), .Y(n870) );
  OAI21X1 U708 ( .A(1'b0), .B(h[0]), .C(n1171), .Y(n867) );
  OAI21X1 U709 ( .A(1'b0), .B(n1170), .C(q[31]), .Y(n864) );
  OAI21X1 U710 ( .A(1'b0), .B(q[29]), .C(n1169), .Y(n861) );
  OAI21X1 U711 ( .A(1'b0), .B(q[28]), .C(n1170), .Y(n858) );
  OAI21X1 U712 ( .A(1'b0), .B(q[26]), .C(n1170), .Y(n855) );
  OAI21X1 U713 ( .A(1'b0), .B(n1171), .C(q[25]), .Y(n852) );
  OAI21X1 U714 ( .A(1'b0), .B(q[24]), .C(n1171), .Y(n849) );
  OAI21X1 U715 ( .A(1'b0), .B(q[22]), .C(n1170), .Y(n846) );
  OAI21X1 U716 ( .A(1'b0), .B(q[20]), .C(n1170), .Y(n843) );
  OAI21X1 U717 ( .A(1'b0), .B(q[19]), .C(n1171), .Y(n840) );
  OAI21X1 U718 ( .A(1'b0), .B(n1169), .C(q[18]), .Y(n837) );
  OAI21X1 U719 ( .A(1'b0), .B(q[17]), .C(n1170), .Y(n834) );
  OAI21X1 U720 ( .A(1'b0), .B(q[16]), .C(n1170), .Y(n831) );
  OAI21X1 U721 ( .A(1'b0), .B(n1170), .C(q[14]), .Y(n828) );
  OAI21X1 U722 ( .A(1'b0), .B(n1170), .C(q[13]), .Y(n825) );
  OAI21X1 U723 ( .A(1'b0), .B(q[12]), .C(n1169), .Y(n822) );
  OAI21X1 U724 ( .A(1'b0), .B(q[10]), .C(n1169), .Y(n819) );
  OAI21X1 U725 ( .A(1'b0), .B(n1169), .C(q[9]), .Y(n816) );
  OAI21X1 U726 ( .A(1'b0), .B(n1171), .C(q[8]), .Y(n813) );
  OAI21X1 U727 ( .A(1'b0), .B(q[7]), .C(n1169), .Y(n810) );
  OAI21X1 U728 ( .A(1'b0), .B(n1171), .C(q[6]), .Y(n807) );
  OAI21X1 U729 ( .A(1'b0), .B(n1171), .C(q[4]), .Y(n804) );
  OAI21X1 U730 ( .A(1'b0), .B(n1169), .C(q[3]), .Y(n801) );
  OAI21X1 U731 ( .A(1'b0), .B(q[2]), .C(n1169), .Y(n798) );
  OAI21X1 U732 ( .A(1'b0), .B(q[1]), .C(n1169), .Y(n795) );
  OAI21X1 U733 ( .A(1'b0), .B(q[0]), .C(n1170), .Y(n792) );
  OAI21X1 U734 ( .A(1'b0), .B(n1376), .C(n1377), .Y(n788) );
  OAI21X1 U735 ( .A(1'b0), .B(N82), .C(n1302), .Y(n753) );
  OAI21X1 U736 ( .A(1'b0), .B(N84), .C(n1302), .Y(n750) );
  OAI21X1 U737 ( .A(1'b0), .B(n630), .C(h1[5]), .Y(n747) );
  OAI21X1 U738 ( .A(1'b0), .B(n630), .C(h1[4]), .Y(n745) );
  OAI21X1 U739 ( .A(1'b0), .B(n630), .C(h1[3]), .Y(n743) );
  OAI21X1 U740 ( .A(1'b0), .B(n630), .C(h1[0]), .Y(n741) );
  OAI21X1 U741 ( .A(1'b0), .B(q[30]), .C(n1169), .Y(n738) );
  OAI21X1 U742 ( .A(1'b0), .B(q[27]), .C(n1171), .Y(n735) );
  OAI21X1 U743 ( .A(1'b0), .B(n1170), .C(q[23]), .Y(n732) );
  OAI21X1 U744 ( .A(1'b0), .B(q[21]), .C(n1169), .Y(n729) );
  OAI21X1 U745 ( .A(1'b0), .B(q[15]), .C(n1169), .Y(n726) );
  OAI21X1 U746 ( .A(1'b0), .B(n1170), .C(q[11]), .Y(n723) );
  OAI21X1 U747 ( .A(1'b0), .B(q[5]), .C(n1171), .Y(n720) );
  OAI21X1 U748 ( .A(1'b0), .B(\DP_OP_19_294_9081/n451 ), .C(
        \DP_OP_19_294_9081/n518 ), .Y(n714) );
  OAI21X1 U749 ( .A(1'b0), .B(n1162), .C(\ashr_28_1/n584 ), .Y(n699) );
  OAI21X1 U750 ( .A(1'b0), .B(\DP_OP_19_294_9081/n448 ), .C(
        \DP_OP_19_294_9081/n517 ), .Y(n692) );
  OAI21X1 U751 ( .A(1'b0), .B(n1163), .C(\ashr_28_1/n585 ), .Y(n684) );
  OAI21X1 U752 ( .A(1'b0), .B(N83), .C(n1302), .Y(n677) );
  OAI21X1 U753 ( .A(1'b0), .B(n1164), .C(\ashr_28_1/n586 ), .Y(n674) );
  INVX2 U754 ( .A(n1166), .Y(n961) );
  BUFX2 U755 ( .A(h2[0]), .Y(n1165) );
  INVX4 U756 ( .A(n1304), .Y(n1302) );
  INVX2 U757 ( .A(n1173), .Y(n1066) );
  INVX4 U758 ( .A(n1173), .Y(n1174) );
  INVX2 U759 ( .A(n1065), .Y(n962) );
  INVX2 U760 ( .A(n1065), .Y(n963) );
  INVX2 U761 ( .A(n1065), .Y(n964) );
  INVX1 U762 ( .A(\ashr_28_1/n584 ), .Y(n672) );
  OAI21X1 U764 ( .A(n1164), .B(n672), .C(n674), .Y(N84) );
  INVX1 U765 ( .A(mulout[2]), .Y(n675) );
  OAI21X1 U767 ( .A(n1066), .B(n675), .C(n677), .Y(\DP_OP_19_294_9081/n655 )
         );
  INVX1 U768 ( .A(push_2), .Y(n678) );
  AOI21X1 U769 ( .A(n1304), .B(n1175), .C(n678), .Y(n1172) );
  OAI21X1 U771 ( .A(\DP_OP_19_294_9081/n447 ), .B(\DP_OP_19_294_9081/n451 ), 
        .C(\DP_OP_19_294_9081/n448 ), .Y(n681) );
  AOI21X1 U772 ( .A(\DP_OP_19_294_9081/n453 ), .B(n680), .C(n681), .Y(
        \DP_OP_19_294_9081/n444 ) );
  INVX1 U773 ( .A(\ashr_28_1/n583 ), .Y(n682) );
  OAI21X1 U775 ( .A(n1163), .B(n682), .C(n684), .Y(N83) );
  INVX1 U776 ( .A(mulout[40]), .Y(n685) );
  INVX1 U777 ( .A(n1161), .Y(n686) );
  OAI21X1 U778 ( .A(\ashr_28_1/n623 ), .B(n1161), .C(n1302), .Y(n687) );
  INVX1 U779 ( .A(n687), .Y(n688) );
  OAI21X1 U780 ( .A(\ashr_28_1/n621 ), .B(n686), .C(n688), .Y(n689) );
  OAI21X1 U781 ( .A(n1174), .B(n685), .C(n689), .Y(\DP_OP_19_294_9081/n693 )
         );
  INVX1 U782 ( .A(n1302), .Y(n690) );
  OAI22X1 U783 ( .A(n1174), .B(n1303), .C(n1090), .D(n690), .Y(
        \DP_OP_19_294_9081/n589 ) );
  OAI21X1 U785 ( .A(push_2), .B(n1299), .C(n1369), .Y(n693) );
  NAND2X1 U786 ( .A(n692), .B(\DP_OP_19_294_9081/n449 ), .Y(n694) );
  OAI21X1 U787 ( .A(n692), .B(\DP_OP_19_294_9081/n449 ), .C(n694), .Y(n695) );
  AOI21X1 U788 ( .A(n1172), .B(n695), .C(n693), .Y(n696) );
  INVX1 U789 ( .A(n696), .Y(n430) );
  INVX1 U790 ( .A(\ashr_28_1/n582 ), .Y(n697) );
  OAI21X1 U792 ( .A(n1162), .B(n697), .C(n699), .Y(N82) );
  INVX1 U793 ( .A(mulout[61]), .Y(n700) );
  INVX1 U794 ( .A(n1161), .Y(n701) );
  OAI21X1 U795 ( .A(\ashr_28_1/n644 ), .B(n1161), .C(n1302), .Y(n702) );
  INVX1 U796 ( .A(n702), .Y(n703) );
  OAI21X1 U797 ( .A(\ashr_28_1/n642 ), .B(n701), .C(n703), .Y(n704) );
  OAI21X1 U798 ( .A(n1174), .B(n700), .C(n704), .Y(\DP_OP_19_294_9081/n714 )
         );
  AND2X2 U800 ( .A(n706), .B(n1304), .Y(n1378) );
  OAI21X1 U802 ( .A(\DP_OP_19_294_9081/n382 ), .B(\DP_OP_19_294_9081/n402 ), 
        .C(\DP_OP_19_294_9081/n383 ), .Y(n709) );
  AOI21X1 U803 ( .A(\DP_OP_19_294_9081/n423 ), .B(n708), .C(n709), .Y(
        \DP_OP_19_294_9081/n1 ) );
  AND2X1 U804 ( .A(\DP_OP_19_294_9081/n479 ), .B(\DP_OP_19_294_9081/n232 ), 
        .Y(n710) );
  NAND2X1 U805 ( .A(\DP_OP_19_294_9081/n233 ), .B(n710), .Y(n711) );
  OAI21X1 U806 ( .A(\DP_OP_19_294_9081/n233 ), .B(n710), .C(n711), .Y(n712) );
  OAI21X1 U807 ( .A(n1176), .B(n712), .C(n1028), .Y(n325) );
  OAI21X1 U809 ( .A(\DP_OP_19_294_9081/n452 ), .B(n714), .C(n1172), .Y(n715)
         );
  AOI21X1 U810 ( .A(\DP_OP_19_294_9081/n452 ), .B(n714), .C(n715), .Y(n716) );
  OAI21X1 U811 ( .A(push_2), .B(n1300), .C(n1370), .Y(n717) );
  OR2X1 U812 ( .A(n716), .B(n717), .Y(n433) );
  INVX1 U813 ( .A(q0[5]), .Y(n718) );
  OAI21X1 U815 ( .A(n1170), .B(n718), .C(n720), .Y(n457) );
  INVX1 U816 ( .A(q0[11]), .Y(n721) );
  OAI21X1 U818 ( .A(n1170), .B(n721), .C(n723), .Y(n469) );
  INVX1 U819 ( .A(q0[15]), .Y(n724) );
  OAI21X1 U821 ( .A(n1171), .B(n724), .C(n726), .Y(n477) );
  INVX1 U822 ( .A(q0[21]), .Y(n727) );
  OAI21X1 U824 ( .A(n1170), .B(n727), .C(n729), .Y(n489) );
  INVX1 U825 ( .A(q0[23]), .Y(n730) );
  OAI21X1 U827 ( .A(n1170), .B(n730), .C(n732), .Y(n493) );
  INVX1 U828 ( .A(q0[27]), .Y(n733) );
  OAI21X1 U830 ( .A(n1169), .B(n733), .C(n735), .Y(n501) );
  INVX1 U831 ( .A(q0[30]), .Y(n736) );
  OAI21X1 U833 ( .A(n1170), .B(n736), .C(n738), .Y(n507) );
  INVX1 U834 ( .A(h2[0]), .Y(n739) );
  OAI21X1 U836 ( .A(n630), .B(n739), .C(n741), .Y(n511) );
  OAI21X1 U838 ( .A(n630), .B(n1168), .C(n743), .Y(n514) );
  OAI21X1 U840 ( .A(n630), .B(n1154), .C(n745), .Y(n515) );
  OAI21X1 U842 ( .A(n630), .B(n1182), .C(n747), .Y(n516) );
  INVX1 U843 ( .A(mulout[3]), .Y(n748) );
  OAI21X1 U845 ( .A(n1066), .B(n748), .C(n750), .Y(\DP_OP_19_294_9081/n656 )
         );
  INVX1 U846 ( .A(mulout[1]), .Y(n751) );
  OAI21X1 U848 ( .A(n1066), .B(n751), .C(n753), .Y(\DP_OP_19_294_9081/n654 )
         );
  INVX1 U849 ( .A(mulout[31]), .Y(n754) );
  INVX1 U850 ( .A(n1163), .Y(n755) );
  OAI21X1 U851 ( .A(\ashr_28_1/n612 ), .B(n1163), .C(n1302), .Y(n756) );
  INVX1 U852 ( .A(n756), .Y(n757) );
  OAI21X1 U853 ( .A(\ashr_28_1/n614 ), .B(n755), .C(n757), .Y(n758) );
  OAI21X1 U854 ( .A(n1066), .B(n754), .C(n758), .Y(\DP_OP_19_294_9081/n684 )
         );
  INVX1 U855 ( .A(mulout[63]), .Y(n759) );
  NAND3X1 U856 ( .A(n1161), .B(n1302), .C(\ashr_28_1/n644 ), .Y(n760) );
  OAI21X1 U857 ( .A(n1066), .B(n759), .C(n760), .Y(\DP_OP_19_294_9081/n716 )
         );
  AND2X1 U858 ( .A(\DP_OP_19_294_9081/n471 ), .B(\DP_OP_19_294_9081/n176 ), 
        .Y(n761) );
  NAND2X1 U859 ( .A(\DP_OP_19_294_9081/n177 ), .B(n761), .Y(n762) );
  OAI21X1 U860 ( .A(\DP_OP_19_294_9081/n177 ), .B(n761), .C(n762), .Y(n763) );
  OAI21X1 U861 ( .A(n1176), .B(n763), .C(n1024), .Y(n309) );
  AND2X1 U862 ( .A(\DP_OP_19_294_9081/n475 ), .B(\DP_OP_19_294_9081/n204 ), 
        .Y(n764) );
  NAND2X1 U863 ( .A(\DP_OP_19_294_9081/n205 ), .B(n764), .Y(n765) );
  OAI21X1 U864 ( .A(\DP_OP_19_294_9081/n205 ), .B(n764), .C(n765), .Y(n766) );
  OAI21X1 U865 ( .A(n1176), .B(n766), .C(n1026), .Y(n317) );
  AND2X1 U866 ( .A(\DP_OP_19_294_9081/n477 ), .B(\DP_OP_19_294_9081/n220 ), 
        .Y(n767) );
  NAND2X1 U867 ( .A(\DP_OP_19_294_9081/n221 ), .B(n767), .Y(n768) );
  OAI21X1 U868 ( .A(\DP_OP_19_294_9081/n221 ), .B(n767), .C(n768), .Y(n769) );
  OAI21X1 U869 ( .A(n1176), .B(n769), .C(n1027), .Y(n321) );
  INVX1 U870 ( .A(\DP_OP_19_294_9081/n234 ), .Y(n770) );
  NAND2X1 U871 ( .A(n770), .B(\DP_OP_19_294_9081/n235 ), .Y(n771) );
  NAND2X1 U872 ( .A(\DP_OP_19_294_9081/n236 ), .B(n771), .Y(n772) );
  OAI21X1 U873 ( .A(\DP_OP_19_294_9081/n236 ), .B(n771), .C(n772), .Y(n773) );
  OAI21X1 U874 ( .A(n1176), .B(n773), .C(n1029), .Y(n327) );
  AND2X1 U875 ( .A(\DP_OP_19_294_9081/n481 ), .B(\DP_OP_19_294_9081/n248 ), 
        .Y(n774) );
  NAND2X1 U876 ( .A(\DP_OP_19_294_9081/n249 ), .B(n774), .Y(n775) );
  OAI21X1 U877 ( .A(\DP_OP_19_294_9081/n249 ), .B(n774), .C(n775), .Y(n776) );
  OAI21X1 U878 ( .A(n1176), .B(n776), .C(n1030), .Y(n329) );
  AND2X1 U879 ( .A(\DP_OP_19_294_9081/n483 ), .B(\DP_OP_19_294_9081/n260 ), 
        .Y(n777) );
  NAND2X1 U880 ( .A(\DP_OP_19_294_9081/n261 ), .B(n777), .Y(n778) );
  OAI21X1 U881 ( .A(\DP_OP_19_294_9081/n261 ), .B(n777), .C(n778), .Y(n779) );
  OAI21X1 U882 ( .A(n1176), .B(n779), .C(n1031), .Y(n333) );
  AND2X1 U883 ( .A(\DP_OP_19_294_9081/n487 ), .B(\DP_OP_19_294_9081/n284 ), 
        .Y(n780) );
  NAND2X1 U884 ( .A(\DP_OP_19_294_9081/n285 ), .B(n780), .Y(n781) );
  OAI21X1 U885 ( .A(\DP_OP_19_294_9081/n285 ), .B(n780), .C(n781), .Y(n782) );
  OAI21X1 U886 ( .A(n1176), .B(n782), .C(n1033), .Y(n341) );
  INVX1 U887 ( .A(n1172), .Y(n783) );
  OAI21X1 U888 ( .A(\DP_OP_19_294_9081/n653 ), .B(\DP_OP_19_294_9081/n589 ), 
        .C(\DP_OP_19_294_9081/n457 ), .Y(n784) );
  OAI21X1 U889 ( .A(n1303), .B(push_2), .C(n1375), .Y(n785) );
  INVX1 U890 ( .A(n785), .Y(n786) );
  OAI21X1 U891 ( .A(n783), .B(n784), .C(n786), .Y(n439) );
  INVX1 U894 ( .A(q0[0]), .Y(n790) );
  OAI21X1 U896 ( .A(n1171), .B(n790), .C(n792), .Y(n447) );
  INVX1 U897 ( .A(q0[1]), .Y(n793) );
  OAI21X1 U899 ( .A(n1171), .B(n793), .C(n795), .Y(n449) );
  INVX1 U900 ( .A(q0[2]), .Y(n796) );
  OAI21X1 U902 ( .A(n1170), .B(n796), .C(n798), .Y(n451) );
  INVX1 U903 ( .A(q0[3]), .Y(n799) );
  OAI21X1 U905 ( .A(n1169), .B(n799), .C(n801), .Y(n453) );
  INVX1 U906 ( .A(q0[4]), .Y(n802) );
  OAI21X1 U908 ( .A(n1171), .B(n802), .C(n804), .Y(n455) );
  INVX1 U909 ( .A(q0[6]), .Y(n805) );
  OAI21X1 U911 ( .A(n1171), .B(n805), .C(n807), .Y(n459) );
  INVX1 U912 ( .A(q0[7]), .Y(n808) );
  OAI21X1 U914 ( .A(n1171), .B(n808), .C(n810), .Y(n461) );
  INVX1 U915 ( .A(q0[8]), .Y(n811) );
  OAI21X1 U917 ( .A(n1171), .B(n811), .C(n813), .Y(n463) );
  INVX1 U918 ( .A(q0[9]), .Y(n814) );
  OAI21X1 U920 ( .A(n1169), .B(n814), .C(n816), .Y(n465) );
  INVX1 U921 ( .A(q0[10]), .Y(n817) );
  OAI21X1 U923 ( .A(n1171), .B(n817), .C(n819), .Y(n467) );
  INVX1 U924 ( .A(q0[12]), .Y(n820) );
  OAI21X1 U926 ( .A(n1171), .B(n820), .C(n822), .Y(n471) );
  INVX1 U927 ( .A(q0[13]), .Y(n823) );
  OAI21X1 U929 ( .A(n1170), .B(n823), .C(n825), .Y(n473) );
  INVX1 U930 ( .A(q0[14]), .Y(n826) );
  OAI21X1 U932 ( .A(n1170), .B(n826), .C(n828), .Y(n475) );
  INVX1 U933 ( .A(q0[16]), .Y(n829) );
  OAI21X1 U935 ( .A(n1169), .B(n829), .C(n831), .Y(n479) );
  INVX1 U936 ( .A(q0[17]), .Y(n832) );
  OAI21X1 U938 ( .A(n1171), .B(n832), .C(n834), .Y(n481) );
  INVX1 U939 ( .A(q0[18]), .Y(n835) );
  OAI21X1 U941 ( .A(n1169), .B(n835), .C(n837), .Y(n483) );
  INVX1 U942 ( .A(q0[19]), .Y(n838) );
  OAI21X1 U944 ( .A(n1170), .B(n838), .C(n840), .Y(n485) );
  INVX1 U945 ( .A(q0[20]), .Y(n841) );
  OAI21X1 U947 ( .A(n1171), .B(n841), .C(n843), .Y(n487) );
  INVX1 U948 ( .A(q0[22]), .Y(n844) );
  OAI21X1 U950 ( .A(n1169), .B(n844), .C(n846), .Y(n491) );
  INVX1 U951 ( .A(q0[24]), .Y(n847) );
  OAI21X1 U953 ( .A(n1169), .B(n847), .C(n849), .Y(n495) );
  INVX1 U954 ( .A(q0[25]), .Y(n850) );
  OAI21X1 U956 ( .A(n1171), .B(n850), .C(n852), .Y(n497) );
  INVX1 U957 ( .A(q0[26]), .Y(n853) );
  OAI21X1 U959 ( .A(n1169), .B(n853), .C(n855), .Y(n499) );
  INVX1 U960 ( .A(q0[28]), .Y(n856) );
  OAI21X1 U962 ( .A(n1169), .B(n856), .C(n858), .Y(n503) );
  INVX1 U963 ( .A(q0[29]), .Y(n859) );
  OAI21X1 U965 ( .A(n1171), .B(n859), .C(n861), .Y(n505) );
  INVX1 U966 ( .A(q0[31]), .Y(n862) );
  OAI21X1 U968 ( .A(n1170), .B(n862), .C(n864), .Y(n509) );
  INVX1 U969 ( .A(h0[0]), .Y(n865) );
  OAI21X1 U971 ( .A(n1169), .B(n865), .C(n867), .Y(n524) );
  INVX1 U972 ( .A(h0[1]), .Y(n868) );
  OAI21X1 U974 ( .A(n1170), .B(n868), .C(n870), .Y(n527) );
  INVX1 U975 ( .A(h0[2]), .Y(n871) );
  OAI21X1 U977 ( .A(n1171), .B(n871), .C(n873), .Y(n530) );
  INVX1 U978 ( .A(h0[3]), .Y(n874) );
  OAI21X1 U980 ( .A(n1171), .B(n874), .C(n876), .Y(n533) );
  INVX1 U981 ( .A(h0[4]), .Y(n877) );
  OAI21X1 U983 ( .A(n1169), .B(n877), .C(n879), .Y(n536) );
  INVX1 U984 ( .A(h0[5]), .Y(n880) );
  OAI21X1 U986 ( .A(n1171), .B(n880), .C(n882), .Y(n539) );
  INVX1 U987 ( .A(h0[6]), .Y(n883) );
  OAI21X1 U989 ( .A(n1171), .B(n883), .C(n885), .Y(n542) );
  INVX1 U990 ( .A(h0[7]), .Y(n886) );
  OAI21X1 U992 ( .A(n1171), .B(n886), .C(n888), .Y(n544) );
  INVX1 U993 ( .A(h0[8]), .Y(n889) );
  OAI21X1 U995 ( .A(n1170), .B(n889), .C(n891), .Y(n546) );
  INVX1 U996 ( .A(h0[9]), .Y(n892) );
  OAI21X1 U998 ( .A(n1170), .B(n892), .C(n894), .Y(n548) );
  INVX1 U999 ( .A(h0[10]), .Y(n895) );
  OAI21X1 U1001 ( .A(n1170), .B(n895), .C(n897), .Y(n550) );
  INVX1 U1002 ( .A(h0[11]), .Y(n898) );
  OAI21X1 U1004 ( .A(n1170), .B(n898), .C(n900), .Y(n552) );
  INVX1 U1005 ( .A(h0[12]), .Y(n901) );
  OAI21X1 U1007 ( .A(n1169), .B(n901), .C(n903), .Y(n554) );
  INVX1 U1008 ( .A(h0[13]), .Y(n904) );
  OAI21X1 U1010 ( .A(n1171), .B(n904), .C(n906), .Y(n556) );
  INVX1 U1011 ( .A(h0[14]), .Y(n907) );
  OAI21X1 U1013 ( .A(n1170), .B(n907), .C(n909), .Y(n558) );
  INVX1 U1014 ( .A(h0[15]), .Y(n910) );
  OAI21X1 U1016 ( .A(n1170), .B(n910), .C(n912), .Y(n560) );
  INVX1 U1017 ( .A(h0[16]), .Y(n913) );
  OAI21X1 U1019 ( .A(n1169), .B(n913), .C(n915), .Y(n562) );
  INVX1 U1020 ( .A(h0[17]), .Y(n916) );
  OAI21X1 U1022 ( .A(n1171), .B(n916), .C(n918), .Y(n564) );
  INVX1 U1023 ( .A(h0[18]), .Y(n919) );
  OAI21X1 U1025 ( .A(n1170), .B(n919), .C(n921), .Y(n566) );
  INVX1 U1026 ( .A(h0[19]), .Y(n922) );
  OAI21X1 U1028 ( .A(n1170), .B(n922), .C(n924), .Y(n568) );
  INVX1 U1029 ( .A(h0[20]), .Y(n925) );
  OAI21X1 U1031 ( .A(n1169), .B(n925), .C(n927), .Y(n570) );
  INVX1 U1032 ( .A(h0[21]), .Y(n928) );
  OAI21X1 U1034 ( .A(n1169), .B(n928), .C(n930), .Y(n572) );
  INVX1 U1035 ( .A(h0[22]), .Y(n931) );
  OAI21X1 U1037 ( .A(n1171), .B(n931), .C(n933), .Y(n574) );
  INVX1 U1038 ( .A(h0[23]), .Y(n934) );
  OAI21X1 U1040 ( .A(n1169), .B(n934), .C(n936), .Y(n576) );
  INVX1 U1041 ( .A(h0[24]), .Y(n937) );
  OAI21X1 U1043 ( .A(n1169), .B(n937), .C(n939), .Y(n578) );
  INVX1 U1044 ( .A(h0[25]), .Y(n940) );
  OAI21X1 U1046 ( .A(n1169), .B(n940), .C(n942), .Y(n580) );
  INVX1 U1047 ( .A(h0[26]), .Y(n943) );
  OAI21X1 U1049 ( .A(n1170), .B(n943), .C(n945), .Y(n582) );
  INVX1 U1050 ( .A(h0[27]), .Y(n946) );
  OAI21X1 U1052 ( .A(n1169), .B(n946), .C(n948), .Y(n584) );
  INVX1 U1053 ( .A(h0[28]), .Y(n949) );
  OAI21X1 U1055 ( .A(n1171), .B(n949), .C(n951), .Y(n586) );
  INVX1 U1056 ( .A(h0[29]), .Y(n952) );
  OAI21X1 U1058 ( .A(n1169), .B(n952), .C(n954), .Y(n588) );
  INVX1 U1059 ( .A(h0[30]), .Y(n955) );
  OAI21X1 U1061 ( .A(n1170), .B(n955), .C(n957), .Y(n590) );
  INVX1 U1062 ( .A(h0[31]), .Y(n958) );
  OAI21X1 U1064 ( .A(n1169), .B(n958), .C(n960), .Y(n592) );
  INVX8 U1065 ( .A(\ashr_28_1/SH[5] ), .Y(n1151) );
  MUX2X1 U1066 ( .B(\ashr_28_1/n649 ), .A(\ashr_28_1/n648 ), .S(n961), .Y(
        \ashr_28_1/n583 ) );
  MUX2X1 U1067 ( .B(\ashr_28_1/n875 ), .A(\ashr_28_1/n859 ), .S(n962), .Y(
        \ashr_28_1/n794 ) );
  MUX2X1 U1068 ( .B(\ashr_28_1/n879 ), .A(\ashr_28_1/n863 ), .S(n963), .Y(
        \ashr_28_1/n798 ) );
  MUX2X1 U1069 ( .B(\ashr_28_1/n877 ), .A(\ashr_28_1/n861 ), .S(n964), .Y(
        \ashr_28_1/n796 ) );
  INVX4 U1070 ( .A(h2[1]), .Y(n1161) );
  BUFX2 U1071 ( .A(pushin), .Y(n1171) );
  BUFX2 U1072 ( .A(pushin), .Y(n1170) );
  BUFX2 U1073 ( .A(pushin), .Y(n1169) );
  XOR2X1 U1074 ( .A(\DP_OP_19_294_9081/n85 ), .B(\DP_OP_19_294_9081/n7 ), .Y(
        n965) );
  XOR2X1 U1075 ( .A(\DP_OP_19_294_9081/n388 ), .B(\DP_OP_19_294_9081/n53 ), 
        .Y(n966) );
  XOR2X1 U1076 ( .A(\DP_OP_19_294_9081/n105 ), .B(\DP_OP_19_294_9081/n9 ), .Y(
        n967) );
  XOR2X1 U1077 ( .A(\DP_OP_19_294_9081/n119 ), .B(\DP_OP_19_294_9081/n11 ), 
        .Y(n968) );
  XOR2X1 U1078 ( .A(\DP_OP_19_294_9081/n135 ), .B(\DP_OP_19_294_9081/n13 ), 
        .Y(n969) );
  XOR2X1 U1079 ( .A(\DP_OP_19_294_9081/n149 ), .B(\DP_OP_19_294_9081/n15 ), 
        .Y(n970) );
  XOR2X1 U1080 ( .A(\DP_OP_19_294_9081/n165 ), .B(\DP_OP_19_294_9081/n17 ), 
        .Y(n971) );
  XOR2X1 U1081 ( .A(\DP_OP_19_294_9081/n193 ), .B(\DP_OP_19_294_9081/n21 ), 
        .Y(n972) );
  XOR2X1 U1082 ( .A(\DP_OP_19_294_9081/n323 ), .B(\DP_OP_19_294_9081/n41 ), 
        .Y(n973) );
  XOR2X1 U1083 ( .A(\DP_OP_19_294_9081/n331 ), .B(\DP_OP_19_294_9081/n43 ), 
        .Y(n974) );
  XOR2X1 U1084 ( .A(\DP_OP_19_294_9081/n346 ), .B(\DP_OP_19_294_9081/n45 ), 
        .Y(n975) );
  XOR2X1 U1085 ( .A(\DP_OP_19_294_9081/n354 ), .B(\DP_OP_19_294_9081/n47 ), 
        .Y(n976) );
  XOR2X1 U1086 ( .A(\DP_OP_19_294_9081/n365 ), .B(\DP_OP_19_294_9081/n49 ), 
        .Y(n977) );
  XOR2X1 U1087 ( .A(\DP_OP_19_294_9081/n300 ), .B(\DP_OP_19_294_9081/n37 ), 
        .Y(n978) );
  XOR2X1 U1088 ( .A(\DP_OP_19_294_9081/n308 ), .B(\DP_OP_19_294_9081/n39 ), 
        .Y(n979) );
  XOR2X1 U1089 ( .A(\DP_OP_19_294_9081/n396 ), .B(\DP_OP_19_294_9081/n55 ), 
        .Y(n980) );
  XOR2X1 U1090 ( .A(\DP_OP_19_294_9081/n430 ), .B(\DP_OP_19_294_9081/n61 ), 
        .Y(n981) );
  XOR2X1 U1091 ( .A(\DP_OP_19_294_9081/n277 ), .B(\DP_OP_19_294_9081/n33 ), 
        .Y(n982) );
  XOR2X1 U1092 ( .A(\DP_OP_19_294_9081/n419 ), .B(\DP_OP_19_294_9081/n59 ), 
        .Y(n983) );
  XOR2X1 U1093 ( .A(\DP_OP_19_294_9081/n412 ), .B(\DP_OP_19_294_9081/n58 ), 
        .Y(n984) );
  XNOR2X1 U1094 ( .A(\DP_OP_19_294_9081/n422 ), .B(\DP_OP_19_294_9081/n60 ), 
        .Y(n985) );
  XOR2X1 U1095 ( .A(\DP_OP_19_294_9081/n443 ), .B(\DP_OP_19_294_9081/n64 ), 
        .Y(n986) );
  XNOR2X1 U1096 ( .A(\DP_OP_19_294_9081/n311 ), .B(\DP_OP_19_294_9081/n40 ), 
        .Y(n987) );
  XNOR2X1 U1097 ( .A(\DP_OP_19_294_9081/n334 ), .B(\DP_OP_19_294_9081/n44 ), 
        .Y(n988) );
  XNOR2X1 U1098 ( .A(\DP_OP_19_294_9081/n357 ), .B(\DP_OP_19_294_9081/n48 ), 
        .Y(n989) );
  XNOR2X1 U1099 ( .A(\DP_OP_19_294_9081/n399 ), .B(\DP_OP_19_294_9081/n56 ), 
        .Y(n990) );
  XNOR2X1 U1100 ( .A(\DP_OP_19_294_9081/n69 ), .B(\DP_OP_19_294_9081/n5 ), .Y(
        n991) );
  XNOR2X1 U1101 ( .A(\DP_OP_19_294_9081/n407 ), .B(\DP_OP_19_294_9081/n57 ), 
        .Y(n992) );
  XNOR2X1 U1102 ( .A(\DP_OP_19_294_9081/n438 ), .B(\DP_OP_19_294_9081/n63 ), 
        .Y(n993) );
  XNOR2X1 U1103 ( .A(\DP_OP_19_294_9081/n373 ), .B(\DP_OP_19_294_9081/n51 ), 
        .Y(n994) );
  XNOR2X1 U1104 ( .A(\DP_OP_19_294_9081/n288 ), .B(\DP_OP_19_294_9081/n36 ), 
        .Y(n995) );
  XNOR2X1 U1105 ( .A(\DP_OP_19_294_9081/n208 ), .B(\DP_OP_19_294_9081/n24 ), 
        .Y(n996) );
  XNOR2X1 U1106 ( .A(\DP_OP_19_294_9081/n264 ), .B(\DP_OP_19_294_9081/n32 ), 
        .Y(n997) );
  XOR2X1 U1107 ( .A(\DP_OP_19_294_9081/n378 ), .B(\DP_OP_19_294_9081/n52 ), 
        .Y(n998) );
  XNOR2X1 U1108 ( .A(\DP_OP_19_294_9081/n196 ), .B(\DP_OP_19_294_9081/n22 ), 
        .Y(n999) );
  XNOR2X1 U1109 ( .A(\DP_OP_19_294_9081/n224 ), .B(\DP_OP_19_294_9081/n26 ), 
        .Y(n1000) );
  XNOR2X1 U1110 ( .A(\DP_OP_19_294_9081/n252 ), .B(\DP_OP_19_294_9081/n30 ), 
        .Y(n1001) );
  XNOR2X1 U1111 ( .A(\DP_OP_19_294_9081/n180 ), .B(\DP_OP_19_294_9081/n20 ), 
        .Y(n1002) );
  XNOR2X1 U1112 ( .A(\DP_OP_19_294_9081/n108 ), .B(\DP_OP_19_294_9081/n10 ), 
        .Y(n1003) );
  XNOR2X1 U1113 ( .A(\DP_OP_19_294_9081/n72 ), .B(\DP_OP_19_294_9081/n6 ), .Y(
        n1004) );
  XNOR2X1 U1114 ( .A(\DP_OP_19_294_9081/n92 ), .B(\DP_OP_19_294_9081/n8 ), .Y(
        n1005) );
  XNOR2X1 U1115 ( .A(\DP_OP_19_294_9081/n122 ), .B(\DP_OP_19_294_9081/n12 ), 
        .Y(n1006) );
  XNOR2X1 U1116 ( .A(\DP_OP_19_294_9081/n138 ), .B(\DP_OP_19_294_9081/n14 ), 
        .Y(n1007) );
  XNOR2X1 U1117 ( .A(\DP_OP_19_294_9081/n152 ), .B(\DP_OP_19_294_9081/n16 ), 
        .Y(n1008) );
  XNOR2X1 U1118 ( .A(\DP_OP_19_294_9081/n168 ), .B(\DP_OP_19_294_9081/n18 ), 
        .Y(n1009) );
  XNOR2X1 U1119 ( .A(\DP_OP_19_294_9081/n280 ), .B(\DP_OP_19_294_9081/n34 ), 
        .Y(n1010) );
  XNOR2X1 U1120 ( .A(\DP_OP_19_294_9081/n303 ), .B(\DP_OP_19_294_9081/n38 ), 
        .Y(n1011) );
  XNOR2X1 U1121 ( .A(\DP_OP_19_294_9081/n326 ), .B(\DP_OP_19_294_9081/n42 ), 
        .Y(n1012) );
  XNOR2X1 U1122 ( .A(\DP_OP_19_294_9081/n349 ), .B(\DP_OP_19_294_9081/n46 ), 
        .Y(n1013) );
  XNOR2X1 U1123 ( .A(\DP_OP_19_294_9081/n391 ), .B(\DP_OP_19_294_9081/n54 ), 
        .Y(n1014) );
  XNOR2X1 U1124 ( .A(\DP_OP_19_294_9081/n433 ), .B(\DP_OP_19_294_9081/n62 ), 
        .Y(n1015) );
  XNOR2X1 U1125 ( .A(\DP_OP_19_294_9081/n368 ), .B(\DP_OP_19_294_9081/n50 ), 
        .Y(n1016) );
  BUFX2 U1126 ( .A(n1307), .Y(n1017) );
  BUFX2 U1127 ( .A(n1309), .Y(n1018) );
  BUFX2 U1128 ( .A(n1311), .Y(n1019) );
  BUFX2 U1129 ( .A(n1313), .Y(n1020) );
  BUFX2 U1130 ( .A(n1315), .Y(n1021) );
  BUFX2 U1131 ( .A(n1317), .Y(n1022) );
  BUFX2 U1132 ( .A(n1319), .Y(n1023) );
  BUFX2 U1133 ( .A(n1321), .Y(n1024) );
  BUFX2 U1134 ( .A(n1323), .Y(n1025) );
  BUFX2 U1135 ( .A(n1325), .Y(n1026) );
  BUFX2 U1136 ( .A(n1327), .Y(n1027) );
  BUFX2 U1137 ( .A(n1329), .Y(n1028) );
  BUFX2 U1138 ( .A(n1330), .Y(n1029) );
  BUFX2 U1139 ( .A(n1331), .Y(n1030) );
  BUFX2 U1140 ( .A(n1333), .Y(n1031) );
  BUFX2 U1141 ( .A(n1335), .Y(n1032) );
  BUFX2 U1142 ( .A(n1337), .Y(n1033) );
  BUFX2 U1143 ( .A(n346), .Y(n1034) );
  BUFX2 U1144 ( .A(n349), .Y(n1035) );
  BUFX2 U1145 ( .A(n352), .Y(n1036) );
  BUFX2 U1146 ( .A(n355), .Y(n1037) );
  BUFX2 U1147 ( .A(n358), .Y(n1038) );
  BUFX2 U1148 ( .A(n361), .Y(n1039) );
  BUFX2 U1149 ( .A(n364), .Y(n1040) );
  BUFX2 U1150 ( .A(n367), .Y(n1041) );
  BUFX2 U1151 ( .A(n370), .Y(n1042) );
  BUFX2 U1152 ( .A(n373), .Y(n1043) );
  BUFX2 U1153 ( .A(n376), .Y(n1044) );
  BUFX2 U1154 ( .A(n379), .Y(n1045) );
  BUFX2 U1155 ( .A(n385), .Y(n1046) );
  BUFX2 U1156 ( .A(n388), .Y(n1047) );
  BUFX2 U1157 ( .A(n391), .Y(n1048) );
  BUFX2 U1158 ( .A(n394), .Y(n1049) );
  BUFX2 U1159 ( .A(n397), .Y(n1050) );
  BUFX2 U1160 ( .A(n400), .Y(n1051) );
  BUFX2 U1161 ( .A(n403), .Y(n1052) );
  BUFX2 U1162 ( .A(n406), .Y(n1053) );
  BUFX2 U1163 ( .A(n409), .Y(n1054) );
  BUFX2 U1164 ( .A(n412), .Y(n1055) );
  BUFX2 U1165 ( .A(n415), .Y(n1056) );
  BUFX2 U1166 ( .A(n418), .Y(n1057) );
  BUFX2 U1167 ( .A(n421), .Y(n1058) );
  BUFX2 U1168 ( .A(n424), .Y(n1059) );
  BUFX2 U1169 ( .A(n427), .Y(n1060) );
  BUFX2 U1170 ( .A(n512), .Y(n1061) );
  BUFX2 U1171 ( .A(n513), .Y(n1062) );
  BUFX2 U1172 ( .A(n517), .Y(n1063) );
  INVX8 U1173 ( .A(n1088), .Y(n1064) );
  AND2X1 U1174 ( .A(n1173), .B(acc[35]), .Y(\C2/Z_35 ) );
  AND2X1 U1175 ( .A(n1173), .B(acc[37]), .Y(\C2/Z_37 ) );
  AND2X1 U1176 ( .A(n1173), .B(acc[38]), .Y(\C2/Z_38 ) );
  AND2X1 U1177 ( .A(n1173), .B(acc[41]), .Y(\C2/Z_41 ) );
  AND2X1 U1178 ( .A(n1173), .B(acc[43]), .Y(\C2/Z_43 ) );
  AND2X1 U1179 ( .A(n1173), .B(acc[33]), .Y(\C2/Z_33 ) );
  AND2X1 U1180 ( .A(n1173), .B(acc[44]), .Y(\C2/Z_44 ) );
  AND2X1 U1181 ( .A(n1173), .B(acc[21]), .Y(\C2/Z_21 ) );
  AND2X1 U1182 ( .A(n1173), .B(acc[45]), .Y(\C2/Z_45 ) );
  AND2X1 U1183 ( .A(n1173), .B(acc[20]), .Y(\C2/Z_20 ) );
  AND2X1 U1184 ( .A(n1173), .B(acc[19]), .Y(\C2/Z_19 ) );
  AND2X1 U1185 ( .A(n1173), .B(acc[18]), .Y(\C2/Z_18 ) );
  AND2X1 U1186 ( .A(n1173), .B(acc[17]), .Y(\C2/Z_17 ) );
  AND2X1 U1187 ( .A(n1173), .B(acc[15]), .Y(\C2/Z_15 ) );
  INVX4 U1188 ( .A(n1177), .Y(n1178) );
  INVX4 U1189 ( .A(h2[4]), .Y(n1154) );
  INVX2 U1190 ( .A(acc[3]), .Y(n1299) );
  INVX2 U1191 ( .A(h2[6]), .Y(n1147) );
  INVX8 U1192 ( .A(n1154), .Y(n1065) );
  INVX8 U1193 ( .A(rst), .Y(n630) );
  INVX2 U1194 ( .A(\DP_OP_19_294_9081/n2 ), .Y(n1088) );
  INVX1 U1195 ( .A(n1373), .Y(n436) );
  INVX1 U1196 ( .A(\DP_OP_19_294_9081/n100 ), .Y(\DP_OP_19_294_9081/n98 ) );
  INVX1 U1197 ( .A(\DP_OP_19_294_9081/n202 ), .Y(\DP_OP_19_294_9081/n200 ) );
  INVX1 U1198 ( .A(\DP_OP_19_294_9081/n174 ), .Y(\DP_OP_19_294_9081/n172 ) );
  INVX1 U1199 ( .A(\DP_OP_19_294_9081/n106 ), .Y(\DP_OP_19_294_9081/n462 ) );
  INVX1 U1200 ( .A(\DP_OP_19_294_9081/n117 ), .Y(\DP_OP_19_294_9081/n463 ) );
  INVX1 U1201 ( .A(\DP_OP_19_294_9081/n120 ), .Y(\DP_OP_19_294_9081/n464 ) );
  INVX1 U1202 ( .A(\DP_OP_19_294_9081/n84 ), .Y(\DP_OP_19_294_9081/n82 ) );
  INVX1 U1203 ( .A(\DP_OP_19_294_9081/n87 ), .Y(\DP_OP_19_294_9081/n89 ) );
  INVX1 U1204 ( .A(\DP_OP_19_294_9081/n86 ), .Y(\DP_OP_19_294_9081/n88 ) );
  INVX1 U1205 ( .A(\DP_OP_19_294_9081/n103 ), .Y(\DP_OP_19_294_9081/n461 ) );
  INVX1 U1206 ( .A(\DP_OP_19_294_9081/n70 ), .Y(\DP_OP_19_294_9081/n458 ) );
  INVX1 U1207 ( .A(n1092), .Y(N91) );
  INVX1 U1208 ( .A(n1104), .Y(N102) );
  INVX1 U1209 ( .A(n1105), .Y(N103) );
  INVX1 U1210 ( .A(n1097), .Y(N96) );
  INVX1 U1211 ( .A(n1144), .Y(N87) );
  INVX1 U1212 ( .A(n1098), .Y(N97) );
  INVX1 U1213 ( .A(n1103), .Y(N101) );
  INVX1 U1214 ( .A(n1143), .Y(N86) );
  INVX1 U1215 ( .A(n1093), .Y(N92) );
  INVX1 U1216 ( .A(n1140), .Y(N85) );
  INVX1 U1217 ( .A(n1102), .Y(N100) );
  INVX1 U1218 ( .A(n1099), .Y(N98) );
  INVX1 U1219 ( .A(n1100), .Y(N99) );
  INVX1 U1220 ( .A(n1146), .Y(N89) );
  INVX1 U1221 ( .A(n1110), .Y(N108) );
  INVX1 U1222 ( .A(n1094), .Y(N93) );
  INVX1 U1223 ( .A(n1111), .Y(N109) );
  INVX1 U1224 ( .A(n1095), .Y(N94) );
  INVX1 U1225 ( .A(n1109), .Y(N107) );
  INVX1 U1226 ( .A(n1112), .Y(N110) );
  INVX1 U1227 ( .A(n1108), .Y(N106) );
  INVX1 U1228 ( .A(n1106), .Y(N104) );
  INVX1 U1229 ( .A(n1145), .Y(N88) );
  INVX1 U1230 ( .A(n1107), .Y(N105) );
  INVX1 U1231 ( .A(n1113), .Y(N111) );
  INVX1 U1232 ( .A(n1091), .Y(N90) );
  INVX1 U1233 ( .A(n1096), .Y(N95) );
  INVX1 U1234 ( .A(n1123), .Y(N123) );
  INVX1 U1235 ( .A(n1131), .Y(N131) );
  INVX1 U1236 ( .A(n1132), .Y(N132) );
  INVX1 U1237 ( .A(n1120), .Y(N119) );
  INVX1 U1238 ( .A(n1118), .Y(N117) );
  INVX1 U1239 ( .A(n1133), .Y(N133) );
  INVX1 U1240 ( .A(n1117), .Y(N116) );
  INVX1 U1241 ( .A(n1119), .Y(N118) );
  INVX1 U1242 ( .A(n1142), .Y(N141) );
  INVX1 U1243 ( .A(n1141), .Y(N140) );
  INVX1 U1244 ( .A(n1122), .Y(N122) );
  INVX1 U1245 ( .A(n1134), .Y(N134) );
  INVX1 U1246 ( .A(n1121), .Y(N120) );
  INVX1 U1247 ( .A(n1116), .Y(N115) );
  INVX1 U1248 ( .A(n1139), .Y(N139) );
  INVX1 U1249 ( .A(n1130), .Y(N130) );
  INVX1 U1250 ( .A(n1138), .Y(N138) );
  INVX1 U1251 ( .A(n1114), .Y(N113) );
  INVX1 U1252 ( .A(n1135), .Y(N135) );
  INVX1 U1253 ( .A(n1137), .Y(N137) );
  INVX1 U1254 ( .A(n1136), .Y(N136) );
  INVX1 U1255 ( .A(n1115), .Y(N114) );
  INVX1 U1256 ( .A(n1128), .Y(N128) );
  INVX1 U1257 ( .A(n1129), .Y(N129) );
  INVX1 U1258 ( .A(n1126), .Y(N126) );
  INVX1 U1259 ( .A(n1125), .Y(N125) );
  INVX1 U1260 ( .A(n1127), .Y(N127) );
  INVX1 U1261 ( .A(n1124), .Y(N124) );
  AND2X1 U1262 ( .A(\ashr_28_1/n643 ), .B(n1161), .Y(N143) );
  AND2X1 U1263 ( .A(n1173), .B(acc[14]), .Y(\C2/Z_14 ) );
  AND2X1 U1264 ( .A(n1173), .B(acc[39]), .Y(\C2/Z_39 ) );
  AND2X1 U1265 ( .A(n1173), .B(acc[59]), .Y(\C2/Z_59 ) );
  AND2X1 U1266 ( .A(n1173), .B(acc[27]), .Y(\C2/Z_27 ) );
  AND2X1 U1267 ( .A(n1173), .B(acc[9]), .Y(\C2/Z_9 ) );
  AND2X1 U1268 ( .A(n1173), .B(acc[26]), .Y(\C2/Z_26 ) );
  AND2X1 U1269 ( .A(n1173), .B(acc[28]), .Y(\C2/Z_28 ) );
  AND2X1 U1270 ( .A(n1173), .B(acc[7]), .Y(\C2/Z_7 ) );
  AND2X1 U1271 ( .A(n1173), .B(acc[16]), .Y(\C2/Z_16 ) );
  AND2X1 U1272 ( .A(n1173), .B(acc[24]), .Y(\C2/Z_24 ) );
  AND2X1 U1273 ( .A(n1173), .B(acc[48]), .Y(\C2/Z_48 ) );
  AND2X1 U1274 ( .A(n1173), .B(acc[61]), .Y(\C2/Z_61 ) );
  AND2X1 U1275 ( .A(n1173), .B(acc[62]), .Y(\C2/Z_62 ) );
  AND2X1 U1276 ( .A(n1173), .B(acc[13]), .Y(\C2/Z_13 ) );
  AND2X1 U1277 ( .A(n1173), .B(acc[60]), .Y(\C2/Z_60 ) );
  AND2X1 U1278 ( .A(n1173), .B(acc[49]), .Y(\C2/Z_49 ) );
  AND2X1 U1279 ( .A(n1173), .B(acc[40]), .Y(\C2/Z_40 ) );
  AND2X1 U1280 ( .A(n1173), .B(acc[6]), .Y(\C2/Z_6 ) );
  AND2X1 U1281 ( .A(n1173), .B(acc[42]), .Y(\C2/Z_42 ) );
  AND2X1 U1282 ( .A(n1173), .B(acc[29]), .Y(\C2/Z_29 ) );
  AND2X1 U1283 ( .A(n1173), .B(acc[46]), .Y(\C2/Z_46 ) );
  AND2X1 U1284 ( .A(n1173), .B(acc[25]), .Y(\C2/Z_25 ) );
  AND2X1 U1285 ( .A(n1173), .B(acc[56]), .Y(\C2/Z_56 ) );
  AND2X1 U1286 ( .A(n1173), .B(acc[32]), .Y(\C2/Z_32 ) );
  AND2X1 U1287 ( .A(n1173), .B(acc[52]), .Y(\C2/Z_52 ) );
  AND2X1 U1288 ( .A(n1173), .B(acc[22]), .Y(\C2/Z_22 ) );
  AND2X1 U1289 ( .A(n1173), .B(acc[51]), .Y(\C2/Z_51 ) );
  AND2X1 U1290 ( .A(n1173), .B(acc[11]), .Y(\C2/Z_11 ) );
  AND2X1 U1291 ( .A(n1173), .B(acc[34]), .Y(\C2/Z_34 ) );
  AND2X1 U1292 ( .A(n1173), .B(acc[36]), .Y(\C2/Z_36 ) );
  AND2X1 U1293 ( .A(n1173), .B(acc[55]), .Y(\C2/Z_55 ) );
  AND2X1 U1294 ( .A(n1173), .B(acc[57]), .Y(\C2/Z_57 ) );
  AND2X1 U1295 ( .A(n1173), .B(acc[31]), .Y(\C2/Z_31 ) );
  AND2X1 U1296 ( .A(n1173), .B(acc[23]), .Y(\C2/Z_23 ) );
  AND2X1 U1297 ( .A(n1173), .B(acc[50]), .Y(\C2/Z_50 ) );
  AND2X1 U1298 ( .A(n1173), .B(acc[53]), .Y(\C2/Z_53 ) );
  AND2X1 U1299 ( .A(n1173), .B(acc[58]), .Y(\C2/Z_58 ) );
  AND2X1 U1300 ( .A(n1173), .B(acc[47]), .Y(\C2/Z_47 ) );
  AND2X1 U1301 ( .A(n1173), .B(acc[10]), .Y(\C2/Z_10 ) );
  AND2X1 U1302 ( .A(n1173), .B(acc[30]), .Y(\C2/Z_30 ) );
  AND2X1 U1303 ( .A(n1173), .B(acc[12]), .Y(\C2/Z_12 ) );
  AND2X1 U1304 ( .A(n1173), .B(acc[54]), .Y(\C2/Z_54 ) );
  INVX2 U1305 ( .A(n1173), .Y(n1175) );
  AND2X1 U1306 ( .A(n1173), .B(acc[8]), .Y(\C2/Z_8 ) );
  INVX2 U1307 ( .A(n1065), .Y(n1167) );
  INVX2 U1308 ( .A(n1156), .Y(n1168) );
  INVX1 U1309 ( .A(mulout[29]), .Y(n1244) );
  INVX1 U1310 ( .A(mulout[58]), .Y(n1190) );
  INVX1 U1311 ( .A(mulout[9]), .Y(n1284) );
  INVX8 U1312 ( .A(n1154), .Y(n1067) );
  INVX1 U1313 ( .A(mulout[6]), .Y(n1290) );
  INVX1 U1314 ( .A(mulout[62]), .Y(n1184) );
  INVX1 U1315 ( .A(mulout[7]), .Y(n1288) );
  INVX1 U1316 ( .A(mulout[60]), .Y(n1186) );
  INVX1 U1317 ( .A(mulout[4]), .Y(n1294) );
  INVX1 U1318 ( .A(mulout[8]), .Y(n1286) );
  INVX1 U1319 ( .A(mulout[59]), .Y(n1188) );
  INVX2 U1320 ( .A(acc[2]), .Y(n1300) );
  INVX1 U1321 ( .A(mulout[5]), .Y(n1292) );
  INVX1 U1322 ( .A(mulout[39]), .Y(n1226) );
  INVX1 U1323 ( .A(mulout[48]), .Y(n1210) );
  INVX1 U1324 ( .A(mulout[49]), .Y(n1208) );
  INVX1 U1325 ( .A(mulout[16]), .Y(n1270) );
  INVX1 U1326 ( .A(mulout[0]), .Y(n1296) );
  INVX1 U1327 ( .A(mulout[23]), .Y(n1256) );
  INVX1 U1328 ( .A(mulout[50]), .Y(n1206) );
  INVX1 U1329 ( .A(mulout[15]), .Y(n1272) );
  INVX1 U1330 ( .A(mulout[51]), .Y(n1204) );
  INVX1 U1331 ( .A(mulout[38]), .Y(n1228) );
  INVX1 U1332 ( .A(mulout[52]), .Y(n1202) );
  INVX1 U1333 ( .A(mulout[24]), .Y(n1254) );
  INVX1 U1334 ( .A(mulout[41]), .Y(n1224) );
  INVX1 U1335 ( .A(mulout[42]), .Y(n1222) );
  INVX2 U1336 ( .A(acc[0]), .Y(n1303) );
  INVX1 U1337 ( .A(mulout[43]), .Y(n1220) );
  INVX1 U1338 ( .A(mulout[20]), .Y(n1262) );
  INVX1 U1339 ( .A(mulout[44]), .Y(n1218) );
  INVX1 U1340 ( .A(mulout[19]), .Y(n1264) );
  INVX1 U1341 ( .A(mulout[22]), .Y(n1258) );
  INVX1 U1342 ( .A(mulout[45]), .Y(n1216) );
  INVX1 U1343 ( .A(mulout[18]), .Y(n1266) );
  INVX1 U1344 ( .A(mulout[46]), .Y(n1214) );
  INVX1 U1345 ( .A(mulout[17]), .Y(n1268) );
  INVX1 U1346 ( .A(mulout[47]), .Y(n1212) );
  INVX1 U1347 ( .A(mulout[57]), .Y(n1192) );
  INVX1 U1348 ( .A(mulout[30]), .Y(n1242) );
  INVX1 U1349 ( .A(mulout[28]), .Y(n1246) );
  INVX1 U1350 ( .A(mulout[10]), .Y(n1282) );
  INVX1 U1351 ( .A(mulout[56]), .Y(n1194) );
  INVX1 U1352 ( .A(mulout[32]), .Y(n1240) );
  INVX1 U1353 ( .A(mulout[27]), .Y(n1248) );
  INVX1 U1354 ( .A(mulout[11]), .Y(n1280) );
  INVX1 U1355 ( .A(mulout[55]), .Y(n1196) );
  INVX1 U1356 ( .A(mulout[33]), .Y(n1238) );
  INVX1 U1357 ( .A(mulout[34]), .Y(n1236) );
  INVX1 U1358 ( .A(mulout[26]), .Y(n1250) );
  INVX1 U1359 ( .A(mulout[12]), .Y(n1278) );
  INVX1 U1360 ( .A(mulout[21]), .Y(n1260) );
  INVX1 U1361 ( .A(mulout[25]), .Y(n1252) );
  INVX1 U1362 ( .A(mulout[35]), .Y(n1234) );
  INVX2 U1363 ( .A(acc[1]), .Y(n1301) );
  INVX1 U1364 ( .A(mulout[54]), .Y(n1198) );
  INVX1 U1365 ( .A(mulout[13]), .Y(n1276) );
  INVX1 U1366 ( .A(mulout[53]), .Y(n1200) );
  INVX1 U1367 ( .A(mulout[36]), .Y(n1232) );
  INVX1 U1368 ( .A(mulout[37]), .Y(n1230) );
  BUFX2 U1369 ( .A(n283), .Y(n1068) );
  BUFX2 U1370 ( .A(n287), .Y(n1069) );
  BUFX2 U1371 ( .A(n291), .Y(n1070) );
  BUFX2 U1372 ( .A(n295), .Y(n1071) );
  BUFX2 U1373 ( .A(n299), .Y(n1072) );
  BUFX2 U1374 ( .A(n303), .Y(n1073) );
  BUFX2 U1375 ( .A(n307), .Y(n1074) );
  BUFX2 U1376 ( .A(n311), .Y(n1075) );
  BUFX2 U1377 ( .A(n315), .Y(n1076) );
  BUFX2 U1378 ( .A(n319), .Y(n1077) );
  BUFX2 U1379 ( .A(n323), .Y(n1078) );
  BUFX2 U1380 ( .A(n331), .Y(n1079) );
  BUFX2 U1381 ( .A(n335), .Y(n1080) );
  BUFX2 U1382 ( .A(n339), .Y(n1081) );
  BUFX2 U1383 ( .A(n343), .Y(n1082) );
  BUFX2 U1384 ( .A(n382), .Y(n1083) );
  BUFX2 U1385 ( .A(push_1), .Y(n1084) );
  BUFX2 U1386 ( .A(push_0), .Y(n1085) );
  BUFX2 U1387 ( .A(cmd0[0]), .Y(n1086) );
  BUFX2 U1388 ( .A(cmd0[1]), .Y(n1087) );
  INVX1 U1389 ( .A(n1064), .Y(\DP_OP_19_294_9081/n288 ) );
  INVX1 U1390 ( .A(\DP_OP_19_294_9081/n417 ), .Y(\DP_OP_19_294_9081/n511 ) );
  INVX1 U1391 ( .A(\DP_OP_19_294_9081/n405 ), .Y(\DP_OP_19_294_9081/n509 ) );
  INVX1 U1392 ( .A(\DP_OP_19_294_9081/n283 ), .Y(\DP_OP_19_294_9081/n487 ) );
  OR2X2 U1393 ( .A(\C2/Z_61 ), .B(\DP_OP_19_294_9081/n714 ), .Y(n1089) );
  INVX1 U1394 ( .A(\DP_OP_19_294_9081/n420 ), .Y(\DP_OP_19_294_9081/n512 ) );
  INVX1 U1395 ( .A(\DP_OP_19_294_9081/n206 ), .Y(\DP_OP_19_294_9081/n476 ) );
  INVX1 U1396 ( .A(\DP_OP_19_294_9081/n317 ), .Y(\DP_OP_19_294_9081/n315 ) );
  INVX1 U1397 ( .A(\DP_OP_19_294_9081/n428 ), .Y(\DP_OP_19_294_9081/n513 ) );
  INVX1 U1398 ( .A(\DP_OP_19_294_9081/n431 ), .Y(\DP_OP_19_294_9081/n514 ) );
  INVX1 U1399 ( .A(\DP_OP_19_294_9081/n247 ), .Y(\DP_OP_19_294_9081/n481 ) );
  INVX1 U1400 ( .A(\DP_OP_19_294_9081/n237 ), .Y(\DP_OP_19_294_9081/n239 ) );
  INVX1 U1401 ( .A(\DP_OP_19_294_9081/n238 ), .Y(\DP_OP_19_294_9081/n240 ) );
  INVX1 U1402 ( .A(\DP_OP_19_294_9081/n222 ), .Y(\DP_OP_19_294_9081/n478 ) );
  INVX1 U1403 ( .A(\DP_OP_19_294_9081/n4 ), .Y(\DP_OP_19_294_9081/n181 ) );
  INVX1 U1404 ( .A(\DP_OP_19_294_9081/n3 ), .Y(\DP_OP_19_294_9081/n182 ) );
  INVX1 U1405 ( .A(\DP_OP_19_294_9081/n178 ), .Y(\DP_OP_19_294_9081/n472 ) );
  INVX1 U1406 ( .A(\DP_OP_19_294_9081/n194 ), .Y(\DP_OP_19_294_9081/n474 ) );
  INVX1 U1407 ( .A(\DP_OP_19_294_9081/n155 ), .Y(\DP_OP_19_294_9081/n157 ) );
  INVX1 U1408 ( .A(\DP_OP_19_294_9081/n219 ), .Y(\DP_OP_19_294_9081/n477 ) );
  INVX1 U1409 ( .A(\DP_OP_19_294_9081/n231 ), .Y(\DP_OP_19_294_9081/n479 ) );
  INVX1 U1410 ( .A(\DP_OP_19_294_9081/n175 ), .Y(\DP_OP_19_294_9081/n471 ) );
  INVX1 U1411 ( .A(\DP_OP_19_294_9081/n250 ), .Y(\DP_OP_19_294_9081/n482 ) );
  INVX1 U1412 ( .A(\DP_OP_19_294_9081/n203 ), .Y(\DP_OP_19_294_9081/n475 ) );
  INVX1 U1413 ( .A(\DP_OP_19_294_9081/n166 ), .Y(\DP_OP_19_294_9081/n470 ) );
  INVX1 U1414 ( .A(\DP_OP_19_294_9081/n442 ), .Y(\DP_OP_19_294_9081/n440 ) );
  INVX1 U1415 ( .A(\DP_OP_19_294_9081/n267 ), .Y(\DP_OP_19_294_9081/n265 ) );
  INVX1 U1416 ( .A(\DP_OP_19_294_9081/n259 ), .Y(\DP_OP_19_294_9081/n483 ) );
  INVX1 U1417 ( .A(\DP_OP_19_294_9081/n275 ), .Y(\DP_OP_19_294_9081/n485 ) );
  INVX1 U1418 ( .A(\DP_OP_19_294_9081/n262 ), .Y(\DP_OP_19_294_9081/n484 ) );
  INVX1 U1419 ( .A(\DP_OP_19_294_9081/n278 ), .Y(\DP_OP_19_294_9081/n486 ) );
  INVX1 U1420 ( .A(\DP_OP_19_294_9081/n363 ), .Y(\DP_OP_19_294_9081/n501 ) );
  INVX1 U1421 ( .A(\DP_OP_19_294_9081/n286 ), .Y(\DP_OP_19_294_9081/n488 ) );
  INVX1 U1422 ( .A(\DP_OP_19_294_9081/n338 ), .Y(\DP_OP_19_294_9081/n336 ) );
  INVX1 U1423 ( .A(\DP_OP_19_294_9081/n339 ), .Y(\DP_OP_19_294_9081/n337 ) );
  INVX1 U1424 ( .A(\DP_OP_19_294_9081/n344 ), .Y(\DP_OP_19_294_9081/n497 ) );
  INVX1 U1425 ( .A(\DP_OP_19_294_9081/n366 ), .Y(\DP_OP_19_294_9081/n502 ) );
  INVX1 U1426 ( .A(\DP_OP_19_294_9081/n386 ), .Y(\DP_OP_19_294_9081/n505 ) );
  INVX1 U1427 ( .A(\DP_OP_19_294_9081/n376 ), .Y(\DP_OP_19_294_9081/n504 ) );
  INVX1 U1428 ( .A(\DP_OP_19_294_9081/n377 ), .Y(\DP_OP_19_294_9081/n375 ) );
  INVX1 U1429 ( .A(\DP_OP_19_294_9081/n371 ), .Y(\DP_OP_19_294_9081/n503 ) );
  INVX1 U1430 ( .A(\DP_OP_19_294_9081/n329 ), .Y(\DP_OP_19_294_9081/n495 ) );
  INVX1 U1431 ( .A(\DP_OP_19_294_9081/n352 ), .Y(\DP_OP_19_294_9081/n499 ) );
  INVX1 U1432 ( .A(\DP_OP_19_294_9081/n306 ), .Y(\DP_OP_19_294_9081/n491 ) );
  INVX1 U1433 ( .A(\DP_OP_19_294_9081/n394 ), .Y(\DP_OP_19_294_9081/n507 ) );
  INVX1 U1434 ( .A(\DP_OP_19_294_9081/n347 ), .Y(\DP_OP_19_294_9081/n498 ) );
  INVX1 U1435 ( .A(\DP_OP_19_294_9081/n324 ), .Y(\DP_OP_19_294_9081/n494 ) );
  INVX1 U1436 ( .A(\DP_OP_19_294_9081/n301 ), .Y(\DP_OP_19_294_9081/n490 ) );
  INVX1 U1437 ( .A(\DP_OP_19_294_9081/n389 ), .Y(\DP_OP_19_294_9081/n506 ) );
  INVX1 U1438 ( .A(\DP_OP_19_294_9081/n309 ), .Y(\DP_OP_19_294_9081/n492 ) );
  INVX1 U1439 ( .A(\DP_OP_19_294_9081/n355 ), .Y(\DP_OP_19_294_9081/n500 ) );
  INVX1 U1440 ( .A(\DP_OP_19_294_9081/n332 ), .Y(\DP_OP_19_294_9081/n496 ) );
  INVX1 U1441 ( .A(\DP_OP_19_294_9081/n397 ), .Y(\DP_OP_19_294_9081/n508 ) );
  INVX2 U1442 ( .A(\DP_OP_19_294_9081/n99 ), .Y(\DP_OP_19_294_9081/n97 ) );
  INVX2 U1443 ( .A(\DP_OP_19_294_9081/n335 ), .Y(\DP_OP_19_294_9081/n334 ) );
  INVX2 U1444 ( .A(\DP_OP_19_294_9081/n358 ), .Y(\DP_OP_19_294_9081/n357 ) );
  INVX2 U1445 ( .A(\DP_OP_19_294_9081/n312 ), .Y(\DP_OP_19_294_9081/n311 ) );
  INVX2 U1446 ( .A(\DP_OP_19_294_9081/n400 ), .Y(\DP_OP_19_294_9081/n399 ) );
  INVX1 U1447 ( .A(\DP_OP_19_294_9081/n450 ), .Y(\DP_OP_19_294_9081/n518 ) );
  INVX1 U1448 ( .A(\DP_OP_19_294_9081/n447 ), .Y(\DP_OP_19_294_9081/n517 ) );
  INVX1 U1449 ( .A(\DP_OP_19_294_9081/n415 ), .Y(\DP_OP_19_294_9081/n413 ) );
  INVX1 U1450 ( .A(\DP_OP_19_294_9081/n416 ), .Y(\DP_OP_19_294_9081/n414 ) );
  INVX1 U1451 ( .A(\DP_OP_19_294_9081/n410 ), .Y(\DP_OP_19_294_9081/n510 ) );
  INVX1 U1452 ( .A(\DP_OP_19_294_9081/n411 ), .Y(\DP_OP_19_294_9081/n409 ) );
  INVX1 U1453 ( .A(\DP_OP_19_294_9081/n163 ), .Y(\DP_OP_19_294_9081/n469 ) );
  INVX1 U1454 ( .A(\DP_OP_19_294_9081/n215 ), .Y(\DP_OP_19_294_9081/n213 ) );
  INVX1 U1455 ( .A(\DP_OP_19_294_9081/n298 ), .Y(\DP_OP_19_294_9081/n489 ) );
  INVX1 U1456 ( .A(\DP_OP_19_294_9081/n257 ), .Y(\DP_OP_19_294_9081/n255 ) );
  INVX1 U1457 ( .A(\DP_OP_19_294_9081/n229 ), .Y(\DP_OP_19_294_9081/n227 ) );
  INVX1 U1458 ( .A(\DP_OP_19_294_9081/n436 ), .Y(\DP_OP_19_294_9081/n515 ) );
  INVX1 U1459 ( .A(\DP_OP_19_294_9081/n268 ), .Y(\DP_OP_19_294_9081/n266 ) );
  INVX1 U1460 ( .A(\DP_OP_19_294_9081/n1 ), .Y(\DP_OP_19_294_9081/n378 ) );
  INVX1 U1461 ( .A(\DP_OP_19_294_9081/n321 ), .Y(\DP_OP_19_294_9081/n493 ) );
  INVX1 U1462 ( .A(\DP_OP_19_294_9081/n454 ), .Y(\DP_OP_19_294_9081/n519 ) );
  INVX1 U1463 ( .A(\DP_OP_19_294_9081/n453 ), .Y(\DP_OP_19_294_9081/n452 ) );
  INVX1 U1464 ( .A(\DP_OP_19_294_9081/n173 ), .Y(\DP_OP_19_294_9081/n171 ) );
  INVX1 U1465 ( .A(\DP_OP_19_294_9081/n211 ), .Y(\DP_OP_19_294_9081/n209 ) );
  INVX1 U1466 ( .A(\DP_OP_19_294_9081/n318 ), .Y(\DP_OP_19_294_9081/n316 ) );
  INVX1 U1467 ( .A(\DP_OP_19_294_9081/n127 ), .Y(\DP_OP_19_294_9081/n125 ) );
  INVX1 U1468 ( .A(\DP_OP_19_294_9081/n201 ), .Y(\DP_OP_19_294_9081/n199 ) );
  INVX1 U1469 ( .A(\DP_OP_19_294_9081/n191 ), .Y(\DP_OP_19_294_9081/n473 ) );
  INVX1 U1470 ( .A(\DP_OP_19_294_9081/n147 ), .Y(\DP_OP_19_294_9081/n467 ) );
  INVX1 U1471 ( .A(\DP_OP_19_294_9081/n216 ), .Y(\DP_OP_19_294_9081/n214 ) );
  INVX1 U1472 ( .A(\DP_OP_19_294_9081/n212 ), .Y(\DP_OP_19_294_9081/n210 ) );
  INVX1 U1473 ( .A(\DP_OP_19_294_9081/n444 ), .Y(\DP_OP_19_294_9081/n443 ) );
  INVX1 U1474 ( .A(\DP_OP_19_294_9081/n128 ), .Y(\DP_OP_19_294_9081/n126 ) );
  INVX1 U1475 ( .A(\DP_OP_19_294_9081/n441 ), .Y(\DP_OP_19_294_9081/n516 ) );
  INVX1 U1476 ( .A(\DP_OP_19_294_9081/n423 ), .Y(\DP_OP_19_294_9081/n422 ) );
  INVX1 U1477 ( .A(\DP_OP_19_294_9081/n258 ), .Y(\DP_OP_19_294_9081/n256 ) );
  INVX1 U1478 ( .A(\DP_OP_19_294_9081/n230 ), .Y(\DP_OP_19_294_9081/n228 ) );
  INVX1 U1479 ( .A(\DP_OP_19_294_9081/n150 ), .Y(\DP_OP_19_294_9081/n468 ) );
  INVX1 U1480 ( .A(\DP_OP_19_294_9081/n156 ), .Y(\DP_OP_19_294_9081/n158 ) );
  INVX1 U1481 ( .A(\DP_OP_19_294_9081/n133 ), .Y(\DP_OP_19_294_9081/n465 ) );
  INVX1 U1482 ( .A(\DP_OP_19_294_9081/n136 ), .Y(\DP_OP_19_294_9081/n466 ) );
  MUX2X1 U1483 ( .B(\ashr_28_1/n582 ), .A(\ashr_28_1/n580 ), .S(n1161), .Y(
        n1090) );
  MUX2X1 U1484 ( .B(\ashr_28_1/n590 ), .A(\ashr_28_1/n592 ), .S(h2[1]), .Y(
        n1091) );
  MUX2X1 U1485 ( .B(\ashr_28_1/n591 ), .A(\ashr_28_1/n593 ), .S(h2[1]), .Y(
        n1092) );
  MUX2X1 U1486 ( .B(\ashr_28_1/n592 ), .A(\ashr_28_1/n594 ), .S(h2[1]), .Y(
        n1093) );
  MUX2X1 U1487 ( .B(\ashr_28_1/n593 ), .A(\ashr_28_1/n595 ), .S(h2[1]), .Y(
        n1094) );
  MUX2X1 U1488 ( .B(\ashr_28_1/n594 ), .A(\ashr_28_1/n596 ), .S(h2[1]), .Y(
        n1095) );
  MUX2X1 U1489 ( .B(\ashr_28_1/n595 ), .A(\ashr_28_1/n597 ), .S(h2[1]), .Y(
        n1096) );
  MUX2X1 U1490 ( .B(\ashr_28_1/n596 ), .A(\ashr_28_1/n598 ), .S(h2[1]), .Y(
        n1097) );
  MUX2X1 U1491 ( .B(\ashr_28_1/n597 ), .A(\ashr_28_1/n599 ), .S(h2[1]), .Y(
        n1098) );
  MUX2X1 U1492 ( .B(\ashr_28_1/n598 ), .A(\ashr_28_1/n600 ), .S(h2[1]), .Y(
        n1099) );
  MUX2X1 U1493 ( .B(\ashr_28_1/n599 ), .A(\ashr_28_1/n601 ), .S(n1162), .Y(
        n1100) );
  MUX2X1 U1494 ( .B(\ashr_28_1/n583 ), .A(\ashr_28_1/n581 ), .S(n1161), .Y(
        n1101) );
  MUX2X1 U1495 ( .B(\ashr_28_1/n600 ), .A(\ashr_28_1/n602 ), .S(n1162), .Y(
        n1102) );
  MUX2X1 U1496 ( .B(\ashr_28_1/n601 ), .A(\ashr_28_1/n603 ), .S(n1162), .Y(
        n1103) );
  MUX2X1 U1497 ( .B(\ashr_28_1/n602 ), .A(\ashr_28_1/n604 ), .S(n1162), .Y(
        n1104) );
  MUX2X1 U1498 ( .B(\ashr_28_1/n603 ), .A(\ashr_28_1/n605 ), .S(n1162), .Y(
        n1105) );
  MUX2X1 U1499 ( .B(\ashr_28_1/n604 ), .A(\ashr_28_1/n606 ), .S(n1162), .Y(
        n1106) );
  MUX2X1 U1500 ( .B(\ashr_28_1/n605 ), .A(\ashr_28_1/n607 ), .S(n1162), .Y(
        n1107) );
  MUX2X1 U1501 ( .B(\ashr_28_1/n606 ), .A(\ashr_28_1/n608 ), .S(n1162), .Y(
        n1108) );
  MUX2X1 U1502 ( .B(\ashr_28_1/n607 ), .A(\ashr_28_1/n609 ), .S(n1162), .Y(
        n1109) );
  MUX2X1 U1503 ( .B(\ashr_28_1/n608 ), .A(\ashr_28_1/n610 ), .S(n1162), .Y(
        n1110) );
  MUX2X1 U1504 ( .B(\ashr_28_1/n609 ), .A(\ashr_28_1/n611 ), .S(n1162), .Y(
        n1111) );
  MUX2X1 U1505 ( .B(\ashr_28_1/n610 ), .A(\ashr_28_1/n612 ), .S(n1163), .Y(
        n1112) );
  MUX2X1 U1506 ( .B(\ashr_28_1/n611 ), .A(\ashr_28_1/n613 ), .S(n1163), .Y(
        n1113) );
  MUX2X1 U1507 ( .B(\ashr_28_1/n615 ), .A(\ashr_28_1/n613 ), .S(n1161), .Y(
        n1114) );
  MUX2X1 U1508 ( .B(\ashr_28_1/n616 ), .A(\ashr_28_1/n614 ), .S(n1161), .Y(
        n1115) );
  MUX2X1 U1509 ( .B(\ashr_28_1/n615 ), .A(\ashr_28_1/n617 ), .S(n1163), .Y(
        n1116) );
  MUX2X1 U1510 ( .B(\ashr_28_1/n616 ), .A(\ashr_28_1/n618 ), .S(n1163), .Y(
        n1117) );
  MUX2X1 U1511 ( .B(\ashr_28_1/n619 ), .A(\ashr_28_1/n617 ), .S(n1161), .Y(
        n1118) );
  MUX2X1 U1512 ( .B(\ashr_28_1/n620 ), .A(\ashr_28_1/n618 ), .S(n1161), .Y(
        n1119) );
  MUX2X1 U1513 ( .B(\ashr_28_1/n619 ), .A(\ashr_28_1/n621 ), .S(n1163), .Y(
        n1120) );
  MUX2X1 U1514 ( .B(\ashr_28_1/n620 ), .A(\ashr_28_1/n622 ), .S(n1163), .Y(
        n1121) );
  MUX2X1 U1515 ( .B(\ashr_28_1/n624 ), .A(\ashr_28_1/n622 ), .S(n1161), .Y(
        n1122) );
  MUX2X1 U1516 ( .B(\ashr_28_1/n623 ), .A(\ashr_28_1/n625 ), .S(n1163), .Y(
        n1123) );
  MUX2X1 U1517 ( .B(\ashr_28_1/n624 ), .A(\ashr_28_1/n626 ), .S(n1163), .Y(
        n1124) );
  MUX2X1 U1518 ( .B(\ashr_28_1/n627 ), .A(\ashr_28_1/n625 ), .S(n1161), .Y(
        n1125) );
  MUX2X1 U1519 ( .B(\ashr_28_1/n628 ), .A(\ashr_28_1/n626 ), .S(n1161), .Y(
        n1126) );
  MUX2X1 U1520 ( .B(\ashr_28_1/n627 ), .A(\ashr_28_1/n629 ), .S(n1163), .Y(
        n1127) );
  MUX2X1 U1521 ( .B(\ashr_28_1/n628 ), .A(\ashr_28_1/n630 ), .S(n1163), .Y(
        n1128) );
  MUX2X1 U1522 ( .B(\ashr_28_1/n631 ), .A(\ashr_28_1/n629 ), .S(n1161), .Y(
        n1129) );
  MUX2X1 U1523 ( .B(\ashr_28_1/n632 ), .A(\ashr_28_1/n630 ), .S(n1161), .Y(
        n1130) );
  MUX2X1 U1524 ( .B(\ashr_28_1/n631 ), .A(\ashr_28_1/n633 ), .S(n1164), .Y(
        n1131) );
  MUX2X1 U1525 ( .B(\ashr_28_1/n632 ), .A(\ashr_28_1/n634 ), .S(n1164), .Y(
        n1132) );
  MUX2X1 U1526 ( .B(\ashr_28_1/n635 ), .A(\ashr_28_1/n633 ), .S(n1161), .Y(
        n1133) );
  MUX2X1 U1527 ( .B(\ashr_28_1/n636 ), .A(\ashr_28_1/n634 ), .S(n1161), .Y(
        n1134) );
  MUX2X1 U1528 ( .B(\ashr_28_1/n635 ), .A(\ashr_28_1/n637 ), .S(n1164), .Y(
        n1135) );
  MUX2X1 U1529 ( .B(\ashr_28_1/n636 ), .A(\ashr_28_1/n638 ), .S(n1164), .Y(
        n1136) );
  MUX2X1 U1530 ( .B(\ashr_28_1/n639 ), .A(\ashr_28_1/n637 ), .S(n1161), .Y(
        n1137) );
  MUX2X1 U1531 ( .B(\ashr_28_1/n640 ), .A(\ashr_28_1/n638 ), .S(n1161), .Y(
        n1138) );
  MUX2X1 U1532 ( .B(\ashr_28_1/n639 ), .A(\ashr_28_1/n641 ), .S(n1164), .Y(
        n1139) );
  MUX2X1 U1533 ( .B(\ashr_28_1/n585 ), .A(\ashr_28_1/n587 ), .S(n1164), .Y(
        n1140) );
  MUX2X1 U1534 ( .B(\ashr_28_1/n640 ), .A(\ashr_28_1/n642 ), .S(n1164), .Y(
        n1141) );
  MUX2X1 U1535 ( .B(\ashr_28_1/n643 ), .A(\ashr_28_1/n641 ), .S(n1161), .Y(
        n1142) );
  MUX2X1 U1536 ( .B(\ashr_28_1/n586 ), .A(\ashr_28_1/n588 ), .S(n1164), .Y(
        n1143) );
  MUX2X1 U1537 ( .B(\ashr_28_1/n587 ), .A(\ashr_28_1/n589 ), .S(n1164), .Y(
        n1144) );
  MUX2X1 U1538 ( .B(\ashr_28_1/n588 ), .A(\ashr_28_1/n590 ), .S(n1164), .Y(
        n1145) );
  MUX2X1 U1539 ( .B(\ashr_28_1/n589 ), .A(\ashr_28_1/n591 ), .S(n1164), .Y(
        n1146) );
  NAND2X1 U1540 ( .A(n1157), .B(\ashr_28_1/n771 ), .Y(\ashr_28_1/n706 ) );
  NAND2X1 U1541 ( .A(n1157), .B(\ashr_28_1/n772 ), .Y(\ashr_28_1/n707 ) );
  NAND2X1 U1542 ( .A(n1157), .B(\ashr_28_1/n773 ), .Y(\ashr_28_1/n708 ) );
  NAND2X1 U1543 ( .A(n1157), .B(\ashr_28_1/n774 ), .Y(\ashr_28_1/n709 ) );
  NAND2X1 U1544 ( .A(n1154), .B(\ashr_28_1/n889 ), .Y(\ashr_28_1/n824 ) );
  NAND2X1 U1545 ( .A(n1154), .B(\ashr_28_1/n890 ), .Y(\ashr_28_1/n825 ) );
  NAND2X1 U1546 ( .A(n1154), .B(\ashr_28_1/n891 ), .Y(\ashr_28_1/n826 ) );
  NAND2X1 U1547 ( .A(n1154), .B(\ashr_28_1/n892 ), .Y(\ashr_28_1/n827 ) );
  NAND2X1 U1548 ( .A(n1154), .B(\ashr_28_1/n893 ), .Y(\ashr_28_1/n828 ) );
  NAND2X1 U1549 ( .A(n1154), .B(\ashr_28_1/n894 ), .Y(\ashr_28_1/n829 ) );
  NAND2X1 U1550 ( .A(n1154), .B(\ashr_28_1/n895 ), .Y(\ashr_28_1/n830 ) );
  NAND2X1 U1551 ( .A(n1154), .B(\ashr_28_1/n896 ), .Y(\ashr_28_1/n831 ) );
  NAND2X1 U1552 ( .A(n1154), .B(\ashr_28_1/n897 ), .Y(\ashr_28_1/n832 ) );
  NAND2X1 U1553 ( .A(n1154), .B(\ashr_28_1/n898 ), .Y(\ashr_28_1/n833 ) );
  NAND2X1 U1554 ( .A(n1154), .B(\ashr_28_1/n899 ), .Y(\ashr_28_1/n834 ) );
  NAND2X1 U1555 ( .A(n1154), .B(\ashr_28_1/n900 ), .Y(\ashr_28_1/n835 ) );
  NAND2X1 U1556 ( .A(n1154), .B(\ashr_28_1/n901 ), .Y(\ashr_28_1/n836 ) );
  NAND2X1 U1557 ( .A(n1154), .B(\ashr_28_1/n902 ), .Y(\ashr_28_1/n837 ) );
  NAND2X1 U1558 ( .A(n1154), .B(\ashr_28_1/n903 ), .Y(\ashr_28_1/n838 ) );
  NAND2X1 U1559 ( .A(n1154), .B(\ashr_28_1/n904 ), .Y(\ashr_28_1/n839 ) );
  NAND2X1 U1560 ( .A(n1150), .B(acc[32]), .Y(\ashr_28_1/n938 ) );
  NAND2X1 U1561 ( .A(n1150), .B(acc[33]), .Y(\ashr_28_1/n939 ) );
  NAND2X1 U1562 ( .A(n1150), .B(acc[34]), .Y(\ashr_28_1/n940 ) );
  NAND2X1 U1563 ( .A(n1150), .B(acc[35]), .Y(\ashr_28_1/n941 ) );
  NAND2X1 U1564 ( .A(n1150), .B(acc[36]), .Y(\ashr_28_1/n942 ) );
  NAND2X1 U1565 ( .A(n1150), .B(acc[37]), .Y(\ashr_28_1/n943 ) );
  NAND2X1 U1566 ( .A(n1150), .B(acc[38]), .Y(\ashr_28_1/n944 ) );
  NAND2X1 U1567 ( .A(n1150), .B(acc[39]), .Y(\ashr_28_1/n945 ) );
  NAND2X1 U1568 ( .A(n1150), .B(acc[40]), .Y(\ashr_28_1/n946 ) );
  NAND2X1 U1569 ( .A(n1150), .B(acc[41]), .Y(\ashr_28_1/n947 ) );
  NAND2X1 U1570 ( .A(n1150), .B(acc[42]), .Y(\ashr_28_1/n948 ) );
  NAND2X1 U1571 ( .A(n1150), .B(acc[43]), .Y(\ashr_28_1/n949 ) );
  NAND2X1 U1572 ( .A(n1150), .B(acc[44]), .Y(\ashr_28_1/n950 ) );
  NAND2X1 U1573 ( .A(n1150), .B(acc[45]), .Y(\ashr_28_1/n951 ) );
  NAND2X1 U1574 ( .A(n1150), .B(acc[46]), .Y(\ashr_28_1/n952 ) );
  NAND2X1 U1575 ( .A(n1150), .B(acc[47]), .Y(\ashr_28_1/n953 ) );
  NAND2X1 U1576 ( .A(n1150), .B(acc[48]), .Y(\ashr_28_1/n954 ) );
  NAND2X1 U1577 ( .A(n1150), .B(acc[49]), .Y(\ashr_28_1/n955 ) );
  NAND2X1 U1578 ( .A(n1150), .B(acc[50]), .Y(\ashr_28_1/n956 ) );
  NAND2X1 U1579 ( .A(n1151), .B(acc[51]), .Y(\ashr_28_1/n957 ) );
  NAND2X1 U1580 ( .A(n1150), .B(acc[52]), .Y(\ashr_28_1/n958 ) );
  NAND2X1 U1581 ( .A(n1150), .B(acc[53]), .Y(\ashr_28_1/n959 ) );
  NAND2X1 U1582 ( .A(n1150), .B(acc[54]), .Y(\ashr_28_1/n960 ) );
  NAND2X1 U1583 ( .A(n1150), .B(acc[55]), .Y(\ashr_28_1/n961 ) );
  NAND2X1 U1584 ( .A(n1150), .B(acc[56]), .Y(\ashr_28_1/n962 ) );
  NAND2X1 U1585 ( .A(n1150), .B(acc[57]), .Y(\ashr_28_1/n963 ) );
  NAND2X1 U1586 ( .A(n1150), .B(acc[58]), .Y(\ashr_28_1/n964 ) );
  NAND2X1 U1587 ( .A(n1150), .B(acc[59]), .Y(\ashr_28_1/n965 ) );
  NAND2X1 U1588 ( .A(n1150), .B(acc[60]), .Y(\ashr_28_1/n966 ) );
  NAND2X1 U1589 ( .A(n1150), .B(acc[61]), .Y(\ashr_28_1/n967 ) );
  NAND2X1 U1590 ( .A(n1150), .B(acc[62]), .Y(\ashr_28_1/n968 ) );
  NAND2X1 U1591 ( .A(acc[63]), .B(n1150), .Y(\ashr_28_1/n969 ) );
  MUX2X1 U1592 ( .B(\ashr_28_1/n864 ), .A(\ashr_28_1/n848 ), .S(n1154), .Y(
        \ashr_28_1/n783 ) );
  INVX2 U1593 ( .A(n1157), .Y(n1158) );
  INVX2 U1594 ( .A(n1161), .Y(n1162) );
  INVX2 U1595 ( .A(n1161), .Y(n1163) );
  INVX2 U1596 ( .A(n1161), .Y(n1164) );
  BUFX4 U1597 ( .A(h2[3]), .Y(n1155) );
  INVX8 U1598 ( .A(n1147), .Y(n1149) );
  INVX4 U1599 ( .A(n1147), .Y(n1148) );
  INVX4 U1600 ( .A(\ashr_28_1/SH[5] ), .Y(n1150) );
  BUFX2 U1601 ( .A(h2[3]), .Y(n1156) );
  INVX8 U1602 ( .A(n1151), .Y(n1153) );
  INVX2 U1603 ( .A(h2[2]), .Y(n1157) );
  INVX2 U1604 ( .A(n1157), .Y(n1160) );
  INVX2 U1605 ( .A(n1157), .Y(n1159) );
  INVX8 U1606 ( .A(n1151), .Y(n1152) );
  BUFX4 U1607 ( .A(h2[0]), .Y(n1166) );
  MUX2X1 U1608 ( .B(\ashr_28_1/n871 ), .A(\ashr_28_1/n855 ), .S(n1167), .Y(
        \ashr_28_1/n790 ) );
  INVX1 U1609 ( .A(n1101), .Y(N81) );
  MUX2X1 U1610 ( .B(\ashr_28_1/n790 ), .A(\ashr_28_1/n782 ), .S(n1168), .Y(
        \ashr_28_1/n717 ) );
  INVX4 U1611 ( .A(h2[5]), .Y(n1182) );
  INVX8 U1612 ( .A(push_2), .Y(n1179) );
  INVX2 U1613 ( .A(n1378), .Y(n1180) );
  INVX2 U1614 ( .A(n1374), .Y(n1177) );
  INVX8 U1615 ( .A(n1182), .Y(\ashr_28_1/SH[5] ) );
  INVX4 U1616 ( .A(n1172), .Y(n1176) );
  INVX1 U1617 ( .A(n629), .Y(n1376) );
  BUFX2 U1618 ( .A(n630), .Y(n1181) );
  INVX1 U1619 ( .A(acc[4]), .Y(n1298) );
  INVX1 U1620 ( .A(acc[5]), .Y(n1297) );
  INVX1 U1621 ( .A(n445), .Y(n1377) );
  INVX8 U1622 ( .A(n1305), .Y(n1173) );
  NAND2X1 U1623 ( .A(n629), .B(n1377), .Y(n1304) );
  NAND2X1 U1624 ( .A(n445), .B(n1376), .Y(n1305) );
  NAND2X1 U1625 ( .A(n1302), .B(N143), .Y(n1183) );
  OAI21X1 U1626 ( .A(n1184), .B(n1174), .C(n1183), .Y(\DP_OP_19_294_9081/n715 ) );
  NAND2X1 U1627 ( .A(n1302), .B(N141), .Y(n1185) );
  OAI21X1 U1628 ( .A(n1186), .B(n1174), .C(n1185), .Y(\DP_OP_19_294_9081/n713 ) );
  NAND2X1 U1629 ( .A(n1302), .B(N140), .Y(n1187) );
  OAI21X1 U1630 ( .A(n1188), .B(n1174), .C(n1187), .Y(\DP_OP_19_294_9081/n712 ) );
  NAND2X1 U1631 ( .A(n1302), .B(N139), .Y(n1189) );
  OAI21X1 U1632 ( .A(n1190), .B(n1174), .C(n1189), .Y(\DP_OP_19_294_9081/n711 ) );
  NAND2X1 U1633 ( .A(n1302), .B(N138), .Y(n1191) );
  OAI21X1 U1634 ( .A(n1192), .B(n1174), .C(n1191), .Y(\DP_OP_19_294_9081/n710 ) );
  NAND2X1 U1635 ( .A(n1302), .B(N137), .Y(n1193) );
  OAI21X1 U1636 ( .A(n1194), .B(n1174), .C(n1193), .Y(\DP_OP_19_294_9081/n709 ) );
  NAND2X1 U1637 ( .A(n1302), .B(N136), .Y(n1195) );
  OAI21X1 U1638 ( .A(n1196), .B(n1174), .C(n1195), .Y(\DP_OP_19_294_9081/n708 ) );
  NAND2X1 U1639 ( .A(n1302), .B(N135), .Y(n1197) );
  OAI21X1 U1640 ( .A(n1198), .B(n1174), .C(n1197), .Y(\DP_OP_19_294_9081/n707 ) );
  NAND2X1 U1641 ( .A(n1302), .B(N134), .Y(n1199) );
  OAI21X1 U1642 ( .A(n1200), .B(n1174), .C(n1199), .Y(\DP_OP_19_294_9081/n706 ) );
  NAND2X1 U1643 ( .A(n1302), .B(N133), .Y(n1201) );
  OAI21X1 U1644 ( .A(n1202), .B(n1174), .C(n1201), .Y(\DP_OP_19_294_9081/n705 ) );
  NAND2X1 U1645 ( .A(n1302), .B(N132), .Y(n1203) );
  OAI21X1 U1646 ( .A(n1204), .B(n1174), .C(n1203), .Y(\DP_OP_19_294_9081/n704 ) );
  NAND2X1 U1647 ( .A(n1302), .B(N131), .Y(n1205) );
  OAI21X1 U1648 ( .A(n1206), .B(n1174), .C(n1205), .Y(\DP_OP_19_294_9081/n703 ) );
  NAND2X1 U1649 ( .A(n1302), .B(N130), .Y(n1207) );
  OAI21X1 U1650 ( .A(n1208), .B(n1174), .C(n1207), .Y(\DP_OP_19_294_9081/n702 ) );
  NAND2X1 U1651 ( .A(n1302), .B(N129), .Y(n1209) );
  OAI21X1 U1652 ( .A(n1210), .B(n1174), .C(n1209), .Y(\DP_OP_19_294_9081/n701 ) );
  NAND2X1 U1653 ( .A(n1302), .B(N128), .Y(n1211) );
  OAI21X1 U1654 ( .A(n1212), .B(n1174), .C(n1211), .Y(\DP_OP_19_294_9081/n700 ) );
  NAND2X1 U1655 ( .A(n1302), .B(N127), .Y(n1213) );
  OAI21X1 U1656 ( .A(n1214), .B(n1174), .C(n1213), .Y(\DP_OP_19_294_9081/n699 ) );
  NAND2X1 U1657 ( .A(n1302), .B(N126), .Y(n1215) );
  OAI21X1 U1658 ( .A(n1216), .B(n1174), .C(n1215), .Y(\DP_OP_19_294_9081/n698 ) );
  NAND2X1 U1659 ( .A(n1302), .B(N125), .Y(n1217) );
  OAI21X1 U1660 ( .A(n1218), .B(n1174), .C(n1217), .Y(\DP_OP_19_294_9081/n697 ) );
  NAND2X1 U1661 ( .A(n1302), .B(N124), .Y(n1219) );
  OAI21X1 U1662 ( .A(n1220), .B(n1174), .C(n1219), .Y(\DP_OP_19_294_9081/n696 ) );
  NAND2X1 U1663 ( .A(n1302), .B(N123), .Y(n1221) );
  OAI21X1 U1664 ( .A(n1222), .B(n1174), .C(n1221), .Y(\DP_OP_19_294_9081/n695 ) );
  NAND2X1 U1665 ( .A(n1302), .B(N122), .Y(n1223) );
  OAI21X1 U1666 ( .A(n1224), .B(n1174), .C(n1223), .Y(\DP_OP_19_294_9081/n694 ) );
  NAND2X1 U1667 ( .A(n1302), .B(N120), .Y(n1225) );
  OAI21X1 U1668 ( .A(n1226), .B(n1174), .C(n1225), .Y(\DP_OP_19_294_9081/n692 ) );
  NAND2X1 U1669 ( .A(n1302), .B(N119), .Y(n1227) );
  OAI21X1 U1670 ( .A(n1228), .B(n1066), .C(n1227), .Y(\DP_OP_19_294_9081/n691 ) );
  NAND2X1 U1671 ( .A(n1302), .B(N118), .Y(n1229) );
  OAI21X1 U1672 ( .A(n1230), .B(n1066), .C(n1229), .Y(\DP_OP_19_294_9081/n690 ) );
  NAND2X1 U1673 ( .A(n1302), .B(N117), .Y(n1231) );
  OAI21X1 U1674 ( .A(n1232), .B(n1066), .C(n1231), .Y(\DP_OP_19_294_9081/n689 ) );
  NAND2X1 U1675 ( .A(n1302), .B(N116), .Y(n1233) );
  OAI21X1 U1676 ( .A(n1234), .B(n1066), .C(n1233), .Y(\DP_OP_19_294_9081/n688 ) );
  NAND2X1 U1677 ( .A(n1302), .B(N115), .Y(n1235) );
  OAI21X1 U1678 ( .A(n1236), .B(n1066), .C(n1235), .Y(\DP_OP_19_294_9081/n687 ) );
  NAND2X1 U1679 ( .A(n1302), .B(N114), .Y(n1237) );
  OAI21X1 U1680 ( .A(n1238), .B(n1066), .C(n1237), .Y(\DP_OP_19_294_9081/n686 ) );
  NAND2X1 U1681 ( .A(n1302), .B(N113), .Y(n1239) );
  OAI21X1 U1682 ( .A(n1240), .B(n1066), .C(n1239), .Y(\DP_OP_19_294_9081/n685 ) );
  NAND2X1 U1683 ( .A(n1302), .B(N111), .Y(n1241) );
  OAI21X1 U1684 ( .A(n1242), .B(n1066), .C(n1241), .Y(\DP_OP_19_294_9081/n683 ) );
  NAND2X1 U1685 ( .A(n1302), .B(N110), .Y(n1243) );
  OAI21X1 U1686 ( .A(n1244), .B(n1066), .C(n1243), .Y(\DP_OP_19_294_9081/n682 ) );
  NAND2X1 U1687 ( .A(n1302), .B(N109), .Y(n1245) );
  OAI21X1 U1688 ( .A(n1246), .B(n1066), .C(n1245), .Y(\DP_OP_19_294_9081/n681 ) );
  NAND2X1 U1689 ( .A(n1302), .B(N108), .Y(n1247) );
  OAI21X1 U1690 ( .A(n1248), .B(n1066), .C(n1247), .Y(\DP_OP_19_294_9081/n680 ) );
  NAND2X1 U1691 ( .A(n1302), .B(N107), .Y(n1249) );
  OAI21X1 U1692 ( .A(n1250), .B(n1174), .C(n1249), .Y(\DP_OP_19_294_9081/n679 ) );
  NAND2X1 U1693 ( .A(n1302), .B(N106), .Y(n1251) );
  OAI21X1 U1694 ( .A(n1252), .B(n1174), .C(n1251), .Y(\DP_OP_19_294_9081/n678 ) );
  NAND2X1 U1695 ( .A(n1302), .B(N105), .Y(n1253) );
  OAI21X1 U1696 ( .A(n1254), .B(n1174), .C(n1253), .Y(\DP_OP_19_294_9081/n677 ) );
  NAND2X1 U1697 ( .A(n1302), .B(N104), .Y(n1255) );
  OAI21X1 U1698 ( .A(n1256), .B(n1174), .C(n1255), .Y(\DP_OP_19_294_9081/n676 ) );
  NAND2X1 U1699 ( .A(n1302), .B(N103), .Y(n1257) );
  OAI21X1 U1700 ( .A(n1258), .B(n1174), .C(n1257), .Y(\DP_OP_19_294_9081/n675 ) );
  NAND2X1 U1701 ( .A(n1302), .B(N102), .Y(n1259) );
  OAI21X1 U1702 ( .A(n1260), .B(n1174), .C(n1259), .Y(\DP_OP_19_294_9081/n674 ) );
  NAND2X1 U1703 ( .A(n1302), .B(N101), .Y(n1261) );
  OAI21X1 U1704 ( .A(n1262), .B(n1174), .C(n1261), .Y(\DP_OP_19_294_9081/n673 ) );
  NAND2X1 U1705 ( .A(n1302), .B(N100), .Y(n1263) );
  OAI21X1 U1706 ( .A(n1264), .B(n1174), .C(n1263), .Y(\DP_OP_19_294_9081/n672 ) );
  NAND2X1 U1707 ( .A(n1302), .B(N99), .Y(n1265) );
  OAI21X1 U1708 ( .A(n1266), .B(n1174), .C(n1265), .Y(\DP_OP_19_294_9081/n671 ) );
  NAND2X1 U1709 ( .A(n1302), .B(N98), .Y(n1267) );
  OAI21X1 U1710 ( .A(n1268), .B(n1174), .C(n1267), .Y(\DP_OP_19_294_9081/n670 ) );
  NAND2X1 U1711 ( .A(n1302), .B(N97), .Y(n1269) );
  OAI21X1 U1712 ( .A(n1270), .B(n1174), .C(n1269), .Y(\DP_OP_19_294_9081/n669 ) );
  NAND2X1 U1713 ( .A(n1302), .B(N96), .Y(n1271) );
  OAI21X1 U1714 ( .A(n1272), .B(n1174), .C(n1271), .Y(\DP_OP_19_294_9081/n668 ) );
  NAND2X1 U1715 ( .A(mulout[14]), .B(n1173), .Y(n1274) );
  NAND2X1 U1716 ( .A(n1302), .B(N95), .Y(n1273) );
  NAND2X1 U1717 ( .A(n1274), .B(n1273), .Y(\DP_OP_19_294_9081/n667 ) );
  NAND2X1 U1718 ( .A(n1302), .B(N94), .Y(n1275) );
  OAI21X1 U1719 ( .A(n1276), .B(n1174), .C(n1275), .Y(\DP_OP_19_294_9081/n666 ) );
  NAND2X1 U1720 ( .A(n1302), .B(N93), .Y(n1277) );
  OAI21X1 U1721 ( .A(n1278), .B(n1066), .C(n1277), .Y(\DP_OP_19_294_9081/n665 ) );
  NAND2X1 U1722 ( .A(n1302), .B(N92), .Y(n1279) );
  OAI21X1 U1723 ( .A(n1280), .B(n1066), .C(n1279), .Y(\DP_OP_19_294_9081/n664 ) );
  NAND2X1 U1724 ( .A(n1302), .B(N91), .Y(n1281) );
  OAI21X1 U1725 ( .A(n1282), .B(n1066), .C(n1281), .Y(\DP_OP_19_294_9081/n663 ) );
  NAND2X1 U1726 ( .A(n1302), .B(N90), .Y(n1283) );
  OAI21X1 U1727 ( .A(n1284), .B(n1066), .C(n1283), .Y(\DP_OP_19_294_9081/n662 ) );
  NAND2X1 U1728 ( .A(n1302), .B(N89), .Y(n1285) );
  OAI21X1 U1729 ( .A(n1286), .B(n1066), .C(n1285), .Y(\DP_OP_19_294_9081/n661 ) );
  NAND2X1 U1730 ( .A(n1302), .B(N88), .Y(n1287) );
  OAI21X1 U1731 ( .A(n1288), .B(n1066), .C(n1287), .Y(\DP_OP_19_294_9081/n660 ) );
  NAND2X1 U1732 ( .A(n1302), .B(N87), .Y(n1289) );
  OAI21X1 U1733 ( .A(n1290), .B(n1066), .C(n1289), .Y(\DP_OP_19_294_9081/n659 ) );
  NAND2X1 U1734 ( .A(n1302), .B(N86), .Y(n1291) );
  OAI21X1 U1735 ( .A(n1292), .B(n1066), .C(n1291), .Y(\DP_OP_19_294_9081/n658 ) );
  NAND2X1 U1736 ( .A(n1302), .B(N85), .Y(n1293) );
  OAI21X1 U1737 ( .A(n1294), .B(n1066), .C(n1293), .Y(\DP_OP_19_294_9081/n657 ) );
  NAND2X1 U1738 ( .A(n1302), .B(N81), .Y(n1295) );
  OAI21X1 U1739 ( .A(n1296), .B(n1066), .C(n1295), .Y(\DP_OP_19_294_9081/n653 ) );
  AND2X2 U1740 ( .A(n1173), .B(acc[63]), .Y(\C2/Z_63 ) );
  NOR2X1 U1741 ( .A(n1297), .B(n1175), .Y(\C2/Z_5 ) );
  NOR2X1 U1742 ( .A(n1298), .B(n1174), .Y(\C2/Z_4 ) );
  NOR2X1 U1743 ( .A(n1299), .B(n1175), .Y(\C2/Z_3 ) );
  NOR2X1 U1744 ( .A(n1300), .B(n1175), .Y(\C2/Z_2 ) );
  NOR2X1 U1745 ( .A(n1301), .B(n1175), .Y(\C2/Z_1 ) );
  NAND2X1 U1746 ( .A(n445), .B(n629), .Y(n1306) );
  NOR2X1 U1747 ( .A(n1179), .B(n1306), .Y(n1374) );
  AOI22X1 U1748 ( .A(acc[63]), .B(n1179), .C(mulout[63]), .D(n1178), .Y(n1307)
         );
  OAI21X1 U1749 ( .A(n1176), .B(n991), .C(n1017), .Y(n281) );
  AOI22X1 U1750 ( .A(acc[62]), .B(n1179), .C(mulout[62]), .D(n1178), .Y(n1308)
         );
  OAI21X1 U1751 ( .A(n1176), .B(n1004), .C(n1308), .Y(n283) );
  AOI22X1 U1752 ( .A(acc[61]), .B(n1179), .C(mulout[61]), .D(n1178), .Y(n1309)
         );
  OAI21X1 U1753 ( .A(n1176), .B(n965), .C(n1018), .Y(n285) );
  AOI22X1 U1754 ( .A(acc[60]), .B(n1179), .C(mulout[60]), .D(n1178), .Y(n1310)
         );
  OAI21X1 U1755 ( .A(n1176), .B(n1005), .C(n1310), .Y(n287) );
  AOI22X1 U1756 ( .A(acc[59]), .B(n1179), .C(mulout[59]), .D(n1178), .Y(n1311)
         );
  OAI21X1 U1757 ( .A(n1176), .B(n967), .C(n1019), .Y(n289) );
  AOI22X1 U1758 ( .A(acc[58]), .B(n1179), .C(mulout[58]), .D(n1178), .Y(n1312)
         );
  OAI21X1 U1759 ( .A(n1176), .B(n1003), .C(n1312), .Y(n291) );
  AOI22X1 U1760 ( .A(acc[57]), .B(n1179), .C(mulout[57]), .D(n1178), .Y(n1313)
         );
  OAI21X1 U1761 ( .A(n1176), .B(n968), .C(n1020), .Y(n293) );
  AOI22X1 U1762 ( .A(acc[56]), .B(n1179), .C(mulout[56]), .D(n1178), .Y(n1314)
         );
  OAI21X1 U1763 ( .A(n1176), .B(n1006), .C(n1314), .Y(n295) );
  AOI22X1 U1764 ( .A(acc[55]), .B(n1179), .C(mulout[55]), .D(n1178), .Y(n1315)
         );
  OAI21X1 U1765 ( .A(n1176), .B(n969), .C(n1021), .Y(n297) );
  AOI22X1 U1766 ( .A(acc[54]), .B(n1179), .C(mulout[54]), .D(n1178), .Y(n1316)
         );
  OAI21X1 U1767 ( .A(n1176), .B(n1007), .C(n1316), .Y(n299) );
  AOI22X1 U1768 ( .A(acc[53]), .B(n1179), .C(mulout[53]), .D(n1178), .Y(n1317)
         );
  OAI21X1 U1769 ( .A(n1176), .B(n970), .C(n1022), .Y(n301) );
  AOI22X1 U1770 ( .A(acc[52]), .B(n1179), .C(mulout[52]), .D(n1178), .Y(n1318)
         );
  OAI21X1 U1771 ( .A(n1176), .B(n1008), .C(n1318), .Y(n303) );
  AOI22X1 U1772 ( .A(acc[51]), .B(n1179), .C(mulout[51]), .D(n1178), .Y(n1319)
         );
  OAI21X1 U1773 ( .A(n1176), .B(n971), .C(n1023), .Y(n305) );
  AOI22X1 U1774 ( .A(acc[50]), .B(n1179), .C(mulout[50]), .D(n1178), .Y(n1320)
         );
  OAI21X1 U1775 ( .A(n1176), .B(n1009), .C(n1320), .Y(n307) );
  AOI22X1 U1776 ( .A(acc[49]), .B(n1179), .C(mulout[49]), .D(n1178), .Y(n1321)
         );
  AOI22X1 U1777 ( .A(acc[48]), .B(n1179), .C(mulout[48]), .D(n1178), .Y(n1322)
         );
  OAI21X1 U1778 ( .A(n1176), .B(n1002), .C(n1322), .Y(n311) );
  AOI22X1 U1779 ( .A(acc[47]), .B(n1179), .C(mulout[47]), .D(n1178), .Y(n1323)
         );
  OAI21X1 U1780 ( .A(n1176), .B(n972), .C(n1025), .Y(n313) );
  AOI22X1 U1781 ( .A(acc[46]), .B(n1179), .C(mulout[46]), .D(n1178), .Y(n1324)
         );
  OAI21X1 U1782 ( .A(n1176), .B(n999), .C(n1324), .Y(n315) );
  AOI22X1 U1783 ( .A(acc[45]), .B(n1179), .C(mulout[45]), .D(n1178), .Y(n1325)
         );
  AOI22X1 U1784 ( .A(acc[44]), .B(n1179), .C(mulout[44]), .D(n1178), .Y(n1326)
         );
  OAI21X1 U1785 ( .A(n1176), .B(n996), .C(n1326), .Y(n319) );
  AOI22X1 U1786 ( .A(acc[43]), .B(n1179), .C(mulout[43]), .D(n1178), .Y(n1327)
         );
  AOI22X1 U1787 ( .A(acc[42]), .B(n1179), .C(mulout[42]), .D(n1178), .Y(n1328)
         );
  OAI21X1 U1788 ( .A(n1176), .B(n1000), .C(n1328), .Y(n323) );
  AOI22X1 U1789 ( .A(acc[41]), .B(n1179), .C(mulout[41]), .D(n1178), .Y(n1329)
         );
  AOI22X1 U1790 ( .A(acc[40]), .B(n1179), .C(mulout[40]), .D(n1178), .Y(n1330)
         );
  AOI22X1 U1791 ( .A(acc[39]), .B(n1179), .C(mulout[39]), .D(n1178), .Y(n1331)
         );
  AOI22X1 U1792 ( .A(acc[38]), .B(n1179), .C(mulout[38]), .D(n1178), .Y(n1332)
         );
  OAI21X1 U1793 ( .A(n1176), .B(n1001), .C(n1332), .Y(n331) );
  AOI22X1 U1794 ( .A(acc[37]), .B(n1179), .C(mulout[37]), .D(n1374), .Y(n1333)
         );
  AOI22X1 U1795 ( .A(acc[36]), .B(n1179), .C(mulout[36]), .D(n1374), .Y(n1334)
         );
  OAI21X1 U1796 ( .A(n1176), .B(n997), .C(n1334), .Y(n335) );
  AOI22X1 U1797 ( .A(acc[35]), .B(n1179), .C(mulout[35]), .D(n1374), .Y(n1335)
         );
  OAI21X1 U1798 ( .A(n1176), .B(n982), .C(n1032), .Y(n337) );
  AOI22X1 U1799 ( .A(acc[34]), .B(n1179), .C(mulout[34]), .D(n1374), .Y(n1336)
         );
  OAI21X1 U1800 ( .A(n1176), .B(n1010), .C(n1336), .Y(n339) );
  AOI22X1 U1801 ( .A(acc[33]), .B(n1179), .C(mulout[33]), .D(n1374), .Y(n1337)
         );
  AOI22X1 U1802 ( .A(acc[32]), .B(n1179), .C(mulout[32]), .D(n1374), .Y(n1338)
         );
  OAI21X1 U1803 ( .A(n1176), .B(n995), .C(n1338), .Y(n343) );
  AOI22X1 U1804 ( .A(acc[31]), .B(n1179), .C(mulout[31]), .D(n1178), .Y(n1339)
         );
  OAI21X1 U1805 ( .A(n1176), .B(n978), .C(n1339), .Y(n346) );
  AOI22X1 U1806 ( .A(acc[30]), .B(n1179), .C(mulout[30]), .D(n1374), .Y(n1340)
         );
  OAI21X1 U1807 ( .A(n1176), .B(n1011), .C(n1340), .Y(n349) );
  AOI22X1 U1808 ( .A(acc[29]), .B(n1179), .C(mulout[29]), .D(n1374), .Y(n1341)
         );
  OAI21X1 U1809 ( .A(n1176), .B(n979), .C(n1341), .Y(n352) );
  AOI22X1 U1810 ( .A(acc[28]), .B(n1179), .C(mulout[28]), .D(n1374), .Y(n1342)
         );
  OAI21X1 U1811 ( .A(n1176), .B(n987), .C(n1342), .Y(n355) );
  AOI22X1 U1812 ( .A(acc[27]), .B(n1179), .C(mulout[27]), .D(n1374), .Y(n1343)
         );
  OAI21X1 U1813 ( .A(n1176), .B(n973), .C(n1343), .Y(n358) );
  AOI22X1 U1814 ( .A(acc[26]), .B(n1179), .C(mulout[26]), .D(n1374), .Y(n1344)
         );
  OAI21X1 U1815 ( .A(n1176), .B(n1012), .C(n1344), .Y(n361) );
  AOI22X1 U1816 ( .A(acc[25]), .B(n1179), .C(mulout[25]), .D(n1374), .Y(n1345)
         );
  OAI21X1 U1817 ( .A(n1176), .B(n974), .C(n1345), .Y(n364) );
  AOI22X1 U1818 ( .A(acc[24]), .B(n1179), .C(mulout[24]), .D(n1374), .Y(n1346)
         );
  OAI21X1 U1819 ( .A(n1176), .B(n988), .C(n1346), .Y(n367) );
  AOI22X1 U1820 ( .A(acc[23]), .B(n1179), .C(mulout[23]), .D(n1374), .Y(n1347)
         );
  OAI21X1 U1821 ( .A(n1176), .B(n975), .C(n1347), .Y(n370) );
  AOI22X1 U1822 ( .A(acc[22]), .B(n1179), .C(mulout[22]), .D(n1374), .Y(n1348)
         );
  OAI21X1 U1823 ( .A(n1176), .B(n1013), .C(n1348), .Y(n373) );
  AOI22X1 U1824 ( .A(acc[21]), .B(n1179), .C(mulout[21]), .D(n1374), .Y(n1349)
         );
  OAI21X1 U1825 ( .A(n1176), .B(n976), .C(n1349), .Y(n376) );
  AOI22X1 U1826 ( .A(acc[20]), .B(n1179), .C(mulout[20]), .D(n1374), .Y(n1350)
         );
  OAI21X1 U1827 ( .A(n1176), .B(n989), .C(n1350), .Y(n379) );
  AOI22X1 U1828 ( .A(acc[19]), .B(n1179), .C(mulout[19]), .D(n1374), .Y(n1351)
         );
  OAI21X1 U1829 ( .A(n1176), .B(n977), .C(n1351), .Y(n382) );
  AOI22X1 U1830 ( .A(acc[18]), .B(n1179), .C(mulout[18]), .D(n1374), .Y(n1352)
         );
  OAI21X1 U1831 ( .A(n1176), .B(n1016), .C(n1352), .Y(n385) );
  AOI22X1 U1832 ( .A(acc[17]), .B(n1179), .C(mulout[17]), .D(n1374), .Y(n1353)
         );
  OAI21X1 U1833 ( .A(n1176), .B(n994), .C(n1353), .Y(n388) );
  AOI22X1 U1834 ( .A(acc[16]), .B(n1179), .C(mulout[16]), .D(n1374), .Y(n1354)
         );
  OAI21X1 U1835 ( .A(n1176), .B(n998), .C(n1354), .Y(n391) );
  AOI22X1 U1836 ( .A(acc[15]), .B(n1179), .C(mulout[15]), .D(n1374), .Y(n1355)
         );
  OAI21X1 U1837 ( .A(n1176), .B(n966), .C(n1355), .Y(n394) );
  AOI22X1 U1838 ( .A(acc[14]), .B(n1179), .C(mulout[14]), .D(n1374), .Y(n1356)
         );
  OAI21X1 U1839 ( .A(n1176), .B(n1014), .C(n1356), .Y(n397) );
  AOI22X1 U1840 ( .A(acc[13]), .B(n1179), .C(mulout[13]), .D(n1374), .Y(n1357)
         );
  OAI21X1 U1841 ( .A(n1176), .B(n980), .C(n1357), .Y(n400) );
  AOI22X1 U1842 ( .A(acc[12]), .B(n1179), .C(mulout[12]), .D(n1374), .Y(n1358)
         );
  OAI21X1 U1843 ( .A(n1176), .B(n990), .C(n1358), .Y(n403) );
  AOI22X1 U1844 ( .A(acc[11]), .B(n1179), .C(mulout[11]), .D(n1178), .Y(n1359)
         );
  OAI21X1 U1845 ( .A(n1176), .B(n992), .C(n1359), .Y(n406) );
  AOI22X1 U1846 ( .A(acc[10]), .B(n1179), .C(mulout[10]), .D(n1178), .Y(n1360)
         );
  OAI21X1 U1847 ( .A(n1176), .B(n984), .C(n1360), .Y(n409) );
  AOI22X1 U1848 ( .A(acc[9]), .B(n1179), .C(mulout[9]), .D(n1178), .Y(n1361)
         );
  OAI21X1 U1849 ( .A(n1176), .B(n983), .C(n1361), .Y(n412) );
  AOI22X1 U1850 ( .A(acc[8]), .B(n1179), .C(mulout[8]), .D(n1178), .Y(n1362)
         );
  OAI21X1 U1851 ( .A(n1176), .B(n985), .C(n1362), .Y(n415) );
  AOI22X1 U1852 ( .A(acc[7]), .B(n1179), .C(mulout[7]), .D(n1178), .Y(n1363)
         );
  OAI21X1 U1853 ( .A(n1176), .B(n981), .C(n1363), .Y(n418) );
  AOI22X1 U1854 ( .A(acc[6]), .B(n1179), .C(mulout[6]), .D(n1178), .Y(n1364)
         );
  OAI21X1 U1855 ( .A(n1176), .B(n1015), .C(n1364), .Y(n421) );
  NOR2X1 U1856 ( .A(n1297), .B(push_2), .Y(n1365) );
  AOI21X1 U1857 ( .A(mulout[5]), .B(n1178), .C(n1365), .Y(n1366) );
  OAI21X1 U1858 ( .A(n1176), .B(n993), .C(n1366), .Y(n424) );
  NOR2X1 U1859 ( .A(n1298), .B(push_2), .Y(n1367) );
  AOI21X1 U1860 ( .A(mulout[4]), .B(n1178), .C(n1367), .Y(n1368) );
  OAI21X1 U1861 ( .A(n1176), .B(n986), .C(n1368), .Y(n427) );
  NAND2X1 U1862 ( .A(mulout[3]), .B(n1178), .Y(n1369) );
  NAND2X1 U1863 ( .A(mulout[2]), .B(n1178), .Y(n1370) );
  NAND2X1 U1864 ( .A(mulout[1]), .B(n1178), .Y(n1371) );
  OAI21X1 U1865 ( .A(push_2), .B(n1301), .C(n1371), .Y(n1372) );
  AOI21X1 U1866 ( .A(n1172), .B(\C2/DATA3_1 ), .C(n1372), .Y(n1373) );
  NAND2X1 U1867 ( .A(mulout[0]), .B(n1178), .Y(n1375) );
  NAND2X1 U1868 ( .A(h1[1]), .B(n630), .Y(n76) );
  NAND2X1 U1869 ( .A(h1[2]), .B(n630), .Y(n74) );
  NAND2X1 U1870 ( .A(h1[6]), .B(n630), .Y(n66) );
endmodule

