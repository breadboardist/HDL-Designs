
module sfilt_DW01_add_2 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n3, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n136, n137, n138, n139, n140, n141, n142,
         n143, n145, n148, n149, n150, n151, n152, n153, n154, n156, n157,
         n158, n159, n160, n161, n162, n163, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n182, n183,
         n184, n185, n186, n187, n188, n189, n191, n194, n195, n196, n197,
         n198, n199, n200, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n238,
         n239, n240, n241, n242, n243, n246, n247, n248, n249, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n270, n271, n272, n273, n274, n275, n276, n277,
         n279, n282, n283, n284, n285, n286, n287, n288, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n326, n327, n328, n329, n330, n331, n334,
         n335, n336, n337, n338, n339, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n354, n355, n356, n357, n358, n359, n360,
         n363, n364, n365, n366, n367, n368, n369, n372, n373, n376, n377,
         n378, n379, n382, n383, n384, n385, n386, n387, n388, n389, n392,
         n393, n394, n395, n397, n400, n401, n402, n404, n405, n406, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n428, n429, n430, n431, n432,
         n433, n434, n435, n437, n440, n441, n442, n443, n444, n445, n446,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n484, n485, n486, n487,
         n488, n489, n492, n493, n494, n495, n496, n497, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n512, n513, n514, n515,
         n516, n517, n518, n521, n522, n523, n524, n525, n526, n527, n530,
         n531, n534, n535, n536, n537, n540, n541, n542, n543, n544, n545,
         n546, n547, n550, n551, n552, n553, n555, n558, n559, n560, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n583, n584, n585, n586,
         n587, n588, n590, n593, n594, n595, n596, n597, n599, n600, n601,
         n602, n603, n604, n605, n606, n609, n610, n611, n612, n613, n614,
         n615, n617, n618, n619, n620, n621, n622, n623, n624, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n648, n649, n650, n651, n653, n656, n657,
         n658, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n940, n941, n942;

  COND1X1 U126 ( .A(n166), .B(n209), .C(n167), .Z(n8) );
  COND1X1 U238 ( .A(n254), .B(n297), .C(n255), .Z(n253) );
  COND1X1 U350 ( .A(n342), .B(n377), .C(n343), .Z(n337) );
  COND1X1 U556 ( .A(n500), .B(n535), .C(n501), .Z(n495) );
  CANR1X1 U647 ( .A(n635), .B(n567), .C(n568), .Z(n566) );
  COND1X1 U740 ( .A(n636), .B(n664), .C(n637), .Z(n635) );
  COND1XL U809 ( .A(n569), .B(n604), .C(n570), .Z(n568) );
  CANR1X1 U810 ( .A(n673), .B(n665), .C(n666), .Z(n664) );
  COND1X1 U811 ( .A(n677), .B(n674), .C(n675), .Z(n673) );
  CANR1XL U812 ( .A(n624), .B(n609), .C(n610), .Z(n604) );
  CIVXL U813 ( .A(n624), .Z(n622) );
  COND1X1 U814 ( .A(n633), .B(n629), .C(n630), .Z(n624) );
  CIVXL U815 ( .A(n604), .Z(n606) );
  CND2XL U816 ( .A(n623), .B(n609), .Z(n603) );
  CNR2X1 U817 ( .A(n632), .B(n629), .Z(n623) );
  CND2XL U818 ( .A(n623), .B(n731), .Z(n614) );
  CIVXL U819 ( .A(n623), .Z(n621) );
  CIVX1 U820 ( .A(n566), .Z(n565) );
  CND2XL U821 ( .A(n177), .B(n210), .Z(n175) );
  CNR2XL U822 ( .A(n225), .B(n216), .Z(n214) );
  CNR2XL U823 ( .A(B[8]), .B(A[8]), .Z(n632) );
  CND2XL U824 ( .A(B[34]), .B(A[34]), .Z(n392) );
  CND2XL U825 ( .A(B[54]), .B(A[54]), .Z(n182) );
  CND2XL U826 ( .A(B[2]), .B(A[2]), .Z(n671) );
  CNR2X1 U827 ( .A(B[24]), .B(A[24]), .Z(n489) );
  CNR2X1 U828 ( .A(B[12]), .B(A[12]), .Z(n600) );
  CNR2X1 U829 ( .A(B[28]), .B(A[28]), .Z(n449) );
  CANR1X1 U830 ( .A(n553), .B(n540), .C(n541), .Z(n535) );
  COND1X1 U831 ( .A(n601), .B(n593), .C(n594), .Z(n588) );
  CNR2XL U832 ( .A(n489), .B(n484), .Z(n478) );
  CNR2XL U833 ( .A(n449), .B(n440), .Z(n434) );
  CNR2XL U834 ( .A(n661), .B(n656), .Z(n650) );
  CNR2XL U835 ( .A(B[4]), .B(A[4]), .Z(n661) );
  CND2XL U836 ( .A(B[46]), .B(A[46]), .Z(n270) );
  CND2XL U837 ( .A(B[58]), .B(A[58]), .Z(n136) );
  CND2X1 U838 ( .A(n336), .B(n252), .Z(n7) );
  CANR1XL U839 ( .A(n360), .B(n379), .C(n363), .Z(n359) );
  CANR1XL U840 ( .A(n495), .B(n410), .C(n411), .Z(n409) );
  CND2X1 U841 ( .A(n423), .B(n456), .Z(n421) );
  CANR1XL U842 ( .A(n277), .B(n256), .C(n257), .Z(n255) );
  CANR1XL U843 ( .A(n143), .B(n122), .C(n123), .Z(n10) );
  COND1XL U844 ( .A(n450), .B(n440), .C(n441), .Z(n435) );
  COND1XL U845 ( .A(n662), .B(n656), .C(n657), .Z(n651) );
  CNR2X1 U846 ( .A(B[40]), .B(A[40]), .Z(n331) );
  CNR2X1 U847 ( .A(B[44]), .B(A[44]), .Z(n291) );
  CND2X1 U848 ( .A(B[36]), .B(A[36]), .Z(n372) );
  CNR2XL U849 ( .A(n7), .B(n162), .Z(n160) );
  CND2XL U850 ( .A(n9), .B(n96), .Z(n94) );
  CND2XL U851 ( .A(n9), .B(n120), .Z(n118) );
  CNR2XL U852 ( .A(n496), .B(n421), .Z(n419) );
  CNR2XL U853 ( .A(n338), .B(n263), .Z(n261) );
  CNIVX2 U854 ( .A(n3), .Z(n942) );
  CND2XL U855 ( .A(n378), .B(n360), .Z(n358) );
  CND2XL U856 ( .A(n536), .B(n518), .Z(n516) );
  CND2XL U857 ( .A(n9), .B(n131), .Z(n129) );
  CND2XL U858 ( .A(n9), .B(n142), .Z(n140) );
  CND2XL U859 ( .A(n9), .B(n685), .Z(n153) );
  CND2XL U860 ( .A(n232), .B(n691), .Z(n221) );
  CND2XL U861 ( .A(n320), .B(n699), .Z(n309) );
  CND2XL U862 ( .A(n478), .B(n715), .Z(n467) );
  CND2XL U863 ( .A(n210), .B(n188), .Z(n186) );
  CND2XL U864 ( .A(n605), .B(n587), .Z(n585) );
  CANR1X1 U865 ( .A(n321), .B(n302), .C(n303), .Z(n297) );
  CANR1X1 U866 ( .A(n395), .B(n382), .C(n383), .Z(n377) );
  CNR2XL U867 ( .A(n670), .B(n667), .Z(n665) );
  CANR1X1 U868 ( .A(n479), .B(n460), .C(n461), .Z(n455) );
  CNR2XL U869 ( .A(n645), .B(n640), .Z(n638) );
  CND2XL U870 ( .A(n650), .B(n638), .Z(n636) );
  CNR2XL U871 ( .A(n547), .B(n542), .Z(n540) );
  CNR2XL U872 ( .A(n471), .B(n462), .Z(n460) );
  CNR2XL U873 ( .A(n618), .B(n611), .Z(n609) );
  CANR1X1 U874 ( .A(n233), .B(n214), .C(n215), .Z(n209) );
  CNR2XL U875 ( .A(n331), .B(n326), .Z(n320) );
  CNR2XL U876 ( .A(n157), .B(n148), .Z(n142) );
  CNR2XL U877 ( .A(n291), .B(n282), .Z(n276) );
  CNR2XL U878 ( .A(n111), .B(n102), .Z(n100) );
  CNR2XL U879 ( .A(n563), .B(n558), .Z(n552) );
  CNR2XL U880 ( .A(n405), .B(n400), .Z(n394) );
  CNR2XL U881 ( .A(n509), .B(n504), .Z(n502) );
  CNR2XL U882 ( .A(n313), .B(n304), .Z(n302) );
  CNR2XL U883 ( .A(n389), .B(n384), .Z(n382) );
  CNR2XL U884 ( .A(n351), .B(n346), .Z(n344) );
  CNR2XL U885 ( .A(n267), .B(n258), .Z(n256) );
  CNR2XL U886 ( .A(n425), .B(n416), .Z(n414) );
  CNR2XL U887 ( .A(n133), .B(n124), .Z(n122) );
  CNR2IXL U888 ( .B(n142), .A(n133), .Z(n131) );
  CND2XL U889 ( .A(B[18]), .B(A[18]), .Z(n550) );
  CND2XL U890 ( .A(B[17]), .B(A[17]), .Z(n559) );
  CND2XL U891 ( .A(B[19]), .B(A[19]), .Z(n543) );
  CND2XL U892 ( .A(B[27]), .B(A[27]), .Z(n463) );
  CND2XL U893 ( .A(B[1]), .B(A[1]), .Z(n675) );
  CEOXL U894 ( .A(n12), .B(n78), .Z(SUM[63]) );
  CEOXL U895 ( .A(n13), .B(n91), .Z(SUM[62]) );
  CND2XL U896 ( .A(n940), .B(n90), .Z(n13) );
  CEOXL U897 ( .A(n14), .B(n104), .Z(SUM[61]) );
  CEOXL U898 ( .A(n15), .B(n115), .Z(SUM[60]) );
  CND2XL U899 ( .A(n681), .B(n114), .Z(n15) );
  CEOXL U900 ( .A(n16), .B(n126), .Z(SUM[59]) );
  CEOXL U901 ( .A(n17), .B(n137), .Z(SUM[58]) );
  CEOXL U902 ( .A(n18), .B(n150), .Z(SUM[57]) );
  CEOXL U903 ( .A(n19), .B(n159), .Z(SUM[56]) );
  CEOXL U904 ( .A(n20), .B(n172), .Z(SUM[55]) );
  CEOXL U905 ( .A(n21), .B(n183), .Z(SUM[54]) );
  CEOXL U906 ( .A(n22), .B(n196), .Z(SUM[53]) );
  CND2XL U907 ( .A(n688), .B(n195), .Z(n22) );
  CEOXL U908 ( .A(n23), .B(n205), .Z(SUM[52]) );
  CEOXL U909 ( .A(n24), .B(n218), .Z(SUM[51]) );
  CEOXL U910 ( .A(n25), .B(n227), .Z(SUM[50]) );
  CEOXL U911 ( .A(n26), .B(n240), .Z(SUM[49]) );
  CEOXL U912 ( .A(n27), .B(n247), .Z(SUM[48]) );
  CND2XL U913 ( .A(n693), .B(n246), .Z(n27) );
  CEOXL U914 ( .A(n28), .B(n260), .Z(SUM[47]) );
  CEOXL U915 ( .A(n29), .B(n271), .Z(SUM[46]) );
  CEOXL U916 ( .A(n30), .B(n284), .Z(SUM[45]) );
  CEOXL U917 ( .A(n31), .B(n293), .Z(SUM[44]) );
  CEOXL U918 ( .A(n32), .B(n306), .Z(SUM[43]) );
  CEOXL U919 ( .A(n33), .B(n315), .Z(SUM[42]) );
  CEOXL U920 ( .A(n34), .B(n328), .Z(SUM[41]) );
  CEOXL U921 ( .A(n35), .B(n335), .Z(SUM[40]) );
  CND2XL U922 ( .A(n701), .B(n334), .Z(n35) );
  CEOXL U923 ( .A(n36), .B(n348), .Z(SUM[39]) );
  CEOXL U924 ( .A(n37), .B(n355), .Z(SUM[38]) );
  CEOXL U925 ( .A(n38), .B(n366), .Z(SUM[37]) );
  CEOXL U926 ( .A(n39), .B(n373), .Z(SUM[36]) );
  CEOXL U927 ( .A(n40), .B(n386), .Z(SUM[35]) );
  CEOXL U928 ( .A(n41), .B(n393), .Z(SUM[34]) );
  CEOXL U929 ( .A(n42), .B(n402), .Z(SUM[33]) );
  CNR2XL U930 ( .A(B[48]), .B(A[48]), .Z(n243) );
  CNR2XL U931 ( .A(B[16]), .B(A[16]), .Z(n563) );
  CNR2XL U932 ( .A(B[32]), .B(A[32]), .Z(n405) );
  CNR2XL U933 ( .A(B[56]), .B(A[56]), .Z(n157) );
  CND2XL U934 ( .A(B[22]), .B(A[22]), .Z(n512) );
  CND2XL U935 ( .A(B[20]), .B(A[20]), .Z(n530) );
  CND2XL U936 ( .A(B[30]), .B(A[30]), .Z(n428) );
  CND2XL U937 ( .A(B[38]), .B(A[38]), .Z(n354) );
  CND2XL U938 ( .A(B[57]), .B(A[57]), .Z(n149) );
  CND2XL U939 ( .A(B[21]), .B(A[21]), .Z(n523) );
  CND2XL U940 ( .A(B[29]), .B(A[29]), .Z(n441) );
  CND2XL U941 ( .A(B[49]), .B(A[49]), .Z(n239) );
  CND2XL U942 ( .A(B[33]), .B(A[33]), .Z(n401) );
  CND2XL U943 ( .A(B[41]), .B(A[41]), .Z(n327) );
  CND2XL U944 ( .A(B[31]), .B(A[31]), .Z(n417) );
  CND2XL U945 ( .A(B[35]), .B(A[35]), .Z(n385) );
  CND2XL U946 ( .A(B[51]), .B(A[51]), .Z(n217) );
  CND2XL U947 ( .A(B[59]), .B(A[59]), .Z(n125) );
  CND2XL U948 ( .A(B[43]), .B(A[43]), .Z(n305) );
  CND2XL U949 ( .A(B[45]), .B(A[45]), .Z(n283) );
  CND2XL U950 ( .A(B[47]), .B(A[47]), .Z(n259) );
  CND2XL U951 ( .A(B[55]), .B(A[55]), .Z(n171) );
  CND2XL U952 ( .A(B[39]), .B(A[39]), .Z(n347) );
  CND2XL U953 ( .A(B[61]), .B(A[61]), .Z(n103) );
  CND2XL U954 ( .A(B[37]), .B(A[37]), .Z(n365) );
  CND2XL U955 ( .A(B[6]), .B(A[6]), .Z(n648) );
  CND2XL U956 ( .A(B[14]), .B(A[14]), .Z(n583) );
  CND2XL U957 ( .A(B[63]), .B(A[63]), .Z(n77) );
  CEOXL U958 ( .A(n52), .B(n506), .Z(SUM[23]) );
  CEOXL U959 ( .A(n53), .B(n513), .Z(SUM[22]) );
  CND2XL U960 ( .A(n719), .B(n512), .Z(n53) );
  CEOXL U961 ( .A(n44), .B(n418), .Z(SUM[31]) );
  CND2XL U962 ( .A(n710), .B(n417), .Z(n44) );
  CEOXL U963 ( .A(n45), .B(n429), .Z(SUM[30]) );
  CND2XL U964 ( .A(n711), .B(n428), .Z(n45) );
  CEOXL U965 ( .A(n46), .B(n442), .Z(SUM[29]) );
  CND2XL U966 ( .A(n712), .B(n441), .Z(n46) );
  CEOXL U967 ( .A(n47), .B(n451), .Z(SUM[28]) );
  CEOXL U968 ( .A(n48), .B(n464), .Z(SUM[27]) );
  CND2XL U969 ( .A(n714), .B(n463), .Z(n48) );
  CEOXL U970 ( .A(n49), .B(n473), .Z(SUM[26]) );
  CEOXL U971 ( .A(n50), .B(n486), .Z(SUM[25]) );
  CEOXL U972 ( .A(n51), .B(n493), .Z(SUM[24]) );
  CEOXL U973 ( .A(n54), .B(n524), .Z(SUM[21]) );
  CND2XL U974 ( .A(n720), .B(n523), .Z(n54) );
  CEOXL U975 ( .A(n55), .B(n531), .Z(SUM[20]) );
  CND2XL U976 ( .A(n721), .B(n530), .Z(n55) );
  CEOXL U977 ( .A(n56), .B(n544), .Z(SUM[19]) );
  CND2XL U978 ( .A(n722), .B(n543), .Z(n56) );
  CEOXL U979 ( .A(n57), .B(n551), .Z(SUM[18]) );
  CND2XL U980 ( .A(n723), .B(n550), .Z(n57) );
  CEOXL U981 ( .A(n58), .B(n560), .Z(SUM[17]) );
  CND2XL U982 ( .A(n724), .B(n559), .Z(n58) );
  CEOXL U983 ( .A(n68), .B(n642), .Z(SUM[7]) );
  CEOXL U984 ( .A(n69), .B(n649), .Z(SUM[6]) );
  CEOXL U985 ( .A(n70), .B(n658), .Z(SUM[5]) );
  CND2IXL U986 ( .B(n676), .A(n677), .Z(n75) );
  CNR2X1 U987 ( .A(n7), .B(n94), .Z(n92) );
  CNR2X1 U988 ( .A(n7), .B(n118), .Z(n116) );
  CNR2XL U989 ( .A(n7), .B(n81), .Z(n79) );
  CNR2X1 U990 ( .A(n208), .B(n166), .Z(n9) );
  CNR2X1 U991 ( .A(n376), .B(n342), .Z(n336) );
  CNR2X1 U992 ( .A(n296), .B(n254), .Z(n252) );
  CNR2X1 U993 ( .A(n534), .B(n500), .Z(n494) );
  CNR2X1 U994 ( .A(n11), .B(n98), .Z(n96) );
  CNR2X1 U995 ( .A(n454), .B(n412), .Z(n410) );
  CNR2XL U996 ( .A(n7), .B(n107), .Z(n105) );
  CNR2XL U997 ( .A(n7), .B(n129), .Z(n127) );
  CNR2XL U998 ( .A(n7), .B(n140), .Z(n138) );
  CNR2XL U999 ( .A(n7), .B(n153), .Z(n151) );
  CNR2XL U1000 ( .A(n7), .B(n175), .Z(n173) );
  CNR2XL U1001 ( .A(n7), .B(n186), .Z(n184) );
  CNR2XL U1002 ( .A(n7), .B(n199), .Z(n197) );
  CNR2XL U1003 ( .A(n7), .B(n208), .Z(n206) );
  CNR2XL U1004 ( .A(n7), .B(n221), .Z(n219) );
  CNR2XL U1005 ( .A(n7), .B(n230), .Z(n228) );
  CNR2XL U1006 ( .A(n338), .B(n274), .Z(n272) );
  CNR2XL U1007 ( .A(n338), .B(n287), .Z(n285) );
  CNR2XL U1008 ( .A(n338), .B(n296), .Z(n294) );
  CNR2XL U1009 ( .A(n338), .B(n309), .Z(n307) );
  CNR2XL U1010 ( .A(n338), .B(n318), .Z(n316) );
  CNR2XL U1011 ( .A(n496), .B(n432), .Z(n430) );
  CNR2XL U1012 ( .A(n496), .B(n445), .Z(n443) );
  CNR2XL U1013 ( .A(n496), .B(n454), .Z(n452) );
  CNR2XL U1014 ( .A(n496), .B(n467), .Z(n465) );
  CNR2XL U1015 ( .A(n496), .B(n476), .Z(n474) );
  CND2XL U1016 ( .A(n9), .B(n83), .Z(n81) );
  CANR1XL U1017 ( .A(n494), .B(n565), .C(n495), .Z(n493) );
  CNR2X1 U1018 ( .A(n603), .B(n569), .Z(n567) );
  CND2X1 U1019 ( .A(n587), .B(n571), .Z(n569) );
  CANR1XL U1020 ( .A(n518), .B(n537), .C(n521), .Z(n517) );
  CANR1XL U1021 ( .A(n587), .B(n606), .C(n588), .Z(n586) );
  COND1XL U1022 ( .A(n408), .B(n566), .C(n409), .Z(n3) );
  CND2XL U1023 ( .A(n494), .B(n410), .Z(n408) );
  CNR2X1 U1024 ( .A(n11), .B(n85), .Z(n83) );
  CND2X1 U1025 ( .A(n142), .B(n122), .Z(n11) );
  COND1XL U1026 ( .A(n94), .B(n5), .C(n95), .Z(n93) );
  CANR1XL U1027 ( .A(n96), .B(n8), .C(n97), .Z(n95) );
  COND1XL U1028 ( .A(n98), .B(n10), .C(n99), .Z(n97) );
  COND1XL U1029 ( .A(n118), .B(n5), .C(n119), .Z(n117) );
  CANR1XL U1030 ( .A(n120), .B(n8), .C(n121), .Z(n119) );
  COND1XL U1031 ( .A(n140), .B(n5), .C(n141), .Z(n139) );
  CANR1XL U1032 ( .A(n142), .B(n8), .C(n143), .Z(n141) );
  COND1XL U1033 ( .A(n162), .B(n5), .C(n163), .Z(n161) );
  COND1XL U1034 ( .A(n186), .B(n5), .C(n187), .Z(n185) );
  CANR1XL U1035 ( .A(n188), .B(n211), .C(n189), .Z(n187) );
  COND1XL U1036 ( .A(n208), .B(n5), .C(n209), .Z(n207) );
  COND1XL U1037 ( .A(n230), .B(n5), .C(n231), .Z(n229) );
  COND1XL U1038 ( .A(n274), .B(n339), .C(n275), .Z(n273) );
  CANR1XL U1039 ( .A(n276), .B(n299), .C(n277), .Z(n275) );
  COND1XL U1040 ( .A(n296), .B(n339), .C(n297), .Z(n295) );
  COND1XL U1041 ( .A(n318), .B(n339), .C(n319), .Z(n317) );
  COND1XL U1042 ( .A(n432), .B(n497), .C(n433), .Z(n431) );
  CANR1XL U1043 ( .A(n434), .B(n457), .C(n435), .Z(n433) );
  COND1XL U1044 ( .A(n454), .B(n497), .C(n455), .Z(n453) );
  COND1XL U1045 ( .A(n476), .B(n497), .C(n477), .Z(n475) );
  CND2X1 U1046 ( .A(n232), .B(n214), .Z(n208) );
  CND2X1 U1047 ( .A(n320), .B(n302), .Z(n296) );
  CND2X1 U1048 ( .A(n478), .B(n460), .Z(n454) );
  CND2X1 U1049 ( .A(n552), .B(n540), .Z(n534) );
  CND2X1 U1050 ( .A(n394), .B(n382), .Z(n376) );
  CND2X1 U1051 ( .A(n518), .B(n502), .Z(n500) );
  CND2X1 U1052 ( .A(n360), .B(n344), .Z(n342) );
  CND2X1 U1053 ( .A(n276), .B(n256), .Z(n254) );
  CND2X1 U1054 ( .A(n188), .B(n168), .Z(n166) );
  CND2X1 U1055 ( .A(n434), .B(n414), .Z(n412) );
  CND2XL U1056 ( .A(n9), .B(n109), .Z(n107) );
  CND2X1 U1057 ( .A(n210), .B(n689), .Z(n199) );
  CND2X1 U1058 ( .A(n298), .B(n276), .Z(n274) );
  CND2X1 U1059 ( .A(n298), .B(n697), .Z(n287) );
  CND2X1 U1060 ( .A(n456), .B(n434), .Z(n432) );
  CND2X1 U1061 ( .A(n456), .B(n713), .Z(n445) );
  CND2X1 U1062 ( .A(n265), .B(n298), .Z(n263) );
  CND2XL U1063 ( .A(n605), .B(n729), .Z(n596) );
  CND2XL U1064 ( .A(n578), .B(n605), .Z(n576) );
  COND1XL U1065 ( .A(n270), .B(n258), .C(n259), .Z(n257) );
  CANR1XL U1066 ( .A(n189), .B(n168), .C(n169), .Z(n167) );
  COND1XL U1067 ( .A(n182), .B(n170), .C(n171), .Z(n169) );
  COND1XL U1068 ( .A(n136), .B(n124), .C(n125), .Z(n123) );
  CANR1XL U1069 ( .A(n363), .B(n344), .C(n345), .Z(n343) );
  COND1XL U1070 ( .A(n354), .B(n346), .C(n347), .Z(n345) );
  CANR1XL U1071 ( .A(n487), .B(n565), .C(n488), .Z(n486) );
  CNR2XL U1072 ( .A(n496), .B(n489), .Z(n487) );
  COND1XL U1073 ( .A(n489), .B(n497), .C(n492), .Z(n488) );
  CANR1XL U1074 ( .A(n507), .B(n565), .C(n508), .Z(n506) );
  CNR2XL U1075 ( .A(n516), .B(n509), .Z(n507) );
  COND1XL U1076 ( .A(n509), .B(n517), .C(n512), .Z(n508) );
  COND1XL U1077 ( .A(n619), .B(n611), .C(n612), .Z(n610) );
  COND1XL U1078 ( .A(n314), .B(n304), .C(n305), .Z(n303) );
  COND1XL U1079 ( .A(n226), .B(n216), .C(n217), .Z(n215) );
  COND1XL U1080 ( .A(n472), .B(n462), .C(n463), .Z(n461) );
  COND1XL U1081 ( .A(n550), .B(n542), .C(n543), .Z(n541) );
  COND1XL U1082 ( .A(n392), .B(n384), .C(n385), .Z(n383) );
  CANR1XL U1083 ( .A(n521), .B(n502), .C(n503), .Z(n501) );
  COND1XL U1084 ( .A(n512), .B(n504), .C(n505), .Z(n503) );
  COND1XL U1085 ( .A(n292), .B(n282), .C(n283), .Z(n277) );
  COND1XL U1086 ( .A(n406), .B(n400), .C(n401), .Z(n395) );
  COND1XL U1087 ( .A(n564), .B(n558), .C(n559), .Z(n553) );
  COND1XL U1088 ( .A(n204), .B(n194), .C(n195), .Z(n189) );
  COND1XL U1089 ( .A(n158), .B(n148), .C(n149), .Z(n143) );
  COND1XL U1090 ( .A(n334), .B(n326), .C(n327), .Z(n321) );
  COND1XL U1091 ( .A(n492), .B(n484), .C(n485), .Z(n479) );
  COND1XL U1092 ( .A(n246), .B(n238), .C(n239), .Z(n233) );
  COND1XL U1093 ( .A(n671), .B(n667), .C(n668), .Z(n666) );
  CNR2X1 U1094 ( .A(n600), .B(n593), .Z(n587) );
  CNR2X1 U1095 ( .A(n203), .B(n194), .Z(n188) );
  CANR1XL U1096 ( .A(n651), .B(n638), .C(n639), .Z(n637) );
  COND1XL U1097 ( .A(n114), .B(n102), .C(n103), .Z(n101) );
  CNR2X1 U1098 ( .A(n243), .B(n238), .Z(n232) );
  CNR2X1 U1099 ( .A(n527), .B(n522), .Z(n518) );
  CNR2X1 U1100 ( .A(n369), .B(n364), .Z(n360) );
  COND1XL U1101 ( .A(n530), .B(n522), .C(n523), .Z(n521) );
  COND1XL U1102 ( .A(n372), .B(n364), .C(n365), .Z(n363) );
  CANR1XL U1103 ( .A(n588), .B(n571), .C(n572), .Z(n570) );
  COND1XL U1104 ( .A(n583), .B(n573), .C(n574), .Z(n572) );
  CANR1XL U1105 ( .A(n606), .B(n578), .C(n579), .Z(n577) );
  COND1XL U1106 ( .A(n580), .B(n590), .C(n583), .Z(n579) );
  CANR1XL U1107 ( .A(n729), .B(n606), .C(n599), .Z(n597) );
  CANR1XL U1108 ( .A(n731), .B(n624), .C(n617), .Z(n615) );
  CNR2X1 U1109 ( .A(n11), .B(n111), .Z(n109) );
  CNR2X1 U1110 ( .A(n580), .B(n573), .Z(n571) );
  CNR2X1 U1111 ( .A(n179), .B(n170), .Z(n168) );
  COND1XL U1112 ( .A(n412), .B(n455), .C(n413), .Z(n411) );
  CANR1XL U1113 ( .A(n435), .B(n414), .C(n415), .Z(n413) );
  COND1XL U1114 ( .A(n428), .B(n416), .C(n417), .Z(n415) );
  COND1XL U1115 ( .A(n648), .B(n640), .C(n641), .Z(n639) );
  COND1XL U1116 ( .A(n81), .B(n5), .C(n82), .Z(n80) );
  CANR1XL U1117 ( .A(n83), .B(n8), .C(n84), .Z(n82) );
  COND1XL U1118 ( .A(n85), .B(n10), .C(n86), .Z(n84) );
  CANR1XL U1119 ( .A(n940), .B(n101), .C(n88), .Z(n86) );
  COND1XL U1120 ( .A(n107), .B(n5), .C(n108), .Z(n106) );
  CANR1XL U1121 ( .A(n109), .B(n8), .C(n110), .Z(n108) );
  COND1XL U1122 ( .A(n111), .B(n10), .C(n114), .Z(n110) );
  COND1XL U1123 ( .A(n129), .B(n5), .C(n130), .Z(n128) );
  CANR1XL U1124 ( .A(n131), .B(n8), .C(n132), .Z(n130) );
  COND1XL U1125 ( .A(n133), .B(n145), .C(n136), .Z(n132) );
  COND1XL U1126 ( .A(n153), .B(n5), .C(n154), .Z(n152) );
  CANR1XL U1127 ( .A(n685), .B(n8), .C(n156), .Z(n154) );
  COND1XL U1128 ( .A(n175), .B(n5), .C(n176), .Z(n174) );
  CANR1XL U1129 ( .A(n211), .B(n177), .C(n178), .Z(n176) );
  COND1XL U1130 ( .A(n179), .B(n191), .C(n182), .Z(n178) );
  COND1XL U1131 ( .A(n199), .B(n5), .C(n200), .Z(n198) );
  CANR1XL U1132 ( .A(n689), .B(n211), .C(n202), .Z(n200) );
  COND1XL U1133 ( .A(n221), .B(n5), .C(n222), .Z(n220) );
  CANR1XL U1134 ( .A(n691), .B(n233), .C(n224), .Z(n222) );
  COND1XL U1135 ( .A(n243), .B(n5), .C(n246), .Z(n242) );
  COND1XL U1136 ( .A(n263), .B(n339), .C(n264), .Z(n262) );
  CANR1XL U1137 ( .A(n299), .B(n265), .C(n266), .Z(n264) );
  COND1XL U1138 ( .A(n267), .B(n279), .C(n270), .Z(n266) );
  COND1XL U1139 ( .A(n287), .B(n339), .C(n288), .Z(n286) );
  CANR1XL U1140 ( .A(n697), .B(n299), .C(n290), .Z(n288) );
  COND1XL U1141 ( .A(n309), .B(n339), .C(n310), .Z(n308) );
  CANR1XL U1142 ( .A(n699), .B(n321), .C(n312), .Z(n310) );
  COND1XL U1143 ( .A(n331), .B(n339), .C(n334), .Z(n330) );
  COND1XL U1144 ( .A(n421), .B(n497), .C(n422), .Z(n420) );
  CANR1XL U1145 ( .A(n457), .B(n423), .C(n424), .Z(n422) );
  COND1XL U1146 ( .A(n425), .B(n437), .C(n428), .Z(n424) );
  COND1XL U1147 ( .A(n445), .B(n497), .C(n446), .Z(n444) );
  CANR1XL U1148 ( .A(n713), .B(n457), .C(n448), .Z(n446) );
  COND1XL U1149 ( .A(n467), .B(n497), .C(n468), .Z(n466) );
  CANR1XL U1150 ( .A(n715), .B(n479), .C(n470), .Z(n468) );
  COND1XL U1151 ( .A(n351), .B(n359), .C(n354), .Z(n350) );
  COND1XL U1152 ( .A(n369), .B(n377), .C(n372), .Z(n368) );
  COND1XL U1153 ( .A(n527), .B(n535), .C(n530), .Z(n526) );
  COND1XL U1154 ( .A(n389), .B(n397), .C(n392), .Z(n388) );
  COND1XL U1155 ( .A(n547), .B(n555), .C(n550), .Z(n546) );
  COND1XL U1156 ( .A(n645), .B(n653), .C(n648), .Z(n644) );
  CNR2IXL U1157 ( .B(n188), .A(n179), .Z(n177) );
  CNR2IXL U1158 ( .B(n276), .A(n267), .Z(n265) );
  CNR2IXL U1159 ( .B(n434), .A(n425), .Z(n423) );
  CNR2IXL U1160 ( .B(n587), .A(n580), .Z(n578) );
  CNR2XL U1161 ( .A(n7), .B(n243), .Z(n241) );
  CNR2XL U1162 ( .A(n338), .B(n331), .Z(n329) );
  CNR2XL U1163 ( .A(n358), .B(n351), .Z(n349) );
  CNR2XL U1164 ( .A(n376), .B(n369), .Z(n367) );
  CNR2XL U1165 ( .A(n534), .B(n527), .Z(n525) );
  CNR2IXL U1166 ( .B(n394), .A(n389), .Z(n387) );
  CNR2IXL U1167 ( .B(n552), .A(n547), .Z(n545) );
  CNR2IXL U1168 ( .B(n650), .A(n645), .Z(n643) );
  CND2X1 U1169 ( .A(n100), .B(n940), .Z(n85) );
  CND2X1 U1170 ( .A(n941), .B(n77), .Z(n12) );
  CANR1XL U1171 ( .A(n79), .B(n942), .C(n80), .Z(n78) );
  CANR1XL U1172 ( .A(n92), .B(n942), .C(n93), .Z(n91) );
  CND2X1 U1173 ( .A(n680), .B(n103), .Z(n14) );
  CANR1XL U1174 ( .A(n105), .B(n942), .C(n106), .Z(n104) );
  CANR1XL U1175 ( .A(n116), .B(n942), .C(n117), .Z(n115) );
  CND2X1 U1176 ( .A(n682), .B(n125), .Z(n16) );
  CANR1XL U1177 ( .A(n127), .B(n942), .C(n128), .Z(n126) );
  CND2X1 U1178 ( .A(n683), .B(n136), .Z(n17) );
  CANR1XL U1179 ( .A(n138), .B(n942), .C(n139), .Z(n137) );
  CND2X1 U1180 ( .A(n684), .B(n149), .Z(n18) );
  CANR1XL U1181 ( .A(n151), .B(n942), .C(n152), .Z(n150) );
  CND2XL U1182 ( .A(n685), .B(n158), .Z(n19) );
  CANR1XL U1183 ( .A(n160), .B(n942), .C(n161), .Z(n159) );
  CND2X1 U1184 ( .A(n686), .B(n171), .Z(n20) );
  CANR1XL U1185 ( .A(n173), .B(n942), .C(n174), .Z(n172) );
  CND2X1 U1186 ( .A(n687), .B(n182), .Z(n21) );
  CANR1XL U1187 ( .A(n184), .B(n942), .C(n185), .Z(n183) );
  CANR1XL U1188 ( .A(n197), .B(n942), .C(n198), .Z(n196) );
  CND2XL U1189 ( .A(n689), .B(n204), .Z(n23) );
  CANR1XL U1190 ( .A(n206), .B(n942), .C(n207), .Z(n205) );
  CND2X1 U1191 ( .A(n690), .B(n217), .Z(n24) );
  CANR1XL U1192 ( .A(n219), .B(n942), .C(n220), .Z(n218) );
  CND2XL U1193 ( .A(n691), .B(n226), .Z(n25) );
  CANR1XL U1194 ( .A(n228), .B(n942), .C(n229), .Z(n227) );
  CND2X1 U1195 ( .A(n692), .B(n239), .Z(n26) );
  CANR1XL U1196 ( .A(n241), .B(n942), .C(n242), .Z(n240) );
  CANR1XL U1197 ( .A(n248), .B(n942), .C(n249), .Z(n247) );
  CND2X1 U1198 ( .A(n694), .B(n259), .Z(n28) );
  CANR1XL U1199 ( .A(n261), .B(n942), .C(n262), .Z(n260) );
  CND2X1 U1200 ( .A(n695), .B(n270), .Z(n29) );
  CANR1XL U1201 ( .A(n272), .B(n942), .C(n273), .Z(n271) );
  CND2X1 U1202 ( .A(n696), .B(n283), .Z(n30) );
  CANR1XL U1203 ( .A(n285), .B(n942), .C(n286), .Z(n284) );
  CND2XL U1204 ( .A(n697), .B(n292), .Z(n31) );
  CANR1XL U1205 ( .A(n294), .B(n942), .C(n295), .Z(n293) );
  CND2X1 U1206 ( .A(n698), .B(n305), .Z(n32) );
  CANR1XL U1207 ( .A(n307), .B(n942), .C(n308), .Z(n306) );
  CND2XL U1208 ( .A(n699), .B(n314), .Z(n33) );
  CANR1XL U1209 ( .A(n316), .B(n942), .C(n317), .Z(n315) );
  CND2X1 U1210 ( .A(n700), .B(n327), .Z(n34) );
  CANR1XL U1211 ( .A(n329), .B(n942), .C(n330), .Z(n328) );
  CANR1XL U1212 ( .A(n336), .B(n942), .C(n337), .Z(n335) );
  CND2X1 U1213 ( .A(n702), .B(n347), .Z(n36) );
  CANR1XL U1214 ( .A(n349), .B(n942), .C(n350), .Z(n348) );
  CND2X1 U1215 ( .A(n703), .B(n354), .Z(n37) );
  CANR1XL U1216 ( .A(n356), .B(n942), .C(n357), .Z(n355) );
  CND2X1 U1217 ( .A(n704), .B(n365), .Z(n38) );
  CANR1XL U1218 ( .A(n367), .B(n942), .C(n368), .Z(n366) );
  CND2X1 U1219 ( .A(n705), .B(n372), .Z(n39) );
  CANR1XL U1220 ( .A(n378), .B(n942), .C(n379), .Z(n373) );
  CND2X1 U1221 ( .A(n706), .B(n385), .Z(n40) );
  CANR1XL U1222 ( .A(n387), .B(n942), .C(n388), .Z(n386) );
  CND2X1 U1223 ( .A(n707), .B(n392), .Z(n41) );
  CANR1XL U1224 ( .A(n394), .B(n942), .C(n395), .Z(n393) );
  CND2X1 U1225 ( .A(n708), .B(n401), .Z(n42) );
  CANR1XL U1226 ( .A(n709), .B(n942), .C(n404), .Z(n402) );
  CANR1XL U1227 ( .A(n419), .B(n565), .C(n420), .Z(n418) );
  CANR1XL U1228 ( .A(n430), .B(n565), .C(n431), .Z(n429) );
  CANR1XL U1229 ( .A(n443), .B(n565), .C(n444), .Z(n442) );
  CND2XL U1230 ( .A(n713), .B(n450), .Z(n47) );
  CANR1XL U1231 ( .A(n452), .B(n565), .C(n453), .Z(n451) );
  CANR1XL U1232 ( .A(n465), .B(n565), .C(n466), .Z(n464) );
  CND2XL U1233 ( .A(n715), .B(n472), .Z(n49) );
  CANR1XL U1234 ( .A(n474), .B(n565), .C(n475), .Z(n473) );
  CANR1XL U1235 ( .A(n514), .B(n565), .C(n515), .Z(n513) );
  CANR1XL U1236 ( .A(n525), .B(n565), .C(n526), .Z(n524) );
  CANR1XL U1237 ( .A(n536), .B(n565), .C(n537), .Z(n531) );
  CANR1XL U1238 ( .A(n545), .B(n565), .C(n546), .Z(n544) );
  CANR1XL U1239 ( .A(n552), .B(n565), .C(n553), .Z(n551) );
  CANR1XL U1240 ( .A(n725), .B(n565), .C(n562), .Z(n560) );
  CNR2X1 U1241 ( .A(B[20]), .B(A[20]), .Z(n527) );
  CNR2X1 U1242 ( .A(B[34]), .B(A[34]), .Z(n389) );
  CNR2X1 U1243 ( .A(B[38]), .B(A[38]), .Z(n351) );
  CNR2X1 U1244 ( .A(B[36]), .B(A[36]), .Z(n369) );
  CNR2X1 U1245 ( .A(B[18]), .B(A[18]), .Z(n547) );
  CNR2X1 U1246 ( .A(B[46]), .B(A[46]), .Z(n267) );
  CNR2X1 U1247 ( .A(B[14]), .B(A[14]), .Z(n580) );
  CNR2X1 U1248 ( .A(B[22]), .B(A[22]), .Z(n509) );
  CNR2X1 U1249 ( .A(B[54]), .B(A[54]), .Z(n179) );
  CNR2X1 U1250 ( .A(B[6]), .B(A[6]), .Z(n645) );
  CNR2X1 U1251 ( .A(B[30]), .B(A[30]), .Z(n425) );
  CNR2X1 U1252 ( .A(B[58]), .B(A[58]), .Z(n133) );
  CNR2X1 U1253 ( .A(B[60]), .B(A[60]), .Z(n111) );
  CNR2X1 U1254 ( .A(B[23]), .B(A[23]), .Z(n504) );
  CNR2X1 U1255 ( .A(B[47]), .B(A[47]), .Z(n258) );
  CNR2X1 U1256 ( .A(B[13]), .B(A[13]), .Z(n593) );
  CNR2X1 U1257 ( .A(B[45]), .B(A[45]), .Z(n282) );
  CNR2X1 U1258 ( .A(B[41]), .B(A[41]), .Z(n326) );
  CNR2X1 U1259 ( .A(B[17]), .B(A[17]), .Z(n558) );
  CNR2X1 U1260 ( .A(B[39]), .B(A[39]), .Z(n346) );
  CNR2X1 U1261 ( .A(B[33]), .B(A[33]), .Z(n400) );
  CNR2X1 U1262 ( .A(B[49]), .B(A[49]), .Z(n238) );
  CNR2X1 U1263 ( .A(B[21]), .B(A[21]), .Z(n522) );
  CNR2X1 U1264 ( .A(B[43]), .B(A[43]), .Z(n304) );
  CNR2X1 U1265 ( .A(B[25]), .B(A[25]), .Z(n484) );
  CNR2X1 U1266 ( .A(B[37]), .B(A[37]), .Z(n364) );
  CNR2X1 U1267 ( .A(B[9]), .B(A[9]), .Z(n629) );
  CNR2X1 U1268 ( .A(B[35]), .B(A[35]), .Z(n384) );
  CNR2X1 U1269 ( .A(B[11]), .B(A[11]), .Z(n611) );
  CNR2X1 U1270 ( .A(B[53]), .B(A[53]), .Z(n194) );
  CNR2X1 U1271 ( .A(B[19]), .B(A[19]), .Z(n542) );
  CNR2X1 U1272 ( .A(B[29]), .B(A[29]), .Z(n440) );
  CNR2X1 U1273 ( .A(B[51]), .B(A[51]), .Z(n216) );
  CNR2X1 U1274 ( .A(B[27]), .B(A[27]), .Z(n462) );
  CNR2X1 U1275 ( .A(B[15]), .B(A[15]), .Z(n573) );
  CNR2X1 U1276 ( .A(B[5]), .B(A[5]), .Z(n656) );
  CNR2X1 U1277 ( .A(B[57]), .B(A[57]), .Z(n148) );
  CNR2X1 U1278 ( .A(B[55]), .B(A[55]), .Z(n170) );
  CNR2X1 U1279 ( .A(B[7]), .B(A[7]), .Z(n640) );
  CNR2X1 U1280 ( .A(B[31]), .B(A[31]), .Z(n416) );
  CNR2X1 U1281 ( .A(B[59]), .B(A[59]), .Z(n124) );
  CNR2X1 U1282 ( .A(B[61]), .B(A[61]), .Z(n102) );
  CNR2X1 U1283 ( .A(B[3]), .B(A[3]), .Z(n667) );
  CNR2X1 U1284 ( .A(B[2]), .B(A[2]), .Z(n670) );
  CNR2X1 U1285 ( .A(B[52]), .B(A[52]), .Z(n203) );
  CNR2X1 U1286 ( .A(B[42]), .B(A[42]), .Z(n313) );
  CNR2X1 U1287 ( .A(B[50]), .B(A[50]), .Z(n225) );
  CNR2X1 U1288 ( .A(B[26]), .B(A[26]), .Z(n471) );
  CNR2X1 U1289 ( .A(B[10]), .B(A[10]), .Z(n618) );
  CND2X1 U1290 ( .A(B[0]), .B(A[0]), .Z(n677) );
  CNR2X1 U1291 ( .A(B[1]), .B(A[1]), .Z(n674) );
  COR2X1 U1292 ( .A(B[62]), .B(A[62]), .Z(n940) );
  CNR2XL U1293 ( .A(B[0]), .B(A[0]), .Z(n676) );
  CND2X1 U1294 ( .A(B[10]), .B(A[10]), .Z(n619) );
  CND2X1 U1295 ( .A(B[4]), .B(A[4]), .Z(n662) );
  CND2X1 U1296 ( .A(B[16]), .B(A[16]), .Z(n564) );
  CND2X1 U1297 ( .A(B[44]), .B(A[44]), .Z(n292) );
  CND2X1 U1298 ( .A(B[32]), .B(A[32]), .Z(n406) );
  CND2X1 U1299 ( .A(B[42]), .B(A[42]), .Z(n314) );
  CND2X1 U1300 ( .A(B[12]), .B(A[12]), .Z(n601) );
  CND2X1 U1301 ( .A(B[26]), .B(A[26]), .Z(n472) );
  CND2X1 U1302 ( .A(B[28]), .B(A[28]), .Z(n450) );
  CND2X1 U1303 ( .A(B[50]), .B(A[50]), .Z(n226) );
  CND2X1 U1304 ( .A(B[52]), .B(A[52]), .Z(n204) );
  CND2X1 U1305 ( .A(B[56]), .B(A[56]), .Z(n158) );
  CND2X1 U1306 ( .A(B[8]), .B(A[8]), .Z(n633) );
  CND2X1 U1307 ( .A(B[40]), .B(A[40]), .Z(n334) );
  CND2X1 U1308 ( .A(B[24]), .B(A[24]), .Z(n492) );
  CND2X1 U1309 ( .A(B[48]), .B(A[48]), .Z(n246) );
  CND2X1 U1310 ( .A(B[60]), .B(A[60]), .Z(n114) );
  CND2X1 U1311 ( .A(B[62]), .B(A[62]), .Z(n90) );
  CND2XL U1312 ( .A(B[23]), .B(A[23]), .Z(n505) );
  CND2XL U1313 ( .A(B[11]), .B(A[11]), .Z(n612) );
  CND2XL U1314 ( .A(B[9]), .B(A[9]), .Z(n630) );
  CND2XL U1315 ( .A(B[5]), .B(A[5]), .Z(n657) );
  CND2XL U1316 ( .A(B[3]), .B(A[3]), .Z(n668) );
  CND2XL U1317 ( .A(B[13]), .B(A[13]), .Z(n594) );
  CND2XL U1318 ( .A(B[25]), .B(A[25]), .Z(n485) );
  CND2XL U1319 ( .A(B[15]), .B(A[15]), .Z(n574) );
  CND2XL U1320 ( .A(B[7]), .B(A[7]), .Z(n641) );
  CND2XL U1321 ( .A(B[53]), .B(A[53]), .Z(n195) );
  CENX1 U1322 ( .A(n942), .B(n43), .Z(SUM[32]) );
  CND2XL U1323 ( .A(n709), .B(n406), .Z(n43) );
  CND2XL U1324 ( .A(n716), .B(n485), .Z(n50) );
  CND2XL U1325 ( .A(n717), .B(n492), .Z(n51) );
  CND2XL U1326 ( .A(n718), .B(n505), .Z(n52) );
  CENX1 U1327 ( .A(n565), .B(n59), .Z(SUM[16]) );
  CND2XL U1328 ( .A(n725), .B(n564), .Z(n59) );
  CENX1 U1329 ( .A(n575), .B(n60), .Z(SUM[15]) );
  CND2XL U1330 ( .A(n726), .B(n574), .Z(n60) );
  COND1XL U1331 ( .A(n576), .B(n634), .C(n577), .Z(n575) );
  CENX1 U1332 ( .A(n584), .B(n61), .Z(SUM[14]) );
  CND2XL U1333 ( .A(n727), .B(n583), .Z(n61) );
  COND1XL U1334 ( .A(n585), .B(n634), .C(n586), .Z(n584) );
  CENX1 U1335 ( .A(n595), .B(n62), .Z(SUM[13]) );
  CND2XL U1336 ( .A(n728), .B(n594), .Z(n62) );
  COND1XL U1337 ( .A(n596), .B(n634), .C(n597), .Z(n595) );
  CENX1 U1338 ( .A(n602), .B(n63), .Z(SUM[12]) );
  CND2XL U1339 ( .A(n729), .B(n601), .Z(n63) );
  COND1XL U1340 ( .A(n603), .B(n634), .C(n604), .Z(n602) );
  CENX1 U1341 ( .A(n613), .B(n64), .Z(SUM[11]) );
  CND2XL U1342 ( .A(n730), .B(n612), .Z(n64) );
  COND1XL U1343 ( .A(n614), .B(n634), .C(n615), .Z(n613) );
  CENX1 U1344 ( .A(n620), .B(n65), .Z(SUM[10]) );
  CND2XL U1345 ( .A(n731), .B(n619), .Z(n65) );
  COND1XL U1346 ( .A(n621), .B(n634), .C(n622), .Z(n620) );
  CENX1 U1347 ( .A(n631), .B(n66), .Z(SUM[9]) );
  CND2XL U1348 ( .A(n732), .B(n630), .Z(n66) );
  COND1XL U1349 ( .A(n632), .B(n634), .C(n633), .Z(n631) );
  CEOXL U1350 ( .A(n67), .B(n634), .Z(SUM[8]) );
  CND2XL U1351 ( .A(n733), .B(n633), .Z(n67) );
  CND2XL U1352 ( .A(n735), .B(n648), .Z(n69) );
  CANR1XL U1353 ( .A(n650), .B(n663), .C(n651), .Z(n649) );
  CND2XL U1354 ( .A(n736), .B(n657), .Z(n70) );
  CANR1XL U1355 ( .A(n737), .B(n663), .C(n660), .Z(n658) );
  CND2XL U1356 ( .A(n734), .B(n641), .Z(n68) );
  CANR1XL U1357 ( .A(n663), .B(n643), .C(n644), .Z(n642) );
  CENX1 U1358 ( .A(n669), .B(n72), .Z(SUM[3]) );
  CND2XL U1359 ( .A(n738), .B(n668), .Z(n72) );
  COND1XL U1360 ( .A(n670), .B(n672), .C(n671), .Z(n669) );
  CENX1 U1361 ( .A(n663), .B(n71), .Z(SUM[4]) );
  CND2XL U1362 ( .A(n737), .B(n662), .Z(n71) );
  CEOXL U1363 ( .A(n73), .B(n672), .Z(SUM[2]) );
  CND2XL U1364 ( .A(n739), .B(n671), .Z(n73) );
  CEOXL U1365 ( .A(n677), .B(n74), .Z(SUM[1]) );
  CND2XL U1366 ( .A(n740), .B(n675), .Z(n74) );
  COR2X1 U1367 ( .A(B[63]), .B(A[63]), .Z(n941) );
  CANR1X2 U1368 ( .A(n337), .B(n252), .C(n253), .Z(n5) );
  CIVX2 U1369 ( .A(n101), .Z(n99) );
  CIVX2 U1370 ( .A(n100), .Z(n98) );
  CIVX2 U1371 ( .A(n90), .Z(n88) );
  CIVX2 U1372 ( .A(n674), .Z(n740) );
  CIVX2 U1373 ( .A(n670), .Z(n739) );
  CIVX2 U1374 ( .A(n667), .Z(n738) );
  CIVX2 U1375 ( .A(n656), .Z(n736) );
  CIVX2 U1376 ( .A(n645), .Z(n735) );
  CIVX2 U1377 ( .A(n640), .Z(n734) );
  CIVX2 U1378 ( .A(n632), .Z(n733) );
  CIVX2 U1379 ( .A(n629), .Z(n732) );
  CIVX2 U1380 ( .A(n611), .Z(n730) );
  CIVX2 U1381 ( .A(n593), .Z(n728) );
  CIVX2 U1382 ( .A(n580), .Z(n727) );
  CIVX2 U1383 ( .A(n573), .Z(n726) );
  CIVX2 U1384 ( .A(n558), .Z(n724) );
  CIVX2 U1385 ( .A(n547), .Z(n723) );
  CIVX2 U1386 ( .A(n542), .Z(n722) );
  CIVX2 U1387 ( .A(n527), .Z(n721) );
  CIVX2 U1388 ( .A(n522), .Z(n720) );
  CIVX2 U1389 ( .A(n509), .Z(n719) );
  CIVX2 U1390 ( .A(n504), .Z(n718) );
  CIVX2 U1391 ( .A(n489), .Z(n717) );
  CIVX2 U1392 ( .A(n484), .Z(n716) );
  CIVX2 U1393 ( .A(n462), .Z(n714) );
  CIVX2 U1394 ( .A(n440), .Z(n712) );
  CIVX2 U1395 ( .A(n425), .Z(n711) );
  CIVX2 U1396 ( .A(n416), .Z(n710) );
  CIVX2 U1397 ( .A(n400), .Z(n708) );
  CIVX2 U1398 ( .A(n389), .Z(n707) );
  CIVX2 U1399 ( .A(n384), .Z(n706) );
  CIVX2 U1400 ( .A(n369), .Z(n705) );
  CIVX2 U1401 ( .A(n364), .Z(n704) );
  CIVX2 U1402 ( .A(n351), .Z(n703) );
  CIVX2 U1403 ( .A(n346), .Z(n702) );
  CIVX2 U1404 ( .A(n331), .Z(n701) );
  CIVX2 U1405 ( .A(n326), .Z(n700) );
  CIVX2 U1406 ( .A(n304), .Z(n698) );
  CIVX2 U1407 ( .A(n282), .Z(n696) );
  CIVX2 U1408 ( .A(n267), .Z(n695) );
  CIVX2 U1409 ( .A(n258), .Z(n694) );
  CIVX2 U1410 ( .A(n243), .Z(n693) );
  CIVX2 U1411 ( .A(n238), .Z(n692) );
  CIVX2 U1412 ( .A(n216), .Z(n690) );
  CIVX2 U1413 ( .A(n194), .Z(n688) );
  CIVX2 U1414 ( .A(n179), .Z(n687) );
  CIVX2 U1415 ( .A(n170), .Z(n686) );
  CIVX2 U1416 ( .A(n148), .Z(n684) );
  CIVX2 U1417 ( .A(n133), .Z(n683) );
  CIVX2 U1418 ( .A(n124), .Z(n682) );
  CIVX2 U1419 ( .A(n111), .Z(n681) );
  CIVX2 U1420 ( .A(n102), .Z(n680) );
  CIVX2 U1421 ( .A(n673), .Z(n672) );
  CIVX2 U1422 ( .A(n664), .Z(n663) );
  CIVX2 U1423 ( .A(n662), .Z(n660) );
  CIVX2 U1424 ( .A(n661), .Z(n737) );
  CIVX2 U1425 ( .A(n651), .Z(n653) );
  CIVX2 U1426 ( .A(n635), .Z(n634) );
  CIVX2 U1427 ( .A(n619), .Z(n617) );
  CIVX2 U1428 ( .A(n618), .Z(n731) );
  CIVX2 U1429 ( .A(n603), .Z(n605) );
  CIVX2 U1430 ( .A(n601), .Z(n599) );
  CIVX2 U1431 ( .A(n600), .Z(n729) );
  CIVX2 U1432 ( .A(n588), .Z(n590) );
  CIVX2 U1433 ( .A(n564), .Z(n562) );
  CIVX2 U1434 ( .A(n563), .Z(n725) );
  CIVX2 U1435 ( .A(n553), .Z(n555) );
  CIVX2 U1436 ( .A(n535), .Z(n537) );
  CIVX2 U1437 ( .A(n534), .Z(n536) );
  CIVX2 U1438 ( .A(n517), .Z(n515) );
  CIVX2 U1439 ( .A(n516), .Z(n514) );
  CIVX2 U1440 ( .A(n495), .Z(n497) );
  CIVX2 U1441 ( .A(n494), .Z(n496) );
  CIVX2 U1442 ( .A(n479), .Z(n477) );
  CIVX2 U1443 ( .A(n478), .Z(n476) );
  CIVX2 U1444 ( .A(n472), .Z(n470) );
  CIVX2 U1445 ( .A(n471), .Z(n715) );
  CIVX2 U1446 ( .A(n455), .Z(n457) );
  CIVX2 U1447 ( .A(n454), .Z(n456) );
  CIVX2 U1448 ( .A(n450), .Z(n448) );
  CIVX2 U1449 ( .A(n449), .Z(n713) );
  CIVX2 U1450 ( .A(n435), .Z(n437) );
  CIVX2 U1451 ( .A(n406), .Z(n404) );
  CIVX2 U1452 ( .A(n405), .Z(n709) );
  CIVX2 U1453 ( .A(n395), .Z(n397) );
  CIVX2 U1454 ( .A(n377), .Z(n379) );
  CIVX2 U1455 ( .A(n376), .Z(n378) );
  CIVX2 U1456 ( .A(n359), .Z(n357) );
  CIVX2 U1457 ( .A(n358), .Z(n356) );
  CIVX2 U1458 ( .A(n337), .Z(n339) );
  CIVX2 U1459 ( .A(n336), .Z(n338) );
  CIVX2 U1460 ( .A(n321), .Z(n319) );
  CIVX2 U1461 ( .A(n320), .Z(n318) );
  CIVX2 U1462 ( .A(n314), .Z(n312) );
  CIVX2 U1463 ( .A(n313), .Z(n699) );
  CIVX2 U1464 ( .A(n297), .Z(n299) );
  CIVX2 U1465 ( .A(n296), .Z(n298) );
  CIVX2 U1466 ( .A(n292), .Z(n290) );
  CIVX2 U1467 ( .A(n291), .Z(n697) );
  CIVX2 U1468 ( .A(n277), .Z(n279) );
  CIVX2 U1469 ( .A(n5), .Z(n249) );
  CIVX2 U1470 ( .A(n7), .Z(n248) );
  CIVX2 U1471 ( .A(n233), .Z(n231) );
  CIVX2 U1472 ( .A(n232), .Z(n230) );
  CIVX2 U1473 ( .A(n226), .Z(n224) );
  CIVX2 U1474 ( .A(n225), .Z(n691) );
  CIVX2 U1475 ( .A(n209), .Z(n211) );
  CIVX2 U1476 ( .A(n208), .Z(n210) );
  CIVX2 U1477 ( .A(n204), .Z(n202) );
  CIVX2 U1478 ( .A(n203), .Z(n689) );
  CIVX2 U1479 ( .A(n189), .Z(n191) );
  CIVX2 U1480 ( .A(n8), .Z(n163) );
  CIVX2 U1481 ( .A(n9), .Z(n162) );
  CIVX2 U1482 ( .A(n158), .Z(n156) );
  CIVX2 U1483 ( .A(n157), .Z(n685) );
  CIVX2 U1484 ( .A(n143), .Z(n145) );
  CIVX2 U1485 ( .A(n10), .Z(n121) );
  CIVX2 U1486 ( .A(n11), .Z(n120) );
  CIVX2 U1487 ( .A(n75), .Z(SUM[0]) );
endmodule


module sfilt_DW01_add_3 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n212, n213, n214, n215,
         n216, n217, n218, n219, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n256, n257, n258, n259, n260, n261, n262,
         n263, n265, n266, n267;
  assign n10 = A[59];
  assign n15 = A[58];
  assign n18 = A[57];
  assign n22 = A[56];
  assign n25 = A[55];
  assign n33 = A[54];
  assign n36 = A[53];
  assign n40 = A[52];
  assign n43 = A[51];
  assign n49 = A[50];
  assign n52 = A[49];
  assign n56 = A[48];
  assign n60 = A[47];
  assign n69 = A[46];
  assign n72 = A[45];
  assign n76 = A[44];
  assign n79 = A[43];
  assign n85 = A[42];
  assign n88 = A[41];
  assign n92 = A[40];
  assign n96 = A[39];
  assign n103 = A[38];
  assign n106 = A[37];
  assign n110 = A[36];
  assign n113 = A[35];
  assign n119 = A[34];
  assign n123 = A[33];
  assign n128 = A[32];
  assign n131 = A[31];
  assign n139 = A[30];
  assign n142 = A[29];
  assign n146 = A[28];
  assign n149 = A[27];
  assign n155 = A[26];
  assign n158 = A[25];
  assign n162 = A[24];
  assign n166 = A[23];
  assign n173 = A[22];
  assign n176 = A[21];
  assign n180 = A[20];
  assign n183 = A[19];
  assign n190 = A[18];
  assign n193 = A[17];
  assign n197 = A[16];
  assign n201 = A[15];
  assign n208 = A[14];
  assign n212 = A[13];
  assign n217 = A[12];
  assign n221 = A[11];
  assign n227 = A[10];
  assign n231 = A[9];
  assign n236 = A[8];
  assign n239 = A[7];
  assign n245 = A[6];
  assign n248 = A[5];
  assign n252 = A[4];
  assign n256 = A[3];
  assign n261 = A[2];
  assign n265 = A[1];

  CHA1X1 U2 ( .A(A[62]), .B(n4), .CO(n3), .S(SUM[62]) );
  CHA1X1 U3 ( .A(A[61]), .B(n5), .CO(n4), .S(SUM[61]) );
  CHA1X1 U4 ( .A(A[60]), .B(n6), .CO(n5), .S(SUM[60]) );
  CIVX1 U333 ( .A(n204), .Z(n203) );
  CIVXL U334 ( .A(n212), .Z(n213) );
  CEOXL U335 ( .A(n156), .B(n157), .Z(SUM[26]) );
  CIVXL U336 ( .A(n208), .Z(n209) );
  CIVXL U337 ( .A(n134), .Z(n133) );
  CIVXL U338 ( .A(n63), .Z(n62) );
  CIVXL U339 ( .A(n99), .Z(n98) );
  CIVXL U340 ( .A(n28), .Z(n27) );
  CIVXL U341 ( .A(n46), .Z(n45) );
  CIVXL U342 ( .A(n82), .Z(n81) );
  CIVXL U343 ( .A(n116), .Z(n115) );
  CIVXL U344 ( .A(n152), .Z(n151) );
  CNR2XL U345 ( .A(n203), .B(n196), .Z(n195) );
  CNR2XL U346 ( .A(n258), .B(n251), .Z(n250) );
  CNR2XL U347 ( .A(n203), .B(n170), .Z(n169) );
  CNR2XL U348 ( .A(n62), .B(n61), .Z(n58) );
  CNR2XL U349 ( .A(n98), .B(n97), .Z(n94) );
  CNR2XL U350 ( .A(n168), .B(n167), .Z(n164) );
  CNR2XL U351 ( .A(n1), .B(n266), .Z(n263) );
  CND2XL U352 ( .A(n133), .B(n126), .Z(n125) );
  CND2XL U353 ( .A(n241), .B(n225), .Z(n224) );
  CIVXL U354 ( .A(n242), .Z(n241) );
  CIVXL U355 ( .A(n259), .Z(n258) );
  CND2XL U356 ( .A(n133), .B(n131), .Z(n130) );
  CND2XL U357 ( .A(n186), .B(n183), .Z(n182) );
  CND2XL U358 ( .A(n195), .B(n193), .Z(n192) );
  CND2XL U359 ( .A(n241), .B(n239), .Z(n238) );
  CND2XL U360 ( .A(n250), .B(n248), .Z(n247) );
  CIVX1 U361 ( .A(n201), .Z(n202) );
  CIVXL U362 ( .A(n231), .Z(n232) );
  CIVXL U363 ( .A(n256), .Z(n257) );
  CIVXL U364 ( .A(n265), .Z(n266) );
  CIVXL U365 ( .A(n221), .Z(n222) );
  CEOXL U366 ( .A(n61), .B(n62), .Z(SUM[47]) );
  CEOXL U367 ( .A(n97), .B(n98), .Z(SUM[39]) );
  CEOXL U368 ( .A(n167), .B(n168), .Z(SUM[23]) );
  CEOXL U369 ( .A(n184), .B(n185), .Z(SUM[19]) );
  CEOXL U370 ( .A(n202), .B(n203), .Z(SUM[15]) );
  CEOXL U371 ( .A(n1), .B(n266), .Z(SUM[1]) );
  CNR2XL U372 ( .A(A[0]), .B(B[0]), .Z(n267) );
  CND2IXL U373 ( .B(n267), .A(n1), .Z(n2) );
  CIVXL U374 ( .A(n236), .Z(n237) );
  CIVXL U375 ( .A(n245), .Z(n246) );
  CIVX1 U376 ( .A(n88), .Z(n89) );
  CIVX1 U377 ( .A(n131), .Z(n132) );
  CIVX1 U378 ( .A(n158), .Z(n159) );
  CIVXL U379 ( .A(n193), .Z(n194) );
  CIVX1 U380 ( .A(n197), .Z(n198) );
  CIVXL U381 ( .A(n217), .Z(n218) );
  CIVXL U382 ( .A(n227), .Z(n228) );
  CIVXL U383 ( .A(n239), .Z(n240) );
  CIVXL U384 ( .A(n248), .Z(n249) );
  CIVXL U385 ( .A(n252), .Z(n253) );
  CIVXL U386 ( .A(n261), .Z(n262) );
  CNR2X1 U387 ( .A(n28), .B(n21), .Z(n20) );
  CNR2X1 U388 ( .A(n46), .B(n39), .Z(n38) );
  CNR2X1 U389 ( .A(n62), .B(n55), .Z(n54) );
  CNR2X1 U390 ( .A(n82), .B(n75), .Z(n74) );
  CNR2X1 U391 ( .A(n98), .B(n91), .Z(n90) );
  CNR2X1 U392 ( .A(n116), .B(n109), .Z(n108) );
  CNR2X1 U393 ( .A(n152), .B(n145), .Z(n144) );
  CNR2X1 U394 ( .A(n168), .B(n161), .Z(n160) );
  CNR2X1 U395 ( .A(n185), .B(n179), .Z(n178) );
  CNR2X1 U396 ( .A(n134), .B(n64), .Z(n63) );
  CNR2X1 U397 ( .A(n125), .B(n124), .Z(n121) );
  CNR2X1 U398 ( .A(n203), .B(n202), .Z(n199) );
  CNR2X1 U399 ( .A(n214), .B(n213), .Z(n210) );
  CNR2X1 U400 ( .A(n224), .B(n222), .Z(n219) );
  CNR2X1 U401 ( .A(n233), .B(n232), .Z(n229) );
  CNR2X1 U402 ( .A(n258), .B(n257), .Z(n254) );
  CNR2X1 U403 ( .A(n134), .B(n100), .Z(n99) );
  CNR2X1 U404 ( .A(n203), .B(n187), .Z(n186) );
  CND2X1 U405 ( .A(n135), .B(n204), .Z(n134) );
  CNR2X1 U406 ( .A(n170), .B(n136), .Z(n135) );
  CND2X1 U407 ( .A(n153), .B(n137), .Z(n136) );
  CNR2X1 U408 ( .A(n145), .B(n138), .Z(n137) );
  CND2X1 U409 ( .A(n223), .B(n215), .Z(n214) );
  CND2X1 U410 ( .A(n241), .B(n234), .Z(n233) );
  CND2X1 U411 ( .A(n63), .B(n29), .Z(n28) );
  CND2X1 U412 ( .A(n63), .B(n47), .Z(n46) );
  CND2X1 U413 ( .A(n99), .B(n83), .Z(n82) );
  CND2X1 U414 ( .A(n133), .B(n117), .Z(n116) );
  CND2X1 U415 ( .A(n169), .B(n153), .Z(n152) );
  CND2X1 U416 ( .A(n27), .B(n13), .Z(n12) );
  CND2X1 U417 ( .A(A[0]), .B(B[0]), .Z(n1) );
  CNR2X1 U418 ( .A(n21), .B(n14), .Z(n13) );
  CND2X1 U419 ( .A(n18), .B(n15), .Z(n14) );
  CNR2X1 U420 ( .A(n127), .B(n118), .Z(n117) );
  CND2X1 U421 ( .A(n123), .B(n119), .Z(n118) );
  CNR2X1 U422 ( .A(n235), .B(n226), .Z(n225) );
  CND2X1 U423 ( .A(n231), .B(n227), .Z(n226) );
  CNR2X1 U424 ( .A(n260), .B(n1), .Z(n259) );
  CND2X1 U425 ( .A(n265), .B(n261), .Z(n260) );
  CNR2X1 U426 ( .A(n205), .B(n242), .Z(n204) );
  CND2X1 U427 ( .A(n225), .B(n206), .Z(n205) );
  CNR2X1 U428 ( .A(n216), .B(n207), .Z(n206) );
  CND2X1 U429 ( .A(n212), .B(n208), .Z(n207) );
  CNR2X1 U430 ( .A(n100), .B(n66), .Z(n65) );
  CND2X1 U431 ( .A(n83), .B(n67), .Z(n66) );
  CNR2X1 U432 ( .A(n75), .B(n68), .Z(n67) );
  CND2X1 U433 ( .A(n72), .B(n69), .Z(n68) );
  CENX1 U434 ( .A(n250), .B(n249), .Z(SUM[5]) );
  CEOX1 U435 ( .A(n11), .B(n12), .Z(SUM[59]) );
  CEOX1 U436 ( .A(n23), .B(n24), .Z(SUM[56]) );
  CEOX1 U437 ( .A(n41), .B(n42), .Z(SUM[52]) );
  CEOX1 U438 ( .A(n50), .B(n51), .Z(SUM[50]) );
  CEOX1 U439 ( .A(n77), .B(n78), .Z(SUM[44]) );
  CEOX1 U440 ( .A(n86), .B(n87), .Z(SUM[42]) );
  CEOX1 U441 ( .A(n111), .B(n112), .Z(SUM[36]) );
  CEOX1 U442 ( .A(n124), .B(n125), .Z(SUM[33]) );
  CEOX1 U443 ( .A(n129), .B(n130), .Z(SUM[32]) );
  CEOX1 U444 ( .A(n147), .B(n148), .Z(SUM[28]) );
  CEOX1 U445 ( .A(n174), .B(n175), .Z(SUM[22]) );
  CEOX1 U446 ( .A(n232), .B(n233), .Z(SUM[9]) );
  CEOX1 U447 ( .A(n246), .B(n247), .Z(SUM[6]) );
  CEOX1 U448 ( .A(A[63]), .B(n3), .Z(SUM[63]) );
  CND2X1 U449 ( .A(n25), .B(n22), .Z(n21) );
  CND2X1 U450 ( .A(n60), .B(n56), .Z(n55) );
  CND2X1 U451 ( .A(n43), .B(n40), .Z(n39) );
  CND2X1 U452 ( .A(n113), .B(n110), .Z(n109) );
  CND2X1 U453 ( .A(n96), .B(n92), .Z(n91) );
  CND2X1 U454 ( .A(n79), .B(n76), .Z(n75) );
  CND2X1 U455 ( .A(n256), .B(n252), .Z(n251) );
  CND2X1 U456 ( .A(n201), .B(n197), .Z(n196) );
  CND2X1 U457 ( .A(n183), .B(n180), .Z(n179) );
  CND2X1 U458 ( .A(n166), .B(n162), .Z(n161) );
  CND2X1 U459 ( .A(n149), .B(n146), .Z(n145) );
  CND2X1 U460 ( .A(n117), .B(n101), .Z(n100) );
  CNR2X1 U461 ( .A(n109), .B(n102), .Z(n101) );
  CND2X1 U462 ( .A(n106), .B(n103), .Z(n102) );
  CND2X1 U463 ( .A(n188), .B(n171), .Z(n170) );
  CNR2X1 U464 ( .A(n179), .B(n172), .Z(n171) );
  CND2X1 U465 ( .A(n176), .B(n173), .Z(n172) );
  CND2X1 U466 ( .A(n243), .B(n259), .Z(n242) );
  CNR2X1 U467 ( .A(n251), .B(n244), .Z(n243) );
  CND2X1 U468 ( .A(n248), .B(n245), .Z(n244) );
  CND2X1 U469 ( .A(n131), .B(n128), .Z(n127) );
  CND2X1 U470 ( .A(n239), .B(n236), .Z(n235) );
  CND2X1 U471 ( .A(n221), .B(n217), .Z(n216) );
  CND2X1 U472 ( .A(n47), .B(n31), .Z(n30) );
  CNR2X1 U473 ( .A(n39), .B(n32), .Z(n31) );
  CND2X1 U474 ( .A(n36), .B(n33), .Z(n32) );
  CND2X1 U475 ( .A(n20), .B(n18), .Z(n17) );
  CND2X1 U476 ( .A(n27), .B(n25), .Z(n24) );
  CND2X1 U477 ( .A(n38), .B(n36), .Z(n35) );
  CND2X1 U478 ( .A(n45), .B(n43), .Z(n42) );
  CND2X1 U479 ( .A(n54), .B(n52), .Z(n51) );
  CND2X1 U480 ( .A(n74), .B(n72), .Z(n71) );
  CND2X1 U481 ( .A(n81), .B(n79), .Z(n78) );
  CND2X1 U482 ( .A(n90), .B(n88), .Z(n87) );
  CND2X1 U483 ( .A(n108), .B(n106), .Z(n105) );
  CND2X1 U484 ( .A(n115), .B(n113), .Z(n112) );
  CND2X1 U485 ( .A(n144), .B(n142), .Z(n141) );
  CND2X1 U486 ( .A(n151), .B(n149), .Z(n148) );
  CND2X1 U487 ( .A(n160), .B(n158), .Z(n157) );
  CND2X1 U488 ( .A(n178), .B(n176), .Z(n175) );
  CNR2X1 U489 ( .A(n7), .B(n134), .Z(n6) );
  CND2X1 U490 ( .A(n65), .B(n8), .Z(n7) );
  CNR2X1 U491 ( .A(n30), .B(n9), .Z(n8) );
  CEOX1 U492 ( .A(n16), .B(n17), .Z(SUM[58]) );
  CENX1 U493 ( .A(n20), .B(n19), .Z(SUM[57]) );
  CENX1 U494 ( .A(n27), .B(n26), .Z(SUM[55]) );
  CEOX1 U495 ( .A(n34), .B(n35), .Z(SUM[54]) );
  CENX1 U496 ( .A(n38), .B(n37), .Z(SUM[53]) );
  CENX1 U497 ( .A(n45), .B(n44), .Z(SUM[51]) );
  CENX1 U498 ( .A(n54), .B(n53), .Z(SUM[49]) );
  CENX1 U499 ( .A(n58), .B(n57), .Z(SUM[48]) );
  CEOX1 U500 ( .A(n70), .B(n71), .Z(SUM[46]) );
  CENX1 U501 ( .A(n74), .B(n73), .Z(SUM[45]) );
  CENX1 U502 ( .A(n81), .B(n80), .Z(SUM[43]) );
  CENX1 U503 ( .A(n90), .B(n89), .Z(SUM[41]) );
  CENX1 U504 ( .A(n94), .B(n93), .Z(SUM[40]) );
  CEOX1 U505 ( .A(n104), .B(n105), .Z(SUM[38]) );
  CENX1 U506 ( .A(n108), .B(n107), .Z(SUM[37]) );
  CENX1 U507 ( .A(n115), .B(n114), .Z(SUM[35]) );
  CENX1 U508 ( .A(n121), .B(n120), .Z(SUM[34]) );
  CENX1 U509 ( .A(n133), .B(n132), .Z(SUM[31]) );
  CEOX1 U510 ( .A(n140), .B(n141), .Z(SUM[30]) );
  CENX1 U511 ( .A(n144), .B(n143), .Z(SUM[29]) );
  CENX1 U512 ( .A(n151), .B(n150), .Z(SUM[27]) );
  CENX1 U513 ( .A(n160), .B(n159), .Z(SUM[25]) );
  CENX1 U514 ( .A(n164), .B(n163), .Z(SUM[24]) );
  CENX1 U515 ( .A(n178), .B(n177), .Z(SUM[21]) );
  CEOX1 U516 ( .A(n181), .B(n182), .Z(SUM[20]) );
  CEOX1 U517 ( .A(n191), .B(n192), .Z(SUM[18]) );
  CENX1 U518 ( .A(n195), .B(n194), .Z(SUM[17]) );
  CENX1 U519 ( .A(n199), .B(n198), .Z(SUM[16]) );
  CENX1 U520 ( .A(n210), .B(n209), .Z(SUM[14]) );
  CEOX1 U521 ( .A(n213), .B(n214), .Z(SUM[13]) );
  CENX1 U522 ( .A(n219), .B(n218), .Z(SUM[12]) );
  CENX1 U523 ( .A(n223), .B(n222), .Z(SUM[11]) );
  CENX1 U524 ( .A(n229), .B(n228), .Z(SUM[10]) );
  CEOX1 U525 ( .A(n237), .B(n238), .Z(SUM[8]) );
  CENX1 U526 ( .A(n241), .B(n240), .Z(SUM[7]) );
  CENX1 U527 ( .A(n254), .B(n253), .Z(SUM[4]) );
  CEOX1 U528 ( .A(n257), .B(n258), .Z(SUM[3]) );
  CENX1 U529 ( .A(n263), .B(n262), .Z(SUM[2]) );
  CND2X1 U530 ( .A(n142), .B(n139), .Z(n138) );
  CNR2X1 U531 ( .A(n55), .B(n48), .Z(n47) );
  CND2X1 U532 ( .A(n52), .B(n49), .Z(n48) );
  CNR2X1 U533 ( .A(n91), .B(n84), .Z(n83) );
  CND2X1 U534 ( .A(n88), .B(n85), .Z(n84) );
  CNR2X1 U535 ( .A(n196), .B(n189), .Z(n188) );
  CND2X1 U536 ( .A(n193), .B(n190), .Z(n189) );
  CNR2X1 U537 ( .A(n161), .B(n154), .Z(n153) );
  CND2X1 U538 ( .A(n158), .B(n155), .Z(n154) );
  CND2X1 U539 ( .A(n13), .B(n10), .Z(n9) );
  CIVX2 U540 ( .A(n96), .Z(n97) );
  CIVX2 U541 ( .A(n92), .Z(n93) );
  CIVX2 U542 ( .A(n85), .Z(n86) );
  CIVX2 U543 ( .A(n79), .Z(n80) );
  CIVX2 U544 ( .A(n76), .Z(n77) );
  CIVX2 U545 ( .A(n72), .Z(n73) );
  CIVX2 U546 ( .A(n69), .Z(n70) );
  CIVX2 U547 ( .A(n65), .Z(n64) );
  CIVX2 U548 ( .A(n60), .Z(n61) );
  CIVX2 U549 ( .A(n56), .Z(n57) );
  CIVX2 U550 ( .A(n52), .Z(n53) );
  CIVX2 U551 ( .A(n49), .Z(n50) );
  CIVX2 U552 ( .A(n43), .Z(n44) );
  CIVX2 U553 ( .A(n40), .Z(n41) );
  CIVX2 U554 ( .A(n36), .Z(n37) );
  CIVX2 U555 ( .A(n33), .Z(n34) );
  CIVX2 U556 ( .A(n30), .Z(n29) );
  CIVX2 U557 ( .A(n25), .Z(n26) );
  CIVX2 U558 ( .A(n235), .Z(n234) );
  CIVX2 U559 ( .A(n22), .Z(n23) );
  CIVX2 U560 ( .A(n224), .Z(n223) );
  CIVX2 U561 ( .A(n216), .Z(n215) );
  CIVX2 U562 ( .A(n190), .Z(n191) );
  CIVX2 U563 ( .A(n18), .Z(n19) );
  CIVX2 U564 ( .A(n188), .Z(n187) );
  CIVX2 U565 ( .A(n186), .Z(n185) );
  CIVX2 U566 ( .A(n183), .Z(n184) );
  CIVX2 U567 ( .A(n180), .Z(n181) );
  CIVX2 U568 ( .A(n176), .Z(n177) );
  CIVX2 U569 ( .A(n173), .Z(n174) );
  CIVX2 U570 ( .A(n169), .Z(n168) );
  CIVX2 U571 ( .A(n166), .Z(n167) );
  CIVX2 U572 ( .A(n162), .Z(n163) );
  CIVX2 U573 ( .A(n15), .Z(n16) );
  CIVX2 U574 ( .A(n155), .Z(n156) );
  CIVX2 U575 ( .A(n149), .Z(n150) );
  CIVX2 U576 ( .A(n146), .Z(n147) );
  CIVX2 U577 ( .A(n142), .Z(n143) );
  CIVX2 U578 ( .A(n139), .Z(n140) );
  CIVX2 U579 ( .A(n128), .Z(n129) );
  CIVX2 U580 ( .A(n127), .Z(n126) );
  CIVX2 U581 ( .A(n123), .Z(n124) );
  CIVX2 U582 ( .A(n119), .Z(n120) );
  CIVX2 U583 ( .A(n113), .Z(n114) );
  CIVX2 U584 ( .A(n110), .Z(n111) );
  CIVX2 U585 ( .A(n10), .Z(n11) );
  CIVX2 U586 ( .A(n106), .Z(n107) );
  CIVX2 U587 ( .A(n103), .Z(n104) );
  CIVX2 U588 ( .A(n2), .Z(SUM[0]) );
endmodule


module sfilt_DW_mult_tc_1 ( a, b, product );
  input [31:0] a;
  input [31:0] b;
  output [63:0] product;
  wire   n3, n6, n12, n18, n21, n24, n27, n30, n33, n36, n39, n42, n45, n48,
         n51, n54, n57, n60, n63, n66, n72, n75, n78, n81, n84, n87, n90, n93,
         n96, n99, n102, n108, n111, n117, n120, n126, n129, n136, n141, n144,
         n145, n149, n150, n151, n153, n154, n155, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n173, n174, n175, n176, n177, n178, n179, n184, n185, n186, n187,
         n188, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n212,
         n213, n214, n216, n218, n219, n220, n221, n222, n223, n224, n225,
         n227, n229, n230, n231, n232, n233, n236, n241, n242, n256, n257,
         n258, n259, n267, n268, n269, n274, n279, n280, n281, n282, n283,
         n286, n291, n292, n304, n305, n306, n317, n318, n319, n320, n324,
         n327, n328, n329, n330, n331, n332, n333, n334, n340, n342, n343,
         n344, n345, n349, n351, n352, n353, n355, n356, n371, n372, n373,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n393,
         n394, n395, n396, n404, n405, n406, n408, n409, n411, n412, n413,
         n414, n415, n416, n418, n424, n425, n426, n427, n428, n432, n434,
         n435, n438, n441, n444, n445, n448, n449, n450, n451, n452, n456,
         n458, n459, n460, n461, n463, n467, n468, n469, n470, n471, n472,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n494, n495, n496, n497, n498, n499, n501, n504,
         n505, n506, n507, n508, n510, n511, n512, n513, n514, n516, n517,
         n520, n524, n525, n526, n528, n529, n530, n531, n532, n533, n534,
         n535, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n559, n560, n561, n562, n564,
         n567, n568, n569, n571, n572, n573, n575, n576, n577, n578, n579,
         n583, n584, n585, n586, n590, n591, n592, n593, n594, n595, n596,
         n597, n601, n602, n603, n604, n605, n606, n608, n613, n614, n616,
         n618, n619, n620, n621, n622, n623, n624, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n639, n641, n642,
         n643, n644, n646, n649, n650, n651, n652, n654, n656, n657, n658,
         n659, n660, n661, n662, n664, n665, n666, n667, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n681, n683, n684,
         n686, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n704, n706, n707, n708, n709, n710,
         n712, n714, n718, n720, n721, n722, n723, n724, n726, n728, n729,
         n730, n731, n741, n748, n749, n751, n753, n754, n755, n756, n757,
         n758, n760, n761, n762, n764, n765, n766, n767, n768, n769, n770,
         n772, n773, n774, n776, n778, n779, n780, n781, n784, n785, n786,
         n788, n791, n793, n794, n795, n796, n797, n800, n803, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n828, n829, n830, n831,
         n832, n833, n835, n838, n839, n840, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n896, n897, n898, n900, n901, n902, n903,
         n904, n905, n910, n911, n914, n915, n918, n919, n920, n921, n922,
         n923, n930, n931, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n965, n966,
         n967, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1842, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1872, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1932, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2314, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         net18489, net18487, net18483, net18495, net18521, net18519, net18517,
         net18515, net18549, net18547, net18561, net18555, net18979, net19062,
         net19068, net19081, net19178, net19189, net19193, net19192, net19191,
         net19216, net19215, net19213, net19268, net19281, net19286, net19302,
         net19309, net19314, net20818, net20981, net20990, net20996, net21177,
         net21206, net21250, net21249, net21248, net21297, net21313, net21312,
         net21311, net21320, net21337, net21344, net21353, net21352, net21375,
         net21389, net21419, net21434, net21433, net21438, net21512, net21591,
         net21590, net21622, net21684, net21683, net21696, net21693, net21725,
         net21744, net21791, net21802, net21801, net21836, net21835, net21846,
         net21859, net21858, net21882, net21892, net21896, net21910, net21909,
         net21948, net21983, net22007, net22006, net22013, net22050, net22097,
         net22186, net22190, net22220, net22242, net22241, net22248, net22262,
         net22304, net22303, net22302, net22301, net22327, net22326, net22344,
         net22351, net22399, net22398, net22439, net22471, net22511, net22590,
         net22599, net22598, net22626, net22642, net22641, n2812, n2270, n2269,
         n410, n403, n359, n747, net20956, n247, n246, n244, n152, n402, n277,
         n275, n272, n266, n265, n261, n745, n744, n417, n399, n397, n392,
         n379, n378, n377, n370, n369, n363, n361, n805, n804, n802, n801,
         n799, n798, n736, n273, n264, n262, n260, n255, n253, n249, n248,
         n1742, n992, n973, n972, n69, n2518, n2517, n1992, n1756, net22004,
         net21472, n929, n925, n924, n907, n906, n971, n970, n969, n968, n964,
         n947, n946, n927, n926, n1933, n1873, n1843, n1815, net22288,
         net22287, net22286, net19171, n933, n932, n928, n917, n916, n913,
         n912, n909, n908, n899, n895, n1931, n1901, n1871, n1841, n1783, n114,
         n738, n307, n297, n296, n295, n156, net22552, n841, n837, n836, n834,
         n827, n826, n366, n364, n362, n360, n354, n323, n740, n739, n316,
         n315, n314, n310, n309, n308, n303, n302, n301, n299, n298, n294,
         n293, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007;
  assign n3 = a[1];
  assign n12 = a[3];
  assign n21 = a[5];
  assign n30 = a[7];
  assign n39 = a[9];
  assign n48 = a[11];
  assign n57 = a[13];
  assign n66 = a[15];
  assign n75 = a[17];
  assign n84 = a[19];
  assign n93 = a[21];
  assign n102 = a[23];
  assign n111 = a[25];
  assign n120 = a[27];
  assign n129 = a[29];
  assign n136 = a[31];
  assign n145 = b[0];
  assign n2780 = b[31];
  assign n2781 = b[30];
  assign n2782 = b[29];
  assign n2783 = b[28];
  assign n2784 = b[27];
  assign n2785 = b[26];
  assign n2786 = b[25];
  assign n2787 = b[24];
  assign n2788 = b[23];
  assign n2789 = b[22];
  assign n2790 = b[21];
  assign n2791 = b[20];
  assign n2792 = b[19];
  assign n2793 = b[18];
  assign n2794 = b[17];
  assign n2795 = b[16];
  assign n2796 = b[15];
  assign n2797 = b[14];
  assign n2798 = b[13];
  assign n2799 = b[12];
  assign n2800 = b[11];
  assign n2801 = b[10];
  assign n2802 = b[9];
  assign n2803 = b[8];
  assign n2804 = b[7];
  assign n2805 = b[6];
  assign n2806 = b[5];
  assign n2807 = b[4];
  assign n2808 = b[3];
  assign n2809 = b[2];
  assign n2810 = b[1];

  COND1X1 U162 ( .A(n220), .B(n3744), .C(n221), .Z(n219) );
  CANR1X1 U168 ( .A(n3223), .B(n236), .C(n227), .Z(n225) );
  CND2X2 U229 ( .A(n283), .B(net20981), .Z(n274) );
  CNR2X2 U243 ( .A(n333), .B(n3910), .Z(n283) );
  COND1X1 U244 ( .A(n3910), .B(n334), .C(n3222), .Z(n286) );
  CNR2X2 U295 ( .A(n835), .B(n844), .Z(n324) );
  CND2X2 U307 ( .A(n3908), .B(n3914), .Z(n333) );
  COND1X1 U328 ( .A(n3238), .B(n3892), .C(net22471), .Z(n352) );
  COND1X1 U350 ( .A(n372), .B(net21389), .C(n373), .Z(n371) );
  COND1X1 U362 ( .A(n381), .B(n3892), .C(n382), .Z(n380) );
  COND1X1 U366 ( .A(n385), .B(n441), .C(n386), .Z(n384) );
  CANR1X1 U368 ( .A(net22590), .B(n387), .C(n388), .Z(n386) );
  COND1X1 U378 ( .A(n394), .B(net21389), .C(n395), .Z(n393) );
  COND1X1 U392 ( .A(n405), .B(n3744), .C(n406), .Z(n404) );
  COND1X1 U402 ( .A(n412), .B(n149), .C(n413), .Z(n411) );
  COND1X1 U406 ( .A(n3335), .B(n441), .C(n3244), .Z(n415) );
  CNR2X2 U417 ( .A(n939), .B(n956), .Z(n424) );
  COND1X1 U420 ( .A(n427), .B(n3892), .C(n428), .Z(n426) );
  COND1X1 U432 ( .A(n3448), .B(n149), .C(n441), .Z(n435) );
  CNR2X2 U447 ( .A(n975), .B(n994), .Z(n448) );
  COND1X1 U450 ( .A(n451), .B(net21389), .C(n452), .Z(n450) );
  COND1X1 U462 ( .A(n3119), .B(n149), .C(net22642), .Z(n459) );
  COND1X1 U476 ( .A(n3902), .B(n3744), .C(n3422), .Z(n470) );
  CNR2X2 U531 ( .A(n1133), .B(n1158), .Z(n511) );
  CNR2X2 U555 ( .A(n1214), .B(n3883), .Z(n529) );
  CNR2X2 U586 ( .A(n1275), .B(n1304), .Z(n551) );
  CNR2X2 U596 ( .A(n3781), .B(n1332), .Z(n556) );
  CNR2X2 U608 ( .A(n1333), .B(n1360), .Z(n567) );
  CNR2X2 U655 ( .A(n1437), .B(n1460), .Z(n602) );
  CNR2X2 U684 ( .A(n1505), .B(n1524), .Z(n622) );
  COND1X1 U767 ( .A(n678), .B(n690), .C(n679), .Z(n677) );
  CFA1X1 U858 ( .A(n800), .B(n1771), .CI(n1741), .CO(n796), .S(n797) );
  CFA1X1 U863 ( .A(n816), .B(n814), .CI(n809), .CO(n806), .S(n807) );
  CFA1X1 U864 ( .A(n1743), .B(n811), .CI(n1804), .CO(n808), .S(n809) );
  CFA1X1 U866 ( .A(n817), .B(n815), .CI(n820), .CO(n812), .S(n813) );
  CFA1X1 U867 ( .A(n1744), .B(n822), .CI(n1834), .CO(n814), .S(n815) );
  CFA1X1 U869 ( .A(n823), .B(n821), .CI(n828), .CO(n818), .S(n819) );
  CFA1X1 U870 ( .A(n825), .B(n830), .CI(n832), .CO(n820), .S(n821) );
  CFA1X1 U871 ( .A(n1745), .B(n1835), .CI(n1775), .CO(n822), .S(n823) );
  CFA1X1 U874 ( .A(n840), .B(n831), .CI(n833), .CO(n828), .S(n829) );
  CFA1X1 U875 ( .A(n1746), .B(n1864), .CI(n1776), .CO(n830), .S(n831) );
  CFA1X1 U876 ( .A(n842), .B(n1836), .CI(n1806), .CO(n832), .S(n833) );
  CFA1X1 U879 ( .A(n1837), .B(n852), .CI(n843), .CO(n838), .S(n839) );
  CFA1X1 U882 ( .A(n849), .B(n847), .CI(n856), .CO(n844), .S(n845) );
  CFA1X1 U883 ( .A(n851), .B(n858), .CI(n853), .CO(n846), .S(n847) );
  CFA1X1 U884 ( .A(n1895), .B(n860), .CI(n862), .CO(n848), .S(n849) );
  CFA1X1 U885 ( .A(n1778), .B(n1838), .CI(n1748), .CO(n850), .S(n851) );
  CFA1X1 U886 ( .A(n864), .B(n1866), .CI(n1807), .CO(n852), .S(n853) );
  CFA1X1 U887 ( .A(n859), .B(n857), .CI(n868), .CO(n854), .S(n855) );
  CFA1X1 U888 ( .A(n861), .B(n870), .CI(n872), .CO(n856), .S(n857) );
  CFA1X1 U889 ( .A(n876), .B(n863), .CI(n874), .CO(n858), .S(n859) );
  CFA1X1 U890 ( .A(n1867), .B(n865), .CI(n1779), .CO(n860), .S(n861) );
  CFA1X1 U891 ( .A(n1808), .B(n1896), .CI(n1749), .CO(n862), .S(n863) );
  CFA1X1 U893 ( .A(n871), .B(n869), .CI(n880), .CO(n866), .S(n867) );
  CFA1X1 U894 ( .A(n884), .B(n882), .CI(n873), .CO(n868), .S(n869) );
  CFA1X1 U895 ( .A(n886), .B(n877), .CI(n875), .CO(n870), .S(n871) );
  CFA1X1 U896 ( .A(n1780), .B(n888), .CI(n1927), .CO(n872), .S(n873) );
  CFA1X1 U897 ( .A(n1839), .B(n1868), .CI(n1750), .CO(n874), .S(n875) );
  CFA1X1 U900 ( .A(n898), .B(n896), .CI(n885), .CO(n880), .S(n881) );
  CFA1X1 U901 ( .A(n900), .B(n889), .CI(n887), .CO(n882), .S(n883) );
  CFA1X1 U902 ( .A(n891), .B(n902), .CI(n904), .CO(n884), .S(n885) );
  CFA1X1 U904 ( .A(n1810), .B(n1928), .CI(n1781), .CO(n888), .S(n889) );
  CFA1X1 U908 ( .A(n905), .B(n914), .CI(n901), .CO(n896), .S(n897) );
  CFA1X1 U910 ( .A(n920), .B(n1958), .CI(n1899), .CO(n900), .S(n901) );
  CFA1X1 U911 ( .A(n1870), .B(n1840), .CI(n1782), .CO(n902), .S(n903) );
  CFA1X1 U912 ( .A(n1752), .B(n1929), .CI(n1811), .CO(n904), .S(n905) );
  CFA1X1 U915 ( .A(n919), .B(n915), .CI(n930), .CO(n910), .S(n911) );
  CFA1X1 U917 ( .A(n3215), .B(n936), .CI(n921), .CO(n914), .S(n915) );
  CFA1X1 U919 ( .A(n1812), .B(n1959), .CI(n1753), .CO(n918), .S(n919) );
  CFA1X1 U925 ( .A(n1990), .B(n950), .CI(n952), .CO(n930), .S(n931) );
  CFA1X1 U928 ( .A(n1754), .B(n1960), .CI(n954), .CO(n936), .S(n937) );
  CFA1X1 U930 ( .A(n945), .B(n960), .CI(n962), .CO(n940), .S(n941) );
  CFA1X1 U932 ( .A(n951), .B(n949), .CI(n953), .CO(n944), .S(n945) );
  CFA1X1 U935 ( .A(n1785), .B(n1902), .CI(n1814), .CO(n950), .S(n951) );
  CFA1X1 U938 ( .A(n961), .B(n959), .CI(n976), .CO(n956), .S(n957) );
  CFA1X1 U940 ( .A(n982), .B(n965), .CI(n967), .CO(n960), .S(n961) );
  CFA1X1 U943 ( .A(n1962), .B(n990), .CI(n2022), .CO(n966), .S(n967) );
  CFA1X1 U949 ( .A(n985), .B(n983), .CI(n1002), .CO(n978), .S(n979) );
  CFA1X1 U950 ( .A(n989), .B(n1004), .CI(n991), .CO(n980), .S(n981) );
  CFA1X1 U951 ( .A(n1008), .B(n987), .CI(n1006), .CO(n982), .S(n983) );
  CFA1X1 U952 ( .A(n993), .B(n1010), .CI(n1012), .CO(n984), .S(n985) );
  CFA1X1 U953 ( .A(n1963), .B(n1934), .CI(n1904), .CO(n986), .S(n987) );
  CFA1X1 U954 ( .A(n1816), .B(n1787), .CI(n1993), .CO(n988), .S(n989) );
  CFA1X1 U955 ( .A(n1844), .B(n2023), .CI(n1757), .CO(n990), .S(n991) );
  CFA1X1 U962 ( .A(n1032), .B(n1030), .CI(n1028), .CO(n1004), .S(n1005) );
  CFA1X1 U963 ( .A(n1994), .B(n2055), .CI(n1964), .CO(n1006), .S(n1007) );
  CFA1X1 U964 ( .A(n1874), .B(n1817), .CI(n1935), .CO(n1008), .S(n1009) );
  CFA1X1 U966 ( .A(n1758), .B(n2024), .CI(n1034), .CO(n1012), .S(n1013) );
  CFA1X1 U970 ( .A(n1048), .B(n1027), .CI(n1046), .CO(n1020), .S(n1021) );
  CFA1X1 U971 ( .A(n1029), .B(n1031), .CI(n1033), .CO(n1022), .S(n1023) );
  CFA1X1 U972 ( .A(n1054), .B(n1052), .CI(n1050), .CO(n1024), .S(n1025) );
  CFA1X1 U973 ( .A(n1965), .B(n1056), .CI(n1035), .CO(n1026), .S(n1027) );
  CFA1X1 U974 ( .A(n1995), .B(n1936), .CI(n1818), .CO(n1028), .S(n1029) );
  CFA1X1 U976 ( .A(n1759), .B(n1875), .CI(n2056), .CO(n1032), .S(n1033) );
  CFA1X1 U980 ( .A(n1047), .B(n1045), .CI(n1066), .CO(n1040), .S(n1041) );
  CFA1X1 U981 ( .A(n1070), .B(n1068), .CI(n1049), .CO(n1042), .S(n1043) );
  CFA1X1 U983 ( .A(n1074), .B(n1051), .CI(n1072), .CO(n1046), .S(n1047) );
  CFA1X1 U984 ( .A(n2088), .B(n1076), .CI(n1078), .CO(n1048), .S(n1049) );
  CFA1X1 U985 ( .A(n1996), .B(n2026), .CI(n1876), .CO(n1050), .S(n1051) );
  CFA1X1 U986 ( .A(n1906), .B(n3497), .CI(n1847), .CO(n1052), .S(n1053) );
  CFA1X1 U987 ( .A(n1937), .B(n1790), .CI(n1819), .CO(n1054), .S(n1055) );
  CFA1X1 U991 ( .A(n1069), .B(n1067), .CI(n1090), .CO(n1062), .S(n1063) );
  CFA1X1 U992 ( .A(n1094), .B(n1071), .CI(n1092), .CO(n1064), .S(n1065) );
  CFA1X1 U993 ( .A(n1079), .B(n1096), .CI(n1073), .CO(n1066), .S(n1067) );
  CFA1X1 U994 ( .A(n1102), .B(n1077), .CI(n1075), .CO(n1068), .S(n1069) );
  CFA1X1 U995 ( .A(n1104), .B(n1100), .CI(n1098), .CO(n1070), .S(n1071) );
  CFA1X1 U996 ( .A(n1967), .B(n1081), .CI(n1848), .CO(n1072), .S(n1073) );
  CFA1X1 U997 ( .A(n1997), .B(n1820), .CI(n1761), .CO(n1074), .S(n1075) );
  CFA1X1 U998 ( .A(n1877), .B(n2027), .CI(n2058), .CO(n1076), .S(n1077) );
  CFA1X1 U999 ( .A(n1907), .B(n2089), .CI(n1791), .CO(n1078), .S(n1079) );
  CFA1X1 U1004 ( .A(n1097), .B(n1095), .CI(n1116), .CO(n1088), .S(n1089) );
  CFA1X1 U1005 ( .A(n1101), .B(n1118), .CI(n1120), .CO(n1090), .S(n1091) );
  CFA1X1 U1006 ( .A(n1099), .B(n1103), .CI(n1105), .CO(n1092), .S(n1093) );
  CFA1X1 U1007 ( .A(n1122), .B(n1126), .CI(n1124), .CO(n1094), .S(n1095) );
  CFA1X1 U1008 ( .A(n2028), .B(n1128), .CI(n2121), .CO(n1096), .S(n1097) );
  CFA1X1 U1009 ( .A(n1998), .B(n1968), .CI(n1130), .CO(n1098), .S(n1099) );
  CFA1X1 U1010 ( .A(n1938), .B(n1878), .CI(n1849), .CO(n1100), .S(n1101) );
  CFA1X1 U1011 ( .A(n1908), .B(n1821), .CI(n1792), .CO(n1102), .S(n1103) );
  CFA1X1 U1012 ( .A(n1762), .B(n2090), .CI(n2059), .CO(n1104), .S(n1105) );
  CFA1X1 U1016 ( .A(n1144), .B(n1142), .CI(n1119), .CO(n1112), .S(n1113) );
  CFA1X1 U1018 ( .A(n1123), .B(n1127), .CI(n1129), .CO(n1116), .S(n1117) );
  CFA1X1 U1019 ( .A(n1150), .B(n1148), .CI(n1152), .CO(n1118), .S(n1119) );
  CFA1X1 U1020 ( .A(n1131), .B(n1154), .CI(n1156), .CO(n1120), .S(n1121) );
  CFA1X1 U1021 ( .A(n2060), .B(n2029), .CI(n1999), .CO(n1122), .S(n1123) );
  CFA1X1 U1022 ( .A(n2091), .B(n1969), .CI(n1850), .CO(n1124), .S(n1125) );
  CFA1X1 U1023 ( .A(n1879), .B(n1822), .CI(n1763), .CO(n1126), .S(n1127) );
  CFA1X1 U1024 ( .A(n1793), .B(n2122), .CI(n1909), .CO(n1128), .S(n1129) );
  CFA1X1 U1029 ( .A(n1147), .B(n1168), .CI(n1145), .CO(n1138), .S(n1139) );
  CFA1X1 U1031 ( .A(n1155), .B(n1149), .CI(n1157), .CO(n1142), .S(n1143) );
  CFA1X1 U1032 ( .A(n1176), .B(n1153), .CI(n1151), .CO(n1144), .S(n1145) );
  CFA1X1 U1033 ( .A(n1178), .B(n1180), .CI(n1182), .CO(n1146), .S(n1147) );
  CFA1X1 U1034 ( .A(n2030), .B(n2154), .CI(n2061), .CO(n1148), .S(n1149) );
  CFA1X1 U1035 ( .A(n1880), .B(n1910), .CI(n2000), .CO(n1150), .S(n1151) );
  CFA1X1 U1037 ( .A(n1794), .B(n1823), .CI(n1939), .CO(n1154), .S(n1155) );
  CFA1X1 U1042 ( .A(n1173), .B(n1171), .CI(n1196), .CO(n1164), .S(n1165) );
  CFA1X1 U1044 ( .A(n1181), .B(n1202), .CI(n1183), .CO(n1168), .S(n1169) );
  CFA1X1 U1045 ( .A(n1208), .B(n1179), .CI(n1177), .CO(n1170), .S(n1171) );
  CFA1X1 U1046 ( .A(n1206), .B(n1204), .CI(n1210), .CO(n1172), .S(n1173) );
  CFA1X1 U1048 ( .A(n2062), .B(n2031), .CI(n2124), .CO(n1176), .S(n1177) );
  CFA1X1 U1050 ( .A(n1911), .B(n1824), .CI(n1795), .CO(n1180), .S(n1181) );
  CFA1X1 U1051 ( .A(n1765), .B(n1940), .CI(n2155), .CO(n1182), .S(n1183) );
  CFA1X1 U1053 ( .A(n1191), .B(n3879), .CI(n1216), .CO(n1186), .S(n1187) );
  CFA1X1 U1054 ( .A(n3196), .B(n1218), .CI(n1193), .CO(n1188), .S(n1189) );
  CFA1X1 U1056 ( .A(n1201), .B(n1224), .CI(n1199), .CO(n1192), .S(n1193) );
  CFA1X1 U1058 ( .A(n1207), .B(n1230), .CI(n1209), .CO(n1196), .S(n1197) );
  CFA1X1 U1060 ( .A(n1236), .B(n1232), .CI(n1234), .CO(n1200), .S(n1201) );
  CFA1X1 U1061 ( .A(n2187), .B(n1238), .CI(n1240), .CO(n1202), .S(n1203) );
  CFA1X1 U1062 ( .A(n1941), .B(n2125), .CI(n2094), .CO(n1204), .S(n1205) );
  CFA1X1 U1063 ( .A(n1825), .B(n2063), .CI(n2032), .CO(n1206), .S(n1207) );
  CFA1X1 U1064 ( .A(n2002), .B(n1912), .CI(n1882), .CO(n1208), .S(n1209) );
  CFA1X1 U1065 ( .A(n1796), .B(n1853), .CI(n1971), .CO(n1210), .S(n1211) );
  CFA1X1 U1066 ( .A(n2156), .B(n1766), .CI(n1242), .CO(n1212), .S(n1213) );
  CFA1X1 U1073 ( .A(n1262), .B(n1233), .CI(n1239), .CO(n1226), .S(n1227) );
  CFA1X1 U1076 ( .A(n2064), .B(n1243), .CI(n2033), .CO(n1232), .S(n1233) );
  CFA1X1 U1077 ( .A(n1972), .B(n2095), .CI(n1883), .CO(n1234), .S(n1235) );
  CFA1X1 U1079 ( .A(n2157), .B(n1797), .CI(n1913), .CO(n1238), .S(n1239) );
  CFA1X1 U1080 ( .A(n1767), .B(n2188), .CI(n1942), .CO(n1240), .S(n1241) );
  CFA1X1 U1087 ( .A(n1267), .B(n1290), .CI(n1263), .CO(n1254), .S(n1255) );
  CFA1X1 U1090 ( .A(n1273), .B(n1296), .CI(n1294), .CO(n1260), .S(n1261) );
  CFA1X1 U1092 ( .A(n2158), .B(n2065), .CI(n2127), .CO(n1264), .S(n1265) );
  CFA1X1 U1098 ( .A(n1279), .B(n1277), .CI(n1306), .CO(n1274), .S(n1275) );
  CFA1X1 U1100 ( .A(n1285), .B(n1310), .CI(n1312), .CO(n1278), .S(n1279) );
  CFA1X1 U1103 ( .A(n1295), .B(n1320), .CI(n1297), .CO(n1284), .S(n1285) );
  CFA1X1 U1104 ( .A(n1301), .B(n1299), .CI(n1293), .CO(n1286), .S(n1287) );
  CFA1X1 U1106 ( .A(n1303), .B(n1328), .CI(n1330), .CO(n1290), .S(n1291) );
  CFA1X1 U1107 ( .A(n1944), .B(n2035), .CI(n1885), .CO(n1292), .S(n1293) );
  CFA1X1 U1109 ( .A(n1915), .B(n2097), .CI(n2128), .CO(n1296), .S(n1297) );
  CFA1X1 U1110 ( .A(n2159), .B(n1974), .CI(n2190), .CO(n1298), .S(n1299) );
  CFA1X1 U1111 ( .A(n2221), .B(n1799), .CI(n2004), .CO(n1300), .S(n1301) );
  CHA1X1 U1112 ( .A(n1724), .B(n1769), .CO(n1302), .S(n1303) );
  CFA1X1 U1117 ( .A(n1346), .B(n1344), .CI(n1321), .CO(n1312), .S(n1313) );
  CFA1X1 U1119 ( .A(n1331), .B(n1329), .CI(n1327), .CO(n1316), .S(n1317) );
  CFA1X1 U1120 ( .A(n1352), .B(n1354), .CI(n1356), .CO(n1318), .S(n1319) );
  CFA1X1 U1121 ( .A(n2129), .B(n1350), .CI(n1358), .CO(n1320), .S(n1321) );
  CFA1X1 U1122 ( .A(n2098), .B(n2067), .CI(n2160), .CO(n1322), .S(n1323) );
  CFA1X1 U1123 ( .A(n1945), .B(n1975), .CI(n1916), .CO(n1324), .S(n1325) );
  CFA1X1 U1124 ( .A(n2191), .B(n1857), .CI(n1886), .CO(n1326), .S(n1327) );
  CFA1X1 U1125 ( .A(n1800), .B(n2222), .CI(n2005), .CO(n1328), .S(n1329) );
  CFA1X1 U1126 ( .A(n1829), .B(n2036), .CI(n1770), .CO(n1330), .S(n1331) );
  CFA1X1 U1131 ( .A(n1374), .B(n1372), .CI(n1349), .CO(n1340), .S(n1341) );
  CFA1X1 U1132 ( .A(n1355), .B(n1357), .CI(n1353), .CO(n1342), .S(n1343) );
  CFA1X1 U1133 ( .A(n1378), .B(n1351), .CI(n1376), .CO(n1344), .S(n1345) );
  CFA1X1 U1134 ( .A(n1384), .B(n1380), .CI(n1382), .CO(n1346), .S(n1347) );
  CFA1X1 U1135 ( .A(n2006), .B(n1359), .CI(n2068), .CO(n1348), .S(n1349) );
  CFA1X1 U1136 ( .A(n2099), .B(n1976), .CI(n1917), .CO(n1350), .S(n1351) );
  CFA1X1 U1137 ( .A(n1887), .B(n1858), .CI(n1830), .CO(n1352), .S(n1353) );
  CFA1X1 U1138 ( .A(n1946), .B(n2130), .CI(n2161), .CO(n1354), .S(n1355) );
  CFA1X1 U1139 ( .A(n2037), .B(n2223), .CI(n2192), .CO(n1356), .S(n1357) );
  CFA1X1 U1142 ( .A(n1392), .B(n1390), .CI(n1367), .CO(n1362), .S(n1363) );
  CFA1X1 U1145 ( .A(n1379), .B(n1398), .CI(n1400), .CO(n1368), .S(n1369) );
  CFA1X1 U1148 ( .A(n1410), .B(n1404), .CI(n1402), .CO(n1374), .S(n1375) );
  CFA1X1 U1150 ( .A(n2131), .B(n1947), .CI(n1918), .CO(n1378), .S(n1379) );
  CFA1X1 U1151 ( .A(n2162), .B(n1888), .CI(n1831), .CO(n1380), .S(n1381) );
  CFA1X1 U1152 ( .A(n2007), .B(n2224), .CI(n2193), .CO(n1382), .S(n1383) );
  CFA1X1 U1153 ( .A(n1802), .B(n2069), .CI(n1859), .CO(n1384), .S(n1385) );
  CFA1X1 U1156 ( .A(n1420), .B(n1418), .CI(n1397), .CO(n1390), .S(n1391) );
  CFA1X1 U1162 ( .A(n1978), .B(n2070), .CI(n2132), .CO(n1402), .S(n1403) );
  CFA1X1 U1163 ( .A(n2163), .B(n1948), .CI(n1919), .CO(n1404), .S(n1405) );
  CFA1X1 U1164 ( .A(n2008), .B(n2194), .CI(n1889), .CO(n1406), .S(n1407) );
  CFA1X1 U1165 ( .A(n1860), .B(n2039), .CI(n2225), .CO(n1408), .S(n1409) );
  CFA1X1 U1167 ( .A(n3393), .B(n1415), .CI(n1438), .CO(n1412), .S(n1413) );
  CFA1X1 U1170 ( .A(n1448), .B(n1444), .CI(n1446), .CO(n1418), .S(n1419) );
  CFA1X1 U1173 ( .A(n1450), .B(n1452), .CI(n1456), .CO(n1424), .S(n1425) );
  CFA1X1 U1174 ( .A(n2133), .B(n1458), .CI(n2102), .CO(n1426), .S(n1427) );
  CFA1X1 U1177 ( .A(n2040), .B(n2226), .CI(n1861), .CO(n1432), .S(n1433) );
  CFA1X1 U1178 ( .A(n1833), .B(n2071), .CI(n1890), .CO(n1434), .S(n1435) );
  CFA1X1 U1182 ( .A(n1472), .B(n1449), .CI(n1470), .CO(n1442), .S(n1443) );
  CFA1X1 U1185 ( .A(n1459), .B(n1478), .CI(n1480), .CO(n1448), .S(n1449) );
  CFA1X1 U1187 ( .A(n2165), .B(n2010), .CI(n1950), .CO(n1452), .S(n1453) );
  CFA1X1 U1188 ( .A(n1891), .B(n1921), .CI(n1980), .CO(n1454), .S(n1455) );
  CFA1X1 U1189 ( .A(n2196), .B(n2227), .CI(n2072), .CO(n1456), .S(n1457) );
  CHA1X1 U1190 ( .A(n1862), .B(n1727), .CO(n1458), .S(n1459) );
  CFA1X1 U1192 ( .A(n1488), .B(n1486), .CI(n1467), .CO(n1462), .S(n1463) );
  CFA1X1 U1193 ( .A(n1490), .B(n1469), .CI(n1471), .CO(n1464), .S(n1465) );
  CFA1X1 U1194 ( .A(n1494), .B(n1473), .CI(n1492), .CO(n1466), .S(n1467) );
  CFA1X1 U1196 ( .A(n1498), .B(n1481), .CI(n1496), .CO(n1470), .S(n1471) );
  CFA1X1 U1197 ( .A(n2104), .B(n1500), .CI(n1502), .CO(n1472), .S(n1473) );
  CFA1X1 U1198 ( .A(n2135), .B(n2011), .CI(n1981), .CO(n1474), .S(n1475) );
  CFA1X1 U1200 ( .A(n2228), .B(n2042), .CI(n1892), .CO(n1478), .S(n1479) );
  CFA1X1 U1201 ( .A(n1863), .B(n1922), .CI(n2073), .CO(n1480), .S(n1481) );
  CFA1X1 U1202 ( .A(n1487), .B(n1485), .CI(n1506), .CO(n1482), .S(n1483) );
  CFA1X1 U1204 ( .A(n1512), .B(n1510), .CI(n1493), .CO(n1486), .S(n1487) );
  CFA1X1 U1205 ( .A(n1501), .B(n1495), .CI(n1514), .CO(n1488), .S(n1489) );
  CFA1X1 U1206 ( .A(n1520), .B(n1499), .CI(n1497), .CO(n1490), .S(n1491) );
  CFA1X1 U1207 ( .A(n1522), .B(n1518), .CI(n1516), .CO(n1492), .S(n1493) );
  CFA1X1 U1208 ( .A(n2105), .B(n1503), .CI(n2043), .CO(n1494), .S(n1495) );
  CFA1X1 U1209 ( .A(n2136), .B(n1982), .CI(n1952), .CO(n1496), .S(n1497) );
  CFA1X1 U1211 ( .A(n2229), .B(n1923), .CI(n2074), .CO(n1500), .S(n1501) );
  CFA1X1 U1214 ( .A(n1513), .B(n1528), .CI(n1511), .CO(n1506), .S(n1507) );
  CFA1X1 U1216 ( .A(n1519), .B(n1534), .CI(n1521), .CO(n1510), .S(n1511) );
  CFA1X1 U1217 ( .A(n1536), .B(n1517), .CI(n1523), .CO(n1512), .S(n1513) );
  CFA1X1 U1218 ( .A(n3214), .B(n1538), .CI(n1540), .CO(n1514), .S(n1515) );
  CFA1X1 U1219 ( .A(n2168), .B(n2137), .CI(n2075), .CO(n1516), .S(n1517) );
  CFA1X1 U1220 ( .A(n2199), .B(n2013), .CI(n1983), .CO(n1518), .S(n1519) );
  CFA1X1 U1221 ( .A(n2044), .B(n2230), .CI(n1924), .CO(n1520), .S(n1521) );
  CFA1X1 U1222 ( .A(n1894), .B(n2106), .CI(n1953), .CO(n1522), .S(n1523) );
  CFA1X1 U1223 ( .A(n1529), .B(n1527), .CI(n1546), .CO(n1524), .S(n1525) );
  CFA1X1 U1224 ( .A(n1533), .B(n1548), .CI(n1531), .CO(n1526), .S(n1527) );
  CFA1X1 U1225 ( .A(n1552), .B(n1550), .CI(n1535), .CO(n1528), .S(n1529) );
  CFA1X1 U1227 ( .A(n1558), .B(n1537), .CI(n1556), .CO(n1532), .S(n1533) );
  CFA1X1 U1228 ( .A(n2045), .B(n1560), .CI(n1543), .CO(n1534), .S(n1535) );
  CFA1X1 U1229 ( .A(n1984), .B(n2107), .CI(n1954), .CO(n1536), .S(n1537) );
  CFA1X1 U1231 ( .A(n2231), .B(n2076), .CI(n2200), .CO(n1540), .S(n1541) );
  CFA1X1 U1234 ( .A(n1553), .B(n1566), .CI(n1551), .CO(n1546), .S(n1547) );
  CFA1X1 U1235 ( .A(n1555), .B(n1568), .CI(n1570), .CO(n1548), .S(n1549) );
  CFA1X1 U1236 ( .A(n1561), .B(n1559), .CI(n1557), .CO(n1550), .S(n1551) );
  CFA1X1 U1237 ( .A(n1576), .B(n1574), .CI(n1572), .CO(n1552), .S(n1553) );
  CFA1X1 U1238 ( .A(n2170), .B(n1578), .CI(n2139), .CO(n1554), .S(n1555) );
  CFA1X1 U1239 ( .A(n2201), .B(n2046), .CI(n2015), .CO(n1556), .S(n1557) );
  CFA1X1 U1240 ( .A(n2077), .B(n3866), .CI(n1955), .CO(n1558), .S(n1559) );
  CFA1X1 U1244 ( .A(n1577), .B(n1586), .CI(n1588), .CO(n1566), .S(n1567) );
  CFA1X1 U1246 ( .A(n1579), .B(n1592), .CI(n1594), .CO(n1570), .S(n1571) );
  CFA1X1 U1247 ( .A(n2171), .B(n2047), .CI(n2140), .CO(n1572), .S(n1573) );
  CFA1X1 U1248 ( .A(n2202), .B(n2016), .CI(n2078), .CO(n1574), .S(n1575) );
  CFA1X1 U1249 ( .A(n2109), .B(n2233), .CI(n1986), .CO(n1576), .S(n1577) );
  CFA1X1 U1251 ( .A(n1585), .B(n1583), .CI(n1598), .CO(n1580), .S(n1581) );
  CFA1X1 U1252 ( .A(n1587), .B(n1600), .CI(n1589), .CO(n1582), .S(n1583) );
  CFA1X1 U1255 ( .A(n2172), .B(n1608), .CI(n1610), .CO(n1588), .S(n1589) );
  CFA1X1 U1256 ( .A(n2203), .B(n2079), .CI(n2048), .CO(n1590), .S(n1591) );
  CFA1X1 U1257 ( .A(n2110), .B(n2234), .CI(n1987), .CO(n1592), .S(n1593) );
  CFA1X1 U1259 ( .A(n1601), .B(n1599), .CI(n1614), .CO(n1596), .S(n1597) );
  CFA1X1 U1260 ( .A(n1605), .B(n1616), .CI(n1603), .CO(n1598), .S(n1599) );
  CFA1X1 U1261 ( .A(n1607), .B(n1618), .CI(n1609), .CO(n1600), .S(n1601) );
  CFA1X1 U1263 ( .A(n2173), .B(n1611), .CI(n2142), .CO(n1604), .S(n1605) );
  CFA1X1 U1264 ( .A(n2049), .B(n2080), .CI(n2018), .CO(n1606), .S(n1607) );
  CFA1X1 U1265 ( .A(n2111), .B(n2235), .CI(n2204), .CO(n1608), .S(n1609) );
  CFA1X1 U1267 ( .A(n1617), .B(n1615), .CI(n1628), .CO(n1612), .S(n1613) );
  CFA1X1 U1268 ( .A(n1632), .B(n1630), .CI(n1619), .CO(n1614), .S(n1615) );
  CFA1X1 U1269 ( .A(n1623), .B(n1625), .CI(n1621), .CO(n1616), .S(n1617) );
  CFA1X1 U1271 ( .A(n2205), .B(n2081), .CI(n2174), .CO(n1620), .S(n1621) );
  CFA1X1 U1273 ( .A(n1989), .B(n2143), .CI(n2050), .CO(n1624), .S(n1625) );
  CFA1X1 U1274 ( .A(n1631), .B(n1629), .CI(n1642), .CO(n1626), .S(n1627) );
  CFA1X1 U1275 ( .A(n1646), .B(n1633), .CI(n1644), .CO(n1628), .S(n1629) );
  CFA1X1 U1276 ( .A(n1648), .B(n1637), .CI(n1635), .CO(n1630), .S(n1631) );
  CFA1X1 U1277 ( .A(n2175), .B(n1650), .CI(n1639), .CO(n1632), .S(n1633) );
  CFA1X1 U1278 ( .A(n2082), .B(n2113), .CI(n2206), .CO(n1634), .S(n1635) );
  CFA1X1 U1281 ( .A(n1645), .B(n1643), .CI(n1654), .CO(n1640), .S(n1641) );
  CFA1X1 U1282 ( .A(n1649), .B(n1656), .CI(n1647), .CO(n1642), .S(n1643) );
  CFA1X1 U1283 ( .A(n1660), .B(n1651), .CI(n1658), .CO(n1644), .S(n1645) );
  CFA1X1 U1284 ( .A(n2207), .B(n1662), .CI(n2114), .CO(n1646), .S(n1647) );
  CFA1X1 U1285 ( .A(n2145), .B(n2238), .CI(n2052), .CO(n1648), .S(n1649) );
  CFA1X1 U1287 ( .A(n1657), .B(n1655), .CI(n1666), .CO(n1652), .S(n1653) );
  CFA1X1 U1288 ( .A(n1659), .B(n1668), .CI(n1661), .CO(n1654), .S(n1655) );
  CFA1X1 U1289 ( .A(n1663), .B(n1670), .CI(n1672), .CO(n1656), .S(n1657) );
  CFA1X1 U1291 ( .A(n2146), .B(n2239), .CI(n2208), .CO(n1660), .S(n1661) );
  CHA1X1 U1292 ( .A(n2084), .B(n2053), .CO(n1662), .S(n1663) );
  CFA1X1 U1293 ( .A(n1676), .B(n1667), .CI(n1669), .CO(n1664), .S(n1665) );
  CFA1X1 U1294 ( .A(n1673), .B(n1678), .CI(n1671), .CO(n1666), .S(n1667) );
  CFA1X1 U1295 ( .A(n2209), .B(n1680), .CI(n1682), .CO(n1668), .S(n1669) );
  CFA1X1 U1296 ( .A(n2085), .B(n3104), .CI(n2147), .CO(n1670), .S(n1671) );
  CFA1X1 U1297 ( .A(n3477), .B(n3106), .CI(n2116), .CO(n1672), .S(n1673) );
  CFA1X1 U1298 ( .A(n1679), .B(n1677), .CI(n1686), .CO(n1674), .S(n1675) );
  CFA1X1 U1299 ( .A(n1690), .B(n1681), .CI(n1688), .CO(n1676), .S(n1677) );
  CFA1X1 U1300 ( .A(n3103), .B(n1683), .CI(n1734), .CO(n1678), .S(n1679) );
  CFA1X1 U1301 ( .A(n2179), .B(n2241), .CI(n2210), .CO(n1680), .S(n1681) );
  CHA1X1 U1302 ( .A(n2117), .B(n2086), .CO(n1682), .S(n1683) );
  CFA1X1 U1303 ( .A(n1689), .B(n1687), .CI(n1694), .CO(n1684), .S(n1685) );
  CFA1X1 U1304 ( .A(n1698), .B(n1691), .CI(n1696), .CO(n1686), .S(n1687) );
  CFA1X1 U1305 ( .A(n2180), .B(n2242), .CI(n2118), .CO(n1688), .S(n1689) );
  CFA1X1 U1306 ( .A(n2087), .B(n2149), .CI(n2211), .CO(n1690), .S(n1691) );
  CFA1X1 U1307 ( .A(n1697), .B(n1695), .CI(n1702), .CO(n1692), .S(n1693) );
  CFA1X1 U1308 ( .A(n2212), .B(n1704), .CI(n1699), .CO(n1694), .S(n1695) );
  CHA1X1 U1310 ( .A(n2150), .B(n2119), .CO(n1698), .S(n1699) );
  CFA1X1 U1311 ( .A(n1708), .B(n1703), .CI(n1705), .CO(n1700), .S(n1701) );
  CFA1X1 U1312 ( .A(n2182), .B(n1710), .CI(n2244), .CO(n1702), .S(n1703) );
  CFA1X1 U1313 ( .A(n2120), .B(n2213), .CI(n2151), .CO(n1704), .S(n1705) );
  CFA1X1 U1314 ( .A(n1711), .B(n1709), .CI(n1714), .CO(n1706), .S(n1707) );
  CFA1X1 U1315 ( .A(n2214), .B(n2245), .CI(n2183), .CO(n1708), .S(n1709) );
  CHA1X1 U1316 ( .A(n1736), .B(n2152), .CO(n1710), .S(n1711) );
  CFA1X1 U1317 ( .A(n2246), .B(n1715), .CI(n1718), .CO(n1712), .S(n1713) );
  CFA1X1 U1319 ( .A(n2216), .B(n1719), .CI(n2247), .CO(n1716), .S(n1717) );
  CHA1X1 U1320 ( .A(n1737), .B(n2185), .CO(n1718), .S(n1719) );
  CFA1X1 U1321 ( .A(n2186), .B(n2248), .CI(n2217), .CO(n1720), .S(n1721) );
  CHA1X1 U1322 ( .A(n1738), .B(n2249), .CO(n1722), .S(n1723) );
  COND2X1 U1335 ( .A(n144), .B(n2263), .C(n3173), .D(n2262), .Z(n1749) );
  COND2X1 U1336 ( .A(n144), .B(n2264), .C(n3086), .D(n2263), .Z(n1750) );
  COND2X1 U1337 ( .A(n144), .B(n2265), .C(n3114), .D(n2264), .Z(n1751) );
  COND2X1 U1338 ( .A(n144), .B(n2266), .C(n3173), .D(n2265), .Z(n1752) );
  COND2X1 U1339 ( .A(n144), .B(n2267), .C(n3085), .D(n2266), .Z(n1753) );
  COND2X1 U1340 ( .A(n2268), .B(net21320), .C(n3114), .D(n2267), .Z(n1754) );
  COND2X1 U1345 ( .A(n144), .B(n2273), .C(n2272), .D(n3114), .Z(n1759) );
  COND2X1 U1346 ( .A(n144), .B(n2274), .C(n3085), .D(n2273), .Z(n1760) );
  COND2X1 U1347 ( .A(n144), .B(n2275), .C(n3173), .D(n2274), .Z(n1761) );
  COND2X1 U1348 ( .A(n144), .B(n2276), .C(n3086), .D(n2275), .Z(n1762) );
  COND2X1 U1349 ( .A(n144), .B(n2277), .C(n3086), .D(n2276), .Z(n1763) );
  COND2X1 U1350 ( .A(net21320), .B(n2278), .C(n2277), .D(n3173), .Z(n1764) );
  COND2X1 U1352 ( .A(n144), .B(n2280), .C(n3173), .D(n2279), .Z(n1766) );
  COND2X1 U1355 ( .A(n2283), .B(n144), .C(n3114), .D(n2282), .Z(n1769) );
  CND2IX1 U1389 ( .B(n3979), .A(net18487), .Z(n2284) );
  COND2X1 U1402 ( .A(net21433), .B(n2296), .C(net19192), .D(n2295), .Z(n1781)
         );
  COND2X1 U1403 ( .A(net21433), .B(n3287), .C(net19192), .D(n2296), .Z(n1782)
         );
  COND2X1 U1406 ( .A(net21434), .B(n2300), .C(net19192), .D(n2299), .Z(n1785)
         );
  COND2X1 U1413 ( .A(net21433), .B(n2307), .C(net19192), .D(n2306), .Z(n1792)
         );
  COND2X1 U1414 ( .A(net21434), .B(n2308), .C(net19192), .D(n2307), .Z(n1793)
         );
  COND2X1 U1415 ( .A(net21433), .B(n2309), .C(net19193), .D(n2308), .Z(n1794)
         );
  COND2X1 U1417 ( .A(net21433), .B(n2311), .C(net19192), .D(n2310), .Z(n1796)
         );
  COND2X1 U1420 ( .A(net21433), .B(n2314), .C(net19193), .D(n3752), .Z(n1799)
         );
  COND2X1 U1421 ( .A(net21434), .B(n3758), .C(net19193), .D(n3750), .Z(n1800)
         );
  COND2X1 U1422 ( .A(n2316), .B(net21434), .C(net19192), .D(n3758), .Z(n1801)
         );
  COND2X1 U1463 ( .A(net21696), .B(n2323), .C(net22006), .D(n2322), .Z(n842)
         );
  COND2X1 U1465 ( .A(net21696), .B(n2325), .C(net22007), .D(n2324), .Z(n1808)
         );
  COND2X1 U1467 ( .A(net21696), .B(n2327), .C(net22007), .D(n2326), .Z(n1810)
         );
  COND2X1 U1468 ( .A(net21696), .B(n2328), .C(net22006), .D(n2327), .Z(n1811)
         );
  COND2X1 U1469 ( .A(net21696), .B(n2329), .C(net22007), .D(n2328), .Z(n1812)
         );
  COND2X1 U1471 ( .A(net21696), .B(n2331), .C(net22007), .D(n2330), .Z(n1814)
         );
  COND2X1 U1473 ( .A(net21696), .B(n2333), .C(net22006), .D(n2332), .Z(n1816)
         );
  COND2X1 U1474 ( .A(net21696), .B(n2334), .C(net22007), .D(n2333), .Z(n1817)
         );
  COND2X1 U1475 ( .A(net21696), .B(n2335), .C(net22007), .D(n2334), .Z(n1818)
         );
  COND2X1 U1476 ( .A(net21696), .B(n2336), .C(net22006), .D(n2335), .Z(n1819)
         );
  COND2X1 U1477 ( .A(net21696), .B(n2337), .C(net22006), .D(n2336), .Z(n1820)
         );
  COND2X1 U1478 ( .A(net21696), .B(n2338), .C(net22006), .D(n2337), .Z(n1821)
         );
  COND2X1 U1480 ( .A(n126), .B(n2340), .C(net22006), .D(n2339), .Z(n1823) );
  COND2X1 U1482 ( .A(n126), .B(n2342), .C(net22007), .D(n2341), .Z(n1825) );
  COND2X1 U1483 ( .A(net21696), .B(n2343), .C(net22006), .D(n2342), .Z(n1826)
         );
  COND2X1 U1484 ( .A(n126), .B(n2344), .C(net22007), .D(n2343), .Z(n1827) );
  COND2X1 U1485 ( .A(net21696), .B(n3782), .C(net22007), .D(n2344), .Z(n1828)
         );
  COND2X1 U1487 ( .A(n126), .B(n2347), .C(net22007), .D(n2346), .Z(n1830) );
  COND2X1 U1488 ( .A(net21696), .B(n2348), .C(net22007), .D(n2347), .Z(n1831)
         );
  CNR2IX2 U1490 ( .B(n3979), .A(net22006), .Z(n1833) );
  COND2X1 U1530 ( .A(net21312), .B(n2356), .C(net21512), .D(n2355), .Z(n864)
         );
  COND2X1 U1532 ( .A(net21311), .B(n2358), .C(net21512), .D(n2357), .Z(n890)
         );
  COND2X1 U1533 ( .A(net21311), .B(n2359), .C(net21512), .D(n2358), .Z(n1840)
         );
  COND2X1 U1536 ( .A(net21311), .B(n2362), .C(net21512), .D(n2361), .Z(n1842)
         );
  COND2X1 U1538 ( .A(net21312), .B(n2364), .C(net21512), .D(n2363), .Z(n1844)
         );
  COND2X1 U1539 ( .A(net21312), .B(n2365), .C(net21512), .D(n2364), .Z(n1845)
         );
  COND2X1 U1542 ( .A(net21311), .B(n2368), .C(net21512), .D(n2367), .Z(n1848)
         );
  COND2X1 U1543 ( .A(net21311), .B(n2369), .C(net21512), .D(n2368), .Z(n1849)
         );
  COND2X1 U1544 ( .A(net21311), .B(n2370), .C(net21512), .D(n2369), .Z(n1850)
         );
  COND2X1 U1545 ( .A(net21312), .B(n2371), .C(net21512), .D(n2370), .Z(n1851)
         );
  COND2X1 U1546 ( .A(n117), .B(n2372), .C(net21512), .D(n2371), .Z(n1852) );
  COND2X1 U1547 ( .A(net21311), .B(n2373), .C(net21512), .D(n2372), .Z(n1853)
         );
  COND2X1 U1548 ( .A(net21312), .B(n2374), .C(net21512), .D(n2373), .Z(n1854)
         );
  COND2X1 U1549 ( .A(n2375), .B(n117), .C(net19281), .D(n2374), .Z(n1855) );
  COND2X1 U1550 ( .A(net21311), .B(n2376), .C(net21512), .D(n2375), .Z(n1856)
         );
  COND2X1 U1551 ( .A(net21311), .B(n2377), .C(net21512), .D(n2376), .Z(n1857)
         );
  COND2X1 U1552 ( .A(net21312), .B(n2378), .C(net21512), .D(n2377), .Z(n1858)
         );
  COND2X1 U1553 ( .A(n117), .B(n2379), .C(net19281), .D(n2378), .Z(n1859) );
  COND2X1 U1554 ( .A(n117), .B(n2380), .C(net19281), .D(n2379), .Z(n1860) );
  COND2X1 U1555 ( .A(net21312), .B(n2381), .C(net21512), .D(n2380), .Z(n1861)
         );
  COND2X1 U1556 ( .A(n2382), .B(n117), .C(net19281), .D(n2381), .Z(n1862) );
  CND2IX1 U1590 ( .B(n3979), .A(net19268), .Z(n2383) );
  COND2X1 U1593 ( .A(n2385), .B(net22344), .C(net21250), .D(n2384), .Z(n1865)
         );
  COND2X1 U1595 ( .A(net22351), .B(n2387), .C(net21250), .D(n2386), .Z(n1867)
         );
  COND2X1 U1597 ( .A(n108), .B(n2389), .C(net21250), .D(n2388), .Z(n1869) );
  COND2X1 U1601 ( .A(n108), .B(n2393), .C(net21248), .D(n2392), .Z(n954) );
  COND2X1 U1605 ( .A(n108), .B(n2397), .C(net21249), .D(n2396), .Z(n1875) );
  COND2X1 U1606 ( .A(n108), .B(n2398), .C(net21250), .D(n2397), .Z(n1876) );
  COND2X1 U1607 ( .A(n108), .B(n2399), .C(net21249), .D(n2398), .Z(n1877) );
  COND2X1 U1609 ( .A(n108), .B(n2401), .C(net21250), .D(n2400), .Z(n1879) );
  COND2X1 U1610 ( .A(n108), .B(n2402), .C(net21248), .D(n2401), .Z(n1880) );
  COND2X1 U1611 ( .A(n108), .B(n2403), .C(net21248), .D(n2402), .Z(n1881) );
  COND2X1 U1612 ( .A(n108), .B(n2404), .C(net21250), .D(n2403), .Z(n1882) );
  COND2X1 U1613 ( .A(n108), .B(n2405), .C(net21248), .D(n2404), .Z(n1883) );
  COND2X1 U1615 ( .A(n108), .B(n2407), .C(net21250), .D(n2406), .Z(n1885) );
  COND2X1 U1616 ( .A(n108), .B(n2408), .C(net21250), .D(n2407), .Z(n1886) );
  COND2X1 U1617 ( .A(n108), .B(n2409), .C(net21250), .D(n2408), .Z(n1887) );
  COND2X1 U1618 ( .A(n108), .B(n2410), .C(net21249), .D(n2409), .Z(n1888) );
  COND2X1 U1619 ( .A(n108), .B(n2411), .C(net21250), .D(n2410), .Z(n1889) );
  COND2X1 U1621 ( .A(n108), .B(n2413), .C(net21248), .D(n2412), .Z(n1891) );
  COND2X1 U1622 ( .A(net22344), .B(n2414), .C(net21250), .D(n2413), .Z(n1892)
         );
  CAOR1X1 U1659 ( .A(net21744), .B(net21344), .C(n2417), .Z(n1895) );
  COND2X1 U1660 ( .A(n2418), .B(n3328), .C(net21744), .D(n2417), .Z(n1896) );
  COND2X1 U1661 ( .A(n2418), .B(net21744), .C(n2419), .D(net21344), .Z(n1897)
         );
  COND2X1 U1663 ( .A(net21344), .B(n2421), .C(net21744), .D(n2420), .Z(n1899)
         );
  COND2X1 U1666 ( .A(net21344), .B(n2424), .C(net21744), .D(n2423), .Z(n1902)
         );
  COND2X1 U1667 ( .A(n3328), .B(n2425), .C(net21744), .D(n2424), .Z(n1903) );
  COND2X1 U1668 ( .A(n3328), .B(n2426), .C(net21744), .D(n2425), .Z(n1904) );
  COND2X1 U1669 ( .A(n3328), .B(n2427), .C(net21744), .D(n2426), .Z(n1905) );
  COND2X1 U1672 ( .A(net21344), .B(n2430), .C(net21744), .D(n2429), .Z(n1907)
         );
  COND2X1 U1673 ( .A(n3328), .B(n2431), .C(net21744), .D(n2430), .Z(n1908) );
  COND2X1 U1674 ( .A(n3328), .B(n2432), .C(net21744), .D(n2431), .Z(n1909) );
  COND2X1 U1676 ( .A(net21344), .B(n2434), .C(net21744), .D(n2433), .Z(n1911)
         );
  COND2X1 U1680 ( .A(net21344), .B(n2438), .C(net21744), .D(n2437), .Z(n1915)
         );
  COND2X1 U1681 ( .A(net21344), .B(n3044), .C(net21744), .D(n2438), .Z(n1916)
         );
  COND2X1 U1682 ( .A(n99), .B(n2440), .C(net21744), .D(n2439), .Z(n1917) );
  COND2X1 U1683 ( .A(net21344), .B(n2441), .C(net21744), .D(n2440), .Z(n1918)
         );
  COND2X1 U1684 ( .A(n3328), .B(n2442), .C(net21744), .D(n2441), .Z(n1919) );
  COND2X1 U1686 ( .A(net21344), .B(n3243), .C(net21744), .D(n2443), .Z(n1921)
         );
  COND2X1 U1687 ( .A(n99), .B(n2445), .C(net21744), .D(n2444), .Z(n1922) );
  COND2X1 U1689 ( .A(n3328), .B(n2447), .C(net21744), .D(n2446), .Z(n1924) );
  COND2X1 U1690 ( .A(n2448), .B(net21344), .C(net21744), .D(n2447), .Z(n1925)
         );
  CND2IX1 U1724 ( .B(n3979), .A(n3925), .Z(n2449) );
  COND2X1 U1727 ( .A(n2451), .B(net21801), .C(n87), .D(n2450), .Z(n1928) );
  COND2X1 U1728 ( .A(n2451), .B(net22326), .C(n2452), .D(net21802), .Z(n1929)
         );
  COND2X1 U1729 ( .A(net21801), .B(n2453), .C(n87), .D(n2452), .Z(n1930) );
  COND2X1 U1733 ( .A(net21802), .B(n2457), .C(net22327), .D(n2456), .Z(n1934)
         );
  COND2X1 U1734 ( .A(net21802), .B(n2458), .C(n87), .D(n2457), .Z(n1935) );
  COND2X1 U1735 ( .A(net21802), .B(n2459), .C(net21846), .D(n2458), .Z(n1936)
         );
  COND2X1 U1736 ( .A(net21802), .B(n2460), .C(net22326), .D(n2459), .Z(n1937)
         );
  COND2X1 U1738 ( .A(net21801), .B(n2462), .C(n87), .D(n2461), .Z(n1938) );
  COND2X1 U1740 ( .A(n90), .B(n2464), .C(net21846), .D(n2463), .Z(n1939) );
  COND2X1 U1742 ( .A(n90), .B(n2466), .C(net21846), .D(n2465), .Z(n1941) );
  COND2X1 U1744 ( .A(n3749), .B(n90), .C(net21846), .D(n2467), .Z(n1943) );
  COND2X1 U1745 ( .A(n3887), .B(n2469), .C(net21846), .D(n2468), .Z(n1944) );
  COND2X1 U1746 ( .A(n3887), .B(n2470), .C(net22326), .D(n2469), .Z(n1945) );
  COND2X1 U1748 ( .A(net21801), .B(n2472), .C(net22327), .D(n2471), .Z(n1947)
         );
  COND2X1 U1749 ( .A(net21801), .B(n2473), .C(net22326), .D(n2472), .Z(n1948)
         );
  COND2X1 U1750 ( .A(net21802), .B(n2474), .C(net22327), .D(n2473), .Z(n1949)
         );
  COND2X1 U1752 ( .A(n2476), .B(net21802), .C(net21846), .D(n2475), .Z(n1951)
         );
  COND2X1 U1754 ( .A(net21802), .B(n2478), .C(net21846), .D(n2477), .Z(n1953)
         );
  COND2X1 U1755 ( .A(net21802), .B(n2479), .C(net22327), .D(n2478), .Z(n1954)
         );
  COND2X1 U1756 ( .A(net21801), .B(n2480), .C(net22326), .D(n2479), .Z(n1955)
         );
  COND2X1 U1795 ( .A(n2484), .B(n3651), .C(n2485), .D(n3871), .Z(n1960) );
  COND2X1 U1798 ( .A(n3871), .B(n2488), .C(n3942), .D(n2487), .Z(n1963) );
  COND2X1 U1799 ( .A(n3344), .B(n2489), .C(n3651), .D(n2488), .Z(n1964) );
  COND2X1 U1802 ( .A(n3344), .B(n2492), .C(n3651), .D(n2491), .Z(n1967) );
  COND2X1 U1803 ( .A(n3871), .B(n2493), .C(n3941), .D(n2492), .Z(n1968) );
  COND2X1 U1805 ( .A(n3871), .B(n2495), .C(n3942), .D(n2494), .Z(n1970) );
  COND2X1 U1807 ( .A(n3871), .B(n2497), .C(n3651), .D(n2496), .Z(n1971) );
  COND2X1 U1812 ( .A(n3231), .B(n2502), .C(n3942), .D(n2501), .Z(n1976) );
  COND2X1 U1815 ( .A(n3344), .B(n2505), .C(n3651), .D(n2504), .Z(n1979) );
  COND2X1 U1816 ( .A(n3871), .B(n2506), .C(n3651), .D(n2505), .Z(n1980) );
  COND2X1 U1817 ( .A(n3871), .B(n2507), .C(n3941), .D(n2506), .Z(n1981) );
  COND2X1 U1819 ( .A(n3871), .B(n2509), .C(n3941), .D(n2508), .Z(n1983) );
  COND2X1 U1820 ( .A(n3871), .B(n2510), .C(n3651), .D(n2509), .Z(n1984) );
  COND2X1 U1821 ( .A(n3871), .B(n2511), .C(n3651), .D(n2510), .Z(n1985) );
  COND2X1 U1865 ( .A(net21353), .B(n2521), .C(net19215), .D(n2520), .Z(n1995)
         );
  COND2X1 U1866 ( .A(net21352), .B(n2522), .C(net19216), .D(n2521), .Z(n1996)
         );
  COND2X1 U1867 ( .A(n2523), .B(net21352), .C(net19216), .D(n2522), .Z(n1997)
         );
  COND2X1 U1868 ( .A(net21352), .B(n2524), .C(net19215), .D(n2523), .Z(n1998)
         );
  COND2X1 U1869 ( .A(net21353), .B(n2525), .C(net19215), .D(n2524), .Z(n1999)
         );
  COND2X1 U1870 ( .A(net21353), .B(n2526), .C(net19216), .D(n2525), .Z(n2000)
         );
  COND2X1 U1874 ( .A(net21353), .B(n2530), .C(net19216), .D(n2529), .Z(n2003)
         );
  COND2X1 U1875 ( .A(net21353), .B(n2531), .C(net19215), .D(n2530), .Z(n2004)
         );
  COND2X1 U1876 ( .A(net21352), .B(n2532), .C(net19215), .D(n2531), .Z(n2005)
         );
  COND2X1 U1878 ( .A(net21352), .B(n2534), .C(net19216), .D(n2533), .Z(n2007)
         );
  COND2X1 U1879 ( .A(net21353), .B(n3617), .C(net19216), .D(n2534), .Z(n2008)
         );
  COND2X1 U1881 ( .A(net21352), .B(n2537), .C(net19216), .D(n2536), .Z(n2010)
         );
  COND2X1 U1882 ( .A(net21352), .B(n2538), .C(net19215), .D(n2537), .Z(n2011)
         );
  COND2X1 U1886 ( .A(net21352), .B(n2542), .C(net19215), .D(n2541), .Z(n2015)
         );
  COND2X1 U1887 ( .A(net21353), .B(n2543), .C(net19215), .D(n2542), .Z(n2016)
         );
  COND2X1 U1889 ( .A(n2545), .B(net21352), .C(net19216), .D(n2544), .Z(n2018)
         );
  COND2X1 U1890 ( .A(net21352), .B(n2546), .C(net19215), .D(n2545), .Z(n2019)
         );
  COND2X1 U1928 ( .A(n2550), .B(n3228), .C(n3660), .D(n2549), .Z(n2023) );
  COND2X1 U1929 ( .A(n2550), .B(n3660), .C(n3550), .D(n2551), .Z(n2024) );
  COND2X1 U1930 ( .A(n3550), .B(n2552), .C(n3660), .D(n3342), .Z(n2025) );
  COND2X1 U1931 ( .A(n3228), .B(n2553), .C(n3618), .D(n2552), .Z(n2026) );
  COND2X1 U1932 ( .A(n3228), .B(n2554), .C(n3660), .D(n2553), .Z(n2027) );
  COND2X1 U1934 ( .A(n3228), .B(n3786), .C(n3618), .D(n2555), .Z(n2029) );
  COND2X1 U1935 ( .A(n3893), .B(n2557), .C(n3618), .D(n2556), .Z(n2030) );
  COND2X1 U1936 ( .A(n3893), .B(n2558), .C(n3660), .D(n2557), .Z(n2031) );
  COND2X1 U1937 ( .A(n3893), .B(n2559), .C(n3660), .D(n2558), .Z(n2032) );
  COND2X1 U1938 ( .A(n63), .B(n2560), .C(n3660), .D(n2559), .Z(n2033) );
  COND2X1 U1940 ( .A(n63), .B(n2562), .C(n3660), .D(n2561), .Z(n2035) );
  COND2X1 U1941 ( .A(n3893), .B(n2563), .C(n3660), .D(n2562), .Z(n2036) );
  COND2X1 U1942 ( .A(n3550), .B(n2564), .C(n3660), .D(n2563), .Z(n2037) );
  COND2X1 U1944 ( .A(n3551), .B(n2566), .C(n3660), .D(n3650), .Z(n2039) );
  COND2X1 U1945 ( .A(n3228), .B(n3623), .C(n3660), .D(n2566), .Z(n2040) );
  COND2X1 U1946 ( .A(n3894), .B(n2568), .C(n3660), .D(n2567), .Z(n2041) );
  COND2X1 U1947 ( .A(n2569), .B(n3893), .C(n3660), .D(n2568), .Z(n2042) );
  COND2X1 U1948 ( .A(n3551), .B(n2570), .C(n3660), .D(n2569), .Z(n2043) );
  COND2X1 U1949 ( .A(n3551), .B(n2571), .C(n3660), .D(n2570), .Z(n2044) );
  COND2X1 U1951 ( .A(n3551), .B(n2573), .C(n3618), .D(n2572), .Z(n2046) );
  COND2X1 U1952 ( .A(n3551), .B(n2574), .C(n3618), .D(n2573), .Z(n2047) );
  COND2X1 U1953 ( .A(n3893), .B(n2575), .C(n3618), .D(n2574), .Z(n2048) );
  COND2X1 U1958 ( .A(n2580), .B(n3550), .C(n3660), .D(n2579), .Z(n2053) );
  COND2X1 U1996 ( .A(n2583), .B(n3145), .C(n2584), .D(n54), .Z(n2057) );
  COND2X1 U1997 ( .A(n3250), .B(n2585), .C(n3145), .D(n2584), .Z(n2058) );
  COND2X1 U1998 ( .A(n3250), .B(n2586), .C(n3145), .D(n2585), .Z(n2059) );
  COND2X1 U1999 ( .A(n54), .B(n2587), .C(n3145), .D(n2586), .Z(n2060) );
  COND2X1 U2000 ( .A(n3250), .B(n2588), .C(n3145), .D(n2587), .Z(n2061) );
  COND2X1 U2005 ( .A(n3250), .B(n3757), .C(n3145), .D(n2592), .Z(n2066) );
  COND2X1 U2006 ( .A(n54), .B(n2594), .C(n3145), .D(n2593), .Z(n2067) );
  COND2X1 U2007 ( .A(n3250), .B(n2595), .C(n3145), .D(n2594), .Z(n2068) );
  COND2X1 U2008 ( .A(n3250), .B(n2596), .C(n3453), .D(n2595), .Z(n2069) );
  COND2X1 U2009 ( .A(n3806), .B(n2597), .C(n3145), .D(n2596), .Z(n2070) );
  COND2X1 U2010 ( .A(n54), .B(n2598), .C(n3145), .D(n2597), .Z(n2071) );
  COND2X1 U2011 ( .A(n3806), .B(n2599), .C(n3145), .D(n2598), .Z(n2072) );
  COND2X1 U2012 ( .A(n3806), .B(n2600), .C(n3145), .D(n2599), .Z(n2073) );
  COND2X1 U2013 ( .A(n54), .B(n2601), .C(n3453), .D(n2600), .Z(n2074) );
  COND2X1 U2014 ( .A(n3250), .B(n2602), .C(n3145), .D(n2601), .Z(n2075) );
  COND2X1 U2015 ( .A(n54), .B(n2603), .C(n3145), .D(n2602), .Z(n2076) );
  COND2X1 U2016 ( .A(n3250), .B(n2604), .C(n3145), .D(n2603), .Z(n2077) );
  COND2X1 U2017 ( .A(n54), .B(n2605), .C(n3145), .D(n2604), .Z(n2078) );
  COND2X1 U2018 ( .A(n3250), .B(n2606), .C(n3145), .D(n2605), .Z(n2079) );
  COND2X1 U2019 ( .A(n3806), .B(n2607), .C(n3145), .D(n2606), .Z(n2080) );
  COND2X1 U2020 ( .A(n54), .B(n2608), .C(n3145), .D(n2607), .Z(n2081) );
  COND2X1 U2021 ( .A(n54), .B(n2609), .C(n3145), .D(n2608), .Z(n2082) );
  COND2X1 U2024 ( .A(n3806), .B(n2612), .C(n3145), .D(n2611), .Z(n2085) );
  COND2X1 U2064 ( .A(n45), .B(n2618), .C(n3938), .D(n2617), .Z(n2091) );
  COND2X1 U2066 ( .A(n45), .B(n3155), .C(n3938), .D(n2619), .Z(n2093) );
  COND2X1 U2067 ( .A(n45), .B(n2621), .C(n3939), .D(n2620), .Z(n2094) );
  COND2X1 U2068 ( .A(n3787), .B(n2622), .C(n3938), .D(n3156), .Z(n2095) );
  COND2X1 U2069 ( .A(n45), .B(n2623), .C(n3938), .D(n2622), .Z(n2096) );
  COND2X1 U2070 ( .A(n45), .B(n2624), .C(n3938), .D(n2623), .Z(n2097) );
  COND2X1 U2071 ( .A(n45), .B(n2625), .C(n3939), .D(n2624), .Z(n2098) );
  COND2X1 U2072 ( .A(n3787), .B(n2626), .C(n3939), .D(n2625), .Z(n2099) );
  COND2X1 U2075 ( .A(n45), .B(n2629), .C(n3939), .D(n2628), .Z(n2102) );
  COND2X1 U2076 ( .A(n45), .B(n2630), .C(n3939), .D(n2629), .Z(n2103) );
  COND2X1 U2079 ( .A(n45), .B(n2633), .C(n3938), .D(n2632), .Z(n2106) );
  COND2X1 U2080 ( .A(n45), .B(n2634), .C(n3939), .D(n2633), .Z(n2107) );
  COND2X1 U2081 ( .A(n45), .B(n2635), .C(n3938), .D(n2634), .Z(n2108) );
  COND2X1 U2083 ( .A(n45), .B(n2637), .C(n3939), .D(n2636), .Z(n2110) );
  COND2X1 U2084 ( .A(n45), .B(n2638), .C(n3938), .D(n2637), .Z(n2111) );
  COND2X1 U2085 ( .A(n45), .B(n2639), .C(n3938), .D(n2638), .Z(n2112) );
  COND2X1 U2086 ( .A(n45), .B(n2640), .C(n3939), .D(n2639), .Z(n2113) );
  COND2X1 U2088 ( .A(n45), .B(n2642), .C(n3939), .D(n2641), .Z(n2115) );
  COND2X1 U2090 ( .A(n45), .B(n2644), .C(n3939), .D(n2643), .Z(n2117) );
  COND2X1 U2091 ( .A(n3787), .B(n2645), .C(n3939), .D(n2644), .Z(n2118) );
  COND2X1 U2129 ( .A(n2649), .B(n3904), .C(n3803), .D(n2648), .Z(n2122) );
  COND2X1 U2130 ( .A(n2649), .B(n3803), .C(n2650), .D(n3954), .Z(n2123) );
  COND2X1 U2131 ( .A(n3904), .B(n2651), .C(n3803), .D(n2650), .Z(n2124) );
  COND2X1 U2133 ( .A(n2653), .B(n3954), .C(n3803), .D(n2652), .Z(n2126) );
  COND2X1 U2135 ( .A(n3953), .B(n2655), .C(n3803), .D(n2654), .Z(n2128) );
  COND2X1 U2137 ( .A(n3904), .B(n2657), .C(n3803), .D(n2656), .Z(n2130) );
  COND2X1 U2138 ( .A(n3905), .B(n2658), .C(n3803), .D(n2657), .Z(n2131) );
  COND2X1 U2140 ( .A(n3905), .B(n2660), .C(n3803), .D(n2659), .Z(n2133) );
  COND2X1 U2143 ( .A(n3953), .B(n2663), .C(n3803), .D(n2662), .Z(n2136) );
  COND2X1 U2144 ( .A(n3905), .B(n2664), .C(n3803), .D(n2663), .Z(n2137) );
  COND2X1 U2145 ( .A(n3904), .B(n2665), .C(n3803), .D(n2664), .Z(n2138) );
  COND2X1 U2147 ( .A(n3953), .B(n2667), .C(n3803), .D(n2666), .Z(n2140) );
  COND2X1 U2148 ( .A(n3904), .B(n2668), .C(n3803), .D(n2667), .Z(n2141) );
  COND2X1 U2150 ( .A(n3953), .B(n3483), .C(n3803), .D(n2669), .Z(n2143) );
  COND2X1 U2153 ( .A(n3953), .B(n2673), .C(n3803), .D(n2672), .Z(n2146) );
  COND2X1 U2154 ( .A(n3905), .B(n2674), .C(n3803), .D(n2673), .Z(n2147) );
  COND2X1 U2156 ( .A(n3905), .B(n2676), .C(n3803), .D(n2675), .Z(n2149) );
  COND2X1 U2200 ( .A(n27), .B(n2686), .C(n3931), .D(n2685), .Z(n2159) );
  COND2X1 U2201 ( .A(n27), .B(n2687), .C(n3930), .D(n2686), .Z(n2160) );
  COND2X1 U2202 ( .A(n27), .B(n2688), .C(n3931), .D(n2687), .Z(n2161) );
  COND2X1 U2203 ( .A(n27), .B(n2689), .C(n3931), .D(n2688), .Z(n2162) );
  COND2X1 U2204 ( .A(n27), .B(n2690), .C(n3931), .D(n2689), .Z(n2163) );
  COND2X1 U2205 ( .A(n27), .B(n2691), .C(n3930), .D(n2690), .Z(n2164) );
  COND2X1 U2206 ( .A(n27), .B(n2692), .C(n3930), .D(n2691), .Z(n2165) );
  COND2X1 U2209 ( .A(n27), .B(n2695), .C(n3931), .D(n2694), .Z(n2168) );
  COND2X1 U2210 ( .A(n27), .B(n2696), .C(n3931), .D(n2695), .Z(n2169) );
  COND2X1 U2211 ( .A(n3885), .B(n2697), .C(n3931), .D(n2696), .Z(n2170) );
  COND2X1 U2212 ( .A(n27), .B(n2698), .C(n3930), .D(n2697), .Z(n2171) );
  COND2X1 U2213 ( .A(n3885), .B(n2699), .C(n3548), .D(n2698), .Z(n2172) );
  COND2X1 U2214 ( .A(n3885), .B(n3108), .C(n3930), .D(n2699), .Z(n2173) );
  COND2X1 U2216 ( .A(n3885), .B(n2702), .C(n3548), .D(n2701), .Z(n2175) );
  COND2X1 U2220 ( .A(n27), .B(n2706), .C(n3931), .D(n2705), .Z(n2179) );
  COND2X1 U2221 ( .A(n3885), .B(n2707), .C(n3931), .D(n2706), .Z(n2180) );
  COND2X1 U2223 ( .A(n3885), .B(n2709), .C(n3548), .D(n2708), .Z(n2182) );
  COND2X1 U2263 ( .A(n2715), .B(n18), .C(n3934), .D(n2714), .Z(n2188) );
  COND2X1 U2265 ( .A(n18), .B(n2717), .C(n3933), .D(n2716), .Z(n2190) );
  COND2X1 U2266 ( .A(n3876), .B(n2718), .C(n3934), .D(n2717), .Z(n2191) );
  COND2X1 U2267 ( .A(n3876), .B(n2719), .C(n3933), .D(n2718), .Z(n2192) );
  COND2X1 U2268 ( .A(n18), .B(n2720), .C(n3933), .D(n2719), .Z(n2193) );
  COND2X1 U2269 ( .A(n3876), .B(n2721), .C(n3934), .D(n2720), .Z(n2194) );
  COND2X1 U2270 ( .A(n18), .B(n2722), .C(n3933), .D(n2721), .Z(n2195) );
  COND2X1 U2271 ( .A(n18), .B(n2723), .C(n3934), .D(n2722), .Z(n2196) );
  COND2X1 U2274 ( .A(n18), .B(n2726), .C(n3933), .D(n2725), .Z(n2199) );
  COND2X1 U2275 ( .A(n18), .B(n2727), .C(n3934), .D(n2726), .Z(n2200) );
  COND2X1 U2276 ( .A(n18), .B(n2728), .C(n3934), .D(n2727), .Z(n2201) );
  COND2X1 U2277 ( .A(n18), .B(n2729), .C(n3934), .D(n2728), .Z(n2202) );
  COND2X1 U2279 ( .A(n18), .B(n2731), .C(n3933), .D(n2730), .Z(n2204) );
  COND2X1 U2280 ( .A(n3876), .B(n2732), .C(n3933), .D(n2731), .Z(n2205) );
  COND2X1 U2281 ( .A(n3876), .B(n2733), .C(n3934), .D(n2732), .Z(n2206) );
  COND2X1 U2283 ( .A(n3876), .B(n2735), .C(n3934), .D(n2734), .Z(n2208) );
  COND2X1 U2285 ( .A(n18), .B(n2737), .C(n3934), .D(n2736), .Z(n2210) );
  COND2X1 U2286 ( .A(n3876), .B(n2738), .C(n3934), .D(n2737), .Z(n2211) );
  COND2X1 U2288 ( .A(n3876), .B(n2740), .C(n3934), .D(n2739), .Z(n2213) );
  COND2X1 U2289 ( .A(n18), .B(n2741), .C(n3933), .D(n2740), .Z(n2214) );
  COND2X1 U2292 ( .A(n3876), .B(n2744), .C(n3934), .D(n2743), .Z(n2217) );
  COND2X1 U2330 ( .A(n2748), .B(n3755), .C(n6), .D(n2747), .Z(n2221) );
  COND2X1 U2332 ( .A(n3880), .B(n2750), .C(n6), .D(n2749), .Z(n2223) );
  COND2X1 U2333 ( .A(n3783), .B(n2751), .C(n6), .D(n2750), .Z(n2224) );
  COND2X1 U2334 ( .A(n3754), .B(n2752), .C(n6), .D(n2751), .Z(n2225) );
  COND2X1 U2336 ( .A(n3880), .B(n2754), .C(n6), .D(n2753), .Z(n2227) );
  COND2X1 U2337 ( .A(n3880), .B(n2755), .C(n6), .D(n2754), .Z(n2228) );
  COND2X1 U2340 ( .A(n3880), .B(n2758), .C(n6), .D(n2757), .Z(n2231) );
  COND2X1 U2342 ( .A(n3880), .B(n2760), .C(n6), .D(n2759), .Z(n2233) );
  COND2X1 U2344 ( .A(n3880), .B(n2762), .C(n6), .D(n2761), .Z(n2235) );
  COND2X1 U2347 ( .A(n3880), .B(n2765), .C(n6), .D(n2764), .Z(n2238) );
  COND2X1 U2350 ( .A(n3880), .B(n2768), .C(n6), .D(n2767), .Z(n2241) );
  COND2X1 U2352 ( .A(n3880), .B(n2770), .C(n6), .D(n2769), .Z(n2243) );
  COND2X1 U2355 ( .A(n3880), .B(n2773), .C(n6), .D(n2772), .Z(n2246) );
  COND2X1 U2356 ( .A(n3880), .B(n2774), .C(n6), .D(n2773), .Z(n2247) );
  COND2X1 U2358 ( .A(n3880), .B(n2776), .C(n6), .D(n2775), .Z(n2249) );
  COND2X1 U2360 ( .A(n2778), .B(n3880), .C(n6), .D(n2777), .Z(n2251) );
  COND2X1 U1341 ( .A(n144), .B(n2269), .C(n3114), .D(n2268), .Z(n1755) );
  COND2X1 U1343 ( .A(n144), .B(n2271), .C(n3086), .D(n2270), .Z(n1757) );
  CND2X2 U400 ( .A(n923), .B(n938), .Z(n410) );
  CND2X2 U333 ( .A(n438), .B(n359), .Z(n353) );
  CNR2X2 U181 ( .A(n274), .B(n3225), .Z(n233) );
  COND1X1 U182 ( .A(n3225), .B(n275), .C(n3378), .Z(n236) );
  CNR2X2 U347 ( .A(n878), .B(n867), .Z(n369) );
  CNR2X2 U359 ( .A(n879), .B(n892), .Z(n378) );
  CNR2X2 U339 ( .A(n389), .B(n3251), .Z(n363) );
  CFA1X1 U861 ( .A(n1803), .B(n805), .CI(n808), .CO(n802), .S(n803) );
  CFA1X1 U862 ( .A(n810), .B(n1773), .CI(n1742), .CO(n804), .S(n805) );
  CFA1X1 U859 ( .A(n1772), .B(n804), .CI(n801), .CO(n798), .S(n799) );
  CANR1X1 U188 ( .A(net20956), .B(n253), .C(n244), .Z(n242) );
  COND2X1 U1863 ( .A(net21353), .B(n2519), .C(net19216), .D(n2518), .Z(n1993)
         );
  COND2X1 U1861 ( .A(n2517), .B(net21352), .C(net19216), .D(n2516), .Z(n1991)
         );
  COND2X1 U1342 ( .A(n144), .B(n2270), .C(n3173), .D(n2269), .Z(n1756) );
  CFA1X1 U946 ( .A(n1992), .B(n1756), .CI(n992), .CO(n972), .S(n973) );
  CFA1X1 U922 ( .A(n944), .B(n942), .CI(n929), .CO(n924), .S(n925) );
  CNR2X2 U375 ( .A(n893), .B(n906), .Z(n389) );
  COND2X1 U1472 ( .A(net21696), .B(n2332), .C(net22007), .D(n2331), .Z(n1815)
         );
  CFA1X1 U941 ( .A(n971), .B(n984), .CI(n973), .CO(n962), .S(n963) );
  CFA1X1 U945 ( .A(n1903), .B(n1786), .CI(n1815), .CO(n970), .S(n971) );
  COND2X1 U1602 ( .A(n108), .B(n2394), .C(net21250), .D(n2393), .Z(n1873) );
  CFA1X1 U942 ( .A(n988), .B(n969), .CI(n986), .CO(n964), .S(n965) );
  CFA1X1 U944 ( .A(n1873), .B(n1843), .CI(n1933), .CO(n968), .S(n969) );
  CFA1X1 U931 ( .A(n966), .B(n947), .CI(n964), .CO(n942), .S(n943) );
  CFA1X1 U933 ( .A(n972), .B(n970), .CI(n968), .CO(n946), .S(n947) );
  CFA1X1 U923 ( .A(n937), .B(n931), .CI(n946), .CO(n926), .S(n927) );
  COND2X1 U1599 ( .A(n108), .B(n2391), .C(net21250), .D(n2390), .Z(n1871) );
  CFA1X1 U909 ( .A(n918), .B(n903), .CI(n916), .CO(n898), .S(n899) );
  COND2X1 U1535 ( .A(net21312), .B(n2361), .C(net21512), .D(n2360), .Z(n1841)
         );
  COND2X1 U1730 ( .A(net21801), .B(n2454), .C(n87), .D(n2453), .Z(n1931) );
  COND2X1 U1665 ( .A(net21344), .B(n2423), .C(net21744), .D(n2422), .Z(n1901)
         );
  CFA1X1 U924 ( .A(n948), .B(n935), .CI(n933), .CO(n928), .S(n929) );
  CFA1X1 U926 ( .A(n1841), .B(n1931), .CI(n1901), .CO(n932), .S(n933) );
  CFA1X1 U916 ( .A(n934), .B(n917), .CI(n932), .CO(n912), .S(n913) );
  CFA1X1 U913 ( .A(n911), .B(n909), .CI(n924), .CO(n906), .S(n907) );
  CFA1X1 U914 ( .A(n928), .B(n926), .CI(n913), .CO(n908), .S(n909) );
  CFA1X1 U880 ( .A(n1777), .B(n1865), .CI(n1747), .CO(n840), .S(n841) );
  CFA1X1 U877 ( .A(n839), .B(n837), .CI(n846), .CO(n834), .S(n835) );
  CFA1X1 U878 ( .A(n850), .B(n848), .CI(n841), .CO(n836), .S(n837) );
  CFA1X1 U873 ( .A(n838), .B(n829), .CI(n836), .CO(n826), .S(n827) );
  CIVXL U2507 ( .A(n3326), .Z(n3022) );
  CIVXL U2508 ( .A(n3022), .Z(n3023) );
  CEOX1 U2509 ( .A(n3181), .B(n1212), .Z(n1175) );
  CND2XL U2510 ( .A(n1212), .B(n2093), .Z(n3183) );
  CIVX1 U2511 ( .A(n469), .Z(n467) );
  CENX2 U2512 ( .A(n3338), .B(n1017), .Z(n1015) );
  CND2X2 U2513 ( .A(n3350), .B(n3351), .Z(n3358) );
  CIVXL U2514 ( .A(net22050), .Z(n3024) );
  CIVX2 U2515 ( .A(net22626), .Z(net22050) );
  COND1X2 U2516 ( .A(n633), .B(n637), .C(n634), .Z(n632) );
  CIVXL U2517 ( .A(n963), .Z(n3308) );
  CEOX2 U2518 ( .A(a[20]), .B(n4002), .Z(n2817) );
  CEOX1 U2519 ( .A(n2096), .B(n2220), .Z(n3025) );
  CEOX2 U2520 ( .A(n3025), .B(n1302), .Z(n1263) );
  CND2X1 U2521 ( .A(n1302), .B(n2220), .Z(n3026) );
  CND2X1 U2522 ( .A(n1302), .B(n2096), .Z(n3027) );
  CND2XL U2523 ( .A(n2220), .B(n2096), .Z(n3028) );
  CND3X1 U2524 ( .A(n3026), .B(n3027), .C(n3028), .Z(n1262) );
  CIVXL U2525 ( .A(n3088), .Z(n3029) );
  CEOX2 U2526 ( .A(n1125), .B(n1146), .Z(n3030) );
  CEOX1 U2527 ( .A(n3030), .B(n1121), .Z(n1115) );
  CND2X1 U2528 ( .A(n1121), .B(n1146), .Z(n3031) );
  CND2X1 U2529 ( .A(n1121), .B(n1125), .Z(n3032) );
  CND2XL U2530 ( .A(n1146), .B(n1125), .Z(n3033) );
  CND3X2 U2531 ( .A(n3031), .B(n3032), .C(n3033), .Z(n1114) );
  CND2X1 U2532 ( .A(n1114), .B(n1093), .Z(n3191) );
  CEOX1 U2533 ( .A(n3958), .B(n3024), .Z(n2476) );
  CIVXL U2534 ( .A(n660), .Z(n778) );
  CND2X1 U2535 ( .A(n3798), .B(n2819), .Z(n3344) );
  CND2X4 U2536 ( .A(n3798), .B(n2819), .Z(n3871) );
  COND2X2 U2537 ( .A(n27), .B(n2685), .C(n3930), .D(n2684), .Z(n2158) );
  CENXL U2538 ( .A(n2798), .B(net21836), .Z(n2468) );
  CENXL U2539 ( .A(n3969), .B(net21836), .Z(n2463) );
  CND2X1 U2540 ( .A(n927), .B(n3035), .Z(n3036) );
  CND2X1 U2541 ( .A(n3034), .B(n940), .Z(n3037) );
  CND2X2 U2542 ( .A(n3036), .B(n3037), .Z(net22301) );
  CIVXL U2543 ( .A(n927), .Z(n3034) );
  CIVX2 U2544 ( .A(n940), .Z(n3035) );
  COND2XL U2545 ( .A(n45), .B(n2628), .C(n3939), .D(n2627), .Z(n2101) );
  CAOR1XL U2546 ( .A(n3938), .B(n45), .C(n2615), .Z(n2088) );
  COND2XL U2547 ( .A(n45), .B(n2632), .C(n3938), .D(n2631), .Z(n2105) );
  COND2XL U2548 ( .A(n45), .B(n2631), .C(n3938), .D(n2630), .Z(n2104) );
  COND2XL U2549 ( .A(n45), .B(n2641), .C(n3938), .D(n2640), .Z(n2114) );
  CNIVX3 U2550 ( .A(n42), .Z(n3939) );
  CIVXL U2551 ( .A(n1252), .Z(n3038) );
  CIVXL U2552 ( .A(n3038), .Z(n3039) );
  CEOX2 U2553 ( .A(n1259), .B(n1257), .Z(n3040) );
  CEOX2 U2554 ( .A(n3040), .B(n1284), .Z(n1251) );
  CND2X1 U2555 ( .A(n1284), .B(n1257), .Z(n3041) );
  CND2X1 U2556 ( .A(n1284), .B(n1259), .Z(n3042) );
  CND2XL U2557 ( .A(n1257), .B(n1259), .Z(n3043) );
  CND3X1 U2558 ( .A(n3041), .B(n3042), .C(n3043), .Z(n1250) );
  CNIVXL U2559 ( .A(n2439), .Z(n3044) );
  CIVX2 U2560 ( .A(n1250), .Z(n3136) );
  CNIVX2 U2561 ( .A(n1278), .Z(n3045) );
  CENX1 U2562 ( .A(n2783), .B(n3984), .Z(n2717) );
  CND2X1 U2563 ( .A(net21419), .B(n3047), .Z(n3048) );
  CND2X2 U2564 ( .A(n3046), .B(a[28]), .Z(n3049) );
  CND2X4 U2565 ( .A(n3048), .B(n3049), .Z(n2813) );
  CIVX2 U2566 ( .A(net21419), .Z(n3046) );
  CIVXL U2567 ( .A(a[28]), .Z(n3047) );
  CIVX2 U2568 ( .A(n3380), .Z(net21419) );
  CND2X4 U2569 ( .A(n2813), .B(net19191), .Z(net21434) );
  COR2X1 U2570 ( .A(n90), .B(n2475), .Z(n3050) );
  COR2X1 U2571 ( .A(net21846), .B(n2474), .Z(n3051) );
  CND2X2 U2572 ( .A(n3050), .B(n3051), .Z(n1950) );
  CEOX2 U2573 ( .A(n3998), .B(a[16]), .Z(n3756) );
  CENX1 U2574 ( .A(n3966), .B(n3998), .Z(n2499) );
  CENX2 U2575 ( .A(n1318), .B(n1291), .Z(n3334) );
  CND2X1 U2576 ( .A(n3271), .B(n3272), .Z(n3052) );
  CNIVXL U2577 ( .A(n1447), .Z(n3053) );
  CEO3X1 U2578 ( .A(n1451), .B(n1474), .C(n1476), .Z(n1447) );
  CEOX2 U2579 ( .A(n912), .B(n899), .Z(n3054) );
  CEOX2 U2580 ( .A(n3054), .B(n910), .Z(n895) );
  CND2X1 U2581 ( .A(n910), .B(n899), .Z(n3055) );
  CND2X1 U2582 ( .A(n910), .B(n912), .Z(n3056) );
  CND2XL U2583 ( .A(n899), .B(n912), .Z(n3057) );
  CND3X2 U2584 ( .A(n3055), .B(n3056), .C(n3057), .Z(n894) );
  CND2XL U2585 ( .A(n894), .B(n883), .Z(n3179) );
  CND2XL U2586 ( .A(n895), .B(n897), .Z(n3122) );
  CAOR1XL U2587 ( .A(n3660), .B(n63), .C(n2549), .Z(n2022) );
  CND3X1 U2588 ( .A(n3524), .B(n3525), .C(n3526), .Z(n1220) );
  CIVXL U2589 ( .A(n992), .Z(n993) );
  CENX4 U2590 ( .A(n3957), .B(net19314), .Z(n2477) );
  CENX1 U2591 ( .A(n3968), .B(net21910), .Z(n2299) );
  COR2X1 U2592 ( .A(n3871), .B(n2501), .Z(n3458) );
  CEO3X2 U2593 ( .A(n1288), .B(n1261), .C(n1286), .Z(n1253) );
  CNIVX4 U2594 ( .A(n4002), .Z(n3926) );
  CIVX2 U2595 ( .A(n3140), .Z(n4002) );
  CEOX2 U2596 ( .A(n1255), .B(n1282), .Z(n3058) );
  CEOX2 U2597 ( .A(n3058), .B(n1280), .Z(n1249) );
  CND2X1 U2598 ( .A(n1280), .B(n1282), .Z(n3059) );
  CND2X1 U2599 ( .A(n1280), .B(n1255), .Z(n3060) );
  CND2X1 U2600 ( .A(n1282), .B(n1255), .Z(n3061) );
  CND3X2 U2601 ( .A(n3059), .B(n3060), .C(n3061), .Z(n1248) );
  CND3X1 U2602 ( .A(n3809), .B(n3810), .C(n3811), .Z(n1282) );
  CIVX2 U2603 ( .A(n1248), .Z(n3670) );
  CNR2X2 U2604 ( .A(n3599), .B(n491), .Z(n3062) );
  CNR2X1 U2605 ( .A(n3599), .B(n491), .Z(n3063) );
  CNR2XL U2606 ( .A(n3599), .B(n491), .Z(n482) );
  CNR2X2 U2607 ( .A(n1693), .B(n1700), .Z(n696) );
  CFA1X1 U2608 ( .A(n2243), .B(n2181), .CI(n1735), .CO(n1696), .S(n1697) );
  COND2X1 U2609 ( .A(n3787), .B(n3995), .C(n3939), .D(n2647), .Z(n1735) );
  CIVX1 U2610 ( .A(n369), .Z(n744) );
  CIVX1 U2611 ( .A(n978), .Z(n3310) );
  CIVX2 U2612 ( .A(n69), .Z(n3376) );
  COND2XL U2613 ( .A(n27), .B(n2710), .C(n3931), .D(n2709), .Z(n2183) );
  COND2XL U2614 ( .A(n27), .B(n2711), .C(n3930), .D(n2710), .Z(n2184) );
  CAOR1XL U2615 ( .A(n3931), .B(n27), .C(n2681), .Z(n2154) );
  CNIVX1 U2616 ( .A(n1445), .Z(n3064) );
  CIVX2 U2617 ( .A(n81), .Z(n3367) );
  CND2X1 U2618 ( .A(n1375), .B(n1396), .Z(n3209) );
  COND2XL U2619 ( .A(net21434), .B(n3424), .C(net19193), .D(n2303), .Z(n1789)
         );
  CND2X1 U2620 ( .A(n1373), .B(n1396), .Z(n3210) );
  CND2XL U2621 ( .A(n1409), .B(n1403), .Z(n3206) );
  CEOX1 U2622 ( .A(n3719), .B(n2012), .Z(n1499) );
  COND2XL U2623 ( .A(net21312), .B(n2367), .C(net21512), .D(n2366), .Z(n1847)
         );
  COND2XL U2624 ( .A(net21312), .B(n2366), .C(net21512), .D(n2365), .Z(n1846)
         );
  COND2X1 U2625 ( .A(net21311), .B(n2360), .C(net21512), .D(n2359), .Z(n920)
         );
  COND2X1 U2626 ( .A(n3904), .B(n2659), .C(n3803), .D(n2658), .Z(n2132) );
  CNR2X2 U2627 ( .A(n3067), .B(n594), .Z(n576) );
  CENX2 U2628 ( .A(n1324), .B(n3065), .Z(n1289) );
  CENX2 U2629 ( .A(n1326), .B(n1322), .Z(n3065) );
  CEO3X2 U2630 ( .A(n1487), .B(n1506), .C(n1485), .Z(n3499) );
  CENX1 U2631 ( .A(n1162), .B(n3288), .Z(n3066) );
  CENX1 U2632 ( .A(n1162), .B(n3288), .Z(n1135) );
  CND2X1 U2633 ( .A(n767), .B(n768), .Z(n3067) );
  CND2XL U2634 ( .A(n767), .B(n768), .Z(n3068) );
  CIVX3 U2635 ( .A(n591), .Z(n768) );
  CENXL U2636 ( .A(n3957), .B(n4005), .Z(n2345) );
  CIVX3 U2637 ( .A(n4007), .Z(n4005) );
  CENX1 U2638 ( .A(n3972), .B(n3984), .Z(n2723) );
  CND2X4 U2639 ( .A(n3936), .B(n2821), .Z(n3228) );
  CENX2 U2640 ( .A(n2785), .B(net19314), .Z(n2455) );
  CEO3X1 U2641 ( .A(n1005), .B(n1003), .C(n1022), .Z(n999) );
  CND2X1 U2642 ( .A(n1005), .B(n1003), .Z(n3069) );
  CND2XL U2643 ( .A(n1005), .B(n1022), .Z(n3070) );
  CND2X1 U2644 ( .A(n1003), .B(n1022), .Z(n3071) );
  CND3X2 U2645 ( .A(n3069), .B(n3070), .C(n3071), .Z(n998) );
  CEOX2 U2646 ( .A(n1000), .B(n981), .Z(n3072) );
  CEOX2 U2647 ( .A(n3072), .B(n998), .Z(n977) );
  CND2XL U2648 ( .A(n1000), .B(n981), .Z(n3073) );
  CND2XL U2649 ( .A(n1000), .B(n998), .Z(n3074) );
  CND2XL U2650 ( .A(n981), .B(n998), .Z(n3075) );
  CND3X1 U2651 ( .A(n3073), .B(n3074), .C(n3075), .Z(n976) );
  CEOX2 U2652 ( .A(n979), .B(n996), .Z(n3076) );
  CEOX2 U2653 ( .A(n3076), .B(n977), .Z(n975) );
  CND2XL U2654 ( .A(n977), .B(n996), .Z(n3077) );
  CND2X1 U2655 ( .A(n977), .B(n979), .Z(n3078) );
  CND2XL U2656 ( .A(n996), .B(n979), .Z(n3079) );
  CND3XL U2657 ( .A(n3077), .B(n3078), .C(n3079), .Z(n974) );
  CENX2 U2658 ( .A(n3956), .B(net19314), .Z(n2478) );
  CND2X1 U2659 ( .A(n1213), .B(n1205), .Z(n3082) );
  CND2X2 U2660 ( .A(n3080), .B(n3081), .Z(n3083) );
  CND2X2 U2661 ( .A(n3082), .B(n3083), .Z(n3408) );
  CIVX1 U2662 ( .A(n1213), .Z(n3080) );
  CIVX2 U2663 ( .A(n1205), .Z(n3081) );
  CANR1X2 U2664 ( .A(n478), .B(net22599), .C(n479), .Z(net19189) );
  CNIVX4 U2665 ( .A(n3864), .Z(n3895) );
  CNIVX4 U2666 ( .A(n48), .Z(n3084) );
  COND1X1 U2667 ( .A(n573), .B(n567), .C(n568), .Z(n562) );
  CENX1 U2668 ( .A(n3157), .B(n1363), .Z(n1361) );
  CENX1 U2669 ( .A(n1388), .B(n1365), .Z(n3157) );
  CENX1 U2670 ( .A(n3387), .B(n1018), .Z(n997) );
  CNR2IX1 U2671 ( .B(n3979), .A(n3173), .Z(n1770) );
  CIVX2 U2672 ( .A(n3113), .Z(n3085) );
  CIVX2 U2673 ( .A(n3113), .Z(n3086) );
  CIVX1 U2674 ( .A(n3113), .Z(net22439) );
  CIVX2 U2675 ( .A(n3997), .Z(n3996) );
  CND2X2 U2676 ( .A(n1258), .B(n3088), .Z(n3089) );
  CND2X1 U2677 ( .A(n3087), .B(n1256), .Z(n3090) );
  CND2X2 U2678 ( .A(n3089), .B(n3090), .Z(n3277) );
  CIVXL U2679 ( .A(n1258), .Z(n3087) );
  CIVX2 U2680 ( .A(n1256), .Z(n3088) );
  CIVX1 U2681 ( .A(net19062), .Z(n87) );
  CIVXL U2682 ( .A(net19062), .Z(net22327) );
  CIVXL U2683 ( .A(net19062), .Z(net22326) );
  CND2X4 U2684 ( .A(n2821), .B(n3660), .Z(n63) );
  CND3X2 U2685 ( .A(n3168), .B(n3169), .C(n3170), .Z(n1288) );
  CENX1 U2686 ( .A(n3973), .B(n3924), .Z(n2590) );
  CND3X1 U2687 ( .A(n3799), .B(n3800), .C(n3801), .Z(n1082) );
  CND2X2 U2688 ( .A(n2823), .B(n3937), .Z(n3787) );
  CND2XL U2689 ( .A(n3966), .B(net21836), .Z(n3093) );
  CND2X2 U2690 ( .A(n3091), .B(n3092), .Z(n3094) );
  CND2X1 U2691 ( .A(n3093), .B(n3094), .Z(n2466) );
  CIVXL U2692 ( .A(n3966), .Z(n3091) );
  CIVX2 U2693 ( .A(net21836), .Z(n3092) );
  CENX2 U2694 ( .A(n1289), .B(n1314), .Z(n3509) );
  COND1X2 U2695 ( .A(n559), .B(n551), .C(n552), .Z(n550) );
  CENX1 U2696 ( .A(n3973), .B(n3984), .Z(n2722) );
  CIVXL U2697 ( .A(n396), .Z(n3095) );
  CIVXL U2698 ( .A(n3095), .Z(n3096) );
  CENX2 U2699 ( .A(n3097), .B(n881), .Z(n3177) );
  CIVX20 U2700 ( .A(n883), .Z(n3097) );
  CENX2 U2701 ( .A(a[20]), .B(net22626), .Z(n3373) );
  CND2X2 U2702 ( .A(n1245), .B(n1274), .Z(n544) );
  COND2XL U2703 ( .A(n126), .B(n3863), .C(net22007), .D(n2350), .Z(n1726) );
  COND2XL U2704 ( .A(n2349), .B(n126), .C(net22007), .D(n2348), .Z(n1832) );
  CENX1 U2705 ( .A(n3976), .B(n3984), .Z(n2718) );
  CND2X2 U2706 ( .A(n1317), .B(n1319), .Z(n3589) );
  CEO3XL U2707 ( .A(n1645), .B(n1643), .C(n1654), .Z(n3098) );
  CEOX1 U2708 ( .A(n3961), .B(n3235), .Z(n2638) );
  CIVX1 U2709 ( .A(n3234), .Z(n3235) );
  CEO3XL U2710 ( .A(n1631), .B(n1629), .C(n1642), .Z(n3099) );
  COND1X1 U2711 ( .A(n628), .B(n622), .C(n623), .Z(n621) );
  CIVXL U2712 ( .A(n628), .Z(n626) );
  CND2X1 U2713 ( .A(n3101), .B(n1544), .Z(n628) );
  CANR1X1 U2714 ( .A(n669), .B(n677), .C(n670), .Z(n3264) );
  COR2X1 U2715 ( .A(n1612), .B(n1597), .Z(n3100) );
  COR2XL U2716 ( .A(n1612), .B(n1597), .Z(n3911) );
  CEO3XL U2717 ( .A(n1529), .B(n1527), .C(n1546), .Z(n3101) );
  CIVXL U2718 ( .A(n3882), .Z(n3102) );
  COND2X1 U2719 ( .A(net21801), .B(net21791), .C(net21846), .D(n2482), .Z(
        n1730) );
  CNIVX2 U2720 ( .A(n2148), .Z(n3103) );
  CENXL U2721 ( .A(n3957), .B(n3991), .Z(n2675) );
  CNIVX1 U2722 ( .A(n2240), .Z(n3104) );
  CIVX1 U2723 ( .A(n2178), .Z(n3105) );
  CIVX2 U2724 ( .A(n3105), .Z(n3106) );
  CENX2 U2725 ( .A(n1443), .B(n3107), .Z(n1439) );
  CENX1 U2726 ( .A(n1466), .B(n1464), .Z(n3107) );
  CNIVXL U2727 ( .A(n2700), .Z(n3108) );
  CND2X1 U2728 ( .A(n1591), .B(n1606), .Z(n3556) );
  CENX1 U2729 ( .A(n3968), .B(n3923), .Z(n2596) );
  CENXL U2730 ( .A(n3970), .B(n3923), .Z(n2593) );
  CND2X1 U2731 ( .A(n51), .B(n2822), .Z(n3806) );
  CIVX4 U2732 ( .A(n3922), .Z(n3932) );
  CENXL U2733 ( .A(n569), .B(n3109), .Z(product[29]) );
  CAN2X2 U2734 ( .A(n765), .B(n568), .Z(n3109) );
  CIVXL U2735 ( .A(net22598), .Z(n3110) );
  CNR2X2 U2736 ( .A(n1387), .B(n1412), .Z(n3886) );
  CNIVX2 U2737 ( .A(n1113), .Z(n3111) );
  CNIVX16 U2738 ( .A(n4003), .Z(n3925) );
  CND2X1 U2739 ( .A(n1339), .B(n1364), .Z(n3404) );
  COND2X1 U2740 ( .A(n54), .B(n2589), .C(n3453), .D(n2588), .Z(n2062) );
  CND2X4 U2741 ( .A(n3472), .B(n3473), .Z(n2822) );
  CND2X2 U2742 ( .A(n3470), .B(a[10]), .Z(n3473) );
  CND2X2 U2743 ( .A(n1059), .B(n1082), .Z(n485) );
  CANR1XL U2744 ( .A(n520), .B(n535), .C(n3023), .Z(n3898) );
  CEO3X1 U2745 ( .A(n1732), .B(n2144), .C(n2237), .Z(n1637) );
  CNIVX1 U2746 ( .A(n1462), .Z(n3112) );
  CENX1 U2747 ( .A(n1462), .B(n1441), .Z(n3462) );
  COND1XL U2748 ( .A(n547), .B(n575), .C(n548), .Z(n3817) );
  COND1X1 U2749 ( .A(n547), .B(n575), .C(n548), .Z(net22598) );
  CIVXL U2750 ( .A(n3565), .Z(n1243) );
  CIVX1 U2751 ( .A(n3955), .Z(n3453) );
  CND2XL U2752 ( .A(n2103), .B(n2041), .Z(n3445) );
  COND2X1 U2753 ( .A(n144), .B(n2279), .C(n3173), .D(n2278), .Z(n1765) );
  CIVDX2 U2754 ( .A(n141), .Z0(n3113), .Z1(n3114) );
  CND2X4 U2755 ( .A(n2812), .B(n3331), .Z(n144) );
  CENX1 U2756 ( .A(n3956), .B(net21910), .Z(n3752) );
  CNIVXL U2757 ( .A(n1224), .Z(n3115) );
  CEO3XL U2758 ( .A(n1311), .B(n1313), .C(n3323), .Z(n1307) );
  CAN2X1 U2759 ( .A(n1167), .B(n3347), .Z(n3116) );
  CND2X2 U2760 ( .A(n745), .B(n744), .Z(n3251) );
  CAN2X1 U2761 ( .A(n3315), .B(n3316), .Z(n3117) );
  CIVDXL U2762 ( .A(n460), .Z0(n3118), .Z1(n3119) );
  CIVX1 U2763 ( .A(n514), .Z(n516) );
  CEOX2 U2764 ( .A(n897), .B(n908), .Z(n3120) );
  CEOX2 U2765 ( .A(n3120), .B(n895), .Z(n893) );
  CND2X1 U2766 ( .A(n895), .B(n908), .Z(n3121) );
  CND2X1 U2767 ( .A(n908), .B(n897), .Z(n3123) );
  CND3X1 U2768 ( .A(n3121), .B(n3122), .C(n3123), .Z(n892) );
  CANR1X1 U2769 ( .A(n363), .B(n397), .C(n364), .Z(n3124) );
  CND2X1 U2770 ( .A(n893), .B(n906), .Z(n392) );
  CANR1X1 U2771 ( .A(n363), .B(n397), .C(n364), .Z(n362) );
  CEO3X1 U2772 ( .A(n1826), .B(n1854), .C(n2126), .Z(n1237) );
  CND2XL U2773 ( .A(n1826), .B(n2126), .Z(n3125) );
  CND2XL U2774 ( .A(n1826), .B(n1854), .Z(n3126) );
  CND2X1 U2775 ( .A(n2126), .B(n1854), .Z(n3127) );
  CND3X1 U2776 ( .A(n3125), .B(n3126), .C(n3127), .Z(n1236) );
  CIVX2 U2777 ( .A(net21859), .Z(n3128) );
  CIVX1 U2778 ( .A(net21859), .Z(n3129) );
  CIVX3 U2779 ( .A(net21859), .Z(net19081) );
  CEOX2 U2780 ( .A(n3504), .B(n1828), .Z(n1295) );
  CIVXL U2781 ( .A(n1199), .Z(n3130) );
  CIVXL U2782 ( .A(n3130), .Z(n3131) );
  CND2X1 U2783 ( .A(a[8]), .B(n30), .Z(n3134) );
  CND2X2 U2784 ( .A(n3132), .B(n3133), .Z(n3135) );
  CND2X2 U2785 ( .A(n3134), .B(n3135), .Z(n42) );
  CIVX2 U2786 ( .A(a[8]), .Z(n3132) );
  CIVX1 U2787 ( .A(n30), .Z(n3133) );
  CND2X1 U2788 ( .A(n1250), .B(n1221), .Z(n3138) );
  CND2X2 U2789 ( .A(n3136), .B(n3137), .Z(n3139) );
  CND2X2 U2790 ( .A(n3138), .B(n3139), .Z(n3685) );
  CIVX2 U2791 ( .A(n1221), .Z(n3137) );
  CND2X1 U2792 ( .A(n3685), .B(n1248), .Z(n3671) );
  CIVX2 U2793 ( .A(n3685), .Z(n3669) );
  CND2X1 U2794 ( .A(n3237), .B(n1198), .Z(n3706) );
  CIVX1 U2795 ( .A(n93), .Z(n3140) );
  CND3X1 U2796 ( .A(n3828), .B(n3829), .C(n3830), .Z(n3141) );
  CND3XL U2797 ( .A(n3828), .B(n3829), .C(n3830), .Z(n1132) );
  CEOXL U2798 ( .A(n1225), .B(n1223), .Z(n3793) );
  CND2X1 U2799 ( .A(n1443), .B(n1464), .Z(n3142) );
  CND2X1 U2800 ( .A(n1443), .B(n1466), .Z(n3143) );
  CND2X1 U2801 ( .A(n1464), .B(n1466), .Z(n3144) );
  CND3X2 U2802 ( .A(n3142), .B(n3143), .C(n3144), .Z(n1438) );
  CNIVX1 U2803 ( .A(n1438), .Z(n3230) );
  CIVX3 U2804 ( .A(n3129), .Z(net21684) );
  CEOX1 U2805 ( .A(n2003), .B(n1884), .Z(n3591) );
  COND2XL U2806 ( .A(n144), .B(n2260), .C(n3085), .D(n2259), .Z(n1746) );
  CIVXL U2807 ( .A(n800), .Z(n801) );
  CEOXL U2808 ( .A(n1842), .B(n1755), .Z(n3151) );
  CND2XL U2809 ( .A(n1991), .B(n1755), .Z(n3152) );
  CENXL U2810 ( .A(n1869), .B(n1751), .Z(n3172) );
  CIVX2 U2811 ( .A(n102), .Z(net19171) );
  CIVX4 U2812 ( .A(n3955), .Z(n3145) );
  CIVX3 U2813 ( .A(n3955), .Z(n51) );
  CENX2 U2814 ( .A(n2810), .B(net19268), .Z(n2381) );
  CND2XL U2815 ( .A(n1167), .B(n1194), .Z(n3356) );
  CND2XL U2816 ( .A(n3331), .B(n2812), .Z(net21320) );
  COND2X2 U2817 ( .A(n3904), .B(n2662), .C(n3803), .D(n2661), .Z(n2135) );
  CIVXL U2818 ( .A(n501), .Z(n3146) );
  CEOX2 U2819 ( .A(n3401), .B(n1364), .Z(n1335) );
  CEOX1 U2820 ( .A(n1117), .B(n1140), .Z(n3147) );
  CEOX1 U2821 ( .A(n3147), .B(n1115), .Z(n1111) );
  CND2X1 U2822 ( .A(n1115), .B(n1140), .Z(n3148) );
  CND2X1 U2823 ( .A(n1115), .B(n1117), .Z(n3149) );
  CND2XL U2824 ( .A(n1140), .B(n1117), .Z(n3150) );
  CND3X2 U2825 ( .A(n3148), .B(n3149), .C(n3150), .Z(n1110) );
  CEOX1 U2826 ( .A(n3151), .B(n1991), .Z(n953) );
  CND2XL U2827 ( .A(n1991), .B(n1842), .Z(n3153) );
  CND2XL U2828 ( .A(n1755), .B(n1842), .Z(n3154) );
  CND3X1 U2829 ( .A(n3152), .B(n3153), .C(n3154), .Z(n952) );
  CIVX8 U2830 ( .A(n3935), .Z(n3660) );
  CEOX2 U2831 ( .A(n1309), .B(n1334), .Z(n3652) );
  CND3X2 U2832 ( .A(n3402), .B(n3403), .C(n3404), .Z(n1334) );
  CND3X2 U2833 ( .A(n3596), .B(n3597), .C(n3598), .Z(n1280) );
  CND2X1 U2834 ( .A(n1314), .B(n1289), .Z(n3598) );
  CND3X2 U2835 ( .A(n3738), .B(n3739), .C(n3740), .Z(n1314) );
  CND2X1 U2836 ( .A(n1325), .B(n1348), .Z(n3739) );
  COND2XL U2837 ( .A(n3876), .B(n2724), .C(n3934), .D(n2723), .Z(n2197) );
  CIVX1 U2838 ( .A(n3833), .Z(n3441) );
  CENXL U2839 ( .A(n2785), .B(n3993), .Z(n3155) );
  CENX1 U2840 ( .A(n3971), .B(net21909), .Z(n2295) );
  CENXL U2841 ( .A(n3975), .B(n3993), .Z(n3156) );
  CIVXL U2842 ( .A(net22050), .Z(n3158) );
  CEOX1 U2843 ( .A(n1241), .B(n1237), .Z(n3624) );
  CIVX3 U2844 ( .A(n3986), .Z(n3985) );
  CEOX2 U2845 ( .A(n1408), .B(n1406), .Z(n3159) );
  CEOX2 U2846 ( .A(n3159), .B(n1385), .Z(n1373) );
  CND2X1 U2847 ( .A(n1385), .B(n1406), .Z(n3160) );
  CND2X1 U2848 ( .A(n1385), .B(n1408), .Z(n3161) );
  CND2X1 U2849 ( .A(n1406), .B(n1408), .Z(n3162) );
  CND3X1 U2850 ( .A(n3160), .B(n3161), .C(n3162), .Z(n1372) );
  CEOX2 U2851 ( .A(n1007), .B(n1026), .Z(n3163) );
  CEOX2 U2852 ( .A(n3163), .B(n1024), .Z(n1001) );
  CND2XL U2853 ( .A(n1024), .B(n1026), .Z(n3164) );
  CND2X1 U2854 ( .A(n1024), .B(n1007), .Z(n3165) );
  CND2XL U2855 ( .A(n1026), .B(n1007), .Z(n3166) );
  CND3X1 U2856 ( .A(n3164), .B(n3165), .C(n3166), .Z(n1000) );
  CENX1 U2857 ( .A(n1020), .B(n1001), .Z(n3387) );
  CIVXL U2858 ( .A(n4003), .Z(n3167) );
  CIVX2 U2859 ( .A(n1165), .Z(n3186) );
  CND2X1 U2860 ( .A(n1324), .B(n1322), .Z(n3168) );
  CND2X1 U2861 ( .A(n1324), .B(n1326), .Z(n3169) );
  CND2X1 U2862 ( .A(n1322), .B(n1326), .Z(n3170) );
  CENX1 U2863 ( .A(n3171), .B(n1195), .Z(n1191) );
  CENX1 U2864 ( .A(n1197), .B(n1222), .Z(n3171) );
  CENX1 U2865 ( .A(n3172), .B(n1898), .Z(n887) );
  CND2X1 U2866 ( .A(n3349), .B(n3361), .Z(n3352) );
  CND2X4 U2867 ( .A(n3807), .B(n3808), .Z(n3869) );
  CIVX8 U2868 ( .A(net22004), .Z(net22006) );
  CIVXL U2869 ( .A(n572), .Z(n766) );
  CENXL U2870 ( .A(n3964), .B(net19309), .Z(n2536) );
  CND2X1 U2871 ( .A(n1203), .B(n1228), .Z(n3283) );
  CNR2IXL U2872 ( .B(n1194), .A(n1169), .Z(n3361) );
  CIVX1 U2873 ( .A(net19171), .Z(net21177) );
  CNIVX4 U2874 ( .A(n141), .Z(n3173) );
  CND2X2 U2875 ( .A(n3174), .B(n3175), .Z(n3176) );
  CND2X2 U2876 ( .A(n3556), .B(n3176), .Z(n3368) );
  CIVXL U2877 ( .A(n1606), .Z(n3174) );
  CIVX2 U2878 ( .A(n1591), .Z(n3175) );
  CENX2 U2879 ( .A(n1337), .B(n1362), .Z(n3337) );
  CENX1 U2880 ( .A(a[14]), .B(n57), .Z(n69) );
  CEOX2 U2881 ( .A(n3177), .B(n894), .Z(n879) );
  CND2XL U2882 ( .A(n894), .B(n881), .Z(n3178) );
  CND2XL U2883 ( .A(n881), .B(n883), .Z(n3180) );
  CND3X1 U2884 ( .A(n3178), .B(n3179), .C(n3180), .Z(n878) );
  CND2X1 U2885 ( .A(n1251), .B(n1253), .Z(n3681) );
  CENXL U2886 ( .A(n3967), .B(n3985), .Z(n2729) );
  CENXL U2887 ( .A(n3966), .B(n3985), .Z(n2730) );
  CEOX2 U2888 ( .A(n2093), .B(n1185), .Z(n3181) );
  CND2XL U2889 ( .A(n1212), .B(n1185), .Z(n3182) );
  CND2XL U2890 ( .A(n1185), .B(n2093), .Z(n3184) );
  CND3X1 U2891 ( .A(n3182), .B(n3183), .C(n3184), .Z(n1174) );
  CENX2 U2892 ( .A(net18979), .B(net21836), .Z(n2467) );
  CIVX2 U2893 ( .A(net19068), .Z(net21835) );
  CND2X2 U2894 ( .A(n1192), .B(n3186), .Z(n3187) );
  CND2X1 U2895 ( .A(n3185), .B(n1165), .Z(n3188) );
  CND2X2 U2896 ( .A(n3187), .B(n3188), .Z(n3613) );
  CIVXL U2897 ( .A(n1192), .Z(n3185) );
  CANR1X1 U2898 ( .A(n745), .B(n384), .C(n377), .Z(n373) );
  CFA1X1 U2899 ( .A(n1930), .B(n1871), .CI(n1783), .CO(n916), .S(n917) );
  COND2X1 U2900 ( .A(net21434), .B(n2298), .C(net19193), .D(n2297), .Z(n1783)
         );
  CND2X1 U2901 ( .A(n3331), .B(n2812), .Z(n3189) );
  CEO3X1 U2902 ( .A(n1114), .B(n1093), .C(n1091), .Z(n1087) );
  CND2X1 U2903 ( .A(n1114), .B(n1091), .Z(n3190) );
  CND2X2 U2904 ( .A(n1091), .B(n1093), .Z(n3192) );
  CND3X2 U2905 ( .A(n3190), .B(n3191), .C(n3192), .Z(n1086) );
  CND2X1 U2906 ( .A(n1086), .B(n1088), .Z(n3254) );
  CENXL U2907 ( .A(n3976), .B(n3926), .Z(n2421) );
  CND2X2 U2908 ( .A(n3193), .B(n3194), .Z(n3195) );
  CND2X2 U2909 ( .A(n3384), .B(n3195), .Z(n3333) );
  CIVXL U2910 ( .A(n999), .Z(n3193) );
  CIVX2 U2911 ( .A(n997), .Z(n3194) );
  CENX1 U2912 ( .A(n3333), .B(n1016), .Z(n995) );
  CND2X1 U2913 ( .A(n999), .B(n997), .Z(n3384) );
  CND2X1 U2914 ( .A(n3458), .B(n3459), .Z(n1975) );
  CEOX1 U2915 ( .A(n3977), .B(net22399), .Z(n2516) );
  CND3X1 U2916 ( .A(n3524), .B(n3525), .C(n3526), .Z(n3196) );
  COND2XL U2917 ( .A(n108), .B(n2400), .C(net21250), .D(n2399), .Z(n1878) );
  COND2X1 U2918 ( .A(n108), .B(n2412), .C(net21248), .D(n2411), .Z(n1890) );
  CNIVX2 U2919 ( .A(n24), .Z(n3929) );
  CNIVX2 U2920 ( .A(n24), .Z(n3930) );
  CNIVX3 U2921 ( .A(n24), .Z(n3931) );
  CIVXL U2922 ( .A(n1013), .Z(n3197) );
  CIVXL U2923 ( .A(n3197), .Z(n3198) );
  CIVXL U2924 ( .A(n399), .Z(n3199) );
  CENX1 U2925 ( .A(n3975), .B(n3926), .Z(n2423) );
  CEO3X1 U2926 ( .A(n1366), .B(n1343), .C(n1368), .Z(n1337) );
  CEOX2 U2927 ( .A(n943), .B(n958), .Z(n3200) );
  CEOX2 U2928 ( .A(n3200), .B(n941), .Z(n939) );
  CND2X1 U2929 ( .A(n941), .B(n958), .Z(n3201) );
  CND2X1 U2930 ( .A(n941), .B(n943), .Z(n3202) );
  CND2XL U2931 ( .A(n958), .B(n943), .Z(n3203) );
  CND3X1 U2932 ( .A(n3201), .B(n3202), .C(n3203), .Z(n938) );
  CND2X2 U2933 ( .A(n3307), .B(n3117), .Z(n958) );
  CEN3X2 U2934 ( .A(n1254), .B(n1229), .C(n3281), .Z(n1221) );
  CND2X4 U2935 ( .A(n3878), .B(n3936), .Z(n3550) );
  CIVDX2 U2936 ( .A(n472), .Z0(n3423), .Z1(n3422) );
  CIVX2 U2937 ( .A(a[26]), .Z(net21683) );
  CIVX2 U2938 ( .A(a[26]), .Z(net21693) );
  CEO3X1 U2939 ( .A(n1426), .B(n1409), .C(n1403), .Z(n1397) );
  CND2XL U2940 ( .A(n1426), .B(n1409), .Z(n3204) );
  CND2XL U2941 ( .A(n1426), .B(n1403), .Z(n3205) );
  CND3X1 U2942 ( .A(n3204), .B(n3205), .C(n3206), .Z(n1396) );
  CEOX2 U2943 ( .A(n1375), .B(n1373), .Z(n3207) );
  CEOX2 U2944 ( .A(n3207), .B(n1396), .Z(n1367) );
  CND2XL U2945 ( .A(n1375), .B(n1373), .Z(n3208) );
  CND3X1 U2946 ( .A(n3208), .B(n3209), .C(n3210), .Z(n1366) );
  CNIVX2 U2947 ( .A(n120), .Z(n3864) );
  CENXL U2948 ( .A(n2809), .B(net21909), .Z(n2314) );
  CENXL U2949 ( .A(n3964), .B(net21909), .Z(n2305) );
  CIVXL U2950 ( .A(n3213), .Z(n3211) );
  CAN2XL U2951 ( .A(net21375), .B(n2816), .Z(n3212) );
  CIVXL U2952 ( .A(n3167), .Z(n3213) );
  CENX2 U2953 ( .A(n1395), .B(n1393), .Z(n3692) );
  CNIVX4 U2954 ( .A(n3864), .Z(n3896) );
  CENXL U2955 ( .A(n2792), .B(net21909), .Z(n2297) );
  CEOX1 U2956 ( .A(n3624), .B(n1260), .Z(n1225) );
  CIVX2 U2957 ( .A(net18561), .Z(net22241) );
  CNIVX4 U2958 ( .A(n2799), .Z(n3965) );
  CNIVX4 U2959 ( .A(n2796), .Z(n3966) );
  CNIVX4 U2960 ( .A(n2803), .Z(n3961) );
  CND2X2 U2961 ( .A(n3683), .B(n3684), .Z(n2821) );
  CND2X1 U2962 ( .A(net22242), .B(n3682), .Z(n3683) );
  CNIVX8 U2963 ( .A(n2808), .Z(n3956) );
  CND2X1 U2964 ( .A(n3527), .B(n1479), .Z(n3530) );
  CENX1 U2965 ( .A(n2810), .B(net18483), .Z(n2282) );
  CENX1 U2966 ( .A(n3961), .B(net21910), .Z(n2308) );
  CENX1 U2967 ( .A(n3967), .B(n3925), .Z(n2432) );
  CENX1 U2968 ( .A(n3970), .B(net19314), .Z(n2461) );
  CENX1 U2969 ( .A(n3968), .B(n3925), .Z(n2431) );
  CENX1 U2970 ( .A(n2809), .B(net19314), .Z(n2479) );
  CIVX1 U2971 ( .A(n3959), .Z(n3508) );
  CND3X1 U2972 ( .A(n3607), .B(n3608), .C(n3609), .Z(n1428) );
  CENX1 U2973 ( .A(n2810), .B(net21910), .Z(n3758) );
  CENX1 U2974 ( .A(n3964), .B(net19314), .Z(n2470) );
  CENX1 U2975 ( .A(n2792), .B(n3923), .Z(n2594) );
  CENX1 U2976 ( .A(n3332), .B(n3158), .Z(n2469) );
  CIVX2 U2977 ( .A(n3965), .Z(n3332) );
  CIVX2 U2978 ( .A(n3376), .Z(net22248) );
  CIVX2 U2979 ( .A(n21), .Z(n3989) );
  CIVX3 U2980 ( .A(n3989), .Z(n3987) );
  CNIVX4 U2981 ( .A(n2789), .Z(n3972) );
  CENX1 U2982 ( .A(n3977), .B(net19314), .Z(n2450) );
  CNR2IX1 U2983 ( .B(n3979), .A(n3145), .Z(n2087) );
  CNR2IX1 U2984 ( .B(n3979), .A(net21248), .Z(n1894) );
  CIVXL U2985 ( .A(n2798), .Z(net22220) );
  CFA1X1 U2986 ( .A(n2195), .B(n1949), .CI(n1920), .CO(n1430), .S(n1431) );
  CEOX1 U2987 ( .A(n3433), .B(n1434), .Z(n1401) );
  CEOX1 U2988 ( .A(n2101), .B(n1411), .Z(n3433) );
  CENX1 U2989 ( .A(n1272), .B(n1266), .Z(n3340) );
  CENX1 U2990 ( .A(n3956), .B(net20996), .Z(n2280) );
  CIVX3 U2991 ( .A(net19213), .Z(net19215) );
  CIVX2 U2992 ( .A(net21206), .Z(net19191) );
  CENX1 U2993 ( .A(n3977), .B(net19302), .Z(n2549) );
  CND2X2 U2994 ( .A(n2827), .B(n6), .Z(n3783) );
  COND2X1 U2995 ( .A(n3876), .B(n2730), .C(n3933), .D(n2729), .Z(n2203) );
  CEOX1 U2996 ( .A(n1435), .B(n1454), .Z(n3743) );
  CND2X1 U2997 ( .A(n1475), .B(n3528), .Z(n3529) );
  CND3XL U2998 ( .A(n3656), .B(n3657), .C(n3658), .Z(n1336) );
  CND2X1 U2999 ( .A(n1369), .B(n1394), .Z(n3400) );
  CEOX1 U3000 ( .A(n3500), .B(n1292), .Z(n1259) );
  CEOX1 U3001 ( .A(n1298), .B(n1300), .Z(n3500) );
  CND2X1 U3002 ( .A(n3352), .B(n3353), .Z(n3359) );
  CENX1 U3003 ( .A(n1112), .B(n1089), .Z(n3240) );
  CND2X1 U3004 ( .A(n3224), .B(net20956), .Z(n241) );
  CND3X1 U3005 ( .A(n3838), .B(n3839), .C(n3840), .Z(n1308) );
  CND2X1 U3006 ( .A(n233), .B(n3223), .Z(n224) );
  CNIVX4 U3007 ( .A(n145), .Z(n3979) );
  CNR2X1 U3008 ( .A(n1713), .B(n1716), .Z(n708) );
  CND2X1 U3009 ( .A(n1015), .B(n1036), .Z(n469) );
  CND2X1 U3010 ( .A(n879), .B(n892), .Z(n379) );
  COND1XL U3011 ( .A(n605), .B(n3102), .C(n606), .Z(n604) );
  CIVX1 U3012 ( .A(n3734), .Z(n3988) );
  CIVX2 U3013 ( .A(n603), .Z(n601) );
  CIVX1 U3014 ( .A(n57), .Z(net18561) );
  CAN2XL U3015 ( .A(n1729), .B(n1925), .Z(n3214) );
  CNIVX1 U3016 ( .A(n1900), .Z(n3215) );
  CAN2X1 U3017 ( .A(n3296), .B(n3297), .Z(n3216) );
  CIVXL U3018 ( .A(net21858), .Z(net21892) );
  CIVX2 U3019 ( .A(n602), .Z(n769) );
  COR2X1 U3020 ( .A(n3499), .B(n1504), .Z(n3217) );
  CAN2XL U3021 ( .A(n1270), .B(n3290), .Z(n3218) );
  CAN2XL U3022 ( .A(n1268), .B(n3291), .Z(n3219) );
  CAN2XL U3023 ( .A(n963), .B(n3309), .Z(n3220) );
  CAN2X1 U3024 ( .A(n1169), .B(n3347), .Z(n3221) );
  COAN1XL U3025 ( .A(n327), .B(n291), .C(n292), .Z(n3222) );
  COR2X1 U3026 ( .A(n796), .B(n795), .Z(n3223) );
  COR2X1 U3027 ( .A(n799), .B(n802), .Z(n3224) );
  COR2X1 U3028 ( .A(n265), .B(n241), .Z(n3225) );
  CNR2X1 U3029 ( .A(n1545), .B(n1562), .Z(n633) );
  CND2XL U3030 ( .A(n1545), .B(n1562), .Z(n634) );
  CENXL U3031 ( .A(n635), .B(n192), .Z(product[20]) );
  CANR1X1 U3032 ( .A(n773), .B(n629), .C(n626), .Z(n624) );
  CENXL U3033 ( .A(n629), .B(n191), .Z(product[21]) );
  CENXL U3034 ( .A(n3226), .B(n619), .Z(product[23]) );
  CAN2XL U3035 ( .A(n3552), .B(n3217), .Z(n3226) );
  CENXL U3036 ( .A(n624), .B(n3227), .Z(product[22]) );
  CAN2XL U3037 ( .A(n772), .B(n623), .Z(n3227) );
  CANR1X1 U3038 ( .A(n608), .B(n769), .C(n601), .Z(n3872) );
  CENX1 U3039 ( .A(n2798), .B(n3985), .Z(n2732) );
  CIVX2 U3040 ( .A(n618), .Z(n616) );
  CND2X2 U3041 ( .A(n1483), .B(n1504), .Z(n618) );
  CND2X2 U3042 ( .A(n2821), .B(n3936), .Z(n3893) );
  CIVXL U3043 ( .A(n671), .Z(n780) );
  CND2X1 U3044 ( .A(n3084), .B(n3471), .Z(n3472) );
  CENXL U3045 ( .A(n185), .B(n584), .Z(product[27]) );
  CENXL U3046 ( .A(n186), .B(n593), .Z(product[26]) );
  CNR2X1 U3047 ( .A(n1525), .B(n1544), .Z(n627) );
  CENXL U3048 ( .A(n187), .B(n604), .Z(product[25]) );
  CENXL U3049 ( .A(n3229), .B(n553), .Z(product[31]) );
  CAN2XL U3050 ( .A(n3881), .B(n552), .Z(n3229) );
  CEOX1 U3051 ( .A(n1729), .B(n1925), .Z(n1543) );
  CANR1XL U3052 ( .A(n766), .B(n3860), .C(n571), .Z(n569) );
  CANR1XL U3053 ( .A(n554), .B(n3860), .C(n555), .Z(n553) );
  CHA1X1 U3054 ( .A(n1730), .B(n1956), .CO(n1578), .S(n1579) );
  CENXL U3055 ( .A(n3969), .B(net19178), .Z(n2562) );
  CENX1 U3056 ( .A(n2782), .B(n3897), .Z(n2683) );
  CENXL U3057 ( .A(n3970), .B(n3897), .Z(n2692) );
  CENX1 U3058 ( .A(n3959), .B(n3923), .Z(n2607) );
  CND2X1 U3059 ( .A(n3798), .B(n3756), .Z(n3231) );
  CND2X1 U3060 ( .A(n3798), .B(n3756), .Z(n81) );
  CND2IX2 U3061 ( .B(n1308), .A(n3610), .Z(n3612) );
  CFA1X1 U3062 ( .A(n2115), .B(n2177), .CI(n1733), .CO(n1658), .S(n1659) );
  CENXL U3063 ( .A(n2792), .B(n3993), .Z(n2627) );
  CENXL U3064 ( .A(n3963), .B(n3993), .Z(n2636) );
  CENXL U3065 ( .A(n2782), .B(n3993), .Z(n2617) );
  CENXL U3066 ( .A(n3973), .B(n3993), .Z(n2623) );
  CENXL U3067 ( .A(n3974), .B(n3993), .Z(n2622) );
  CENXL U3068 ( .A(n2785), .B(n3993), .Z(n2620) );
  CENXL U3069 ( .A(n3975), .B(n3993), .Z(n2621) );
  CENXL U3070 ( .A(n3965), .B(n3993), .Z(n2634) );
  CENX1 U3071 ( .A(n3976), .B(n3993), .Z(n2619) );
  CENX1 U3072 ( .A(n3971), .B(n3993), .Z(n2625) );
  CENX1 U3073 ( .A(n2783), .B(n3993), .Z(n2618) );
  CENX1 U3074 ( .A(n3960), .B(n3993), .Z(n2639) );
  CIVX2 U3075 ( .A(n36), .Z(n3232) );
  CIVX1 U3076 ( .A(n36), .Z(n3233) );
  CIVX2 U3077 ( .A(n36), .Z(n3952) );
  CIVXL U3078 ( .A(n627), .Z(n773) );
  COND1X2 U3079 ( .A(n613), .B(n630), .C(n614), .Z(n3882) );
  CND2X1 U3080 ( .A(n1143), .B(n1141), .Z(n3710) );
  CND2XL U3081 ( .A(n1113), .B(n1136), .Z(n3266) );
  CIVX2 U3082 ( .A(n30), .Z(n3946) );
  CNR2X2 U3083 ( .A(n636), .B(n633), .Z(n631) );
  CIVXL U3084 ( .A(n3498), .Z(n3234) );
  CIVX4 U3085 ( .A(n3371), .Z(net21512) );
  CIVXL U3086 ( .A(n1200), .Z(n3236) );
  CIVXL U3087 ( .A(n3236), .Z(n3237) );
  CIVXL U3088 ( .A(n415), .Z(n413) );
  CENX1 U3089 ( .A(n1084), .B(n1063), .Z(n3425) );
  CNR2X2 U3090 ( .A(n3945), .B(n543), .Z(n534) );
  CNR2X1 U3091 ( .A(n1274), .B(n1245), .Z(n543) );
  CND2XL U3092 ( .A(n414), .B(n748), .Z(n405) );
  CND2X1 U3093 ( .A(n1161), .B(n3441), .Z(n3848) );
  CIVX2 U3094 ( .A(n3940), .Z(n3942) );
  CIVXL U3095 ( .A(n355), .Z(n3238) );
  COAN1X1 U3096 ( .A(n458), .B(n448), .C(n449), .Z(n3239) );
  CND2IX2 U3097 ( .B(n3832), .A(n3833), .Z(n3834) );
  COND1X2 U3098 ( .A(n530), .B(n3741), .C(n3797), .Z(n3326) );
  CND2X1 U3099 ( .A(n1162), .B(n1164), .Z(n3644) );
  CENX1 U3100 ( .A(n3240), .B(n1110), .Z(n1085) );
  CENX1 U3101 ( .A(n3241), .B(n3388), .Z(n1257) );
  CENX1 U3102 ( .A(n1265), .B(n1269), .Z(n3241) );
  CND2XL U3103 ( .A(n1244), .B(n1215), .Z(n3242) );
  CENX2 U3104 ( .A(n3968), .B(n3992), .Z(n2662) );
  CENXL U3105 ( .A(n2792), .B(net18547), .Z(n2528) );
  CNIVXL U3106 ( .A(n2444), .Z(n3243) );
  CND2X1 U3107 ( .A(n1109), .B(n1134), .Z(n3949) );
  CENXL U3108 ( .A(n3963), .B(n4005), .Z(n2339) );
  CENXL U3109 ( .A(n3959), .B(n3984), .Z(n2739) );
  CENXL U3110 ( .A(n3958), .B(n3984), .Z(n2740) );
  CENXL U3111 ( .A(n2810), .B(n3985), .Z(n2744) );
  CENXL U3112 ( .A(n2809), .B(n3985), .Z(n2743) );
  CENXL U3113 ( .A(n3962), .B(n3984), .Z(n2736) );
  CENXL U3114 ( .A(n3956), .B(n3984), .Z(n2742) );
  CENXL U3115 ( .A(n3961), .B(n3984), .Z(n2737) );
  CENXL U3116 ( .A(n3957), .B(n3985), .Z(n2741) );
  CENXL U3117 ( .A(n3977), .B(n3985), .Z(n2714) );
  CENXL U3118 ( .A(n3965), .B(n3985), .Z(n2733) );
  CIVX1 U3119 ( .A(n353), .Z(n355) );
  CND2XL U3120 ( .A(n3237), .B(n1175), .Z(n3707) );
  CIVXL U3121 ( .A(n666), .Z(n664) );
  CND2X1 U3122 ( .A(n779), .B(n666), .Z(n197) );
  COND1X1 U3123 ( .A(n666), .B(n660), .C(n661), .Z(n659) );
  CIVXL U3124 ( .A(net22590), .Z(n3244) );
  COAN1X1 U3125 ( .A(n434), .B(n424), .C(n425), .Z(n417) );
  CND2X1 U3126 ( .A(n3449), .B(n974), .Z(n434) );
  CND2X1 U3127 ( .A(n1254), .B(n1229), .Z(n3525) );
  CIVX3 U3128 ( .A(net19171), .Z(net18517) );
  CENX1 U3129 ( .A(n3959), .B(n3991), .Z(n2673) );
  CHA1XL U3130 ( .A(n1731), .B(n1988), .CO(n1610), .S(n1611) );
  CND2XL U3131 ( .A(n2782), .B(n3990), .Z(n3247) );
  CND2X1 U3132 ( .A(n3245), .B(n3246), .Z(n3248) );
  CND2X1 U3133 ( .A(n3247), .B(n3248), .Z(n2650) );
  CIVXL U3134 ( .A(n2782), .Z(n3245) );
  CIVXL U3135 ( .A(n3990), .Z(n3246) );
  CEOX1 U3136 ( .A(n3429), .B(n1547), .Z(n1545) );
  CNR2X1 U3137 ( .A(n1333), .B(n1360), .Z(n3249) );
  CENX2 U3138 ( .A(n3337), .B(n1335), .Z(n1333) );
  CND2X1 U3139 ( .A(n878), .B(n867), .Z(n370) );
  CND2X2 U3140 ( .A(n51), .B(n2822), .Z(n3250) );
  COAN1X1 U3141 ( .A(n592), .B(n3886), .C(n583), .Z(n579) );
  CIVXL U3142 ( .A(n592), .Z(n590) );
  CIVX3 U3143 ( .A(net18547), .Z(net22399) );
  CEOX2 U3144 ( .A(n1088), .B(n1065), .Z(n3252) );
  CEOX2 U3145 ( .A(n3252), .B(n1086), .Z(n1061) );
  CND2XL U3146 ( .A(n1086), .B(n1065), .Z(n3253) );
  CND2XL U3147 ( .A(n1065), .B(n1088), .Z(n3255) );
  CND3X1 U3148 ( .A(n3253), .B(n3254), .C(n3255), .Z(n1060) );
  CND2X1 U3149 ( .A(n3661), .B(n3257), .Z(n3258) );
  CND2X1 U3150 ( .A(n3256), .B(n1039), .Z(n3259) );
  CND2X2 U3151 ( .A(n3258), .B(n3259), .Z(n1037) );
  CIVX2 U3152 ( .A(n3661), .Z(n3256) );
  CIVXL U3153 ( .A(n1039), .Z(n3257) );
  CIVXL U3154 ( .A(n379), .Z(n377) );
  CENXL U3155 ( .A(n3969), .B(n3985), .Z(n2727) );
  CENXL U3156 ( .A(n3968), .B(n3985), .Z(n2728) );
  CENXL U3157 ( .A(net18979), .B(n3985), .Z(n2731) );
  COND2XL U3158 ( .A(n3550), .B(n2555), .C(n3660), .D(n2554), .Z(n2028) );
  CIVXL U3159 ( .A(n1530), .Z(n3260) );
  CIVX1 U3160 ( .A(n3260), .Z(n3261) );
  CENX1 U3161 ( .A(n3956), .B(n3923), .Z(n2610) );
  CENX1 U3162 ( .A(n2781), .B(n3923), .Z(n2583) );
  CENX2 U3163 ( .A(n1414), .B(n1391), .Z(n3590) );
  CIVXL U3164 ( .A(n3380), .Z(n3262) );
  COND2XL U3165 ( .A(net21433), .B(n2289), .C(net19192), .D(n2288), .Z(n1774)
         );
  COND2XL U3166 ( .A(net21433), .B(n2291), .C(net19192), .D(n2290), .Z(n1776)
         );
  CNR2X1 U3167 ( .A(n361), .B(n416), .Z(n3263) );
  CNR2X2 U3168 ( .A(n361), .B(n416), .Z(n359) );
  CIVX4 U3169 ( .A(n3734), .Z(n3897) );
  CIVX4 U3170 ( .A(n75), .Z(n3659) );
  CEOX2 U3171 ( .A(n1138), .B(n1136), .Z(n3265) );
  CEOX2 U3172 ( .A(n3265), .B(n3111), .Z(n1109) );
  CND2X1 U3173 ( .A(n1113), .B(n1138), .Z(n3267) );
  CND2X1 U3174 ( .A(n1138), .B(n1136), .Z(n3268) );
  CND3X1 U3175 ( .A(n3266), .B(n3267), .C(n3268), .Z(n1108) );
  CND2X1 U3176 ( .A(n3603), .B(n1419), .Z(n3271) );
  CND2X2 U3177 ( .A(n3269), .B(n3270), .Z(n3272) );
  CND2X2 U3178 ( .A(n3271), .B(n3272), .Z(n1415) );
  CIVX2 U3179 ( .A(n3603), .Z(n3269) );
  CIVXL U3180 ( .A(n1419), .Z(n3270) );
  CND2X1 U3181 ( .A(n3983), .B(a[2]), .Z(n3275) );
  CND2X2 U3182 ( .A(n3273), .B(n3274), .Z(n3276) );
  CND2X4 U3183 ( .A(n3275), .B(n3276), .Z(n3922) );
  CIVX2 U3184 ( .A(n3983), .Z(n3273) );
  CIVX2 U3185 ( .A(a[2]), .Z(n3274) );
  CIVX3 U3186 ( .A(n3922), .Z(n3933) );
  CIVX4 U3187 ( .A(n3922), .Z(n3934) );
  CEOX2 U3188 ( .A(n3277), .B(n1231), .Z(n1223) );
  CND2XL U3189 ( .A(n1231), .B(n3029), .Z(n3278) );
  CND2X1 U3190 ( .A(n1231), .B(n1258), .Z(n3279) );
  CND2XL U3191 ( .A(n3029), .B(n1258), .Z(n3280) );
  CND3X1 U3192 ( .A(n3278), .B(n3279), .C(n3280), .Z(n1222) );
  CENX1 U3193 ( .A(n3340), .B(n1264), .Z(n1231) );
  CND2X1 U3194 ( .A(n1223), .B(n1252), .Z(n3796) );
  CENX1 U3195 ( .A(n1174), .B(n1172), .Z(n3322) );
  CENX2 U3196 ( .A(n1416), .B(n3692), .Z(n1389) );
  CENX1 U3197 ( .A(n1064), .B(n1043), .Z(n3324) );
  CIVX2 U3198 ( .A(n1163), .Z(n3832) );
  CIVXL U3199 ( .A(n1227), .Z(n3281) );
  COND2X1 U3200 ( .A(n72), .B(net21948), .C(net19215), .D(n2548), .Z(n1732) );
  CEO3X2 U3201 ( .A(n1203), .B(n1228), .C(n1226), .Z(n1195) );
  CND2X1 U3202 ( .A(n1203), .B(n1226), .Z(n3282) );
  CND2X1 U3203 ( .A(n1226), .B(n1228), .Z(n3284) );
  CND3X2 U3204 ( .A(n3282), .B(n3283), .C(n3284), .Z(n1194) );
  CENX2 U3205 ( .A(a[22]), .B(n4003), .Z(n3285) );
  CENX2 U3206 ( .A(a[22]), .B(n4003), .Z(net21375) );
  CND3X1 U3207 ( .A(n3517), .B(n3518), .C(n3519), .Z(n1504) );
  CENX1 U3208 ( .A(n3966), .B(net21909), .Z(n2301) );
  CENX1 U3209 ( .A(n3969), .B(net21909), .Z(n2298) );
  CFA1XL U3210 ( .A(n890), .B(n1897), .CI(n1809), .CO(n876), .S(n877) );
  COND2X2 U3211 ( .A(n126), .B(n2346), .C(net22007), .D(n3782), .Z(n1829) );
  CNIVX2 U3212 ( .A(n2345), .Z(n3782) );
  CNR2XL U3213 ( .A(n3068), .B(n594), .Z(n3286) );
  CENXL U3214 ( .A(n2792), .B(net21909), .Z(n3287) );
  CEOX1 U3215 ( .A(n3967), .B(net21622), .Z(n2564) );
  CENXL U3216 ( .A(n3958), .B(n3770), .Z(n2443) );
  CENXL U3217 ( .A(n3977), .B(n3770), .Z(n2417) );
  CENXL U3218 ( .A(n3963), .B(n3770), .Z(n2438) );
  CENX2 U3219 ( .A(n1164), .B(n1139), .Z(n3288) );
  CENX2 U3220 ( .A(net22241), .B(n3682), .Z(n3878) );
  CIVX1 U3221 ( .A(a[12]), .Z(n3682) );
  CIVX1 U3222 ( .A(n1268), .Z(n3290) );
  CIVX1 U3223 ( .A(n1270), .Z(n3291) );
  CIVXL U3224 ( .A(n1235), .Z(n3292) );
  CND2X1 U3225 ( .A(n3291), .B(n3294), .Z(n3293) );
  CND2X1 U3226 ( .A(n3292), .B(n3218), .Z(n3295) );
  CND2X1 U3227 ( .A(n3292), .B(n3219), .Z(n3296) );
  CND2X1 U3228 ( .A(n1268), .B(n3298), .Z(n3297) );
  CND2X1 U3229 ( .A(n1270), .B(n1268), .Z(n3299) );
  CND2X1 U3230 ( .A(n1235), .B(n1268), .Z(n3300) );
  CND2XL U3231 ( .A(n1235), .B(n3290), .Z(n3301) );
  CIVX1 U3232 ( .A(n3301), .Z(n3294) );
  CND2X1 U3233 ( .A(n1235), .B(n1270), .Z(n3302) );
  CIVX2 U3234 ( .A(n3302), .Z(n3298) );
  CND2X1 U3235 ( .A(n3293), .B(n3295), .Z(n3303) );
  CND2X1 U3236 ( .A(n3299), .B(n3300), .Z(n3304) );
  CIVX2 U3237 ( .A(n3304), .Z(n3289) );
  CND2IX2 U3238 ( .B(n3298), .A(n3289), .Z(n1228) );
  CND2IX2 U3239 ( .B(n3303), .A(n3216), .Z(n1229) );
  CND3X1 U3240 ( .A(n3510), .B(n3511), .C(n3512), .Z(n1268) );
  CENX2 U3241 ( .A(n3970), .B(n3925), .Z(n2428) );
  CND2X1 U3242 ( .A(n1315), .B(n1338), .Z(n3838) );
  CND2XL U3243 ( .A(n1789), .B(n2025), .Z(n3428) );
  CND2XL U3244 ( .A(n1846), .B(n1789), .Z(n3426) );
  CENX2 U3245 ( .A(n3971), .B(n3925), .Z(n2427) );
  CND2X2 U3246 ( .A(n3305), .B(n3306), .Z(n959) );
  CIVX1 U3247 ( .A(n980), .Z(n3309) );
  CND2X1 U3248 ( .A(n3310), .B(n3319), .Z(n3312) );
  CND2X1 U3249 ( .A(n3310), .B(n3220), .Z(n3313) );
  CND2XL U3250 ( .A(n980), .B(n963), .Z(n3315) );
  CND2XL U3251 ( .A(n978), .B(n963), .Z(n3316) );
  CND2XL U3252 ( .A(n978), .B(n980), .Z(n3307) );
  CND2X1 U3253 ( .A(n3311), .B(n3312), .Z(n3317) );
  CIVX2 U3254 ( .A(n3317), .Z(n3305) );
  CND2X1 U3255 ( .A(n3313), .B(n3314), .Z(n3318) );
  CIVX2 U3256 ( .A(n3318), .Z(n3306) );
  CNR2XL U3257 ( .A(n3309), .B(n963), .Z(n3319) );
  CND2XL U3258 ( .A(n978), .B(n3320), .Z(n3314) );
  CNR2IXL U3259 ( .B(n980), .A(n3308), .Z(n3320) );
  CND2X1 U3260 ( .A(n978), .B(n3321), .Z(n3311) );
  CNR2XL U3261 ( .A(n963), .B(n980), .Z(n3321) );
  COND2X1 U3262 ( .A(net21802), .B(n2456), .C(net21846), .D(n2455), .Z(n1933)
         );
  CENX1 U3263 ( .A(n3723), .B(net21622), .Z(n2563) );
  CIVX1 U3264 ( .A(n3968), .Z(n3723) );
  CENX1 U3265 ( .A(n1170), .B(n3322), .Z(n1141) );
  CND3X1 U3266 ( .A(n3656), .B(n3657), .C(n3658), .Z(n3323) );
  CND2XL U3267 ( .A(n1336), .B(n1313), .Z(n3586) );
  CENX1 U3268 ( .A(n3324), .B(n1062), .Z(n1039) );
  CND2X2 U3269 ( .A(n1037), .B(n1058), .Z(n472) );
  CNR2X1 U3270 ( .A(n1037), .B(n1058), .Z(n471) );
  CND3X1 U3271 ( .A(n3693), .B(n3694), .C(n3695), .Z(n1058) );
  CEOXL U3272 ( .A(n3957), .B(n3380), .Z(n2312) );
  CND2X2 U3273 ( .A(n3581), .B(n3582), .Z(n3325) );
  CND2X1 U3274 ( .A(n3581), .B(n3582), .Z(n1059) );
  COND2X1 U3275 ( .A(n3755), .B(n2757), .C(n6), .D(n2756), .Z(n2230) );
  CIVXL U3276 ( .A(n528), .Z(n3327) );
  CND2X2 U3277 ( .A(n2817), .B(n96), .Z(n3328) );
  CND2X1 U3278 ( .A(n2817), .B(n96), .Z(n99) );
  CND2X2 U3279 ( .A(n2817), .B(n96), .Z(net21344) );
  COND2XL U3280 ( .A(n99), .B(n2428), .C(net21744), .D(n2427), .Z(n3329) );
  CND2XL U3281 ( .A(n1170), .B(n1174), .Z(n3819) );
  COND2X1 U3282 ( .A(n144), .B(net18489), .C(net22439), .D(n2284), .Z(n1724)
         );
  CENX2 U3283 ( .A(n2798), .B(n3926), .Z(n2435) );
  CIVX1 U3284 ( .A(n3895), .Z(n3863) );
  CND2X2 U3285 ( .A(n3895), .B(net21693), .Z(n3804) );
  COND2XL U3286 ( .A(n81), .B(n2499), .C(n3651), .D(n2498), .Z(n3330) );
  CENX2 U3287 ( .A(a[30]), .B(n3379), .Z(n3331) );
  CENX2 U3288 ( .A(a[30]), .B(n3379), .Z(n141) );
  CENX2 U3289 ( .A(n2798), .B(n3923), .Z(n2600) );
  CIVXL U3290 ( .A(n3264), .Z(n667) );
  CND3X2 U3291 ( .A(n3413), .B(n3414), .C(n3415), .Z(n1018) );
  CND2X1 U3292 ( .A(n1023), .B(n1025), .Z(n3415) );
  COND1X1 U3293 ( .A(n410), .B(n402), .C(n403), .Z(n397) );
  CENX2 U3294 ( .A(n3334), .B(n3751), .Z(n1283) );
  COR2X2 U3295 ( .A(n3651), .B(n2500), .Z(n3459) );
  CND2X1 U3296 ( .A(net20990), .B(n749), .Z(n3335) );
  CND3X2 U3297 ( .A(n3620), .B(n3621), .C(n3622), .Z(n1460) );
  CND2XL U3298 ( .A(n1484), .B(n1465), .Z(n3622) );
  COND2X1 U3299 ( .A(n3887), .B(n2461), .C(net21846), .D(n2460), .Z(n1080) );
  CENX2 U3300 ( .A(n3971), .B(net19314), .Z(n2460) );
  CND2IX1 U3301 ( .B(n3864), .A(a[26]), .Z(n3805) );
  COND2X1 U3302 ( .A(n144), .B(n2262), .C(n3173), .D(n2261), .Z(n1748) );
  COND2XL U3303 ( .A(n144), .B(n2259), .C(n3173), .D(n2258), .Z(n1745) );
  COND2XL U3304 ( .A(n144), .B(n2261), .C(n3173), .D(n2260), .Z(n1747) );
  CENX1 U3305 ( .A(a[28]), .B(n4007), .Z(n3336) );
  CENX1 U3306 ( .A(a[28]), .B(n4007), .Z(net21206) );
  COND2X2 U3307 ( .A(n2583), .B(n54), .C(n3145), .D(n2582), .Z(n2056) );
  CND3X2 U3308 ( .A(n3949), .B(n3950), .C(n3951), .Z(n1106) );
  CND2X1 U3309 ( .A(n1139), .B(n1164), .Z(n3645) );
  CENX2 U3310 ( .A(n1019), .B(n1038), .Z(n3338) );
  CENX2 U3311 ( .A(n3956), .B(net19268), .Z(n2379) );
  COND1X1 U3312 ( .A(n361), .B(n417), .C(n3124), .Z(n3339) );
  COND1X1 U3313 ( .A(n361), .B(n417), .C(n362), .Z(n360) );
  CNR2X1 U3314 ( .A(n907), .B(n922), .Z(n3341) );
  CNR2X1 U3315 ( .A(n907), .B(n922), .Z(n402) );
  CND3X1 U3316 ( .A(net22302), .B(net22303), .C(net22304), .Z(n922) );
  CIVX1 U3317 ( .A(n920), .Z(n921) );
  CENXL U3318 ( .A(n2782), .B(net19178), .Z(n3342) );
  CIVX3 U3319 ( .A(net21438), .Z(net19178) );
  CIVX2 U3320 ( .A(net18561), .Z(net18555) );
  CND2X1 U3321 ( .A(n1221), .B(n1250), .Z(n3737) );
  CENX2 U3322 ( .A(n3957), .B(net19268), .Z(n2378) );
  CND2X1 U3323 ( .A(n2237), .B(n2144), .Z(n3463) );
  CENX2 U3324 ( .A(n3973), .B(net19314), .Z(n2458) );
  CND2IX1 U3325 ( .B(n1041), .A(n1060), .Z(n3486) );
  CNR2X2 U3326 ( .A(n511), .B(n3637), .Z(n3343) );
  CNR2X1 U3327 ( .A(n511), .B(n3637), .Z(n498) );
  CND2X1 U3328 ( .A(n498), .B(n3062), .Z(n480) );
  CENX1 U3329 ( .A(n3976), .B(net19314), .Z(n2454) );
  CIVXL U3330 ( .A(n954), .Z(n955) );
  COND1X1 U3331 ( .A(n547), .B(n575), .C(n548), .Z(net22599) );
  CNR2X2 U3332 ( .A(n1685), .B(n1692), .Z(n693) );
  CND2X1 U3333 ( .A(n1685), .B(n1692), .Z(n694) );
  CND2XL U3334 ( .A(n1292), .B(n1300), .Z(n3501) );
  CHA1X1 U3335 ( .A(n2051), .B(n2020), .CO(n1638), .S(n1639) );
  COND2X1 U3336 ( .A(n2547), .B(net21352), .C(net19215), .D(n2546), .Z(n2020)
         );
  CENX2 U3337 ( .A(n3974), .B(n3923), .Z(n2589) );
  COND2X1 U3338 ( .A(n3953), .B(n2661), .C(n3803), .D(n2660), .Z(n2134) );
  COND2X1 U3339 ( .A(n3953), .B(n2666), .C(n3803), .D(n2665), .Z(n2139) );
  CEOXL U3340 ( .A(n3960), .B(n3167), .Z(n2441) );
  CENX2 U3341 ( .A(n3963), .B(net19314), .Z(n2471) );
  COND2XL U3342 ( .A(n3328), .B(n2429), .C(net21744), .D(n2428), .Z(n1906) );
  CENX2 U3343 ( .A(n3966), .B(net19302), .Z(n3650) );
  CENX2 U3344 ( .A(n3958), .B(net19302), .Z(n2575) );
  CND2X2 U3345 ( .A(n3346), .B(n3345), .Z(n1163) );
  CIVX2 U3346 ( .A(n1194), .Z(n3347) );
  CIVX2 U3347 ( .A(n1169), .Z(n3348) );
  CIVX1 U3348 ( .A(n1167), .Z(n3349) );
  CND2X1 U3349 ( .A(n3348), .B(n3116), .Z(n3350) );
  CND2X1 U3350 ( .A(n3349), .B(n3221), .Z(n3351) );
  CND2XL U3351 ( .A(n1169), .B(n1194), .Z(n3355) );
  CND2X1 U3352 ( .A(n1167), .B(n1169), .Z(n3357) );
  CIVX2 U3353 ( .A(n3357), .Z(n3354) );
  CIVX2 U3354 ( .A(n3358), .Z(n3345) );
  CIVX2 U3355 ( .A(n3359), .Z(n3346) );
  CND2IX2 U3356 ( .B(n3354), .A(n3360), .Z(n1162) );
  CAN2X1 U3357 ( .A(n3355), .B(n3356), .Z(n3360) );
  CND2IX1 U3358 ( .B(n3347), .A(n3354), .Z(n3353) );
  CEO3X2 U3359 ( .A(n1200), .B(n1175), .C(n1198), .Z(n1167) );
  CENX1 U3360 ( .A(n2792), .B(n3926), .Z(n2429) );
  CND2X2 U3361 ( .A(n3362), .B(n3363), .Z(n1978) );
  CIVX1 U3362 ( .A(n2503), .Z(n3364) );
  CIVX1 U3363 ( .A(n3942), .Z(n3365) );
  CIVX1 U3364 ( .A(n2504), .Z(n3366) );
  CND2X1 U3365 ( .A(n3364), .B(n3365), .Z(n3362) );
  CND2X2 U3366 ( .A(n3366), .B(n3367), .Z(n3363) );
  CENX1 U3367 ( .A(n2782), .B(n3923), .Z(n2584) );
  CND2XL U3368 ( .A(n757), .B(n505), .Z(n175) );
  CND2X1 U3369 ( .A(n1217), .B(n1246), .Z(n3666) );
  CEOX1 U3370 ( .A(n3960), .B(net21892), .Z(n2375) );
  CNR2X2 U3371 ( .A(n3325), .B(n1082), .Z(n484) );
  CENX1 U3372 ( .A(n3967), .B(net20996), .Z(n2267) );
  COND2X2 U3373 ( .A(n3887), .B(n2471), .C(n87), .D(n2470), .Z(n1946) );
  CIVX4 U3374 ( .A(net21835), .Z(net21836) );
  COND2X1 U3375 ( .A(n2481), .B(net21801), .C(n87), .D(n2480), .Z(n1956) );
  CENX2 U3376 ( .A(n1595), .B(n3368), .Z(n1587) );
  CND2XL U3377 ( .A(n1283), .B(n1308), .Z(n3842) );
  COND2X1 U3378 ( .A(n3228), .B(n2578), .C(n3618), .D(n2577), .Z(n2051) );
  CND2IX1 U3379 ( .B(n3989), .A(n3478), .Z(n3480) );
  CENX2 U3380 ( .A(n3369), .B(n1217), .Z(n1215) );
  CENX2 U3381 ( .A(n1219), .B(n1246), .Z(n3369) );
  CIVX3 U3382 ( .A(n3232), .Z(n3904) );
  CIVX3 U3383 ( .A(n3952), .Z(n3954) );
  CIVX2 U3384 ( .A(n3233), .Z(n3953) );
  CND2X4 U3385 ( .A(net21846), .B(n2818), .Z(n90) );
  CANR1X1 U3386 ( .A(n3263), .B(net22552), .C(n360), .Z(n3370) );
  CANR1X1 U3387 ( .A(n3263), .B(net22552), .C(n3339), .Z(n354) );
  CIVX1 U3388 ( .A(n3370), .Z(n356) );
  CANR1X1 U3389 ( .A(n739), .B(n308), .C(n301), .Z(n299) );
  COND1XL U3390 ( .A(n298), .B(net19189), .C(n299), .Z(n297) );
  CIVX2 U3391 ( .A(n303), .Z(n301) );
  CIVX2 U3392 ( .A(n302), .Z(n739) );
  CND2XL U3393 ( .A(n307), .B(n739), .Z(n298) );
  CND2XL U3394 ( .A(n739), .B(n303), .Z(n157) );
  COND1X1 U3395 ( .A(n309), .B(n354), .C(n310), .Z(n308) );
  CIVXL U3396 ( .A(n308), .Z(n306) );
  CANR1XL U3397 ( .A(n740), .B(n323), .C(n314), .Z(n310) );
  CIVX2 U3398 ( .A(n316), .Z(n314) );
  CANR1XL U3399 ( .A(n314), .B(n293), .C(n294), .Z(n292) );
  CIVX2 U3400 ( .A(n315), .Z(n740) );
  CND2XL U3401 ( .A(n320), .B(n740), .Z(n309) );
  CND2XL U3402 ( .A(n740), .B(n316), .Z(n158) );
  CND2X1 U3403 ( .A(n293), .B(n740), .Z(n291) );
  CNR2X1 U3404 ( .A(n827), .B(n834), .Z(n315) );
  CND2X1 U3405 ( .A(n826), .B(n819), .Z(n303) );
  COND1XL U3406 ( .A(n295), .B(n303), .C(n296), .Z(n294) );
  CNR2X1 U3407 ( .A(n826), .B(n819), .Z(n302) );
  CNR2X1 U3408 ( .A(n302), .B(n295), .Z(n293) );
  CNR2X1 U3409 ( .A(n353), .B(n309), .Z(n307) );
  COND1X1 U3410 ( .A(n261), .B(n354), .C(n262), .Z(n260) );
  COND1XL U3411 ( .A(n224), .B(n3370), .C(n225), .Z(n223) );
  CANR1XL U3412 ( .A(n320), .B(n356), .C(n323), .Z(n319) );
  CND2X1 U3413 ( .A(n827), .B(n834), .Z(n316) );
  COND1X1 U3414 ( .A(n392), .B(n3251), .C(n366), .Z(n364) );
  COAN1X1 U3415 ( .A(n369), .B(n379), .C(n370), .Z(n366) );
  COND1X1 U3416 ( .A(net22511), .B(n461), .C(n445), .Z(net22552) );
  COND1XL U3417 ( .A(n324), .B(n334), .C(n327), .Z(n323) );
  CENXL U3418 ( .A(n297), .B(n156), .Z(product[56]) );
  CND2X1 U3419 ( .A(n738), .B(n296), .Z(n156) );
  CIVX2 U3420 ( .A(n295), .Z(n738) );
  CND2X1 U3421 ( .A(n813), .B(n818), .Z(n296) );
  CNR2X1 U3422 ( .A(n813), .B(n818), .Z(n295) );
  CIVXL U3423 ( .A(n307), .Z(n305) );
  CANR1X1 U3424 ( .A(n478), .B(n3817), .C(n479), .Z(net21297) );
  CANR1X1 U3425 ( .A(net21983), .B(net22598), .C(net21313), .Z(net21389) );
  CIVX4 U3426 ( .A(n3373), .Z(net21744) );
  CIVX2 U3427 ( .A(n84), .Z(net22626) );
  CIVX8 U3428 ( .A(net19062), .Z(net21846) );
  CIVX4 U3429 ( .A(n114), .Z(n3371) );
  CIVX8 U3430 ( .A(n3371), .Z(net19281) );
  CND2X2 U3431 ( .A(net22288), .B(n3372), .Z(n114) );
  CND2X1 U3432 ( .A(net22286), .B(net19171), .Z(n3372) );
  CIVX2 U3433 ( .A(net19171), .Z(net22287) );
  CIVX2 U3434 ( .A(a[24]), .Z(net22286) );
  CND2X2 U3435 ( .A(a[24]), .B(net22287), .Z(net22288) );
  CIVX2 U3436 ( .A(n3336), .Z(net19193) );
  CND2XL U3437 ( .A(n940), .B(n927), .Z(net22304) );
  CND2X1 U3438 ( .A(n925), .B(n927), .Z(net22303) );
  COND2X1 U3439 ( .A(net21311), .B(n2363), .C(net21512), .D(n2362), .Z(n1843)
         );
  CNIVX4 U3440 ( .A(net21375), .Z(net21250) );
  CIVX8 U3441 ( .A(net22004), .Z(net22007) );
  CIVX8 U3442 ( .A(net21472), .Z(net22004) );
  CND2X1 U3443 ( .A(n907), .B(n922), .Z(n403) );
  CND2XL U3444 ( .A(n925), .B(n940), .Z(net22302) );
  CEOX2 U3445 ( .A(net22301), .B(n925), .Z(n923) );
  CENX4 U3446 ( .A(a[26]), .B(net19081), .Z(net21472) );
  COND2X1 U3447 ( .A(n2517), .B(net19216), .C(n2518), .D(net21353), .Z(n1992)
         );
  CIVX4 U3448 ( .A(n3377), .Z(net19216) );
  CIVX1 U3449 ( .A(n69), .Z(n3377) );
  COND2X1 U3450 ( .A(n108), .B(n2395), .C(net21250), .D(n2394), .Z(n992) );
  CENXL U3451 ( .A(n2781), .B(net18547), .Z(n2517) );
  CIVX3 U3452 ( .A(n3374), .Z(net18547) );
  CIVX2 U3453 ( .A(n66), .Z(n3374) );
  CIVX3 U3454 ( .A(n3374), .Z(net18549) );
  CENXL U3455 ( .A(n2782), .B(net18547), .Z(n2518) );
  CND2X4 U3456 ( .A(net21896), .B(n3375), .Z(net21353) );
  CIVX2 U3457 ( .A(n3376), .Z(n3375) );
  CIVX1 U3458 ( .A(n69), .Z(net19213) );
  CIVX2 U3459 ( .A(n57), .Z(net21438) );
  CANR1X1 U3460 ( .A(n3224), .B(n260), .C(n253), .Z(n249) );
  COND1XL U3461 ( .A(n248), .B(net19189), .C(n249), .Z(n247) );
  CIVX2 U3462 ( .A(n255), .Z(n253) );
  CND2XL U3463 ( .A(n259), .B(n3224), .Z(n248) );
  CND2XL U3464 ( .A(n3224), .B(n255), .Z(n153) );
  CIVXL U3465 ( .A(n260), .Z(n258) );
  CANR1X1 U3466 ( .A(n736), .B(n273), .C(n264), .Z(n262) );
  CIVX2 U3467 ( .A(n266), .Z(n264) );
  CIVX1 U3468 ( .A(n275), .Z(n273) );
  CANR1XL U3469 ( .A(n272), .B(n356), .C(n273), .Z(n269) );
  CIVX2 U3470 ( .A(n265), .Z(n736) );
  CND2X1 U3471 ( .A(n272), .B(n736), .Z(n261) );
  CND2XL U3472 ( .A(n736), .B(n266), .Z(n154) );
  CND2X1 U3473 ( .A(n799), .B(n802), .Z(n255) );
  COR2X1 U3474 ( .A(n798), .B(n797), .Z(net20956) );
  CND2X1 U3475 ( .A(n798), .B(n797), .Z(n246) );
  COND2XL U3476 ( .A(n144), .B(n2256), .C(n3331), .D(n2255), .Z(n1742) );
  CND2X2 U3477 ( .A(n363), .B(n396), .Z(n361) );
  CIVXL U3478 ( .A(n397), .Z(n399) );
  CANR1XL U3479 ( .A(n3096), .B(n415), .C(n3199), .Z(n395) );
  CND2IXL U3480 ( .B(n389), .A(n392), .Z(n164) );
  COND1XL U3481 ( .A(n389), .B(n399), .C(n392), .Z(n388) );
  CND2XL U3482 ( .A(n744), .B(n370), .Z(n162) );
  CIVX2 U3483 ( .A(n378), .Z(n745) );
  CND2XL U3484 ( .A(n745), .B(n383), .Z(n372) );
  CND2XL U3485 ( .A(n745), .B(n379), .Z(n163) );
  COND1XL U3486 ( .A(n434), .B(n424), .C(n425), .Z(net22590) );
  CND2XL U3487 ( .A(net20990), .B(n434), .Z(n168) );
  CNR2X1 U3488 ( .A(n353), .B(n261), .Z(n259) );
  CIVX2 U3489 ( .A(n274), .Z(n272) );
  CND2XL U3490 ( .A(n355), .B(n272), .Z(n268) );
  CND2X1 U3491 ( .A(n806), .B(n803), .Z(n266) );
  COAN1X1 U3492 ( .A(n266), .B(n241), .C(n242), .Z(n3378) );
  CANR1X2 U3493 ( .A(net20981), .B(n286), .C(n277), .Z(n275) );
  CIVX2 U3494 ( .A(n279), .Z(n277) );
  CNR2X1 U3495 ( .A(n806), .B(n803), .Z(n265) );
  CIVXL U3496 ( .A(n3341), .Z(n747) );
  CNR2X2 U3497 ( .A(n409), .B(n3341), .Z(n396) );
  CENXL U3498 ( .A(n247), .B(n152), .Z(product[60]) );
  CND2XL U3499 ( .A(net20956), .B(n246), .Z(n152) );
  CIVX2 U3500 ( .A(n246), .Z(n244) );
  CNR2IX1 U3501 ( .B(n396), .A(n389), .Z(n387) );
  CND2XL U3502 ( .A(n748), .B(n410), .Z(n166) );
  CIVX2 U3503 ( .A(n410), .Z(n408) );
  CND2XL U3504 ( .A(n747), .B(n403), .Z(n165) );
  CNR2X2 U3505 ( .A(n923), .B(n938), .Z(n409) );
  CIVDX2 U3506 ( .A(n129), .Z0(n3380), .Z1(n3379) );
  CIVX2 U3507 ( .A(n3380), .Z(net18495) );
  COND2X1 U3508 ( .A(net21433), .B(n3380), .C(net19193), .D(n2317), .Z(n1725)
         );
  CENX2 U3509 ( .A(net18489), .B(a[30]), .Z(n2812) );
  CENXL U3510 ( .A(n2798), .B(net20996), .Z(n2270) );
  CNIVX3 U3511 ( .A(n136), .Z(net20996) );
  CENXL U3512 ( .A(net18979), .B(net20996), .Z(n2269) );
  CNIVX4 U3513 ( .A(n2797), .Z(net18979) );
  CIVX4 U3514 ( .A(n136), .Z(net18489) );
  CEO3X2 U3515 ( .A(n1042), .B(n1040), .C(n1021), .Z(n1017) );
  CND2X1 U3516 ( .A(n1042), .B(n1040), .Z(n3381) );
  CND2X1 U3517 ( .A(n1042), .B(n1021), .Z(n3382) );
  CND2X1 U3518 ( .A(n1040), .B(n1021), .Z(n3383) );
  CND3X2 U3519 ( .A(n3381), .B(n3382), .C(n3383), .Z(n1016) );
  CND2X1 U3520 ( .A(n999), .B(n1016), .Z(n3385) );
  CND2XL U3521 ( .A(n997), .B(n1016), .Z(n3386) );
  CND3X1 U3522 ( .A(n3384), .B(n3385), .C(n3386), .Z(n994) );
  CND2X1 U3523 ( .A(n1288), .B(n1286), .Z(n3790) );
  CNIVXL U3524 ( .A(n1271), .Z(n3388) );
  CEO3X1 U3525 ( .A(n1973), .B(n2189), .C(n1768), .Z(n1271) );
  CEOX2 U3526 ( .A(n1491), .B(n1508), .Z(n3389) );
  CEOX2 U3527 ( .A(n3389), .B(n1489), .Z(n1485) );
  CND2XL U3528 ( .A(n1508), .B(n1489), .Z(n3390) );
  CND2X1 U3529 ( .A(n1489), .B(n1491), .Z(n3391) );
  CND2XL U3530 ( .A(n1508), .B(n1491), .Z(n3392) );
  CND3X2 U3531 ( .A(n3390), .B(n3391), .C(n3392), .Z(n1484) );
  CND2X1 U3532 ( .A(n1463), .B(n1484), .Z(n3620) );
  CNIVX2 U3533 ( .A(n1417), .Z(n3393) );
  CEOX2 U3534 ( .A(n1433), .B(n1431), .Z(n3394) );
  CEOX2 U3535 ( .A(n3394), .B(n1427), .Z(n1421) );
  CND2X1 U3536 ( .A(n1427), .B(n1431), .Z(n3395) );
  CND2XL U3537 ( .A(n1427), .B(n1433), .Z(n3396) );
  CND2XL U3538 ( .A(n1431), .B(n1433), .Z(n3397) );
  CND3XL U3539 ( .A(n3395), .B(n3396), .C(n3397), .Z(n1420) );
  CEO3XL U3540 ( .A(n1425), .B(n1421), .C(n1423), .Z(n1417) );
  COND2X1 U3541 ( .A(n144), .B(n2282), .C(n2281), .D(n3173), .Z(n1768) );
  CND3X2 U3542 ( .A(n3666), .B(n3667), .C(n3668), .Z(n1214) );
  CND2X1 U3543 ( .A(n1286), .B(n1261), .Z(n3792) );
  CND2X1 U3544 ( .A(n1089), .B(n1112), .Z(n3578) );
  CENX1 U3545 ( .A(n3976), .B(n3924), .Z(n2586) );
  CENX1 U3546 ( .A(n2785), .B(n3924), .Z(n2587) );
  CEOX2 U3547 ( .A(n3678), .B(n3045), .Z(n1247) );
  CND2X1 U3548 ( .A(n1278), .B(n1251), .Z(n3679) );
  CEO3X1 U3549 ( .A(n1371), .B(n1369), .C(n1394), .Z(n1365) );
  CND2X1 U3550 ( .A(n1371), .B(n1369), .Z(n3398) );
  CND2XL U3551 ( .A(n1371), .B(n1394), .Z(n3399) );
  CND3X2 U3552 ( .A(n3398), .B(n3399), .C(n3400), .Z(n1364) );
  CEOX2 U3553 ( .A(n1341), .B(n1339), .Z(n3401) );
  CND2XL U3554 ( .A(n1341), .B(n1339), .Z(n3402) );
  CND2X1 U3555 ( .A(n1341), .B(n1364), .Z(n3403) );
  CND2XL U3556 ( .A(n1335), .B(n1362), .Z(n3405) );
  CND2XL U3557 ( .A(n1335), .B(n1337), .Z(n3406) );
  CND2XL U3558 ( .A(n1362), .B(n1337), .Z(n3407) );
  CND3X1 U3559 ( .A(n3405), .B(n3406), .C(n3407), .Z(n1332) );
  CND2X2 U3560 ( .A(n1333), .B(n1360), .Z(n568) );
  CEO3X2 U3561 ( .A(n1309), .B(n1334), .C(n1307), .Z(n3781) );
  CENX1 U3562 ( .A(n3975), .B(n3897), .Z(n2687) );
  CENX2 U3563 ( .A(n3408), .B(n1211), .Z(n1199) );
  CND2XL U3564 ( .A(n3878), .B(n3660), .Z(n3894) );
  CNR2X1 U3565 ( .A(n671), .B(n674), .Z(n669) );
  CENXL U3566 ( .A(n3964), .B(n3985), .Z(n2734) );
  COND2X1 U3567 ( .A(net21352), .B(n2540), .C(net19215), .D(n2539), .Z(n2013)
         );
  CND2X1 U3568 ( .A(n1278), .B(n1253), .Z(n3680) );
  CEOX2 U3569 ( .A(n1407), .B(n1405), .Z(n3409) );
  CEOX2 U3570 ( .A(n3409), .B(n1424), .Z(n1395) );
  CND2X1 U3571 ( .A(n1424), .B(n1405), .Z(n3410) );
  CND2X1 U3572 ( .A(n1424), .B(n1407), .Z(n3411) );
  CND2XL U3573 ( .A(n1405), .B(n1407), .Z(n3412) );
  CND3X1 U3574 ( .A(n3410), .B(n3411), .C(n3412), .Z(n1394) );
  CND2X2 U3575 ( .A(n1083), .B(n1106), .Z(n494) );
  CEO3X2 U3576 ( .A(n1044), .B(n1023), .C(n1025), .Z(n1019) );
  CND2XL U3577 ( .A(n1044), .B(n1023), .Z(n3413) );
  CND2X1 U3578 ( .A(n1044), .B(n1025), .Z(n3414) );
  CND2XL U3579 ( .A(n1020), .B(n1001), .Z(n3416) );
  CND2XL U3580 ( .A(n1020), .B(n1018), .Z(n3417) );
  CND2XL U3581 ( .A(n1001), .B(n1018), .Z(n3418) );
  CND3X1 U3582 ( .A(n3416), .B(n3417), .C(n3418), .Z(n996) );
  CEO3X2 U3583 ( .A(n1457), .B(n1453), .C(n1455), .Z(n1445) );
  CND2XL U3584 ( .A(n1457), .B(n1455), .Z(n3419) );
  CND2XL U3585 ( .A(n1457), .B(n1453), .Z(n3420) );
  CND2X1 U3586 ( .A(n1455), .B(n1453), .Z(n3421) );
  CND3X1 U3587 ( .A(n3419), .B(n3420), .C(n3421), .Z(n1444) );
  CFA1X1 U3588 ( .A(n2021), .B(n2176), .CI(n2083), .CO(n1650), .S(n1651) );
  CNR2IX1 U3589 ( .B(n3979), .A(net19216), .Z(n2021) );
  CND2XL U3590 ( .A(n1419), .B(n1442), .Z(n3675) );
  CND2XL U3591 ( .A(n1134), .B(n1111), .Z(n3951) );
  CANR1X2 U3592 ( .A(n686), .B(n3915), .C(n681), .Z(n679) );
  COND2XL U3593 ( .A(net21344), .B(n2422), .C(net21744), .D(n2421), .Z(n1900)
         );
  CENXL U3594 ( .A(n3965), .B(net21909), .Z(n3424) );
  COND2XL U3595 ( .A(net21696), .B(n2326), .C(net22007), .D(n2325), .Z(n1809)
         );
  CENX1 U3596 ( .A(n1063), .B(n1084), .Z(n3673) );
  CIVXL U3597 ( .A(n3329), .Z(n1035) );
  COND2XL U3598 ( .A(net21696), .B(n2330), .C(net22006), .D(n2329), .Z(n1813)
         );
  CFA1XL U3599 ( .A(n824), .B(n1805), .CI(n1774), .CO(n816), .S(n817) );
  CIVX1 U3600 ( .A(n824), .Z(n825) );
  CENX1 U3601 ( .A(n3967), .B(n3999), .Z(n2498) );
  CIVXL U3602 ( .A(n1966), .Z(n3496) );
  CIVX1 U3603 ( .A(a[10]), .Z(n3471) );
  CEO3X1 U3604 ( .A(n1789), .B(n2025), .C(n1846), .Z(n1031) );
  CND2XL U3605 ( .A(n1846), .B(n2025), .Z(n3427) );
  CND3X1 U3606 ( .A(n3426), .B(n3427), .C(n3428), .Z(n1030) );
  CND2X1 U3607 ( .A(n1217), .B(n1219), .Z(n3667) );
  CEOX2 U3608 ( .A(n1549), .B(n1564), .Z(n3429) );
  CND2XL U3609 ( .A(n1547), .B(n1564), .Z(n3430) );
  CND2XL U3610 ( .A(n1547), .B(n1549), .Z(n3431) );
  CND2X1 U3611 ( .A(n1564), .B(n1549), .Z(n3432) );
  CND3XL U3612 ( .A(n3430), .B(n3431), .C(n3432), .Z(n1544) );
  CENX1 U3613 ( .A(n2785), .B(n3897), .Z(n2686) );
  CND2XL U3614 ( .A(n1434), .B(n1411), .Z(n3434) );
  CND2X1 U3615 ( .A(n1434), .B(n2101), .Z(n3435) );
  CND2XL U3616 ( .A(n1411), .B(n2101), .Z(n3436) );
  CND3X1 U3617 ( .A(n3434), .B(n3435), .C(n3436), .Z(n1400) );
  CNIVX4 U3618 ( .A(n48), .Z(n3437) );
  CIVXL U3619 ( .A(n48), .Z(n3997) );
  CENX2 U3620 ( .A(n1283), .B(n1281), .Z(n3638) );
  CENX2 U3621 ( .A(n3986), .B(a[2]), .Z(n2826) );
  CIVX4 U3622 ( .A(n3986), .Z(n3984) );
  CEO3X2 U3623 ( .A(n1532), .B(n1515), .C(n3261), .Z(n1509) );
  CND2XL U3624 ( .A(n1532), .B(n1530), .Z(n3438) );
  CND2XL U3625 ( .A(n1532), .B(n1515), .Z(n3439) );
  CND2XL U3626 ( .A(n1530), .B(n1515), .Z(n3440) );
  CND3X1 U3627 ( .A(n3438), .B(n3439), .C(n3440), .Z(n1508) );
  CENX1 U3628 ( .A(n3967), .B(n3924), .Z(n2597) );
  CENX1 U3629 ( .A(n3966), .B(n3924), .Z(n2598) );
  COND2X1 U3630 ( .A(n99), .B(n2428), .C(net21744), .D(n2427), .Z(n1034) );
  CIVX1 U3631 ( .A(n1188), .Z(n3833) );
  CIVXL U3632 ( .A(n764), .Z(n3442) );
  CEO3X1 U3633 ( .A(n2134), .B(n2041), .C(n2103), .Z(n1451) );
  CND2XL U3634 ( .A(n3446), .B(n2103), .Z(n3443) );
  CND2XL U3635 ( .A(n3446), .B(n2041), .Z(n3444) );
  CND3X1 U3636 ( .A(n3443), .B(n3444), .C(n3445), .Z(n1450) );
  COND2XL U3637 ( .A(n3953), .B(n2661), .C(n3803), .D(n2660), .Z(n3446) );
  CND2X1 U3638 ( .A(n3804), .B(n3805), .Z(n3447) );
  CND2X2 U3639 ( .A(n3804), .B(n3805), .Z(n2814) );
  CND2XL U3640 ( .A(n1827), .B(n1855), .Z(n3512) );
  CND2IXL U3641 ( .B(n3979), .A(n3923), .Z(n2614) );
  COND2X1 U3642 ( .A(net21344), .B(n2443), .C(net21744), .D(n2442), .Z(n1920)
         );
  CIVX3 U3643 ( .A(n12), .Z(n3986) );
  CIVX1 U3644 ( .A(a[18]), .Z(n3703) );
  COR2X1 U3645 ( .A(n460), .B(n444), .Z(n3448) );
  CND2X2 U3646 ( .A(n754), .B(n753), .Z(n460) );
  CEO3XL U3647 ( .A(n961), .B(n959), .C(n976), .Z(n3449) );
  CND2X1 U3648 ( .A(n1161), .B(n1163), .Z(n3849) );
  COND2X1 U3649 ( .A(n3328), .B(n2435), .C(net21744), .D(n2434), .Z(n1912) );
  CENX1 U3650 ( .A(n2798), .B(net21909), .Z(n2303) );
  CIVX2 U3651 ( .A(n3940), .Z(n3941) );
  COND1X2 U3652 ( .A(n544), .B(n3945), .C(n541), .Z(n535) );
  CND2X1 U3653 ( .A(n1062), .B(n1043), .Z(n3450) );
  CND2X1 U3654 ( .A(n1062), .B(n1064), .Z(n3451) );
  CND2X1 U3655 ( .A(n1043), .B(n1064), .Z(n3452) );
  CND3X2 U3656 ( .A(n3450), .B(n3451), .C(n3452), .Z(n1038) );
  CEO3X2 U3657 ( .A(n1970), .B(n1851), .C(n1184), .Z(n1153) );
  CFA1X1 U3658 ( .A(n2092), .B(n2123), .CI(n1764), .CO(n1156), .S(n1157) );
  CENX1 U3659 ( .A(n3975), .B(n3990), .Z(n2654) );
  CENX1 U3660 ( .A(n2810), .B(net19302), .Z(n2579) );
  COND2X1 U3661 ( .A(n3228), .B(n2579), .C(n3660), .D(n2578), .Z(n2052) );
  CNR2IXL U3662 ( .B(n3979), .A(n33), .Z(n2153) );
  COR2X1 U3663 ( .A(n2670), .B(n33), .Z(n3482) );
  CENXL U3664 ( .A(n3967), .B(net21419), .Z(n2300) );
  CENXL U3665 ( .A(n3973), .B(net21419), .Z(n2293) );
  CND2X1 U3666 ( .A(n3574), .B(n3575), .Z(n1893) );
  CENXL U3667 ( .A(n3958), .B(net18517), .Z(n2410) );
  CENXL U3668 ( .A(n3965), .B(net18517), .Z(n2403) );
  CENXL U3669 ( .A(n3959), .B(net18517), .Z(n2409) );
  CENXL U3670 ( .A(n3961), .B(net18517), .Z(n2407) );
  CENXL U3671 ( .A(n2809), .B(net18517), .Z(n2413) );
  CENXL U3672 ( .A(n3962), .B(net18517), .Z(n2406) );
  CENXL U3673 ( .A(n3963), .B(net18517), .Z(n2405) );
  CENXL U3674 ( .A(n3964), .B(net18517), .Z(n2404) );
  CND2XL U3675 ( .A(n774), .B(n634), .Z(n192) );
  CNR2IXL U3676 ( .B(n561), .A(n3442), .Z(n554) );
  CND2X1 U3677 ( .A(n1347), .B(n1370), .Z(n3649) );
  CND2XL U3678 ( .A(n3509), .B(n1287), .Z(n3456) );
  CND2X1 U3679 ( .A(n3454), .B(n3455), .Z(n3457) );
  CND2X2 U3680 ( .A(n3456), .B(n3457), .Z(n1281) );
  CIVX1 U3681 ( .A(n3509), .Z(n3454) );
  CIVXL U3682 ( .A(n1287), .Z(n3455) );
  CIVXL U3683 ( .A(n461), .Z(net22641) );
  CIVX1 U3684 ( .A(net22641), .Z(net22642) );
  CANR1X2 U3685 ( .A(n753), .B(n3423), .C(n467), .Z(n461) );
  CENX2 U3686 ( .A(n3066), .B(n3628), .Z(n1133) );
  CANR1XL U3687 ( .A(n561), .B(n3860), .C(n3784), .Z(n560) );
  COND2X1 U3688 ( .A(net21312), .B(n2357), .C(net21512), .D(n2356), .Z(n1839)
         );
  CIVX1 U3689 ( .A(n3335), .Z(n418) );
  COND2XL U3690 ( .A(net21434), .B(n2292), .C(net19192), .D(n2291), .Z(n1777)
         );
  COND1X1 U3691 ( .A(net22511), .B(n461), .C(n3239), .Z(n3460) );
  CIVXL U3692 ( .A(n384), .Z(n382) );
  COND2X1 U3693 ( .A(n3954), .B(n2652), .C(n3803), .D(n2651), .Z(n2125) );
  COND2X2 U3694 ( .A(n3954), .B(n2654), .C(n3803), .D(n2653), .Z(n2127) );
  CIVX2 U3695 ( .A(n84), .Z(net20818) );
  COND2X1 U3696 ( .A(net21801), .B(n2477), .C(net21846), .D(n2476), .Z(n1952)
         );
  COND1X1 U3697 ( .A(n504), .B(n512), .C(n505), .Z(n3461) );
  COND1X1 U3698 ( .A(n504), .B(n512), .C(n505), .Z(n499) );
  CENX1 U3699 ( .A(n3965), .B(net18555), .Z(n2568) );
  CIVX1 U3700 ( .A(n1061), .Z(n3580) );
  CENX1 U3701 ( .A(n3462), .B(n1439), .Z(n1437) );
  COND2X1 U3702 ( .A(n3344), .B(n2494), .C(n3941), .D(n2493), .Z(n1969) );
  CND2XL U3703 ( .A(n2237), .B(n1732), .Z(n3464) );
  CND2X1 U3704 ( .A(n2144), .B(n1732), .Z(n3465) );
  CND3X2 U3705 ( .A(n3463), .B(n3464), .C(n3465), .Z(n1636) );
  CEOX2 U3706 ( .A(n1638), .B(n1634), .Z(n3466) );
  CEOX2 U3707 ( .A(n3466), .B(n1636), .Z(n1619) );
  CND2XL U3708 ( .A(n1638), .B(n1634), .Z(n3467) );
  CND2XL U3709 ( .A(n1638), .B(n1636), .Z(n3468) );
  CND2XL U3710 ( .A(n1634), .B(n1636), .Z(n3469) );
  CND3X1 U3711 ( .A(n3467), .B(n3468), .C(n3469), .Z(n1618) );
  COND2X1 U3712 ( .A(n3551), .B(net22186), .C(n3660), .D(n2581), .Z(n1733) );
  CIVXL U3713 ( .A(n690), .Z(n689) );
  CND2X2 U3714 ( .A(n751), .B(n3906), .Z(n444) );
  COND2XL U3715 ( .A(n3228), .B(n2572), .C(n3618), .D(n2571), .Z(n2045) );
  CENX1 U3716 ( .A(n3966), .B(net20996), .Z(n2268) );
  CNR2X2 U3717 ( .A(n3325), .B(n1082), .Z(n3599) );
  CIVX1 U3718 ( .A(n3084), .Z(n3470) );
  CND2XL U3719 ( .A(n1451), .B(n1476), .Z(n3474) );
  CND2XL U3720 ( .A(n1451), .B(n1474), .Z(n3475) );
  CND2X1 U3721 ( .A(n1476), .B(n1474), .Z(n3476) );
  CND3X1 U3722 ( .A(n3474), .B(n3475), .C(n3476), .Z(n1446) );
  CFA1XL U3723 ( .A(n2197), .B(n2166), .CI(n1951), .CO(n1476), .S(n1477) );
  CND2X1 U3724 ( .A(n1361), .B(n1386), .Z(n573) );
  CENXL U3725 ( .A(n2792), .B(n3998), .Z(n2495) );
  CNIVX2 U3726 ( .A(n2054), .Z(n3477) );
  CND2X2 U3727 ( .A(n776), .B(n3909), .Z(n636) );
  CND2XL U3728 ( .A(n3989), .B(a[4]), .Z(n3479) );
  CND2X2 U3729 ( .A(n3479), .B(n3480), .Z(n2825) );
  CIVXL U3730 ( .A(a[4]), .Z(n3478) );
  COR2X1 U3731 ( .A(n3954), .B(n2671), .Z(n3481) );
  CND2X2 U3732 ( .A(n3481), .B(n3482), .Z(n2144) );
  CENXL U3733 ( .A(n3962), .B(n3991), .Z(n3483) );
  CENX1 U3734 ( .A(n3961), .B(n3991), .Z(n2671) );
  COND2XL U3735 ( .A(net21312), .B(n2354), .C(net21512), .D(n2353), .Z(n1837)
         );
  CAOR1XL U3736 ( .A(net21512), .B(net21311), .C(n2351), .Z(n1834) );
  COND2XL U3737 ( .A(net21311), .B(n2355), .C(net21512), .D(n2354), .Z(n1838)
         );
  COND2XL U3738 ( .A(n2352), .B(net21512), .C(n2353), .D(net21311), .Z(n1836)
         );
  COND2XL U3739 ( .A(n2352), .B(net21312), .C(net21512), .D(n2351), .Z(n1835)
         );
  CNR2IX1 U3740 ( .B(n3979), .A(net21512), .Z(n1863) );
  CND2X2 U3741 ( .A(n1041), .B(n3484), .Z(n3485) );
  CND2X2 U3742 ( .A(n3485), .B(n3486), .Z(n3661) );
  CIVX2 U3743 ( .A(n1060), .Z(n3484) );
  CIVX8 U3744 ( .A(n3935), .Z(n3936) );
  CDLY1XL U3745 ( .A(n633), .Z(n3487) );
  CIVX2 U3746 ( .A(n1479), .Z(n3528) );
  CFA1X1 U3747 ( .A(n1760), .B(n2057), .CI(n1080), .CO(n1056), .S(n1057) );
  CND2XL U3748 ( .A(n1213), .B(n1211), .Z(n3488) );
  CND2XL U3749 ( .A(n1211), .B(n1205), .Z(n3489) );
  CND2XL U3750 ( .A(n1213), .B(n1205), .Z(n3490) );
  CND3X1 U3751 ( .A(n3488), .B(n3489), .C(n3490), .Z(n1198) );
  CND2X1 U3752 ( .A(n1198), .B(n1175), .Z(n3708) );
  CENX1 U3753 ( .A(n2782), .B(net19314), .Z(n2452) );
  CEOX1 U3754 ( .A(n1430), .B(n1428), .Z(n3491) );
  CEOX1 U3755 ( .A(n3491), .B(n1432), .Z(n1399) );
  CND2XL U3756 ( .A(n1432), .B(n1428), .Z(n3492) );
  CND2XL U3757 ( .A(n1432), .B(n1430), .Z(n3493) );
  CND2XL U3758 ( .A(n1428), .B(n1430), .Z(n3494) );
  CND3X1 U3759 ( .A(n3492), .B(n3493), .C(n3494), .Z(n1398) );
  CENX2 U3760 ( .A(n3975), .B(net19314), .Z(n2456) );
  COND2XL U3761 ( .A(n3749), .B(n90), .C(net22327), .D(n2467), .Z(n3495) );
  CIVX2 U3762 ( .A(n3496), .Z(n3497) );
  CHA1X1 U3763 ( .A(n1726), .B(n1832), .CO(n1410), .S(n1411) );
  CIVX3 U3764 ( .A(n39), .Z(n3498) );
  CIVX3 U3765 ( .A(n39), .Z(n3995) );
  CND2X1 U3766 ( .A(n1305), .B(n1332), .Z(n559) );
  CENX1 U3767 ( .A(n2798), .B(n3994), .Z(n2633) );
  COND2XL U3768 ( .A(n3876), .B(n2742), .C(n3934), .D(n2741), .Z(n2215) );
  COND2XL U3769 ( .A(n3876), .B(n2734), .C(n3934), .D(n2733), .Z(n2207) );
  CAOR1XL U3770 ( .A(n3934), .B(n3876), .C(n2714), .Z(n2187) );
  COND2XL U3771 ( .A(n18), .B(n2736), .C(n3934), .D(n2735), .Z(n2209) );
  COND2XL U3772 ( .A(n18), .B(n2739), .C(n3933), .D(n2738), .Z(n2212) );
  COND2XL U3773 ( .A(n3876), .B(n2743), .C(n3933), .D(n2742), .Z(n2216) );
  COND2XL U3774 ( .A(n2745), .B(n3876), .C(n3933), .D(n2744), .Z(n2218) );
  COND2X1 U3775 ( .A(n2715), .B(n3933), .C(n2716), .D(n3876), .Z(n2189) );
  CFA1XL U3776 ( .A(n2153), .B(n2215), .CI(n2184), .CO(n1714), .S(n1715) );
  CND2XL U3777 ( .A(n1292), .B(n1298), .Z(n3502) );
  CND2XL U3778 ( .A(n1300), .B(n1298), .Z(n3503) );
  CND3X1 U3779 ( .A(n3501), .B(n3502), .C(n3503), .Z(n1258) );
  CENXL U3780 ( .A(n3963), .B(n3996), .Z(n2603) );
  CENXL U3781 ( .A(n3965), .B(n3996), .Z(n2601) );
  CENXL U3782 ( .A(n3957), .B(n3996), .Z(n2609) );
  CENXL U3783 ( .A(n3969), .B(n3996), .Z(n2595) );
  CENXL U3784 ( .A(net18979), .B(n3996), .Z(n2599) );
  CNIVX12 U3785 ( .A(n3084), .Z(n3923) );
  CND2XL U3786 ( .A(n1264), .B(n1266), .Z(n3560) );
  CND2XL U3787 ( .A(net22050), .B(n3703), .Z(n3705) );
  CEOX1 U3788 ( .A(n1856), .B(n2066), .Z(n3504) );
  CND2X1 U3789 ( .A(n1828), .B(n2066), .Z(n3505) );
  CND2X1 U3790 ( .A(n1828), .B(n1856), .Z(n3506) );
  CND2X1 U3791 ( .A(n2066), .B(n1856), .Z(n3507) );
  CND3X2 U3792 ( .A(n3505), .B(n3506), .C(n3507), .Z(n1294) );
  CND2X1 U3793 ( .A(n1135), .B(n1137), .Z(n3829) );
  COND2X1 U3794 ( .A(n3328), .B(n2433), .C(net21744), .D(n2432), .Z(n1910) );
  COND2X1 U3795 ( .A(n18), .B(n2725), .C(n3933), .D(n2724), .Z(n2198) );
  CND2XL U3796 ( .A(n1170), .B(n1172), .Z(n3818) );
  CENX1 U3797 ( .A(n2798), .B(net19309), .Z(n2534) );
  CENXL U3798 ( .A(n3962), .B(net18555), .Z(n2571) );
  CND2IXL U3799 ( .B(n3979), .A(net19302), .Z(n2581) );
  CENXL U3800 ( .A(n3966), .B(net19302), .Z(n2565) );
  CENX1 U3801 ( .A(n2798), .B(net19302), .Z(n3623) );
  CEOX2 U3802 ( .A(n3508), .B(net19314), .Z(n2475) );
  CNR2X1 U3803 ( .A(n3448), .B(n3335), .Z(n414) );
  CNR2XL U3804 ( .A(n353), .B(n224), .Z(n222) );
  CND2X2 U3805 ( .A(n3906), .B(n751), .Z(net22511) );
  COR2X2 U3806 ( .A(n995), .B(n1014), .Z(n3906) );
  CND2X1 U3807 ( .A(n1979), .B(n2009), .Z(n3607) );
  CEO3X2 U3808 ( .A(n1943), .B(n1855), .C(n1827), .Z(n1269) );
  CND2XL U3809 ( .A(n3495), .B(n1827), .Z(n3510) );
  CND2XL U3810 ( .A(n3495), .B(n1855), .Z(n3511) );
  COND2X1 U3811 ( .A(n2613), .B(n3250), .C(n3145), .D(n2612), .Z(n2086) );
  COND2X1 U3812 ( .A(n90), .B(n2465), .C(n87), .D(n2464), .Z(n1940) );
  CND2X1 U3813 ( .A(n1195), .B(n1222), .Z(n3513) );
  CND2X1 U3814 ( .A(n1195), .B(n1197), .Z(n3514) );
  CND2XL U3815 ( .A(n1222), .B(n1197), .Z(n3515) );
  CND3X2 U3816 ( .A(n3513), .B(n3514), .C(n3515), .Z(n1190) );
  CEOX2 U3817 ( .A(n1509), .B(n1526), .Z(n3516) );
  CEOX2 U3818 ( .A(n3516), .B(n1507), .Z(n1505) );
  CND2XL U3819 ( .A(n1507), .B(n1526), .Z(n3517) );
  CND2XL U3820 ( .A(n1507), .B(n1509), .Z(n3518) );
  CND2XL U3821 ( .A(n1526), .B(n1509), .Z(n3519) );
  CEOX2 U3822 ( .A(n1926), .B(n2108), .Z(n3520) );
  CEOX2 U3823 ( .A(n3520), .B(n1985), .Z(n1561) );
  CND2XL U3824 ( .A(n1985), .B(n2108), .Z(n3521) );
  CND2X1 U3825 ( .A(n1985), .B(n1926), .Z(n3522) );
  CND2X1 U3826 ( .A(n2108), .B(n1926), .Z(n3523) );
  CND3X1 U3827 ( .A(n3521), .B(n3522), .C(n3523), .Z(n1560) );
  CNR2IX1 U3828 ( .B(n3979), .A(net21744), .Z(n1926) );
  COND2X1 U3829 ( .A(n3344), .B(n2512), .C(n3941), .D(n2511), .Z(n1986) );
  COND2X1 U3830 ( .A(n3871), .B(n2513), .C(n3651), .D(n2512), .Z(n1987) );
  COND2XL U3831 ( .A(n3344), .B(n2491), .C(n3942), .D(n2490), .Z(n1966) );
  CND2XL U3832 ( .A(n1254), .B(n1227), .Z(n3524) );
  CND2X1 U3833 ( .A(n1227), .B(n1229), .Z(n3526) );
  CND2X2 U3834 ( .A(n3529), .B(n3530), .Z(n3762) );
  CIVX2 U3835 ( .A(n1475), .Z(n3527) );
  CIVXL U3836 ( .A(n356), .Z(net22471) );
  CEO3X2 U3837 ( .A(n2014), .B(n2138), .C(n2169), .Z(n1539) );
  CEOX2 U3838 ( .A(n1554), .B(n1541), .Z(n3531) );
  CEOX2 U3839 ( .A(n3531), .B(n1539), .Z(n1531) );
  CND2XL U3840 ( .A(n3538), .B(n2138), .Z(n3532) );
  CND2XL U3841 ( .A(n3538), .B(n2169), .Z(n3533) );
  CND2X1 U3842 ( .A(n2138), .B(n2169), .Z(n3534) );
  CND3X1 U3843 ( .A(n3532), .B(n3533), .C(n3534), .Z(n1538) );
  CND2XL U3844 ( .A(n1554), .B(n1541), .Z(n3535) );
  CND2XL U3845 ( .A(n1554), .B(n1539), .Z(n3536) );
  CND2X1 U3846 ( .A(n1541), .B(n1539), .Z(n3537) );
  CND3X1 U3847 ( .A(n3535), .B(n3536), .C(n3537), .Z(n1530) );
  COND2XL U3848 ( .A(n2541), .B(net21353), .C(net19216), .D(n2540), .Z(n3538)
         );
  COND2XL U3849 ( .A(net21353), .B(n2541), .C(net19216), .D(n2540), .Z(n2014)
         );
  CEO3X1 U3850 ( .A(n1055), .B(n1057), .C(n1053), .Z(n1045) );
  CND2XL U3851 ( .A(n1055), .B(n1053), .Z(n3539) );
  CND2XL U3852 ( .A(n1055), .B(n1057), .Z(n3540) );
  CND2X1 U3853 ( .A(n1053), .B(n1057), .Z(n3541) );
  CND3X1 U3854 ( .A(n3539), .B(n3540), .C(n3541), .Z(n1044) );
  CNIVX1 U3855 ( .A(n3285), .Z(net21249) );
  CND2XL U3856 ( .A(n1898), .B(n1751), .Z(n3542) );
  CND2XL U3857 ( .A(n1898), .B(n1869), .Z(n3543) );
  CND2XL U3858 ( .A(n1751), .B(n1869), .Z(n3544) );
  CND3XL U3859 ( .A(n3542), .B(n3543), .C(n3544), .Z(n886) );
  CNR2XL U3860 ( .A(n3328), .B(n2420), .Z(n3545) );
  CNR2XL U3861 ( .A(net21744), .B(n2419), .Z(n3546) );
  COR2X1 U3862 ( .A(n3545), .B(n3546), .Z(n1898) );
  CENXL U3863 ( .A(n2782), .B(n3925), .Z(n2419) );
  CIVXL U3864 ( .A(n3931), .Z(n3547) );
  CIVX1 U3865 ( .A(n3547), .Z(n3548) );
  CENX1 U3866 ( .A(n3972), .B(n3926), .Z(n2426) );
  CENX1 U3867 ( .A(n3971), .B(n3988), .Z(n2691) );
  CENXL U3868 ( .A(n3970), .B(net19309), .Z(n2527) );
  CIVX2 U3869 ( .A(n3659), .Z(n4000) );
  CND2X1 U3870 ( .A(n855), .B(n866), .Z(n351) );
  CIVXL U3871 ( .A(n3990), .Z(n3549) );
  CIVX2 U3872 ( .A(n3946), .Z(n3990) );
  CND3X2 U3873 ( .A(n3689), .B(n3690), .C(n3691), .Z(n1256) );
  CND2X1 U3874 ( .A(n1269), .B(n1265), .Z(n3689) );
  CND2X2 U3875 ( .A(n3878), .B(n3660), .Z(n3551) );
  CND2XL U3876 ( .A(n3499), .B(n1504), .Z(n3552) );
  CEO3X2 U3877 ( .A(n1957), .B(n2141), .C(n3559), .Z(n1595) );
  CND2X1 U3878 ( .A(n1957), .B(n2141), .Z(n3553) );
  CND2X1 U3879 ( .A(n1957), .B(n3559), .Z(n3554) );
  CND2X1 U3880 ( .A(n2141), .B(n3559), .Z(n3555) );
  CND3X2 U3881 ( .A(n3553), .B(n3554), .C(n3555), .Z(n1594) );
  CND2X1 U3882 ( .A(n1606), .B(n1595), .Z(n3557) );
  CND2XL U3883 ( .A(n1591), .B(n1595), .Z(n3558) );
  CND3X1 U3884 ( .A(n3556), .B(n3558), .C(n3557), .Z(n1586) );
  CNIVX2 U3885 ( .A(n2017), .Z(n3559) );
  COND2XL U3886 ( .A(net21352), .B(n2544), .C(net19215), .D(n2543), .Z(n2017)
         );
  CND2X1 U3887 ( .A(n1264), .B(n1272), .Z(n3561) );
  CND2XL U3888 ( .A(n1266), .B(n1272), .Z(n3562) );
  CND3X1 U3889 ( .A(n3560), .B(n3561), .C(n3562), .Z(n1230) );
  COND2X1 U3890 ( .A(n3755), .B(n2759), .C(n6), .D(n2758), .Z(n2232) );
  CND3X1 U3891 ( .A(n3662), .B(n3663), .C(n3664), .Z(n1036) );
  CND2X2 U3892 ( .A(a[14]), .B(net22399), .Z(n3563) );
  CND2X1 U3893 ( .A(net18547), .B(net22398), .Z(n3564) );
  CND2X2 U3894 ( .A(n3563), .B(n3564), .Z(net21896) );
  CIVXL U3895 ( .A(a[14]), .Z(net22398) );
  COND2XL U3896 ( .A(n72), .B(n2529), .C(net19215), .D(n2528), .Z(n3565) );
  CND2X1 U3897 ( .A(n1159), .B(n1186), .Z(n3797) );
  CNIVXL U3898 ( .A(net18547), .Z(net22262) );
  CEOX2 U3899 ( .A(n1567), .B(n1582), .Z(n3566) );
  CEOX2 U3900 ( .A(n3566), .B(n1565), .Z(n1563) );
  CND2XL U3901 ( .A(n1565), .B(n1582), .Z(n3567) );
  CND2X1 U3902 ( .A(n1565), .B(n1567), .Z(n3568) );
  CND2XL U3903 ( .A(n1582), .B(n1567), .Z(n3569) );
  CND3XL U3904 ( .A(n3567), .B(n3568), .C(n3569), .Z(n1562) );
  CEO3X1 U3905 ( .A(n1573), .B(n1590), .C(n1575), .Z(n1569) );
  CND2XL U3906 ( .A(n1573), .B(n1575), .Z(n3570) );
  CND2XL U3907 ( .A(n1573), .B(n1590), .Z(n3571) );
  CND2X1 U3908 ( .A(n1575), .B(n1590), .Z(n3572) );
  CND3X1 U3909 ( .A(n3570), .B(n3571), .C(n3572), .Z(n1568) );
  CND2X1 U3910 ( .A(n3631), .B(n3632), .Z(n1565) );
  CIVX1 U3911 ( .A(n1569), .Z(n3634) );
  CNR2X2 U3912 ( .A(n1107), .B(n3141), .Z(n504) );
  CENX2 U3913 ( .A(n3907), .B(n1109), .Z(n1107) );
  CENX2 U3914 ( .A(n1111), .B(n1134), .Z(n3907) );
  CENXL U3915 ( .A(n3967), .B(n3994), .Z(n2630) );
  CENX1 U3916 ( .A(n3977), .B(n3923), .Z(n2582) );
  COND2X2 U3917 ( .A(n3189), .B(n2272), .C(net22439), .D(n2271), .Z(n1758) );
  CENX1 U3918 ( .A(n3966), .B(n3897), .Z(n2697) );
  CEOXL U3919 ( .A(n2198), .B(n2167), .Z(n3719) );
  COND2X1 U3920 ( .A(n27), .B(n2694), .C(n3930), .D(n2693), .Z(n2167) );
  CEOX2 U3921 ( .A(n1728), .B(n1893), .Z(n1503) );
  CIVX2 U3922 ( .A(n3573), .Z(n1502) );
  CND2X1 U3923 ( .A(n1728), .B(n1893), .Z(n3573) );
  COR2XL U3924 ( .A(n2415), .B(n108), .Z(n3574) );
  COR2XL U3925 ( .A(net21248), .B(n2414), .Z(n3575) );
  COND2X1 U3926 ( .A(n108), .B(net18521), .C(net21248), .D(n2416), .Z(n1728)
         );
  CENXL U3927 ( .A(n2810), .B(net18517), .Z(n2414) );
  CND3X1 U3928 ( .A(n3814), .B(n3815), .C(n3816), .Z(n1244) );
  CENX1 U3929 ( .A(n3976), .B(n3897), .Z(n2685) );
  CIVX2 U3930 ( .A(net18521), .Z(net18519) );
  CIVX2 U3931 ( .A(net18521), .Z(net18515) );
  CENX2 U3932 ( .A(n1137), .B(n1160), .Z(n3628) );
  COND2X1 U3933 ( .A(n3755), .B(n2763), .C(n6), .D(n2762), .Z(n2236) );
  CND2X1 U3934 ( .A(n1641), .B(n1652), .Z(n672) );
  COND2X1 U3935 ( .A(n3953), .B(n2672), .C(n3803), .D(n2671), .Z(n2145) );
  CND2X1 U3936 ( .A(n1110), .B(n1089), .Z(n3576) );
  CND2X1 U3937 ( .A(n1110), .B(n1112), .Z(n3577) );
  CND3X2 U3938 ( .A(n3576), .B(n3577), .C(n3578), .Z(n1084) );
  CND2X1 U3939 ( .A(n3425), .B(n1061), .Z(n3581) );
  CND2X2 U3940 ( .A(n3579), .B(n3580), .Z(n3582) );
  CIVX2 U3941 ( .A(n3673), .Z(n3579) );
  CND2X2 U3942 ( .A(net21683), .B(net21684), .Z(n3808) );
  CIVXL U3943 ( .A(n3212), .Z(net22351) );
  CANR1XL U3944 ( .A(n658), .B(n667), .C(n659), .Z(n657) );
  CIVXL U3945 ( .A(n3988), .Z(n3583) );
  CIVX1 U3946 ( .A(n424), .Z(n749) );
  CND2X1 U3947 ( .A(n939), .B(n956), .Z(n425) );
  CIVXL U3948 ( .A(n3212), .Z(net22344) );
  CND2XL U3949 ( .A(n1311), .B(n1336), .Z(n3584) );
  CND2XL U3950 ( .A(n1311), .B(n1313), .Z(n3585) );
  CND3X1 U3951 ( .A(n3584), .B(n3586), .C(n3585), .Z(n1306) );
  CEO3X2 U3952 ( .A(n1342), .B(n1319), .C(n1317), .Z(n1311) );
  CND2X1 U3953 ( .A(n1342), .B(n1317), .Z(n3587) );
  CND2XL U3954 ( .A(n1342), .B(n1319), .Z(n3588) );
  CND3X2 U3955 ( .A(n3587), .B(n3588), .C(n3589), .Z(n1310) );
  CENX2 U3956 ( .A(n3590), .B(n1389), .Z(n1387) );
  CIVX2 U3957 ( .A(net22241), .Z(net22097) );
  CND2X1 U3958 ( .A(a[26]), .B(n3129), .Z(n3807) );
  CFA1X1 U3959 ( .A(n2112), .B(n2019), .CI(n2236), .CO(n1622), .S(n1623) );
  COND2X1 U3960 ( .A(n27), .B(n2701), .C(n3931), .D(n2700), .Z(n2174) );
  CIVXL U3961 ( .A(n458), .Z(n456) );
  CND2X2 U3962 ( .A(n1133), .B(n1158), .Z(n512) );
  CENX1 U3963 ( .A(n3963), .B(net19268), .Z(n2372) );
  CIVX2 U3964 ( .A(n21), .Z(n3734) );
  CENXL U3965 ( .A(n3969), .B(n3998), .Z(n2496) );
  CENXL U3966 ( .A(n3963), .B(n3999), .Z(n2504) );
  CENXL U3967 ( .A(n2798), .B(n3999), .Z(n2501) );
  CENXL U3968 ( .A(net18979), .B(n3999), .Z(n2500) );
  CENXL U3969 ( .A(n2785), .B(n3999), .Z(n2488) );
  CIVX2 U3970 ( .A(n643), .Z(n776) );
  COND1X1 U3971 ( .A(n643), .B(n649), .C(n3875), .Z(n642) );
  CNR2X2 U3972 ( .A(n1581), .B(n1596), .Z(n643) );
  COND2X1 U3973 ( .A(n27), .B(n2703), .C(n3931), .D(n2702), .Z(n2176) );
  COND2X1 U3974 ( .A(n3905), .B(n2678), .C(n3803), .D(n2677), .Z(n2151) );
  COND2X1 U3975 ( .A(net21344), .B(n2437), .C(n96), .D(n2436), .Z(n1914) );
  CND2XL U3976 ( .A(n2827), .B(n6), .Z(n3754) );
  CEOX1 U3977 ( .A(n3591), .B(n3595), .Z(n1267) );
  CND2XL U3978 ( .A(n1914), .B(n1884), .Z(n3592) );
  CND2XL U3979 ( .A(n1914), .B(n2003), .Z(n3593) );
  CND2XL U3980 ( .A(n1884), .B(n2003), .Z(n3594) );
  CND3X1 U3981 ( .A(n3592), .B(n3593), .C(n3594), .Z(n1266) );
  CNIVX1 U3982 ( .A(n1914), .Z(n3595) );
  COND2X1 U3983 ( .A(net21353), .B(n2527), .C(net19216), .D(n2526), .Z(n2001)
         );
  CND2X1 U3984 ( .A(n1287), .B(n1314), .Z(n3596) );
  CND2X1 U3985 ( .A(n1287), .B(n1289), .Z(n3597) );
  CEO3X1 U3986 ( .A(n1585), .B(n1583), .C(n1598), .Z(n3874) );
  COR2XL U3987 ( .A(net19215), .B(n3617), .Z(n3746) );
  CEO3X1 U3988 ( .A(n1013), .B(n1011), .C(n1009), .Z(n1003) );
  CND2XL U3989 ( .A(n3198), .B(n1009), .Z(n3600) );
  CND2XL U3990 ( .A(n3198), .B(n1011), .Z(n3601) );
  CND2X1 U3991 ( .A(n1009), .B(n1011), .Z(n3602) );
  CND3X1 U3992 ( .A(n3600), .B(n3601), .C(n3602), .Z(n1002) );
  CIVX1 U3993 ( .A(n4007), .Z(n4006) );
  CIVX3 U3994 ( .A(n3940), .Z(n3651) );
  CNR2X2 U3995 ( .A(n3098), .B(n1652), .Z(n671) );
  CIVX2 U3996 ( .A(n641), .Z(n639) );
  CENX1 U3997 ( .A(n3962), .B(n3923), .Z(n2604) );
  CEO3X1 U3998 ( .A(n1220), .B(n1218), .C(n3665), .Z(n3879) );
  CENX1 U3999 ( .A(n3973), .B(n3925), .Z(n2425) );
  CENXL U4000 ( .A(n3972), .B(n3990), .Z(n2657) );
  CENXL U4001 ( .A(n3973), .B(n3990), .Z(n2656) );
  CENXL U4002 ( .A(n3974), .B(n3990), .Z(n2655) );
  CENXL U4003 ( .A(n3970), .B(n3990), .Z(n2659) );
  CENXL U4004 ( .A(n3976), .B(n3990), .Z(n2652) );
  CENXL U4005 ( .A(n2792), .B(n3990), .Z(n2660) );
  CENXL U4006 ( .A(n3971), .B(n3990), .Z(n2658) );
  CENXL U4007 ( .A(n2783), .B(n3990), .Z(n2651) );
  CENX1 U4008 ( .A(n2785), .B(n3990), .Z(n2653) );
  COND2XL U4009 ( .A(net21802), .B(n2455), .C(net21846), .D(n2454), .Z(n1932)
         );
  CND3X2 U4010 ( .A(n3706), .B(n3707), .C(n3708), .Z(n1166) );
  CIVX1 U4011 ( .A(n644), .Z(n646) );
  CND2IXL U4012 ( .B(n3979), .A(n3982), .Z(n2779) );
  CENXL U4013 ( .A(n2798), .B(n3982), .Z(n2765) );
  CENXL U4014 ( .A(n3968), .B(n3982), .Z(n2761) );
  CENXL U4015 ( .A(n3964), .B(n3982), .Z(n2767) );
  CENXL U4016 ( .A(net18979), .B(n3982), .Z(n2764) );
  CENXL U4017 ( .A(n3965), .B(n3982), .Z(n2766) );
  CENXL U4018 ( .A(n3969), .B(n3982), .Z(n2760) );
  CENXL U4019 ( .A(n3966), .B(n3982), .Z(n2763) );
  CENX2 U4020 ( .A(n1442), .B(n1440), .Z(n3603) );
  CND2XL U4021 ( .A(n1391), .B(n1389), .Z(n3604) );
  CND2X1 U4022 ( .A(n1389), .B(n1414), .Z(n3605) );
  CND2XL U4023 ( .A(n1391), .B(n1414), .Z(n3606) );
  CND3XL U4024 ( .A(n3604), .B(n3605), .C(n3606), .Z(n1386) );
  CEO3X1 U4025 ( .A(n1979), .B(n2164), .C(n2009), .Z(n1429) );
  CND2XL U4026 ( .A(n1979), .B(n2164), .Z(n3608) );
  CND2X1 U4027 ( .A(n2009), .B(n2164), .Z(n3609) );
  CNR2X1 U4028 ( .A(n1361), .B(n1386), .Z(n572) );
  CND2X1 U4029 ( .A(n3745), .B(n3746), .Z(n2009) );
  CFA1XL U4030 ( .A(n1961), .B(n955), .CI(n1932), .CO(n948), .S(n949) );
  CND2X1 U4031 ( .A(n1221), .B(n1248), .Z(n3735) );
  CIVXL U4032 ( .A(n491), .Z(n756) );
  CND2X1 U4033 ( .A(n3638), .B(n1308), .Z(n3611) );
  CND2X2 U4034 ( .A(n3611), .B(n3612), .Z(n1277) );
  CIVX2 U4035 ( .A(n3638), .Z(n3610) );
  CENX1 U4036 ( .A(n3965), .B(n3991), .Z(n2667) );
  CNR2X2 U4037 ( .A(n1159), .B(n1186), .Z(n3741) );
  COND2XL U4038 ( .A(n3953), .B(n2669), .C(n3803), .D(n2668), .Z(n2142) );
  COND2XL U4039 ( .A(n3905), .B(n2675), .C(n3803), .D(n2674), .Z(n2148) );
  COND2XL U4040 ( .A(n2679), .B(n3904), .C(n3803), .D(n2678), .Z(n2152) );
  COND2XL U4041 ( .A(n3953), .B(n2656), .C(n3803), .D(n2655), .Z(n2129) );
  COND2XL U4042 ( .A(n3953), .B(n2677), .C(n3803), .D(n2676), .Z(n2150) );
  CND2XL U4043 ( .A(n1160), .B(n1137), .Z(n3830) );
  COND2X1 U4044 ( .A(n54), .B(n2590), .C(n3453), .D(n2589), .Z(n2063) );
  CEOX2 U4045 ( .A(n3613), .B(n1190), .Z(n1161) );
  CND2X1 U4046 ( .A(n1190), .B(n1165), .Z(n3614) );
  CND2X1 U4047 ( .A(n1190), .B(n1192), .Z(n3615) );
  CND2XL U4048 ( .A(n1165), .B(n1192), .Z(n3616) );
  CND3X2 U4049 ( .A(n3614), .B(n3615), .C(n3616), .Z(n1160) );
  CND2X1 U4050 ( .A(n1160), .B(n1135), .Z(n3828) );
  CENXL U4051 ( .A(n3965), .B(net19309), .Z(n3617) );
  CIVX4 U4052 ( .A(n3868), .Z(n3991) );
  CIVX2 U4053 ( .A(n3935), .Z(n3618) );
  CND2XL U4054 ( .A(n1425), .B(n1421), .Z(n3713) );
  CND3X1 U4055 ( .A(n3713), .B(n3714), .C(n3715), .Z(n1416) );
  COND1X1 U4056 ( .A(n697), .B(n693), .C(n694), .Z(n692) );
  CND2XL U4057 ( .A(n1245), .B(n1274), .Z(n3852) );
  COND2XL U4058 ( .A(n3871), .B(n2486), .C(n3941), .D(n2485), .Z(n1961) );
  CIVX2 U4059 ( .A(net21438), .Z(net22242) );
  COND2X1 U4060 ( .A(n63), .B(n2577), .C(n3660), .D(n2576), .Z(n2050) );
  CND2X1 U4061 ( .A(n975), .B(n994), .Z(n449) );
  CEOX2 U4062 ( .A(n1465), .B(n1484), .Z(n3619) );
  CEOX2 U4063 ( .A(n3619), .B(n1463), .Z(n1461) );
  CND2X1 U4064 ( .A(n1463), .B(n1465), .Z(n3621) );
  CND2X2 U4065 ( .A(n1437), .B(n1460), .Z(n603) );
  COND2XL U4066 ( .A(n2484), .B(n3871), .C(n3941), .D(n2483), .Z(n1959) );
  CENXL U4067 ( .A(n3965), .B(n3769), .Z(n2436) );
  CENXL U4068 ( .A(n3957), .B(n3769), .Z(n2444) );
  CEOX1 U4069 ( .A(n3743), .B(n1429), .Z(n1423) );
  CND3X1 U4070 ( .A(n3821), .B(n3822), .C(n3823), .Z(n1422) );
  CND2XL U4071 ( .A(n1421), .B(n1423), .Z(n3715) );
  CND3X2 U4072 ( .A(n3766), .B(n3767), .C(n3768), .Z(n1436) );
  CND2X1 U4073 ( .A(n1439), .B(n1441), .Z(n3767) );
  CIVX4 U4074 ( .A(net20818), .Z(net19068) );
  CENXL U4075 ( .A(n3977), .B(n3897), .Z(n2681) );
  CENX1 U4076 ( .A(n3963), .B(net21910), .Z(n2306) );
  CFA1XL U4077 ( .A(n1872), .B(n1813), .CI(n1784), .CO(n934), .S(n935) );
  CENXL U4078 ( .A(net22220), .B(net21622), .Z(n2567) );
  COND2X1 U4079 ( .A(net21344), .B(n2446), .C(net21744), .D(n2445), .Z(n1923)
         );
  CND2X1 U4080 ( .A(n1260), .B(n1237), .Z(n3625) );
  CND2X1 U4081 ( .A(n1260), .B(n1241), .Z(n3626) );
  CND2XL U4082 ( .A(n1237), .B(n1241), .Z(n3627) );
  CND3X2 U4083 ( .A(n3625), .B(n3626), .C(n3627), .Z(n1224) );
  COND2XL U4084 ( .A(n54), .B(n2611), .C(n3145), .D(n2610), .Z(n2084) );
  CAOR1XL U4085 ( .A(n3453), .B(n54), .C(n2582), .Z(n2055) );
  CIVX2 U4086 ( .A(n3831), .Z(n3868) );
  COND2X1 U4087 ( .A(n3871), .B(n2500), .C(n3941), .D(n2499), .Z(n1974) );
  CIVX1 U4088 ( .A(n1184), .Z(n1185) );
  CEOX1 U4089 ( .A(n1143), .B(n1141), .Z(n3709) );
  CENXL U4090 ( .A(n2781), .B(n3896), .Z(n2319) );
  CENXL U4091 ( .A(n3974), .B(n3896), .Z(n2325) );
  CENXL U4092 ( .A(n3970), .B(n3896), .Z(n2329) );
  CENXL U4093 ( .A(n2785), .B(n3896), .Z(n2323) );
  CENXL U4094 ( .A(n3975), .B(n3896), .Z(n2324) );
  CENXL U4095 ( .A(n2782), .B(n3896), .Z(n2320) );
  CENXL U4096 ( .A(n3971), .B(n3896), .Z(n2328) );
  CENXL U4097 ( .A(n3972), .B(n3896), .Z(n2327) );
  CENXL U4098 ( .A(n3973), .B(n3896), .Z(n2326) );
  CENXL U4099 ( .A(n3976), .B(n3896), .Z(n2322) );
  CENXL U4100 ( .A(n2783), .B(n3896), .Z(n2321) );
  CANR1X2 U4101 ( .A(n349), .B(n3914), .C(n340), .Z(n334) );
  CIVXL U4102 ( .A(n334), .Z(n332) );
  CENXL U4103 ( .A(n3968), .B(n4000), .Z(n2497) );
  CENXL U4104 ( .A(n3957), .B(n4000), .Z(n2510) );
  CENXL U4105 ( .A(n3964), .B(n4000), .Z(n2503) );
  CND2X1 U4106 ( .A(n3677), .B(n1584), .Z(n3631) );
  CND2X2 U4107 ( .A(n3629), .B(n3630), .Z(n3632) );
  CIVX2 U4108 ( .A(n3677), .Z(n3629) );
  CIVXL U4109 ( .A(n1584), .Z(n3630) );
  CND2X1 U4110 ( .A(n1571), .B(n1569), .Z(n3635) );
  CND2X2 U4111 ( .A(n3633), .B(n3634), .Z(n3636) );
  CND2X2 U4112 ( .A(n3635), .B(n3636), .Z(n3677) );
  CIVXL U4113 ( .A(n1571), .Z(n3633) );
  CIVX1 U4114 ( .A(n511), .Z(n758) );
  CND2X1 U4115 ( .A(n1613), .B(n1626), .Z(n661) );
  CND2X1 U4116 ( .A(n1338), .B(n1340), .Z(n3840) );
  CND3X2 U4117 ( .A(n3647), .B(n3648), .C(n3649), .Z(n1338) );
  COND2X1 U4118 ( .A(n3228), .B(n2561), .C(n3618), .D(n2560), .Z(n2034) );
  COND2X1 U4119 ( .A(net21433), .B(n3752), .C(net19193), .D(n2312), .Z(n1798)
         );
  CNR2X1 U4120 ( .A(n1107), .B(n3141), .Z(n3637) );
  CNIVX2 U4121 ( .A(a[14]), .Z(net22190) );
  CAOR1XL U4122 ( .A(n3085), .B(n144), .C(n2252), .Z(n1740) );
  COND2XL U4123 ( .A(n2253), .B(n3189), .C(n3086), .D(n2252), .Z(n794) );
  COND2XL U4124 ( .A(n2253), .B(n3085), .C(n2254), .D(n144), .Z(n1741) );
  COND2XL U4125 ( .A(n144), .B(n2255), .C(n3086), .D(n2254), .Z(n800) );
  COND2XL U4126 ( .A(n144), .B(n2257), .C(n3085), .D(n2256), .Z(n1743) );
  COND2XL U4127 ( .A(n144), .B(n2258), .C(n3086), .D(n2257), .Z(n1744) );
  CIVXL U4128 ( .A(net19302), .Z(net22186) );
  CIVX8 U4129 ( .A(net21622), .Z(net19302) );
  CEO3X1 U4130 ( .A(n2038), .B(n1977), .C(n2100), .Z(n3639) );
  CEO3X1 U4131 ( .A(n2038), .B(n1977), .C(n2100), .Z(n1377) );
  COND2X1 U4132 ( .A(n81), .B(n2503), .C(n3651), .D(n2502), .Z(n1977) );
  CIVX12 U4133 ( .A(n3802), .Z(n3803) );
  CENX2 U4134 ( .A(n3969), .B(n3992), .Z(n2661) );
  CND2X2 U4135 ( .A(n3785), .B(net21846), .Z(n3887) );
  CND2XL U4136 ( .A(n1017), .B(n1038), .Z(n3640) );
  CND2X1 U4137 ( .A(n1017), .B(n1019), .Z(n3641) );
  CND2XL U4138 ( .A(n1038), .B(n1019), .Z(n3642) );
  CND3XL U4139 ( .A(n3640), .B(n3641), .C(n3642), .Z(n1014) );
  CND2X1 U4140 ( .A(n995), .B(n1014), .Z(n458) );
  CND2X1 U4141 ( .A(n1162), .B(n1139), .Z(n3643) );
  CND3X2 U4142 ( .A(n3643), .B(n3644), .C(n3645), .Z(n1134) );
  CEOX2 U4143 ( .A(n1370), .B(n1347), .Z(n3646) );
  CEOX2 U4144 ( .A(n3646), .B(n1345), .Z(n1339) );
  CND2X1 U4145 ( .A(n1345), .B(n1347), .Z(n3647) );
  CND2X1 U4146 ( .A(n1345), .B(n1370), .Z(n3648) );
  CND3X2 U4147 ( .A(n3853), .B(n3854), .C(n3855), .Z(n1370) );
  CEO3X2 U4148 ( .A(n1315), .B(n1338), .C(n1340), .Z(n1309) );
  CENXL U4149 ( .A(n3979), .B(n3988), .Z(n2712) );
  CENXL U4150 ( .A(n2792), .B(n3897), .Z(n2693) );
  CENXL U4151 ( .A(n3974), .B(n3897), .Z(n2688) );
  CENXL U4152 ( .A(n3969), .B(n3897), .Z(n2694) );
  CANR1X1 U4153 ( .A(n3100), .B(n659), .C(n654), .Z(n652) );
  CIVX2 U4154 ( .A(n78), .Z(n3940) );
  CENX2 U4155 ( .A(net18979), .B(net19302), .Z(n2566) );
  CEOX1 U4156 ( .A(n3652), .B(n3748), .Z(n1305) );
  CND2XL U4157 ( .A(n3748), .B(n1334), .Z(n3653) );
  CND2XL U4158 ( .A(n3748), .B(n1309), .Z(n3654) );
  CND2XL U4159 ( .A(n1334), .B(n1309), .Z(n3655) );
  CND3X1 U4160 ( .A(n3653), .B(n3654), .C(n3655), .Z(n1304) );
  CND2XL U4161 ( .A(n1366), .B(n1368), .Z(n3656) );
  CND2XL U4162 ( .A(n1366), .B(n1343), .Z(n3657) );
  CND2X1 U4163 ( .A(n1368), .B(n1343), .Z(n3658) );
  CEO3X1 U4164 ( .A(n1313), .B(n3323), .C(n1311), .Z(n3748) );
  CIVX2 U4165 ( .A(n75), .Z(n4001) );
  COND2X2 U4166 ( .A(n3189), .B(n2281), .C(n3085), .D(n2280), .Z(n1767) );
  CENXL U4167 ( .A(n2783), .B(n3980), .Z(n2750) );
  CENXL U4168 ( .A(n2782), .B(n3980), .Z(n2749) );
  CENXL U4169 ( .A(n3975), .B(n3980), .Z(n2753) );
  CENXL U4170 ( .A(n3974), .B(n3980), .Z(n2754) );
  CENXL U4171 ( .A(n3971), .B(n3980), .Z(n2757) );
  CENXL U4172 ( .A(n2785), .B(n3980), .Z(n2752) );
  CENXL U4173 ( .A(n3972), .B(n3980), .Z(n2756) );
  CENX1 U4174 ( .A(n3962), .B(net19286), .Z(n2307) );
  CND3X1 U4175 ( .A(n3730), .B(n3731), .C(n3732), .Z(n1360) );
  CND2XL U4176 ( .A(n1039), .B(n1060), .Z(n3662) );
  CND2X1 U4177 ( .A(n1039), .B(n1041), .Z(n3663) );
  CND2XL U4178 ( .A(n1060), .B(n1041), .Z(n3664) );
  CIVX4 U4179 ( .A(n3995), .Z(n3993) );
  CND2X2 U4180 ( .A(n1461), .B(n1482), .Z(n606) );
  CEO3XL U4181 ( .A(n1201), .B(n3115), .C(n3131), .Z(n3665) );
  CNR2IX1 U4182 ( .B(n3979), .A(n3941), .Z(n1989) );
  CND2XL U4183 ( .A(n1246), .B(n1219), .Z(n3668) );
  CND2X2 U4184 ( .A(n3669), .B(n3670), .Z(n3672) );
  CND2X2 U4185 ( .A(n3671), .B(n3672), .Z(n1217) );
  CND3X2 U4186 ( .A(n3679), .B(n3680), .C(n3681), .Z(n1246) );
  CIVXL U4187 ( .A(n3487), .Z(n774) );
  CAOR1XL U4188 ( .A(net22006), .B(net21696), .C(n2318), .Z(n1803) );
  COND2XL U4189 ( .A(n2319), .B(net21696), .C(net22007), .D(n2318), .Z(n1804)
         );
  COND2XL U4190 ( .A(n2319), .B(net22006), .C(n2320), .D(net21696), .Z(n1805)
         );
  COND2XL U4191 ( .A(net21696), .B(n2321), .C(net22007), .D(n2320), .Z(n824)
         );
  COND2XL U4192 ( .A(net21696), .B(n2324), .C(net22006), .D(n2323), .Z(n1807)
         );
  COND2XL U4193 ( .A(net21696), .B(n2322), .C(net22007), .D(n2321), .Z(n1806)
         );
  CENXL U4194 ( .A(n2809), .B(n3788), .Z(n2446) );
  CENXL U4195 ( .A(n3961), .B(n4003), .Z(n2440) );
  CIVX2 U4196 ( .A(n1080), .Z(n1081) );
  CENX1 U4197 ( .A(n2781), .B(n3984), .Z(n2715) );
  CND2XL U4198 ( .A(n1440), .B(n1419), .Z(n3674) );
  CND2XL U4199 ( .A(n1440), .B(n1442), .Z(n3676) );
  CND3X1 U4200 ( .A(n3674), .B(n3675), .C(n3676), .Z(n1414) );
  CEOX2 U4201 ( .A(n1253), .B(n1251), .Z(n3678) );
  COND2X1 U4202 ( .A(net21353), .B(n2520), .C(net19216), .D(n2519), .Z(n1994)
         );
  CAOR1XL U4203 ( .A(n3803), .B(n3905), .C(n2648), .Z(n2121) );
  CND2X2 U4204 ( .A(net22097), .B(a[12]), .Z(n3684) );
  CNR2X1 U4205 ( .A(n627), .B(n622), .Z(n620) );
  CIVXL U4206 ( .A(n622), .Z(n772) );
  CND2XL U4207 ( .A(n3330), .B(n2189), .Z(n3686) );
  CND2XL U4208 ( .A(n3330), .B(n1768), .Z(n3687) );
  CND2XL U4209 ( .A(n2189), .B(n1768), .Z(n3688) );
  CND3X1 U4210 ( .A(n3686), .B(n3687), .C(n3688), .Z(n1270) );
  CND2X1 U4211 ( .A(n1265), .B(n1271), .Z(n3690) );
  CND2X1 U4212 ( .A(n1269), .B(n1271), .Z(n3691) );
  CENX1 U4213 ( .A(a[4]), .B(n12), .Z(n24) );
  CEO3X2 U4214 ( .A(n1881), .B(n1852), .C(n2001), .Z(n1179) );
  CIVX2 U4215 ( .A(n471), .Z(n754) );
  COR2X1 U4216 ( .A(net21434), .B(n2312), .Z(n3900) );
  COND2X1 U4217 ( .A(n3871), .B(n2508), .C(n3651), .D(n2507), .Z(n1982) );
  CIVXL U4218 ( .A(n3140), .Z(n3788) );
  COAN1X1 U4219 ( .A(n458), .B(n448), .C(n449), .Z(n445) );
  CND2IXL U4220 ( .B(n3979), .A(net18495), .Z(n2317) );
  CND3X2 U4221 ( .A(n3735), .B(n3736), .C(n3737), .Z(n1216) );
  CND2X4 U4222 ( .A(n2822), .B(n51), .Z(n54) );
  COND2X1 U4223 ( .A(n3228), .B(n2576), .C(n3660), .D(n2575), .Z(n2049) );
  CND2X1 U4224 ( .A(n1468), .B(n1445), .Z(n3760) );
  CENX1 U4225 ( .A(n1798), .B(n2034), .Z(n1273) );
  CND2XL U4226 ( .A(n1061), .B(n1084), .Z(n3693) );
  CND2X1 U4227 ( .A(n1061), .B(n1063), .Z(n3694) );
  CND2XL U4228 ( .A(n1084), .B(n1063), .Z(n3695) );
  CND2XL U4229 ( .A(n1401), .B(n1399), .Z(n3698) );
  CND2X2 U4230 ( .A(n3696), .B(n3697), .Z(n3699) );
  CND2X2 U4231 ( .A(n3698), .B(n3699), .Z(n3789) );
  CIVXL U4232 ( .A(n1401), .Z(n3696) );
  CIVX1 U4233 ( .A(n1399), .Z(n3697) );
  CAOR1XL U4234 ( .A(n87), .B(n90), .C(n2450), .Z(n1927) );
  COND2X1 U4235 ( .A(n90), .B(n2467), .C(net21846), .D(n2466), .Z(n1942) );
  CND2XL U4236 ( .A(n1970), .B(n1184), .Z(n3700) );
  CND2XL U4237 ( .A(n1970), .B(n1851), .Z(n3701) );
  CND2XL U4238 ( .A(n1184), .B(n1851), .Z(n3702) );
  CND3X1 U4239 ( .A(n3700), .B(n3701), .C(n3702), .Z(n1152) );
  COND2X1 U4240 ( .A(n3231), .B(n2496), .C(n3941), .D(n2495), .Z(n1184) );
  CANR1X1 U4241 ( .A(n3916), .B(n707), .C(n704), .Z(n702) );
  CND2XL U4242 ( .A(net22626), .B(a[18]), .Z(n3704) );
  CND2X1 U4243 ( .A(n3704), .B(n3705), .Z(n2818) );
  CND2XL U4244 ( .A(n3793), .B(n3727), .Z(n3728) );
  COND2X1 U4245 ( .A(n3228), .B(n2565), .C(n3618), .D(n2564), .Z(n2038) );
  CEOX2 U4246 ( .A(n3709), .B(n1166), .Z(n1137) );
  CND2X1 U4247 ( .A(n1143), .B(n1166), .Z(n3711) );
  CND2X1 U4248 ( .A(n1141), .B(n1166), .Z(n3712) );
  CND3X2 U4249 ( .A(n3710), .B(n3711), .C(n3712), .Z(n1136) );
  COND1X1 U4250 ( .A(n3264), .B(n651), .C(n652), .Z(n650) );
  CND2X1 U4251 ( .A(n1425), .B(n1423), .Z(n3714) );
  CND2XL U4252 ( .A(n1395), .B(n1393), .Z(n3716) );
  CND2XL U4253 ( .A(n1395), .B(n1416), .Z(n3717) );
  CND2XL U4254 ( .A(n1393), .B(n1416), .Z(n3718) );
  CND3X1 U4255 ( .A(n3716), .B(n3717), .C(n3718), .Z(n1388) );
  CENX2 U4256 ( .A(n3960), .B(net19314), .Z(n2474) );
  CND2X4 U4257 ( .A(n2815), .B(net19281), .Z(net21312) );
  CND2XL U4258 ( .A(n2167), .B(n2012), .Z(n3720) );
  CND2XL U4259 ( .A(n2012), .B(n2198), .Z(n3721) );
  CND2XL U4260 ( .A(n2167), .B(n2198), .Z(n3722) );
  CND3X1 U4261 ( .A(n3720), .B(n3721), .C(n3722), .Z(n1498) );
  COND2X1 U4262 ( .A(net21352), .B(n2528), .C(net19216), .D(n2527), .Z(n2002)
         );
  CNR2X2 U4263 ( .A(n1083), .B(n1106), .Z(n491) );
  CND2XL U4264 ( .A(n3968), .B(net19068), .Z(n3724) );
  CND2X1 U4265 ( .A(n3723), .B(net22013), .Z(n3725) );
  CND2X1 U4266 ( .A(n3724), .B(n3725), .Z(n2464) );
  CIVXL U4267 ( .A(net19068), .Z(net22013) );
  CNIVX4 U4268 ( .A(n2794), .Z(n3968) );
  CIVX3 U4269 ( .A(n3659), .Z(n3999) );
  CENXL U4270 ( .A(n3970), .B(n3999), .Z(n2494) );
  CNR2X1 U4271 ( .A(n514), .B(n3742), .Z(net21983) );
  CND2X2 U4272 ( .A(n3726), .B(n3039), .Z(n3729) );
  CND2X2 U4273 ( .A(n3728), .B(n3729), .Z(n1219) );
  CIVX1 U4274 ( .A(n3793), .Z(n3726) );
  CIVXL U4275 ( .A(n1252), .Z(n3727) );
  CND3X2 U4276 ( .A(n3790), .B(n3791), .C(n3792), .Z(n1252) );
  CND2XL U4277 ( .A(n1363), .B(n1365), .Z(n3730) );
  CND2XL U4278 ( .A(n1363), .B(n1388), .Z(n3731) );
  CND2X1 U4279 ( .A(n1365), .B(n1388), .Z(n3732) );
  CNR2X2 U4280 ( .A(n514), .B(n3742), .Z(n478) );
  CNR2IX1 U4281 ( .B(n3979), .A(net21846), .Z(n1957) );
  CENXL U4282 ( .A(n3974), .B(net18547), .Z(n2523) );
  CNR2X1 U4283 ( .A(n514), .B(n3742), .Z(n3733) );
  CND2X1 U4284 ( .A(n1439), .B(n3112), .Z(n3766) );
  CND2X2 U4285 ( .A(n3447), .B(n3869), .Z(n126) );
  CND2X1 U4286 ( .A(n1248), .B(n1250), .Z(n3736) );
  CEO3X1 U4287 ( .A(n1191), .B(n1189), .C(n1216), .Z(n3883) );
  CNIVX4 U4288 ( .A(n2787), .Z(n3974) );
  CENXL U4289 ( .A(n3956), .B(n3897), .Z(n2709) );
  CND2IXL U4290 ( .B(n3979), .A(n3897), .Z(n2713) );
  CENXL U4291 ( .A(n3957), .B(n3897), .Z(n2708) );
  CENXL U4292 ( .A(n3964), .B(n3897), .Z(n2701) );
  CENXL U4293 ( .A(n3962), .B(n3897), .Z(n2703) );
  CENXL U4294 ( .A(n3958), .B(n3897), .Z(n2707) );
  CENXL U4295 ( .A(n2810), .B(n3897), .Z(n2711) );
  CENXL U4296 ( .A(n3965), .B(n3897), .Z(n2700) );
  CENX1 U4297 ( .A(n2783), .B(n3897), .Z(n2684) );
  CEO3X1 U4298 ( .A(n1325), .B(n1323), .C(n1348), .Z(n1315) );
  CND2XL U4299 ( .A(n1325), .B(n1323), .Z(n3738) );
  CND2X1 U4300 ( .A(n1323), .B(n1348), .Z(n3740) );
  CIVXL U4301 ( .A(net19309), .Z(net21948) );
  CIVX4 U4302 ( .A(n4004), .Z(n4003) );
  CNIVX4 U4303 ( .A(net21375), .Z(net21248) );
  CENXL U4304 ( .A(n2810), .B(n3769), .Z(n2447) );
  CENXL U4305 ( .A(n3962), .B(n3769), .Z(n2439) );
  CENXL U4306 ( .A(n2809), .B(net21910), .Z(n3750) );
  CND2X2 U4307 ( .A(n3343), .B(n3062), .Z(n3742) );
  CND2XL U4308 ( .A(n1085), .B(n1087), .Z(n3801) );
  CANR1X1 U4309 ( .A(n3733), .B(n546), .C(n3903), .Z(n3744) );
  COR2X1 U4310 ( .A(net21353), .B(n2536), .Z(n3745) );
  CANR1X1 U4311 ( .A(net21983), .B(net22598), .C(n3903), .Z(n3892) );
  CIVX2 U4312 ( .A(n3460), .Z(n441) );
  CND2X4 U4313 ( .A(n3285), .B(n2816), .Z(n108) );
  CENXL U4314 ( .A(n3969), .B(net21836), .Z(n3747) );
  CIVXL U4315 ( .A(n677), .Z(n676) );
  COND2X1 U4316 ( .A(n3787), .B(n2643), .C(n3938), .D(n2642), .Z(n2116) );
  COND2XL U4317 ( .A(net21353), .B(n2539), .C(net19215), .D(n2538), .Z(n2012)
         );
  CAOR1XL U4318 ( .A(n3941), .B(n3871), .C(n2483), .Z(n1958) );
  CIVX1 U4319 ( .A(n3983), .Z(n3981) );
  CNIVX20 U4320 ( .A(net19068), .Z(net19314) );
  CNIVX4 U4321 ( .A(net18495), .Z(net21909) );
  CNIVX4 U4322 ( .A(net18495), .Z(net21910) );
  CNIVX1 U4323 ( .A(net18495), .Z(net19286) );
  CIVX2 U4324 ( .A(n3812), .Z(n3982) );
  CENXL U4325 ( .A(n2798), .B(net21836), .Z(n3749) );
  COND2X1 U4326 ( .A(n3328), .B(n3211), .C(net21744), .D(n2449), .Z(n1729) );
  CIVX12 U4327 ( .A(net21725), .Z(net19268) );
  CNIVX4 U4328 ( .A(n2786), .Z(n3975) );
  CNIVX2 U4329 ( .A(n1316), .Z(n3751) );
  CENX1 U4330 ( .A(n3753), .B(n1247), .Z(n1245) );
  CENX1 U4331 ( .A(n1249), .B(n1276), .Z(n3753) );
  CEOX2 U4332 ( .A(net22190), .B(net18547), .Z(n2820) );
  CND2X2 U4333 ( .A(n2827), .B(n6), .Z(n3755) );
  COND1X1 U4334 ( .A(n710), .B(n708), .C(n709), .Z(n707) );
  CANR1X1 U4335 ( .A(n3912), .B(n3917), .C(n712), .Z(n710) );
  CIVXL U4336 ( .A(net19268), .Z(net21882) );
  CAOR1XL U4337 ( .A(net19216), .B(net21353), .C(n2516), .Z(n1990) );
  CND2X4 U4338 ( .A(n2823), .B(n3937), .Z(n45) );
  CEOX2 U4339 ( .A(n3998), .B(a[16]), .Z(n2819) );
  CIVX4 U4340 ( .A(n4001), .Z(n3998) );
  CENXL U4341 ( .A(n3970), .B(n3923), .Z(n3757) );
  CENX1 U4342 ( .A(n3959), .B(net21909), .Z(n2310) );
  CENXL U4343 ( .A(n3971), .B(net18547), .Z(n2526) );
  CNR2X2 U4344 ( .A(n1015), .B(n1036), .Z(n468) );
  CIVDX2 U4345 ( .A(n111), .Z0(net21859), .Z1(net21858) );
  CIVX1 U4346 ( .A(n3232), .Z(n3905) );
  CIVX4 U4347 ( .A(net21858), .Z(net21725) );
  CENXL U4348 ( .A(n2782), .B(n3984), .Z(n2716) );
  CENXL U4349 ( .A(n3975), .B(n3984), .Z(n2720) );
  CENXL U4350 ( .A(n3971), .B(n3984), .Z(n2724) );
  CENXL U4351 ( .A(n3970), .B(n3984), .Z(n2725) );
  CENXL U4352 ( .A(n2785), .B(n3984), .Z(n2719) );
  CENXL U4353 ( .A(n2792), .B(n3984), .Z(n2726) );
  COND2X1 U4354 ( .A(n27), .B(n2684), .C(n3930), .D(n2683), .Z(n2157) );
  COND2XL U4355 ( .A(n2712), .B(n27), .C(n3931), .D(n2711), .Z(n2185) );
  COND2XL U4356 ( .A(n27), .B(n2708), .C(n3931), .D(n2707), .Z(n2181) );
  COND2XL U4357 ( .A(n27), .B(n2705), .C(n3931), .D(n2704), .Z(n2178) );
  COND2XL U4358 ( .A(n27), .B(n2704), .C(n3931), .D(n2703), .Z(n2177) );
  COND2XL U4359 ( .A(n45), .B(n2636), .C(n3938), .D(n2635), .Z(n2109) );
  COND2X1 U4360 ( .A(n81), .B(n2498), .C(n3942), .D(n2497), .Z(n1972) );
  COND2XL U4361 ( .A(n2514), .B(n3871), .C(n3651), .D(n2513), .Z(n1988) );
  COND2XL U4362 ( .A(n3344), .B(n2490), .C(n3651), .D(n2489), .Z(n1965) );
  COND2XL U4363 ( .A(n3344), .B(n2487), .C(n3651), .D(n2486), .Z(n1962) );
  CND2XL U4364 ( .A(n2100), .B(n1977), .Z(n3858) );
  CEO3X2 U4365 ( .A(n1468), .B(n3064), .C(n3053), .Z(n1441) );
  CND2X1 U4366 ( .A(n1468), .B(n1447), .Z(n3759) );
  CND2X1 U4367 ( .A(n1447), .B(n1445), .Z(n3761) );
  CND3X2 U4368 ( .A(n3761), .B(n3760), .C(n3759), .Z(n1440) );
  CEOX2 U4369 ( .A(n3762), .B(n1477), .Z(n1469) );
  CND2XL U4370 ( .A(n1477), .B(n1479), .Z(n3763) );
  CND2XL U4371 ( .A(n1477), .B(n1475), .Z(n3764) );
  CND2XL U4372 ( .A(n1479), .B(n1475), .Z(n3765) );
  CND3X1 U4373 ( .A(n3763), .B(n3764), .C(n3765), .Z(n1468) );
  COND2X1 U4374 ( .A(n2616), .B(n3787), .C(n3938), .D(n2615), .Z(n2089) );
  CND2IXL U4375 ( .B(n3979), .A(net22262), .Z(n2548) );
  CENXL U4376 ( .A(net18979), .B(net19309), .Z(n2533) );
  CENX1 U4377 ( .A(n3967), .B(net19309), .Z(n2531) );
  CNIVX4 U4378 ( .A(net18549), .Z(net19309) );
  CND2XL U4379 ( .A(n1462), .B(n1441), .Z(n3768) );
  CIVXL U4380 ( .A(n3140), .Z(n3769) );
  CIVXL U4381 ( .A(n3140), .Z(n3770) );
  CIVX2 U4382 ( .A(n93), .Z(n4004) );
  CAOR1XL U4383 ( .A(net19192), .B(net21433), .C(n2285), .Z(n1771) );
  COND2XL U4384 ( .A(net21434), .B(n2294), .C(net19192), .D(n2293), .Z(n1779)
         );
  COND2XL U4385 ( .A(n2286), .B(net19192), .C(n2287), .D(net21434), .Z(n1773)
         );
  CIVXL U4386 ( .A(n810), .Z(n811) );
  CEO3X1 U4387 ( .A(n1620), .B(n1624), .C(n1622), .Z(n1603) );
  CND2XL U4388 ( .A(n1624), .B(n1622), .Z(n3771) );
  CND2XL U4389 ( .A(n1624), .B(n1620), .Z(n3772) );
  CND2X1 U4390 ( .A(n1622), .B(n1620), .Z(n3773) );
  CND3X1 U4391 ( .A(n3771), .B(n3772), .C(n3773), .Z(n1602) );
  CEO3X2 U4392 ( .A(n1593), .B(n1602), .C(n1604), .Z(n1585) );
  CND2X1 U4393 ( .A(n1593), .B(n1602), .Z(n3774) );
  CND2X1 U4394 ( .A(n1593), .B(n1604), .Z(n3775) );
  CND2X1 U4395 ( .A(n1602), .B(n1604), .Z(n3776) );
  CND3X2 U4396 ( .A(n3774), .B(n3775), .C(n3776), .Z(n1584) );
  CND2XL U4397 ( .A(n1571), .B(n1569), .Z(n3777) );
  CND2XL U4398 ( .A(n1571), .B(n1584), .Z(n3778) );
  CND2XL U4399 ( .A(n1569), .B(n1584), .Z(n3779) );
  CND3X1 U4400 ( .A(n3777), .B(n3778), .C(n3779), .Z(n1564) );
  CIVXL U4401 ( .A(n3996), .Z(n3780) );
  CND2X2 U4402 ( .A(n3785), .B(net21846), .Z(net21801) );
  CND2X2 U4403 ( .A(net21846), .B(n3785), .Z(net21802) );
  CENX1 U4404 ( .A(n3960), .B(net18515), .Z(n2408) );
  CNIVX4 U4405 ( .A(n2804), .Z(n3960) );
  CIVXL U4406 ( .A(net21337), .Z(net21791) );
  CND2X1 U4407 ( .A(n3877), .B(n1436), .Z(n592) );
  CND2X1 U4408 ( .A(net22248), .B(net21896), .Z(n72) );
  CIVX1 U4409 ( .A(n3867), .Z(n3947) );
  CIVX4 U4410 ( .A(n3947), .Z(n3992) );
  CNIVX4 U4411 ( .A(n2791), .Z(n3970) );
  CIVX3 U4412 ( .A(n3983), .Z(n3980) );
  CNR2X2 U4413 ( .A(n1613), .B(n1626), .Z(n660) );
  COND2X1 U4414 ( .A(n3783), .B(n2764), .C(n6), .D(n2763), .Z(n2237) );
  CIVXL U4415 ( .A(n564), .Z(n3784) );
  CENXL U4416 ( .A(n3977), .B(n3999), .Z(n2483) );
  CENXL U4417 ( .A(n3979), .B(n3999), .Z(n2514) );
  CENXL U4418 ( .A(n3959), .B(n4000), .Z(n2508) );
  CENXL U4419 ( .A(n2809), .B(n3999), .Z(n2512) );
  CENXL U4420 ( .A(n3958), .B(n3999), .Z(n2509) );
  CENXL U4421 ( .A(n2810), .B(n3999), .Z(n2513) );
  CENXL U4422 ( .A(n3965), .B(n4000), .Z(n2502) );
  CND2IXL U4423 ( .B(n3979), .A(n3999), .Z(n2515) );
  CENXL U4424 ( .A(n3961), .B(n3998), .Z(n2506) );
  CENXL U4425 ( .A(n3956), .B(n3998), .Z(n2511) );
  CENXL U4426 ( .A(n3962), .B(n3998), .Z(n2505) );
  CENX1 U4427 ( .A(a[18]), .B(net22626), .Z(n3785) );
  CENX2 U4428 ( .A(net18521), .B(a[22]), .Z(n2816) );
  CND2IXL U4429 ( .B(n3979), .A(net21836), .Z(n2482) );
  CENXL U4430 ( .A(n3967), .B(net19068), .Z(n2465) );
  CENXL U4431 ( .A(n3974), .B(net19178), .Z(n3786) );
  CNIVX4 U4432 ( .A(n42), .Z(n3937) );
  COND2X1 U4433 ( .A(n126), .B(n2341), .C(net22006), .D(n2340), .Z(n1824) );
  CENX2 U4434 ( .A(n3789), .B(n1422), .Z(n1393) );
  CND2X1 U4435 ( .A(n1288), .B(n1261), .Z(n3791) );
  CND2X1 U4436 ( .A(n1225), .B(n1223), .Z(n3794) );
  CND2X1 U4437 ( .A(n1225), .B(n1252), .Z(n3795) );
  CND3X2 U4438 ( .A(n3794), .B(n3795), .C(n3796), .Z(n1218) );
  CENX2 U4439 ( .A(a[20]), .B(net19068), .Z(n96) );
  CENX2 U4440 ( .A(n3995), .B(a[8]), .Z(n2823) );
  CNIVX4 U4441 ( .A(n2795), .Z(n3967) );
  CENXL U4442 ( .A(n2792), .B(net22242), .Z(n2561) );
  CENXL U4443 ( .A(n3971), .B(net18555), .Z(n2559) );
  CENXL U4444 ( .A(n2783), .B(net22242), .Z(n2552) );
  CENXL U4445 ( .A(n3974), .B(net19178), .Z(n2556) );
  CENXL U4446 ( .A(n3970), .B(net18555), .Z(n2560) );
  CENXL U4447 ( .A(n3975), .B(net19178), .Z(n2555) );
  CENXL U4448 ( .A(n2782), .B(net19178), .Z(n2551) );
  CENXL U4449 ( .A(n2785), .B(net19178), .Z(n2554) );
  CENXL U4450 ( .A(n2781), .B(net19178), .Z(n2550) );
  COND2X1 U4451 ( .A(n2616), .B(n3939), .C(n2617), .D(n3787), .Z(n2090) );
  CNIVX4 U4452 ( .A(n78), .Z(n3798) );
  COND1X1 U4453 ( .A(n675), .B(n671), .C(n672), .Z(n670) );
  CNIVX4 U4454 ( .A(n2801), .Z(n3963) );
  COND2X2 U4455 ( .A(n90), .B(n3747), .C(n87), .D(n2462), .Z(n1130) );
  CND2XL U4456 ( .A(n1247), .B(n1249), .Z(n3815) );
  CFA1X1 U4457 ( .A(n1905), .B(n1845), .CI(n1788), .CO(n1010), .S(n1011) );
  CANR1XL U4458 ( .A(n748), .B(n415), .C(n408), .Z(n406) );
  COND2X1 U4459 ( .A(net21433), .B(n2303), .C(net19193), .D(n2302), .Z(n1788)
         );
  CND2X2 U4460 ( .A(n1187), .B(n1214), .Z(n530) );
  CEO3X2 U4461 ( .A(n1108), .B(n1087), .C(n1085), .Z(n1083) );
  CND2XL U4462 ( .A(n1108), .B(n1085), .Z(n3799) );
  CND2XL U4463 ( .A(n1108), .B(n1087), .Z(n3800) );
  CNIVX4 U4464 ( .A(n2790), .Z(n3971) );
  COND1X1 U4465 ( .A(n305), .B(net21297), .C(n306), .Z(n304) );
  COND1X1 U4466 ( .A(n257), .B(net21297), .C(n258), .Z(n256) );
  CENXL U4467 ( .A(n3978), .B(net19268), .Z(n2382) );
  CENX1 U4468 ( .A(n3971), .B(net18515), .Z(n2394) );
  CIVX8 U4469 ( .A(n3943), .Z(n3802) );
  COND2X1 U4470 ( .A(n2682), .B(n27), .C(n3930), .D(n2681), .Z(n2155) );
  CNIVX4 U4471 ( .A(n2788), .Z(n3973) );
  COND2X2 U4472 ( .A(n3787), .B(n2619), .C(n3938), .D(n2618), .Z(n2092) );
  CND2X4 U4473 ( .A(n2814), .B(n3869), .Z(net21696) );
  CENX1 U4474 ( .A(n3956), .B(n4005), .Z(n2346) );
  CENXL U4475 ( .A(n3963), .B(n3928), .Z(n2768) );
  CENXL U4476 ( .A(n3963), .B(n3985), .Z(n2735) );
  CENXL U4477 ( .A(n3963), .B(n3988), .Z(n2702) );
  COND2X1 U4478 ( .A(net21696), .B(n2339), .C(net22006), .D(n2338), .Z(n1822)
         );
  CENXL U4479 ( .A(n3963), .B(net18483), .Z(n2273) );
  CND2X1 U4480 ( .A(n1316), .B(n1291), .Z(n3809) );
  CND2X1 U4481 ( .A(n1316), .B(n1318), .Z(n3810) );
  CND2XL U4482 ( .A(n1291), .B(n1318), .Z(n3811) );
  CIVXL U4483 ( .A(n3), .Z(n3812) );
  CENXL U4484 ( .A(n3960), .B(n3924), .Z(n2606) );
  CENXL U4485 ( .A(n3960), .B(n3982), .Z(n2771) );
  CENXL U4486 ( .A(n3960), .B(n3897), .Z(n2705) );
  CENXL U4487 ( .A(n3960), .B(n3984), .Z(n2738) );
  CENXL U4488 ( .A(n3960), .B(n3990), .Z(n2672) );
  CENXL U4489 ( .A(n3960), .B(net22242), .Z(n2573) );
  CENXL U4490 ( .A(n3960), .B(net18483), .Z(n2276) );
  CENXL U4491 ( .A(n3960), .B(n4000), .Z(n2507) );
  CENX1 U4492 ( .A(n3960), .B(net21419), .Z(n2309) );
  CIVXL U4493 ( .A(n761), .Z(n3813) );
  CAOR1X1 U4494 ( .A(n6), .B(n3880), .C(n2747), .Z(n2220) );
  CND3X1 U4495 ( .A(n3848), .B(n3849), .C(n3850), .Z(n1158) );
  CND2X2 U4496 ( .A(n2824), .B(n33), .Z(n36) );
  CENX1 U4497 ( .A(a[6]), .B(n3946), .Z(n2824) );
  CND2XL U4498 ( .A(n1247), .B(n1276), .Z(n3814) );
  CND2XL U4499 ( .A(n1276), .B(n1249), .Z(n3816) );
  COND1X1 U4500 ( .A(n547), .B(n575), .C(n548), .Z(n546) );
  COND2X1 U4501 ( .A(n108), .B(n2390), .C(net21249), .D(n2389), .Z(n1870) );
  CENXL U4502 ( .A(n3975), .B(net18517), .Z(n2390) );
  CIVXL U4503 ( .A(n562), .Z(n564) );
  CND2XL U4504 ( .A(n1172), .B(n1174), .Z(n3820) );
  CND3X1 U4505 ( .A(n3818), .B(n3819), .C(n3820), .Z(n1140) );
  CIVXL U4506 ( .A(n543), .Z(n762) );
  CND3X1 U4507 ( .A(n3856), .B(n3857), .C(n3858), .Z(n1376) );
  COND2X1 U4508 ( .A(n3787), .B(n2627), .C(n3939), .D(n2626), .Z(n2100) );
  CENX1 U4509 ( .A(n3970), .B(n3993), .Z(n2626) );
  CND2XL U4510 ( .A(n2001), .B(n1852), .Z(n3846) );
  CND2XL U4511 ( .A(n1454), .B(n1429), .Z(n3821) );
  CND2XL U4512 ( .A(n1454), .B(n1435), .Z(n3822) );
  CND2XL U4513 ( .A(n1429), .B(n1435), .Z(n3823) );
  CND2XL U4514 ( .A(n1401), .B(n1399), .Z(n3824) );
  CND2X1 U4515 ( .A(n1401), .B(n1422), .Z(n3825) );
  CND2XL U4516 ( .A(n1399), .B(n1422), .Z(n3826) );
  CND3X1 U4517 ( .A(n3824), .B(n3825), .C(n3826), .Z(n1392) );
  CNIVX4 U4518 ( .A(a[6]), .Z(n3827) );
  CIVXL U4519 ( .A(n3946), .Z(n3831) );
  CND2X4 U4520 ( .A(net22248), .B(n2820), .Z(net21352) );
  CNIVX4 U4521 ( .A(net21438), .Z(net21622) );
  CENXL U4522 ( .A(n2809), .B(n3996), .Z(n2611) );
  CENXL U4523 ( .A(n2810), .B(n3996), .Z(n2612) );
  CENXL U4524 ( .A(n3961), .B(n3996), .Z(n2605) );
  CENXL U4525 ( .A(n3964), .B(n3996), .Z(n2602) );
  CENXL U4526 ( .A(n3958), .B(n3996), .Z(n2608) );
  CEOX4 U4527 ( .A(n3128), .B(a[24]), .Z(n2815) );
  CND2X1 U4528 ( .A(n1188), .B(n3832), .Z(n3835) );
  CND2X2 U4529 ( .A(n3835), .B(n3834), .Z(n3847) );
  COND2XL U4530 ( .A(net21434), .B(n2302), .C(net19192), .D(n2301), .Z(n1787)
         );
  CENXL U4531 ( .A(n2781), .B(n3993), .Z(n2616) );
  CND2XL U4532 ( .A(net18979), .B(net18519), .Z(n3836) );
  CND2X1 U4533 ( .A(net21590), .B(net21591), .Z(n3837) );
  CND2X1 U4534 ( .A(n3836), .B(n3837), .Z(n2401) );
  CIVXL U4535 ( .A(net18979), .Z(net21590) );
  CIVXL U4536 ( .A(net18519), .Z(net21591) );
  CND2X2 U4537 ( .A(n767), .B(n768), .Z(n578) );
  CND2X1 U4538 ( .A(n1315), .B(n1340), .Z(n3839) );
  CND2XL U4539 ( .A(n1283), .B(n1281), .Z(n3841) );
  CND2XL U4540 ( .A(n1281), .B(n1308), .Z(n3843) );
  CND3X1 U4541 ( .A(n3841), .B(n3842), .C(n3843), .Z(n1276) );
  CNIVX4 U4542 ( .A(n2784), .Z(n3976) );
  COND1XL U4543 ( .A(n3442), .B(n564), .C(n559), .Z(n555) );
  CAN2X1 U4544 ( .A(n764), .B(n559), .Z(n3862) );
  CND2XL U4545 ( .A(n1881), .B(n2001), .Z(n3844) );
  CND2XL U4546 ( .A(n1881), .B(n1852), .Z(n3845) );
  CND3X1 U4547 ( .A(n3844), .B(n3845), .C(n3846), .Z(n1178) );
  CIVX2 U4548 ( .A(n102), .Z(net18521) );
  CIVXL U4549 ( .A(n556), .Z(n764) );
  CEOX2 U4550 ( .A(n3847), .B(n1161), .Z(n1159) );
  CND2XL U4551 ( .A(n3441), .B(n1163), .Z(n3850) );
  CENXL U4552 ( .A(n2783), .B(n4000), .Z(n2486) );
  CENXL U4553 ( .A(n3975), .B(n4000), .Z(n2489) );
  CENXL U4554 ( .A(n2781), .B(n3999), .Z(n2484) );
  CENXL U4555 ( .A(n2782), .B(n3999), .Z(n2485) );
  CENXL U4556 ( .A(n3971), .B(n4000), .Z(n2493) );
  CENXL U4557 ( .A(n3974), .B(n4000), .Z(n2490) );
  CENXL U4558 ( .A(n3973), .B(n3999), .Z(n2491) );
  CENXL U4559 ( .A(n3972), .B(n3999), .Z(n2492) );
  CENXL U4560 ( .A(n3976), .B(n4000), .Z(n2487) );
  CIVXL U4561 ( .A(n756), .Z(n3851) );
  CNIVX4 U4562 ( .A(n2802), .Z(n3962) );
  CENXL U4563 ( .A(n3972), .B(net22242), .Z(n2558) );
  CNIVX4 U4564 ( .A(n3084), .Z(n3924) );
  COND2X1 U4565 ( .A(n108), .B(n2406), .C(net21248), .D(n2405), .Z(n1884) );
  CENX1 U4566 ( .A(a[6]), .B(n21), .Z(n33) );
  CNIVX3 U4567 ( .A(n42), .Z(n3938) );
  CIVXL U4568 ( .A(n259), .Z(n257) );
  COND2X1 U4569 ( .A(n108), .B(n2396), .C(net21249), .D(n2395), .Z(n1874) );
  CENXL U4570 ( .A(n3976), .B(n3981), .Z(n2751) );
  CENXL U4571 ( .A(n2781), .B(n3980), .Z(n2748) );
  CENXL U4572 ( .A(n3970), .B(n3980), .Z(n2758) );
  CEO3X2 U4573 ( .A(n1377), .B(n1381), .C(n1383), .Z(n1371) );
  CND2XL U4574 ( .A(n3639), .B(n1383), .Z(n3853) );
  CND2XL U4575 ( .A(n3639), .B(n1381), .Z(n3854) );
  CND2X1 U4576 ( .A(n1383), .B(n1381), .Z(n3855) );
  CND2XL U4577 ( .A(n2038), .B(n2100), .Z(n3856) );
  CND2XL U4578 ( .A(n2038), .B(n1977), .Z(n3857) );
  CENXL U4579 ( .A(n3859), .B(n3110), .Z(product[32]) );
  CAN2XL U4580 ( .A(n762), .B(n3852), .Z(n3859) );
  CAOR1XL U4581 ( .A(n3286), .B(n3882), .C(n577), .Z(n3860) );
  CIVXL U4582 ( .A(n212), .Z(product[63]) );
  CENXL U4583 ( .A(n3861), .B(net21297), .Z(product[40]) );
  CAN2XL U4584 ( .A(n754), .B(n3422), .Z(n3861) );
  CENXL U4585 ( .A(n3860), .B(n184), .Z(product[28]) );
  CENXL U4586 ( .A(n3862), .B(n560), .Z(product[30]) );
  CENXL U4587 ( .A(n3972), .B(net20996), .Z(n2261) );
  CENXL U4588 ( .A(n3973), .B(net20996), .Z(n2260) );
  CENXL U4589 ( .A(n3975), .B(net20996), .Z(n2258) );
  CENXL U4590 ( .A(n3974), .B(net20996), .Z(n2259) );
  CENXL U4591 ( .A(n3970), .B(net20996), .Z(n2263) );
  CENXL U4592 ( .A(n3971), .B(net20996), .Z(n2262) );
  CENXL U4593 ( .A(n3968), .B(net20996), .Z(n2266) );
  CENXL U4594 ( .A(n3969), .B(net20996), .Z(n2265) );
  CENXL U4595 ( .A(n2792), .B(net20996), .Z(n2264) );
  COND2X1 U4596 ( .A(n3231), .B(n2499), .C(n3942), .D(n2498), .Z(n1973) );
  CENX2 U4597 ( .A(a[16]), .B(net18549), .Z(n78) );
  CHA1X1 U4598 ( .A(n1801), .B(n1725), .CO(n1358), .S(n1359) );
  COND2X1 U4599 ( .A(n2436), .B(n99), .C(net21744), .D(n2435), .Z(n1913) );
  CENXL U4600 ( .A(n3958), .B(n3993), .Z(n2641) );
  CENXL U4601 ( .A(n2810), .B(n3993), .Z(n2645) );
  CENXL U4602 ( .A(n2809), .B(n3994), .Z(n2644) );
  CENXL U4603 ( .A(n3959), .B(n3993), .Z(n2640) );
  CENXL U4604 ( .A(n3962), .B(n3993), .Z(n2637) );
  CENXL U4605 ( .A(n3957), .B(n3993), .Z(n2642) );
  CENXL U4606 ( .A(n3956), .B(n3994), .Z(n2643) );
  CENXL U4607 ( .A(n3964), .B(n3993), .Z(n2635) );
  COND2XL U4608 ( .A(n27), .B(n2693), .C(n3930), .D(n2692), .Z(n2166) );
  CENXL U4609 ( .A(n3959), .B(net18555), .Z(n2574) );
  CENXL U4610 ( .A(n175), .B(n506), .Z(product[37]) );
  COND1XL U4611 ( .A(n507), .B(n545), .C(n508), .Z(n506) );
  CIVX1 U4612 ( .A(n546), .Z(n545) );
  CIVXL U4613 ( .A(n2232), .Z(n3865) );
  CIVX1 U4614 ( .A(n3865), .Z(n3866) );
  CIVXL U4615 ( .A(n3946), .Z(n3867) );
  CENX1 U4616 ( .A(n3964), .B(n3926), .Z(n2437) );
  COND2X1 U4617 ( .A(n3783), .B(n2756), .C(n6), .D(n2755), .Z(n2229) );
  CIVXL U4618 ( .A(n223), .Z(n221) );
  CND2X2 U4619 ( .A(n3900), .B(n3901), .Z(n1797) );
  CIVXL U4620 ( .A(n3599), .Z(n755) );
  COND1X1 U4621 ( .A(n494), .B(n484), .C(n485), .Z(n3870) );
  COND1X1 U4622 ( .A(n494), .B(n484), .C(n485), .Z(n483) );
  COND2X1 U4623 ( .A(n3250), .B(n2591), .C(n3145), .D(n2590), .Z(n2064) );
  CIVXL U4624 ( .A(n650), .Z(n649) );
  COND2X1 U4625 ( .A(n3783), .B(n2753), .C(n6), .D(n2752), .Z(n2226) );
  CENXL U4626 ( .A(n2798), .B(n3897), .Z(n2699) );
  CENXL U4627 ( .A(n3961), .B(n3897), .Z(n2704) );
  CENXL U4628 ( .A(n3959), .B(n3988), .Z(n2706) );
  CENXL U4629 ( .A(n3967), .B(n3897), .Z(n2696) );
  CENXL U4630 ( .A(n2809), .B(n3897), .Z(n2710) );
  CENXL U4631 ( .A(net18979), .B(n3897), .Z(n2698) );
  CENXL U4632 ( .A(n3968), .B(n3897), .Z(n2695) );
  CENXL U4633 ( .A(n3973), .B(n3897), .Z(n2689) );
  CND2X2 U4634 ( .A(n2813), .B(net19191), .Z(net21433) );
  CND2X4 U4635 ( .A(net19281), .B(n2815), .Z(n117) );
  COR2X1 U4636 ( .A(n1563), .B(n1580), .Z(n3873) );
  COR2XL U4637 ( .A(n1580), .B(n1563), .Z(n3909) );
  CIVXL U4638 ( .A(n573), .Z(n571) );
  CENX1 U4639 ( .A(n3969), .B(net19309), .Z(n2529) );
  COR2X1 U4640 ( .A(n1798), .B(n2034), .Z(n1272) );
  CIVXL U4641 ( .A(n646), .Z(n3875) );
  CND2X1 U4642 ( .A(n3874), .B(n1596), .Z(n644) );
  CND2X4 U4643 ( .A(n2826), .B(n3932), .Z(n3876) );
  CNR2X2 U4644 ( .A(n1413), .B(n1436), .Z(n591) );
  CEO3XL U4645 ( .A(n1417), .B(n3052), .C(n3230), .Z(n3877) );
  CND2XL U4646 ( .A(n3909), .B(n641), .Z(n193) );
  CENXL U4647 ( .A(n2810), .B(n4005), .Z(n2348) );
  CENXL U4648 ( .A(n2792), .B(n3981), .Z(n2759) );
  CANR1X2 U4649 ( .A(n3217), .B(n621), .C(n616), .Z(n614) );
  COND2XL U4650 ( .A(n3783), .B(n2771), .C(n6), .D(n2770), .Z(n2244) );
  COND2XL U4651 ( .A(n3783), .B(n2769), .C(n6), .D(n2768), .Z(n2242) );
  COND2XL U4652 ( .A(n3783), .B(n2766), .C(n6), .D(n2765), .Z(n2239) );
  COND2XL U4653 ( .A(n3783), .B(n2772), .C(n6), .D(n2771), .Z(n2245) );
  COND2XL U4654 ( .A(n3783), .B(n2761), .C(n6), .D(n2760), .Z(n2234) );
  COND2XL U4655 ( .A(n3783), .B(n2767), .C(n6), .D(n2766), .Z(n2240) );
  COND2XL U4656 ( .A(n3783), .B(n2777), .C(n6), .D(n2776), .Z(n2250) );
  CENXL U4657 ( .A(n3973), .B(net22242), .Z(n2557) );
  CENXL U4658 ( .A(n3976), .B(net22242), .Z(n2553) );
  CIVX1 U4659 ( .A(n3995), .Z(n3994) );
  CIVX2 U4660 ( .A(n120), .Z(n4007) );
  CANR1X1 U4661 ( .A(n3733), .B(net22598), .C(net21313), .Z(n149) );
  CNR2X2 U4662 ( .A(n3249), .B(n572), .Z(n561) );
  COND2XL U4663 ( .A(net21353), .B(n2533), .C(net19216), .D(n2532), .Z(n2006)
         );
  COR2X1 U4664 ( .A(net19192), .B(n2311), .Z(n3901) );
  CND2XL U4665 ( .A(n776), .B(n3875), .Z(n194) );
  CENXL U4666 ( .A(n3970), .B(net18515), .Z(n2395) );
  CENXL U4667 ( .A(n2785), .B(net18515), .Z(n2389) );
  CENXL U4668 ( .A(n2792), .B(net18515), .Z(n2396) );
  CENXL U4669 ( .A(n3973), .B(net18515), .Z(n2392) );
  CENX1 U4670 ( .A(n2783), .B(net19314), .Z(n2453) );
  CNIVX3 U4671 ( .A(n145), .Z(n3978) );
  CENXL U4672 ( .A(n3957), .B(net22242), .Z(n2576) );
  CENXL U4673 ( .A(n3956), .B(net19178), .Z(n2577) );
  CENXL U4674 ( .A(n3964), .B(net19178), .Z(n2569) );
  CENXL U4675 ( .A(n2809), .B(net19178), .Z(n2578) );
  CENXL U4676 ( .A(n3961), .B(net19178), .Z(n2572) );
  CENXL U4677 ( .A(n3963), .B(net19178), .Z(n2570) );
  CND2X4 U4678 ( .A(n2827), .B(n6), .Z(n3880) );
  COR2XL U4679 ( .A(n1304), .B(n1275), .Z(n3881) );
  CIVXL U4680 ( .A(n567), .Z(n765) );
  CIVXL U4681 ( .A(n27), .Z(n3884) );
  CIVX1 U4682 ( .A(n3884), .Z(n3885) );
  CND2X2 U4683 ( .A(n549), .B(n561), .Z(n547) );
  CENXL U4684 ( .A(n2809), .B(net19309), .Z(n2545) );
  CENXL U4685 ( .A(n3959), .B(net19309), .Z(n2541) );
  CENXL U4686 ( .A(n2810), .B(net19309), .Z(n2546) );
  CENXL U4687 ( .A(n3958), .B(net19309), .Z(n2542) );
  CENXL U4688 ( .A(n3962), .B(net19309), .Z(n2538) );
  CENXL U4689 ( .A(n3961), .B(net19309), .Z(n2539) );
  CENXL U4690 ( .A(n3963), .B(net19309), .Z(n2537) );
  CENXL U4691 ( .A(n3966), .B(net19309), .Z(n2532) );
  CENXL U4692 ( .A(n2781), .B(n3990), .Z(n2649) );
  COND2XL U4693 ( .A(n2385), .B(net21249), .C(n2386), .D(n108), .Z(n1866) );
  CAOR1XL U4694 ( .A(net21249), .B(n108), .C(n2384), .Z(n1864) );
  COND2XL U4695 ( .A(n108), .B(n2388), .C(net21249), .D(n2387), .Z(n1868) );
  COND2XL U4696 ( .A(n108), .B(n2392), .C(net21248), .D(n2391), .Z(n1872) );
  CIVXL U4697 ( .A(n530), .Z(n528) );
  CIVX2 U4698 ( .A(n3886), .Z(n767) );
  CIVXL U4699 ( .A(n529), .Z(n760) );
  CENXL U4700 ( .A(n2783), .B(net18547), .Z(n2519) );
  CENXL U4701 ( .A(n2785), .B(net18547), .Z(n2521) );
  CENXL U4702 ( .A(n3976), .B(net18547), .Z(n2520) );
  CIVXL U4703 ( .A(net22626), .Z(net21337) );
  CND2XL U4704 ( .A(n760), .B(n3327), .Z(n178) );
  CANR1X1 U4705 ( .A(n482), .B(n3461), .C(n483), .Z(n3888) );
  CANR1X1 U4706 ( .A(n3461), .B(n3063), .C(n483), .Z(n481) );
  CANR1XL U4707 ( .A(n646), .B(n3873), .C(n639), .Z(n3889) );
  COND1X2 U4708 ( .A(n578), .B(n595), .C(n579), .Z(n577) );
  CANR1X2 U4709 ( .A(n520), .B(n535), .C(n3326), .Z(n3890) );
  CANR1X1 U4710 ( .A(n520), .B(n535), .C(n3326), .Z(n3899) );
  CND2X4 U4711 ( .A(n2815), .B(net19281), .Z(net21311) );
  COND1X1 U4712 ( .A(n3742), .B(n3890), .C(n3888), .Z(net21313) );
  COND1X1 U4713 ( .A(n3742), .B(n3899), .C(n481), .Z(n3903) );
  CENXL U4714 ( .A(n3977), .B(n4005), .Z(n2318) );
  CENXL U4715 ( .A(n3964), .B(n4005), .Z(n2338) );
  CENXL U4716 ( .A(n3965), .B(n4005), .Z(n2337) );
  CENXL U4717 ( .A(n3961), .B(n4005), .Z(n2341) );
  CENXL U4718 ( .A(n3958), .B(n4005), .Z(n2344) );
  CENXL U4719 ( .A(n3962), .B(n4005), .Z(n2340) );
  CENXL U4720 ( .A(n2809), .B(n4005), .Z(n2347) );
  CENXL U4721 ( .A(n3959), .B(n4005), .Z(n2343) );
  CENXL U4722 ( .A(n3977), .B(net21909), .Z(n2285) );
  CENXL U4723 ( .A(n2781), .B(n3262), .Z(n2286) );
  CENXL U4724 ( .A(n2782), .B(net21909), .Z(n2287) );
  CENXL U4725 ( .A(n2783), .B(n3262), .Z(n2288) );
  CENXL U4726 ( .A(n3975), .B(net21909), .Z(n2291) );
  CENXL U4727 ( .A(n2785), .B(net21910), .Z(n2290) );
  CENXL U4728 ( .A(n3974), .B(n3262), .Z(n2292) );
  CENXL U4729 ( .A(n3976), .B(net21909), .Z(n2289) );
  CENXL U4730 ( .A(n3972), .B(net21909), .Z(n2294) );
  CENXL U4731 ( .A(n3970), .B(net21910), .Z(n2296) );
  CENXL U4732 ( .A(n3978), .B(net21910), .Z(n2316) );
  CENXL U4733 ( .A(net18979), .B(net21910), .Z(n2302) );
  CANR1X2 U4734 ( .A(n499), .B(n3063), .C(n3870), .Z(n3891) );
  COND2X1 U4735 ( .A(net21434), .B(n2310), .C(net19193), .D(n2309), .Z(n1795)
         );
  CND2X2 U4736 ( .A(n520), .B(n534), .Z(n514) );
  COND1X2 U4737 ( .A(n480), .B(n3890), .C(n3891), .Z(n479) );
  CENXL U4738 ( .A(n176), .B(n513), .Z(product[36]) );
  CENXL U4739 ( .A(n177), .B(n524), .Z(product[35]) );
  CENXL U4740 ( .A(n178), .B(n531), .Z(product[34]) );
  CENXL U4741 ( .A(n179), .B(n542), .Z(product[33]) );
  COND2X1 U4742 ( .A(net21434), .B(n2306), .C(net19193), .D(n2305), .Z(n1791)
         );
  CIVXL U4743 ( .A(n461), .Z(n463) );
  CND2IXL U4744 ( .B(n3979), .A(n3994), .Z(n2647) );
  CENXL U4745 ( .A(n3968), .B(n3994), .Z(n2629) );
  CENXL U4746 ( .A(net18979), .B(n3994), .Z(n2632) );
  CENXL U4747 ( .A(n470), .B(n171), .Z(product[41]) );
  COND2XL U4748 ( .A(n2286), .B(net21434), .C(net19192), .D(n2285), .Z(n1772)
         );
  COND2XL U4749 ( .A(net21433), .B(n2288), .C(net19193), .D(n2287), .Z(n810)
         );
  COND2XL U4750 ( .A(net21433), .B(n2293), .C(net19193), .D(n2292), .Z(n1778)
         );
  COND2XL U4751 ( .A(net21434), .B(n2290), .C(net19193), .D(n2289), .Z(n1775)
         );
  COND2XL U4752 ( .A(net21434), .B(n2295), .C(net19193), .D(n2294), .Z(n1780)
         );
  COND2XL U4753 ( .A(net21433), .B(n2299), .C(net19193), .D(n2298), .Z(n1784)
         );
  COND2XL U4754 ( .A(net21433), .B(n2301), .C(net19193), .D(n2300), .Z(n1786)
         );
  COND2XL U4755 ( .A(net21433), .B(n2305), .C(net19193), .D(n3424), .Z(n1790)
         );
  CENXL U4756 ( .A(n459), .B(n170), .Z(product[42]) );
  CENXL U4757 ( .A(n435), .B(n168), .Z(product[44]) );
  CENXL U4758 ( .A(n411), .B(n166), .Z(product[46]) );
  CENXL U4759 ( .A(n393), .B(n164), .Z(product[48]) );
  CENXL U4760 ( .A(n371), .B(n162), .Z(product[50]) );
  CENXL U4761 ( .A(n3972), .B(net18547), .Z(n2525) );
  CENXL U4762 ( .A(n3973), .B(net18547), .Z(n2524) );
  CENXL U4763 ( .A(n3960), .B(net19309), .Z(n2540) );
  CENXL U4764 ( .A(n3975), .B(net18547), .Z(n2522) );
  COND2X1 U4765 ( .A(n72), .B(n2529), .C(net19215), .D(n2528), .Z(n1242) );
  CENXL U4766 ( .A(n3969), .B(net18519), .Z(n2397) );
  CENXL U4767 ( .A(n2798), .B(net18519), .Z(n2402) );
  CENXL U4768 ( .A(n3968), .B(net18519), .Z(n2398) );
  CENXL U4769 ( .A(n450), .B(n169), .Z(product[43]) );
  CENXL U4770 ( .A(n426), .B(n167), .Z(product[45]) );
  CENXL U4771 ( .A(n404), .B(n165), .Z(product[47]) );
  CENXL U4772 ( .A(n380), .B(n163), .Z(product[49]) );
  CENXL U4773 ( .A(n352), .B(n161), .Z(product[51]) );
  CANR1X2 U4774 ( .A(n646), .B(n3873), .C(n639), .Z(n637) );
  CENXL U4775 ( .A(n219), .B(n150), .Z(product[62]) );
  CENXL U4776 ( .A(n343), .B(n160), .Z(product[52]) );
  CENXL U4777 ( .A(n328), .B(n159), .Z(product[53]) );
  CENXL U4778 ( .A(n317), .B(n158), .Z(product[54]) );
  CENXL U4779 ( .A(n304), .B(n157), .Z(product[55]) );
  CENXL U4780 ( .A(n280), .B(n155), .Z(product[57]) );
  CENXL U4781 ( .A(n267), .B(n154), .Z(product[58]) );
  CENXL U4782 ( .A(n256), .B(n153), .Z(product[59]) );
  CENXL U4783 ( .A(n230), .B(n151), .Z(product[61]) );
  CNIVX16 U4784 ( .A(n2806), .Z(n3958) );
  CENXL U4785 ( .A(n3958), .B(n3991), .Z(n2674) );
  CENXL U4786 ( .A(n3964), .B(n3991), .Z(n2668) );
  CENXL U4787 ( .A(n3963), .B(n3991), .Z(n2669) );
  CENXL U4788 ( .A(n3956), .B(n3991), .Z(n2676) );
  CENXL U4789 ( .A(n2810), .B(n3991), .Z(n2678) );
  CENXL U4790 ( .A(n3977), .B(n3991), .Z(n2648) );
  CENXL U4791 ( .A(n3962), .B(n3991), .Z(n2670) );
  CNIVX16 U4792 ( .A(n2805), .Z(n3959) );
  CNIVX16 U4793 ( .A(n2807), .Z(n3957) );
  CENXL U4794 ( .A(n2809), .B(n3991), .Z(n2677) );
  CENXL U4795 ( .A(n3978), .B(n3991), .Z(n2679) );
  CENXL U4796 ( .A(n3978), .B(n3984), .Z(n2745) );
  CENXL U4797 ( .A(n3978), .B(n3993), .Z(n2646) );
  CENXL U4798 ( .A(n3978), .B(net22262), .Z(n2547) );
  CENXL U4799 ( .A(n3978), .B(net19314), .Z(n2481) );
  CENXL U4800 ( .A(n3978), .B(net18517), .Z(n2415) );
  CENXL U4801 ( .A(n3978), .B(n3928), .Z(n2778) );
  CENXL U4802 ( .A(n3978), .B(n3788), .Z(n2448) );
  CENXL U4803 ( .A(n3957), .B(net18547), .Z(n2543) );
  CENXL U4804 ( .A(n3956), .B(net19309), .Z(n2544) );
  CIVX2 U4805 ( .A(n3336), .Z(net19192) );
  CNR2IX1 U4806 ( .B(n3979), .A(n3931), .Z(n2186) );
  CIVX8 U4807 ( .A(a[0]), .Z(n6) );
  CENX1 U4808 ( .A(n3957), .B(net18483), .Z(n2279) );
  CENX1 U4809 ( .A(n3957), .B(net18517), .Z(n2411) );
  CENX1 U4810 ( .A(n3957), .B(n3928), .Z(n2774) );
  CNR2X2 U4811 ( .A(n460), .B(n444), .Z(n438) );
  CENX1 U4812 ( .A(n3958), .B(net19286), .Z(n2311) );
  COND1XL U4813 ( .A(n329), .B(net19189), .C(n330), .Z(n328) );
  COND1XL U4814 ( .A(n318), .B(net19189), .C(n319), .Z(n317) );
  COND1XL U4815 ( .A(n344), .B(net19189), .C(n345), .Z(n343) );
  COND1XL U4816 ( .A(n268), .B(net19189), .C(n269), .Z(n267) );
  COND1XL U4817 ( .A(n281), .B(net19189), .C(n282), .Z(n280) );
  CIVXL U4818 ( .A(n754), .Z(n3902) );
  CND2X2 U4819 ( .A(n769), .B(n770), .Z(n594) );
  COND2X1 U4820 ( .A(n3783), .B(n2775), .C(n6), .D(n2774), .Z(n2248) );
  CENX1 U4821 ( .A(n3966), .B(net19268), .Z(n2367) );
  CNIVX8 U4822 ( .A(n2800), .Z(n3964) );
  COND2X1 U4823 ( .A(n3250), .B(n2610), .C(n3145), .D(n2609), .Z(n2083) );
  CNR2X1 U4824 ( .A(n3448), .B(n385), .Z(n383) );
  CND2X1 U4825 ( .A(n387), .B(n418), .Z(n385) );
  CND2XL U4826 ( .A(n414), .B(n3096), .Z(n394) );
  CND2X2 U4827 ( .A(net20990), .B(n749), .Z(n416) );
  CANR1X1 U4828 ( .A(n699), .B(n691), .C(n692), .Z(n690) );
  CNR2XL U4829 ( .A(n693), .B(n696), .Z(n691) );
  CND2XL U4830 ( .A(n1723), .B(n2218), .Z(n723) );
  CENXL U4831 ( .A(n3978), .B(n4005), .Z(n2349) );
  CNR2X1 U4832 ( .A(n3099), .B(n1640), .Z(n665) );
  CND2X1 U4833 ( .A(n1505), .B(n1524), .Z(n623) );
  CND2X1 U4834 ( .A(n1701), .B(n1706), .Z(n701) );
  CANR1XL U4835 ( .A(n729), .B(n3918), .C(n726), .Z(n724) );
  CENX1 U4836 ( .A(n3974), .B(net19314), .Z(n2457) );
  CENX1 U4837 ( .A(n3972), .B(net19314), .Z(n2459) );
  CENX1 U4838 ( .A(n2792), .B(net19314), .Z(n2462) );
  CENX1 U4839 ( .A(n3961), .B(net19314), .Z(n2473) );
  CENX1 U4840 ( .A(n3962), .B(net19314), .Z(n2472) );
  COND2XL U4841 ( .A(n27), .B(n3583), .C(n3930), .D(n2713), .Z(n1737) );
  CENXL U4842 ( .A(n174), .B(n495), .Z(product[38]) );
  CENXL U4843 ( .A(n486), .B(n173), .Z(product[39]) );
  CND2X1 U4844 ( .A(n620), .B(n3217), .Z(n613) );
  CND2XL U4845 ( .A(n3906), .B(n3118), .Z(n451) );
  CND2XL U4846 ( .A(n355), .B(n331), .Z(n329) );
  CIVXL U4847 ( .A(n3872), .Z(n597) );
  CND2XL U4848 ( .A(n3911), .B(n658), .Z(n651) );
  CIVX1 U4849 ( .A(n656), .Z(n654) );
  CIVXL U4850 ( .A(n383), .Z(n381) );
  CIVXL U4851 ( .A(n414), .Z(n412) );
  CEOXL U4852 ( .A(n196), .B(n662), .Z(product[16]) );
  CEOXL U4853 ( .A(n195), .B(n657), .Z(product[17]) );
  CND2XL U4854 ( .A(n3100), .B(n656), .Z(n195) );
  COND1X1 U4855 ( .A(n700), .B(n702), .C(n701), .Z(n699) );
  CND2XL U4856 ( .A(n3915), .B(n3913), .Z(n678) );
  CND2XL U4857 ( .A(n355), .B(n320), .Z(n318) );
  CND2XL U4858 ( .A(n741), .B(n327), .Z(n159) );
  CND2XL U4859 ( .A(n355), .B(n3908), .Z(n344) );
  CND2XL U4860 ( .A(n3914), .B(n342), .Z(n160) );
  CND2XL U4861 ( .A(n355), .B(n283), .Z(n281) );
  CND2XL U4862 ( .A(net20981), .B(n279), .Z(n155) );
  CEOXL U4863 ( .A(n200), .B(n684), .Z(product[12]) );
  CND2XL U4864 ( .A(n3915), .B(n683), .Z(n200) );
  CND2XL U4865 ( .A(n781), .B(n675), .Z(n199) );
  CND2XL U4866 ( .A(n785), .B(n697), .Z(n203) );
  CND2XL U4867 ( .A(n3913), .B(n688), .Z(n201) );
  CEOXL U4868 ( .A(n702), .B(n204), .Z(product[8]) );
  COND1X1 U4869 ( .A(n724), .B(n722), .C(n723), .Z(n721) );
  CIVXL U4870 ( .A(n222), .Z(n220) );
  CND2XL U4871 ( .A(n3917), .B(n714), .Z(n207) );
  CND2XL U4872 ( .A(n3918), .B(n728), .Z(n210) );
  CND2XL U4873 ( .A(n3919), .B(n720), .Z(n208) );
  CENXL U4874 ( .A(n2781), .B(net21337), .Z(n2451) );
  COND2XL U4875 ( .A(n2646), .B(n45), .C(n3938), .D(n2645), .Z(n2119) );
  CENX1 U4876 ( .A(n3968), .B(net19268), .Z(n2365) );
  CENX1 U4877 ( .A(n3967), .B(net19268), .Z(n2366) );
  CENXL U4878 ( .A(n2785), .B(n3925), .Z(n2422) );
  CENXL U4879 ( .A(n3966), .B(n3994), .Z(n2631) );
  CENXL U4880 ( .A(n3969), .B(n3994), .Z(n2628) );
  CENXL U4881 ( .A(n3974), .B(n3925), .Z(n2424) );
  CENXL U4882 ( .A(n2783), .B(n3926), .Z(n2420) );
  CENXL U4883 ( .A(n3977), .B(n3993), .Z(n2615) );
  CNIVX4 U4884 ( .A(n2793), .Z(n3969) );
  CND2XL U4885 ( .A(n516), .B(n758), .Z(n507) );
  CND2XL U4886 ( .A(n516), .B(n3343), .Z(n496) );
  CND2XL U4887 ( .A(n489), .B(n516), .Z(n487) );
  CND2XL U4888 ( .A(n751), .B(n449), .Z(n169) );
  CND2XL U4889 ( .A(n753), .B(n469), .Z(n171) );
  CANR1XL U4890 ( .A(n768), .B(n597), .C(n590), .Z(n586) );
  COND1XL U4891 ( .A(n496), .B(n545), .C(n497), .Z(n495) );
  CND2XL U4892 ( .A(n485), .B(n755), .Z(n173) );
  COND1XL U4893 ( .A(n487), .B(n545), .C(n488), .Z(n486) );
  COND1XL U4894 ( .A(n543), .B(n545), .C(n3852), .Z(n542) );
  COND1XL U4895 ( .A(n532), .B(n545), .C(n533), .Z(n531) );
  CND2XL U4896 ( .A(n768), .B(n592), .Z(n186) );
  CND2XL U4897 ( .A(n766), .B(n573), .Z(n184) );
  CND2XL U4898 ( .A(n769), .B(n603), .Z(n187) );
  CND2XL U4899 ( .A(n767), .B(n583), .Z(n185) );
  COND1XL U4900 ( .A(n585), .B(n3102), .C(n586), .Z(n584) );
  CND2XL U4901 ( .A(n596), .B(n768), .Z(n585) );
  CANR1XL U4902 ( .A(n620), .B(n629), .C(n621), .Z(n619) );
  CEOXL U4903 ( .A(n3102), .B(n188), .Z(product[24]) );
  CND2XL U4904 ( .A(n770), .B(n606), .Z(n188) );
  CNR2IXL U4905 ( .B(n3343), .A(n3851), .Z(n489) );
  CND2XL U4906 ( .A(n3906), .B(n458), .Z(n170) );
  CANR1XL U4907 ( .A(n3906), .B(n463), .C(n456), .Z(n452) );
  CND2XL U4908 ( .A(n3908), .B(n351), .Z(n161) );
  CND2XL U4909 ( .A(n749), .B(n425), .Z(n167) );
  CND2XL U4910 ( .A(net20990), .B(n438), .Z(n427) );
  CANR1XL U4911 ( .A(net20990), .B(n3460), .C(n432), .Z(n428) );
  CANR1XL U4912 ( .A(n283), .B(n356), .C(n286), .Z(n282) );
  CANR1XL U4913 ( .A(n331), .B(n356), .C(n332), .Z(n330) );
  CANR1XL U4914 ( .A(n3908), .B(n356), .C(n349), .Z(n345) );
  CND2XL U4915 ( .A(n3948), .B(n3797), .Z(n177) );
  COND1XL U4916 ( .A(n525), .B(n545), .C(n526), .Z(n524) );
  CND2XL U4917 ( .A(n773), .B(n628), .Z(n191) );
  CENX1 U4918 ( .A(n642), .B(n193), .Z(product[19]) );
  COND1XL U4919 ( .A(n636), .B(n649), .C(n3889), .Z(n635) );
  CENX1 U4920 ( .A(n667), .B(n197), .Z(product[15]) );
  CEOXL U4921 ( .A(n194), .B(n649), .Z(product[18]) );
  CND2X1 U4922 ( .A(n778), .B(n661), .Z(n196) );
  CANR1XL U4923 ( .A(n779), .B(n667), .C(n664), .Z(n662) );
  CNR2X1 U4924 ( .A(n660), .B(n665), .Z(n658) );
  CND2X1 U4925 ( .A(n1275), .B(n1304), .Z(n552) );
  CND2X1 U4926 ( .A(n1107), .B(n1132), .Z(n505) );
  CND2X1 U4927 ( .A(n1387), .B(n1412), .Z(n583) );
  CND2X1 U4928 ( .A(n1244), .B(n1215), .Z(n541) );
  CNR2XL U4929 ( .A(n333), .B(n324), .Z(n320) );
  CANR1XL U4930 ( .A(n233), .B(n356), .C(n236), .Z(n232) );
  CENX1 U4931 ( .A(n673), .B(n198), .Z(product[14]) );
  CND2X1 U4932 ( .A(n780), .B(n672), .Z(n198) );
  COND1XL U4933 ( .A(n674), .B(n676), .C(n675), .Z(n673) );
  COR2X1 U4934 ( .A(n855), .B(n866), .Z(n3908) );
  COR2X1 U4935 ( .A(n957), .B(n974), .Z(net20990) );
  COR2X1 U4936 ( .A(n291), .B(n324), .Z(n3910) );
  CND2X1 U4937 ( .A(n1627), .B(n1640), .Z(n666) );
  CND2X1 U4938 ( .A(n1563), .B(n1580), .Z(n641) );
  CND2X1 U4939 ( .A(n1597), .B(n1612), .Z(n656) );
  CENX1 U4940 ( .A(n202), .B(n695), .Z(product[10]) );
  CND2X1 U4941 ( .A(n784), .B(n694), .Z(n202) );
  COND1XL U4942 ( .A(n696), .B(n698), .C(n697), .Z(n695) );
  CENX1 U4943 ( .A(n689), .B(n201), .Z(product[11]) );
  CANR1XL U4944 ( .A(n3913), .B(n689), .C(n686), .Z(n684) );
  CEOXL U4945 ( .A(n199), .B(n676), .Z(product[13]) );
  CEOXL U4946 ( .A(n698), .B(n203), .Z(product[9]) );
  CND2X1 U4947 ( .A(n786), .B(n701), .Z(n204) );
  CND2XL U4948 ( .A(n222), .B(n3920), .Z(n213) );
  CANR1XL U4949 ( .A(n3920), .B(n223), .C(n216), .Z(n214) );
  CNR2X1 U4950 ( .A(n1653), .B(n1664), .Z(n674) );
  CND2X1 U4951 ( .A(n3920), .B(n218), .Z(n150) );
  CND2X1 U4952 ( .A(n3223), .B(n229), .Z(n151) );
  COND1XL U4953 ( .A(n231), .B(net19189), .C(n232), .Z(n230) );
  CND2X1 U4954 ( .A(n355), .B(n233), .Z(n231) );
  CNR2X1 U4955 ( .A(n1701), .B(n1706), .Z(n700) );
  CAOR1X1 U4956 ( .A(n721), .B(n3919), .C(n718), .Z(n3912) );
  COR2X1 U4957 ( .A(n1675), .B(n1684), .Z(n3913) );
  COR2X1 U4958 ( .A(n845), .B(n854), .Z(n3914) );
  COR2X1 U4959 ( .A(n1674), .B(n1665), .Z(n3915) );
  CND2X1 U4960 ( .A(n835), .B(n844), .Z(n327) );
  CND2X1 U4961 ( .A(n1653), .B(n1664), .Z(n675) );
  CND2X1 U4962 ( .A(n1693), .B(n1700), .Z(n697) );
  CND2X1 U4963 ( .A(n1675), .B(n1684), .Z(n688) );
  CND2X1 U4964 ( .A(n845), .B(n854), .Z(n342) );
  CND2X1 U4965 ( .A(n1665), .B(n1674), .Z(n683) );
  CENX1 U4966 ( .A(n205), .B(n707), .Z(product[7]) );
  CND2X1 U4967 ( .A(n3916), .B(n706), .Z(n205) );
  CENX1 U4968 ( .A(n210), .B(n729), .Z(product[2]) );
  CENX1 U4969 ( .A(n208), .B(n721), .Z(product[4]) );
  CEOXL U4970 ( .A(n710), .B(n206), .Z(product[6]) );
  CND2X1 U4971 ( .A(n788), .B(n709), .Z(n206) );
  CEOXL U4972 ( .A(n724), .B(n209), .Z(product[3]) );
  CND2X1 U4973 ( .A(n791), .B(n723), .Z(n209) );
  COR2X1 U4974 ( .A(n807), .B(n812), .Z(net20981) );
  CENX1 U4975 ( .A(n207), .B(n3912), .Z(product[5]) );
  CND2X1 U4976 ( .A(n807), .B(n812), .Z(n279) );
  CNR2IXL U4977 ( .B(n3979), .A(n3933), .Z(n2219) );
  CNR2X1 U4978 ( .A(n1723), .B(n2218), .Z(n722) );
  COR2X1 U4979 ( .A(n1707), .B(n1712), .Z(n3916) );
  CND2X1 U4980 ( .A(n1713), .B(n1716), .Z(n709) );
  CND2X1 U4981 ( .A(n2250), .B(n2219), .Z(n728) );
  CND2X1 U4982 ( .A(n1721), .B(n1722), .Z(n720) );
  CND2X1 U4983 ( .A(n1707), .B(n1712), .Z(n706) );
  COR2X1 U4984 ( .A(n1717), .B(n1720), .Z(n3917) );
  CND2X1 U4985 ( .A(n1717), .B(n1720), .Z(n714) );
  COR2X1 U4986 ( .A(n2250), .B(n2219), .Z(n3918) );
  COR2X1 U4987 ( .A(n1721), .B(n1722), .Z(n3919) );
  COR2X1 U4988 ( .A(n1740), .B(n794), .Z(n3920) );
  CND2X1 U4989 ( .A(n796), .B(n795), .Z(n229) );
  CND2X1 U4990 ( .A(n1740), .B(n794), .Z(n218) );
  CAN2XL U4991 ( .A(n793), .B(n731), .Z(product[1]) );
  CENX1 U4992 ( .A(n2781), .B(n3897), .Z(n2682) );
  CENX1 U4993 ( .A(n3965), .B(net18483), .Z(n2271) );
  CENX1 U4994 ( .A(n3964), .B(net18483), .Z(n2272) );
  CENX1 U4995 ( .A(n2792), .B(n3896), .Z(n2330) );
  CENX1 U4996 ( .A(n3974), .B(n3984), .Z(n2721) );
  CENX1 U4997 ( .A(n3959), .B(n3925), .Z(n2442) );
  CENX1 U4998 ( .A(n3972), .B(n3897), .Z(n2690) );
  CENX1 U4999 ( .A(n3959), .B(net18483), .Z(n2277) );
  CENX1 U5000 ( .A(n3962), .B(net18483), .Z(n2274) );
  CENX1 U5001 ( .A(n3961), .B(net18483), .Z(n2275) );
  CENX1 U5002 ( .A(n3958), .B(net18483), .Z(n2278) );
  CENX1 U5003 ( .A(net18979), .B(n3992), .Z(n2665) );
  CENX1 U5004 ( .A(n2809), .B(net18483), .Z(n2281) );
  CENX1 U5005 ( .A(n3956), .B(net18517), .Z(n2412) );
  CENX1 U5006 ( .A(n3966), .B(n3992), .Z(n2664) );
  CENX1 U5007 ( .A(n2798), .B(n3992), .Z(n2666) );
  CENX1 U5008 ( .A(n3960), .B(n3896), .Z(n2342) );
  CENX1 U5009 ( .A(n3956), .B(n3788), .Z(n2445) );
  CENX1 U5010 ( .A(n2781), .B(net21177), .Z(n2385) );
  CENX1 U5011 ( .A(n3977), .B(net18519), .Z(n2384) );
  CIVX1 U5012 ( .A(net18489), .Z(net18487) );
  CIVX4 U5013 ( .A(n3927), .Z(n3928) );
  CENX1 U5014 ( .A(n3971), .B(n3923), .Z(n2592) );
  CENX1 U5015 ( .A(n3972), .B(n3924), .Z(n2591) );
  CENX1 U5016 ( .A(n2782), .B(net19268), .Z(n2353) );
  CENXL U5017 ( .A(n3969), .B(net19268), .Z(n2364) );
  CENX1 U5018 ( .A(n2792), .B(net19268), .Z(n2363) );
  CENX1 U5019 ( .A(n3970), .B(net19268), .Z(n2362) );
  CENXL U5020 ( .A(net18979), .B(net19268), .Z(n2368) );
  CENX1 U5021 ( .A(n3971), .B(net19268), .Z(n2361) );
  CENX1 U5022 ( .A(n3974), .B(net19268), .Z(n2358) );
  CENX1 U5023 ( .A(n3972), .B(net19268), .Z(n2360) );
  CENX1 U5024 ( .A(n3973), .B(net19268), .Z(n2359) );
  CENX1 U5025 ( .A(n3975), .B(net19268), .Z(n2357) );
  CENX1 U5026 ( .A(n3969), .B(n3925), .Z(n2430) );
  CENX1 U5027 ( .A(n2798), .B(net19268), .Z(n2369) );
  CENX1 U5028 ( .A(n3965), .B(net19268), .Z(n2370) );
  CENX1 U5029 ( .A(n2809), .B(net19268), .Z(n2380) );
  CENX1 U5030 ( .A(n3964), .B(net19268), .Z(n2371) );
  CENX1 U5031 ( .A(n3966), .B(n3925), .Z(n2433) );
  CENX1 U5032 ( .A(n3958), .B(net19268), .Z(n2377) );
  CENX1 U5033 ( .A(net18979), .B(n3925), .Z(n2434) );
  CENX1 U5034 ( .A(n3973), .B(n3981), .Z(n2755) );
  CENX1 U5035 ( .A(n2785), .B(net19268), .Z(n2356) );
  CENX1 U5036 ( .A(n3962), .B(net19268), .Z(n2373) );
  CENX1 U5037 ( .A(n3961), .B(net19268), .Z(n2374) );
  CENX1 U5038 ( .A(n3968), .B(net19309), .Z(n2530) );
  CENX1 U5039 ( .A(n3959), .B(net19268), .Z(n2376) );
  CENX1 U5040 ( .A(n3972), .B(n3993), .Z(n2624) );
  CENX1 U5041 ( .A(n2783), .B(net19268), .Z(n2354) );
  CENX1 U5042 ( .A(n2810), .B(net19314), .Z(n2480) );
  CENX1 U5043 ( .A(n3976), .B(net19268), .Z(n2355) );
  CENX1 U5044 ( .A(n3967), .B(n3982), .Z(n2762) );
  CENX1 U5045 ( .A(n3975), .B(n3924), .Z(n2588) );
  CENX1 U5046 ( .A(n2783), .B(n3923), .Z(n2585) );
  CENX1 U5047 ( .A(n2810), .B(n3928), .Z(n2777) );
  CENX1 U5048 ( .A(n2809), .B(n3928), .Z(n2776) );
  CENX1 U5049 ( .A(n3956), .B(n3928), .Z(n2775) );
  CENX1 U5050 ( .A(n3961), .B(n3928), .Z(n2770) );
  CENX1 U5051 ( .A(n3962), .B(n3928), .Z(n2769) );
  CENX1 U5052 ( .A(n3958), .B(n3928), .Z(n2773) );
  CENX1 U5053 ( .A(n3959), .B(n3928), .Z(n2772) );
  CENX1 U5054 ( .A(n2781), .B(n3213), .Z(n2418) );
  CENX1 U5055 ( .A(n2781), .B(net19268), .Z(n2352) );
  CENX1 U5056 ( .A(n3977), .B(n3982), .Z(n2747) );
  CENX1 U5057 ( .A(n3977), .B(net19268), .Z(n2351) );
  CNR2IXL U5058 ( .B(n3979), .A(n3660), .Z(n2054) );
  COND2X1 U5059 ( .A(n2748), .B(n6), .C(n2749), .D(n3880), .Z(n2222) );
  COND2X1 U5060 ( .A(n2592), .B(n54), .C(n3145), .D(n2591), .Z(n2065) );
  CNR2IXL U5061 ( .B(n3979), .A(n3939), .Z(n2120) );
  CENX1 U5062 ( .A(n3978), .B(net18483), .Z(n2283) );
  CENX1 U5063 ( .A(n3977), .B(net18483), .Z(n2252) );
  CENX1 U5064 ( .A(n2782), .B(net18487), .Z(n2254) );
  CENX1 U5065 ( .A(n2785), .B(net18487), .Z(n2257) );
  CENX1 U5066 ( .A(n3976), .B(net18487), .Z(n2256) );
  CENX1 U5067 ( .A(n2783), .B(net18487), .Z(n2255) );
  CENX1 U5068 ( .A(n2781), .B(net18487), .Z(n2253) );
  CNR2IXL U5069 ( .B(n3979), .A(n6), .Z(product[0]) );
  CNIVX8 U5070 ( .A(n2780), .Z(n3977) );
  CND2IXL U5071 ( .B(n3979), .A(n3985), .Z(n2746) );
  COND2X2 U5072 ( .A(n2682), .B(n3931), .C(n2683), .D(n27), .Z(n2156) );
  CENXL U5073 ( .A(n3978), .B(n3923), .Z(n2613) );
  CIVX2 U5074 ( .A(n3), .Z(n3983) );
  COND2XL U5075 ( .A(n3871), .B(n3659), .C(n3941), .D(n2515), .Z(n1731) );
  CNR2X2 U5076 ( .A(n551), .B(n556), .Z(n549) );
  CEOX4 U5077 ( .A(a[0]), .B(n3980), .Z(n2827) );
  CNR2IX1 U5078 ( .B(n3979), .A(net19192), .Z(n1802) );
  CND2X1 U5079 ( .A(n2251), .B(n1739), .Z(n731) );
  CNR2XL U5080 ( .A(n2251), .B(n1739), .Z(n730) );
  CIVX2 U5081 ( .A(n3981), .Z(n3927) );
  CNR2X2 U5082 ( .A(n3741), .B(n529), .Z(n520) );
  CIVX8 U5083 ( .A(n60), .Z(n3935) );
  CENX4 U5084 ( .A(n3827), .B(n3987), .Z(n3943) );
  COND1XL U5085 ( .A(n213), .B(net19189), .C(n214), .Z(n212) );
  CIVXL U5086 ( .A(n630), .Z(n629) );
  COND2X1 U5087 ( .A(n117), .B(net21882), .C(net19281), .D(n2383), .Z(n1727)
         );
  COND1XL U5088 ( .A(n514), .B(n545), .C(n3898), .Z(n513) );
  CANR1XL U5089 ( .A(n758), .B(n517), .C(n510), .Z(n508) );
  CANR1XL U5090 ( .A(n3343), .B(n517), .C(n3146), .Z(n497) );
  CANR1XL U5091 ( .A(n489), .B(n517), .C(n490), .Z(n488) );
  COND1XL U5092 ( .A(n3852), .B(n3813), .C(n3242), .Z(n3944) );
  CNR2X1 U5093 ( .A(n1461), .B(n1482), .Z(n605) );
  CIVXL U5094 ( .A(n3944), .Z(n533) );
  CND2XL U5095 ( .A(n534), .B(n760), .Z(n525) );
  CIVXL U5096 ( .A(n534), .Z(n532) );
  CNR2X2 U5097 ( .A(n1215), .B(n1244), .Z(n3945) );
  CENX1 U5098 ( .A(n3967), .B(n3992), .Z(n2663) );
  CND2IXL U5099 ( .B(n3979), .A(n3992), .Z(n2680) );
  CENXL U5100 ( .A(n3966), .B(net18519), .Z(n2400) );
  CENXL U5101 ( .A(n3967), .B(net18519), .Z(n2399) );
  CND2IXL U5102 ( .B(n3979), .A(net18519), .Z(n2416) );
  CENX1 U5103 ( .A(n2782), .B(net21177), .Z(n2386) );
  CENX1 U5104 ( .A(n2783), .B(net21177), .Z(n2387) );
  CENX1 U5105 ( .A(n3976), .B(net21177), .Z(n2388) );
  CENX1 U5106 ( .A(n3974), .B(net21177), .Z(n2391) );
  CENX1 U5107 ( .A(n3972), .B(net18515), .Z(n2393) );
  CND2X1 U5108 ( .A(n756), .B(n494), .Z(n174) );
  COND1XL U5109 ( .A(n3851), .B(n501), .C(n494), .Z(n490) );
  CIVXL U5110 ( .A(n3945), .Z(n761) );
  COND2XL U5111 ( .A(n3880), .B(n3812), .C(n6), .D(n2779), .Z(n1739) );
  CIVXL U5112 ( .A(n512), .Z(n510) );
  CND2XL U5113 ( .A(n758), .B(n512), .Z(n176) );
  CIVXL U5114 ( .A(n3899), .Z(n517) );
  COR2XL U5115 ( .A(n1186), .B(n1159), .Z(n3948) );
  CND2XL U5116 ( .A(n3242), .B(n761), .Z(n179) );
  CENXL U5117 ( .A(n3968), .B(n4006), .Z(n2332) );
  CND2X1 U5118 ( .A(n1109), .B(n1111), .Z(n3950) );
  CENXL U5119 ( .A(n3966), .B(n4006), .Z(n2334) );
  CENXL U5120 ( .A(n2798), .B(n4006), .Z(n2336) );
  CENXL U5121 ( .A(net18979), .B(n4006), .Z(n2335) );
  CENXL U5122 ( .A(n3969), .B(n4006), .Z(n2331) );
  CENXL U5123 ( .A(n3967), .B(n4006), .Z(n2333) );
  CND2IXL U5124 ( .B(n3979), .A(n4006), .Z(n2350) );
  CANR1XL U5125 ( .A(n760), .B(n3944), .C(n528), .Z(n526) );
  CANR1X2 U5126 ( .A(n631), .B(n650), .C(n632), .Z(n630) );
  CENXL U5127 ( .A(n3979), .B(net19302), .Z(n2580) );
  CANR1X2 U5128 ( .A(n608), .B(n769), .C(n601), .Z(n595) );
  CANR1X2 U5129 ( .A(n562), .B(n549), .C(n550), .Z(n548) );
  CENX4 U5130 ( .A(a[10]), .B(n3498), .Z(n3955) );
  CENX4 U5131 ( .A(a[18]), .B(n3659), .Z(net19062) );
  COND2XL U5132 ( .A(n54), .B(n3780), .C(n3145), .D(n2614), .Z(n1734) );
  COND2XL U5133 ( .A(n18), .B(n3986), .C(n3933), .D(n2746), .Z(n1738) );
  COND2XL U5134 ( .A(n3904), .B(n3549), .C(n33), .D(n2680), .Z(n1736) );
  COND1XL U5135 ( .A(n594), .B(n3102), .C(n3872), .Z(n593) );
  CIVXL U5136 ( .A(n504), .Z(n757) );
  CIVXL U5137 ( .A(n3461), .Z(n501) );
  CIVXL U5138 ( .A(n714), .Z(n712) );
  CANR1X2 U5139 ( .A(n576), .B(n3882), .C(n577), .Z(n575) );
  CIVX8 U5140 ( .A(net18489), .Z(net18483) );
  CND2X4 U5141 ( .A(n2826), .B(n3932), .Z(n18) );
  CND2X4 U5142 ( .A(n3929), .B(n2825), .Z(n27) );
  CENX4 U5143 ( .A(a[12]), .B(n3437), .Z(n60) );
  CIVX2 U5144 ( .A(n890), .Z(n891) );
  CIVX2 U5145 ( .A(n864), .Z(n865) );
  CIVX2 U5146 ( .A(n842), .Z(n843) );
  CIVX2 U5147 ( .A(n794), .Z(n795) );
  CIVX2 U5148 ( .A(n730), .Z(n793) );
  CIVX2 U5149 ( .A(n722), .Z(n791) );
  CIVX2 U5150 ( .A(n708), .Z(n788) );
  CIVX2 U5151 ( .A(n700), .Z(n786) );
  CIVX2 U5152 ( .A(n696), .Z(n785) );
  CIVX2 U5153 ( .A(n693), .Z(n784) );
  CIVX2 U5154 ( .A(n674), .Z(n781) );
  CIVX2 U5155 ( .A(n324), .Z(n741) );
  CIVX2 U5156 ( .A(n731), .Z(n729) );
  CIVX2 U5157 ( .A(n728), .Z(n726) );
  CIVX2 U5158 ( .A(n720), .Z(n718) );
  CIVX2 U5159 ( .A(n706), .Z(n704) );
  CIVX2 U5160 ( .A(n699), .Z(n698) );
  CIVX2 U5161 ( .A(n688), .Z(n686) );
  CIVX2 U5162 ( .A(n683), .Z(n681) );
  CIVX2 U5163 ( .A(n665), .Z(n779) );
  CIVX2 U5164 ( .A(n606), .Z(n608) );
  CIVX2 U5165 ( .A(n605), .Z(n770) );
  CIVX2 U5166 ( .A(n594), .Z(n596) );
  CIVX2 U5167 ( .A(n468), .Z(n753) );
  CIVX2 U5168 ( .A(n448), .Z(n751) );
  CIVX2 U5169 ( .A(n434), .Z(n432) );
  CIVX2 U5170 ( .A(n409), .Z(n748) );
  CIVX2 U5171 ( .A(n351), .Z(n349) );
  CIVX2 U5172 ( .A(n342), .Z(n340) );
  CIVX2 U5173 ( .A(n333), .Z(n331) );
  CIVX2 U5174 ( .A(n229), .Z(n227) );
  CIVX2 U5175 ( .A(n218), .Z(n216) );
  CIVX2 U5176 ( .A(n1130), .Z(n1131) );
endmodule


module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push0, cmd0_en_0, cmd1_en_0, cmd0_en_1, cmd1_en_1, push0_0,
         cmd0_en_2_d, cmd1_en_2_d, push0_2, push0_1, cmd2_en_1, cmd2_en_2,
         cmd0_en_2, cmd1_en_2, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, roundit, _pushout_d,
         N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428,
         N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439,
         N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450,
         N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461,
         N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472,
         N473, N474, N475, N476, N477, N478, N479, N480, N481, n12, n215, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467;
  wire   [1:0] cmd0;
  wire   [1:0] cmd0_0;
  wire   [1:0] cmd0_2;
  wire   [1:0] cmd0_1;
  wire   [63:0] out0_0;
  wire   [63:0] out0_2;
  wire   [63:0] out0_1;
  wire   [31:0] q0;
  wire   [31:0] h0;
  wire   [63:0] acc_cmd1;
  wire   [63:0] acc;
  wire   [63:0] out1_2;
  wire   [63:0] out1_0;
  wire   [63:0] out1_1;
  wire   [63:0] out2_2;
  wire   [6:0] h0_1;
  wire   [6:0] h0_0;

  CFD2QX2 cmd0_en_2_d_reg ( .D(n1389), .CP(clk), .CD(n1442), .Q(cmd0_en_2_d)
         );
  CFD2QX2 \q0_reg[30]  ( .D(n688), .CP(clk), .CD(n1450), .Q(q0[30]) );
  CFD2QX2 \q0_reg[28]  ( .D(n686), .CP(clk), .CD(n1450), .Q(q0[28]) );
  CFD2QX2 \q0_reg[24]  ( .D(n682), .CP(clk), .CD(n1450), .Q(q0[24]) );
  CFD2QX2 \q0_reg[22]  ( .D(n680), .CP(clk), .CD(n1450), .Q(q0[22]) );
  CFD2QX2 \q0_reg[16]  ( .D(n1184), .CP(clk), .CD(n1451), .Q(q0[16]) );
  CFD2QX2 \q0_reg[10]  ( .D(n668), .CP(clk), .CD(n1451), .Q(q0[10]) );
  CFD2QX2 \q0_reg[8]  ( .D(n1183), .CP(clk), .CD(n1451), .Q(q0[8]) );
  CFD2QX2 \q0_reg[2]  ( .D(n1180), .CP(clk), .CD(n1452), .Q(q0[2]) );
  CFD2QX2 \q0_reg[0]  ( .D(n658), .CP(clk), .CD(n1452), .Q(q0[0]) );
  CFD2QX2 \h0_reg[15]  ( .D(n1175), .CP(clk), .CD(n1453), .Q(h0[15]) );
  sfilt_DW01_add_2 add_117 ( .A(out1_1), .B(acc_cmd1), .CI(1'b0), .SUM({N272, 
        N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209}) );
  sfilt_DW01_add_3 add_183 ( .A(out2_2), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, roundit}), 
        .CI(1'b0), .SUM({N481, N480, N479, N478, N477, N476, N475, N474, N473, 
        N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, 
        N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, 
        N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, 
        N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, 
        N424, N423, N422, N421, N420, N419, N418}) );
  sfilt_DW_mult_tc_1 r304 ( .a(q0), .b(h0), .product({N78, N77, N76, N75, N74, 
        N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, 
        N17, N16, N15}) );
  CFD2QX1 \q0_reg[1]  ( .D(n659), .CP(clk), .CD(n1437), .Q(q0[1]) );
  CFD2QX1 \q0_reg[27]  ( .D(n685), .CP(clk), .CD(n1437), .Q(q0[27]) );
  CFD2QX1 \q0_reg[15]  ( .D(n673), .CP(clk), .CD(n1451), .Q(q0[15]) );
  CFD2QX1 \q0_reg[13]  ( .D(n671), .CP(clk), .CD(n1451), .Q(q0[13]) );
  CFD2QX1 \q0_reg[29]  ( .D(n687), .CP(clk), .CD(n1437), .Q(q0[29]) );
  CFD2QX1 \q0_reg[7]  ( .D(n665), .CP(clk), .CD(n1451), .Q(q0[7]) );
  CFD2QX1 \q0_reg[23]  ( .D(n681), .CP(clk), .CD(n1437), .Q(q0[23]) );
  CFD2QX1 \q0_reg[25]  ( .D(n683), .CP(clk), .CD(n1450), .Q(q0[25]) );
  CFD2QXL \out0_0_reg[42]  ( .D(N57), .CP(clk), .CD(n1472), .Q(out0_0[42]) );
  CFD2QXL \out1_0_reg[42]  ( .D(N57), .CP(clk), .CD(n1459), .Q(out1_0[42]) );
  CFD2QXL \out0_0_reg[43]  ( .D(N58), .CP(clk), .CD(n1472), .Q(out0_0[43]) );
  CFD2QXL \out1_0_reg[43]  ( .D(N58), .CP(clk), .CD(n1459), .Q(out1_0[43]) );
  CFD2QXL \out0_0_reg[44]  ( .D(N59), .CP(clk), .CD(n1449), .Q(out0_0[44]) );
  CFD2QXL \out1_0_reg[44]  ( .D(N59), .CP(clk), .CD(n1459), .Q(out1_0[44]) );
  CFD2QXL \out0_0_reg[45]  ( .D(N60), .CP(clk), .CD(n1448), .Q(out0_0[45]) );
  CFD2QXL \out1_0_reg[45]  ( .D(N60), .CP(clk), .CD(n1459), .Q(out1_0[45]) );
  CFD2QXL \out0_0_reg[46]  ( .D(N61), .CP(clk), .CD(n1448), .Q(out0_0[46]) );
  CFD2QXL \out1_0_reg[46]  ( .D(N61), .CP(clk), .CD(n1459), .Q(out1_0[46]) );
  CFD2QXL \out0_0_reg[47]  ( .D(N62), .CP(clk), .CD(n1448), .Q(out0_0[47]) );
  CFD2QXL \out1_0_reg[47]  ( .D(N62), .CP(clk), .CD(n1458), .Q(out1_0[47]) );
  CFD2QXL \out0_0_reg[48]  ( .D(N63), .CP(clk), .CD(n1447), .Q(out0_0[48]) );
  CFD2QXL \out1_0_reg[48]  ( .D(N63), .CP(clk), .CD(n1458), .Q(out1_0[48]) );
  CFD2QXL \out0_0_reg[49]  ( .D(N64), .CP(clk), .CD(n1447), .Q(out0_0[49]) );
  CFD2QXL \out1_0_reg[49]  ( .D(N64), .CP(clk), .CD(n1458), .Q(out1_0[49]) );
  CFD2QXL \out0_0_reg[50]  ( .D(N65), .CP(clk), .CD(n1447), .Q(out0_0[50]) );
  CFD2QXL \out1_0_reg[50]  ( .D(N65), .CP(clk), .CD(n1458), .Q(out1_0[50]) );
  CFD2QXL \out0_0_reg[51]  ( .D(N66), .CP(clk), .CD(n1446), .Q(out0_0[51]) );
  CFD2QXL \out1_0_reg[51]  ( .D(N66), .CP(clk), .CD(n1458), .Q(out1_0[51]) );
  CFD2QXL \out0_0_reg[52]  ( .D(N67), .CP(clk), .CD(n1446), .Q(out0_0[52]) );
  CFD2QXL \out1_0_reg[52]  ( .D(N67), .CP(clk), .CD(n1458), .Q(out1_0[52]) );
  CFD2QXL \out0_0_reg[53]  ( .D(N68), .CP(clk), .CD(n1445), .Q(out0_0[53]) );
  CFD2QXL \out1_0_reg[53]  ( .D(N68), .CP(clk), .CD(n1458), .Q(out1_0[53]) );
  CFD2QXL \out0_0_reg[54]  ( .D(N69), .CP(clk), .CD(n1445), .Q(out0_0[54]) );
  CFD2QXL \out1_0_reg[54]  ( .D(N69), .CP(clk), .CD(n1457), .Q(out1_0[54]) );
  CFD2QXL \out0_0_reg[55]  ( .D(N70), .CP(clk), .CD(n1445), .Q(out0_0[55]) );
  CFD2QXL \out1_0_reg[55]  ( .D(N70), .CP(clk), .CD(n1457), .Q(out1_0[55]) );
  CFD2QXL \out0_0_reg[56]  ( .D(N71), .CP(clk), .CD(n1444), .Q(out0_0[56]) );
  CFD2QXL \out1_0_reg[56]  ( .D(N71), .CP(clk), .CD(n1457), .Q(out1_0[56]) );
  CFD2QXL \out0_0_reg[57]  ( .D(N72), .CP(clk), .CD(n1444), .Q(out0_0[57]) );
  CFD2QXL \out1_0_reg[57]  ( .D(N72), .CP(clk), .CD(n1457), .Q(out1_0[57]) );
  CFD2QXL \out0_0_reg[58]  ( .D(N73), .CP(clk), .CD(n1443), .Q(out0_0[58]) );
  CFD2QXL \out1_0_reg[58]  ( .D(N73), .CP(clk), .CD(n1457), .Q(out1_0[58]) );
  CFD2QXL \out0_0_reg[59]  ( .D(N74), .CP(clk), .CD(n1443), .Q(out0_0[59]) );
  CFD2QXL \out1_0_reg[59]  ( .D(N74), .CP(clk), .CD(n1457), .Q(out1_0[59]) );
  CFD2QXL \out0_0_reg[60]  ( .D(N75), .CP(clk), .CD(n1443), .Q(out0_0[60]) );
  CFD2QXL \out1_0_reg[60]  ( .D(N75), .CP(clk), .CD(n1456), .Q(out1_0[60]) );
  CFD2QXL \out0_0_reg[61]  ( .D(N76), .CP(clk), .CD(n1442), .Q(out0_0[61]) );
  CFD2QXL \out1_0_reg[61]  ( .D(N76), .CP(clk), .CD(n1456), .Q(out1_0[61]) );
  CFD2QXL \out0_0_reg[62]  ( .D(N77), .CP(clk), .CD(n1442), .Q(out0_0[62]) );
  CFD2QXL \out1_0_reg[62]  ( .D(N77), .CP(clk), .CD(n1456), .Q(out1_0[62]) );
  CFD2QX1 \q0_reg[21]  ( .D(n679), .CP(clk), .CD(n1437), .Q(q0[21]) );
  CFD2QXL \out1_0_reg[41]  ( .D(N56), .CP(clk), .CD(n1459), .Q(out1_0[41]) );
  CFD2QXL \out1_1_reg[41]  ( .D(n1157), .CP(clk), .CD(n1459), .Q(out1_1[41])
         );
  CFD2QXL \out0_1_reg[63]  ( .D(n1155), .CP(clk), .CD(n1456), .Q(out0_1[63])
         );
  CFD2QXL \out0_1_reg[62]  ( .D(n1153), .CP(clk), .CD(n1442), .Q(out0_1[62])
         );
  CFD2QXL \out0_1_reg[61]  ( .D(n1151), .CP(clk), .CD(n1442), .Q(out0_1[61])
         );
  CFD2QXL \out0_1_reg[60]  ( .D(n1149), .CP(clk), .CD(n1443), .Q(out0_1[60])
         );
  CFD2QXL \out0_1_reg[59]  ( .D(n1147), .CP(clk), .CD(n1443), .Q(out0_1[59])
         );
  CFD2QXL \out0_1_reg[58]  ( .D(n1145), .CP(clk), .CD(n1444), .Q(out0_1[58])
         );
  CFD2QXL \out0_1_reg[57]  ( .D(n1143), .CP(clk), .CD(n1444), .Q(out0_1[57])
         );
  CFD2QXL \out0_1_reg[56]  ( .D(n1141), .CP(clk), .CD(n1444), .Q(out0_1[56])
         );
  CFD2QXL \out0_1_reg[55]  ( .D(n1139), .CP(clk), .CD(n1445), .Q(out0_1[55])
         );
  CFD2QXL \out0_1_reg[54]  ( .D(n1137), .CP(clk), .CD(n1445), .Q(out0_1[54])
         );
  CFD2QXL \out0_1_reg[53]  ( .D(n1135), .CP(clk), .CD(n1445), .Q(out0_1[53])
         );
  CFD2QXL \out0_1_reg[52]  ( .D(n1133), .CP(clk), .CD(n1446), .Q(out0_1[52])
         );
  CFD2QXL \out0_1_reg[51]  ( .D(n1131), .CP(clk), .CD(n1446), .Q(out0_1[51])
         );
  CFD2QXL \out0_1_reg[50]  ( .D(n1129), .CP(clk), .CD(n1447), .Q(out0_1[50])
         );
  CFD2QXL \out0_1_reg[49]  ( .D(n1127), .CP(clk), .CD(n1447), .Q(out0_1[49])
         );
  CFD2QXL \out0_1_reg[48]  ( .D(n1125), .CP(clk), .CD(n1447), .Q(out0_1[48])
         );
  CFD2QXL \out0_1_reg[47]  ( .D(n1123), .CP(clk), .CD(n1448), .Q(out0_1[47])
         );
  CFD2QXL \out0_1_reg[46]  ( .D(n1121), .CP(clk), .CD(n1448), .Q(out0_1[46])
         );
  CFD2QXL \out0_1_reg[45]  ( .D(n1119), .CP(clk), .CD(n1449), .Q(out0_1[45])
         );
  CFD2QXL \out0_1_reg[44]  ( .D(n1117), .CP(clk), .CD(n1449), .Q(out0_1[44])
         );
  CFD2QXL \out0_1_reg[43]  ( .D(n1115), .CP(clk), .CD(n1472), .Q(out0_1[43])
         );
  CFD2QXL \out0_1_reg[42]  ( .D(n1113), .CP(clk), .CD(n1472), .Q(out0_1[42])
         );
  CFD2QXL \out0_1_reg[41]  ( .D(n1111), .CP(clk), .CD(n1472), .Q(out0_1[41])
         );
  CFD2QXL \out0_1_reg[40]  ( .D(n1109), .CP(clk), .CD(n1473), .Q(out0_1[40])
         );
  CFD2QXL \out0_1_reg[39]  ( .D(n1107), .CP(clk), .CD(n1473), .Q(out0_1[39])
         );
  CFD2QXL \out0_1_reg[38]  ( .D(n1105), .CP(clk), .CD(n1474), .Q(out0_1[38])
         );
  CFD2QXL \out0_1_reg[37]  ( .D(n1103), .CP(clk), .CD(n1474), .Q(out0_1[37])
         );
  CFD2QXL \out0_1_reg[36]  ( .D(n1101), .CP(clk), .CD(n1474), .Q(out0_1[36])
         );
  CFD2QXL \out0_1_reg[35]  ( .D(n1099), .CP(clk), .CD(n1475), .Q(out0_1[35])
         );
  CFD2QXL \out0_1_reg[34]  ( .D(n1097), .CP(clk), .CD(n1475), .Q(out0_1[34])
         );
  CFD2QXL \out0_1_reg[33]  ( .D(n1095), .CP(clk), .CD(n1476), .Q(out0_1[33])
         );
  CFD2QXL \out0_1_reg[32]  ( .D(n1093), .CP(clk), .CD(n1476), .Q(out0_1[32])
         );
  CFD2QXL \out0_1_reg[31]  ( .D(n1091), .CP(clk), .CD(n1476), .Q(out0_1[31])
         );
  CFD2QXL \out0_1_reg[30]  ( .D(n1089), .CP(clk), .CD(n1477), .Q(out0_1[30])
         );
  CFD2QXL \out0_1_reg[29]  ( .D(n1087), .CP(clk), .CD(n1477), .Q(out0_1[29])
         );
  CFD2QXL \out0_1_reg[28]  ( .D(n1085), .CP(clk), .CD(n1477), .Q(out0_1[28])
         );
  CFD2QXL \out0_1_reg[27]  ( .D(n1083), .CP(clk), .CD(n1478), .Q(out0_1[27])
         );
  CFD2QXL \out0_1_reg[26]  ( .D(n1081), .CP(clk), .CD(n1478), .Q(out0_1[26])
         );
  CFD2QXL \out0_1_reg[25]  ( .D(n1079), .CP(clk), .CD(n1479), .Q(out0_1[25])
         );
  CFD2QXL \out0_1_reg[24]  ( .D(n1077), .CP(clk), .CD(n1479), .Q(out0_1[24])
         );
  CFD2QXL \out0_1_reg[23]  ( .D(n1075), .CP(clk), .CD(n1480), .Q(out0_1[23])
         );
  CFD2QXL \out0_1_reg[22]  ( .D(n1073), .CP(clk), .CD(n1480), .Q(out0_1[22])
         );
  CFD2QXL \out0_1_reg[21]  ( .D(n1071), .CP(clk), .CD(n1480), .Q(out0_1[21])
         );
  CFD2QXL \out0_1_reg[20]  ( .D(n1069), .CP(clk), .CD(n1481), .Q(out0_1[20])
         );
  CFD2QXL \out0_1_reg[19]  ( .D(n1067), .CP(clk), .CD(n1481), .Q(out0_1[19])
         );
  CFD2QXL \out0_1_reg[18]  ( .D(n1065), .CP(clk), .CD(n1481), .Q(out0_1[18])
         );
  CFD2QXL \out0_1_reg[17]  ( .D(n1063), .CP(clk), .CD(n1482), .Q(out0_1[17])
         );
  CFD2QXL \out0_1_reg[16]  ( .D(n1061), .CP(clk), .CD(n1482), .Q(out0_1[16])
         );
  CFD2QXL \out0_1_reg[15]  ( .D(n1059), .CP(clk), .CD(n1481), .Q(out0_1[15])
         );
  CFD2QXL \out0_1_reg[14]  ( .D(n1057), .CP(clk), .CD(n1483), .Q(out0_1[14])
         );
  CFD2QXL \out0_1_reg[13]  ( .D(n1055), .CP(clk), .CD(n1483), .Q(out0_1[13])
         );
  CFD2QXL \out0_1_reg[12]  ( .D(n1053), .CP(clk), .CD(n1483), .Q(out0_1[12])
         );
  CFD2QXL \out0_1_reg[11]  ( .D(n1051), .CP(clk), .CD(n1461), .Q(out0_1[11])
         );
  CFD2QXL \out0_1_reg[10]  ( .D(n1049), .CP(clk), .CD(n1462), .Q(out0_1[10])
         );
  CFD2QXL \out0_1_reg[9]  ( .D(n1047), .CP(clk), .CD(n1462), .Q(out0_1[9]) );
  CFD2QXL \out0_1_reg[8]  ( .D(n1045), .CP(clk), .CD(n1463), .Q(out0_1[8]) );
  CFD2QXL \out0_1_reg[7]  ( .D(n1043), .CP(clk), .CD(n1463), .Q(out0_1[7]) );
  CFD2QXL \out0_1_reg[6]  ( .D(n1041), .CP(clk), .CD(n1463), .Q(out0_1[6]) );
  CFD2QXL \out0_1_reg[5]  ( .D(n1039), .CP(clk), .CD(n1464), .Q(out0_1[5]) );
  CFD2QXL \out0_1_reg[4]  ( .D(n1037), .CP(clk), .CD(n1464), .Q(out0_1[4]) );
  CFD2QXL \out0_1_reg[3]  ( .D(n1035), .CP(clk), .CD(n1465), .Q(out0_1[3]) );
  CFD2QXL \out0_1_reg[2]  ( .D(n1033), .CP(clk), .CD(n1465), .Q(out0_1[2]) );
  CFD2QXL \out0_1_reg[1]  ( .D(n1031), .CP(clk), .CD(n1465), .Q(out0_1[1]) );
  CFD2QXL \out0_1_reg[0]  ( .D(n1029), .CP(clk), .CD(n1455), .Q(out0_1[0]) );
  CFD2QXL cmd1_en_1_reg ( .D(cmd1_en_0), .CP(clk), .CD(n1442), .Q(cmd1_en_1)
         );
  CFD2QXL cmd0_en_1_reg ( .D(cmd0_en_0), .CP(clk), .CD(n1437), .Q(cmd0_en_1)
         );
  CFD2QXL \h0_0_reg[6]  ( .D(n631), .CP(clk), .CD(n1455), .Q(h0_0[6]) );
  CFD2QXL \h0_0_reg[5]  ( .D(n628), .CP(clk), .CD(n1455), .Q(h0_0[5]) );
  CFD2QXL \h0_0_reg[4]  ( .D(n625), .CP(clk), .CD(n1455), .Q(h0_0[4]) );
  CFD2QXL \h0_0_reg[3]  ( .D(n622), .CP(clk), .CD(n1466), .Q(h0_0[3]) );
  CFD2QXL \h0_0_reg[2]  ( .D(n619), .CP(clk), .CD(n1456), .Q(h0_0[2]) );
  CFD2QXL \h0_0_reg[1]  ( .D(n616), .CP(clk), .CD(n1455), .Q(h0_0[1]) );
  CFD2QXL \h0_0_reg[0]  ( .D(n613), .CP(clk), .CD(n1455), .Q(h0_0[0]) );
  CFD2QXL \dout_reg[31]  ( .D(n789), .CP(clk), .CD(n1471), .Q(z[31]) );
  CFD2QXL \dout_reg[30]  ( .D(n788), .CP(clk), .CD(n1471), .Q(z[30]) );
  CFD2QXL \dout_reg[29]  ( .D(n1028), .CP(clk), .CD(n1471), .Q(z[29]) );
  CFD2QXL \dout_reg[28]  ( .D(n1027), .CP(clk), .CD(n1471), .Q(z[28]) );
  CFD2QXL \dout_reg[27]  ( .D(n1026), .CP(clk), .CD(n1471), .Q(z[27]) );
  CFD2QXL \dout_reg[26]  ( .D(n1025), .CP(clk), .CD(n1471), .Q(z[26]) );
  CFD2QXL \dout_reg[25]  ( .D(n1024), .CP(clk), .CD(n1471), .Q(z[25]) );
  CFD2QXL \dout_reg[24]  ( .D(n1023), .CP(clk), .CD(n1471), .Q(z[24]) );
  CFD2QXL \dout_reg[23]  ( .D(n781), .CP(clk), .CD(n1471), .Q(z[23]) );
  CFD2QXL \dout_reg[22]  ( .D(n780), .CP(clk), .CD(n1471), .Q(z[22]) );
  CFD2QXL \dout_reg[21]  ( .D(n1022), .CP(clk), .CD(n1471), .Q(z[21]) );
  CFD2QXL \dout_reg[20]  ( .D(n778), .CP(clk), .CD(n1471), .Q(z[20]) );
  CFD2QXL \dout_reg[19]  ( .D(n1021), .CP(clk), .CD(n1470), .Q(z[19]) );
  CFD2QXL \dout_reg[18]  ( .D(n1020), .CP(clk), .CD(n1470), .Q(z[18]) );
  CFD2QXL \dout_reg[17]  ( .D(n1019), .CP(clk), .CD(n1470), .Q(z[17]) );
  CFD2QXL \dout_reg[16]  ( .D(n1018), .CP(clk), .CD(n1470), .Q(z[16]) );
  CFD2QXL \dout_reg[15]  ( .D(n1017), .CP(clk), .CD(n1470), .Q(z[15]) );
  CFD2QXL \dout_reg[14]  ( .D(n1016), .CP(clk), .CD(n1470), .Q(z[14]) );
  CFD2QXL \dout_reg[13]  ( .D(n1015), .CP(clk), .CD(n1470), .Q(z[13]) );
  CFD2QXL \dout_reg[12]  ( .D(n1014), .CP(clk), .CD(n1470), .Q(z[12]) );
  CFD2QXL \dout_reg[11]  ( .D(n1013), .CP(clk), .CD(n1470), .Q(z[11]) );
  CFD2QXL \dout_reg[10]  ( .D(n1012), .CP(clk), .CD(n1470), .Q(z[10]) );
  CFD2QXL \dout_reg[9]  ( .D(n1011), .CP(clk), .CD(n1470), .Q(z[9]) );
  CFD2QXL \dout_reg[8]  ( .D(n1010), .CP(clk), .CD(n1470), .Q(z[8]) );
  CFD2QXL \dout_reg[7]  ( .D(n1009), .CP(clk), .CD(n1470), .Q(z[7]) );
  CFD2QXL \dout_reg[6]  ( .D(n1008), .CP(clk), .CD(n1469), .Q(z[6]) );
  CFD2QXL \dout_reg[5]  ( .D(n1007), .CP(clk), .CD(n1469), .Q(z[5]) );
  CFD2QXL \dout_reg[4]  ( .D(n1006), .CP(clk), .CD(n1469), .Q(z[4]) );
  CFD2QXL \dout_reg[3]  ( .D(n1005), .CP(clk), .CD(n1469), .Q(z[3]) );
  CFD2QXL \dout_reg[2]  ( .D(n1004), .CP(clk), .CD(n1469), .Q(z[2]) );
  CFD2QXL \dout_reg[1]  ( .D(n1003), .CP(clk), .CD(n1469), .Q(z[1]) );
  CFD2QXL \dout_reg[0]  ( .D(n1002), .CP(clk), .CD(n1469), .Q(z[0]) );
  CFD2QXL \out2_2_reg[62]  ( .D(n1001), .CP(clk), .CD(n1466), .Q(out2_2[62])
         );
  CFD2QXL \out1_1_reg[63]  ( .D(n999), .CP(clk), .CD(n1456), .Q(out1_1[63]) );
  CFD2QXL push0_reg ( .D(n1501), .CP(clk), .CD(n1449), .Q(push0) );
  CFD2QXL \out2_2_reg[63]  ( .D(n547), .CP(clk), .CD(n1466), .Q(out2_2[63]) );
  CFD2QXL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n1450), .Q(cmd0[0]) );
  CFD2QXL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n1450), .Q(cmd0[1]) );
  CFD2QXL cmd2_en_1_reg ( .D(n2465), .CP(clk), .CD(n1455), .Q(cmd2_en_1) );
  CFD2QXL \h0_1_reg[6]  ( .D(n630), .CP(clk), .CD(n1455), .Q(h0_1[6]) );
  CFD2QXL \h0_1_reg[5]  ( .D(n627), .CP(clk), .CD(n1455), .Q(h0_1[5]) );
  CFD2QXL \acc_reg[63]  ( .D(n546), .CP(clk), .CD(n1466), .Q(acc[63]) );
  CFD2QXL \acc_reg[52]  ( .D(n440), .CP(clk), .CD(n1446), .Q(acc[52]) );
  CFD2QXL \acc_reg[54]  ( .D(n436), .CP(clk), .CD(n1445), .Q(acc[54]) );
  CFD2QXL \acc_reg[58]  ( .D(n428), .CP(clk), .CD(n1444), .Q(acc[58]) );
  CFD2QXL \acc_reg[60]  ( .D(n424), .CP(clk), .CD(n1443), .Q(acc[60]) );
  CFD2QXL \acc_reg[61]  ( .D(n422), .CP(clk), .CD(n1443), .Q(acc[61]) );
  CFD2QXL \acc_reg[62]  ( .D(n420), .CP(clk), .CD(n1442), .Q(acc[62]) );
  CFD2QXL \acc_reg[32]  ( .D(n480), .CP(clk), .CD(n1476), .Q(acc[32]) );
  CFD2QXL \acc_reg[43]  ( .D(n458), .CP(clk), .CD(n1472), .Q(acc[43]) );
  CFD2QXL \acc_reg[41]  ( .D(n462), .CP(clk), .CD(n1473), .Q(acc[41]) );
  CFD2QXL \acc_reg[35]  ( .D(n474), .CP(clk), .CD(n1475), .Q(acc[35]) );
  CFD2QXL \acc_reg[33]  ( .D(n478), .CP(clk), .CD(n1476), .Q(acc[33]) );
  CFD2QXL \acc_reg[59]  ( .D(n426), .CP(clk), .CD(n1443), .Q(acc[59]) );
  CFD2QXL \acc_reg[55]  ( .D(n434), .CP(clk), .CD(n1445), .Q(acc[55]) );
  CFD2QXL \acc_reg[56]  ( .D(n432), .CP(clk), .CD(n1445), .Q(acc[56]) );
  CFD2QXL \acc_reg[57]  ( .D(n430), .CP(clk), .CD(n1444), .Q(acc[57]) );
  CFD2QXL \acc_reg[37]  ( .D(n470), .CP(clk), .CD(n1474), .Q(acc[37]) );
  CFD2QXL \acc_reg[51]  ( .D(n442), .CP(clk), .CD(n1446), .Q(acc[51]) );
  CFD2QXL \acc_reg[50]  ( .D(n444), .CP(clk), .CD(n1447), .Q(acc[50]) );
  CFD2QXL \acc_reg[53]  ( .D(n438), .CP(clk), .CD(n1446), .Q(acc[53]) );
  CFD2QXL \acc_reg[44]  ( .D(n456), .CP(clk), .CD(n1472), .Q(acc[44]) );
  CFD2QXL \acc_reg[42]  ( .D(n460), .CP(clk), .CD(n1472), .Q(acc[42]) );
  CFD2QXL \acc_reg[49]  ( .D(n446), .CP(clk), .CD(n1447), .Q(acc[49]) );
  CFD2QXL \acc_reg[39]  ( .D(n466), .CP(clk), .CD(n1473), .Q(acc[39]) );
  CFD2QXL \acc_reg[47]  ( .D(n450), .CP(clk), .CD(n1448), .Q(acc[47]) );
  CFD2QXL \acc_reg[45]  ( .D(n454), .CP(clk), .CD(n1449), .Q(acc[45]) );
  CFD2QXL \acc_reg[38]  ( .D(n468), .CP(clk), .CD(n1474), .Q(acc[38]) );
  CFD2QXL \acc_reg[48]  ( .D(n448), .CP(clk), .CD(n1448), .Q(acc[48]) );
  CFD2QXL \acc_reg[40]  ( .D(n464), .CP(clk), .CD(n1473), .Q(acc[40]) );
  CFD2QXL \acc_reg[36]  ( .D(n472), .CP(clk), .CD(n1475), .Q(acc[36]) );
  CFD2QXL \acc_reg[34]  ( .D(n476), .CP(clk), .CD(n1475), .Q(acc[34]) );
  CFD2QXL \acc_reg[46]  ( .D(n452), .CP(clk), .CD(n1448), .Q(acc[46]) );
  CFD2QXL \h0_1_reg[4]  ( .D(n624), .CP(clk), .CD(n1455), .Q(h0_1[4]) );
  CFD2QXL \out1_1_reg[62]  ( .D(n996), .CP(clk), .CD(n1456), .Q(out1_1[62]) );
  CFD2QXL \out1_1_reg[61]  ( .D(n994), .CP(clk), .CD(n1456), .Q(out1_1[61]) );
  CFD2QXL \out1_1_reg[60]  ( .D(n992), .CP(clk), .CD(n1457), .Q(out1_1[60]) );
  CFD2QXL \out1_1_reg[59]  ( .D(n990), .CP(clk), .CD(n1457), .Q(out1_1[59]) );
  CFD2QXL \out1_1_reg[58]  ( .D(n988), .CP(clk), .CD(n1457), .Q(out1_1[58]) );
  CFD2QXL \out1_1_reg[57]  ( .D(n986), .CP(clk), .CD(n1457), .Q(out1_1[57]) );
  CFD2QXL \out1_1_reg[56]  ( .D(n984), .CP(clk), .CD(n1457), .Q(out1_1[56]) );
  CFD2QXL \out1_1_reg[55]  ( .D(n982), .CP(clk), .CD(n1457), .Q(out1_1[55]) );
  CFD2QXL \out1_1_reg[54]  ( .D(n980), .CP(clk), .CD(n1457), .Q(out1_1[54]) );
  CFD2QXL \out1_1_reg[53]  ( .D(n978), .CP(clk), .CD(n1458), .Q(out1_1[53]) );
  CFD2QXL \out1_1_reg[52]  ( .D(n976), .CP(clk), .CD(n1458), .Q(out1_1[52]) );
  CFD2QXL \out1_1_reg[51]  ( .D(n974), .CP(clk), .CD(n1458), .Q(out1_1[51]) );
  CFD2QXL \out1_1_reg[50]  ( .D(n972), .CP(clk), .CD(n1458), .Q(out1_1[50]) );
  CFD2QXL \out1_1_reg[49]  ( .D(n970), .CP(clk), .CD(n1458), .Q(out1_1[49]) );
  CFD2QXL \out1_1_reg[48]  ( .D(n968), .CP(clk), .CD(n1458), .Q(out1_1[48]) );
  CFD2QXL \out1_1_reg[47]  ( .D(n966), .CP(clk), .CD(n1459), .Q(out1_1[47]) );
  CFD2QXL \out1_1_reg[46]  ( .D(n964), .CP(clk), .CD(n1459), .Q(out1_1[46]) );
  CFD2QXL \out1_1_reg[45]  ( .D(n962), .CP(clk), .CD(n1459), .Q(out1_1[45]) );
  CFD2QXL \out1_1_reg[44]  ( .D(n960), .CP(clk), .CD(n1459), .Q(out1_1[44]) );
  CFD2QXL \out1_1_reg[43]  ( .D(n958), .CP(clk), .CD(n1459), .Q(out1_1[43]) );
  CFD2QXL \out1_1_reg[42]  ( .D(n956), .CP(clk), .CD(n1459), .Q(out1_1[42]) );
  CFD2QXL \out1_1_reg[40]  ( .D(n954), .CP(clk), .CD(n1460), .Q(out1_1[40]) );
  CFD2QXL \out1_1_reg[39]  ( .D(n952), .CP(clk), .CD(n1460), .Q(out1_1[39]) );
  CFD2QXL \out1_1_reg[38]  ( .D(n950), .CP(clk), .CD(n1460), .Q(out1_1[38]) );
  CFD2QXL \out1_1_reg[37]  ( .D(n948), .CP(clk), .CD(n1460), .Q(out1_1[37]) );
  CFD2QXL \out1_1_reg[36]  ( .D(n946), .CP(clk), .CD(n1460), .Q(out1_1[36]) );
  CFD2QXL \out1_1_reg[35]  ( .D(n944), .CP(clk), .CD(n1460), .Q(out1_1[35]) );
  CFD2QXL \out1_1_reg[34]  ( .D(n942), .CP(clk), .CD(n1461), .Q(out1_1[34]) );
  CFD2QXL \out1_1_reg[33]  ( .D(n940), .CP(clk), .CD(n1461), .Q(out1_1[33]) );
  CFD2QXL \out1_1_reg[32]  ( .D(n938), .CP(clk), .CD(n1461), .Q(out1_1[32]) );
  CFD2QXL \out1_1_reg[31]  ( .D(n936), .CP(clk), .CD(n1461), .Q(out1_1[31]) );
  CFD2QXL \out1_1_reg[30]  ( .D(n934), .CP(clk), .CD(n1443), .Q(out1_1[30]) );
  CFD2QXL \out1_1_reg[29]  ( .D(n932), .CP(clk), .CD(n1437), .Q(out1_1[29]) );
  CFD2QXL \out1_1_reg[28]  ( .D(n930), .CP(clk), .CD(n1437), .Q(out1_1[28]) );
  CFD2QXL \out1_1_reg[27]  ( .D(n928), .CP(clk), .CD(n1437), .Q(out1_1[27]) );
  CFD2QXL \out1_1_reg[26]  ( .D(n926), .CP(clk), .CD(n1437), .Q(out1_1[26]) );
  CFD2QXL \out1_1_reg[25]  ( .D(n924), .CP(clk), .CD(n1438), .Q(out1_1[25]) );
  CFD2QXL \out1_1_reg[24]  ( .D(n922), .CP(clk), .CD(n1438), .Q(out1_1[24]) );
  CFD2QXL \out1_1_reg[23]  ( .D(n920), .CP(clk), .CD(n1438), .Q(out1_1[23]) );
  CFD2QXL \out1_1_reg[22]  ( .D(n918), .CP(clk), .CD(n1438), .Q(out1_1[22]) );
  CFD2QXL \out1_1_reg[21]  ( .D(n916), .CP(clk), .CD(n1438), .Q(out1_1[21]) );
  CFD2QXL \out1_1_reg[20]  ( .D(n914), .CP(clk), .CD(n1438), .Q(out1_1[20]) );
  CFD2QXL \out1_1_reg[19]  ( .D(n912), .CP(clk), .CD(n1439), .Q(out1_1[19]) );
  CFD2QXL \out1_1_reg[18]  ( .D(n910), .CP(clk), .CD(n1439), .Q(out1_1[18]) );
  CFD2QXL \out1_1_reg[17]  ( .D(n908), .CP(clk), .CD(n1439), .Q(out1_1[17]) );
  CFD2QXL \out1_1_reg[16]  ( .D(n906), .CP(clk), .CD(n1439), .Q(out1_1[16]) );
  CFD2QXL \out1_1_reg[15]  ( .D(n904), .CP(clk), .CD(n1439), .Q(out1_1[15]) );
  CFD2QXL \out1_1_reg[14]  ( .D(n902), .CP(clk), .CD(n1439), .Q(out1_1[14]) );
  CFD2QXL \out1_1_reg[13]  ( .D(n900), .CP(clk), .CD(n1439), .Q(out1_1[13]) );
  CFD2QXL \out1_1_reg[12]  ( .D(n898), .CP(clk), .CD(n1440), .Q(out1_1[12]) );
  CFD2QXL \out1_1_reg[11]  ( .D(n896), .CP(clk), .CD(n1440), .Q(out1_1[11]) );
  CFD2QXL \out1_1_reg[10]  ( .D(n894), .CP(clk), .CD(n1440), .Q(out1_1[10]) );
  CFD2QXL \out1_1_reg[9]  ( .D(n892), .CP(clk), .CD(n1440), .Q(out1_1[9]) );
  CFD2QXL \out1_1_reg[8]  ( .D(n890), .CP(clk), .CD(n1440), .Q(out1_1[8]) );
  CFD2QXL \out1_1_reg[7]  ( .D(n888), .CP(clk), .CD(n1440), .Q(out1_1[7]) );
  CFD2QXL \out1_1_reg[6]  ( .D(n886), .CP(clk), .CD(n1441), .Q(out1_1[6]) );
  CFD2QXL \out1_1_reg[5]  ( .D(n884), .CP(clk), .CD(n1441), .Q(out1_1[5]) );
  CFD2QXL \out1_1_reg[4]  ( .D(n882), .CP(clk), .CD(n1441), .Q(out1_1[4]) );
  CFD2QXL \out1_1_reg[3]  ( .D(n880), .CP(clk), .CD(n1441), .Q(out1_1[3]) );
  CFD2QXL \out1_1_reg[2]  ( .D(n878), .CP(clk), .CD(n1441), .Q(out1_1[2]) );
  CFD2QXL \out1_1_reg[1]  ( .D(n876), .CP(clk), .CD(n1441), .Q(out1_1[1]) );
  CFD2QXL \out1_1_reg[0]  ( .D(n874), .CP(clk), .CD(n1442), .Q(out1_1[0]) );
  CFD2QXL \out0_2_reg[60]  ( .D(n694), .CP(clk), .CD(n1443), .Q(out0_2[60]) );
  CFD2QXL \out0_2_reg[61]  ( .D(n693), .CP(clk), .CD(n1442), .Q(out0_2[61]) );
  CFD2QXL \out0_2_reg[62]  ( .D(n692), .CP(clk), .CD(n1442), .Q(out0_2[62]) );
  CFD2QXL \out0_2_reg[63]  ( .D(n691), .CP(clk), .CD(n1456), .Q(out0_2[63]) );
  CFD2QXL \out0_2_reg[39]  ( .D(n873), .CP(clk), .CD(n1473), .Q(out0_2[39]) );
  CFD2QXL \out0_2_reg[45]  ( .D(n871), .CP(clk), .CD(n1449), .Q(out0_2[45]) );
  CFD2QXL \out0_2_reg[7]  ( .D(n870), .CP(clk), .CD(n1463), .Q(out0_2[7]) );
  CFD2QXL \out0_2_reg[15]  ( .D(n869), .CP(clk), .CD(n1483), .Q(out0_2[15]) );
  CFD2QXL \out0_2_reg[42]  ( .D(n868), .CP(clk), .CD(n1472), .Q(out0_2[42]) );
  CFD2QXL \out0_2_reg[27]  ( .D(n867), .CP(clk), .CD(n1478), .Q(out0_2[27]) );
  CFD2QXL \out0_2_reg[40]  ( .D(n866), .CP(clk), .CD(n1473), .Q(out0_2[40]) );
  CFD2QXL \out0_2_reg[0]  ( .D(n865), .CP(clk), .CD(n1455), .Q(out0_2[0]) );
  CFD2QXL \out0_2_reg[5]  ( .D(n864), .CP(clk), .CD(n1464), .Q(out0_2[5]) );
  CFD2QXL \out0_2_reg[25]  ( .D(n863), .CP(clk), .CD(n1479), .Q(out0_2[25]) );
  CFD2QXL \out0_2_reg[13]  ( .D(n862), .CP(clk), .CD(n1483), .Q(out0_2[13]) );
  CFD2QXL \out0_2_reg[34]  ( .D(n861), .CP(clk), .CD(n1475), .Q(out0_2[34]) );
  CFD2QXL \out0_2_reg[19]  ( .D(n860), .CP(clk), .CD(n1481), .Q(out0_2[19]) );
  CFD2QXL \out0_2_reg[10]  ( .D(n859), .CP(clk), .CD(n1462), .Q(out0_2[10]) );
  CFD2QXL \out0_2_reg[3]  ( .D(n858), .CP(clk), .CD(n1465), .Q(out0_2[3]) );
  CFD2QXL \out0_2_reg[32]  ( .D(n856), .CP(clk), .CD(n1476), .Q(out0_2[32]) );
  CFD2QXL \out0_2_reg[17]  ( .D(n855), .CP(clk), .CD(n1482), .Q(out0_2[17]) );
  CFD2QXL \out0_2_reg[43]  ( .D(n854), .CP(clk), .CD(n1472), .Q(out0_2[43]) );
  CFD2QXL \out0_2_reg[41]  ( .D(n853), .CP(clk), .CD(n1473), .Q(out0_2[41]) );
  CFD2QXL \out0_2_reg[35]  ( .D(n852), .CP(clk), .CD(n1475), .Q(out0_2[35]) );
  CFD2QXL \out0_2_reg[11]  ( .D(n851), .CP(clk), .CD(n1462), .Q(out0_2[11]) );
  CFD2QXL \out0_2_reg[33]  ( .D(n850), .CP(clk), .CD(n1476), .Q(out0_2[33]) );
  CFD2QXL \out0_2_reg[9]  ( .D(n849), .CP(clk), .CD(n1462), .Q(out0_2[9]) );
  CFD2QXL \out0_2_reg[59]  ( .D(n848), .CP(clk), .CD(n1443), .Q(out0_2[59]) );
  CFD2QXL \out1_2_reg[0]  ( .D(n545), .CP(clk), .CD(n1466), .Q(out1_2[0]) );
  CFD2QXL \out0_2_reg[2]  ( .D(n847), .CP(clk), .CD(n1465), .Q(out0_2[2]) );
  CFD2QXL \out0_2_reg[31]  ( .D(n846), .CP(clk), .CD(n1476), .Q(out0_2[31]) );
  CFD2QXL \out0_2_reg[4]  ( .D(n845), .CP(clk), .CD(n1464), .Q(out0_2[4]) );
  CFD2QXL \out0_2_reg[55]  ( .D(n844), .CP(clk), .CD(n1445), .Q(out0_2[55]) );
  CFD2QXL \out0_2_reg[56]  ( .D(n843), .CP(clk), .CD(n1444), .Q(out0_2[56]) );
  CFD2QXL \out0_2_reg[57]  ( .D(n842), .CP(clk), .CD(n1444), .Q(out0_2[57]) );
  CFD2QXL \out0_2_reg[26]  ( .D(n841), .CP(clk), .CD(n1478), .Q(out0_2[26]) );
  CFD2QXL \out0_2_reg[29]  ( .D(n840), .CP(clk), .CD(n1477), .Q(out0_2[29]) );
  CFD2QXL \out0_2_reg[37]  ( .D(n839), .CP(clk), .CD(n1474), .Q(out0_2[37]) );
  CFD2QXL \out0_2_reg[51]  ( .D(n838), .CP(clk), .CD(n1446), .Q(out0_2[51]) );
  CFD2QXL \out0_2_reg[50]  ( .D(n837), .CP(clk), .CD(n1447), .Q(out0_2[50]) );
  CFD2QXL \out0_2_reg[21]  ( .D(n836), .CP(clk), .CD(n1480), .Q(out0_2[21]) );
  CFD2QXL \out0_2_reg[53]  ( .D(n835), .CP(clk), .CD(n1446), .Q(out0_2[53]) );
  CFD2QXL \out0_2_reg[12]  ( .D(n834), .CP(clk), .CD(n1467), .Q(out0_2[12]) );
  CFD2QXL \out0_2_reg[44]  ( .D(n833), .CP(clk), .CD(n1449), .Q(out0_2[44]) );
  CFD2QXL \out0_2_reg[28]  ( .D(n832), .CP(clk), .CD(n1478), .Q(out0_2[28]) );
  CFD2QXL \out0_2_reg[6]  ( .D(n831), .CP(clk), .CD(n1463), .Q(out0_2[6]) );
  CFD2QXL \out0_2_reg[58]  ( .D(n830), .CP(clk), .CD(n1444), .Q(out0_2[58]) );
  CFD2QXL \out0_2_reg[30]  ( .D(n829), .CP(clk), .CD(n1477), .Q(out0_2[30]) );
  CFD2QXL \out0_2_reg[24]  ( .D(n828), .CP(clk), .CD(n1479), .Q(out0_2[24]) );
  CFD2QXL \out0_2_reg[49]  ( .D(n827), .CP(clk), .CD(n1447), .Q(out0_2[49]) );
  CFD2QXL \out0_2_reg[14]  ( .D(n826), .CP(clk), .CD(n1483), .Q(out0_2[14]) );
  CFD2QXL \out0_2_reg[52]  ( .D(n825), .CP(clk), .CD(n1446), .Q(out0_2[52]) );
  CFD2QXL \out0_2_reg[47]  ( .D(n824), .CP(clk), .CD(n1448), .Q(out0_2[47]) );
  CFD2QXL \out0_2_reg[18]  ( .D(n823), .CP(clk), .CD(n1482), .Q(out0_2[18]) );
  CFD2QXL \out0_2_reg[54]  ( .D(n822), .CP(clk), .CD(n1445), .Q(out0_2[54]) );
  CFD2QXL \out0_2_reg[38]  ( .D(n821), .CP(clk), .CD(n1474), .Q(out0_2[38]) );
  CFD2QXL \out0_2_reg[48]  ( .D(n820), .CP(clk), .CD(n1447), .Q(out0_2[48]) );
  CFD2QXL \out0_2_reg[20]  ( .D(n819), .CP(clk), .CD(n1481), .Q(out0_2[20]) );
  CFD2QXL \out0_2_reg[36]  ( .D(n818), .CP(clk), .CD(n1474), .Q(out0_2[36]) );
  CFD2QXL \out0_2_reg[23]  ( .D(n817), .CP(clk), .CD(n1480), .Q(out0_2[23]) );
  CFD2QXL \out0_2_reg[22]  ( .D(n816), .CP(clk), .CD(n1480), .Q(out0_2[22]) );
  CFD2QXL \out0_2_reg[46]  ( .D(n815), .CP(clk), .CD(n1448), .Q(out0_2[46]) );
  CFD2QXL \out1_2_reg[1]  ( .D(n543), .CP(clk), .CD(n1465), .Q(out1_2[1]) );
  CFD2QXL \out1_2_reg[3]  ( .D(n539), .CP(clk), .CD(n1465), .Q(out1_2[3]) );
  CFD2QXL \out1_2_reg[2]  ( .D(n541), .CP(clk), .CD(n1465), .Q(out1_2[2]) );
  CFD2QXL \out1_2_reg[4]  ( .D(n537), .CP(clk), .CD(n1464), .Q(out1_2[4]) );
  CFD2QXL \out1_2_reg[21]  ( .D(n503), .CP(clk), .CD(n1480), .Q(out1_2[21]) );
  CFD2QXL \out1_2_reg[19]  ( .D(n507), .CP(clk), .CD(n1481), .Q(out1_2[19]) );
  CFD2QXL \out1_2_reg[18]  ( .D(n509), .CP(clk), .CD(n1482), .Q(out1_2[18]) );
  CFD2QXL \out1_2_reg[17]  ( .D(n511), .CP(clk), .CD(n1482), .Q(out1_2[17]) );
  CFD2QXL \out1_2_reg[20]  ( .D(n505), .CP(clk), .CD(n1481), .Q(out1_2[20]) );
  CFD2QXL \acc_reg[5]  ( .D(n534), .CP(clk), .CD(n1464), .Q(acc[5]) );
  CFD2QXL \acc_reg[25]  ( .D(n494), .CP(clk), .CD(n1479), .Q(acc[25]) );
  CFD2QXL \acc_reg[13]  ( .D(n518), .CP(clk), .CD(n1484), .Q(acc[13]) );
  CFD2QXL \acc_reg[19]  ( .D(n506), .CP(clk), .CD(n1481), .Q(acc[19]) );
  CFD2QXL \acc_reg[10]  ( .D(n524), .CP(clk), .CD(n1462), .Q(acc[10]) );
  CFD2QXL \acc_reg[8]  ( .D(n528), .CP(clk), .CD(n1463), .Q(acc[8]) );
  CFD2QXL \acc_reg[3]  ( .D(n538), .CP(clk), .CD(n1465), .Q(acc[3]) );
  CFD2QXL \acc_reg[17]  ( .D(n510), .CP(clk), .CD(n1482), .Q(acc[17]) );
  CFD2QXL \acc_reg[11]  ( .D(n522), .CP(clk), .CD(n1462), .Q(acc[11]) );
  CFD2QXL \acc_reg[9]  ( .D(n526), .CP(clk), .CD(n1462), .Q(acc[9]) );
  CFD2QXL \acc_reg[1]  ( .D(n542), .CP(clk), .CD(n1466), .Q(acc[1]) );
  CFD2QXL \acc_reg[2]  ( .D(n540), .CP(clk), .CD(n1465), .Q(acc[2]) );
  CFD2QXL \acc_reg[31]  ( .D(n482), .CP(clk), .CD(n1477), .Q(acc[31]) );
  CFD2QXL \acc_reg[4]  ( .D(n536), .CP(clk), .CD(n1464), .Q(acc[4]) );
  CFD2QXL \acc_reg[7]  ( .D(n530), .CP(clk), .CD(n1463), .Q(acc[7]) );
  CFD2QXL \acc_reg[26]  ( .D(n492), .CP(clk), .CD(n1479), .Q(acc[26]) );
  CFD2QXL \acc_reg[29]  ( .D(n486), .CP(clk), .CD(n1477), .Q(acc[29]) );
  CFD2QXL \acc_reg[15]  ( .D(n514), .CP(clk), .CD(n1483), .Q(acc[15]) );
  CFD2QXL \acc_reg[27]  ( .D(n490), .CP(clk), .CD(n1478), .Q(acc[27]) );
  CFD2QXL \acc_reg[21]  ( .D(n502), .CP(clk), .CD(n1481), .Q(acc[21]) );
  CFD2QXL \acc_reg[12]  ( .D(n520), .CP(clk), .CD(n1461), .Q(acc[12]) );
  CFD2QXL \acc_reg[28]  ( .D(n488), .CP(clk), .CD(n1478), .Q(acc[28]) );
  CFD2QXL \acc_reg[6]  ( .D(n532), .CP(clk), .CD(n1464), .Q(acc[6]) );
  CFD2QXL \acc_reg[16]  ( .D(n512), .CP(clk), .CD(n1482), .Q(acc[16]) );
  CFD2QXL \acc_reg[30]  ( .D(n484), .CP(clk), .CD(n1477), .Q(acc[30]) );
  CFD2QXL \acc_reg[24]  ( .D(n496), .CP(clk), .CD(n1479), .Q(acc[24]) );
  CFD2QXL \acc_reg[14]  ( .D(n516), .CP(clk), .CD(n1483), .Q(acc[14]) );
  CFD2QXL \acc_reg[18]  ( .D(n508), .CP(clk), .CD(n1482), .Q(acc[18]) );
  CFD2QXL \acc_reg[20]  ( .D(n504), .CP(clk), .CD(n1481), .Q(acc[20]) );
  CFD2QXL \acc_reg[23]  ( .D(n498), .CP(clk), .CD(n1480), .Q(acc[23]) );
  CFD2QXL \acc_reg[22]  ( .D(n500), .CP(clk), .CD(n1479), .Q(acc[22]) );
  CFD2QXL \cmd0_2_reg[0]  ( .D(n812), .CP(clk), .CD(n1449), .Q(cmd0_2[0]) );
  CFD2QXL \acc_reg[0]  ( .D(n544), .CP(clk), .CD(n1469), .Q(acc[0]) );
  CFD2QXL \cmd0_2_reg[1]  ( .D(n810), .CP(clk), .CD(n1450), .Q(cmd0_2[1]) );
  CFD2QXL \out2_2_reg[3]  ( .D(n607), .CP(clk), .CD(n1469), .Q(out2_2[3]) );
  CFD2QXL \out2_2_reg[5]  ( .D(n807), .CP(clk), .CD(n1468), .Q(out2_2[5]) );
  CFD2QXL _pushout_reg ( .D(n798), .CP(clk), .CD(n1455), .Q(pushout) );
  CFD2QXL \out0_0_reg[63]  ( .D(N78), .CP(clk), .CD(n1456), .Q(out0_0[63]) );
  CFD2QXL \out0_0_reg[41]  ( .D(N56), .CP(clk), .CD(n1472), .Q(out0_0[41]) );
  CFD2QXL \out0_0_reg[40]  ( .D(N55), .CP(clk), .CD(n1473), .Q(out0_0[40]) );
  CFD2QXL \out0_0_reg[39]  ( .D(N54), .CP(clk), .CD(n1473), .Q(out0_0[39]) );
  CFD2QXL \out0_0_reg[38]  ( .D(N53), .CP(clk), .CD(n1474), .Q(out0_0[38]) );
  CFD2QXL \out0_0_reg[37]  ( .D(N52), .CP(clk), .CD(n1474), .Q(out0_0[37]) );
  CFD2QXL \out0_0_reg[36]  ( .D(N51), .CP(clk), .CD(n1474), .Q(out0_0[36]) );
  CFD2QXL \out0_0_reg[35]  ( .D(N50), .CP(clk), .CD(n1475), .Q(out0_0[35]) );
  CFD2QXL \out0_0_reg[34]  ( .D(N49), .CP(clk), .CD(n1475), .Q(out0_0[34]) );
  CFD2QXL \out0_0_reg[33]  ( .D(N48), .CP(clk), .CD(n1475), .Q(out0_0[33]) );
  CFD2QXL \out0_0_reg[32]  ( .D(N47), .CP(clk), .CD(n1476), .Q(out0_0[32]) );
  CFD2QXL \out0_0_reg[31]  ( .D(N46), .CP(clk), .CD(n1476), .Q(out0_0[31]) );
  CFD2QXL \out0_0_reg[30]  ( .D(N45), .CP(clk), .CD(n1477), .Q(out0_0[30]) );
  CFD2QXL \out0_0_reg[29]  ( .D(N44), .CP(clk), .CD(n1477), .Q(out0_0[29]) );
  CFD2QXL \out0_0_reg[28]  ( .D(N43), .CP(clk), .CD(n1477), .Q(out0_0[28]) );
  CFD2QXL \out0_0_reg[27]  ( .D(N42), .CP(clk), .CD(n1478), .Q(out0_0[27]) );
  CFD2QXL \out0_0_reg[26]  ( .D(N41), .CP(clk), .CD(n1478), .Q(out0_0[26]) );
  CFD2QXL \out0_0_reg[25]  ( .D(N40), .CP(clk), .CD(n1479), .Q(out0_0[25]) );
  CFD2QXL \out0_0_reg[24]  ( .D(N39), .CP(clk), .CD(n1479), .Q(out0_0[24]) );
  CFD2QXL \out0_0_reg[23]  ( .D(N38), .CP(clk), .CD(n1479), .Q(out0_0[23]) );
  CFD2QXL \out0_0_reg[22]  ( .D(N37), .CP(clk), .CD(n1480), .Q(out0_0[22]) );
  CFD2QXL \out0_0_reg[21]  ( .D(N36), .CP(clk), .CD(n1480), .Q(out0_0[21]) );
  CFD2QXL \out0_0_reg[20]  ( .D(N35), .CP(clk), .CD(n1481), .Q(out0_0[20]) );
  CFD2QXL \out0_0_reg[19]  ( .D(N34), .CP(clk), .CD(n1481), .Q(out0_0[19]) );
  CFD2QXL \out0_0_reg[18]  ( .D(N33), .CP(clk), .CD(n1480), .Q(out0_0[18]) );
  CFD2QXL \out0_0_reg[17]  ( .D(N32), .CP(clk), .CD(n1482), .Q(out0_0[17]) );
  CFD2QXL \out0_0_reg[16]  ( .D(N31), .CP(clk), .CD(n1482), .Q(out0_0[16]) );
  CFD2QXL \out0_0_reg[14]  ( .D(N29), .CP(clk), .CD(n1483), .Q(out0_0[14]) );
  CFD2QXL \out0_0_reg[7]  ( .D(N22), .CP(clk), .CD(n1463), .Q(out0_0[7]) );
  CFD2QXL \out0_0_reg[6]  ( .D(N21), .CP(clk), .CD(n1463), .Q(out0_0[6]) );
  CFD2QXL \out0_0_reg[5]  ( .D(N20), .CP(clk), .CD(n1464), .Q(out0_0[5]) );
  CFD2QXL \out0_0_reg[4]  ( .D(N19), .CP(clk), .CD(n1464), .Q(out0_0[4]) );
  CFD2QXL \out0_0_reg[3]  ( .D(N18), .CP(clk), .CD(n1464), .Q(out0_0[3]) );
  CFD2QXL \out0_0_reg[2]  ( .D(N17), .CP(clk), .CD(n1465), .Q(out0_0[2]) );
  CFD2QXL \out0_0_reg[1]  ( .D(N16), .CP(clk), .CD(n1465), .Q(out0_0[1]) );
  CFD2QXL \out0_0_reg[0]  ( .D(N15), .CP(clk), .CD(n1454), .Q(out0_0[0]) );
  CFD2QXL \out1_0_reg[63]  ( .D(N78), .CP(clk), .CD(n1456), .Q(out1_0[63]) );
  CFD2QXL \out1_0_reg[40]  ( .D(N55), .CP(clk), .CD(n1460), .Q(out1_0[40]) );
  CFD2QXL \out1_0_reg[39]  ( .D(N54), .CP(clk), .CD(n1460), .Q(out1_0[39]) );
  CFD2QXL \out1_0_reg[38]  ( .D(N53), .CP(clk), .CD(n1460), .Q(out1_0[38]) );
  CFD2QXL \out1_0_reg[37]  ( .D(N52), .CP(clk), .CD(n1460), .Q(out1_0[37]) );
  CFD2QXL \out1_0_reg[36]  ( .D(N51), .CP(clk), .CD(n1460), .Q(out1_0[36]) );
  CFD2QXL \out1_0_reg[35]  ( .D(N50), .CP(clk), .CD(n1460), .Q(out1_0[35]) );
  CFD2QXL \out1_0_reg[34]  ( .D(N49), .CP(clk), .CD(n1460), .Q(out1_0[34]) );
  CFD2QXL \out1_0_reg[33]  ( .D(N48), .CP(clk), .CD(n1461), .Q(out1_0[33]) );
  CFD2QXL \out1_0_reg[32]  ( .D(N47), .CP(clk), .CD(n1461), .Q(out1_0[32]) );
  CFD2QXL \out1_0_reg[31]  ( .D(N46), .CP(clk), .CD(n1461), .Q(out1_0[31]) );
  CFD2QXL \out1_0_reg[30]  ( .D(N45), .CP(clk), .CD(n1461), .Q(out1_0[30]) );
  CFD2QXL \out1_0_reg[29]  ( .D(N44), .CP(clk), .CD(n1437), .Q(out1_0[29]) );
  CFD2QXL \out1_0_reg[28]  ( .D(N43), .CP(clk), .CD(n1437), .Q(out1_0[28]) );
  CFD2QXL \out1_0_reg[27]  ( .D(N42), .CP(clk), .CD(n1437), .Q(out1_0[27]) );
  CFD2QXL \out1_0_reg[26]  ( .D(N41), .CP(clk), .CD(n1438), .Q(out1_0[26]) );
  CFD2QXL \out1_0_reg[25]  ( .D(N40), .CP(clk), .CD(n1438), .Q(out1_0[25]) );
  CFD2QXL \out1_0_reg[24]  ( .D(N39), .CP(clk), .CD(n1438), .Q(out1_0[24]) );
  CFD2QXL \out1_0_reg[23]  ( .D(N38), .CP(clk), .CD(n1438), .Q(out1_0[23]) );
  CFD2QXL \out1_0_reg[22]  ( .D(N37), .CP(clk), .CD(n1438), .Q(out1_0[22]) );
  CFD2QXL \out1_0_reg[21]  ( .D(N36), .CP(clk), .CD(n1438), .Q(out1_0[21]) );
  CFD2QXL \out1_0_reg[20]  ( .D(N35), .CP(clk), .CD(n1438), .Q(out1_0[20]) );
  CFD2QXL \out1_0_reg[19]  ( .D(N34), .CP(clk), .CD(n1439), .Q(out1_0[19]) );
  CFD2QXL \out1_0_reg[18]  ( .D(N33), .CP(clk), .CD(n1439), .Q(out1_0[18]) );
  CFD2QXL \out1_0_reg[17]  ( .D(N32), .CP(clk), .CD(n1439), .Q(out1_0[17]) );
  CFD2QXL \out1_0_reg[16]  ( .D(N31), .CP(clk), .CD(n1439), .Q(out1_0[16]) );
  CFD2QXL \out1_0_reg[14]  ( .D(N29), .CP(clk), .CD(n1439), .Q(out1_0[14]) );
  CFD2QXL \out1_0_reg[7]  ( .D(N22), .CP(clk), .CD(n1440), .Q(out1_0[7]) );
  CFD2QXL \out1_0_reg[6]  ( .D(N21), .CP(clk), .CD(n1441), .Q(out1_0[6]) );
  CFD2QXL \out1_0_reg[5]  ( .D(N20), .CP(clk), .CD(n1441), .Q(out1_0[5]) );
  CFD2QXL \out1_0_reg[4]  ( .D(N19), .CP(clk), .CD(n1441), .Q(out1_0[4]) );
  CFD2QXL \out1_0_reg[3]  ( .D(N18), .CP(clk), .CD(n1441), .Q(out1_0[3]) );
  CFD2QXL \out1_0_reg[2]  ( .D(N17), .CP(clk), .CD(n1441), .Q(out1_0[2]) );
  CFD2QXL \out1_0_reg[1]  ( .D(N16), .CP(clk), .CD(n1441), .Q(out1_0[1]) );
  CFD2QXL \out1_0_reg[0]  ( .D(N15), .CP(clk), .CD(n1441), .Q(out1_0[0]) );
  CFD2QXL \cmd0_0_reg[1]  ( .D(n1211), .CP(clk), .CD(n1450), .Q(cmd0_0[1]) );
  CFD2QXL \cmd0_1_reg[1]  ( .D(n1235), .CP(clk), .CD(n1450), .Q(cmd0_1[1]) );
  CFD2QXL \cmd0_0_reg[0]  ( .D(n1213), .CP(clk), .CD(n1449), .Q(cmd0_0[0]) );
  CFD2QXL \cmd0_1_reg[0]  ( .D(n1237), .CP(clk), .CD(n1449), .Q(cmd0_1[0]) );
  CFD2QXL push0_0_reg ( .D(n1215), .CP(clk), .CD(n1449), .Q(push0_0) );
  CFD2QXL push0_1_reg ( .D(n1239), .CP(clk), .CD(n1449), .Q(push0_1) );
  CFD2QX1 \h0_1_reg[3]  ( .D(n621), .CP(clk), .CD(n1466), .Q(h0_1[3]) );
  CFD2QXL \h0_1_reg[0]  ( .D(n1223), .CP(clk), .CD(n1456), .Q(h0_1[0]) );
  CFD2QXL \out0_2_reg[8]  ( .D(n1222), .CP(clk), .CD(n1463), .Q(out0_2[8]) );
  CFD2QXL \out0_2_reg[16]  ( .D(n1221), .CP(clk), .CD(n1482), .Q(out0_2[16])
         );
  CFD2QXL \h0_1_reg[1]  ( .D(n615), .CP(clk), .CD(n1455), .Q(h0_1[1]) );
  CFD2QX1 \q0_reg[19]  ( .D(n677), .CP(clk), .CD(n1451), .Q(q0[19]) );
  CFD2QX2 \h0_1_reg[2]  ( .D(n618), .CP(clk), .CD(n1456), .Q(h0_1[2]) );
  CFD2QX2 \q0_reg[20]  ( .D(n1163), .CP(clk), .CD(n1450), .Q(q0[20]) );
  CFD2QXL cmd1_en_2_d_reg ( .D(n1429), .CP(clk), .CD(n1442), .Q(cmd1_en_2_d)
         );
  CFD2QX2 \h0_reg[2]  ( .D(n620), .CP(clk), .CD(n1454), .Q(h0[2]) );
  CFD2QX2 \h0_reg[4]  ( .D(n626), .CP(clk), .CD(n1454), .Q(h0[4]) );
  CFD2QX4 \h0_reg[1]  ( .D(n617), .CP(clk), .CD(n1454), .Q(h0[1]) );
  CFD2QX1 \h0_reg[0]  ( .D(n614), .CP(clk), .CD(n1454), .Q(h0[0]) );
  CFD2QX4 \h0_reg[26]  ( .D(n652), .CP(clk), .CD(n1452), .Q(h0[26]) );
  CFD2QX2 \h0_reg[18]  ( .D(n1202), .CP(clk), .CD(n1453), .Q(h0[18]) );
  CFD2QX4 \h0_reg[30]  ( .D(n656), .CP(clk), .CD(n1452), .Q(h0[30]) );
  CFD2QX4 \h0_reg[29]  ( .D(n655), .CP(clk), .CD(n1452), .Q(h0[29]) );
  CFD2QX4 \h0_reg[13]  ( .D(n639), .CP(clk), .CD(n1453), .Q(h0[13]) );
  CFD2QX4 \h0_reg[19]  ( .D(n645), .CP(clk), .CD(n1453), .Q(h0[19]) );
  CFD2QX1 \h0_reg[8]  ( .D(n634), .CP(clk), .CD(n1454), .Q(h0[8]) );
  CFD2QX1 \h0_reg[31]  ( .D(n1200), .CP(clk), .CD(n1452), .Q(h0[31]) );
  CFD2QX1 \h0_reg[9]  ( .D(n1199), .CP(clk), .CD(n1454), .Q(h0[9]) );
  CFD2QX1 \h0_reg[17]  ( .D(n1198), .CP(clk), .CD(n1453), .Q(h0[17]) );
  CFD2QX1 \h0_reg[27]  ( .D(n1197), .CP(clk), .CD(n1452), .Q(h0[27]) );
  CFD2QX1 \h0_reg[22]  ( .D(n1196), .CP(clk), .CD(n1453), .Q(h0[22]) );
  CFD2QX4 \h0_reg[28]  ( .D(n654), .CP(clk), .CD(n1452), .Q(h0[28]) );
  CFD2QX1 \h0_reg[23]  ( .D(n1193), .CP(clk), .CD(n1453), .Q(h0[23]) );
  CFD2QX1 \h0_reg[21]  ( .D(n1192), .CP(clk), .CD(n1453), .Q(h0[21]) );
  CFD2QX1 \h0_reg[14]  ( .D(n1191), .CP(clk), .CD(n1453), .Q(h0[14]) );
  CFD2QX1 \q0_reg[11]  ( .D(n669), .CP(clk), .CD(n1451), .Q(q0[11]) );
  CFD2QX1 \h0_reg[10]  ( .D(n1190), .CP(clk), .CD(n1454), .Q(h0[10]) );
  CFD2QX1 \h0_reg[16]  ( .D(n1189), .CP(clk), .CD(n1453), .Q(h0[16]) );
  CFD2QX1 \h0_reg[20]  ( .D(n1188), .CP(clk), .CD(n1453), .Q(h0[20]) );
  CFD2QX1 \h0_reg[7]  ( .D(n1187), .CP(clk), .CD(n1454), .Q(h0[7]) );
  CFD2QX1 \h0_reg[11]  ( .D(n998), .CP(clk), .CD(n1454), .Q(h0[11]) );
  CFD2QX1 \h0_reg[25]  ( .D(n857), .CP(clk), .CD(n1452), .Q(h0[25]) );
  CFD2QX1 \q0_reg[31]  ( .D(n872), .CP(clk), .CD(n1450), .Q(q0[31]) );
  CFD2QX1 \h0_reg[24]  ( .D(n814), .CP(clk), .CD(n1453), .Q(h0[24]) );
  CFD2QX2 \q0_reg[5]  ( .D(n808), .CP(clk), .CD(n1452), .Q(q0[5]) );
  CFD2QX2 \q0_reg[3]  ( .D(n661), .CP(clk), .CD(n1452), .Q(q0[3]) );
  CFD2QX2 \q0_reg[9]  ( .D(n667), .CP(clk), .CD(n1451), .Q(q0[9]) );
  CFD2QX2 \q0_reg[17]  ( .D(n675), .CP(clk), .CD(n1451), .Q(q0[17]) );
  CFD2QX2 \q0_reg[18]  ( .D(n676), .CP(clk), .CD(n1451), .Q(q0[18]) );
  CFD2QX2 \q0_reg[12]  ( .D(n670), .CP(clk), .CD(n1451), .Q(q0[12]) );
  CFD1XL cmd0_en_2_reg ( .D(n755), .CP(clk), .Q(cmd0_en_2), .QN(n1362) );
  CFD1XL cmd2_en_2_reg ( .D(n690), .CP(clk), .Q(cmd2_en_2), .QN(n1495) );
  CFD2XL \out0_2_reg[1]  ( .D(n1160), .CP(clk), .CD(n2462), .Q(out0_2[1]), 
        .QN(n2392) );
  CFD2XL \out1_0_reg[8]  ( .D(N23), .CP(clk), .CD(n2462), .Q(out1_0[8]) );
  CFD2XL \out0_0_reg[8]  ( .D(N23), .CP(clk), .CD(n2462), .Q(out0_0[8]) );
  CFD2XL \out2_2_reg[60]  ( .D(n1185), .CP(clk), .CD(n2462), .Q(out2_2[60]), 
        .QN(n1800) );
  CFD2XL \out2_2_reg[61]  ( .D(n1186), .CP(clk), .CD(n2462), .Q(out2_2[61]), 
        .QN(n1790) );
  CFD2XL \out1_2_reg[8]  ( .D(n529), .CP(clk), .CD(n2462), .Q(out1_2[8]), .QN(
        n1740) );
  CFD2XL \out1_2_reg[6]  ( .D(n533), .CP(clk), .CD(n2462), .Q(out1_2[6]), .QN(
        n1748) );
  CFD2XL \out1_2_reg[5]  ( .D(n535), .CP(clk), .CD(n2462), .Q(out1_2[5]), .QN(
        n1752) );
  CFD2XL \out1_2_reg[7]  ( .D(n531), .CP(clk), .CD(n2462), .Q(out1_2[7]), .QN(
        n1744) );
  CFD2XL \out1_0_reg[9]  ( .D(N24), .CP(clk), .CD(n2462), .Q(out1_0[9]) );
  CFD2XL \out0_0_reg[9]  ( .D(N24), .CP(clk), .CD(n2462), .Q(out0_0[9]) );
  CFD2XL \out2_2_reg[58]  ( .D(n1171), .CP(clk), .CD(n2462), .Q(out2_2[58]), 
        .QN(n1815) );
  CFD2XL \out2_2_reg[50]  ( .D(n1170), .CP(clk), .CD(n2462), .Q(out2_2[50]), 
        .QN(n1872) );
  CFD2XL \out1_2_reg[15]  ( .D(n515), .CP(clk), .CD(n2462), .Q(out1_2[15]), 
        .QN(n1712) );
  CFD2XL \out1_2_reg[14]  ( .D(n517), .CP(clk), .CD(n2462), .Q(out1_2[14]), 
        .QN(n1716) );
  CFD2XL \out1_2_reg[13]  ( .D(n519), .CP(clk), .CD(n2462), .Q(out1_2[13]), 
        .QN(n1720) );
  CFD2XL \out1_2_reg[12]  ( .D(n521), .CP(clk), .CD(n2462), .Q(out1_2[12]), 
        .QN(n1724) );
  CFD2XL \out1_2_reg[11]  ( .D(n523), .CP(clk), .CD(n2462), .Q(out1_2[11]), 
        .QN(n1728) );
  CFD2XL \out1_2_reg[10]  ( .D(n525), .CP(clk), .CD(n2462), .Q(out1_2[10]), 
        .QN(n1732) );
  CFD2XL \out1_2_reg[9]  ( .D(n527), .CP(clk), .CD(n2462), .Q(out1_2[9]), .QN(
        n1736) );
  CFD2XL \out2_2_reg[59]  ( .D(n1162), .CP(clk), .CD(n2462), .Q(out2_2[59]), 
        .QN(n1808) );
  CFD2XL \out2_2_reg[55]  ( .D(n1165), .CP(clk), .CD(n2462), .Q(out2_2[55]), 
        .QN(n1833) );
  CFD2XL \out2_2_reg[51]  ( .D(n1167), .CP(clk), .CD(n2462), .Q(out2_2[51]), 
        .QN(n1863) );
  CFD2XL \out2_2_reg[56]  ( .D(n1161), .CP(clk), .CD(n2462), .Q(out2_2[56]), 
        .QN(n1827) );
  CFD2XL \out2_2_reg[48]  ( .D(n1168), .CP(clk), .CD(n2462), .Q(out2_2[48]), 
        .QN(n1886) );
  CFD2XL \out2_2_reg[54]  ( .D(n1166), .CP(clk), .CD(n2462), .Q(out2_2[54]), 
        .QN(n1840) );
  CFD2XL \out2_2_reg[57]  ( .D(n1164), .CP(clk), .CD(n2462), .Q(out2_2[57]), 
        .QN(n1821) );
  CFD2XL \out2_2_reg[30]  ( .D(n580), .CP(clk), .CD(n2462), .Q(out2_2[30]) );
  CFD2XL \out2_2_reg[29]  ( .D(n581), .CP(clk), .CD(n2462), .Q(out2_2[29]) );
  CFD2XL \out2_2_reg[28]  ( .D(n582), .CP(clk), .CD(n2462), .Q(out2_2[28]) );
  CFD2XL \out2_2_reg[49]  ( .D(n1177), .CP(clk), .CD(n2462), .Q(out2_2[49]), 
        .QN(n1879) );
  CFD2XL \out2_2_reg[52]  ( .D(n1176), .CP(clk), .CD(n2462), .Q(out2_2[52]), 
        .QN(n1855) );
  CFD2XL \out2_2_reg[31]  ( .D(n579), .CP(clk), .CD(n2462), .Q(out2_2[31]) );
  CFD2XL \out1_0_reg[11]  ( .D(N26), .CP(clk), .CD(n2462), .Q(out1_0[11]) );
  CFD2XL \out0_0_reg[11]  ( .D(N26), .CP(clk), .CD(n2462), .Q(out0_0[11]) );
  CFD2XL \out2_2_reg[23]  ( .D(n587), .CP(clk), .CD(n2462), .Q(out2_2[23]) );
  CFD2XL \out2_2_reg[27]  ( .D(n583), .CP(clk), .CD(n2462), .Q(out2_2[27]) );
  CFD2XL \out1_0_reg[10]  ( .D(N25), .CP(clk), .CD(n2462), .Q(out1_0[10]) );
  CFD2XL \out0_0_reg[10]  ( .D(N25), .CP(clk), .CD(n2462), .Q(out0_0[10]) );
  CFD2XL \out2_2_reg[24]  ( .D(n586), .CP(clk), .CD(n2462), .Q(out2_2[24]) );
  CFD2XL \out2_2_reg[26]  ( .D(n584), .CP(clk), .CD(n2462), .Q(out2_2[26]) );
  CFD2XL \out2_2_reg[25]  ( .D(n585), .CP(clk), .CD(n2462), .Q(out2_2[25]) );
  CFD2XL \out2_2_reg[22]  ( .D(n588), .CP(clk), .CD(n2462), .Q(out2_2[22]) );
  CFD2XL \out2_2_reg[19]  ( .D(n591), .CP(clk), .CD(n2462), .Q(out2_2[19]) );
  CFD2XL \out2_2_reg[18]  ( .D(n592), .CP(clk), .CD(n2462), .Q(out2_2[18]) );
  CFD2XL \out2_2_reg[16]  ( .D(n594), .CP(clk), .CD(n2462), .Q(out2_2[16]) );
  CFD2XL \out2_2_reg[17]  ( .D(n593), .CP(clk), .CD(n2462), .Q(out2_2[17]) );
  CFD2XL \out2_2_reg[53]  ( .D(n1234), .CP(clk), .CD(n2462), .Q(out2_2[53]), 
        .QN(n1847) );
  CFD2XL \out1_2_reg[32]  ( .D(n481), .CP(clk), .CD(n2462), .Q(out1_2[32]), 
        .QN(n1644) );
  CFD2XL \out2_2_reg[47]  ( .D(n1233), .CP(clk), .CD(n2462), .Q(out2_2[47]), 
        .QN(n1896) );
  CFD2XL \out1_2_reg[16]  ( .D(n513), .CP(clk), .CD(n2462), .Q(out1_2[16]), 
        .QN(n1708) );
  CFD2XL \out2_2_reg[43]  ( .D(n799), .CP(clk), .CD(n2462), .Q(out2_2[43]), 
        .QN(n1933) );
  CFD2XL \out2_2_reg[20]  ( .D(n590), .CP(clk), .CD(n2462), .Q(out2_2[20]) );
  CFD2XL \out2_2_reg[46]  ( .D(n805), .CP(clk), .CD(n2462), .Q(out2_2[46]), 
        .QN(n1904) );
  CFD2XL \out2_2_reg[45]  ( .D(n806), .CP(clk), .CD(n2462), .Q(out2_2[45]), 
        .QN(n1913) );
  CFD2XL \out2_2_reg[44]  ( .D(n800), .CP(clk), .CD(n2462), .Q(out2_2[44]), 
        .QN(n1923) );
  CFD2XL \out2_2_reg[40]  ( .D(n804), .CP(clk), .CD(n2462), .Q(out2_2[40]), 
        .QN(n1960) );
  CFD2XL \out2_2_reg[42]  ( .D(n801), .CP(clk), .CD(n2462), .Q(out2_2[42]), 
        .QN(n1942) );
  CFD2XL \out2_2_reg[34]  ( .D(n803), .CP(clk), .CD(n2462), .Q(out2_2[34]), 
        .QN(n2014) );
  CFD2XL \out2_2_reg[32]  ( .D(n802), .CP(clk), .CD(n2462), .Q(out2_2[32]), 
        .QN(n2032) );
  CFD2XL \out2_2_reg[39]  ( .D(n1173), .CP(clk), .CD(n2462), .Q(out2_2[39]), 
        .QN(n1969) );
  CFD2XL \out2_2_reg[35]  ( .D(n1174), .CP(clk), .CD(n2462), .Q(out2_2[35]), 
        .QN(n2005) );
  CFD2XL \out2_2_reg[41]  ( .D(n1172), .CP(clk), .CD(n2462), .Q(out2_2[41]), 
        .QN(n1951) );
  CFD2XL \out2_2_reg[21]  ( .D(n589), .CP(clk), .CD(n2462), .Q(out2_2[21]) );
  CFD2XL \out2_2_reg[38]  ( .D(n1182), .CP(clk), .CD(n2462), .Q(out2_2[38]), 
        .QN(n1978) );
  CFD2XL \out2_2_reg[33]  ( .D(n1179), .CP(clk), .CD(n2462), .Q(out2_2[33]), 
        .QN(n2023) );
  CFD2XL \out2_2_reg[15]  ( .D(n595), .CP(clk), .CD(n2462), .Q(out2_2[15]) );
  CFD2XL \out2_2_reg[36]  ( .D(n1178), .CP(clk), .CD(n2462), .Q(out2_2[36]), 
        .QN(n1996) );
  CFD2XL \out2_2_reg[37]  ( .D(n1225), .CP(clk), .CD(n2462), .Q(out2_2[37]), 
        .QN(n1987) );
  CFD2XL \out1_0_reg[13]  ( .D(N28), .CP(clk), .CD(n2462), .Q(out1_0[13]) );
  CFD2XL \out0_0_reg[13]  ( .D(N28), .CP(clk), .CD(n2462), .Q(out0_0[13]) );
  CFD2XL \out1_0_reg[12]  ( .D(N27), .CP(clk), .CD(n2462), .Q(out1_0[12]) );
  CFD2XL \out0_0_reg[12]  ( .D(N27), .CP(clk), .CD(n2462), .Q(out0_0[12]) );
  CFD2XL \out2_2_reg[14]  ( .D(n1194), .CP(clk), .CD(n2462), .Q(out2_2[14]), 
        .QN(n2230) );
  CFD2XL \out2_2_reg[13]  ( .D(n1159), .CP(clk), .CD(n2462), .Q(out2_2[13]), 
        .QN(n2242) );
  CFD2XL \out2_2_reg[12]  ( .D(n1195), .CP(clk), .CD(n2462), .Q(out2_2[12]), 
        .QN(n2254) );
  CFD2XL \out2_2_reg[11]  ( .D(n1227), .CP(clk), .CD(n2462), .Q(out2_2[11]), 
        .QN(n2267) );
  CFD2XL \out2_2_reg[10]  ( .D(n1209), .CP(clk), .CD(n2462), .Q(out2_2[10]), 
        .QN(n2280) );
  CFD2XL \out2_2_reg[9]  ( .D(n1231), .CP(clk), .CD(n2462), .Q(out2_2[9]), 
        .QN(n2293) );
  CFD2XL \out2_2_reg[8]  ( .D(n1230), .CP(clk), .CD(n2462), .Q(out2_2[8]), 
        .QN(n2306) );
  CFD2XL \out2_2_reg[7]  ( .D(n1226), .CP(clk), .CD(n2462), .Q(out2_2[7]), 
        .QN(n2319) );
  CFD2XL \out2_2_reg[6]  ( .D(n1232), .CP(clk), .CD(n2462), .Q(out2_2[6]), 
        .QN(n2332) );
  CFD2XL \out2_2_reg[2]  ( .D(n1228), .CP(clk), .CD(n2462), .Q(out2_2[2]), 
        .QN(n2389) );
  CFD2XL \out2_2_reg[1]  ( .D(n1229), .CP(clk), .CD(n2462), .Q(out2_2[1]), 
        .QN(n2403) );
  CFD2XL \out2_2_reg[0]  ( .D(n1210), .CP(clk), .CD(n2462), .Q(out2_2[0]), 
        .QN(n2425) );
  CFD2XL \out1_0_reg[15]  ( .D(N30), .CP(clk), .CD(n2462), .Q(out1_0[15]) );
  CFD2XL \out0_0_reg[15]  ( .D(N30), .CP(clk), .CD(n2462), .Q(out0_0[15]) );
  CFD2XL \out1_2_reg[63]  ( .D(n419), .CP(clk), .CD(n2462), .Q(out1_2[63]), 
        .QN(n1518) );
  CFD2XL \out1_2_reg[62]  ( .D(n421), .CP(clk), .CD(n2462), .Q(out1_2[62]), 
        .QN(n1524) );
  CFD2XL \out1_2_reg[61]  ( .D(n423), .CP(clk), .CD(n2462), .Q(out1_2[61]), 
        .QN(n1528) );
  CFD2XL \out1_2_reg[60]  ( .D(n425), .CP(clk), .CD(n2462), .Q(out1_2[60]), 
        .QN(n1532) );
  CFD2XL \out1_2_reg[59]  ( .D(n427), .CP(clk), .CD(n2462), .Q(out1_2[59]), 
        .QN(n1536) );
  CFD2XL \out1_2_reg[58]  ( .D(n429), .CP(clk), .CD(n2462), .Q(out1_2[58]), 
        .QN(n1540) );
  CFD2XL \out1_2_reg[57]  ( .D(n431), .CP(clk), .CD(n2462), .Q(out1_2[57]), 
        .QN(n1544) );
  CFD2XL \out1_2_reg[56]  ( .D(n433), .CP(clk), .CD(n2462), .Q(out1_2[56]), 
        .QN(n1548) );
  CFD2XL \out1_2_reg[55]  ( .D(n435), .CP(clk), .CD(n2462), .Q(out1_2[55]), 
        .QN(n1552) );
  CFD2XL \out1_2_reg[54]  ( .D(n437), .CP(clk), .CD(n2462), .Q(out1_2[54]), 
        .QN(n1556) );
  CFD2XL \out1_2_reg[53]  ( .D(n439), .CP(clk), .CD(n2462), .Q(out1_2[53]), 
        .QN(n1560) );
  CFD2XL \out1_2_reg[52]  ( .D(n441), .CP(clk), .CD(n2462), .Q(out1_2[52]), 
        .QN(n1564) );
  CFD2XL \out1_2_reg[51]  ( .D(n443), .CP(clk), .CD(n2462), .Q(out1_2[51]), 
        .QN(n1568) );
  CFD2XL \out1_2_reg[50]  ( .D(n445), .CP(clk), .CD(n2462), .Q(out1_2[50]), 
        .QN(n1572) );
  CFD2XL \out1_2_reg[49]  ( .D(n447), .CP(clk), .CD(n2462), .Q(out1_2[49]), 
        .QN(n1576) );
  CFD2XL \out1_2_reg[48]  ( .D(n449), .CP(clk), .CD(n2462), .Q(out1_2[48]), 
        .QN(n1580) );
  CFD2XL \out1_2_reg[47]  ( .D(n451), .CP(clk), .CD(n2462), .Q(out1_2[47]), 
        .QN(n1584) );
  CFD2XL \out1_2_reg[46]  ( .D(n453), .CP(clk), .CD(n2462), .Q(out1_2[46]), 
        .QN(n1588) );
  CFD2XL \out1_2_reg[45]  ( .D(n455), .CP(clk), .CD(n2462), .Q(out1_2[45]), 
        .QN(n1592) );
  CFD2XL \out1_2_reg[44]  ( .D(n457), .CP(clk), .CD(n2462), .Q(out1_2[44]), 
        .QN(n1596) );
  CFD2XL \out1_2_reg[43]  ( .D(n459), .CP(clk), .CD(n2462), .Q(out1_2[43]), 
        .QN(n1600) );
  CFD2XL \out1_2_reg[42]  ( .D(n461), .CP(clk), .CD(n2462), .Q(out1_2[42]), 
        .QN(n1604) );
  CFD2XL \out1_2_reg[41]  ( .D(n463), .CP(clk), .CD(n2462), .Q(out1_2[41]), 
        .QN(n1608) );
  CFD2XL \out1_2_reg[40]  ( .D(n465), .CP(clk), .CD(n2462), .Q(out1_2[40]), 
        .QN(n1612) );
  CFD2XL \out1_2_reg[39]  ( .D(n467), .CP(clk), .CD(n2462), .Q(out1_2[39]), 
        .QN(n1616) );
  CFD2XL \out1_2_reg[38]  ( .D(n469), .CP(clk), .CD(n2462), .Q(out1_2[38]), 
        .QN(n1620) );
  CFD2XL \out1_2_reg[37]  ( .D(n471), .CP(clk), .CD(n2462), .Q(out1_2[37]), 
        .QN(n1624) );
  CFD2XL \out1_2_reg[36]  ( .D(n473), .CP(clk), .CD(n2462), .Q(out1_2[36]), 
        .QN(n1628) );
  CFD2XL \out1_2_reg[35]  ( .D(n475), .CP(clk), .CD(n2462), .Q(out1_2[35]), 
        .QN(n1632) );
  CFD2XL \out1_2_reg[34]  ( .D(n477), .CP(clk), .CD(n2462), .Q(out1_2[34]), 
        .QN(n1636) );
  CFD2XL \out1_2_reg[33]  ( .D(n479), .CP(clk), .CD(n2462), .Q(out1_2[33]), 
        .QN(n1640) );
  CFD2XL \out2_2_reg[4]  ( .D(n1224), .CP(clk), .CD(n2462), .Q(out2_2[4]), 
        .QN(n2358) );
  CFD2XL \out1_2_reg[31]  ( .D(n483), .CP(clk), .CD(n2462), .Q(out1_2[31]), 
        .QN(n1648) );
  CFD2XL \out1_2_reg[30]  ( .D(n485), .CP(clk), .CD(n2462), .Q(out1_2[30]), 
        .QN(n1652) );
  CFD2XL \out1_2_reg[29]  ( .D(n487), .CP(clk), .CD(n2462), .Q(out1_2[29]), 
        .QN(n1656) );
  CFD2XL \out1_2_reg[28]  ( .D(n489), .CP(clk), .CD(n2462), .Q(out1_2[28]), 
        .QN(n1660) );
  CFD2XL \out1_2_reg[27]  ( .D(n491), .CP(clk), .CD(n2462), .Q(out1_2[27]), 
        .QN(n1664) );
  CFD2XL \out1_2_reg[26]  ( .D(n493), .CP(clk), .CD(n2462), .Q(out1_2[26]), 
        .QN(n1668) );
  CFD2XL \out1_2_reg[25]  ( .D(n495), .CP(clk), .CD(n2462), .Q(out1_2[25]), 
        .QN(n1672) );
  CFD2XL \out1_2_reg[24]  ( .D(n497), .CP(clk), .CD(n2462), .Q(out1_2[24]), 
        .QN(n1676) );
  CFD2XL \out1_2_reg[23]  ( .D(n499), .CP(clk), .CD(n2462), .Q(out1_2[23]), 
        .QN(n1680) );
  CFD2XL \out1_2_reg[22]  ( .D(n501), .CP(clk), .CD(n2462), .Q(out1_2[22]), 
        .QN(n1684) );
  CFD1XL roundit_reg ( .D(n1217), .CP(clk), .Q(roundit), .QN(n2455) );
  CFD2X1 push0_2_reg ( .D(n1219), .CP(clk), .CD(n2462), .Q(push0_2), .QN(n2461) );
  CFD1X1 cmd1_en_2_reg ( .D(n756), .CP(clk), .Q(cmd1_en_2), .QN(n1395) );
  CFD2QX1 \q0_reg[4]  ( .D(n1181), .CP(clk), .CD(n1452), .Q(q0[4]) );
  CFD2QX1 \h0_reg[6]  ( .D(n632), .CP(clk), .CD(n1454), .Q(h0[6]) );
  CFD2QX1 \h0_reg[3]  ( .D(n623), .CP(clk), .CD(n1454), .Q(h0[3]) );
  CFD2QX1 \h0_reg[5]  ( .D(n629), .CP(clk), .CD(n1454), .Q(h0[5]) );
  CFD2QX1 \h0_reg[12]  ( .D(n1201), .CP(clk), .CD(n1453), .Q(h0[12]) );
  CFD2QX1 \q0_reg[6]  ( .D(n664), .CP(clk), .CD(n1452), .Q(q0[6]) );
  CFD2QX4 \q0_reg[26]  ( .D(n684), .CP(clk), .CD(n1450), .Q(q0[26]) );
  CFD2QX2 \q0_reg[14]  ( .D(n791), .CP(clk), .CD(n1451), .Q(q0[14]) );
  CDLY1XL U921 ( .A(q0[5]), .Z(n790) );
  CIVXL U922 ( .A(cmd1_en_2), .Z(n1400) );
  CNIVX1 U923 ( .A(n672), .Z(n791) );
  CNIVXL U924 ( .A(n1395), .Z(n792) );
  CDLY1XL U925 ( .A(q0[8]), .Z(n793) );
  CIVDXL U926 ( .A(cmd2_en_2), .Z0(n794), .Z1(n795) );
  CAN4X1 U927 ( .A(n2460), .B(push0_2), .C(n2459), .D(n2458), .Z(n796) );
  CMX2XL U928 ( .A0(q0[20]), .A1(q[20]), .S(n1496), .Z(n678) );
  CDLY1XL U929 ( .A(q0[24]), .Z(n797) );
  CNIVX1 U930 ( .A(_pushout_d), .Z(n798) );
  CNIVX1 U931 ( .A(n567), .Z(n799) );
  CNIVX1 U932 ( .A(n566), .Z(n800) );
  CNIVX1 U933 ( .A(n568), .Z(n801) );
  CNIVX1 U934 ( .A(n578), .Z(n802) );
  CNIVX1 U935 ( .A(n576), .Z(n803) );
  CNIVX1 U936 ( .A(n570), .Z(n804) );
  CNIVX1 U937 ( .A(n564), .Z(n805) );
  CNIVX1 U938 ( .A(n565), .Z(n806) );
  CNIVX1 U939 ( .A(n605), .Z(n807) );
  CNIVX1 U940 ( .A(n663), .Z(n808) );
  CIVXL U941 ( .A(out2_2[3]), .Z(n2375) );
  CNIVX1 U942 ( .A(n2375), .Z(n809) );
  CIVDX1 U943 ( .A(cmd0_1[1]), .Z1(n811) );
  CNIVX1 U944 ( .A(n811), .Z(n810) );
  CIVDX1 U945 ( .A(cmd0_1[0]), .Z1(n813) );
  CNIVX1 U946 ( .A(n813), .Z(n812) );
  CANR2XL U947 ( .A(out1_2[22]), .B(n1299), .C(acc[22]), .D(n2461), .Z(n1681)
         );
  CANR2XL U948 ( .A(out1_2[23]), .B(n1299), .C(acc[23]), .D(n2461), .Z(n1677)
         );
  CANR2XL U949 ( .A(out1_2[14]), .B(n1299), .C(acc[14]), .D(n2461), .Z(n1713)
         );
  CANR2XL U950 ( .A(out1_2[24]), .B(n1299), .C(acc[24]), .D(n2461), .Z(n1673)
         );
  CANR2XL U951 ( .A(out1_2[30]), .B(n1299), .C(acc[30]), .D(n2461), .Z(n1649)
         );
  CANR2XL U952 ( .A(out1_2[16]), .B(n1299), .C(acc[16]), .D(n2461), .Z(n1705)
         );
  CANR2XL U953 ( .A(out1_2[6]), .B(n1299), .C(acc[6]), .D(n2461), .Z(n1745) );
  CANR2XL U954 ( .A(out1_2[28]), .B(n1299), .C(acc[28]), .D(n2461), .Z(n1657)
         );
  CANR2XL U955 ( .A(out1_2[12]), .B(n1299), .C(acc[12]), .D(n2461), .Z(n1721)
         );
  CANR2XL U956 ( .A(out1_2[27]), .B(n1299), .C(acc[27]), .D(n2461), .Z(n1661)
         );
  CANR2XL U957 ( .A(out1_2[15]), .B(n1299), .C(acc[15]), .D(n2461), .Z(n1709)
         );
  CANR2XL U958 ( .A(out1_2[29]), .B(n1299), .C(acc[29]), .D(n2461), .Z(n1653)
         );
  CANR2XL U959 ( .A(out1_2[26]), .B(n1299), .C(acc[26]), .D(n2461), .Z(n1665)
         );
  CANR2XL U960 ( .A(out1_2[7]), .B(n1299), .C(acc[7]), .D(n2461), .Z(n1741) );
  CANR2XL U961 ( .A(out1_2[31]), .B(n1299), .C(acc[31]), .D(n2461), .Z(n1645)
         );
  CANR2XL U962 ( .A(out1_2[9]), .B(n1299), .C(acc[9]), .D(n2461), .Z(n1733) );
  CANR2XL U963 ( .A(out1_2[11]), .B(n1299), .C(acc[11]), .D(n2461), .Z(n1725)
         );
  CANR2XL U964 ( .A(out1_2[8]), .B(n1299), .C(acc[8]), .D(n2461), .Z(n1737) );
  CANR2XL U965 ( .A(out1_2[10]), .B(n1299), .C(acc[10]), .D(n2461), .Z(n1729)
         );
  CANR2XL U966 ( .A(out1_2[13]), .B(n1299), .C(acc[13]), .D(n2461), .Z(n1717)
         );
  CANR2XL U967 ( .A(out1_2[25]), .B(n1299), .C(acc[25]), .D(n2461), .Z(n1669)
         );
  CANR2XL U968 ( .A(out1_2[5]), .B(n1299), .C(acc[5]), .D(n2461), .Z(n1749) );
  CNIVX1 U969 ( .A(n650), .Z(n814) );
  CNIVX1 U970 ( .A(n708), .Z(n815) );
  CMX2XL U971 ( .A0(out0_2[46]), .A1(out0_1[46]), .S(n1383), .Z(n708) );
  CNIVX1 U972 ( .A(n732), .Z(n816) );
  CMX2XL U973 ( .A0(out0_2[22]), .A1(out0_1[22]), .S(n1368), .Z(n732) );
  CNIVX1 U974 ( .A(n731), .Z(n817) );
  CMX2XL U975 ( .A0(out0_2[23]), .A1(out0_1[23]), .S(n1368), .Z(n731) );
  CNIVX1 U976 ( .A(n718), .Z(n818) );
  CMX2XL U977 ( .A0(out0_2[36]), .A1(out0_1[36]), .S(n1393), .Z(n718) );
  CNIVX1 U978 ( .A(n734), .Z(n819) );
  CMX2XL U979 ( .A0(out0_2[20]), .A1(out0_1[20]), .S(n1368), .Z(n734) );
  CNIVX1 U980 ( .A(n706), .Z(n820) );
  CMX2XL U981 ( .A0(out0_2[48]), .A1(out0_1[48]), .S(n1381), .Z(n706) );
  CNIVX1 U982 ( .A(n716), .Z(n821) );
  CMX2XL U983 ( .A0(out0_2[38]), .A1(out0_1[38]), .S(n1391), .Z(n716) );
  CNIVX1 U984 ( .A(n700), .Z(n822) );
  CMX2XL U985 ( .A0(out0_2[54]), .A1(out0_1[54]), .S(n1375), .Z(n700) );
  CNIVX1 U986 ( .A(n736), .Z(n823) );
  CMX2XL U987 ( .A0(out0_2[18]), .A1(out0_1[18]), .S(n1370), .Z(n736) );
  CNIVX1 U988 ( .A(n707), .Z(n824) );
  CMX2XL U989 ( .A0(out0_2[47]), .A1(out0_1[47]), .S(n1382), .Z(n707) );
  CNIVX1 U990 ( .A(n702), .Z(n825) );
  CMX2XL U991 ( .A0(out0_2[52]), .A1(out0_1[52]), .S(n1377), .Z(n702) );
  CNIVX1 U992 ( .A(n740), .Z(n826) );
  CMX2XL U993 ( .A0(out0_2[14]), .A1(out0_1[14]), .S(n1374), .Z(n740) );
  CNIVX1 U994 ( .A(n705), .Z(n827) );
  CMX2XL U995 ( .A0(out0_2[49]), .A1(out0_1[49]), .S(n1380), .Z(n705) );
  CNIVX1 U996 ( .A(n730), .Z(n828) );
  CMX2XL U997 ( .A0(out0_2[24]), .A1(out0_1[24]), .S(n1368), .Z(n730) );
  CNIVX1 U998 ( .A(n724), .Z(n829) );
  CMX2XL U999 ( .A0(out0_2[30]), .A1(out0_1[30]), .S(n1390), .Z(n724) );
  CNIVX1 U1000 ( .A(n696), .Z(n830) );
  CMX2XL U1001 ( .A0(out0_2[58]), .A1(out0_1[58]), .S(n1371), .Z(n696) );
  CNIVX1 U1002 ( .A(n748), .Z(n831) );
  CMX2XL U1003 ( .A0(out0_2[6]), .A1(out0_1[6]), .S(n1382), .Z(n748) );
  CNIVX1 U1004 ( .A(n726), .Z(n832) );
  CNIVX1 U1005 ( .A(n710), .Z(n833) );
  CMX2XL U1006 ( .A0(out0_2[44]), .A1(out0_1[44]), .S(n1385), .Z(n710) );
  CNIVX1 U1007 ( .A(n742), .Z(n834) );
  CMX2XL U1008 ( .A0(out0_2[12]), .A1(out0_1[12]), .S(n1376), .Z(n742) );
  CNIVX1 U1009 ( .A(n701), .Z(n835) );
  CMX2XL U1010 ( .A0(out0_2[53]), .A1(out0_1[53]), .S(n1376), .Z(n701) );
  CNIVX1 U1011 ( .A(n733), .Z(n836) );
  CMX2XL U1012 ( .A0(out0_2[21]), .A1(out0_1[21]), .S(n1368), .Z(n733) );
  CNIVX1 U1013 ( .A(n704), .Z(n837) );
  CMX2XL U1014 ( .A0(out0_2[50]), .A1(out0_1[50]), .S(n1379), .Z(n704) );
  CNIVX1 U1015 ( .A(n703), .Z(n838) );
  CMX2XL U1016 ( .A0(out0_2[51]), .A1(out0_1[51]), .S(n1378), .Z(n703) );
  CNIVX1 U1017 ( .A(n717), .Z(n839) );
  CMX2XL U1018 ( .A0(out0_2[37]), .A1(out0_1[37]), .S(n1392), .Z(n717) );
  CNIVX1 U1019 ( .A(n725), .Z(n840) );
  CMX2XL U1020 ( .A0(out0_2[29]), .A1(out0_1[29]), .S(n1394), .Z(n725) );
  CNIVX1 U1021 ( .A(n728), .Z(n841) );
  CNIVX1 U1022 ( .A(n697), .Z(n842) );
  CMX2XL U1023 ( .A0(out0_2[57]), .A1(out0_1[57]), .S(n1372), .Z(n697) );
  CNIVX1 U1024 ( .A(n698), .Z(n843) );
  CMX2XL U1025 ( .A0(out0_2[56]), .A1(out0_1[56]), .S(n1373), .Z(n698) );
  CNIVX1 U1026 ( .A(n699), .Z(n844) );
  CMX2XL U1027 ( .A0(out0_2[55]), .A1(out0_1[55]), .S(n1374), .Z(n699) );
  CNIVX1 U1028 ( .A(n750), .Z(n845) );
  CMX2XL U1029 ( .A0(out0_2[4]), .A1(out0_1[4]), .S(n1384), .Z(n750) );
  CNIVX1 U1030 ( .A(n723), .Z(n846) );
  CMX2XL U1031 ( .A0(out0_2[31]), .A1(out0_1[31]), .S(n1388), .Z(n723) );
  CNIVX1 U1032 ( .A(n752), .Z(n847) );
  CMX2XL U1033 ( .A0(out0_2[2]), .A1(out0_1[2]), .S(n1386), .Z(n752) );
  CNIVX1 U1034 ( .A(n695), .Z(n848) );
  CMX2XL U1035 ( .A0(out0_2[59]), .A1(out0_1[59]), .S(n1370), .Z(n695) );
  CNIVX1 U1036 ( .A(n745), .Z(n849) );
  CMX2XL U1037 ( .A0(out0_2[9]), .A1(out0_1[9]), .S(n1379), .Z(n745) );
  CNIVX1 U1038 ( .A(n721), .Z(n850) );
  CMX2XL U1039 ( .A0(out0_2[33]), .A1(out0_1[33]), .S(n1393), .Z(n721) );
  CNIVX1 U1040 ( .A(n743), .Z(n851) );
  CMX2XL U1041 ( .A0(out0_2[11]), .A1(out0_1[11]), .S(n1377), .Z(n743) );
  CNIVX1 U1042 ( .A(n719), .Z(n852) );
  CMX2XL U1043 ( .A0(out0_2[35]), .A1(out0_1[35]), .S(n1391), .Z(n719) );
  CNIVX1 U1044 ( .A(n713), .Z(n853) );
  CMX2XL U1045 ( .A0(out0_2[41]), .A1(out0_1[41]), .S(n1388), .Z(n713) );
  CNIVX1 U1046 ( .A(n711), .Z(n854) );
  CMX2XL U1047 ( .A0(out0_2[43]), .A1(out0_1[43]), .S(n1386), .Z(n711) );
  CNIVX1 U1048 ( .A(n737), .Z(n855) );
  CMX2XL U1049 ( .A0(out0_2[17]), .A1(out0_1[17]), .S(n1371), .Z(n737) );
  CNIVX1 U1050 ( .A(n722), .Z(n856) );
  CMX2XL U1051 ( .A0(out0_2[32]), .A1(out0_1[32]), .S(n1394), .Z(n722) );
  CNIVX1 U1052 ( .A(n651), .Z(n857) );
  CNIVX1 U1053 ( .A(n751), .Z(n858) );
  CMX2XL U1054 ( .A0(out0_2[3]), .A1(out0_1[3]), .S(n1385), .Z(n751) );
  CNIVX1 U1055 ( .A(n744), .Z(n859) );
  CMX2XL U1056 ( .A0(out0_2[10]), .A1(out0_1[10]), .S(n1378), .Z(n744) );
  CNIVX1 U1057 ( .A(n735), .Z(n860) );
  CMX2XL U1058 ( .A0(out0_2[19]), .A1(out0_1[19]), .S(n1369), .Z(n735) );
  CNIVX1 U1059 ( .A(n720), .Z(n861) );
  CMX2XL U1060 ( .A0(out0_2[34]), .A1(out0_1[34]), .S(n1392), .Z(n720) );
  CNIVX1 U1061 ( .A(n741), .Z(n862) );
  CMX2XL U1062 ( .A0(out0_2[13]), .A1(out0_1[13]), .S(n1375), .Z(n741) );
  CNIVX1 U1063 ( .A(n729), .Z(n863) );
  CNIVX1 U1064 ( .A(n749), .Z(n864) );
  CMX2XL U1065 ( .A0(out0_2[5]), .A1(out0_1[5]), .S(n1383), .Z(n749) );
  CNIVX1 U1066 ( .A(n754), .Z(n865) );
  CMX2XL U1067 ( .A0(out0_2[0]), .A1(out0_1[0]), .S(n1368), .Z(n754) );
  CNIVX1 U1068 ( .A(n714), .Z(n866) );
  CMX2XL U1069 ( .A0(out0_2[40]), .A1(out0_1[40]), .S(n1389), .Z(n714) );
  CNIVX1 U1070 ( .A(n727), .Z(n867) );
  CNIVX1 U1071 ( .A(n712), .Z(n868) );
  CMX2XL U1072 ( .A0(out0_2[42]), .A1(out0_1[42]), .S(n1387), .Z(n712) );
  CNIVX1 U1073 ( .A(n739), .Z(n869) );
  CMX2XL U1074 ( .A0(out0_2[15]), .A1(out0_1[15]), .S(n1373), .Z(n739) );
  CNIVX1 U1075 ( .A(n747), .Z(n870) );
  CMX2XL U1076 ( .A0(out0_2[7]), .A1(out0_1[7]), .S(n1381), .Z(n747) );
  CNIVX1 U1077 ( .A(n709), .Z(n871) );
  CMX2XL U1078 ( .A0(out0_2[45]), .A1(out0_1[45]), .S(n1384), .Z(n709) );
  CNIVX1 U1079 ( .A(n689), .Z(n872) );
  CNIVX1 U1080 ( .A(n715), .Z(n873) );
  CMX2XL U1081 ( .A0(out0_2[39]), .A1(out0_1[39]), .S(n1390), .Z(n715) );
  CMX2X2 U1082 ( .A0(out0_2[63]), .A1(out0_1[63]), .S(n1368), .Z(n691) );
  CMX2X2 U1083 ( .A0(out0_2[62]), .A1(out0_1[62]), .S(n1368), .Z(n692) );
  CMX2X2 U1084 ( .A0(out0_2[61]), .A1(out0_1[61]), .S(n1368), .Z(n693) );
  CMX2X2 U1085 ( .A0(out0_2[60]), .A1(out0_1[60]), .S(n1369), .Z(n694) );
  CIVDX1 U1086 ( .A(out1_0[0]), .Z1(n875) );
  CNIVX1 U1087 ( .A(n875), .Z(n874) );
  CIVDX1 U1088 ( .A(out1_0[1]), .Z1(n877) );
  CNIVX1 U1089 ( .A(n877), .Z(n876) );
  CIVDX1 U1090 ( .A(out1_0[2]), .Z1(n879) );
  CNIVX1 U1091 ( .A(n879), .Z(n878) );
  CIVDX1 U1092 ( .A(out1_0[3]), .Z1(n881) );
  CNIVX1 U1093 ( .A(n881), .Z(n880) );
  CIVDX1 U1094 ( .A(out1_0[4]), .Z1(n883) );
  CNIVX1 U1095 ( .A(n883), .Z(n882) );
  CIVDX1 U1096 ( .A(out1_0[5]), .Z1(n885) );
  CNIVX1 U1097 ( .A(n885), .Z(n884) );
  CIVDX1 U1098 ( .A(out1_0[6]), .Z1(n887) );
  CNIVX1 U1099 ( .A(n887), .Z(n886) );
  CIVDX1 U1100 ( .A(out1_0[7]), .Z1(n889) );
  CNIVX1 U1101 ( .A(n889), .Z(n888) );
  CIVDX1 U1102 ( .A(out1_0[8]), .Z1(n891) );
  CNIVX1 U1103 ( .A(n891), .Z(n890) );
  CIVDX1 U1104 ( .A(out1_0[9]), .Z1(n893) );
  CNIVX1 U1105 ( .A(n893), .Z(n892) );
  CIVDX1 U1106 ( .A(out1_0[10]), .Z1(n895) );
  CNIVX1 U1107 ( .A(n895), .Z(n894) );
  CIVDX1 U1108 ( .A(out1_0[11]), .Z1(n897) );
  CNIVX1 U1109 ( .A(n897), .Z(n896) );
  CIVDX1 U1110 ( .A(out1_0[12]), .Z1(n899) );
  CNIVX1 U1111 ( .A(n899), .Z(n898) );
  CIVDX1 U1112 ( .A(out1_0[13]), .Z1(n901) );
  CNIVX1 U1113 ( .A(n901), .Z(n900) );
  CIVDX1 U1114 ( .A(out1_0[14]), .Z1(n903) );
  CNIVX1 U1115 ( .A(n903), .Z(n902) );
  CIVDX1 U1116 ( .A(out1_0[15]), .Z1(n905) );
  CNIVX1 U1117 ( .A(n905), .Z(n904) );
  CIVDX1 U1118 ( .A(out1_0[16]), .Z1(n907) );
  CNIVX1 U1119 ( .A(n907), .Z(n906) );
  CIVDX1 U1120 ( .A(out1_0[17]), .Z1(n909) );
  CNIVX1 U1121 ( .A(n909), .Z(n908) );
  CIVDX1 U1122 ( .A(out1_0[18]), .Z1(n911) );
  CNIVX1 U1123 ( .A(n911), .Z(n910) );
  CIVDX1 U1124 ( .A(out1_0[19]), .Z1(n913) );
  CNIVX1 U1125 ( .A(n913), .Z(n912) );
  CIVDX1 U1126 ( .A(out1_0[20]), .Z1(n915) );
  CNIVX1 U1127 ( .A(n915), .Z(n914) );
  CIVDX1 U1128 ( .A(out1_0[21]), .Z1(n917) );
  CNIVX1 U1129 ( .A(n917), .Z(n916) );
  CIVDX1 U1130 ( .A(out1_0[22]), .Z1(n919) );
  CNIVX1 U1131 ( .A(n919), .Z(n918) );
  CIVDX1 U1132 ( .A(out1_0[23]), .Z1(n921) );
  CNIVX1 U1133 ( .A(n921), .Z(n920) );
  CIVDX1 U1134 ( .A(out1_0[24]), .Z1(n923) );
  CNIVX1 U1135 ( .A(n923), .Z(n922) );
  CIVDX1 U1136 ( .A(out1_0[25]), .Z1(n925) );
  CNIVX1 U1137 ( .A(n925), .Z(n924) );
  CIVDX1 U1138 ( .A(out1_0[26]), .Z1(n927) );
  CNIVX1 U1139 ( .A(n927), .Z(n926) );
  CIVDX1 U1140 ( .A(out1_0[27]), .Z1(n929) );
  CNIVX1 U1141 ( .A(n929), .Z(n928) );
  CIVDX1 U1142 ( .A(out1_0[28]), .Z1(n931) );
  CNIVX1 U1143 ( .A(n931), .Z(n930) );
  CIVDX1 U1144 ( .A(out1_0[29]), .Z1(n933) );
  CNIVX1 U1145 ( .A(n933), .Z(n932) );
  CIVDX1 U1146 ( .A(out1_0[30]), .Z1(n935) );
  CNIVX1 U1147 ( .A(n935), .Z(n934) );
  CIVDX1 U1148 ( .A(out1_0[31]), .Z1(n937) );
  CNIVX1 U1149 ( .A(n937), .Z(n936) );
  CIVDX1 U1150 ( .A(out1_0[32]), .Z1(n939) );
  CNIVX1 U1151 ( .A(n939), .Z(n938) );
  CIVDX1 U1152 ( .A(out1_0[33]), .Z1(n941) );
  CNIVX1 U1153 ( .A(n941), .Z(n940) );
  CIVDX1 U1154 ( .A(out1_0[34]), .Z1(n943) );
  CNIVX1 U1155 ( .A(n943), .Z(n942) );
  CIVDX1 U1156 ( .A(out1_0[35]), .Z1(n945) );
  CNIVX1 U1157 ( .A(n945), .Z(n944) );
  CIVDX1 U1158 ( .A(out1_0[36]), .Z1(n947) );
  CNIVX1 U1159 ( .A(n947), .Z(n946) );
  CIVDX1 U1160 ( .A(out1_0[37]), .Z1(n949) );
  CNIVX1 U1161 ( .A(n949), .Z(n948) );
  CIVDX1 U1162 ( .A(out1_0[38]), .Z1(n951) );
  CNIVX1 U1163 ( .A(n951), .Z(n950) );
  CIVDX1 U1164 ( .A(out1_0[39]), .Z1(n953) );
  CNIVX1 U1165 ( .A(n953), .Z(n952) );
  CIVDX1 U1166 ( .A(out1_0[40]), .Z1(n955) );
  CNIVX1 U1167 ( .A(n955), .Z(n954) );
  CIVDX1 U1168 ( .A(out1_0[42]), .Z1(n957) );
  CNIVX1 U1169 ( .A(n957), .Z(n956) );
  CIVDX1 U1170 ( .A(out1_0[43]), .Z1(n959) );
  CNIVX1 U1171 ( .A(n959), .Z(n958) );
  CIVDX1 U1172 ( .A(out1_0[44]), .Z1(n961) );
  CNIVX1 U1173 ( .A(n961), .Z(n960) );
  CIVDX1 U1174 ( .A(out1_0[45]), .Z1(n963) );
  CNIVX1 U1175 ( .A(n963), .Z(n962) );
  CIVDX1 U1176 ( .A(out1_0[46]), .Z1(n965) );
  CNIVX1 U1177 ( .A(n965), .Z(n964) );
  CIVDX1 U1178 ( .A(out1_0[47]), .Z1(n967) );
  CNIVX1 U1179 ( .A(n967), .Z(n966) );
  CIVDX1 U1180 ( .A(out1_0[48]), .Z1(n969) );
  CNIVX1 U1181 ( .A(n969), .Z(n968) );
  CIVDX1 U1182 ( .A(out1_0[49]), .Z1(n971) );
  CNIVX1 U1183 ( .A(n971), .Z(n970) );
  CIVDX1 U1184 ( .A(out1_0[50]), .Z1(n973) );
  CNIVX1 U1185 ( .A(n973), .Z(n972) );
  CIVDX1 U1186 ( .A(out1_0[51]), .Z1(n975) );
  CNIVX1 U1187 ( .A(n975), .Z(n974) );
  CIVDX1 U1188 ( .A(out1_0[52]), .Z1(n977) );
  CNIVX1 U1189 ( .A(n977), .Z(n976) );
  CIVDX1 U1190 ( .A(out1_0[53]), .Z1(n979) );
  CNIVX1 U1191 ( .A(n979), .Z(n978) );
  CIVDX1 U1192 ( .A(out1_0[54]), .Z1(n981) );
  CNIVX1 U1193 ( .A(n981), .Z(n980) );
  CIVDX1 U1194 ( .A(out1_0[55]), .Z1(n983) );
  CNIVX1 U1195 ( .A(n983), .Z(n982) );
  CIVDX1 U1196 ( .A(out1_0[56]), .Z1(n985) );
  CNIVX1 U1197 ( .A(n985), .Z(n984) );
  CIVDX1 U1198 ( .A(out1_0[57]), .Z1(n987) );
  CNIVX1 U1199 ( .A(n987), .Z(n986) );
  CIVDX1 U1200 ( .A(out1_0[58]), .Z1(n989) );
  CNIVX1 U1201 ( .A(n989), .Z(n988) );
  CIVDX1 U1202 ( .A(out1_0[59]), .Z1(n991) );
  CNIVX1 U1203 ( .A(n991), .Z(n990) );
  CIVDX1 U1204 ( .A(out1_0[60]), .Z1(n993) );
  CNIVX1 U1205 ( .A(n993), .Z(n992) );
  CIVDX1 U1206 ( .A(out1_0[61]), .Z1(n995) );
  CNIVX1 U1207 ( .A(n995), .Z(n994) );
  CIVDX1 U1208 ( .A(out1_0[62]), .Z1(n997) );
  CNIVX1 U1209 ( .A(n997), .Z(n996) );
  CANR2XL U1210 ( .A(out1_2[46]), .B(n1299), .C(acc[46]), .D(n2461), .Z(n1585)
         );
  CANR2XL U1211 ( .A(out1_2[34]), .B(n1299), .C(acc[34]), .D(n2461), .Z(n1633)
         );
  CANR2XL U1212 ( .A(out1_2[36]), .B(n1299), .C(acc[36]), .D(n2461), .Z(n1625)
         );
  CANR2XL U1213 ( .A(out1_2[40]), .B(n1299), .C(acc[40]), .D(n2461), .Z(n1609)
         );
  CANR2XL U1214 ( .A(out1_2[48]), .B(n1299), .C(acc[48]), .D(n2461), .Z(n1577)
         );
  CANR2XL U1215 ( .A(out1_2[38]), .B(n1299), .C(acc[38]), .D(n2461), .Z(n1617)
         );
  CANR2XL U1216 ( .A(out1_2[45]), .B(n1299), .C(acc[45]), .D(n2461), .Z(n1589)
         );
  CANR2XL U1217 ( .A(out1_2[47]), .B(n1299), .C(acc[47]), .D(n2461), .Z(n1581)
         );
  CANR2XL U1218 ( .A(out1_2[39]), .B(n1299), .C(acc[39]), .D(n2461), .Z(n1613)
         );
  CANR2XL U1219 ( .A(out1_2[49]), .B(n1299), .C(acc[49]), .D(n2461), .Z(n1573)
         );
  CANR2XL U1220 ( .A(out1_2[42]), .B(n1299), .C(acc[42]), .D(n2461), .Z(n1601)
         );
  CANR2XL U1221 ( .A(out1_2[44]), .B(n1299), .C(acc[44]), .D(n2461), .Z(n1593)
         );
  CANR2XL U1222 ( .A(out1_2[53]), .B(n1299), .C(acc[53]), .D(n2461), .Z(n1557)
         );
  CANR2XL U1223 ( .A(out1_2[50]), .B(n1299), .C(acc[50]), .D(n2461), .Z(n1569)
         );
  CANR2XL U1224 ( .A(out1_2[51]), .B(n1299), .C(acc[51]), .D(n2461), .Z(n1565)
         );
  CANR2XL U1225 ( .A(out1_2[37]), .B(n1299), .C(acc[37]), .D(n2461), .Z(n1621)
         );
  CANR2XL U1226 ( .A(out1_2[57]), .B(n1299), .C(acc[57]), .D(n2461), .Z(n1541)
         );
  CANR2XL U1227 ( .A(out1_2[56]), .B(n1299), .C(acc[56]), .D(n2461), .Z(n1545)
         );
  CANR2XL U1228 ( .A(out1_2[55]), .B(n1299), .C(acc[55]), .D(n2461), .Z(n1549)
         );
  CANR2XL U1229 ( .A(out1_2[59]), .B(n1299), .C(acc[59]), .D(n2461), .Z(n1533)
         );
  CANR2XL U1230 ( .A(out1_2[33]), .B(n1299), .C(acc[33]), .D(n2461), .Z(n1637)
         );
  CANR2XL U1231 ( .A(out1_2[35]), .B(n1299), .C(acc[35]), .D(n2461), .Z(n1629)
         );
  CANR2XL U1232 ( .A(out1_2[41]), .B(n1299), .C(acc[41]), .D(n2461), .Z(n1605)
         );
  CANR2XL U1233 ( .A(out1_2[43]), .B(n1299), .C(acc[43]), .D(n2461), .Z(n1597)
         );
  CANR2XL U1234 ( .A(out1_2[32]), .B(n1299), .C(acc[32]), .D(n2461), .Z(n1641)
         );
  CND2X2 U1235 ( .A(n1522), .B(n1521), .Z(n420) );
  CANR2XL U1236 ( .A(out1_2[61]), .B(n1299), .C(acc[61]), .D(n2461), .Z(n1525)
         );
  CANR2XL U1237 ( .A(out1_2[60]), .B(n1299), .C(acc[60]), .D(n2461), .Z(n1529)
         );
  CANR2XL U1238 ( .A(out1_2[58]), .B(n1299), .C(acc[58]), .D(n2461), .Z(n1537)
         );
  CANR2XL U1239 ( .A(out1_2[54]), .B(n1299), .C(acc[54]), .D(n2461), .Z(n1553)
         );
  CANR2XL U1240 ( .A(out1_2[52]), .B(n1299), .C(acc[52]), .D(n2461), .Z(n1561)
         );
  CNIVX1 U1241 ( .A(n637), .Z(n998) );
  CIVXL U1242 ( .A(h0_1[5]), .Z(n2426) );
  CIVXL U1243 ( .A(h0_1[6]), .Z(n2033) );
  CIVX3 U1244 ( .A(out2_2[63]), .Z(n1781) );
  CIVDX1 U1245 ( .A(out1_0[63]), .Z1(n1000) );
  CNIVX1 U1246 ( .A(n1000), .Z(n999) );
  CNIVX1 U1247 ( .A(n548), .Z(n1001) );
  CNIVX1 U1248 ( .A(n758), .Z(n1002) );
  CNIVX1 U1249 ( .A(n759), .Z(n1003) );
  CNIVX1 U1250 ( .A(n760), .Z(n1004) );
  CNIVX1 U1251 ( .A(n761), .Z(n1005) );
  CNIVX1 U1252 ( .A(n762), .Z(n1006) );
  CNIVX1 U1253 ( .A(n763), .Z(n1007) );
  CNIVX1 U1254 ( .A(n764), .Z(n1008) );
  CNIVX1 U1255 ( .A(n765), .Z(n1009) );
  CNIVX1 U1256 ( .A(n766), .Z(n1010) );
  CNIVX1 U1257 ( .A(n767), .Z(n1011) );
  CNIVX1 U1258 ( .A(n768), .Z(n1012) );
  CNIVX1 U1259 ( .A(n769), .Z(n1013) );
  CNIVX1 U1260 ( .A(n770), .Z(n1014) );
  CNIVX1 U1261 ( .A(n771), .Z(n1015) );
  CNIVX1 U1262 ( .A(n772), .Z(n1016) );
  CNIVX1 U1263 ( .A(n773), .Z(n1017) );
  CNIVX1 U1264 ( .A(n774), .Z(n1018) );
  CNIVX1 U1265 ( .A(n775), .Z(n1019) );
  CNIVX1 U1266 ( .A(n776), .Z(n1020) );
  CNIVX1 U1267 ( .A(n777), .Z(n1021) );
  CMX2X2 U1268 ( .A0(z[20]), .A1(acc[20]), .S(n796), .Z(n778) );
  CNIVX1 U1269 ( .A(n779), .Z(n1022) );
  CMX2X2 U1270 ( .A0(z[22]), .A1(acc[22]), .S(n796), .Z(n780) );
  CMX2X2 U1271 ( .A0(z[23]), .A1(acc[23]), .S(n796), .Z(n781) );
  CNIVX1 U1272 ( .A(n782), .Z(n1023) );
  CNIVX1 U1273 ( .A(n783), .Z(n1024) );
  CNIVX1 U1274 ( .A(n784), .Z(n1025) );
  CNIVX1 U1275 ( .A(n785), .Z(n1026) );
  CNIVX1 U1276 ( .A(n786), .Z(n1027) );
  CNIVX1 U1277 ( .A(n787), .Z(n1028) );
  CMX2X2 U1278 ( .A0(z[30]), .A1(acc[30]), .S(n796), .Z(n788) );
  CMX2X2 U1279 ( .A0(z[31]), .A1(acc[31]), .S(n796), .Z(n789) );
  CMXI2X2 U1280 ( .A0(n1489), .A1(n1511), .S(n215), .Z(n613) );
  CMXI2X2 U1281 ( .A0(n1776), .A1(n1777), .S(n215), .Z(n622) );
  CIVX4 U1282 ( .A(h0_0[4]), .Z(n1508) );
  CIVX4 U1283 ( .A(h0_0[5]), .Z(n1506) );
  CIVX4 U1284 ( .A(h0_0[6]), .Z(n1504) );
  CIVDX1 U1285 ( .A(out0_0[0]), .Z1(n1030) );
  CNIVX1 U1286 ( .A(n1030), .Z(n1029) );
  CIVDX1 U1287 ( .A(out0_0[1]), .Z1(n1032) );
  CNIVX1 U1288 ( .A(n1032), .Z(n1031) );
  CIVDX1 U1289 ( .A(out0_0[2]), .Z1(n1034) );
  CNIVX1 U1290 ( .A(n1034), .Z(n1033) );
  CIVDX1 U1291 ( .A(out0_0[3]), .Z1(n1036) );
  CNIVX1 U1292 ( .A(n1036), .Z(n1035) );
  CIVDX1 U1293 ( .A(out0_0[4]), .Z1(n1038) );
  CNIVX1 U1294 ( .A(n1038), .Z(n1037) );
  CIVDX1 U1295 ( .A(out0_0[5]), .Z1(n1040) );
  CNIVX1 U1296 ( .A(n1040), .Z(n1039) );
  CIVDX1 U1297 ( .A(out0_0[6]), .Z1(n1042) );
  CNIVX1 U1298 ( .A(n1042), .Z(n1041) );
  CIVDX1 U1299 ( .A(out0_0[7]), .Z1(n1044) );
  CNIVX1 U1300 ( .A(n1044), .Z(n1043) );
  CIVDX1 U1301 ( .A(out0_0[8]), .Z1(n1046) );
  CNIVX1 U1302 ( .A(n1046), .Z(n1045) );
  CIVDX1 U1303 ( .A(out0_0[9]), .Z1(n1048) );
  CNIVX1 U1304 ( .A(n1048), .Z(n1047) );
  CIVDX1 U1305 ( .A(out0_0[10]), .Z1(n1050) );
  CNIVX1 U1306 ( .A(n1050), .Z(n1049) );
  CIVDX1 U1307 ( .A(out0_0[11]), .Z1(n1052) );
  CNIVX1 U1308 ( .A(n1052), .Z(n1051) );
  CIVDX1 U1309 ( .A(out0_0[12]), .Z1(n1054) );
  CNIVX1 U1310 ( .A(n1054), .Z(n1053) );
  CIVDX1 U1311 ( .A(out0_0[13]), .Z1(n1056) );
  CNIVX1 U1312 ( .A(n1056), .Z(n1055) );
  CIVDX1 U1313 ( .A(out0_0[14]), .Z1(n1058) );
  CNIVX1 U1314 ( .A(n1058), .Z(n1057) );
  CIVDX1 U1315 ( .A(out0_0[15]), .Z1(n1060) );
  CNIVX1 U1316 ( .A(n1060), .Z(n1059) );
  CIVDX1 U1317 ( .A(out0_0[16]), .Z1(n1062) );
  CNIVX1 U1318 ( .A(n1062), .Z(n1061) );
  CIVDX1 U1319 ( .A(out0_0[17]), .Z1(n1064) );
  CNIVX1 U1320 ( .A(n1064), .Z(n1063) );
  CIVDX1 U1321 ( .A(out0_0[18]), .Z1(n1066) );
  CNIVX1 U1322 ( .A(n1066), .Z(n1065) );
  CIVDX1 U1323 ( .A(out0_0[19]), .Z1(n1068) );
  CNIVX1 U1324 ( .A(n1068), .Z(n1067) );
  CIVDX1 U1325 ( .A(out0_0[20]), .Z1(n1070) );
  CNIVX1 U1326 ( .A(n1070), .Z(n1069) );
  CIVDX1 U1327 ( .A(out0_0[21]), .Z1(n1072) );
  CNIVX1 U1328 ( .A(n1072), .Z(n1071) );
  CIVDX1 U1329 ( .A(out0_0[22]), .Z1(n1074) );
  CNIVX1 U1330 ( .A(n1074), .Z(n1073) );
  CIVDX1 U1331 ( .A(out0_0[23]), .Z1(n1076) );
  CNIVX1 U1332 ( .A(n1076), .Z(n1075) );
  CIVDX1 U1333 ( .A(out0_0[24]), .Z1(n1078) );
  CNIVX1 U1334 ( .A(n1078), .Z(n1077) );
  CIVDX1 U1335 ( .A(out0_0[25]), .Z1(n1080) );
  CNIVX1 U1336 ( .A(n1080), .Z(n1079) );
  CIVDX1 U1337 ( .A(out0_0[26]), .Z1(n1082) );
  CNIVX1 U1338 ( .A(n1082), .Z(n1081) );
  CIVDX1 U1339 ( .A(out0_0[27]), .Z1(n1084) );
  CNIVX1 U1340 ( .A(n1084), .Z(n1083) );
  CIVDX1 U1341 ( .A(out0_0[28]), .Z1(n1086) );
  CNIVX1 U1342 ( .A(n1086), .Z(n1085) );
  CIVDX1 U1343 ( .A(out0_0[29]), .Z1(n1088) );
  CNIVX1 U1344 ( .A(n1088), .Z(n1087) );
  CIVDX1 U1345 ( .A(out0_0[30]), .Z1(n1090) );
  CNIVX1 U1346 ( .A(n1090), .Z(n1089) );
  CIVDX1 U1347 ( .A(out0_0[31]), .Z1(n1092) );
  CNIVX1 U1348 ( .A(n1092), .Z(n1091) );
  CIVDX1 U1349 ( .A(out0_0[32]), .Z1(n1094) );
  CNIVX1 U1350 ( .A(n1094), .Z(n1093) );
  CIVDX1 U1351 ( .A(out0_0[33]), .Z1(n1096) );
  CNIVX1 U1352 ( .A(n1096), .Z(n1095) );
  CIVDX1 U1353 ( .A(out0_0[34]), .Z1(n1098) );
  CNIVX1 U1354 ( .A(n1098), .Z(n1097) );
  CIVDX1 U1355 ( .A(out0_0[35]), .Z1(n1100) );
  CNIVX1 U1356 ( .A(n1100), .Z(n1099) );
  CIVDX1 U1357 ( .A(out0_0[36]), .Z1(n1102) );
  CNIVX1 U1358 ( .A(n1102), .Z(n1101) );
  CIVDX1 U1359 ( .A(out0_0[37]), .Z1(n1104) );
  CNIVX1 U1360 ( .A(n1104), .Z(n1103) );
  CIVDX1 U1361 ( .A(out0_0[38]), .Z1(n1106) );
  CNIVX1 U1362 ( .A(n1106), .Z(n1105) );
  CIVDX1 U1363 ( .A(out0_0[39]), .Z1(n1108) );
  CNIVX1 U1364 ( .A(n1108), .Z(n1107) );
  CIVDX1 U1365 ( .A(out0_0[40]), .Z1(n1110) );
  CNIVX1 U1366 ( .A(n1110), .Z(n1109) );
  CIVDX1 U1367 ( .A(out0_0[41]), .Z1(n1112) );
  CNIVX1 U1368 ( .A(n1112), .Z(n1111) );
  CIVDX1 U1369 ( .A(out0_0[42]), .Z1(n1114) );
  CNIVX1 U1370 ( .A(n1114), .Z(n1113) );
  CIVDX1 U1371 ( .A(out0_0[43]), .Z1(n1116) );
  CNIVX1 U1372 ( .A(n1116), .Z(n1115) );
  CIVDX1 U1373 ( .A(out0_0[44]), .Z1(n1118) );
  CNIVX1 U1374 ( .A(n1118), .Z(n1117) );
  CIVDX1 U1375 ( .A(out0_0[45]), .Z1(n1120) );
  CNIVX1 U1376 ( .A(n1120), .Z(n1119) );
  CIVDX1 U1377 ( .A(out0_0[46]), .Z1(n1122) );
  CNIVX1 U1378 ( .A(n1122), .Z(n1121) );
  CIVDX1 U1379 ( .A(out0_0[47]), .Z1(n1124) );
  CNIVX1 U1380 ( .A(n1124), .Z(n1123) );
  CIVDX1 U1381 ( .A(out0_0[48]), .Z1(n1126) );
  CNIVX1 U1382 ( .A(n1126), .Z(n1125) );
  CIVDX1 U1383 ( .A(out0_0[49]), .Z1(n1128) );
  CNIVX1 U1384 ( .A(n1128), .Z(n1127) );
  CIVDX1 U1385 ( .A(out0_0[50]), .Z1(n1130) );
  CNIVX1 U1386 ( .A(n1130), .Z(n1129) );
  CIVDX1 U1387 ( .A(out0_0[51]), .Z1(n1132) );
  CNIVX1 U1388 ( .A(n1132), .Z(n1131) );
  CIVDX1 U1389 ( .A(out0_0[52]), .Z1(n1134) );
  CNIVX1 U1390 ( .A(n1134), .Z(n1133) );
  CIVDX1 U1391 ( .A(out0_0[53]), .Z1(n1136) );
  CNIVX1 U1392 ( .A(n1136), .Z(n1135) );
  CIVDX1 U1393 ( .A(out0_0[54]), .Z1(n1138) );
  CNIVX1 U1394 ( .A(n1138), .Z(n1137) );
  CIVDX1 U1395 ( .A(out0_0[55]), .Z1(n1140) );
  CNIVX1 U1396 ( .A(n1140), .Z(n1139) );
  CIVDX1 U1397 ( .A(out0_0[56]), .Z1(n1142) );
  CNIVX1 U1398 ( .A(n1142), .Z(n1141) );
  CIVDX1 U1399 ( .A(out0_0[57]), .Z1(n1144) );
  CNIVX1 U1400 ( .A(n1144), .Z(n1143) );
  CIVDX1 U1401 ( .A(out0_0[58]), .Z1(n1146) );
  CNIVX1 U1402 ( .A(n1146), .Z(n1145) );
  CIVDX1 U1403 ( .A(out0_0[59]), .Z1(n1148) );
  CNIVX1 U1404 ( .A(n1148), .Z(n1147) );
  CIVDX1 U1405 ( .A(out0_0[60]), .Z1(n1150) );
  CNIVX1 U1406 ( .A(n1150), .Z(n1149) );
  CIVDX1 U1407 ( .A(out0_0[61]), .Z1(n1152) );
  CNIVX1 U1408 ( .A(n1152), .Z(n1151) );
  CIVDX1 U1409 ( .A(out0_0[62]), .Z1(n1154) );
  CNIVX1 U1410 ( .A(n1154), .Z(n1153) );
  CIVDX1 U1411 ( .A(out0_0[63]), .Z1(n1156) );
  CNIVX1 U1412 ( .A(n1156), .Z(n1155) );
  CIVDX1 U1413 ( .A(out1_0[41]), .Z1(n1158) );
  CNIVX1 U1414 ( .A(n1158), .Z(n1157) );
  CNIVX1 U1415 ( .A(n597), .Z(n1159) );
  CNIVX1 U1416 ( .A(n753), .Z(n1160) );
  CMX2XL U1417 ( .A0(out0_2[1]), .A1(out0_1[1]), .S(n1387), .Z(n753) );
  CNIVX1 U1418 ( .A(n554), .Z(n1161) );
  CNIVX1 U1419 ( .A(n551), .Z(n1162) );
  CNIVX1 U1420 ( .A(n678), .Z(n1163) );
  CNIVX1 U1421 ( .A(n553), .Z(n1164) );
  CNIVX1 U1422 ( .A(n555), .Z(n1165) );
  CNIVX1 U1423 ( .A(n556), .Z(n1166) );
  CNIVX1 U1424 ( .A(n559), .Z(n1167) );
  CNIVX1 U1425 ( .A(n562), .Z(n1168) );
  CNIVX1 U1426 ( .A(n1495), .Z(n1169) );
  CNIVX1 U1427 ( .A(n560), .Z(n1170) );
  CNIVX1 U1428 ( .A(n552), .Z(n1171) );
  CNIVX1 U1429 ( .A(n569), .Z(n1172) );
  CIVX4 U1430 ( .A(h0_0[2]), .Z(n1513) );
  CNIVX1 U1431 ( .A(n571), .Z(n1173) );
  CNIVX1 U1432 ( .A(n575), .Z(n1174) );
  CNIVX1 U1433 ( .A(n641), .Z(n1175) );
  CMX2XL U1434 ( .A0(h0[15]), .A1(h[15]), .S(n1500), .Z(n641) );
  CNIVX1 U1435 ( .A(n558), .Z(n1176) );
  CNIVX1 U1436 ( .A(n561), .Z(n1177) );
  CNIVX1 U1437 ( .A(n574), .Z(n1178) );
  CNIVX1 U1438 ( .A(n577), .Z(n1179) );
  CNIVX1 U1439 ( .A(n660), .Z(n1180) );
  CNIVX1 U1440 ( .A(n662), .Z(n1181) );
  CMX2XL U1441 ( .A0(q0[4]), .A1(q[4]), .S(n1498), .Z(n662) );
  CNIVX1 U1442 ( .A(n572), .Z(n1182) );
  CNIVX1 U1443 ( .A(n666), .Z(n1183) );
  CNIVX1 U1444 ( .A(n674), .Z(n1184) );
  CNIVX1 U1445 ( .A(n550), .Z(n1185) );
  CNIVX1 U1446 ( .A(n549), .Z(n1186) );
  CNIVX1 U1447 ( .A(n633), .Z(n1187) );
  CNIVX1 U1448 ( .A(n646), .Z(n1188) );
  CNIVX1 U1449 ( .A(n642), .Z(n1189) );
  CNIVX1 U1450 ( .A(n636), .Z(n1190) );
  CNIVX1 U1451 ( .A(n640), .Z(n1191) );
  CNIVX1 U1452 ( .A(n647), .Z(n1192) );
  CNIVX1 U1453 ( .A(n649), .Z(n1193) );
  CNIVX1 U1454 ( .A(n596), .Z(n1194) );
  CNIVX1 U1455 ( .A(n598), .Z(n1195) );
  CNIVX1 U1456 ( .A(n648), .Z(n1196) );
  CNIVX1 U1457 ( .A(n653), .Z(n1197) );
  CNIVX1 U1458 ( .A(n643), .Z(n1198) );
  CNIVX1 U1459 ( .A(n635), .Z(n1199) );
  CNIVX1 U1460 ( .A(n657), .Z(n1200) );
  CNIVX1 U1461 ( .A(n638), .Z(n1201) );
  CMX2XL U1462 ( .A0(h0[12]), .A1(h[12]), .S(n1500), .Z(n638) );
  CNIVX1 U1463 ( .A(n644), .Z(n1202) );
  CMX2XL U1464 ( .A0(h0[18]), .A1(h[18]), .S(n1499), .Z(n644) );
  CNIVX1 U1465 ( .A(h0[0]), .Z(n1203) );
  CNIVX1 U1466 ( .A(h0[5]), .Z(n1204) );
  CNIVX1 U1467 ( .A(h0[3]), .Z(n1205) );
  CNIVX1 U1468 ( .A(h0[6]), .Z(n1206) );
  CNIVX1 U1469 ( .A(h0[4]), .Z(n1207) );
  CNIVX1 U1470 ( .A(h0[2]), .Z(n1208) );
  CNIVX1 U1471 ( .A(n600), .Z(n1209) );
  CNIVX1 U1472 ( .A(n610), .Z(n1210) );
  CNIVX1 U1473 ( .A(n1212), .Z(n1211) );
  CNIVX1 U1474 ( .A(cmd0[1]), .Z(n1212) );
  CNIVX1 U1475 ( .A(n1214), .Z(n1213) );
  CNIVX1 U1476 ( .A(cmd0[0]), .Z(n1214) );
  CNIVX1 U1477 ( .A(n1216), .Z(n1215) );
  CNIVX1 U1478 ( .A(push0), .Z(n1216) );
  CNIVX1 U1479 ( .A(n1218), .Z(n1217) );
  CNIVX1 U1480 ( .A(n611), .Z(n1218) );
  CNIVX1 U1481 ( .A(n1220), .Z(n1219) );
  CNIVX1 U1482 ( .A(push0_1), .Z(n1220) );
  CIVX4 U1483 ( .A(h0_0[1]), .Z(n1510) );
  CNIVX1 U1484 ( .A(n738), .Z(n1221) );
  CMX2XL U1485 ( .A0(out0_2[16]), .A1(out0_1[16]), .S(n1372), .Z(n738) );
  CNIVX1 U1486 ( .A(n746), .Z(n1222) );
  CMX2XL U1487 ( .A0(out0_2[8]), .A1(out0_1[8]), .S(n1380), .Z(n746) );
  CNIVX1 U1488 ( .A(n612), .Z(n1223) );
  CNIVX1 U1489 ( .A(n606), .Z(n1224) );
  CNIVX1 U1490 ( .A(n573), .Z(n1225) );
  CNIVX1 U1491 ( .A(n603), .Z(n1226) );
  CNIVX1 U1492 ( .A(n599), .Z(n1227) );
  CNIVX1 U1493 ( .A(n608), .Z(n1228) );
  CNIVX1 U1494 ( .A(n609), .Z(n1229) );
  CNIVX1 U1495 ( .A(n602), .Z(n1230) );
  CNIVX1 U1496 ( .A(n601), .Z(n1231) );
  CNIVX1 U1497 ( .A(n604), .Z(n1232) );
  CNIVX1 U1498 ( .A(n563), .Z(n1233) );
  CNIVX1 U1499 ( .A(n557), .Z(n1234) );
  CIVDX1 U1500 ( .A(cmd0_0[1]), .Z1(n1236) );
  CNIVX1 U1501 ( .A(n1236), .Z(n1235) );
  CIVDX1 U1502 ( .A(cmd0_0[0]), .Z1(n1238) );
  CNIVX1 U1503 ( .A(n1238), .Z(n1237) );
  CIVDX1 U1504 ( .A(push0_0), .Z1(n1240) );
  CNIVX1 U1505 ( .A(n1240), .Z(n1239) );
  CIVX4 U1506 ( .A(rst), .Z(n2462) );
  CDLY1XL U1507 ( .A(q0[9]), .Z(n1241) );
  CMX2XL U1508 ( .A0(q0[18]), .A1(q[18]), .S(n1497), .Z(n676) );
  CMX2XL U1509 ( .A0(n797), .A1(q[24]), .S(n1496), .Z(n682) );
  CMX2XL U1510 ( .A0(q0[12]), .A1(q[12]), .S(n1497), .Z(n670) );
  CDLY1XL U1511 ( .A(q0[29]), .Z(n1242) );
  CMX2XL U1512 ( .A0(q0[14]), .A1(q[14]), .S(n1497), .Z(n672) );
  CMX2XL U1513 ( .A0(h0[24]), .A1(h[24]), .S(n1499), .Z(n650) );
  CDLY1XL U1514 ( .A(q0[28]), .Z(n1243) );
  CDLY1XL U1515 ( .A(q0[15]), .Z(n1244) );
  CMX2XL U1516 ( .A0(q0[31]), .A1(q[31]), .S(n1496), .Z(n689) );
  CMX2XL U1517 ( .A0(h0[25]), .A1(h[25]), .S(n1499), .Z(n651) );
  CDLY1XL U1518 ( .A(q0[17]), .Z(n1245) );
  CDLY1XL U1519 ( .A(q0[25]), .Z(n1246) );
  CDLY1XL U1520 ( .A(q0[11]), .Z(n1247) );
  CMX2XL U1521 ( .A0(h0[20]), .A1(h[20]), .S(n1499), .Z(n646) );
  CMX2XL U1522 ( .A0(h0[16]), .A1(h[16]), .S(n1499), .Z(n642) );
  CMX2XL U1523 ( .A0(n1247), .A1(q[11]), .S(n1497), .Z(n669) );
  CMX2XL U1524 ( .A0(h0[21]), .A1(h[21]), .S(n1499), .Z(n647) );
  CMX2XL U1525 ( .A0(h0[10]), .A1(h[10]), .S(n1500), .Z(n636) );
  CMX2XL U1526 ( .A0(h0[7]), .A1(h[7]), .S(n1500), .Z(n633) );
  CDLY1XL U1527 ( .A(q0[1]), .Z(n1248) );
  CDLY1XL U1528 ( .A(q0[6]), .Z(n1249) );
  CMX2XL U1529 ( .A0(h0[22]), .A1(h[22]), .S(n1499), .Z(n648) );
  CDLY1XL U1530 ( .A(q0[3]), .Z(n1250) );
  CMX2XL U1531 ( .A0(n1241), .A1(q[9]), .S(n1497), .Z(n667) );
  CMX2XL U1532 ( .A0(h0[27]), .A1(h[27]), .S(n1499), .Z(n653) );
  CDLY1XL U1533 ( .A(q0[23]), .Z(n1359) );
  CMX2XL U1534 ( .A0(h0[17]), .A1(h[17]), .S(n1499), .Z(n643) );
  CMX2XL U1535 ( .A0(h0[9]), .A1(h[9]), .S(n1500), .Z(n635) );
  CMX2XL U1536 ( .A0(h0[31]), .A1(h[31]), .S(n1498), .Z(n657) );
  CDLY1XL U1537 ( .A(h0[8]), .Z(n1251) );
  CMX2XL U1538 ( .A0(n793), .A1(q[8]), .S(n1497), .Z(n666) );
  CDLY1XL U1539 ( .A(q0[21]), .Z(n1252) );
  CDLY1XL U1540 ( .A(q0[13]), .Z(n1253) );
  CDLY1XL U1541 ( .A(q0[19]), .Z(n1254) );
  CDLY1XL U1542 ( .A(q0[7]), .Z(n1358) );
  CDLY1XL U1543 ( .A(q0[27]), .Z(n1360) );
  CMX2XL U1544 ( .A0(n1204), .A1(h[5]), .S(n1500), .Z(n629) );
  CIVXL U1545 ( .A(n1204), .Z(n1505) );
  CMX2XL U1546 ( .A0(n1205), .A1(h[3]), .S(n1501), .Z(n623) );
  CIVXL U1547 ( .A(n1205), .Z(n1776) );
  CMX2XL U1548 ( .A0(n1206), .A1(h[6]), .S(n1500), .Z(n632) );
  CIVXL U1549 ( .A(n1206), .Z(n1503) );
  CMX2XL U1550 ( .A0(n1207), .A1(h[4]), .S(n1500), .Z(n626) );
  CIVXL U1551 ( .A(n1207), .Z(n1507) );
  CMX2XL U1552 ( .A0(n1208), .A1(h[2]), .S(n1501), .Z(n620) );
  CIVXL U1553 ( .A(n1208), .Z(n1512) );
  CAN2XL U1554 ( .A(n1778), .B(n2408), .Z(n1257) );
  CANR2XL U1555 ( .A(n1770), .B(acc[8]), .C(n1769), .D(out0_2[8]), .Z(n1739)
         );
  CIVX2 U1556 ( .A(h0_1[2]), .Z(n1864) );
  CMX2XL U1557 ( .A0(z[6]), .A1(acc[6]), .S(n796), .Z(n764) );
  CMX2XL U1558 ( .A0(z[14]), .A1(acc[14]), .S(n796), .Z(n772) );
  CMX2XL U1559 ( .A0(z[15]), .A1(acc[15]), .S(n796), .Z(n773) );
  CIVX2 U1560 ( .A(n1789), .Z(n2410) );
  CIVX2 U1561 ( .A(n1853), .Z(n2207) );
  CAN2XL U1562 ( .A(n2169), .B(n2168), .Z(n1268) );
  CIVX2 U1563 ( .A(n2437), .Z(n2405) );
  CIVX2 U1564 ( .A(n2435), .Z(n2406) );
  CIVX2 U1565 ( .A(n1794), .Z(n2441) );
  CAN2X1 U1566 ( .A(n2207), .B(n1488), .Z(n1258) );
  CNIVX1 U1567 ( .A(n2450), .Z(n1361) );
  CND3XL U1568 ( .A(cmd2_en_2), .B(n2033), .C(n2426), .Z(n2450) );
  CND2X1 U1569 ( .A(n2422), .B(n1488), .Z(n1887) );
  CAN2XL U1570 ( .A(n2003), .B(n2002), .Z(n1287) );
  CAN2XL U1571 ( .A(n2012), .B(n2011), .Z(n1286) );
  CAN2XL U1572 ( .A(n1940), .B(n1939), .Z(n1285) );
  CAN2XL U1573 ( .A(n1967), .B(n1966), .Z(n1282) );
  CAN2XL U1574 ( .A(n2030), .B(n2029), .Z(n1283) );
  CAN2XL U1575 ( .A(n1985), .B(n1984), .Z(n1288) );
  CAN2XL U1576 ( .A(n2021), .B(n2020), .Z(n1289) );
  CAN2XL U1577 ( .A(n1976), .B(n1975), .Z(n1291) );
  CAN2XL U1578 ( .A(n1949), .B(n1948), .Z(n1290) );
  CAN2XL U1579 ( .A(n1931), .B(n1930), .Z(n1281) );
  CAN2XL U1580 ( .A(n1958), .B(n1957), .Z(n1284) );
  CAN2XL U1581 ( .A(n1994), .B(n1993), .Z(n1292) );
  CAN2X1 U1582 ( .A(cmd1_en_2_d), .B(n2408), .Z(n1297) );
  COND3X1 U1583 ( .A(n2430), .B(n2289), .C(n2288), .D(n2287), .Z(n2290) );
  CIVX3 U1584 ( .A(h0_1[3]), .Z(n1861) );
  CANR2XL U1585 ( .A(out0_2[60]), .B(n1357), .C(N478), .D(n1298), .Z(n1530) );
  CND2XL U1586 ( .A(n1487), .B(n2207), .Z(n1922) );
  CIVXL U1587 ( .A(n2430), .Z(n2416) );
  COND1X1 U1588 ( .A(n1862), .B(n1861), .C(n1860), .Z(n2004) );
  COND1X1 U1589 ( .A(n1293), .B(n1861), .C(n1832), .Z(n1968) );
  CANR2XL U1590 ( .A(n2218), .B(n2001), .C(n2207), .D(n2127), .Z(n2002) );
  CANR2XL U1591 ( .A(n1296), .B(n2001), .C(n1295), .D(n2038), .Z(n1967) );
  CANR2XL U1592 ( .A(n2218), .B(n1929), .C(n2207), .D(n2038), .Z(n1930) );
  CANR2XL U1593 ( .A(n2218), .B(n2010), .C(n2207), .D(n2137), .Z(n2011) );
  CANR2XL U1594 ( .A(n2218), .B(n1938), .C(n2207), .D(n2051), .Z(n1939) );
  CANR2XL U1595 ( .A(n2218), .B(n2028), .C(n2207), .D(n2157), .Z(n2029) );
  CANR2XL U1596 ( .A(n2218), .B(n1947), .C(n2207), .D(n2064), .Z(n1948) );
  CANR2XL U1597 ( .A(n2218), .B(n2019), .C(n2207), .D(n2147), .Z(n2020) );
  CANR2XL U1598 ( .A(n2218), .B(n1983), .C(n2207), .D(n2107), .Z(n1984) );
  CANR2XL U1599 ( .A(n2218), .B(n1974), .C(n2207), .D(n2097), .Z(n1975) );
  CANR2XL U1600 ( .A(n2218), .B(n1956), .C(n2207), .D(n2077), .Z(n1957) );
  CANR2XL U1601 ( .A(n2218), .B(n1992), .C(n2207), .D(n2117), .Z(n1993) );
  CANR2XL U1602 ( .A(n1305), .B(n2441), .C(n1318), .D(n2410), .Z(n2222) );
  CANR2XL U1603 ( .A(n1311), .B(n2441), .C(n1319), .D(n2410), .Z(n2234) );
  CANR2XL U1604 ( .A(n1303), .B(n2441), .C(n1320), .D(n2410), .Z(n2246) );
  CANR2XL U1605 ( .A(n1319), .B(n2441), .C(n1322), .D(n2410), .Z(n2272) );
  CANR2XL U1606 ( .A(n1320), .B(n2441), .C(n1323), .D(n2410), .Z(n2285) );
  CANR2XL U1607 ( .A(n1317), .B(n2441), .C(n1324), .D(n2410), .Z(n2298) );
  CND2XL U1608 ( .A(n1295), .B(n1488), .Z(n2420) );
  CND2XL U1609 ( .A(n1296), .B(n1488), .Z(n2443) );
  CANR2XL U1610 ( .A(n2218), .B(n2167), .C(n2207), .D(n2315), .Z(n2168) );
  CAN2XL U1611 ( .A(n1258), .B(n1300), .Z(n1255) );
  CAN3XL U1612 ( .A(n2410), .B(n1864), .C(n1806), .Z(n1293) );
  CIVXL U1613 ( .A(n1169), .Z(n1490) );
  CANR2XL U1614 ( .A(n1770), .B(acc[13]), .C(n1769), .D(out0_2[13]), .Z(n1719)
         );
  CANR2XL U1615 ( .A(n1770), .B(acc[18]), .C(n1769), .D(out0_2[18]), .Z(n1699)
         );
  CANR2XL U1616 ( .A(n1770), .B(acc[12]), .C(n1769), .D(out0_2[12]), .Z(n1723)
         );
  CANR2XL U1617 ( .A(n1770), .B(acc[24]), .C(n1769), .D(out0_2[24]), .Z(n1675)
         );
  CANR2XL U1618 ( .A(n1770), .B(acc[26]), .C(n1769), .D(out0_2[26]), .Z(n1667)
         );
  CANR2XL U1619 ( .A(n1770), .B(acc[19]), .C(n1769), .D(out0_2[19]), .Z(n1695)
         );
  CANR2XL U1620 ( .A(n1770), .B(acc[25]), .C(n1769), .D(out0_2[25]), .Z(n1671)
         );
  CANR2XL U1621 ( .A(n1770), .B(acc[27]), .C(n1769), .D(out0_2[27]), .Z(n1663)
         );
  CANR2XL U1622 ( .A(n1770), .B(acc[2]), .C(n1769), .D(out0_2[2]), .Z(n1763)
         );
  CANR2XL U1623 ( .A(n1770), .B(acc[41]), .C(n1769), .D(out0_2[41]), .Z(n1607)
         );
  CANR2XL U1624 ( .A(n1770), .B(acc[10]), .C(n1769), .D(out0_2[10]), .Z(n1731)
         );
  CANR2XL U1625 ( .A(n1770), .B(acc[11]), .C(n1769), .D(out0_2[11]), .Z(n1727)
         );
  CANR2XL U1626 ( .A(n1770), .B(acc[16]), .C(n1769), .D(out0_2[16]), .Z(n1707)
         );
  CANR2XL U1627 ( .A(n1770), .B(acc[33]), .C(n1769), .D(out0_2[33]), .Z(n1639)
         );
  CANR2XL U1628 ( .A(n1770), .B(acc[5]), .C(n1769), .D(out0_2[5]), .Z(n1751)
         );
  CANR2XL U1629 ( .A(n1770), .B(acc[4]), .C(n1769), .D(out0_2[4]), .Z(n1755)
         );
  CANR2XL U1630 ( .A(n1770), .B(acc[1]), .C(n1769), .D(out0_2[1]), .Z(n1767)
         );
  CANR2XL U1631 ( .A(n1770), .B(acc[0]), .C(n1769), .D(out0_2[0]), .Z(n1771)
         );
  CANR2XL U1632 ( .A(n1770), .B(acc[3]), .C(n1769), .D(out0_2[3]), .Z(n1759)
         );
  CANR2XL U1633 ( .A(n1770), .B(acc[63]), .C(n1769), .D(out0_2[63]), .Z(n1517)
         );
  COAN1XL U1634 ( .A(n2408), .B(n1783), .C(n1782), .Z(n1301) );
  CANR2XL U1635 ( .A(acc[62]), .B(n1257), .C(out1_2[62]), .D(n1297), .Z(n1782)
         );
  COAN1XL U1636 ( .A(n2408), .B(n1857), .C(n1856), .Z(n1337) );
  CANR2XL U1637 ( .A(acc[51]), .B(n1257), .C(out1_2[51]), .D(n1297), .Z(n1856)
         );
  COAN1XL U1638 ( .A(n2408), .B(n1842), .C(n1841), .Z(n1338) );
  CANR2XL U1639 ( .A(acc[53]), .B(n1257), .C(out1_2[53]), .D(n1297), .Z(n1841)
         );
  COAN1XL U1640 ( .A(n2408), .B(n1889), .C(n1888), .Z(n1335) );
  CANR2XL U1641 ( .A(acc[47]), .B(n1257), .C(out1_2[47]), .D(n1297), .Z(n1888)
         );
  COAN1XL U1642 ( .A(n2408), .B(n1874), .C(n1873), .Z(n1336) );
  CANR2XL U1643 ( .A(acc[49]), .B(n1257), .C(out1_2[49]), .D(n1297), .Z(n1873)
         );
  COAN1XL U1644 ( .A(n2408), .B(n1829), .C(n1828), .Z(n1343) );
  CANR2XL U1645 ( .A(acc[55]), .B(n1257), .C(out1_2[55]), .D(n1297), .Z(n1828)
         );
  COAN1XL U1646 ( .A(n2408), .B(n1817), .C(n1816), .Z(n1344) );
  CANR2XL U1647 ( .A(acc[57]), .B(n1257), .C(out1_2[57]), .D(n1297), .Z(n1816)
         );
  COAN1XL U1648 ( .A(n2408), .B(n1803), .C(n1802), .Z(n1316) );
  CANR2XL U1649 ( .A(acc[59]), .B(n1257), .C(out1_2[59]), .D(n1297), .Z(n1802)
         );
  COAN1XL U1650 ( .A(n2408), .B(n1796), .C(n1795), .Z(n1326) );
  CANR2XL U1651 ( .A(acc[60]), .B(n1257), .C(out1_2[60]), .D(n1297), .Z(n1795)
         );
  COAN1XL U1652 ( .A(n2408), .B(n1867), .C(n1866), .Z(n1350) );
  CANR2XL U1653 ( .A(acc[50]), .B(n1257), .C(out1_2[50]), .D(n1297), .Z(n1866)
         );
  COAN1XL U1654 ( .A(n2408), .B(n1881), .C(n1880), .Z(n1351) );
  CANR2XL U1655 ( .A(acc[48]), .B(n1257), .C(out1_2[48]), .D(n1297), .Z(n1880)
         );
  COAN1XL U1656 ( .A(n2408), .B(n2144), .C(n2143), .Z(n1304) );
  CANR2XL U1657 ( .A(acc[21]), .B(n1257), .C(out1_2[21]), .D(n1297), .Z(n2143)
         );
  COAN1XL U1658 ( .A(n2408), .B(n2134), .C(n2133), .Z(n1306) );
  CANR2XL U1659 ( .A(acc[22]), .B(n1257), .C(out1_2[22]), .D(n1297), .Z(n2133)
         );
  COAN1XL U1660 ( .A(n2408), .B(n1835), .C(n1834), .Z(n1348) );
  CANR2XL U1661 ( .A(acc[54]), .B(n1257), .C(out1_2[54]), .D(n1297), .Z(n1834)
         );
  COAN1XL U1662 ( .A(n2408), .B(n2164), .C(n2163), .Z(n1302) );
  CANR2XL U1663 ( .A(acc[19]), .B(n1257), .C(out1_2[19]), .D(n1297), .Z(n2163)
         );
  COAN1XL U1664 ( .A(n2408), .B(n2104), .C(n2103), .Z(n1328) );
  CANR2XL U1665 ( .A(acc[25]), .B(n1257), .C(out1_2[25]), .D(n1297), .Z(n2103)
         );
  COAN1XL U1666 ( .A(n2408), .B(n1849), .C(n1848), .Z(n1349) );
  CANR2XL U1667 ( .A(acc[52]), .B(n1257), .C(out1_2[52]), .D(n1297), .Z(n1848)
         );
  COAN1XL U1668 ( .A(n2408), .B(n2174), .C(n2173), .Z(n1308) );
  CANR2XL U1669 ( .A(acc[18]), .B(n1257), .C(out1_2[18]), .D(n1297), .Z(n2173)
         );
  COAN1XL U1670 ( .A(n2408), .B(n2204), .C(n2203), .Z(n1303) );
  CANR2XL U1671 ( .A(acc[15]), .B(n1257), .C(out1_2[15]), .D(n1297), .Z(n2203)
         );
  COAN1XL U1672 ( .A(n2408), .B(n2154), .C(n2153), .Z(n1309) );
  CANR2XL U1673 ( .A(acc[20]), .B(n1257), .C(out1_2[20]), .D(n1297), .Z(n2153)
         );
  COAN1XL U1674 ( .A(n2408), .B(n2195), .C(n2194), .Z(n1311) );
  CANR2XL U1675 ( .A(acc[16]), .B(n1257), .C(out1_2[16]), .D(n1297), .Z(n2194)
         );
  COAN1XL U1676 ( .A(n2408), .B(n2184), .C(n2183), .Z(n1305) );
  CANR2XL U1677 ( .A(acc[17]), .B(n1257), .C(out1_2[17]), .D(n1297), .Z(n2183)
         );
  COAN1XL U1678 ( .A(n2408), .B(n2061), .C(n2060), .Z(n1310) );
  CANR2XL U1679 ( .A(acc[29]), .B(n1257), .C(out1_2[29]), .D(n1297), .Z(n2060)
         );
  COAN1XL U1680 ( .A(n2408), .B(n2124), .C(n2123), .Z(n1312) );
  CANR2XL U1681 ( .A(acc[23]), .B(n1257), .C(out1_2[23]), .D(n1297), .Z(n2123)
         );
  COAN1XL U1682 ( .A(n2408), .B(n2084), .C(n2083), .Z(n1307) );
  CANR2XL U1683 ( .A(acc[27]), .B(n1257), .C(out1_2[27]), .D(n1297), .Z(n2083)
         );
  COAN1XL U1684 ( .A(n2408), .B(n2114), .C(n2113), .Z(n1327) );
  CANR2XL U1685 ( .A(acc[24]), .B(n1257), .C(out1_2[24]), .D(n1297), .Z(n2113)
         );
  COAN1XL U1686 ( .A(n2408), .B(n2007), .C(n2006), .Z(n1331) );
  CANR2XL U1687 ( .A(acc[34]), .B(n1257), .C(out1_2[34]), .D(n1297), .Z(n2006)
         );
  COAN1XL U1688 ( .A(n2408), .B(n2016), .C(n2015), .Z(n1332) );
  CANR2XL U1689 ( .A(acc[33]), .B(n1257), .C(out1_2[33]), .D(n1297), .Z(n2015)
         );
  COAN1XL U1690 ( .A(n2408), .B(n1998), .C(n1997), .Z(n1333) );
  CANR2XL U1691 ( .A(acc[35]), .B(n1257), .C(out1_2[35]), .D(n1297), .Z(n1997)
         );
  COAN1XL U1692 ( .A(n2408), .B(n1989), .C(n1988), .Z(n1334) );
  CANR2XL U1693 ( .A(acc[36]), .B(n1257), .C(out1_2[36]), .D(n1297), .Z(n1988)
         );
  COAN1XL U1694 ( .A(n2408), .B(n2035), .C(n2034), .Z(n1329) );
  CANR2XL U1695 ( .A(acc[31]), .B(n1257), .C(out1_2[31]), .D(n1297), .Z(n2034)
         );
  COAN1XL U1696 ( .A(n2408), .B(n2025), .C(n2024), .Z(n1330) );
  CANR2XL U1697 ( .A(acc[32]), .B(n1257), .C(out1_2[32]), .D(n1297), .Z(n2024)
         );
  COAN1XL U1698 ( .A(n2408), .B(n2048), .C(n2047), .Z(n1314) );
  CANR2XL U1699 ( .A(acc[30]), .B(n1257), .C(out1_2[30]), .D(n1297), .Z(n2047)
         );
  COAN1XL U1700 ( .A(n2408), .B(n1971), .C(n1970), .Z(n1339) );
  CANR2XL U1701 ( .A(acc[38]), .B(n1257), .C(out1_2[38]), .D(n1297), .Z(n1970)
         );
  COAN1XL U1702 ( .A(n2408), .B(n1980), .C(n1979), .Z(n1340) );
  CANR2XL U1703 ( .A(acc[37]), .B(n1257), .C(out1_2[37]), .D(n1297), .Z(n1979)
         );
  COAN1XL U1704 ( .A(n2408), .B(n1962), .C(n1961), .Z(n1355) );
  CANR2XL U1705 ( .A(acc[39]), .B(n1257), .C(out1_2[39]), .D(n1297), .Z(n1961)
         );
  COAN1XL U1706 ( .A(n2408), .B(n1916), .C(n1915), .Z(n1341) );
  CANR2XL U1707 ( .A(acc[44]), .B(n1257), .C(out1_2[44]), .D(n1297), .Z(n1915)
         );
  COAN1XL U1708 ( .A(n2408), .B(n1926), .C(n1925), .Z(n1342) );
  CANR2XL U1709 ( .A(acc[43]), .B(n1257), .C(out1_2[43]), .D(n1297), .Z(n1925)
         );
  COAN1XL U1710 ( .A(n2408), .B(n1935), .C(n1934), .Z(n1353) );
  CANR2XL U1711 ( .A(acc[42]), .B(n1257), .C(out1_2[42]), .D(n1297), .Z(n1934)
         );
  COAN1XL U1712 ( .A(n2408), .B(n2074), .C(n2073), .Z(n1313) );
  CANR2XL U1713 ( .A(acc[28]), .B(n1257), .C(out1_2[28]), .D(n1297), .Z(n2073)
         );
  COAN1XL U1714 ( .A(n2408), .B(n2094), .C(n2093), .Z(n1315) );
  CANR2XL U1715 ( .A(acc[26]), .B(n1257), .C(out1_2[26]), .D(n1297), .Z(n2093)
         );
  COAN1XL U1716 ( .A(n2408), .B(n1898), .C(n1897), .Z(n1352) );
  CANR2XL U1717 ( .A(acc[46]), .B(n1257), .C(out1_2[46]), .D(n1297), .Z(n1897)
         );
  COAN1XL U1718 ( .A(n2408), .B(n1810), .C(n1809), .Z(n1345) );
  CANR2XL U1719 ( .A(acc[58]), .B(n1257), .C(out1_2[58]), .D(n1297), .Z(n1809)
         );
  COAN1XL U1720 ( .A(n2408), .B(n1823), .C(n1822), .Z(n1346) );
  CANR2XL U1721 ( .A(acc[56]), .B(n1257), .C(out1_2[56]), .D(n1297), .Z(n1822)
         );
  COAN1XL U1722 ( .A(n2408), .B(n1953), .C(n1952), .Z(n1354) );
  CANR2XL U1723 ( .A(acc[40]), .B(n1257), .C(out1_2[40]), .D(n1297), .Z(n1952)
         );
  COAN1XL U1724 ( .A(n2408), .B(n1944), .C(n1943), .Z(n1356) );
  CANR2XL U1725 ( .A(acc[41]), .B(n1257), .C(out1_2[41]), .D(n1297), .Z(n1943)
         );
  COAN1XL U1726 ( .A(n2408), .B(n1907), .C(n1906), .Z(n1347) );
  CANR2XL U1727 ( .A(acc[45]), .B(n1257), .C(out1_2[45]), .D(n1297), .Z(n1906)
         );
  COAN1XL U1728 ( .A(n2408), .B(n2258), .C(n2257), .Z(n1317) );
  CANR2XL U1729 ( .A(acc[11]), .B(n1257), .C(out1_2[11]), .D(n1297), .Z(n2257)
         );
  COAN1XL U1730 ( .A(n2408), .B(n2310), .C(n2309), .Z(n1321) );
  CANR2XL U1731 ( .A(acc[7]), .B(n1257), .C(out1_2[7]), .D(n1297), .Z(n2309)
         );
  COAN1XL U1732 ( .A(n2408), .B(n2233), .C(n2232), .Z(n1319) );
  CANR2XL U1733 ( .A(acc[13]), .B(n1257), .C(out1_2[13]), .D(n1297), .Z(n2232)
         );
  COAN1XL U1734 ( .A(n2408), .B(n2284), .C(n2283), .Z(n1323) );
  CANR2XL U1735 ( .A(acc[9]), .B(n1257), .C(out1_2[9]), .D(n1297), .Z(n2283)
         );
  COAN1XL U1736 ( .A(n2408), .B(n2221), .C(n2220), .Z(n1318) );
  CANR2XL U1737 ( .A(acc[14]), .B(n1257), .C(out1_2[14]), .D(n1297), .Z(n2220)
         );
  COAN1XL U1738 ( .A(n2408), .B(n2271), .C(n2270), .Z(n1322) );
  CANR2XL U1739 ( .A(acc[10]), .B(n1257), .C(out1_2[10]), .D(n1297), .Z(n2270)
         );
  COAN1XL U1740 ( .A(n2408), .B(n2245), .C(n2244), .Z(n1320) );
  CANR2XL U1741 ( .A(acc[12]), .B(n1257), .C(out1_2[12]), .D(n1297), .Z(n2244)
         );
  COAN1XL U1742 ( .A(n2408), .B(n2297), .C(n2296), .Z(n1324) );
  CANR2XL U1743 ( .A(acc[8]), .B(n1257), .C(out1_2[8]), .D(n1297), .Z(n2296)
         );
  COAN1XL U1744 ( .A(n2408), .B(n2322), .C(n2321), .Z(n1325) );
  CANR2XL U1745 ( .A(acc[6]), .B(n1257), .C(out1_2[6]), .D(n1297), .Z(n2321)
         );
  CND2XL U1746 ( .A(h0_1[2]), .B(h0_1[3]), .Z(n1865) );
  CANR2XL U1747 ( .A(out0_2[26]), .B(n1357), .C(N444), .D(n1298), .Z(n1666) );
  CANR2XL U1748 ( .A(acc[61]), .B(n1257), .C(out1_2[61]), .D(n1297), .Z(n1786)
         );
  CANR2XL U1749 ( .A(n1770), .B(acc[23]), .C(n1769), .D(out0_2[23]), .Z(n1679)
         );
  CANR2XL U1750 ( .A(n1770), .B(acc[22]), .C(n1769), .D(out0_2[22]), .Z(n1683)
         );
  CANR2XL U1751 ( .A(n1770), .B(acc[20]), .C(n1769), .D(out0_2[20]), .Z(n1691)
         );
  CANR2XL U1752 ( .A(n1770), .B(acc[21]), .C(n1769), .D(out0_2[21]), .Z(n1687)
         );
  CANR2XL U1753 ( .A(n1770), .B(acc[29]), .C(n1769), .D(out0_2[29]), .Z(n1655)
         );
  CANR2XL U1754 ( .A(n1770), .B(acc[28]), .C(n1769), .D(out0_2[28]), .Z(n1659)
         );
  CANR2XL U1755 ( .A(n1770), .B(acc[30]), .C(n1769), .D(out0_2[30]), .Z(n1651)
         );
  CANR2XL U1756 ( .A(n1770), .B(acc[49]), .C(n1769), .D(out0_2[49]), .Z(n1575)
         );
  CANR2XL U1757 ( .A(n1770), .B(acc[58]), .C(n1769), .D(out0_2[58]), .Z(n1539)
         );
  CANR2XL U1758 ( .A(n1770), .B(acc[35]), .C(n1769), .D(out0_2[35]), .Z(n1631)
         );
  CANR2XL U1759 ( .A(n1770), .B(acc[34]), .C(n1769), .D(out0_2[34]), .Z(n1635)
         );
  CANR2XL U1760 ( .A(n1770), .B(acc[14]), .C(n1769), .D(out0_2[14]), .Z(n1715)
         );
  CANR2XL U1761 ( .A(n1770), .B(acc[40]), .C(n1769), .D(out0_2[40]), .Z(n1611)
         );
  CANR2XL U1762 ( .A(n1770), .B(acc[57]), .C(n1769), .D(out0_2[57]), .Z(n1543)
         );
  CANR2XL U1763 ( .A(n1770), .B(acc[43]), .C(n1769), .D(out0_2[43]), .Z(n1599)
         );
  CANR2XL U1764 ( .A(n1770), .B(acc[6]), .C(n1769), .D(out0_2[6]), .Z(n1747)
         );
  CANR2XL U1765 ( .A(n1770), .B(acc[51]), .C(n1769), .D(out0_2[51]), .Z(n1567)
         );
  CANR2XL U1766 ( .A(n1770), .B(acc[31]), .C(n1769), .D(out0_2[31]), .Z(n1647)
         );
  CANR2XL U1767 ( .A(n1770), .B(acc[48]), .C(n1769), .D(out0_2[48]), .Z(n1579)
         );
  CANR2XL U1768 ( .A(n1770), .B(acc[50]), .C(n1769), .D(out0_2[50]), .Z(n1571)
         );
  CANR2XL U1769 ( .A(n1770), .B(acc[42]), .C(n1769), .D(out0_2[42]), .Z(n1603)
         );
  CANR2XL U1770 ( .A(n1770), .B(acc[45]), .C(n1769), .D(out0_2[45]), .Z(n1591)
         );
  CANR2XL U1771 ( .A(n1770), .B(acc[56]), .C(n1769), .D(out0_2[56]), .Z(n1547)
         );
  CANR2XL U1772 ( .A(n1770), .B(acc[32]), .C(n1769), .D(out0_2[32]), .Z(n1643)
         );
  CANR2XL U1773 ( .A(n1770), .B(acc[47]), .C(n1769), .D(out0_2[47]), .Z(n1583)
         );
  CANR2XL U1774 ( .A(n1770), .B(acc[15]), .C(n1769), .D(out0_2[15]), .Z(n1711)
         );
  CANR2XL U1775 ( .A(n1770), .B(acc[59]), .C(n1769), .D(out0_2[59]), .Z(n1535)
         );
  CANR2XL U1776 ( .A(n1770), .B(acc[39]), .C(n1769), .D(out0_2[39]), .Z(n1615)
         );
  CANR2XL U1777 ( .A(n1770), .B(acc[7]), .C(n1769), .D(out0_2[7]), .Z(n1743)
         );
  CANR2XL U1778 ( .A(n1770), .B(acc[52]), .C(n1769), .D(out0_2[52]), .Z(n1563)
         );
  CANR2XL U1779 ( .A(n1770), .B(acc[44]), .C(n1769), .D(out0_2[44]), .Z(n1595)
         );
  CANR2XL U1780 ( .A(n1770), .B(acc[53]), .C(n1769), .D(out0_2[53]), .Z(n1559)
         );
  CANR2XL U1781 ( .A(n1770), .B(acc[54]), .C(n1769), .D(out0_2[54]), .Z(n1555)
         );
  CANR2XL U1782 ( .A(n1770), .B(acc[46]), .C(n1769), .D(out0_2[46]), .Z(n1587)
         );
  CANR2XL U1783 ( .A(n1770), .B(acc[55]), .C(n1769), .D(out0_2[55]), .Z(n1551)
         );
  CANR2XL U1784 ( .A(n1770), .B(acc[38]), .C(n1769), .D(out0_2[38]), .Z(n1619)
         );
  CANR2XL U1785 ( .A(n1770), .B(acc[60]), .C(n1769), .D(out0_2[60]), .Z(n1531)
         );
  CANR2XL U1786 ( .A(n1770), .B(acc[37]), .C(n1769), .D(out0_2[37]), .Z(n1623)
         );
  CANR2XL U1787 ( .A(acc[3]), .B(n1257), .C(out1_2[3]), .D(n1297), .Z(n2364)
         );
  CANR2XL U1788 ( .A(n1770), .B(acc[36]), .C(n1769), .D(out0_2[36]), .Z(n1627)
         );
  CANR2XL U1789 ( .A(acc[1]), .B(n1257), .C(out1_2[1]), .D(n1297), .Z(n2391)
         );
  CANR2XL U1790 ( .A(n1770), .B(acc[61]), .C(n1769), .D(out0_2[61]), .Z(n1527)
         );
  CANR2XL U1791 ( .A(acc[4]), .B(n1257), .C(out1_2[4]), .D(n1297), .Z(n2347)
         );
  CANR2XL U1792 ( .A(acc[2]), .B(n1257), .C(out1_2[2]), .D(n1297), .Z(n2377)
         );
  CANR2XL U1793 ( .A(acc[5]), .B(n1257), .C(out1_2[5]), .D(n1297), .Z(n2334)
         );
  CIVX1 U1794 ( .A(n2376), .Z(n2387) );
  CIVX1 U1795 ( .A(n2404), .Z(n2423) );
  CIVX1 U1796 ( .A(n2268), .Z(n2278) );
  CIVX1 U1797 ( .A(n2294), .Z(n2304) );
  CIVX1 U1798 ( .A(n2255), .Z(n2265) );
  CANR2XL U1799 ( .A(n1257), .B(acc[0]), .C(n1297), .D(out1_2[0]), .Z(n2407)
         );
  CANR2XL U1800 ( .A(n1770), .B(acc[62]), .C(n1769), .D(out0_2[62]), .Z(n1523)
         );
  CMXI2XL U1801 ( .A0(n1861), .A1(n1777), .S(cmd2_en_1), .Z(n621) );
  CANR2XL U1802 ( .A(out0_2[61]), .B(n1357), .C(N479), .D(n1298), .Z(n1526) );
  CANR2XL U1803 ( .A(out0_2[57]), .B(n1357), .C(N475), .D(n1298), .Z(n1542) );
  CANR2XL U1804 ( .A(out0_2[55]), .B(n1357), .C(N473), .D(n1298), .Z(n1550) );
  CANR2XL U1805 ( .A(out0_2[53]), .B(n1357), .C(N471), .D(n1298), .Z(n1558) );
  CANR2XL U1806 ( .A(out0_2[51]), .B(n1357), .C(N469), .D(n1298), .Z(n1566) );
  CANR2XL U1807 ( .A(out0_2[49]), .B(n1357), .C(N467), .D(n1298), .Z(n1574) );
  CANR2XL U1808 ( .A(out0_2[47]), .B(n1357), .C(N465), .D(n1298), .Z(n1582) );
  CANR2XL U1809 ( .A(out0_2[45]), .B(n1357), .C(N463), .D(n1298), .Z(n1590) );
  CANR2XL U1810 ( .A(out0_2[43]), .B(n1357), .C(N461), .D(n1298), .Z(n1598) );
  CANR2XL U1811 ( .A(out0_2[41]), .B(n1357), .C(N459), .D(n1298), .Z(n1606) );
  CANR2XL U1812 ( .A(out0_2[40]), .B(n1357), .C(N458), .D(n1298), .Z(n1610) );
  CANR2XL U1813 ( .A(out0_2[39]), .B(n1357), .C(N457), .D(n1298), .Z(n1614) );
  CANR2XL U1814 ( .A(out0_2[37]), .B(n1357), .C(N455), .D(n1298), .Z(n1622) );
  CANR2XL U1815 ( .A(out0_2[35]), .B(n1357), .C(N453), .D(n1298), .Z(n1630) );
  CANR2XL U1816 ( .A(out0_2[34]), .B(n1357), .C(N452), .D(n1298), .Z(n1634) );
  CANR2XL U1817 ( .A(out0_2[33]), .B(n1357), .C(N451), .D(n1298), .Z(n1638) );
  CANR2XL U1818 ( .A(out0_2[32]), .B(n1357), .C(N450), .D(n1298), .Z(n1642) );
  CANR2XL U1819 ( .A(out0_2[31]), .B(n1357), .C(N449), .D(n1298), .Z(n1646) );
  CANR2XL U1820 ( .A(out0_2[29]), .B(n1357), .C(N447), .D(n1298), .Z(n1654) );
  CANR2XL U1821 ( .A(out0_2[27]), .B(n1357), .C(N445), .D(n1298), .Z(n1662) );
  CANR2XL U1822 ( .A(out0_2[25]), .B(n1357), .C(N443), .D(n1298), .Z(n1670) );
  CANR2XL U1823 ( .A(out0_2[24]), .B(n1357), .C(N442), .D(n1298), .Z(n1674) );
  CANR2XL U1824 ( .A(out0_2[23]), .B(n1357), .C(N441), .D(n1298), .Z(n1678) );
  CANR2XL U1825 ( .A(out0_2[21]), .B(n1357), .C(N439), .D(n1298), .Z(n1686) );
  CANR2XL U1826 ( .A(out0_2[20]), .B(n1357), .C(N438), .D(n1298), .Z(n1690) );
  CANR2XL U1827 ( .A(out0_2[19]), .B(n1357), .C(N437), .D(n1298), .Z(n1694) );
  CANR2XL U1828 ( .A(out0_2[18]), .B(n1357), .C(N436), .D(n1298), .Z(n1698) );
  CANR2XL U1829 ( .A(out0_2[17]), .B(n1357), .C(N435), .D(n1298), .Z(n1702) );
  CANR2XL U1830 ( .A(out0_2[16]), .B(n1357), .C(N434), .D(n1298), .Z(n1706) );
  CANR2XL U1831 ( .A(out0_2[15]), .B(n1357), .C(N433), .D(n1298), .Z(n1710) );
  CANR2XL U1832 ( .A(out0_2[14]), .B(n1357), .C(N432), .D(n1298), .Z(n1714) );
  CANR2XL U1833 ( .A(out0_2[13]), .B(n1357), .C(N431), .D(n1298), .Z(n1718) );
  CANR2XL U1834 ( .A(out0_2[12]), .B(n1357), .C(N430), .D(n1298), .Z(n1722) );
  CANR2XL U1835 ( .A(out0_2[11]), .B(n1357), .C(N429), .D(n1298), .Z(n1726) );
  CANR2XL U1836 ( .A(out0_2[10]), .B(n1357), .C(N428), .D(n1298), .Z(n1730) );
  CANR2XL U1837 ( .A(out0_2[9]), .B(n1357), .C(N427), .D(n1298), .Z(n1734) );
  CANR2XL U1838 ( .A(out0_2[8]), .B(n1357), .C(N426), .D(n1298), .Z(n1738) );
  CANR2XL U1839 ( .A(out0_2[7]), .B(n1357), .C(N425), .D(n1298), .Z(n1742) );
  CANR2XL U1840 ( .A(out0_2[6]), .B(n1357), .C(N424), .D(n1298), .Z(n1746) );
  CANR2XL U1841 ( .A(out0_2[5]), .B(n1357), .C(N423), .D(n1298), .Z(n1750) );
  CANR2XL U1842 ( .A(out0_2[4]), .B(n1357), .C(N422), .D(n1298), .Z(n1754) );
  CANR2XL U1843 ( .A(out0_2[3]), .B(n1357), .C(N421), .D(n1298), .Z(n1758) );
  CANR2XL U1844 ( .A(out0_2[2]), .B(n1357), .C(N420), .D(n1298), .Z(n1762) );
  CANR2XL U1845 ( .A(out0_2[1]), .B(n1357), .C(N419), .D(n1298), .Z(n1766) );
  CMX2XL U1846 ( .A0(z[0]), .A1(acc[0]), .S(n796), .Z(n758) );
  CMX2XL U1847 ( .A0(z[1]), .A1(acc[1]), .S(n796), .Z(n759) );
  CMX2XL U1848 ( .A0(z[2]), .A1(acc[2]), .S(n796), .Z(n760) );
  CMX2XL U1849 ( .A0(z[3]), .A1(acc[3]), .S(n796), .Z(n761) );
  CMX2XL U1850 ( .A0(z[4]), .A1(acc[4]), .S(n796), .Z(n762) );
  CMX2XL U1851 ( .A0(z[5]), .A1(acc[5]), .S(n796), .Z(n763) );
  CMX2XL U1852 ( .A0(z[7]), .A1(acc[7]), .S(n796), .Z(n765) );
  CMX2XL U1853 ( .A0(z[8]), .A1(acc[8]), .S(n796), .Z(n766) );
  CMX2XL U1854 ( .A0(z[9]), .A1(acc[9]), .S(n796), .Z(n767) );
  CMX2XL U1855 ( .A0(z[10]), .A1(acc[10]), .S(n796), .Z(n768) );
  CMX2XL U1856 ( .A0(z[11]), .A1(acc[11]), .S(n796), .Z(n769) );
  CMX2XL U1857 ( .A0(z[12]), .A1(acc[12]), .S(n796), .Z(n770) );
  CMX2XL U1858 ( .A0(z[13]), .A1(acc[13]), .S(n796), .Z(n771) );
  CMX2XL U1859 ( .A0(z[16]), .A1(acc[16]), .S(n796), .Z(n774) );
  CMX2XL U1860 ( .A0(z[17]), .A1(acc[17]), .S(n796), .Z(n775) );
  CMX2XL U1861 ( .A0(z[18]), .A1(acc[18]), .S(n796), .Z(n776) );
  CMX2XL U1862 ( .A0(z[19]), .A1(acc[19]), .S(n796), .Z(n777) );
  CMX2XL U1863 ( .A0(z[21]), .A1(acc[21]), .S(n796), .Z(n779) );
  CMX2XL U1864 ( .A0(z[24]), .A1(acc[24]), .S(n796), .Z(n782) );
  CMX2XL U1865 ( .A0(z[25]), .A1(acc[25]), .S(n796), .Z(n783) );
  CMX2XL U1866 ( .A0(z[26]), .A1(acc[26]), .S(n796), .Z(n784) );
  CMX2XL U1867 ( .A0(z[27]), .A1(acc[27]), .S(n796), .Z(n785) );
  CMX2XL U1868 ( .A0(z[28]), .A1(acc[28]), .S(n796), .Z(n786) );
  CMX2XL U1869 ( .A0(z[29]), .A1(acc[29]), .S(n796), .Z(n787) );
  CIVXL U1870 ( .A(cmd2_en_2), .Z(n1494) );
  CIVXL U1871 ( .A(cmd2_en_2), .Z(n1493) );
  CIVXL U1872 ( .A(cmd2_en_2), .Z(n1492) );
  CIVXL U1873 ( .A(cmd2_en_2), .Z(n1491) );
  CMX2XL U1874 ( .A0(out0_1[28]), .A1(out0_2[28]), .S(n1365), .Z(n726) );
  CMX2XL U1875 ( .A0(out0_1[27]), .A1(out0_2[27]), .S(n1364), .Z(n727) );
  CMX2XL U1876 ( .A0(out0_1[26]), .A1(out0_2[26]), .S(n1365), .Z(n728) );
  CMX2XL U1877 ( .A0(out0_1[25]), .A1(out0_2[25]), .S(n1364), .Z(n729) );
  CAN2X1 U1878 ( .A(n2422), .B(n1486), .Z(n1256) );
  CIVX2 U1879 ( .A(n2443), .Z(n2414) );
  CIVX2 U1880 ( .A(n1361), .Z(n2422) );
  CIVX2 U1881 ( .A(n2420), .Z(n2447) );
  CIVX2 U1882 ( .A(n2448), .Z(n2192) );
  CIVX2 U1883 ( .A(n1887), .Z(n2212) );
  CIVX2 U1884 ( .A(n1865), .Z(n2218) );
  CIVX4 U1885 ( .A(n1514), .Z(n1773) );
  CIVX4 U1886 ( .A(n1515), .Z(n1770) );
  COND1XL U1887 ( .A(n2444), .B(n2443), .C(n2442), .Z(n2445) );
  CIVX2 U1888 ( .A(n1488), .Z(n1486) );
  CIVX2 U1889 ( .A(n1488), .Z(n1485) );
  CND2X1 U1890 ( .A(n2218), .B(n1488), .Z(n2430) );
  CAN2X1 U1891 ( .A(n2223), .B(n2222), .Z(n1259) );
  CAN2X1 U1892 ( .A(n2235), .B(n2234), .Z(n1260) );
  CAN2X1 U1893 ( .A(n2247), .B(n2246), .Z(n1261) );
  CAN2X1 U1894 ( .A(n2273), .B(n2272), .Z(n1262) );
  CAN2X1 U1895 ( .A(n2286), .B(n2285), .Z(n1263) );
  CAN2X1 U1896 ( .A(n2299), .B(n2298), .Z(n1264) );
  CAN2X1 U1897 ( .A(n1894), .B(n1893), .Z(n1265) );
  CAN2X1 U1898 ( .A(n2089), .B(n2088), .Z(n1266) );
  CAN2X1 U1899 ( .A(n2200), .B(n2199), .Z(n1267) );
  CAN2X1 U1900 ( .A(n2179), .B(n2178), .Z(n1269) );
  CAN2X1 U1901 ( .A(n2129), .B(n2128), .Z(n1270) );
  CAN2X1 U1902 ( .A(n2119), .B(n2118), .Z(n1271) );
  CAN2X1 U1903 ( .A(n2099), .B(n2098), .Z(n1272) );
  CAN2X1 U1904 ( .A(n2139), .B(n2138), .Z(n1273) );
  CAN2X1 U1905 ( .A(n2149), .B(n2148), .Z(n1274) );
  CAN2X1 U1906 ( .A(n2159), .B(n2158), .Z(n1275) );
  CAN2X1 U1907 ( .A(n2189), .B(n2188), .Z(n1276) );
  CAN2X1 U1908 ( .A(n2053), .B(n2052), .Z(n1277) );
  CAN2X1 U1909 ( .A(n2066), .B(n2065), .Z(n1278) );
  CAN2X1 U1910 ( .A(n2079), .B(n2078), .Z(n1279) );
  CAN2X1 U1911 ( .A(n2109), .B(n2108), .Z(n1280) );
  CAN2X1 U1912 ( .A(n2368), .B(n2367), .Z(n1294) );
  CNR3XL U1913 ( .A(n2461), .B(n2463), .C(n2464), .Z(_pushout_d) );
  CNIVX1 U1914 ( .A(n2462), .Z(n1470) );
  CNIVX1 U1915 ( .A(n2462), .Z(n1471) );
  CNIVX1 U1916 ( .A(n2462), .Z(n1468) );
  CNIVX1 U1917 ( .A(n2462), .Z(n1469) );
  CNIVX1 U1918 ( .A(n2462), .Z(n1466) );
  CNIVX1 U1919 ( .A(n2462), .Z(n1453) );
  CNIVX1 U1920 ( .A(n2462), .Z(n1467) );
  CNIVX1 U1921 ( .A(n2462), .Z(n1441) );
  CNIVX1 U1922 ( .A(n2462), .Z(n1440) );
  CNIVX1 U1923 ( .A(n2462), .Z(n1439) );
  CNIVX1 U1924 ( .A(n2462), .Z(n1438) );
  CNIVX1 U1925 ( .A(n2462), .Z(n1460) );
  CNIVX1 U1926 ( .A(n2462), .Z(n1455) );
  CNIVX1 U1927 ( .A(n2462), .Z(n1454) );
  CNIVX1 U1928 ( .A(n2462), .Z(n1465) );
  CNIVX1 U1929 ( .A(n2462), .Z(n1464) );
  CNIVX1 U1930 ( .A(n2462), .Z(n1463) );
  CNIVX1 U1931 ( .A(n2462), .Z(n1462) );
  CNIVX1 U1932 ( .A(n2462), .Z(n1461) );
  CNIVX1 U1933 ( .A(n2462), .Z(n1483) );
  CNIVX1 U1934 ( .A(n2462), .Z(n1482) );
  CNIVX1 U1935 ( .A(n2462), .Z(n1481) );
  CNIVX1 U1936 ( .A(n2462), .Z(n1480) );
  CNIVX1 U1937 ( .A(n2462), .Z(n1479) );
  CNIVX1 U1938 ( .A(n2462), .Z(n1478) );
  CNIVX1 U1939 ( .A(n2462), .Z(n1477) );
  CNIVX1 U1940 ( .A(n2462), .Z(n1476) );
  CNIVX1 U1941 ( .A(n2462), .Z(n1475) );
  CNIVX1 U1942 ( .A(n2462), .Z(n1474) );
  CNIVX1 U1943 ( .A(n2462), .Z(n1473) );
  CNIVX1 U1944 ( .A(n2462), .Z(n1452) );
  CNIVX1 U1945 ( .A(n2462), .Z(n1450) );
  CNIVX1 U1946 ( .A(n2462), .Z(n1451) );
  CNIVX1 U1947 ( .A(n2462), .Z(n1437) );
  CNIVX1 U1948 ( .A(n2462), .Z(n1449) );
  CNIVX1 U1949 ( .A(n2462), .Z(n1446) );
  CNIVX1 U1950 ( .A(n2462), .Z(n1444) );
  CNIVX1 U1951 ( .A(n2462), .Z(n1442) );
  CNIVX1 U1952 ( .A(n2462), .Z(n1472) );
  CNIVX1 U1953 ( .A(n2462), .Z(n1448) );
  CNIVX1 U1954 ( .A(n2462), .Z(n1447) );
  CNIVX1 U1955 ( .A(n2462), .Z(n1445) );
  CNIVX1 U1956 ( .A(n2462), .Z(n1443) );
  CNIVX1 U1957 ( .A(n2462), .Z(n1456) );
  CNIVX1 U1958 ( .A(n2462), .Z(n1457) );
  CNIVX1 U1959 ( .A(n2462), .Z(n1459) );
  CNIVX1 U1960 ( .A(n2462), .Z(n1458) );
  CNIVX1 U1961 ( .A(n2462), .Z(n1484) );
  COND1XL U1962 ( .A(n2408), .B(n1780), .C(n1779), .Z(n1806) );
  COND1XL U1963 ( .A(n2408), .B(n2365), .C(n2364), .Z(n2411) );
  CAN2X1 U1964 ( .A(h0_1[2]), .B(n1861), .Z(n1295) );
  COND1XL U1965 ( .A(n1773), .B(n1692), .C(n1691), .Z(acc_cmd1[20]) );
  COND1XL U1966 ( .A(n1773), .B(n1580), .C(n1579), .Z(acc_cmd1[48]) );
  COND1XL U1967 ( .A(n1773), .B(n1684), .C(n1683), .Z(acc_cmd1[22]) );
  COND1XL U1968 ( .A(n1773), .B(n1676), .C(n1675), .Z(acc_cmd1[24]) );
  COND1XL U1969 ( .A(n1773), .B(n1740), .C(n1739), .Z(acc_cmd1[8]) );
  COND1XL U1970 ( .A(n1773), .B(n1724), .C(n1723), .Z(acc_cmd1[12]) );
  COND1XL U1971 ( .A(n1773), .B(n1556), .C(n1555), .Z(acc_cmd1[54]) );
  COND1XL U1972 ( .A(n1773), .B(n1688), .C(n1687), .Z(acc_cmd1[21]) );
  COND1XL U1973 ( .A(n1773), .B(n1708), .C(n1707), .Z(acc_cmd1[16]) );
  COND1XL U1974 ( .A(n1773), .B(n1564), .C(n1563), .Z(acc_cmd1[52]) );
  COND1XL U1975 ( .A(n1773), .B(n1660), .C(n1659), .Z(acc_cmd1[28]) );
  COND1XL U1976 ( .A(n1773), .B(n1560), .C(n1559), .Z(acc_cmd1[53]) );
  COND1XL U1977 ( .A(n1773), .B(n1572), .C(n1571), .Z(acc_cmd1[50]) );
  COND1XL U1978 ( .A(n1773), .B(n1756), .C(n1755), .Z(acc_cmd1[4]) );
  COND1XL U1979 ( .A(n1773), .B(n1764), .C(n1763), .Z(acc_cmd1[2]) );
  COND1XL U1980 ( .A(n1773), .B(n1772), .C(n1771), .Z(acc_cmd1[0]) );
  COND1XL U1981 ( .A(n1773), .B(n1518), .C(n1517), .Z(acc_cmd1[63]) );
  COND1XL U1982 ( .A(n2408), .B(n2378), .C(n2377), .Z(n2440) );
  COND1XL U1983 ( .A(n2408), .B(n2348), .C(n2347), .Z(n2393) );
  CIVX4 U1984 ( .A(n1516), .Z(n1769) );
  CAN2X1 U1985 ( .A(h0_1[3]), .B(n1864), .Z(n1296) );
  CAN2X1 U1986 ( .A(n1519), .B(push0_2), .Z(n1298) );
  CAN2X1 U1987 ( .A(n1520), .B(push0_2), .Z(n1299) );
  COND1XL U1988 ( .A(n2409), .B(n2408), .C(n2407), .Z(n2434) );
  COND1XL U1989 ( .A(n2408), .B(n2335), .C(n2334), .Z(n2379) );
  COND1XL U1990 ( .A(n2408), .B(n1787), .C(n1786), .Z(n1791) );
  CND2XL U1991 ( .A(n2410), .B(n1806), .Z(n1807) );
  CAN3X2 U1992 ( .A(h0_1[5]), .B(cmd2_en_2), .C(n2033), .Z(n1300) );
  COND1XL U1993 ( .A(n1773), .B(n1680), .C(n1679), .Z(acc_cmd1[23]) );
  COND1XL U1994 ( .A(n1773), .B(n1588), .C(n1587), .Z(acc_cmd1[46]) );
  COND1XL U1995 ( .A(n1773), .B(n1636), .C(n1635), .Z(acc_cmd1[34]) );
  COND1XL U1996 ( .A(n1773), .B(n1620), .C(n1619), .Z(acc_cmd1[38]) );
  COND1XL U1997 ( .A(n1773), .B(n1700), .C(n1699), .Z(acc_cmd1[18]) );
  COND1XL U1998 ( .A(n1773), .B(n1584), .C(n1583), .Z(acc_cmd1[47]) );
  COND1XL U1999 ( .A(n1773), .B(n1628), .C(n1627), .Z(acc_cmd1[36]) );
  COND1XL U2000 ( .A(n1773), .B(n1612), .C(n1611), .Z(acc_cmd1[40]) );
  COND1XL U2001 ( .A(n1773), .B(n1716), .C(n1715), .Z(acc_cmd1[14]) );
  COND1XL U2002 ( .A(n1773), .B(n1592), .C(n1591), .Z(acc_cmd1[45]) );
  COND1XL U2003 ( .A(n1773), .B(n1720), .C(n1719), .Z(acc_cmd1[13]) );
  COND1XL U2004 ( .A(n1773), .B(n1616), .C(n1615), .Z(acc_cmd1[39]) );
  COND1XL U2005 ( .A(n1773), .B(n1748), .C(n1747), .Z(acc_cmd1[6]) );
  COND1XL U2006 ( .A(n1773), .B(n1704), .C(n1703), .Z(acc_cmd1[17]) );
  COND1XL U2007 ( .A(n1773), .B(n1728), .C(n1727), .Z(acc_cmd1[11]) );
  COND1XL U2008 ( .A(n1773), .B(n1640), .C(n1639), .Z(acc_cmd1[33]) );
  COND1XL U2009 ( .A(n1773), .B(n1600), .C(n1599), .Z(acc_cmd1[43]) );
  COND1XL U2010 ( .A(n1773), .B(n1596), .C(n1595), .Z(acc_cmd1[44]) );
  COND1XL U2011 ( .A(n1773), .B(n1736), .C(n1735), .Z(acc_cmd1[9]) );
  COND1XL U2012 ( .A(n1773), .B(n1672), .C(n1671), .Z(acc_cmd1[25]) );
  COND1XL U2013 ( .A(n1773), .B(n1604), .C(n1603), .Z(acc_cmd1[42]) );
  COND1XL U2014 ( .A(n1773), .B(n1576), .C(n1575), .Z(acc_cmd1[49]) );
  COND1XL U2015 ( .A(n1773), .B(n1632), .C(n1631), .Z(acc_cmd1[35]) );
  COND1XL U2016 ( .A(n1773), .B(n1652), .C(n1651), .Z(acc_cmd1[30]) );
  COND1XL U2017 ( .A(n1773), .B(n1624), .C(n1623), .Z(acc_cmd1[37]) );
  COND1XL U2018 ( .A(n1773), .B(n1696), .C(n1695), .Z(acc_cmd1[19]) );
  COND1XL U2019 ( .A(n1773), .B(n1732), .C(n1731), .Z(acc_cmd1[10]) );
  COND1XL U2020 ( .A(n1773), .B(n1656), .C(n1655), .Z(acc_cmd1[29]) );
  COND1XL U2021 ( .A(n1773), .B(n1664), .C(n1663), .Z(acc_cmd1[27]) );
  COND1XL U2022 ( .A(n1773), .B(n1668), .C(n1667), .Z(acc_cmd1[26]) );
  COND1XL U2023 ( .A(n1773), .B(n1752), .C(n1751), .Z(acc_cmd1[5]) );
  COND1XL U2024 ( .A(n1773), .B(n1568), .C(n1567), .Z(acc_cmd1[51]) );
  COND1XL U2025 ( .A(n1773), .B(n1712), .C(n1711), .Z(acc_cmd1[15]) );
  COND1XL U2026 ( .A(n1773), .B(n1540), .C(n1539), .Z(acc_cmd1[58]) );
  COND1XL U2027 ( .A(n1773), .B(n1644), .C(n1643), .Z(acc_cmd1[32]) );
  COND1XL U2028 ( .A(n1773), .B(n1544), .C(n1543), .Z(acc_cmd1[57]) );
  COND1XL U2029 ( .A(n1773), .B(n1548), .C(n1547), .Z(acc_cmd1[56]) );
  COND1XL U2030 ( .A(n1773), .B(n1552), .C(n1551), .Z(acc_cmd1[55]) );
  COND1XL U2031 ( .A(n1773), .B(n1608), .C(n1607), .Z(acc_cmd1[41]) );
  COND1XL U2032 ( .A(n1773), .B(n1744), .C(n1743), .Z(acc_cmd1[7]) );
  COND1XL U2033 ( .A(n1773), .B(n1648), .C(n1647), .Z(acc_cmd1[31]) );
  COND1XL U2034 ( .A(n1773), .B(n1532), .C(n1531), .Z(acc_cmd1[60]) );
  COND1XL U2035 ( .A(n1773), .B(n1536), .C(n1535), .Z(acc_cmd1[59]) );
  COND1XL U2036 ( .A(n1773), .B(n1760), .C(n1759), .Z(acc_cmd1[3]) );
  COND1XL U2037 ( .A(n1773), .B(n1768), .C(n1767), .Z(acc_cmd1[1]) );
  COND1XL U2038 ( .A(n1773), .B(n1528), .C(n1527), .Z(acc_cmd1[61]) );
  COND1XL U2039 ( .A(n1773), .B(n1524), .C(n1523), .Z(acc_cmd1[62]) );
  COND1XL U2040 ( .A(n2408), .B(n2392), .C(n2391), .Z(n2433) );
  CNIVX1 U2041 ( .A(pushin), .Z(n1500) );
  CNIVX1 U2042 ( .A(pushin), .Z(n1499) );
  COND1XL U2043 ( .A(n2453), .B(n2452), .C(n1484), .Z(n2454) );
  CNIVX1 U2044 ( .A(pushin), .Z(n1498) );
  CNIVX1 U2045 ( .A(pushin), .Z(n1497) );
  CNIVX1 U2046 ( .A(pushin), .Z(n1496) );
  COND1XL U2047 ( .A(n795), .B(n2345), .C(n2344), .Z(n605) );
  COND1XL U2048 ( .A(n795), .B(n2403), .C(n2402), .Z(n609) );
  COND1XL U2049 ( .A(n795), .B(n2293), .C(n2292), .Z(n601) );
  COND1XL U2050 ( .A(n795), .B(n2332), .C(n2331), .Z(n604) );
  COND1XL U2051 ( .A(n795), .B(n2358), .C(n2357), .Z(n606) );
  COND1XL U2052 ( .A(n795), .B(n809), .C(n2374), .Z(n607) );
  COND1XL U2053 ( .A(n795), .B(n2389), .C(n2388), .Z(n608) );
  COND1XL U2054 ( .A(n795), .B(n2425), .C(n2424), .Z(n610) );
  COND1XL U2055 ( .A(n1490), .B(n2230), .C(n2229), .Z(n596) );
  COND1XL U2056 ( .A(n795), .B(n2242), .C(n2241), .Z(n597) );
  COND1XL U2057 ( .A(n795), .B(n2254), .C(n2253), .Z(n598) );
  COND1XL U2058 ( .A(n795), .B(n2267), .C(n2266), .Z(n599) );
  COND1XL U2059 ( .A(n1490), .B(n2280), .C(n2279), .Z(n600) );
  COND1XL U2060 ( .A(n795), .B(n2306), .C(n2305), .Z(n602) );
  COND1XL U2061 ( .A(n795), .B(n2319), .C(n2318), .Z(n603) );
  CNIVX1 U2062 ( .A(pushin), .Z(n1501) );
  CND3XL U2063 ( .A(cmd0[1]), .B(n2466), .C(push0), .Z(n215) );
  CAN2X1 U2064 ( .A(n12), .B(push0_2), .Z(n1357) );
  CNR3XL U2065 ( .A(n2467), .B(n1212), .C(n1214), .Z(cmd0_en_0) );
  CNR3XL U2066 ( .A(n2466), .B(n1212), .C(n2467), .Z(cmd1_en_0) );
  CNR2X1 U2067 ( .A(cmd0_2[0]), .B(cmd0_2[1]), .Z(n12) );
  CMX2XL U2068 ( .A0(q0[30]), .A1(q[30]), .S(n1496), .Z(n688) );
  CMX2XL U2069 ( .A0(n1245), .A1(q[17]), .S(n1497), .Z(n675) );
  CMX2XL U2070 ( .A0(n1246), .A1(q[25]), .S(n1496), .Z(n683) );
  CMX2XL U2071 ( .A0(n1250), .A1(q[3]), .S(n1498), .Z(n661) );
  CMX2XL U2072 ( .A0(n1254), .A1(q[19]), .S(n1497), .Z(n677) );
  CMX2XL U2073 ( .A0(n790), .A1(q[5]), .S(n1498), .Z(n663) );
  CMX2XL U2074 ( .A0(n1244), .A1(q[15]), .S(n1497), .Z(n673) );
  CMX2XL U2075 ( .A0(n1359), .A1(q[23]), .S(n1496), .Z(n681) );
  CMX2XL U2076 ( .A0(n1358), .A1(q[7]), .S(n1498), .Z(n665) );
  CMX2XL U2077 ( .A0(n1252), .A1(q[21]), .S(n1496), .Z(n679) );
  CMX2XL U2078 ( .A0(n1242), .A1(q[29]), .S(n1496), .Z(n687) );
  CMX2XL U2079 ( .A0(n1248), .A1(q[1]), .S(n1498), .Z(n659) );
  CMX2XL U2080 ( .A0(n1253), .A1(q[13]), .S(n1497), .Z(n671) );
  CIVX8 U2081 ( .A(cmd0_en_2_d), .Z(n2408) );
  CIVX1 U2082 ( .A(cmd0_en_2), .Z(n1363) );
  CIVX1 U2083 ( .A(cmd0_en_2), .Z(n1364) );
  CIVX1 U2084 ( .A(cmd0_en_2), .Z(n1365) );
  CIVX1 U2085 ( .A(cmd0_en_2), .Z(n1366) );
  CIVX1 U2086 ( .A(cmd0_en_2), .Z(n1367) );
  CIVXL U2087 ( .A(n1362), .Z(n1368) );
  CIVX1 U2088 ( .A(n1363), .Z(n1369) );
  CIVX1 U2089 ( .A(n1363), .Z(n1370) );
  CIVX1 U2090 ( .A(n1363), .Z(n1371) );
  CIVX1 U2091 ( .A(n1363), .Z(n1372) );
  CIVX1 U2092 ( .A(n1363), .Z(n1373) );
  CIVX1 U2093 ( .A(n1364), .Z(n1374) );
  CIVX1 U2094 ( .A(n1364), .Z(n1375) );
  CIVX1 U2095 ( .A(n1364), .Z(n1376) );
  CIVX1 U2096 ( .A(n1364), .Z(n1377) );
  CIVX1 U2097 ( .A(n1364), .Z(n1378) );
  CIVX1 U2098 ( .A(n1365), .Z(n1379) );
  CIVX1 U2099 ( .A(n1365), .Z(n1380) );
  CIVX1 U2100 ( .A(n1365), .Z(n1381) );
  CIVX1 U2101 ( .A(n1365), .Z(n1382) );
  CIVX1 U2102 ( .A(n1365), .Z(n1383) );
  CIVX1 U2103 ( .A(n1366), .Z(n1384) );
  CIVX1 U2104 ( .A(n1366), .Z(n1385) );
  CIVX1 U2105 ( .A(n1366), .Z(n1386) );
  CIVX1 U2106 ( .A(n1366), .Z(n1387) );
  CIVX1 U2107 ( .A(n1366), .Z(n1388) );
  CIVXL U2108 ( .A(n1367), .Z(n1389) );
  CIVX1 U2109 ( .A(n1367), .Z(n1390) );
  CIVX1 U2110 ( .A(n1367), .Z(n1391) );
  CIVX1 U2111 ( .A(n1367), .Z(n1392) );
  CIVX1 U2112 ( .A(n1367), .Z(n1393) );
  CIVX1 U2113 ( .A(n1366), .Z(n1394) );
  CIVX1 U2114 ( .A(cmd1_en_2), .Z(n1396) );
  CIVX1 U2115 ( .A(cmd1_en_2), .Z(n1397) );
  CIVX1 U2116 ( .A(cmd1_en_2), .Z(n1398) );
  CIVX1 U2117 ( .A(cmd1_en_2), .Z(n1399) );
  CIVX1 U2118 ( .A(cmd1_en_2), .Z(n1401) );
  CIVX2 U2119 ( .A(n792), .Z(n1402) );
  CIVXL U2120 ( .A(n792), .Z(n1403) );
  CIVXL U2121 ( .A(n792), .Z(n1404) );
  CIVXL U2122 ( .A(n792), .Z(n1405) );
  CIVXL U2123 ( .A(n792), .Z(n1406) );
  CIVX1 U2124 ( .A(n1396), .Z(n1407) );
  CIVX1 U2125 ( .A(n1396), .Z(n1408) );
  CIVX1 U2126 ( .A(n1396), .Z(n1409) );
  CIVX1 U2127 ( .A(n1396), .Z(n1410) );
  CIVX1 U2128 ( .A(n1396), .Z(n1411) );
  CIVX1 U2129 ( .A(n1397), .Z(n1412) );
  CIVX1 U2130 ( .A(n1397), .Z(n1413) );
  CIVX1 U2131 ( .A(n1397), .Z(n1414) );
  CIVX1 U2132 ( .A(n1397), .Z(n1415) );
  CIVX1 U2133 ( .A(n1397), .Z(n1416) );
  CIVX1 U2134 ( .A(n1398), .Z(n1417) );
  CIVX1 U2135 ( .A(n1398), .Z(n1418) );
  CIVX1 U2136 ( .A(n1398), .Z(n1419) );
  CIVX1 U2137 ( .A(n1398), .Z(n1420) );
  CIVX1 U2138 ( .A(n1398), .Z(n1421) );
  CIVX1 U2139 ( .A(n1399), .Z(n1422) );
  CIVX1 U2140 ( .A(n1399), .Z(n1423) );
  CIVX1 U2141 ( .A(n1399), .Z(n1424) );
  CIVX1 U2142 ( .A(n1399), .Z(n1425) );
  CIVXL U2143 ( .A(n1399), .Z(n1426) );
  CIVX1 U2144 ( .A(n1400), .Z(n1427) );
  CIVX1 U2145 ( .A(n1400), .Z(n1428) );
  CIVXL U2146 ( .A(n1400), .Z(n1429) );
  CIVX1 U2147 ( .A(n1400), .Z(n1430) );
  CIVX1 U2148 ( .A(n1400), .Z(n1431) );
  CIVX1 U2149 ( .A(n1401), .Z(n1432) );
  CIVX1 U2150 ( .A(n1401), .Z(n1433) );
  CIVXL U2151 ( .A(n1401), .Z(n1434) );
  CIVXL U2152 ( .A(n1401), .Z(n1435) );
  CIVXL U2153 ( .A(n1401), .Z(n1436) );
  CIVXL U2154 ( .A(n1488), .Z(n1487) );
  CIVX1 U2155 ( .A(h0_1[4]), .Z(n1488) );
  CIVXL U2156 ( .A(n1203), .Z(n1489) );
  CIVX2 U2157 ( .A(cmd0_2[1]), .Z(n2463) );
  CIVX2 U2158 ( .A(cmd0_2[0]), .Z(n2464) );
  CMX2X1 U2159 ( .A0(n1243), .A1(q[28]), .S(n1496), .Z(n686) );
  CMX2X1 U2160 ( .A0(n1360), .A1(q[27]), .S(n1496), .Z(n685) );
  CMX2X1 U2161 ( .A0(q0[26]), .A1(q[26]), .S(n1496), .Z(n684) );
  CMX2X1 U2162 ( .A0(q0[22]), .A1(q[22]), .S(n1496), .Z(n680) );
  CMX2X1 U2163 ( .A0(q0[16]), .A1(q[16]), .S(n1497), .Z(n674) );
  CMX2X1 U2164 ( .A0(q0[10]), .A1(q[10]), .S(n1497), .Z(n668) );
  CMX2X1 U2165 ( .A0(n1249), .A1(q[6]), .S(n1498), .Z(n664) );
  CMX2X1 U2166 ( .A0(q0[2]), .A1(q[2]), .S(n1498), .Z(n660) );
  CMX2X1 U2167 ( .A0(q0[0]), .A1(q[0]), .S(n1498), .Z(n658) );
  CMX2X1 U2168 ( .A0(h0[30]), .A1(h[30]), .S(n1498), .Z(n656) );
  CMX2X1 U2169 ( .A0(h0[29]), .A1(h[29]), .S(n1498), .Z(n655) );
  CMX2X1 U2170 ( .A0(h0[28]), .A1(h[28]), .S(n1498), .Z(n654) );
  CMX2X1 U2171 ( .A0(h0[26]), .A1(h[26]), .S(n1499), .Z(n652) );
  CMX2X1 U2172 ( .A0(h0[23]), .A1(h[23]), .S(n1499), .Z(n649) );
  CMX2X1 U2173 ( .A0(h0[19]), .A1(h[19]), .S(n1499), .Z(n645) );
  CMX2X1 U2174 ( .A0(h0[14]), .A1(h[14]), .S(n1500), .Z(n640) );
  CMX2X1 U2175 ( .A0(h0[13]), .A1(h[13]), .S(n1500), .Z(n639) );
  CMX2X1 U2176 ( .A0(h0[11]), .A1(h[11]), .S(n1500), .Z(n637) );
  CMX2X1 U2177 ( .A0(n1251), .A1(h[8]), .S(n1500), .Z(n634) );
  CMX2X1 U2178 ( .A0(h0[1]), .A1(h[1]), .S(n1501), .Z(n617) );
  CMX2X1 U2179 ( .A0(n1203), .A1(h[0]), .S(n1501), .Z(n614) );
  CMX2X1 U2180 ( .A0(cmd0_en_1), .A1(n1368), .S(rst), .Z(n755) );
  CIVX2 U2181 ( .A(n215), .Z(n2465) );
  CIVX2 U2182 ( .A(cmd2_en_1), .Z(n1502) );
  CMXI2X1 U2183 ( .A0(n1502), .A1(n794), .S(rst), .Z(n690) );
  CMXI2X1 U2184 ( .A0(n1503), .A1(n1504), .S(n215), .Z(n631) );
  CMXI2X1 U2185 ( .A0(n2033), .A1(n1504), .S(cmd2_en_1), .Z(n630) );
  CMXI2X1 U2186 ( .A0(n1505), .A1(n1506), .S(n215), .Z(n628) );
  CMXI2X1 U2187 ( .A0(n2426), .A1(n1506), .S(cmd2_en_1), .Z(n627) );
  CMXI2X1 U2188 ( .A0(n1507), .A1(n1508), .S(n215), .Z(n625) );
  CMXI2X1 U2189 ( .A0(n1488), .A1(n1508), .S(cmd2_en_1), .Z(n624) );
  CIVX2 U2190 ( .A(h0[1]), .Z(n1509) );
  CMXI2X1 U2191 ( .A0(n1509), .A1(n1510), .S(n215), .Z(n616) );
  CIVX2 U2192 ( .A(h0_1[1]), .Z(n1792) );
  CMXI2X1 U2193 ( .A0(n1792), .A1(n1510), .S(cmd2_en_1), .Z(n615) );
  CIVX2 U2194 ( .A(h0_0[0]), .Z(n1511) );
  CIVX2 U2195 ( .A(h0_1[0]), .Z(n1793) );
  CMXI2X1 U2196 ( .A0(n1793), .A1(n1511), .S(cmd2_en_1), .Z(n612) );
  CMXI2X1 U2197 ( .A0(n1512), .A1(n1513), .S(n215), .Z(n619) );
  CMXI2X1 U2198 ( .A0(n1864), .A1(n1513), .S(cmd2_en_1), .Z(n618) );
  CMX2X1 U2199 ( .A0(cmd1_en_1), .A1(n1402), .S(rst), .Z(n756) );
  CIVX2 U2200 ( .A(cmd1_en_2_d), .Z(n1778) );
  CND2X1 U2201 ( .A(n1426), .B(n1778), .Z(n1514) );
  CND2X1 U2202 ( .A(n1773), .B(n2408), .Z(n1515) );
  CND2X1 U2203 ( .A(n1773), .B(cmd0_en_2_d), .Z(n1516) );
  CMX2X1 U2204 ( .A0(out1_2[62]), .A1(N271), .S(n1403), .Z(n421) );
  CND2X1 U2205 ( .A(cmd0_2[1]), .B(n2464), .Z(n2460) );
  CIVX2 U2206 ( .A(n2460), .Z(n1519) );
  CANR2X1 U2207 ( .A(out0_2[62]), .B(n1357), .C(N480), .D(n1298), .Z(n1522) );
  CND2X1 U2208 ( .A(cmd0_2[0]), .B(n2463), .Z(n2459) );
  CIVX2 U2209 ( .A(n2459), .Z(n1520) );
  CANR2X1 U2210 ( .A(out1_2[62]), .B(n1299), .C(acc[62]), .D(n2461), .Z(n1521)
         );
  CMX2X1 U2211 ( .A0(out1_2[61]), .A1(N270), .S(n1404), .Z(n423) );
  CND2X1 U2212 ( .A(n1526), .B(n1525), .Z(n422) );
  CMX2X1 U2213 ( .A0(out1_2[60]), .A1(N269), .S(n1405), .Z(n425) );
  CND2X1 U2214 ( .A(n1530), .B(n1529), .Z(n424) );
  CMX2X1 U2215 ( .A0(out1_2[59]), .A1(N268), .S(n1406), .Z(n427) );
  CANR2X1 U2216 ( .A(out0_2[59]), .B(n1357), .C(N477), .D(n1298), .Z(n1534) );
  CND2X1 U2217 ( .A(n1534), .B(n1533), .Z(n426) );
  CMX2X1 U2218 ( .A0(out1_2[58]), .A1(N267), .S(n1407), .Z(n429) );
  CANR2X1 U2219 ( .A(out0_2[58]), .B(n1357), .C(N476), .D(n1298), .Z(n1538) );
  CND2X1 U2220 ( .A(n1538), .B(n1537), .Z(n428) );
  CMX2X1 U2221 ( .A0(out1_2[57]), .A1(N266), .S(n1408), .Z(n431) );
  CND2X1 U2222 ( .A(n1542), .B(n1541), .Z(n430) );
  CMX2X1 U2223 ( .A0(out1_2[56]), .A1(N265), .S(n1409), .Z(n433) );
  CANR2X1 U2224 ( .A(out0_2[56]), .B(n1357), .C(N474), .D(n1298), .Z(n1546) );
  CND2X1 U2225 ( .A(n1546), .B(n1545), .Z(n432) );
  CMX2X1 U2226 ( .A0(out1_2[55]), .A1(N264), .S(n1410), .Z(n435) );
  CND2X1 U2227 ( .A(n1550), .B(n1549), .Z(n434) );
  CMX2X1 U2228 ( .A0(out1_2[54]), .A1(N263), .S(n1411), .Z(n437) );
  CANR2X1 U2229 ( .A(out0_2[54]), .B(n1357), .C(N472), .D(n1298), .Z(n1554) );
  CND2X1 U2230 ( .A(n1554), .B(n1553), .Z(n436) );
  CMX2X1 U2231 ( .A0(out1_2[53]), .A1(N262), .S(n1412), .Z(n439) );
  CND2X1 U2232 ( .A(n1558), .B(n1557), .Z(n438) );
  CMX2X1 U2233 ( .A0(out1_2[52]), .A1(N261), .S(n1413), .Z(n441) );
  CANR2X1 U2234 ( .A(out0_2[52]), .B(n1357), .C(N470), .D(n1298), .Z(n1562) );
  CND2X1 U2235 ( .A(n1562), .B(n1561), .Z(n440) );
  CMX2X1 U2236 ( .A0(out1_2[51]), .A1(N260), .S(n1414), .Z(n443) );
  CND2X1 U2237 ( .A(n1566), .B(n1565), .Z(n442) );
  CMX2X1 U2238 ( .A0(out1_2[50]), .A1(N259), .S(n1415), .Z(n445) );
  CANR2X1 U2239 ( .A(out0_2[50]), .B(n1357), .C(N468), .D(n1298), .Z(n1570) );
  CND2X1 U2240 ( .A(n1570), .B(n1569), .Z(n444) );
  CMX2X1 U2241 ( .A0(out1_2[49]), .A1(N258), .S(n1416), .Z(n447) );
  CND2X1 U2242 ( .A(n1574), .B(n1573), .Z(n446) );
  CMX2X1 U2243 ( .A0(out1_2[48]), .A1(N257), .S(n1417), .Z(n449) );
  CANR2X1 U2244 ( .A(out0_2[48]), .B(n1357), .C(N466), .D(n1298), .Z(n1578) );
  CND2X1 U2245 ( .A(n1578), .B(n1577), .Z(n448) );
  CMX2X1 U2246 ( .A0(out1_2[47]), .A1(N256), .S(n1418), .Z(n451) );
  CND2X1 U2247 ( .A(n1582), .B(n1581), .Z(n450) );
  CMX2X1 U2248 ( .A0(out1_2[46]), .A1(N255), .S(n1419), .Z(n453) );
  CANR2X1 U2249 ( .A(out0_2[46]), .B(n1357), .C(N464), .D(n1298), .Z(n1586) );
  CND2X1 U2250 ( .A(n1586), .B(n1585), .Z(n452) );
  CMX2X1 U2251 ( .A0(out1_2[45]), .A1(N254), .S(n1420), .Z(n455) );
  CND2X1 U2252 ( .A(n1590), .B(n1589), .Z(n454) );
  CMX2X1 U2253 ( .A0(out1_2[44]), .A1(N253), .S(n1421), .Z(n457) );
  CANR2X1 U2254 ( .A(out0_2[44]), .B(n1357), .C(N462), .D(n1298), .Z(n1594) );
  CND2X1 U2255 ( .A(n1594), .B(n1593), .Z(n456) );
  CMX2X1 U2256 ( .A0(out1_2[43]), .A1(N252), .S(n1422), .Z(n459) );
  CND2X1 U2257 ( .A(n1598), .B(n1597), .Z(n458) );
  CMX2X1 U2258 ( .A0(out1_2[42]), .A1(N251), .S(n1423), .Z(n461) );
  CANR2X1 U2259 ( .A(out0_2[42]), .B(n1357), .C(N460), .D(n1298), .Z(n1602) );
  CND2X1 U2260 ( .A(n1602), .B(n1601), .Z(n460) );
  CMX2X1 U2261 ( .A0(out1_2[41]), .A1(N250), .S(n1424), .Z(n463) );
  CND2X1 U2262 ( .A(n1606), .B(n1605), .Z(n462) );
  CMX2X1 U2263 ( .A0(out1_2[40]), .A1(N249), .S(n1425), .Z(n465) );
  CND2X1 U2264 ( .A(n1610), .B(n1609), .Z(n464) );
  CMX2X1 U2265 ( .A0(out1_2[39]), .A1(N248), .S(n1426), .Z(n467) );
  CND2X1 U2266 ( .A(n1614), .B(n1613), .Z(n466) );
  CMX2X1 U2267 ( .A0(out1_2[38]), .A1(N247), .S(n1427), .Z(n469) );
  CANR2X1 U2268 ( .A(out0_2[38]), .B(n1357), .C(N456), .D(n1298), .Z(n1618) );
  CND2X1 U2269 ( .A(n1618), .B(n1617), .Z(n468) );
  CMX2X1 U2270 ( .A0(out1_2[37]), .A1(N246), .S(n1428), .Z(n471) );
  CND2X1 U2271 ( .A(n1622), .B(n1621), .Z(n470) );
  CMX2X1 U2272 ( .A0(out1_2[36]), .A1(N245), .S(n1429), .Z(n473) );
  CANR2X1 U2273 ( .A(out0_2[36]), .B(n1357), .C(N454), .D(n1298), .Z(n1626) );
  CND2X1 U2274 ( .A(n1626), .B(n1625), .Z(n472) );
  CMX2X1 U2275 ( .A0(out1_2[35]), .A1(N244), .S(n1430), .Z(n475) );
  CND2X1 U2276 ( .A(n1630), .B(n1629), .Z(n474) );
  CMX2X1 U2277 ( .A0(out1_2[34]), .A1(N243), .S(n1431), .Z(n477) );
  CND2X1 U2278 ( .A(n1634), .B(n1633), .Z(n476) );
  CMX2X1 U2279 ( .A0(out1_2[33]), .A1(N242), .S(n1431), .Z(n479) );
  CND2X1 U2280 ( .A(n1638), .B(n1637), .Z(n478) );
  CMX2X1 U2281 ( .A0(out1_2[32]), .A1(N241), .S(n1432), .Z(n481) );
  CND2X1 U2282 ( .A(n1642), .B(n1641), .Z(n480) );
  CMX2X1 U2283 ( .A0(out1_2[31]), .A1(N240), .S(n1433), .Z(n483) );
  CND2X1 U2284 ( .A(n1646), .B(n1645), .Z(n482) );
  CMX2X1 U2285 ( .A0(out1_2[30]), .A1(N239), .S(n1428), .Z(n485) );
  CANR2X1 U2286 ( .A(out0_2[30]), .B(n1357), .C(N448), .D(n1298), .Z(n1650) );
  CND2X1 U2287 ( .A(n1650), .B(n1649), .Z(n484) );
  CMX2X1 U2288 ( .A0(out1_2[29]), .A1(N238), .S(n1430), .Z(n487) );
  CND2X1 U2289 ( .A(n1654), .B(n1653), .Z(n486) );
  CMX2X1 U2290 ( .A0(out1_2[28]), .A1(N237), .S(n1427), .Z(n489) );
  CANR2X1 U2291 ( .A(out0_2[28]), .B(n1357), .C(N446), .D(n1298), .Z(n1658) );
  CND2X1 U2292 ( .A(n1658), .B(n1657), .Z(n488) );
  CMX2X1 U2293 ( .A0(out1_2[27]), .A1(N236), .S(n1432), .Z(n491) );
  CND2X1 U2294 ( .A(n1662), .B(n1661), .Z(n490) );
  CMX2X1 U2295 ( .A0(out1_2[26]), .A1(N235), .S(n1433), .Z(n493) );
  CND2X1 U2296 ( .A(n1666), .B(n1665), .Z(n492) );
  CMX2X1 U2297 ( .A0(out1_2[25]), .A1(N234), .S(n1434), .Z(n495) );
  CND2X1 U2298 ( .A(n1670), .B(n1669), .Z(n494) );
  CMX2X1 U2299 ( .A0(out1_2[24]), .A1(N233), .S(n1435), .Z(n497) );
  CND2X1 U2300 ( .A(n1674), .B(n1673), .Z(n496) );
  CMX2X1 U2301 ( .A0(out1_2[23]), .A1(N232), .S(n1436), .Z(n499) );
  CND2X1 U2302 ( .A(n1678), .B(n1677), .Z(n498) );
  CMX2X1 U2303 ( .A0(out1_2[22]), .A1(N231), .S(n1402), .Z(n501) );
  CANR2X1 U2304 ( .A(out0_2[22]), .B(n1357), .C(N440), .D(n1298), .Z(n1682) );
  CND2X1 U2305 ( .A(n1682), .B(n1681), .Z(n500) );
  CMX2X1 U2306 ( .A0(out1_2[21]), .A1(N230), .S(n1403), .Z(n503) );
  CANR2X1 U2307 ( .A(out1_2[21]), .B(n1299), .C(acc[21]), .D(n2461), .Z(n1685)
         );
  CND2X1 U2308 ( .A(n1686), .B(n1685), .Z(n502) );
  CIVX2 U2309 ( .A(out1_2[21]), .Z(n1688) );
  CMX2X1 U2310 ( .A0(out1_2[20]), .A1(N229), .S(n1404), .Z(n505) );
  CANR2X1 U2311 ( .A(out1_2[20]), .B(n1299), .C(acc[20]), .D(n2461), .Z(n1689)
         );
  CND2X1 U2312 ( .A(n1690), .B(n1689), .Z(n504) );
  CIVX2 U2313 ( .A(out1_2[20]), .Z(n1692) );
  CMX2X1 U2314 ( .A0(out1_2[19]), .A1(N228), .S(n1405), .Z(n507) );
  CANR2X1 U2315 ( .A(out1_2[19]), .B(n1299), .C(acc[19]), .D(n2461), .Z(n1693)
         );
  CND2X1 U2316 ( .A(n1694), .B(n1693), .Z(n506) );
  CIVX2 U2317 ( .A(out1_2[19]), .Z(n1696) );
  CMX2X1 U2318 ( .A0(out1_2[18]), .A1(N227), .S(n1406), .Z(n509) );
  CANR2X1 U2319 ( .A(out1_2[18]), .B(n1299), .C(acc[18]), .D(n2461), .Z(n1697)
         );
  CND2X1 U2320 ( .A(n1698), .B(n1697), .Z(n508) );
  CIVX2 U2321 ( .A(out1_2[18]), .Z(n1700) );
  CMX2X1 U2322 ( .A0(out1_2[17]), .A1(N226), .S(n1407), .Z(n511) );
  CANR2X1 U2323 ( .A(out1_2[17]), .B(n1299), .C(acc[17]), .D(n2461), .Z(n1701)
         );
  CND2X1 U2324 ( .A(n1702), .B(n1701), .Z(n510) );
  CIVX2 U2325 ( .A(out1_2[17]), .Z(n1704) );
  CANR2X1 U2326 ( .A(n1770), .B(acc[17]), .C(n1769), .D(out0_2[17]), .Z(n1703)
         );
  CMX2X1 U2327 ( .A0(out1_2[16]), .A1(N225), .S(n1408), .Z(n513) );
  CND2X1 U2328 ( .A(n1706), .B(n1705), .Z(n512) );
  CMX2X1 U2329 ( .A0(out1_2[15]), .A1(N224), .S(n1409), .Z(n515) );
  CND2X1 U2330 ( .A(n1710), .B(n1709), .Z(n514) );
  CMX2X1 U2331 ( .A0(out1_2[14]), .A1(N223), .S(n1410), .Z(n517) );
  CND2X1 U2332 ( .A(n1714), .B(n1713), .Z(n516) );
  CMX2X1 U2333 ( .A0(out1_2[13]), .A1(N222), .S(n1411), .Z(n519) );
  CND2X1 U2334 ( .A(n1718), .B(n1717), .Z(n518) );
  CMX2X1 U2335 ( .A0(out1_2[12]), .A1(N221), .S(n1412), .Z(n521) );
  CND2X1 U2336 ( .A(n1722), .B(n1721), .Z(n520) );
  CMX2X1 U2337 ( .A0(out1_2[11]), .A1(N220), .S(n1413), .Z(n523) );
  CND2X1 U2338 ( .A(n1726), .B(n1725), .Z(n522) );
  CMX2X1 U2339 ( .A0(out1_2[10]), .A1(N219), .S(n1414), .Z(n525) );
  CND2X1 U2340 ( .A(n1730), .B(n1729), .Z(n524) );
  CMX2X1 U2341 ( .A0(out1_2[9]), .A1(N218), .S(n1415), .Z(n527) );
  CND2X1 U2342 ( .A(n1734), .B(n1733), .Z(n526) );
  CANR2X1 U2343 ( .A(n1770), .B(acc[9]), .C(n1769), .D(out0_2[9]), .Z(n1735)
         );
  CMX2X1 U2344 ( .A0(out1_2[8]), .A1(N217), .S(n1416), .Z(n529) );
  CND2X1 U2345 ( .A(n1738), .B(n1737), .Z(n528) );
  CMX2X1 U2346 ( .A0(out1_2[7]), .A1(N216), .S(n1417), .Z(n531) );
  CND2X1 U2347 ( .A(n1742), .B(n1741), .Z(n530) );
  CMX2X1 U2348 ( .A0(out1_2[6]), .A1(N215), .S(n1418), .Z(n533) );
  CND2X1 U2349 ( .A(n1746), .B(n1745), .Z(n532) );
  CMX2X1 U2350 ( .A0(out1_2[5]), .A1(N214), .S(n1419), .Z(n535) );
  CND2X1 U2351 ( .A(n1750), .B(n1749), .Z(n534) );
  CMX2X1 U2352 ( .A0(out1_2[4]), .A1(N213), .S(n1420), .Z(n537) );
  CANR2X1 U2353 ( .A(out1_2[4]), .B(n1299), .C(acc[4]), .D(n2461), .Z(n1753)
         );
  CND2X1 U2354 ( .A(n1754), .B(n1753), .Z(n536) );
  CIVX2 U2355 ( .A(out1_2[4]), .Z(n1756) );
  CMX2X1 U2356 ( .A0(out1_2[3]), .A1(N212), .S(n1421), .Z(n539) );
  CANR2X1 U2357 ( .A(out1_2[3]), .B(n1299), .C(acc[3]), .D(n2461), .Z(n1757)
         );
  CND2X1 U2358 ( .A(n1758), .B(n1757), .Z(n538) );
  CIVX2 U2359 ( .A(out1_2[3]), .Z(n1760) );
  CMX2X1 U2360 ( .A0(out1_2[2]), .A1(N211), .S(n1422), .Z(n541) );
  CANR2X1 U2361 ( .A(out1_2[2]), .B(n1299), .C(acc[2]), .D(n2461), .Z(n1761)
         );
  CND2X1 U2362 ( .A(n1762), .B(n1761), .Z(n540) );
  CIVX2 U2363 ( .A(out1_2[2]), .Z(n1764) );
  CMX2X1 U2364 ( .A0(out1_2[1]), .A1(N210), .S(n1423), .Z(n543) );
  CANR2X1 U2365 ( .A(out1_2[1]), .B(n1299), .C(acc[1]), .D(n2461), .Z(n1765)
         );
  CND2X1 U2366 ( .A(n1766), .B(n1765), .Z(n542) );
  CIVX2 U2367 ( .A(out1_2[1]), .Z(n1768) );
  CMX2X1 U2368 ( .A0(out1_2[0]), .A1(N209), .S(n1424), .Z(n545) );
  CIVX2 U2369 ( .A(out1_2[0]), .Z(n1772) );
  CMX2X1 U2370 ( .A0(out1_2[63]), .A1(N272), .S(n1425), .Z(n419) );
  CANR2X1 U2371 ( .A(out0_2[63]), .B(n1357), .C(N481), .D(n1298), .Z(n1775) );
  CANR2X1 U2372 ( .A(out1_2[63]), .B(n1299), .C(acc[63]), .D(n2461), .Z(n1774)
         );
  CND2X1 U2373 ( .A(n1775), .B(n1774), .Z(n546) );
  CIVX2 U2374 ( .A(h0_0[3]), .Z(n1777) );
  CND2X1 U2375 ( .A(n1792), .B(n1793), .Z(n1789) );
  CIVX2 U2376 ( .A(out0_2[63]), .Z(n1780) );
  CANR2X1 U2377 ( .A(acc[63]), .B(n1257), .C(out1_2[63]), .D(n1297), .Z(n1779)
         );
  CND2X1 U2378 ( .A(n1293), .B(n1861), .Z(n1895) );
  COND2X1 U2379 ( .A(n1895), .B(n1887), .C(n795), .D(n1781), .Z(n547) );
  CIVX2 U2380 ( .A(out0_2[62]), .Z(n1783) );
  CIVX2 U2381 ( .A(n1806), .Z(n1797) );
  CMXI2X1 U2382 ( .A0(n1301), .A1(n1797), .S(h0_1[0]), .Z(n1784) );
  CND2X1 U2383 ( .A(n1784), .B(n1792), .Z(n2043) );
  CND2X1 U2384 ( .A(n1864), .B(n1861), .Z(n1853) );
  CND2X1 U2385 ( .A(n2212), .B(n2207), .Z(n1801) );
  CIVX2 U2386 ( .A(out2_2[62]), .Z(n1785) );
  COND2X1 U2387 ( .A(n2043), .B(n1801), .C(n1490), .D(n1785), .Z(n548) );
  CIVX2 U2388 ( .A(out0_2[61]), .Z(n1787) );
  CND2X1 U2389 ( .A(h0_1[1]), .B(h0_1[0]), .Z(n1794) );
  CANR2X1 U2390 ( .A(n1301), .B(h0_1[0]), .C(n1797), .D(h0_1[1]), .Z(n1788) );
  COND3X1 U2391 ( .A(n1789), .B(n1791), .C(n1794), .D(n1788), .Z(n2056) );
  COND2X1 U2392 ( .A(n2056), .B(n1801), .C(n1490), .D(n1790), .Z(n549) );
  CIVX2 U2393 ( .A(n1791), .Z(n1811) );
  CND2X1 U2394 ( .A(h0_1[0]), .B(n1792), .Z(n2435) );
  CND2X1 U2395 ( .A(h0_1[1]), .B(n1793), .Z(n2437) );
  CANR2X1 U2396 ( .A(n1811), .B(n2406), .C(n1301), .D(n2405), .Z(n1799) );
  CIVX2 U2397 ( .A(out0_2[60]), .Z(n1796) );
  CANR2X1 U2398 ( .A(n1797), .B(n2441), .C(n1326), .D(n2410), .Z(n1798) );
  CND2X1 U2399 ( .A(n1799), .B(n1798), .Z(n2069) );
  COND2X1 U2400 ( .A(n2069), .B(n1801), .C(n795), .D(n1800), .Z(n550) );
  CANR2X1 U2401 ( .A(n1326), .B(n2406), .C(n1811), .D(n2405), .Z(n1805) );
  CIVX2 U2402 ( .A(out0_2[59]), .Z(n1803) );
  CANR2X1 U2403 ( .A(n1301), .B(n2441), .C(n1316), .D(n2410), .Z(n1804) );
  CND2X1 U2404 ( .A(n1805), .B(n1804), .Z(n1892) );
  CMXI2X1 U2405 ( .A0(n1892), .A1(n1807), .S(h0_1[2]), .Z(n1862) );
  CND2X1 U2406 ( .A(n1862), .B(n1861), .Z(n1932) );
  COND2X1 U2407 ( .A(n1887), .B(n1932), .C(n795), .D(n1808), .Z(n551) );
  CANR2X1 U2408 ( .A(n1316), .B(n2406), .C(n1326), .D(n2405), .Z(n1813) );
  CIVX2 U2409 ( .A(out0_2[58]), .Z(n1810) );
  CANR2X1 U2410 ( .A(n1811), .B(n2441), .C(n1345), .D(n2410), .Z(n1812) );
  CND2X1 U2411 ( .A(n1813), .B(n1812), .Z(n1901) );
  CMXI2X1 U2412 ( .A0(n1901), .A1(n2043), .S(h0_1[2]), .Z(n1814) );
  CND2X1 U2413 ( .A(n1814), .B(n1861), .Z(n1941) );
  COND2X1 U2414 ( .A(n1887), .B(n1941), .C(n1490), .D(n1815), .Z(n552) );
  CANR2X1 U2415 ( .A(n1345), .B(n2406), .C(n1316), .D(n2405), .Z(n1819) );
  CIVX2 U2416 ( .A(out0_2[57]), .Z(n1817) );
  CANR2X1 U2417 ( .A(n1326), .B(n2441), .C(n1344), .D(n2410), .Z(n1818) );
  CND2X1 U2418 ( .A(n1819), .B(n1818), .Z(n1910) );
  CMXI2X1 U2419 ( .A0(n1910), .A1(n2056), .S(h0_1[2]), .Z(n1820) );
  CND2X1 U2420 ( .A(n1820), .B(n1861), .Z(n1950) );
  COND2X1 U2421 ( .A(n1887), .B(n1950), .C(n1490), .D(n1821), .Z(n553) );
  CANR2X1 U2422 ( .A(n1344), .B(n2406), .C(n1345), .D(n2405), .Z(n1825) );
  CIVX2 U2423 ( .A(out0_2[56]), .Z(n1823) );
  CANR2X1 U2424 ( .A(n1316), .B(n2441), .C(n1346), .D(n2410), .Z(n1824) );
  CND2X1 U2425 ( .A(n1825), .B(n1824), .Z(n1919) );
  CMXI2X1 U2426 ( .A0(n1919), .A1(n2069), .S(h0_1[2]), .Z(n1826) );
  CND2X1 U2427 ( .A(n1826), .B(n1861), .Z(n1959) );
  COND2X1 U2428 ( .A(n1887), .B(n1959), .C(n1490), .D(n1827), .Z(n554) );
  CANR2X1 U2429 ( .A(n1346), .B(n2406), .C(n1344), .D(n2405), .Z(n1831) );
  CIVX2 U2430 ( .A(out0_2[55]), .Z(n1829) );
  CANR2X1 U2431 ( .A(n1345), .B(n2441), .C(n1343), .D(n2410), .Z(n1830) );
  CND2X1 U2432 ( .A(n1831), .B(n1830), .Z(n1929) );
  CANR2X1 U2433 ( .A(n1295), .B(n1892), .C(n2207), .D(n1929), .Z(n1832) );
  COND2X1 U2434 ( .A(n1887), .B(n1968), .C(n1490), .D(n1833), .Z(n555) );
  CANR2X1 U2435 ( .A(n1343), .B(n2406), .C(n1346), .D(n2405), .Z(n1837) );
  CIVX2 U2436 ( .A(out0_2[54]), .Z(n1835) );
  CANR2X1 U2437 ( .A(n1344), .B(n2441), .C(n1348), .D(n2410), .Z(n1836) );
  CND2X1 U2438 ( .A(n1837), .B(n1836), .Z(n1938) );
  CIVX2 U2439 ( .A(n1938), .Z(n1839) );
  CANR2X1 U2440 ( .A(h0_1[2]), .B(n1901), .C(h0_1[3]), .D(n2043), .Z(n1838) );
  COND3X1 U2441 ( .A(n1839), .B(n1853), .C(n1865), .D(n1838), .Z(n1977) );
  COND2X1 U2442 ( .A(n1887), .B(n1977), .C(n1490), .D(n1840), .Z(n556) );
  CANR2X1 U2443 ( .A(n1348), .B(n2406), .C(n1343), .D(n2405), .Z(n1844) );
  CIVX2 U2444 ( .A(out0_2[53]), .Z(n1842) );
  CANR2X1 U2445 ( .A(n1346), .B(n2441), .C(n1338), .D(n2410), .Z(n1843) );
  CND2X1 U2446 ( .A(n1844), .B(n1843), .Z(n1947) );
  CIVX2 U2447 ( .A(n1947), .Z(n1846) );
  CANR2X1 U2448 ( .A(h0_1[2]), .B(n1910), .C(h0_1[3]), .D(n2056), .Z(n1845) );
  COND3X1 U2449 ( .A(n1846), .B(n1853), .C(n1865), .D(n1845), .Z(n1986) );
  COND2X1 U2450 ( .A(n1887), .B(n1986), .C(n1490), .D(n1847), .Z(n557) );
  CANR2X1 U2451 ( .A(n1338), .B(n2406), .C(n1348), .D(n2405), .Z(n1851) );
  CIVX2 U2452 ( .A(out0_2[52]), .Z(n1849) );
  CANR2X1 U2453 ( .A(n1343), .B(n2441), .C(n1349), .D(n2410), .Z(n1850) );
  CND2X1 U2454 ( .A(n1851), .B(n1850), .Z(n1956) );
  CIVX2 U2455 ( .A(n1956), .Z(n1854) );
  CANR2X1 U2456 ( .A(h0_1[2]), .B(n1919), .C(h0_1[3]), .D(n2069), .Z(n1852) );
  COND3X1 U2457 ( .A(n1854), .B(n1853), .C(n1865), .D(n1852), .Z(n1995) );
  COND2X1 U2458 ( .A(n1887), .B(n1995), .C(n1490), .D(n1855), .Z(n558) );
  CANR2X1 U2459 ( .A(n1349), .B(n2406), .C(n1338), .D(n2405), .Z(n1859) );
  CIVX2 U2460 ( .A(out0_2[51]), .Z(n1857) );
  CANR2X1 U2461 ( .A(n1348), .B(n2441), .C(n1337), .D(n2410), .Z(n1858) );
  CND2X1 U2462 ( .A(n1859), .B(n1858), .Z(n1965) );
  CANR2X1 U2463 ( .A(n1295), .B(n1929), .C(n2207), .D(n1965), .Z(n1860) );
  COND2X1 U2464 ( .A(n1887), .B(n2004), .C(n1490), .D(n1863), .Z(n559) );
  CANR2X1 U2465 ( .A(n1296), .B(n1901), .C(n1295), .D(n1938), .Z(n1871) );
  CANR2X1 U2466 ( .A(n1337), .B(n2406), .C(n1349), .D(n2405), .Z(n1869) );
  CIVX2 U2467 ( .A(out0_2[50]), .Z(n1867) );
  CANR2X1 U2468 ( .A(n1338), .B(n2441), .C(n1350), .D(n2410), .Z(n1868) );
  CND2X1 U2469 ( .A(n1869), .B(n1868), .Z(n1974) );
  CANR2X1 U2470 ( .A(n2218), .B(n2043), .C(n2207), .D(n1974), .Z(n1870) );
  CND2X1 U2471 ( .A(n1871), .B(n1870), .Z(n2013) );
  COND2X1 U2472 ( .A(n1887), .B(n2013), .C(n1490), .D(n1872), .Z(n560) );
  CANR2X1 U2473 ( .A(n1296), .B(n1910), .C(n1295), .D(n1947), .Z(n1878) );
  CANR2X1 U2474 ( .A(n1350), .B(n2406), .C(n1337), .D(n2405), .Z(n1876) );
  CIVX2 U2475 ( .A(out0_2[49]), .Z(n1874) );
  CANR2X1 U2476 ( .A(n1349), .B(n2441), .C(n1336), .D(n2410), .Z(n1875) );
  CND2X1 U2477 ( .A(n1876), .B(n1875), .Z(n1983) );
  CANR2X1 U2478 ( .A(n2218), .B(n2056), .C(n2207), .D(n1983), .Z(n1877) );
  CND2X1 U2479 ( .A(n1878), .B(n1877), .Z(n2022) );
  COND2X1 U2480 ( .A(n1887), .B(n2022), .C(n1490), .D(n1879), .Z(n561) );
  CANR2X1 U2481 ( .A(n1296), .B(n1919), .C(n1295), .D(n1956), .Z(n1885) );
  CANR2X1 U2482 ( .A(n1336), .B(n2406), .C(n1350), .D(n2405), .Z(n1883) );
  CIVX2 U2483 ( .A(out0_2[48]), .Z(n1881) );
  CANR2X1 U2484 ( .A(n1337), .B(n2441), .C(n1351), .D(n2410), .Z(n1882) );
  CND2X1 U2485 ( .A(n1883), .B(n1882), .Z(n1992) );
  CANR2X1 U2486 ( .A(n2218), .B(n2069), .C(n2207), .D(n1992), .Z(n1884) );
  CND2X1 U2487 ( .A(n1885), .B(n1884), .Z(n2031) );
  COND2X1 U2488 ( .A(n1887), .B(n2031), .C(n1490), .D(n1886), .Z(n562) );
  CANR2X1 U2489 ( .A(n1296), .B(n1929), .C(n1295), .D(n1965), .Z(n1894) );
  CANR2X1 U2490 ( .A(n1351), .B(n2406), .C(n1336), .D(n2405), .Z(n1891) );
  CIVX2 U2491 ( .A(out0_2[47]), .Z(n1889) );
  CANR2X1 U2492 ( .A(n1350), .B(n2441), .C(n1335), .D(n2410), .Z(n1890) );
  CND2X1 U2493 ( .A(n1891), .B(n1890), .Z(n2001) );
  CANR2X1 U2494 ( .A(n2218), .B(n1892), .C(n2207), .D(n2001), .Z(n1893) );
  CIVX2 U2495 ( .A(n1895), .Z(n2427) );
  CMXI2X1 U2496 ( .A0(n1265), .A1(n2427), .S(n1485), .Z(n2214) );
  COND2X1 U2497 ( .A(n2214), .B(n1361), .C(n1490), .D(n1896), .Z(n563) );
  CANR2X1 U2498 ( .A(n1296), .B(n1938), .C(n1295), .D(n1974), .Z(n1903) );
  CANR2X1 U2499 ( .A(n1335), .B(n2406), .C(n1351), .D(n2405), .Z(n1900) );
  CIVX2 U2500 ( .A(out0_2[46]), .Z(n1898) );
  CANR2X1 U2501 ( .A(n1336), .B(n2441), .C(n1352), .D(n2410), .Z(n1899) );
  CND2X1 U2502 ( .A(n1900), .B(n1899), .Z(n2010) );
  CANR2X1 U2503 ( .A(n2218), .B(n1901), .C(n2207), .D(n2010), .Z(n1902) );
  CND2X1 U2504 ( .A(n1903), .B(n1902), .Z(n2044) );
  COND2X1 U2505 ( .A(n1487), .B(n2044), .C(n1922), .D(n2043), .Z(n2228) );
  CIVX2 U2506 ( .A(n2228), .Z(n1905) );
  COND2X1 U2507 ( .A(n1905), .B(n1361), .C(n1490), .D(n1904), .Z(n564) );
  CANR2X1 U2508 ( .A(n1296), .B(n1947), .C(n1295), .D(n1983), .Z(n1912) );
  CANR2X1 U2509 ( .A(n1352), .B(n2406), .C(n1335), .D(n2405), .Z(n1909) );
  CIVX2 U2510 ( .A(out0_2[45]), .Z(n1907) );
  CANR2X1 U2511 ( .A(n1351), .B(n2441), .C(n1347), .D(n2410), .Z(n1908) );
  CND2X1 U2512 ( .A(n1909), .B(n1908), .Z(n2019) );
  CANR2X1 U2513 ( .A(n2218), .B(n1910), .C(n2207), .D(n2019), .Z(n1911) );
  CND2X1 U2514 ( .A(n1912), .B(n1911), .Z(n2057) );
  COND2X1 U2515 ( .A(n1486), .B(n2057), .C(n1922), .D(n2056), .Z(n2240) );
  CIVX2 U2516 ( .A(n2240), .Z(n1914) );
  COND2X1 U2517 ( .A(n1914), .B(n1361), .C(n1490), .D(n1913), .Z(n565) );
  CANR2X1 U2518 ( .A(n1296), .B(n1956), .C(n1295), .D(n1992), .Z(n1921) );
  CANR2X1 U2519 ( .A(n1347), .B(n2406), .C(n1352), .D(n2405), .Z(n1918) );
  CIVX2 U2520 ( .A(out0_2[44]), .Z(n1916) );
  CANR2X1 U2521 ( .A(n1335), .B(n2441), .C(n1341), .D(n2410), .Z(n1917) );
  CND2X1 U2522 ( .A(n1918), .B(n1917), .Z(n2028) );
  CANR2X1 U2523 ( .A(n2218), .B(n1919), .C(n2207), .D(n2028), .Z(n1920) );
  CND2X1 U2524 ( .A(n1921), .B(n1920), .Z(n2070) );
  COND2X1 U2525 ( .A(n1486), .B(n2070), .C(n1922), .D(n2069), .Z(n2252) );
  CIVX2 U2526 ( .A(n2252), .Z(n1924) );
  COND2X1 U2527 ( .A(n1924), .B(n1361), .C(n795), .D(n1923), .Z(n566) );
  CANR2X1 U2528 ( .A(n1296), .B(n1965), .C(n1295), .D(n2001), .Z(n1931) );
  CANR2X1 U2529 ( .A(n1341), .B(n2406), .C(n1347), .D(n2405), .Z(n1928) );
  CIVX2 U2530 ( .A(out0_2[43]), .Z(n1926) );
  CANR2X1 U2531 ( .A(n1352), .B(n2441), .C(n1342), .D(n2410), .Z(n1927) );
  CND2X1 U2532 ( .A(n1928), .B(n1927), .Z(n2038) );
  CIVX2 U2533 ( .A(n1932), .Z(n2082) );
  CMXI2X1 U2534 ( .A0(n1281), .A1(n2082), .S(n1486), .Z(n2255) );
  COND2X1 U2535 ( .A(n2255), .B(n1361), .C(n795), .D(n1933), .Z(n567) );
  CANR2X1 U2536 ( .A(n1296), .B(n1974), .C(n1295), .D(n2010), .Z(n1940) );
  CANR2X1 U2537 ( .A(n1342), .B(n2406), .C(n1341), .D(n2405), .Z(n1937) );
  CIVX2 U2538 ( .A(out0_2[42]), .Z(n1935) );
  CANR2X1 U2539 ( .A(n1347), .B(n2441), .C(n2410), .D(n1353), .Z(n1936) );
  CND2X1 U2540 ( .A(n1937), .B(n1936), .Z(n2051) );
  CIVX2 U2541 ( .A(n1941), .Z(n2092) );
  CMXI2X1 U2542 ( .A0(n1285), .A1(n2092), .S(n1486), .Z(n2268) );
  COND2X1 U2543 ( .A(n2268), .B(n1361), .C(n795), .D(n1942), .Z(n568) );
  CANR2X1 U2544 ( .A(n1296), .B(n1983), .C(n1295), .D(n2019), .Z(n1949) );
  CANR2X1 U2545 ( .A(n1353), .B(n2406), .C(n1342), .D(n2405), .Z(n1946) );
  CIVX2 U2546 ( .A(out0_2[41]), .Z(n1944) );
  CANR2X1 U2547 ( .A(n1341), .B(n2441), .C(n2410), .D(n1356), .Z(n1945) );
  CND2X1 U2548 ( .A(n1946), .B(n1945), .Z(n2064) );
  CIVX2 U2549 ( .A(n1950), .Z(n2102) );
  CMXI2X1 U2550 ( .A0(n1290), .A1(n2102), .S(n1485), .Z(n2281) );
  COND2X1 U2551 ( .A(n2281), .B(n1361), .C(n795), .D(n1951), .Z(n569) );
  CANR2X1 U2552 ( .A(n1296), .B(n1992), .C(n1295), .D(n2028), .Z(n1958) );
  CANR2X1 U2553 ( .A(n1356), .B(n2406), .C(n1353), .D(n2405), .Z(n1955) );
  CIVX2 U2554 ( .A(out0_2[40]), .Z(n1953) );
  CANR2X1 U2555 ( .A(n1342), .B(n2441), .C(n2410), .D(n1354), .Z(n1954) );
  CND2X1 U2556 ( .A(n1955), .B(n1954), .Z(n2077) );
  CIVX2 U2557 ( .A(n1959), .Z(n2112) );
  CMXI2X1 U2558 ( .A0(n1284), .A1(n2112), .S(n1485), .Z(n2294) );
  COND2X1 U2559 ( .A(n2294), .B(n1361), .C(n795), .D(n1960), .Z(n570) );
  CANR2X1 U2560 ( .A(n2406), .B(n1354), .C(n2405), .D(n1356), .Z(n1964) );
  CIVX2 U2561 ( .A(out0_2[39]), .Z(n1962) );
  CANR2X1 U2562 ( .A(n2441), .B(n1353), .C(n2410), .D(n1355), .Z(n1963) );
  CND2X1 U2563 ( .A(n1964), .B(n1963), .Z(n2087) );
  CANR2X1 U2564 ( .A(n2218), .B(n1965), .C(n2207), .D(n2087), .Z(n1966) );
  CIVX2 U2565 ( .A(n1968), .Z(n2122) );
  CMXI2X1 U2566 ( .A0(n1282), .A1(n2122), .S(n1485), .Z(n2307) );
  COND2X1 U2567 ( .A(n2307), .B(n1361), .C(n795), .D(n1969), .Z(n571) );
  CANR2X1 U2568 ( .A(n1296), .B(n2010), .C(n1295), .D(n2051), .Z(n1976) );
  CANR2X1 U2569 ( .A(n1355), .B(n2406), .C(n2405), .D(n1354), .Z(n1973) );
  CIVX2 U2570 ( .A(out0_2[38]), .Z(n1971) );
  CANR2X1 U2571 ( .A(n2441), .B(n1356), .C(n1339), .D(n2410), .Z(n1972) );
  CND2X1 U2572 ( .A(n1973), .B(n1972), .Z(n2097) );
  CIVX2 U2573 ( .A(n1977), .Z(n2132) );
  CMXI2X1 U2574 ( .A0(n1291), .A1(n2132), .S(n1485), .Z(n2320) );
  COND2X1 U2575 ( .A(n2320), .B(n1361), .C(n795), .D(n1978), .Z(n572) );
  CANR2X1 U2576 ( .A(n1296), .B(n2019), .C(n1295), .D(n2064), .Z(n1985) );
  CANR2X1 U2577 ( .A(n1339), .B(n2406), .C(n1355), .D(n2405), .Z(n1982) );
  CIVX2 U2578 ( .A(out0_2[37]), .Z(n1980) );
  CANR2X1 U2579 ( .A(n2441), .B(n1354), .C(n1340), .D(n2410), .Z(n1981) );
  CND2X1 U2580 ( .A(n1982), .B(n1981), .Z(n2107) );
  CIVX2 U2581 ( .A(n1986), .Z(n2142) );
  CMXI2X1 U2582 ( .A0(n1288), .A1(n2142), .S(n1485), .Z(n2333) );
  COND2X1 U2583 ( .A(n2333), .B(n1361), .C(n795), .D(n1987), .Z(n573) );
  CANR2X1 U2584 ( .A(n1296), .B(n2028), .C(n1295), .D(n2077), .Z(n1994) );
  CANR2X1 U2585 ( .A(n1340), .B(n2406), .C(n1339), .D(n2405), .Z(n1991) );
  CIVX2 U2586 ( .A(out0_2[36]), .Z(n1989) );
  CANR2X1 U2587 ( .A(n1355), .B(n2441), .C(n1334), .D(n2410), .Z(n1990) );
  CND2X1 U2588 ( .A(n1991), .B(n1990), .Z(n2117) );
  CIVX2 U2589 ( .A(n1995), .Z(n2152) );
  CMXI2X1 U2590 ( .A0(n1292), .A1(n2152), .S(n1485), .Z(n2346) );
  COND2X1 U2591 ( .A(n2346), .B(n1361), .C(n795), .D(n1996), .Z(n574) );
  CANR2X1 U2592 ( .A(n1296), .B(n2038), .C(n1295), .D(n2087), .Z(n2003) );
  CANR2X1 U2593 ( .A(n1334), .B(n2406), .C(n1340), .D(n2405), .Z(n2000) );
  CIVX2 U2594 ( .A(out0_2[35]), .Z(n1998) );
  CANR2X1 U2595 ( .A(n1339), .B(n2441), .C(n1333), .D(n2410), .Z(n1999) );
  CND2X1 U2596 ( .A(n2000), .B(n1999), .Z(n2127) );
  CIVX2 U2597 ( .A(n2004), .Z(n2162) );
  CMXI2X1 U2598 ( .A0(n1287), .A1(n2162), .S(n1485), .Z(n2359) );
  COND2X1 U2599 ( .A(n2359), .B(n1361), .C(n795), .D(n2005), .Z(n575) );
  CANR2X1 U2600 ( .A(n1296), .B(n2051), .C(n1295), .D(n2097), .Z(n2012) );
  CANR2X1 U2601 ( .A(n1333), .B(n2406), .C(n1334), .D(n2405), .Z(n2009) );
  CIVX2 U2602 ( .A(out0_2[34]), .Z(n2007) );
  CANR2X1 U2603 ( .A(n1340), .B(n2441), .C(n1331), .D(n2410), .Z(n2008) );
  CND2X1 U2604 ( .A(n2009), .B(n2008), .Z(n2137) );
  CIVX2 U2605 ( .A(n2013), .Z(n2172) );
  CMXI2X1 U2606 ( .A0(n1286), .A1(n2172), .S(n1485), .Z(n2376) );
  COND2X1 U2607 ( .A(n2376), .B(n1361), .C(n795), .D(n2014), .Z(n576) );
  CANR2X1 U2608 ( .A(n1296), .B(n2064), .C(n1295), .D(n2107), .Z(n2021) );
  CANR2X1 U2609 ( .A(n1331), .B(n2406), .C(n1333), .D(n2405), .Z(n2018) );
  CIVX2 U2610 ( .A(out0_2[33]), .Z(n2016) );
  CANR2X1 U2611 ( .A(n1334), .B(n2441), .C(n1332), .D(n2410), .Z(n2017) );
  CND2X1 U2612 ( .A(n2018), .B(n2017), .Z(n2147) );
  CIVX2 U2613 ( .A(n2022), .Z(n2182) );
  CMXI2X1 U2614 ( .A0(n1289), .A1(n2182), .S(n1485), .Z(n2390) );
  COND2X1 U2615 ( .A(n2390), .B(n1361), .C(n795), .D(n2023), .Z(n577) );
  CANR2X1 U2616 ( .A(n1296), .B(n2077), .C(n1295), .D(n2117), .Z(n2030) );
  CANR2X1 U2617 ( .A(n1332), .B(n2406), .C(n1331), .D(n2405), .Z(n2027) );
  CIVX2 U2618 ( .A(out0_2[32]), .Z(n2025) );
  CANR2X1 U2619 ( .A(n1333), .B(n2441), .C(n1330), .D(n2410), .Z(n2026) );
  CND2X1 U2620 ( .A(n2027), .B(n2026), .Z(n2157) );
  CIVX2 U2621 ( .A(n2031), .Z(n2193) );
  CMXI2X1 U2622 ( .A0(n1283), .A1(n2193), .S(n1485), .Z(n2404) );
  COND2X1 U2623 ( .A(n2404), .B(n1361), .C(n795), .D(n2032), .Z(n578) );
  CND2X1 U2624 ( .A(n1300), .B(n1488), .Z(n2448) );
  CANR2X1 U2625 ( .A(n2427), .B(n2192), .C(n1256), .D(n1265), .Z(n2042) );
  CANR2X1 U2626 ( .A(n1296), .B(n2087), .C(n1295), .D(n2127), .Z(n2040) );
  CANR2X1 U2627 ( .A(n1330), .B(n2406), .C(n1332), .D(n2405), .Z(n2037) );
  CIVX2 U2628 ( .A(out0_2[31]), .Z(n2035) );
  CANR2X1 U2629 ( .A(n1331), .B(n2441), .C(n1329), .D(n2410), .Z(n2036) );
  CND2X1 U2630 ( .A(n2037), .B(n2036), .Z(n2167) );
  CANR2X1 U2631 ( .A(n2218), .B(n2038), .C(n2207), .D(n2167), .Z(n2039) );
  CND2X1 U2632 ( .A(n2040), .B(n2039), .Z(n2449) );
  CIVX2 U2633 ( .A(n2449), .Z(n2213) );
  CANR2X1 U2634 ( .A(n2212), .B(n2213), .C(out2_2[31]), .D(n794), .Z(n2041) );
  CND2X1 U2635 ( .A(n2042), .B(n2041), .Z(n579) );
  CIVX2 U2636 ( .A(n2043), .Z(n2046) );
  CIVX2 U2637 ( .A(n2044), .Z(n2045) );
  CANR2X1 U2638 ( .A(n1255), .B(n2046), .C(n1256), .D(n2045), .Z(n2055) );
  CANR2X1 U2639 ( .A(n1296), .B(n2097), .C(n1295), .D(n2137), .Z(n2053) );
  CANR2X1 U2640 ( .A(n1329), .B(n2406), .C(n1330), .D(n2405), .Z(n2050) );
  CIVX2 U2641 ( .A(out0_2[30]), .Z(n2048) );
  CANR2X1 U2642 ( .A(n1332), .B(n2441), .C(n1314), .D(n2410), .Z(n2049) );
  CND2X1 U2643 ( .A(n2050), .B(n2049), .Z(n2177) );
  CANR2X1 U2644 ( .A(n2218), .B(n2051), .C(n2207), .D(n2177), .Z(n2052) );
  CANR2X1 U2645 ( .A(n2212), .B(n1277), .C(out2_2[30]), .D(n794), .Z(n2054) );
  CND2X1 U2646 ( .A(n2055), .B(n2054), .Z(n580) );
  CIVX2 U2647 ( .A(n2056), .Z(n2059) );
  CIVX2 U2648 ( .A(n2057), .Z(n2058) );
  CANR2X1 U2649 ( .A(n1255), .B(n2059), .C(n1256), .D(n2058), .Z(n2068) );
  CANR2X1 U2650 ( .A(n1296), .B(n2107), .C(n1295), .D(n2147), .Z(n2066) );
  CANR2X1 U2651 ( .A(n1314), .B(n2406), .C(n1329), .D(n2405), .Z(n2063) );
  CIVX2 U2652 ( .A(out0_2[29]), .Z(n2061) );
  CANR2X1 U2653 ( .A(n1330), .B(n2441), .C(n1310), .D(n2410), .Z(n2062) );
  CND2X1 U2654 ( .A(n2063), .B(n2062), .Z(n2187) );
  CANR2X1 U2655 ( .A(n2218), .B(n2064), .C(n2207), .D(n2187), .Z(n2065) );
  CANR2X1 U2656 ( .A(n2212), .B(n1278), .C(out2_2[29]), .D(n1169), .Z(n2067)
         );
  CND2X1 U2657 ( .A(n2068), .B(n2067), .Z(n581) );
  CIVX2 U2658 ( .A(n2069), .Z(n2072) );
  CIVX2 U2659 ( .A(n2070), .Z(n2071) );
  CANR2X1 U2660 ( .A(n1255), .B(n2072), .C(n1256), .D(n2071), .Z(n2081) );
  CANR2X1 U2661 ( .A(n1296), .B(n2117), .C(n1295), .D(n2157), .Z(n2079) );
  CANR2X1 U2662 ( .A(n1310), .B(n2406), .C(n1314), .D(n2405), .Z(n2076) );
  CIVX2 U2663 ( .A(out0_2[28]), .Z(n2074) );
  CANR2X1 U2664 ( .A(n1329), .B(n2441), .C(n1313), .D(n2410), .Z(n2075) );
  CND2X1 U2665 ( .A(n2076), .B(n2075), .Z(n2198) );
  CANR2X1 U2666 ( .A(n2218), .B(n2077), .C(n2207), .D(n2198), .Z(n2078) );
  CANR2X1 U2667 ( .A(n2212), .B(n1279), .C(out2_2[28]), .D(n1169), .Z(n2080)
         );
  CND2X1 U2668 ( .A(n2081), .B(n2080), .Z(n582) );
  CANR2X1 U2669 ( .A(n2082), .B(n2192), .C(n1281), .D(n1256), .Z(n2091) );
  CANR2X1 U2670 ( .A(n1296), .B(n2127), .C(n1295), .D(n2167), .Z(n2089) );
  CANR2X1 U2671 ( .A(n1313), .B(n2406), .C(n1310), .D(n2405), .Z(n2086) );
  CIVX2 U2672 ( .A(out0_2[27]), .Z(n2084) );
  CANR2X1 U2673 ( .A(n1314), .B(n2441), .C(n1307), .D(n2410), .Z(n2085) );
  CND2X1 U2674 ( .A(n2086), .B(n2085), .Z(n2208) );
  CANR2X1 U2675 ( .A(n2218), .B(n2087), .C(n2207), .D(n2208), .Z(n2088) );
  CANR2X1 U2676 ( .A(n2212), .B(n1266), .C(out2_2[27]), .D(n1169), .Z(n2090)
         );
  CND2X1 U2677 ( .A(n2091), .B(n2090), .Z(n583) );
  CANR2X1 U2678 ( .A(n2092), .B(n2192), .C(n1285), .D(n1256), .Z(n2101) );
  CANR2X1 U2679 ( .A(n1296), .B(n2137), .C(n1295), .D(n2177), .Z(n2099) );
  CANR2X1 U2680 ( .A(n1307), .B(n2406), .C(n1313), .D(n2405), .Z(n2096) );
  CIVX2 U2681 ( .A(out0_2[26]), .Z(n2094) );
  CANR2X1 U2682 ( .A(n1310), .B(n2441), .C(n1315), .D(n2410), .Z(n2095) );
  CND2X1 U2683 ( .A(n2096), .B(n2095), .Z(n2226) );
  CANR2X1 U2684 ( .A(n2218), .B(n2097), .C(n2207), .D(n2226), .Z(n2098) );
  CANR2X1 U2685 ( .A(n2212), .B(n1272), .C(out2_2[26]), .D(n1494), .Z(n2100)
         );
  CND2X1 U2686 ( .A(n2101), .B(n2100), .Z(n584) );
  CANR2X1 U2687 ( .A(n2102), .B(n2192), .C(n1290), .D(n1256), .Z(n2111) );
  CANR2X1 U2688 ( .A(n1296), .B(n2147), .C(n1295), .D(n2187), .Z(n2109) );
  CANR2X1 U2689 ( .A(n1315), .B(n2406), .C(n1307), .D(n2405), .Z(n2106) );
  CIVX2 U2690 ( .A(out0_2[25]), .Z(n2104) );
  CANR2X1 U2691 ( .A(n1313), .B(n2441), .C(n1328), .D(n2410), .Z(n2105) );
  CND2X1 U2692 ( .A(n2106), .B(n2105), .Z(n2238) );
  CANR2X1 U2693 ( .A(n2218), .B(n2107), .C(n2207), .D(n2238), .Z(n2108) );
  CANR2X1 U2694 ( .A(n2212), .B(n1280), .C(out2_2[25]), .D(n1494), .Z(n2110)
         );
  CND2X1 U2695 ( .A(n2111), .B(n2110), .Z(n585) );
  CANR2X1 U2696 ( .A(n2112), .B(n2192), .C(n1284), .D(n1256), .Z(n2121) );
  CANR2X1 U2697 ( .A(n1296), .B(n2157), .C(n1295), .D(n2198), .Z(n2119) );
  CANR2X1 U2698 ( .A(n1328), .B(n2406), .C(n1315), .D(n2405), .Z(n2116) );
  CIVX2 U2699 ( .A(out0_2[24]), .Z(n2114) );
  CANR2X1 U2700 ( .A(n1307), .B(n2441), .C(n1327), .D(n2410), .Z(n2115) );
  CND2X1 U2701 ( .A(n2116), .B(n2115), .Z(n2250) );
  CANR2X1 U2702 ( .A(n2218), .B(n2117), .C(n2207), .D(n2250), .Z(n2118) );
  CANR2X1 U2703 ( .A(n2212), .B(n1271), .C(out2_2[24]), .D(n1494), .Z(n2120)
         );
  CND2X1 U2704 ( .A(n2121), .B(n2120), .Z(n586) );
  CANR2X1 U2705 ( .A(n2122), .B(n2192), .C(n1282), .D(n1256), .Z(n2131) );
  CANR2X1 U2706 ( .A(n1296), .B(n2167), .C(n1295), .D(n2208), .Z(n2129) );
  CANR2X1 U2707 ( .A(n1327), .B(n2406), .C(n1328), .D(n2405), .Z(n2126) );
  CIVX2 U2708 ( .A(out0_2[23]), .Z(n2124) );
  CANR2X1 U2709 ( .A(n1315), .B(n2441), .C(n1312), .D(n2410), .Z(n2125) );
  CND2X1 U2710 ( .A(n2126), .B(n2125), .Z(n2263) );
  CANR2X1 U2711 ( .A(n2218), .B(n2127), .C(n2207), .D(n2263), .Z(n2128) );
  CANR2X1 U2712 ( .A(n2212), .B(n1270), .C(out2_2[23]), .D(n1493), .Z(n2130)
         );
  CND2X1 U2713 ( .A(n2131), .B(n2130), .Z(n587) );
  CANR2X1 U2714 ( .A(n2132), .B(n2192), .C(n1291), .D(n1256), .Z(n2141) );
  CANR2X1 U2715 ( .A(n1296), .B(n2177), .C(n1295), .D(n2226), .Z(n2139) );
  CANR2X1 U2716 ( .A(n1312), .B(n2406), .C(n1327), .D(n2405), .Z(n2136) );
  CIVX2 U2717 ( .A(out0_2[22]), .Z(n2134) );
  CANR2X1 U2718 ( .A(n1328), .B(n2441), .C(n1306), .D(n2410), .Z(n2135) );
  CND2X1 U2719 ( .A(n2136), .B(n2135), .Z(n2276) );
  CANR2X1 U2720 ( .A(n2218), .B(n2137), .C(n2207), .D(n2276), .Z(n2138) );
  CANR2X1 U2721 ( .A(n2212), .B(n1273), .C(out2_2[22]), .D(n1493), .Z(n2140)
         );
  CND2X1 U2722 ( .A(n2141), .B(n2140), .Z(n588) );
  CANR2X1 U2723 ( .A(n2142), .B(n2192), .C(n1288), .D(n1256), .Z(n2151) );
  CANR2X1 U2724 ( .A(n1296), .B(n2187), .C(n1295), .D(n2238), .Z(n2149) );
  CANR2X1 U2725 ( .A(n1306), .B(n2406), .C(n1312), .D(n2405), .Z(n2146) );
  CIVX2 U2726 ( .A(out0_2[21]), .Z(n2144) );
  CANR2X1 U2727 ( .A(n1327), .B(n2441), .C(n1304), .D(n2410), .Z(n2145) );
  CND2X1 U2728 ( .A(n2146), .B(n2145), .Z(n2289) );
  CANR2X1 U2729 ( .A(n2218), .B(n2147), .C(n2207), .D(n2289), .Z(n2148) );
  CANR2X1 U2730 ( .A(n2212), .B(n1274), .C(out2_2[21]), .D(n1493), .Z(n2150)
         );
  CND2X1 U2731 ( .A(n2151), .B(n2150), .Z(n589) );
  CANR2X1 U2732 ( .A(n2152), .B(n2192), .C(n1292), .D(n1256), .Z(n2161) );
  CANR2X1 U2733 ( .A(n1296), .B(n2198), .C(n1295), .D(n2250), .Z(n2159) );
  CANR2X1 U2734 ( .A(n1304), .B(n2406), .C(n1306), .D(n2405), .Z(n2156) );
  CIVX2 U2735 ( .A(out0_2[20]), .Z(n2154) );
  CANR2X1 U2736 ( .A(n1312), .B(n2441), .C(n1309), .D(n2410), .Z(n2155) );
  CND2X1 U2737 ( .A(n2156), .B(n2155), .Z(n2302) );
  CANR2X1 U2738 ( .A(n2218), .B(n2157), .C(n2207), .D(n2302), .Z(n2158) );
  CANR2X1 U2739 ( .A(n2212), .B(n1275), .C(out2_2[20]), .D(n1492), .Z(n2160)
         );
  CND2X1 U2740 ( .A(n2161), .B(n2160), .Z(n590) );
  CANR2X1 U2741 ( .A(n2162), .B(n2192), .C(n1287), .D(n1256), .Z(n2171) );
  CANR2X1 U2742 ( .A(n1296), .B(n2208), .C(n1295), .D(n2263), .Z(n2169) );
  CANR2X1 U2743 ( .A(n1309), .B(n2406), .C(n1304), .D(n2405), .Z(n2166) );
  CIVX2 U2744 ( .A(out0_2[19]), .Z(n2164) );
  CANR2X1 U2745 ( .A(n1306), .B(n2441), .C(n1302), .D(n2410), .Z(n2165) );
  CND2X1 U2746 ( .A(n2166), .B(n2165), .Z(n2315) );
  CANR2X1 U2747 ( .A(n2212), .B(n1268), .C(out2_2[19]), .D(n1492), .Z(n2170)
         );
  CND2X1 U2748 ( .A(n2171), .B(n2170), .Z(n591) );
  CANR2X1 U2749 ( .A(n2172), .B(n2192), .C(n1286), .D(n1256), .Z(n2181) );
  CANR2X1 U2750 ( .A(n1296), .B(n2226), .C(n1295), .D(n2276), .Z(n2179) );
  CANR2X1 U2751 ( .A(n1302), .B(n2406), .C(n1309), .D(n2405), .Z(n2176) );
  CIVX2 U2752 ( .A(out0_2[18]), .Z(n2174) );
  CANR2X1 U2753 ( .A(n1304), .B(n2441), .C(n1308), .D(n2410), .Z(n2175) );
  CND2X1 U2754 ( .A(n2176), .B(n2175), .Z(n2328) );
  CANR2X1 U2755 ( .A(n2218), .B(n2177), .C(n2207), .D(n2328), .Z(n2178) );
  CANR2X1 U2756 ( .A(n2212), .B(n1269), .C(out2_2[18]), .D(n1492), .Z(n2180)
         );
  CND2X1 U2757 ( .A(n2181), .B(n2180), .Z(n592) );
  CANR2X1 U2758 ( .A(n2182), .B(n2192), .C(n1289), .D(n1256), .Z(n2191) );
  CANR2X1 U2759 ( .A(n1296), .B(n2238), .C(n1295), .D(n2289), .Z(n2189) );
  CANR2X1 U2760 ( .A(n1308), .B(n2406), .C(n1302), .D(n2405), .Z(n2186) );
  CIVX2 U2761 ( .A(out0_2[17]), .Z(n2184) );
  CANR2X1 U2762 ( .A(n1309), .B(n2441), .C(n1305), .D(n2410), .Z(n2185) );
  CND2X1 U2763 ( .A(n2186), .B(n2185), .Z(n2341) );
  CANR2X1 U2764 ( .A(n2218), .B(n2187), .C(n2207), .D(n2341), .Z(n2188) );
  CANR2X1 U2765 ( .A(n2212), .B(n1276), .C(out2_2[17]), .D(n1491), .Z(n2190)
         );
  CND2X1 U2766 ( .A(n2191), .B(n2190), .Z(n593) );
  CANR2X1 U2767 ( .A(n2193), .B(n2192), .C(n1283), .D(n1256), .Z(n2202) );
  CANR2X1 U2768 ( .A(n1296), .B(n2250), .C(n1295), .D(n2302), .Z(n2200) );
  CANR2X1 U2769 ( .A(n1305), .B(n2406), .C(n1308), .D(n2405), .Z(n2197) );
  CIVX2 U2770 ( .A(out0_2[16]), .Z(n2195) );
  CANR2X1 U2771 ( .A(n1302), .B(n2441), .C(n1311), .D(n2410), .Z(n2196) );
  CND2X1 U2772 ( .A(n2197), .B(n2196), .Z(n2354) );
  CANR2X1 U2773 ( .A(n2218), .B(n2198), .C(n2207), .D(n2354), .Z(n2199) );
  CANR2X1 U2774 ( .A(n2212), .B(n1267), .C(out2_2[16]), .D(n1491), .Z(n2201)
         );
  CND2X1 U2775 ( .A(n2202), .B(n2201), .Z(n594) );
  CANR2X1 U2776 ( .A(n1296), .B(n2263), .C(n1295), .D(n2315), .Z(n2210) );
  CANR2X1 U2777 ( .A(n1311), .B(n2406), .C(n1305), .D(n2405), .Z(n2206) );
  CIVX2 U2778 ( .A(out0_2[15]), .Z(n2204) );
  CANR2X1 U2779 ( .A(n1308), .B(n2441), .C(n1303), .D(n2410), .Z(n2205) );
  CND2X1 U2780 ( .A(n2206), .B(n2205), .Z(n2371) );
  CANR2X1 U2781 ( .A(n2218), .B(n2208), .C(n2207), .D(n2371), .Z(n2209) );
  CND2X1 U2782 ( .A(n2210), .B(n2209), .Z(n2432) );
  CIVX2 U2783 ( .A(n2432), .Z(n2211) );
  CANR2X1 U2784 ( .A(n1256), .B(n2213), .C(n2212), .D(n2211), .Z(n2217) );
  CIVX2 U2785 ( .A(n2214), .Z(n2215) );
  CANR2X1 U2786 ( .A(n1300), .B(n2215), .C(out2_2[15]), .D(n1491), .Z(n2216)
         );
  CND2X1 U2787 ( .A(n2217), .B(n2216), .Z(n595) );
  CIVX2 U2788 ( .A(n2276), .Z(n2219) );
  CIVX2 U2789 ( .A(n2328), .Z(n2269) );
  CANR2X1 U2790 ( .A(n2219), .B(n2414), .C(n2269), .D(n2447), .Z(n2225) );
  CANR2X1 U2791 ( .A(n1303), .B(n2406), .C(n1311), .D(n2405), .Z(n2223) );
  CIVX2 U2792 ( .A(out0_2[14]), .Z(n2221) );
  CANR2X1 U2793 ( .A(n1259), .B(n1258), .C(n1277), .D(n1486), .Z(n2224) );
  COND3X1 U2794 ( .A(n2430), .B(n2226), .C(n2225), .D(n2224), .Z(n2227) );
  CANR2X1 U2795 ( .A(n1300), .B(n2228), .C(n2422), .D(n2227), .Z(n2229) );
  CIVX2 U2796 ( .A(n2289), .Z(n2231) );
  CIVX2 U2797 ( .A(n2341), .Z(n2282) );
  CANR2X1 U2798 ( .A(n2231), .B(n2414), .C(n2282), .D(n2447), .Z(n2237) );
  CANR2X1 U2799 ( .A(n1318), .B(n2406), .C(n1303), .D(n2405), .Z(n2235) );
  CIVX2 U2800 ( .A(out0_2[13]), .Z(n2233) );
  CANR2X1 U2801 ( .A(n1260), .B(n1258), .C(n1278), .D(n1486), .Z(n2236) );
  COND3X1 U2802 ( .A(n2430), .B(n2238), .C(n2237), .D(n2236), .Z(n2239) );
  CANR2X1 U2803 ( .A(n1300), .B(n2240), .C(n2422), .D(n2239), .Z(n2241) );
  CIVX2 U2804 ( .A(n2302), .Z(n2243) );
  CIVX2 U2805 ( .A(n2354), .Z(n2295) );
  CANR2X1 U2806 ( .A(n2243), .B(n2414), .C(n2295), .D(n2447), .Z(n2249) );
  CANR2X1 U2807 ( .A(n1319), .B(n2406), .C(n1318), .D(n2405), .Z(n2247) );
  CIVX2 U2808 ( .A(out0_2[12]), .Z(n2245) );
  CANR2X1 U2809 ( .A(n1261), .B(n1258), .C(n1279), .D(n1486), .Z(n2248) );
  COND3X1 U2810 ( .A(n2430), .B(n2250), .C(n2249), .D(n2248), .Z(n2251) );
  CANR2X1 U2811 ( .A(n1300), .B(n2252), .C(n2422), .D(n2251), .Z(n2253) );
  CIVX2 U2812 ( .A(n2315), .Z(n2256) );
  CIVX2 U2813 ( .A(n2371), .Z(n2308) );
  CANR2X1 U2814 ( .A(n2256), .B(n2414), .C(n2308), .D(n2447), .Z(n2262) );
  CANR2X1 U2815 ( .A(n1320), .B(n2406), .C(n1319), .D(n2405), .Z(n2260) );
  CIVX2 U2816 ( .A(out0_2[11]), .Z(n2258) );
  CANR2X1 U2817 ( .A(n1318), .B(n2441), .C(n1317), .D(n2410), .Z(n2259) );
  CND2X1 U2818 ( .A(n2260), .B(n2259), .Z(n2431) );
  CIVX2 U2819 ( .A(n2431), .Z(n2361) );
  CANR2X1 U2820 ( .A(n2361), .B(n1258), .C(n1266), .D(n1486), .Z(n2261) );
  COND3X1 U2821 ( .A(n2430), .B(n2263), .C(n2262), .D(n2261), .Z(n2264) );
  CANR2X1 U2822 ( .A(n1300), .B(n2265), .C(n2422), .D(n2264), .Z(n2266) );
  CANR2X1 U2823 ( .A(n2269), .B(n2414), .C(n1259), .D(n2447), .Z(n2275) );
  CANR2X1 U2824 ( .A(n1317), .B(n2406), .C(n1320), .D(n2405), .Z(n2273) );
  CIVX2 U2825 ( .A(out0_2[10]), .Z(n2271) );
  CANR2X1 U2826 ( .A(n1262), .B(n1258), .C(n1272), .D(n1486), .Z(n2274) );
  COND3X1 U2827 ( .A(n2430), .B(n2276), .C(n2275), .D(n2274), .Z(n2277) );
  CANR2X1 U2828 ( .A(n1300), .B(n2278), .C(n2422), .D(n2277), .Z(n2279) );
  CIVX2 U2829 ( .A(n2281), .Z(n2291) );
  CANR2X1 U2830 ( .A(n2282), .B(n2414), .C(n1260), .D(n2447), .Z(n2288) );
  CANR2X1 U2831 ( .A(n1322), .B(n2406), .C(n1317), .D(n2405), .Z(n2286) );
  CIVX2 U2832 ( .A(out0_2[9]), .Z(n2284) );
  CANR2X1 U2833 ( .A(n1263), .B(n1258), .C(n1280), .D(n1486), .Z(n2287) );
  CANR2X1 U2834 ( .A(n1300), .B(n2291), .C(n2422), .D(n2290), .Z(n2292) );
  CANR2X1 U2835 ( .A(n2295), .B(n2414), .C(n1261), .D(n2447), .Z(n2301) );
  CANR2X1 U2836 ( .A(n1323), .B(n2406), .C(n1322), .D(n2405), .Z(n2299) );
  CIVX2 U2837 ( .A(out0_2[8]), .Z(n2297) );
  CANR2X1 U2838 ( .A(n1264), .B(n1258), .C(n1271), .D(n1486), .Z(n2300) );
  COND3X1 U2839 ( .A(n2430), .B(n2302), .C(n2301), .D(n2300), .Z(n2303) );
  CANR2X1 U2840 ( .A(n1300), .B(n2304), .C(n2422), .D(n2303), .Z(n2305) );
  CIVX2 U2841 ( .A(n2307), .Z(n2317) );
  CANR2X1 U2842 ( .A(n2308), .B(n2414), .C(n2361), .D(n2447), .Z(n2314) );
  CANR2X1 U2843 ( .A(n1324), .B(n2406), .C(n1323), .D(n2405), .Z(n2312) );
  CIVX2 U2844 ( .A(out0_2[7]), .Z(n2310) );
  CANR2X1 U2845 ( .A(n1322), .B(n2441), .C(n1321), .D(n2410), .Z(n2311) );
  CND2X1 U2846 ( .A(n2312), .B(n2311), .Z(n2444) );
  CIVX2 U2847 ( .A(n2444), .Z(n2360) );
  CANR2X1 U2848 ( .A(n2360), .B(n1258), .C(n1270), .D(n1486), .Z(n2313) );
  COND3X1 U2849 ( .A(n2430), .B(n2315), .C(n2314), .D(n2313), .Z(n2316) );
  CANR2X1 U2850 ( .A(n1300), .B(n2317), .C(n2422), .D(n2316), .Z(n2318) );
  CIVX2 U2851 ( .A(n2320), .Z(n2330) );
  CANR2X1 U2852 ( .A(n1259), .B(n2414), .C(n1262), .D(n2447), .Z(n2327) );
  CANR2X1 U2853 ( .A(n1321), .B(n2406), .C(n1324), .D(n2405), .Z(n2324) );
  CIVX2 U2854 ( .A(out0_2[6]), .Z(n2322) );
  CANR2X1 U2855 ( .A(n1323), .B(n2441), .C(n1325), .D(n2410), .Z(n2323) );
  CND2X1 U2856 ( .A(n2324), .B(n2323), .Z(n2385) );
  CIVX2 U2857 ( .A(n2385), .Z(n2325) );
  CANR2X1 U2858 ( .A(n2325), .B(n1258), .C(n1273), .D(n1486), .Z(n2326) );
  COND3X1 U2859 ( .A(n2430), .B(n2328), .C(n2327), .D(n2326), .Z(n2329) );
  CANR2X1 U2860 ( .A(n1300), .B(n2330), .C(n2422), .D(n2329), .Z(n2331) );
  CIVX2 U2861 ( .A(out2_2[5]), .Z(n2345) );
  CIVX2 U2862 ( .A(n2333), .Z(n2343) );
  CANR2X1 U2863 ( .A(n1260), .B(n2414), .C(n1263), .D(n2447), .Z(n2340) );
  CANR2X1 U2864 ( .A(n1325), .B(n2406), .C(n1321), .D(n2405), .Z(n2337) );
  CIVX2 U2865 ( .A(out0_2[5]), .Z(n2335) );
  CIVX2 U2866 ( .A(n2379), .Z(n2362) );
  CANR2X1 U2867 ( .A(n1324), .B(n2441), .C(n2362), .D(n2410), .Z(n2336) );
  CND2X1 U2868 ( .A(n2337), .B(n2336), .Z(n2399) );
  CIVX2 U2869 ( .A(n2399), .Z(n2338) );
  CANR2X1 U2870 ( .A(n2338), .B(n1258), .C(n1274), .D(n1486), .Z(n2339) );
  COND3X1 U2871 ( .A(n2430), .B(n2341), .C(n2340), .D(n2339), .Z(n2342) );
  CANR2X1 U2872 ( .A(n1300), .B(n2343), .C(n2422), .D(n2342), .Z(n2344) );
  CIVX2 U2873 ( .A(n2346), .Z(n2356) );
  CANR2X1 U2874 ( .A(n1261), .B(n2414), .C(n1264), .D(n2447), .Z(n2353) );
  CANR2X1 U2875 ( .A(n2362), .B(n2406), .C(n1325), .D(n2405), .Z(n2350) );
  CIVX2 U2876 ( .A(out0_2[4]), .Z(n2348) );
  CIVX2 U2877 ( .A(n2393), .Z(n2363) );
  CANR2X1 U2878 ( .A(n1321), .B(n2441), .C(n2363), .D(n2410), .Z(n2349) );
  CND2X1 U2879 ( .A(n2350), .B(n2349), .Z(n2419) );
  CIVX2 U2880 ( .A(n2419), .Z(n2351) );
  CANR2X1 U2881 ( .A(n2351), .B(n1258), .C(n1275), .D(n1486), .Z(n2352) );
  COND3X1 U2882 ( .A(n2430), .B(n2354), .C(n2353), .D(n2352), .Z(n2355) );
  CANR2X1 U2883 ( .A(n1300), .B(n2356), .C(n2422), .D(n2355), .Z(n2357) );
  CIVX2 U2884 ( .A(n2359), .Z(n2373) );
  CANR2X1 U2885 ( .A(n2361), .B(n2414), .C(n2447), .D(n2360), .Z(n2370) );
  CANR2X1 U2886 ( .A(n2363), .B(n2406), .C(n2362), .D(n2405), .Z(n2368) );
  CIVX2 U2887 ( .A(out0_2[3]), .Z(n2365) );
  CIVX2 U2888 ( .A(n2411), .Z(n2366) );
  CANR2X1 U2889 ( .A(n1325), .B(n2441), .C(n2366), .D(n2410), .Z(n2367) );
  CANR2X1 U2890 ( .A(n1294), .B(n1258), .C(n1268), .D(n1486), .Z(n2369) );
  COND3X1 U2891 ( .A(n2430), .B(n2371), .C(n2370), .D(n2369), .Z(n2372) );
  CANR2X1 U2892 ( .A(n1300), .B(n2373), .C(n2422), .D(n2372), .Z(n2374) );
  CANR2X1 U2893 ( .A(n2406), .B(n2411), .C(n2405), .D(n2393), .Z(n2381) );
  CIVX2 U2894 ( .A(out0_2[2]), .Z(n2378) );
  CANR2X1 U2895 ( .A(n2441), .B(n2379), .C(n2410), .D(n2440), .Z(n2380) );
  CND2X1 U2896 ( .A(n2381), .B(n2380), .Z(n2382) );
  CANR2X1 U2897 ( .A(n1258), .B(n2382), .C(n1262), .D(n2414), .Z(n2384) );
  CANR2X1 U2898 ( .A(n1259), .B(n2416), .C(n1269), .D(n1486), .Z(n2383) );
  COND3X1 U2899 ( .A(n2420), .B(n2385), .C(n2384), .D(n2383), .Z(n2386) );
  CANR2X1 U2900 ( .A(n1300), .B(n2387), .C(n2422), .D(n2386), .Z(n2388) );
  CIVX2 U2901 ( .A(n2390), .Z(n2401) );
  CANR2X1 U2902 ( .A(n2406), .B(n2440), .C(n2405), .D(n2411), .Z(n2395) );
  CANR2X1 U2903 ( .A(n2441), .B(n2393), .C(n2410), .D(n2433), .Z(n2394) );
  CND2X1 U2904 ( .A(n2395), .B(n2394), .Z(n2396) );
  CANR2X1 U2905 ( .A(n1258), .B(n2396), .C(n1263), .D(n2414), .Z(n2398) );
  CANR2X1 U2906 ( .A(n1260), .B(n2416), .C(n1276), .D(n1486), .Z(n2397) );
  COND3X1 U2907 ( .A(n2420), .B(n2399), .C(n2398), .D(n2397), .Z(n2400) );
  CANR2X1 U2908 ( .A(n1300), .B(n2401), .C(n2422), .D(n2400), .Z(n2402) );
  CANR2X1 U2909 ( .A(n2406), .B(n2433), .C(n2405), .D(n2440), .Z(n2413) );
  CIVX2 U2910 ( .A(out0_2[0]), .Z(n2409) );
  CANR2X1 U2911 ( .A(n2441), .B(n2411), .C(n2410), .D(n2434), .Z(n2412) );
  CND2X1 U2912 ( .A(n2413), .B(n2412), .Z(n2415) );
  CANR2X1 U2913 ( .A(n1258), .B(n2415), .C(n1264), .D(n2414), .Z(n2418) );
  CANR2X1 U2914 ( .A(n1261), .B(n2416), .C(n1267), .D(n1486), .Z(n2417) );
  COND3X1 U2915 ( .A(n2420), .B(n2419), .C(n2418), .D(n2417), .Z(n2421) );
  CANR2X1 U2916 ( .A(n1300), .B(n2423), .C(n2422), .D(n2421), .Z(n2424) );
  CND4X1 U2917 ( .A(h0_1[6]), .B(n1490), .C(n2427), .D(n2426), .Z(n2429) );
  CND2X1 U2918 ( .A(n1265), .B(n1300), .Z(n2428) );
  CMXI2X1 U2919 ( .A0(n2429), .A1(n2428), .S(n1485), .Z(n2453) );
  COND2X1 U2920 ( .A(n2432), .B(n1488), .C(n2431), .D(n2430), .Z(n2446) );
  CIVX2 U2921 ( .A(n2433), .Z(n2438) );
  CIVX2 U2922 ( .A(n2434), .Z(n2436) );
  COND2X1 U2923 ( .A(n2438), .B(n2437), .C(n2436), .D(n2435), .Z(n2439) );
  COND4CX1 U2924 ( .A(n2441), .B(n2440), .C(n2439), .D(n1258), .Z(n2442) );
  CANR3X1 U2925 ( .A(n2447), .B(n1294), .C(n2446), .D(n2445), .Z(n2451) );
  COND2X1 U2926 ( .A(n2451), .B(n1361), .C(n2449), .D(n2448), .Z(n2452) );
  COND4CX1 U2927 ( .A(n795), .B(n1484), .C(n2455), .D(n2454), .Z(n611) );
  CANR2X1 U2928 ( .A(out0_2[0]), .B(n1357), .C(N418), .D(n1298), .Z(n2457) );
  CANR2X1 U2929 ( .A(out1_2[0]), .B(n1299), .C(acc[0]), .D(n2461), .Z(n2456)
         );
  CND2X1 U2930 ( .A(n2457), .B(n2456), .Z(n544) );
  CIVX2 U2931 ( .A(n12), .Z(n2458) );
  CIVX2 U2932 ( .A(n1213), .Z(n2466) );
  CIVX2 U2933 ( .A(n1215), .Z(n2467) );
endmodule

