
module bits ( clk, rst, pushin, datain, reqin, reqlen, pushout, lenout, 
        dataout );
  input [31:0] datain;
  input [3:0] reqlen;
  output [3:0] lenout;
  output [14:0] dataout;
  input clk, rst, pushin, reqin;
  output pushout;
  wire   N111, N112, N113, N114, pushout_stg_1, N118, N119, N120, N121, N16590,
         N16591, N16592, N16593, N16594, N16595, N16596, N16597, N16598,
         N16599, n4, n5, n8, n9, n10, n11, n12, n13, n14, n16, n17, n19, n20,
         n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n38, n39, n40, n41, n44, n46, n48, n49, n50, n52, n54, n56, n57,
         n58, n60, n61, n62, n64, n65, n67, n68, n69, n70, n71, n72, n75, n76,
         n78, n79, n80, n84, n86, n89, n90, n92, n93, n94, n96, n97, n99, n100,
         n101, n102, n104, n105, n107, n108, n109, n111, n112, n113, n114,
         n115, n116, n117, n118, n120, n124, n125, n126, n127, n129, n130,
         n131, n132, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n172, n173, n174, n175, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n195, n197, n198, n199, n201, n202, n203, n204,
         n205, n206, n207, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n221, n222, n223, n224, n225, n226, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n243, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n262, n263, n264, n265,
         n266, n267, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n281, n282, n284, n285, n286, n287, n288, n289, n290,
         n291, n293, n294, n295, n296, n297, n298, n299, n300, n301, n303,
         n304, n306, n307, n308, n310, n311, n312, n313, n314, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n328, n329,
         n330, n331, n332, n333, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n348, n349, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n384, n385, n386, n387, n388, n390,
         n391, n392, n393, n394, n395, n396, n409, n410, n411, n412, n421,
         n422, n423, n424, n433, n434, n435, n436, n437, n438, n439, n440,
         n449, n450, n451, n452, n461, n462, n463, n464, n465, n466, n475,
         n476, n477, n478, n488, n490, n491, n492, n493, n495, n496, n497,
         n498, n499, n500, n509, n510, n511, n512, n513, n522, n523, n524,
         n525, n534, n535, n536, n537, n538, n539, n540, n541, n550, n551,
         n552, n553, n562, n563, n564, n565, n566, n567, n576, n577, n578,
         n579, n588, n589, n590, n591, n592, n593, n594, n596, n597, n598,
         n599, n600, n601, n610, n611, n612, n613, n622, n623, n624, n625,
         n634, n635, n636, n637, n638, n639, n640, n641, n650, n651, n652,
         n653, n662, n663, n664, n665, n666, n667, n676, n677, n678, n679,
         n688, n689, n690, n691, n692, n694, n695, n697, n699, n700, n701,
         n702, n703, n712, n713, n714, n715, n724, n725, n726, n727, n736,
         n737, n738, n739, n740, n741, n742, n743, n752, n753, n754, n755,
         n764, n765, n766, n767, n768, n769, n778, n779, n780, n781, n790,
         n791, n792, n793, n794, n795, n797, n798, n799, n800, n801, n802,
         n811, n812, n813, n814, n823, n824, n825, n826, n835, n836, n837,
         n838, n839, n840, n841, n842, n851, n852, n853, n854, n863, n864,
         n865, n866, n867, n868, n877, n878, n879, n880, n889, n890, n891,
         n892, n893, n894, n895, n897, n899, n900, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n920, n921, n926, n927, n928,
         n929, n938, n940, n941, n942, n945, n946, n947, n948, n949, n950,
         n959, n960, n961, n962, n971, n972, n973, n974, n975, n976, n985,
         n986, n987, n988, n997, n998, n999, n1000, n1001, n1002, n1003, n1005,
         n1006, n1007, n1008, n1009, n1010, n1019, n1020, n1021, n1022, n1031,
         n1032, n1033, n1034, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1059, n1060, n1061, n1062, n1071, n1072, n1073, n1074, n1075,
         n1076, n1085, n1086, n1087, n1088, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1113, n1114, n1115, n1116, n1125, n1126, n1127,
         n1128, n1129, n1130, n1139, n1140, n1141, n1142, n1152, n1153, n1154,
         n1156, n1157, n1158, n1159, n1160, n1161, n1170, n1171, n1172, n1173,
         n1174, n1183, n1184, n1185, n1186, n1195, n1196, n1198, n1200, n1202,
         n1204, n1205, n1206, n1207, n1208, n1210, n1211, n1212, n1213, n1214,
         n1215, n1224, n1225, n1226, n1227, n1236, n1237, n1238, n1239, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1264, n1265, n1266,
         n1267, n1276, n1277, n1278, n1279, n1280, n1281, n1290, n1291, n1292,
         n1293, n1302, n1303, n1304, n1305, n1306, n1307, n1309, n1310, n1311,
         n1312, n1313, n1314, n1323, n1324, n1325, n1326, n1335, n1336, n1337,
         n1338, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1363,
         n1364, n1365, n1366, n1375, n1376, n1377, n1378, n1379, n1380, n1389,
         n1390, n1391, n1392, n1401, n1402, n1403, n1404, n1405, n1406, n1408,
         n1409, n1410, n1411, n1412, n1413, n1422, n1423, n1424, n1425, n1434,
         n1435, n1436, n1437, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1462, n1463, n1464, n1465, n1474, n1475, n1476, n1477, n1478,
         n1479, n1488, n1489, n1490, n1491, n1500, n1501, n1502, n1504, n1505,
         n1506, n1507, n1518, n1519, n1520, n1521, n1523, n1524, n1525, n1526,
         n1527, n1528, n1537, n1538, n1539, n1540, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1565, n1566, n1567, n1568, n1577, n1578,
         n1579, n1580, n1581, n1582, n1591, n1592, n1593, n1594, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1611, n1612, n1613, n1614, n1615,
         n1616, n1625, n1626, n1627, n1628, n1637, n1638, n1639, n1640, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1665, n1666, n1667,
         n1668, n1677, n1678, n1679, n1680, n1681, n1682, n1691, n1692, n1693,
         n1694, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1719,
         n1720, n1721, n1722, n1731, n1732, n1733, n1734, n1735, n1736, n1745,
         n1746, n1747, n1748, n1758, n1759, n1760, n1762, n1763, n1764, n1765,
         n1766, n1767, n1776, n1777, n1778, n1779, n1780, n1789, n1790, n1791,
         n1792, n1801, n1802, n1803, n1804, n1805, n1806, n1808, n1809, n1811,
         n1812, n1813, n1814, n1823, n1824, n1825, n1826, n1835, n1836, n1837,
         n1838, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1863,
         n1864, n1865, n1866, n1875, n1876, n1877, n1878, n1879, n1880, n1889,
         n1890, n1891, n1892, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1909, n1911, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1931, n1932, n1937, n1938, n1939, n1940, n1949, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1967, n1968, n1969,
         n1970, n1979, n1980, n1981, n1982, n1983, n1984, n1993, n1994, n1995,
         n1996, n2007, n2008, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2066, n2067, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2093, n2094, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2116, n2117, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2140, n2141, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2164, n2165, n2168, n2169, n2171, n2172, n2173,
         n2174, n2176, n2177, n2191, n2192, n2193, n2194, n2195, n2196, n2198,
         n2199, n2214, n2215, n2216, n2217, n2218, n2219, n2234, n2235, n2292,
         n2381, n2383, n2384, n2385, n2387, n2388, n2401, n2404, n2453, n2502,
         n2567, n2624, n2714, n2755, n2844, n2846, n2847, n2848, n2850, n2851,
         n2864, n2867, n2916, n2965, n3030, n3047, n3136, n3162, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311;
  wire   [4:0] wrt_ptr;
  wire   [14:0] dataout_stg_1;
  wire   [3:0] lenout_stg_1;
  wire   [1037:0] buffer;
  wire   [9:0] rd_ptr;
  wire   [9:1] \add_121/carry ;
  wire   [4:2] \add_44/carry ;

  CAOR2X1 U3 ( .A(wrt_ptr[4]), .B(n7174), .C(pushin), .D(N114), .Z(n3164) );
  CAOR2X1 U4 ( .A(wrt_ptr[3]), .B(n7174), .C(N113), .D(pushin), .Z(n3165) );
  CAOR2X1 U6 ( .A(wrt_ptr[2]), .B(n7174), .C(N112), .D(pushin), .Z(n3166) );
  CAOR2X1 U7 ( .A(wrt_ptr[1]), .B(n7174), .C(N111), .D(pushin), .Z(n3167) );
  CAOR2X1 U8 ( .A(wrt_ptr[0]), .B(n7174), .C(n7220), .D(pushin), .Z(n3168) );
  CAOR2X1 U9 ( .A(n4267), .B(n4), .C(n5), .D(n7218), .Z(n3175) );
  CAOR2X1 U22 ( .A(n44), .B(n8295), .C(n46), .D(n8291), .Z(n24) );
  CAOR1X1 U38 ( .A(n8302), .B(n89), .C(n90), .Z(n71) );
  CAOR2X1 U52 ( .A(n8016), .B(n7097), .C(n7760), .D(n40), .Z(n117) );
  CAOR2X1 U58 ( .A(n101), .B(n7171), .C(n131), .D(n7172), .Z(n130) );
  CAOR2X1 U66 ( .A(n144), .B(n8303), .C(n145), .D(n39), .Z(n140) );
  CAOR1X1 U85 ( .A(n4269), .B(n7092), .C(n170), .Z(n3180) );
  CAOR1X1 U103 ( .A(n4268), .B(n7092), .C(n7169), .Z(n3181) );
  COAN1X1 U110 ( .A(rd_ptr[3]), .B(n7247), .C(n209), .Z(n13) );
  CAN4X1 U163 ( .A(n272), .B(n273), .C(n274), .D(n275), .Z(n68) );
  CAOR1X1 U179 ( .A(n8293), .B(n290), .C(n291), .Z(n155) );
  CAN4X1 U181 ( .A(n293), .B(n294), .C(n295), .D(n296), .Z(n111) );
  CAOR1X1 U215 ( .A(n8293), .B(n332), .C(n333), .Z(n207) );
  CAN4X1 U257 ( .A(n376), .B(n377), .C(n378), .D(n379), .Z(n375) );
  COR4X1 U264 ( .A(n392), .B(n393), .C(n394), .D(n395), .Z(n340) );
  COR4X1 U270 ( .A(n409), .B(n410), .C(n411), .D(n412), .Z(n342) );
  COR4X1 U275 ( .A(n421), .B(n422), .C(n423), .D(n424), .Z(n341) );
  COR4X1 U283 ( .A(n437), .B(n438), .C(n439), .D(n440), .Z(n436) );
  COR4X1 U288 ( .A(n449), .B(n450), .C(n451), .D(n452), .Z(n435) );
  COR4X1 U294 ( .A(n463), .B(n464), .C(n465), .D(n466), .Z(n462) );
  COR4X1 U299 ( .A(n475), .B(n476), .C(n477), .D(n478), .Z(n461) );
  COAN1X1 U304 ( .A(n8296), .B(n160), .C(n488), .Z(n332) );
  COR4X1 U313 ( .A(n497), .B(n498), .C(n499), .D(n500), .Z(n166) );
  COR4X1 U332 ( .A(n538), .B(n539), .C(n540), .D(n541), .Z(n537) );
  COR4X1 U337 ( .A(n550), .B(n551), .C(n552), .D(n553), .Z(n536) );
  COR4X1 U343 ( .A(n564), .B(n565), .C(n566), .D(n567), .Z(n563) );
  COR4X1 U348 ( .A(n576), .B(n577), .C(n578), .D(n579), .Z(n562) );
  CAOR1X1 U355 ( .A(rd_ptr[3]), .B(n290), .C(n589), .Z(n588) );
  COR4X1 U364 ( .A(n598), .B(n599), .C(n600), .D(n601), .Z(n298) );
  COR4X1 U370 ( .A(n610), .B(n611), .C(n612), .D(n613), .Z(n300) );
  COR4X1 U375 ( .A(n622), .B(n623), .C(n624), .D(n625), .Z(n299) );
  COR4X1 U383 ( .A(n638), .B(n639), .C(n640), .D(n641), .Z(n637) );
  COR4X1 U388 ( .A(n650), .B(n651), .C(n652), .D(n653), .Z(n636) );
  COR4X1 U394 ( .A(n664), .B(n665), .C(n666), .D(n667), .Z(n663) );
  COR4X1 U399 ( .A(n676), .B(n677), .C(n678), .D(n679), .Z(n662) );
  CAOR2X1 U404 ( .A(n115), .B(rd_ptr[4]), .C(n8296), .D(n688), .Z(n290) );
  COR4X1 U426 ( .A(n724), .B(n725), .C(n726), .D(n727), .Z(n126) );
  COR4X1 U434 ( .A(n740), .B(n741), .C(n742), .D(n743), .Z(n739) );
  COR4X1 U439 ( .A(n752), .B(n753), .C(n754), .D(n755), .Z(n738) );
  COR4X1 U445 ( .A(n766), .B(n767), .C(n768), .D(n769), .Z(n765) );
  COR4X1 U450 ( .A(n778), .B(n779), .C(n780), .D(n781), .Z(n764) );
  COR4X1 U464 ( .A(n799), .B(n800), .C(n801), .D(n802), .Z(n217) );
  COR4X1 U470 ( .A(n811), .B(n812), .C(n813), .D(n814), .Z(n219) );
  COR4X1 U475 ( .A(n823), .B(n824), .C(n825), .D(n826), .Z(n218) );
  COR4X1 U482 ( .A(n839), .B(n840), .C(n841), .D(n842), .Z(n838) );
  COR4X1 U487 ( .A(n851), .B(n852), .C(n853), .D(n854), .Z(n837) );
  COR4X1 U493 ( .A(n865), .B(n866), .C(n867), .D(n868), .Z(n864) );
  COR4X1 U498 ( .A(n877), .B(n878), .C(n879), .D(n880), .Z(n863) );
  COR4X1 U521 ( .A(n926), .B(n927), .C(n928), .D(n929), .Z(n904) );
  COR4X1 U531 ( .A(n947), .B(n948), .C(n949), .D(n950), .Z(n946) );
  COR4X1 U536 ( .A(n959), .B(n960), .C(n961), .D(n962), .Z(n945) );
  COR4X1 U542 ( .A(n973), .B(n974), .C(n975), .D(n976), .Z(n972) );
  COR4X1 U547 ( .A(n985), .B(n986), .C(n987), .D(n988), .Z(n971) );
  COR4X1 U562 ( .A(n1007), .B(n1008), .C(n1009), .D(n1010), .Z(n255) );
  COR4X1 U568 ( .A(n1019), .B(n1020), .C(n1021), .D(n1022), .Z(n257) );
  COR4X1 U573 ( .A(n1031), .B(n1032), .C(n1033), .D(n1034), .Z(n256) );
  COR4X1 U580 ( .A(n1047), .B(n1048), .C(n1049), .D(n1050), .Z(n1046) );
  COR4X1 U585 ( .A(n1059), .B(n1060), .C(n1061), .D(n1062), .Z(n1045) );
  COR4X1 U591 ( .A(n1073), .B(n1074), .C(n1075), .D(n1076), .Z(n1072) );
  COR4X1 U596 ( .A(n1085), .B(n1086), .C(n1087), .D(n1088), .Z(n1071) );
  COR4X1 U604 ( .A(n1101), .B(n1102), .C(n1103), .D(n1104), .Z(n1100) );
  COR4X1 U609 ( .A(n1113), .B(n1114), .C(n1115), .D(n1116), .Z(n1099) );
  COR4X1 U615 ( .A(n1127), .B(n1128), .C(n1129), .D(n1130), .Z(n1126) );
  COR4X1 U620 ( .A(n1139), .B(n1140), .C(n1141), .D(n1142), .Z(n1125) );
  COR4X1 U632 ( .A(n1158), .B(n1159), .C(n1160), .D(n1161), .Z(n36) );
  CAN4X1 U662 ( .A(n1205), .B(n1206), .C(n1207), .D(n1208), .Z(n1204) );
  COR4X1 U669 ( .A(n1212), .B(n1213), .C(n1214), .D(n1215), .Z(n363) );
  COR4X1 U675 ( .A(n1224), .B(n1225), .C(n1226), .D(n1227), .Z(n364) );
  COR4X1 U680 ( .A(n1236), .B(n1237), .C(n1238), .D(n1239), .Z(n362) );
  COR4X1 U688 ( .A(n1252), .B(n1253), .C(n1254), .D(n1255), .Z(n1251) );
  COR4X1 U693 ( .A(n1264), .B(n1265), .C(n1266), .D(n1267), .Z(n1250) );
  COR4X1 U699 ( .A(n1278), .B(n1279), .C(n1280), .D(n1281), .Z(n1277) );
  COR4X1 U704 ( .A(n1290), .B(n1291), .C(n1292), .D(n1293), .Z(n1276) );
  COR4X1 U719 ( .A(n1311), .B(n1312), .C(n1313), .D(n1314), .Z(n193) );
  COR4X1 U725 ( .A(n1323), .B(n1324), .C(n1325), .D(n1326), .Z(n197) );
  COR4X1 U730 ( .A(n1335), .B(n1336), .C(n1337), .D(n1338), .Z(n195) );
  COR4X1 U737 ( .A(n1351), .B(n1352), .C(n1353), .D(n1354), .Z(n1350) );
  COR4X1 U742 ( .A(n1363), .B(n1364), .C(n1365), .D(n1366), .Z(n1349) );
  COR4X1 U748 ( .A(n1377), .B(n1378), .C(n1379), .D(n1380), .Z(n1376) );
  COR4X1 U753 ( .A(n1389), .B(n1390), .C(n1391), .D(n1392), .Z(n1375) );
  CAOR2X1 U761 ( .A(n8292), .B(n271), .C(n8291), .D(n1402), .Z(n1401) );
  COR4X1 U769 ( .A(n1410), .B(n1411), .C(n1412), .D(n1413), .Z(n277) );
  COR4X1 U775 ( .A(n1422), .B(n1423), .C(n1424), .D(n1425), .Z(n279) );
  COR4X1 U780 ( .A(n1434), .B(n1435), .C(n1436), .D(n1437), .Z(n278) );
  COR4X1 U787 ( .A(n1450), .B(n1451), .C(n1452), .D(n1453), .Z(n1449) );
  COR4X1 U792 ( .A(n1462), .B(n1463), .C(n1464), .D(n1465), .Z(n1448) );
  COR4X1 U798 ( .A(n1476), .B(n1477), .C(n1478), .D(n1479), .Z(n1475) );
  COR4X1 U803 ( .A(n1488), .B(n1489), .C(n1490), .D(n1491), .Z(n1474) );
  COR4X1 U836 ( .A(n1553), .B(n1554), .C(n1555), .D(n1556), .Z(n1552) );
  COR4X1 U841 ( .A(n1565), .B(n1566), .C(n1567), .D(n1568), .Z(n1551) );
  COR4X1 U847 ( .A(n1579), .B(n1580), .C(n1581), .D(n1582), .Z(n1578) );
  COR4X1 U852 ( .A(n1591), .B(n1592), .C(n1593), .D(n1594), .Z(n1577) );
  COR4X1 U867 ( .A(n1613), .B(n1614), .C(n1615), .D(n1616), .Z(n324) );
  COR4X1 U873 ( .A(n1625), .B(n1626), .C(n1627), .D(n1628), .Z(n326) );
  COR4X1 U878 ( .A(n1637), .B(n1638), .C(n1639), .D(n1640), .Z(n325) );
  COR4X1 U885 ( .A(n1653), .B(n1654), .C(n1655), .D(n1656), .Z(n1652) );
  COR4X1 U890 ( .A(n1665), .B(n1666), .C(n1667), .D(n1668), .Z(n1651) );
  COR4X1 U896 ( .A(n1679), .B(n1680), .C(n1681), .D(n1682), .Z(n1678) );
  COR4X1 U901 ( .A(n1691), .B(n1692), .C(n1693), .D(n1694), .Z(n1677) );
  COR4X1 U909 ( .A(n1707), .B(n1708), .C(n1709), .D(n1710), .Z(n1706) );
  COR4X1 U914 ( .A(n1719), .B(n1720), .C(n1721), .D(n1722), .Z(n1705) );
  COR4X1 U920 ( .A(n1733), .B(n1734), .C(n1735), .D(n1736), .Z(n1732) );
  COR4X1 U925 ( .A(n1745), .B(n1746), .C(n1747), .D(n1748), .Z(n1731) );
  COR4X1 U939 ( .A(n1764), .B(n1765), .C(n1766), .D(n1767), .Z(n144) );
  COR4X1 U971 ( .A(n1811), .B(n1812), .C(n1813), .D(n1814), .Z(n236) );
  COR4X1 U977 ( .A(n1823), .B(n1824), .C(n1825), .D(n1826), .Z(n238) );
  COR4X1 U982 ( .A(n1835), .B(n1836), .C(n1837), .D(n1838), .Z(n237) );
  COR4X1 U991 ( .A(n1851), .B(n1852), .C(n1853), .D(n1854), .Z(n1850) );
  COR4X1 U996 ( .A(n1863), .B(n1864), .C(n1865), .D(n1866), .Z(n1849) );
  COR4X1 U1002 ( .A(n1877), .B(n1878), .C(n1879), .D(n1880), .Z(n1876) );
  COR4X1 U1007 ( .A(n1889), .B(n1890), .C(n1891), .D(n1892), .Z(n1875) );
  COR4X1 U1041 ( .A(n1937), .B(n1938), .C(n1939), .D(n1940), .Z(n1915) );
  COR4X1 U1057 ( .A(n1955), .B(n1956), .C(n1957), .D(n1958), .Z(n1954) );
  COR4X1 U1064 ( .A(n1967), .B(n1968), .C(n1969), .D(n1970), .Z(n1953) );
  COR4X1 U1073 ( .A(n1981), .B(n1982), .C(n1983), .D(n1984), .Z(n1980) );
  COR4X1 U1081 ( .A(n1993), .B(n1994), .C(n1995), .D(n1996), .Z(n1979) );
  CAOR2X1 U1111 ( .A(N16596), .B(n3173), .C(n4), .D(rd_ptr[6]), .Z(n3193) );
  CAOR2X1 U1112 ( .A(N16595), .B(n6164), .C(n7092), .D(rd_ptr[5]), .Z(n3194)
         );
  CAOR2X1 U1113 ( .A(N16594), .B(n6165), .C(n7091), .D(rd_ptr[4]), .Z(n3195)
         );
  CAOR2X1 U1114 ( .A(N16593), .B(n3173), .C(n4), .D(rd_ptr[3]), .Z(n3196) );
  CAOR2X1 U1115 ( .A(N16592), .B(n6164), .C(n7092), .D(rd_ptr[2]), .Z(n3197)
         );
  CAOR2X1 U1116 ( .A(N16591), .B(n6165), .C(n4), .D(rd_ptr[1]), .Z(n3198) );
  CAOR2X1 U1117 ( .A(N16590), .B(n3173), .C(n4), .D(rd_ptr[0]), .Z(n3199) );
  CAN3X2 U2833 ( .A(n7221), .B(n7222), .C(wrt_ptr[3]), .Z(n2107) );
  CAN3X2 U2966 ( .A(wrt_ptr[3]), .B(n7222), .C(wrt_ptr[1]), .Z(n2112) );
  CAN3X2 U3100 ( .A(wrt_ptr[3]), .B(n7221), .C(wrt_ptr[2]), .Z(n2130) );
  CAN3X2 U3168 ( .A(pushin), .B(n7220), .C(wrt_ptr[4]), .Z(n2155) );
  CAN3X2 U3254 ( .A(wrt_ptr[2]), .B(wrt_ptr[3]), .C(wrt_ptr[1]), .Z(n2135) );
  CAN3X2 U3255 ( .A(wrt_ptr[4]), .B(pushin), .C(wrt_ptr[0]), .Z(n2158) );
  CFA1X1 \add_121/U1_1  ( .A(rd_ptr[1]), .B(n6161), .CI(\add_121/carry [1]), 
        .CO(\add_121/carry [2]), .S(N16591) );
  CFA1X1 \add_121/U1_2  ( .A(rd_ptr[2]), .B(n6162), .CI(\add_121/carry [2]), 
        .CO(\add_121/carry [3]), .S(N16592) );
  CFA1X1 \add_121/U1_3  ( .A(rd_ptr[3]), .B(n6163), .CI(\add_121/carry [3]), 
        .CO(\add_121/carry [4]), .S(N16593) );
  CHA1X1 \add_44/U1_1_1  ( .A(wrt_ptr[1]), .B(wrt_ptr[0]), .CO(
        \add_44/carry [2]), .S(N111) );
  CHA1X1 \add_44/U1_1_2  ( .A(wrt_ptr[2]), .B(\add_44/carry [2]), .CO(
        \add_44/carry [3]), .S(N112) );
  CHA1X1 \add_44/U1_1_3  ( .A(wrt_ptr[3]), .B(\add_44/carry [3]), .CO(
        \add_44/carry [4]), .S(N113) );
  CFD1QXL \dataout_stg_1_reg[9]  ( .D(n3180), .CP(clk), .Q(dataout_stg_1[9])
         );
  CFD1QXL \dataout_stg_1_reg[8]  ( .D(n3181), .CP(clk), .Q(dataout_stg_1[8])
         );
  CFD1QXL \dataout_stg_1_reg[14]  ( .D(n3175), .CP(clk), .Q(dataout_stg_1[14])
         );
  CFD1QXL \dataout_stg_1_reg[12]  ( .D(n3177), .CP(clk), .Q(dataout_stg_1[12])
         );
  CFD1QXL \dataout_stg_1_reg[11]  ( .D(n3178), .CP(clk), .Q(dataout_stg_1[11])
         );
  CFD1QXL \dataout_stg_1_reg[13]  ( .D(n3176), .CP(clk), .Q(dataout_stg_1[13])
         );
  CFD1QXL \dataout_stg_1_reg[10]  ( .D(n3179), .CP(clk), .Q(dataout_stg_1[10])
         );
  CFD1QXL \dataout_stg_1_reg[7]  ( .D(n3182), .CP(clk), .Q(dataout_stg_1[7])
         );
  CFD1QXL \dataout_stg_1_reg[2]  ( .D(n3187), .CP(clk), .Q(dataout_stg_1[2])
         );
  CFD1QXL \dataout_stg_1_reg[6]  ( .D(n3183), .CP(clk), .Q(dataout_stg_1[6])
         );
  CFD1QXL \dataout_stg_1_reg[5]  ( .D(n3184), .CP(clk), .Q(dataout_stg_1[5])
         );
  CFD1QXL \dataout_stg_1_reg[4]  ( .D(n3185), .CP(clk), .Q(dataout_stg_1[4])
         );
  CFD1QXL \dataout_stg_1_reg[3]  ( .D(n3186), .CP(clk), .Q(dataout_stg_1[3])
         );
  CFD1QXL \dataout_stg_1_reg[1]  ( .D(n3188), .CP(clk), .Q(dataout_stg_1[1])
         );
  CFD1QXL \buffer_reg[1037]  ( .D(n4237), .CP(clk), .Q(buffer[1037]) );
  CFD2QXL \lenout_stg_2_reg[3]  ( .D(n4260), .CP(clk), .CD(n7173), .Q(
        lenout[3]) );
  CFD2QXL \lenout_stg_2_reg[2]  ( .D(n4258), .CP(clk), .CD(n7173), .Q(
        lenout[2]) );
  CFD2QXL \lenout_stg_2_reg[1]  ( .D(n4256), .CP(clk), .CD(n7173), .Q(
        lenout[1]) );
  CFD2QXL \lenout_stg_2_reg[0]  ( .D(n4254), .CP(clk), .CD(n7173), .Q(
        lenout[0]) );
  CFD1QXL \dataout_stg_1_reg[0]  ( .D(n3189), .CP(clk), .Q(dataout_stg_1[0])
         );
  CFD1QXL \buffer_reg[908]  ( .D(n4108), .CP(clk), .Q(buffer[908]) );
  CFD1QXL \buffer_reg[653]  ( .D(n3853), .CP(clk), .Q(buffer[653]) );
  CFD1QXL \buffer_reg[652]  ( .D(n3852), .CP(clk), .Q(buffer[652]) );
  CFD1QXL \buffer_reg[651]  ( .D(n3851), .CP(clk), .Q(buffer[651]) );
  CFD1QXL \buffer_reg[650]  ( .D(n3850), .CP(clk), .Q(buffer[650]) );
  CFD1QXL \buffer_reg[649]  ( .D(n3849), .CP(clk), .Q(buffer[649]) );
  CFD1QXL \buffer_reg[648]  ( .D(n3848), .CP(clk), .Q(buffer[648]) );
  CFD1QXL \buffer_reg[647]  ( .D(n3847), .CP(clk), .Q(buffer[647]) );
  CFD1QXL \buffer_reg[646]  ( .D(n3846), .CP(clk), .Q(buffer[646]) );
  CFD1QXL \buffer_reg[645]  ( .D(n3845), .CP(clk), .Q(buffer[645]) );
  CFD1QXL \buffer_reg[644]  ( .D(n3844), .CP(clk), .Q(buffer[644]) );
  CFD1QXL \buffer_reg[643]  ( .D(n3843), .CP(clk), .Q(buffer[643]) );
  CFD1QXL \buffer_reg[642]  ( .D(n3842), .CP(clk), .Q(buffer[642]) );
  CFD1QXL \buffer_reg[641]  ( .D(n3841), .CP(clk), .Q(buffer[641]) );
  CFD1QXL \buffer_reg[640]  ( .D(n3840), .CP(clk), .Q(buffer[640]) );
  CFD1QXL \buffer_reg[140]  ( .D(n3340), .CP(clk), .Q(buffer[140]) );
  CFD1QXL \buffer_reg[397]  ( .D(n3597), .CP(clk), .Q(buffer[397]) );
  CFD1QXL \buffer_reg[395]  ( .D(n3595), .CP(clk), .Q(buffer[395]) );
  CFD1QXL \buffer_reg[394]  ( .D(n3594), .CP(clk), .Q(buffer[394]) );
  CFD1QXL \buffer_reg[392]  ( .D(n3592), .CP(clk), .Q(buffer[392]) );
  CFD1QXL \buffer_reg[391]  ( .D(n3591), .CP(clk), .Q(buffer[391]) );
  CFD1QXL \buffer_reg[390]  ( .D(n3590), .CP(clk), .Q(buffer[390]) );
  CFD1QXL \buffer_reg[389]  ( .D(n3589), .CP(clk), .Q(buffer[389]) );
  CFD1QXL \buffer_reg[388]  ( .D(n3588), .CP(clk), .Q(buffer[388]) );
  CFD1QXL \buffer_reg[387]  ( .D(n3587), .CP(clk), .Q(buffer[387]) );
  CFD1QXL \buffer_reg[386]  ( .D(n3586), .CP(clk), .Q(buffer[386]) );
  CFD1QXL \buffer_reg[385]  ( .D(n3585), .CP(clk), .Q(buffer[385]) );
  CFD1QXL \buffer_reg[384]  ( .D(n3584), .CP(clk), .Q(buffer[384]) );
  CFD1QXL \buffer_reg[141]  ( .D(n3341), .CP(clk), .Q(buffer[141]) );
  CFD1QXL \buffer_reg[139]  ( .D(n3339), .CP(clk), .Q(buffer[139]) );
  CFD1QXL \buffer_reg[138]  ( .D(n3338), .CP(clk), .Q(buffer[138]) );
  CFD1QXL \buffer_reg[136]  ( .D(n3336), .CP(clk), .Q(buffer[136]) );
  CFD1QXL \buffer_reg[135]  ( .D(n3335), .CP(clk), .Q(buffer[135]) );
  CFD1QXL \buffer_reg[134]  ( .D(n3334), .CP(clk), .Q(buffer[134]) );
  CFD1QXL \buffer_reg[133]  ( .D(n3333), .CP(clk), .Q(buffer[133]) );
  CFD1QXL \buffer_reg[132]  ( .D(n3332), .CP(clk), .Q(buffer[132]) );
  CFD1QXL \buffer_reg[131]  ( .D(n3331), .CP(clk), .Q(buffer[131]) );
  CFD1QXL \buffer_reg[130]  ( .D(n3330), .CP(clk), .Q(buffer[130]) );
  CFD1QXL \buffer_reg[128]  ( .D(n3328), .CP(clk), .Q(buffer[128]) );
  CFD1QXL \buffer_reg[1025]  ( .D(n4225), .CP(clk), .Q(buffer[1025]) );
  CFD1QXL \buffer_reg[393]  ( .D(n3593), .CP(clk), .Q(buffer[393]) );
  CFD1QXL \buffer_reg[396]  ( .D(n3596), .CP(clk), .Q(buffer[396]) );
  CFD1QXL \buffer_reg[909]  ( .D(n4109), .CP(clk), .Q(buffer[909]) );
  CFD1QXL \buffer_reg[907]  ( .D(n4107), .CP(clk), .Q(buffer[907]) );
  CFD1QXL \buffer_reg[906]  ( .D(n4106), .CP(clk), .Q(buffer[906]) );
  CFD1QXL \buffer_reg[905]  ( .D(n4105), .CP(clk), .Q(buffer[905]) );
  CFD1QXL \buffer_reg[904]  ( .D(n4104), .CP(clk), .Q(buffer[904]) );
  CFD1QXL \buffer_reg[903]  ( .D(n4103), .CP(clk), .Q(buffer[903]) );
  CFD1QXL \buffer_reg[902]  ( .D(n4102), .CP(clk), .Q(buffer[902]) );
  CFD1QXL \buffer_reg[901]  ( .D(n4101), .CP(clk), .Q(buffer[901]) );
  CFD1QXL \buffer_reg[900]  ( .D(n4100), .CP(clk), .Q(buffer[900]) );
  CFD1QXL \buffer_reg[899]  ( .D(n4099), .CP(clk), .Q(buffer[899]) );
  CFD1QXL \buffer_reg[898]  ( .D(n4098), .CP(clk), .Q(buffer[898]) );
  CFD1QXL \buffer_reg[897]  ( .D(n4097), .CP(clk), .Q(buffer[897]) );
  CFD1QXL \buffer_reg[896]  ( .D(n4096), .CP(clk), .Q(buffer[896]) );
  CFD1QXL \buffer_reg[1034]  ( .D(n4234), .CP(clk), .Q(buffer[1034]) );
  CFD1QXL \buffer_reg[1033]  ( .D(n4233), .CP(clk), .Q(buffer[1033]) );
  CFD1QXL \buffer_reg[1032]  ( .D(n4232), .CP(clk), .Q(buffer[1032]) );
  CFD1QXL \buffer_reg[1031]  ( .D(n4231), .CP(clk), .Q(buffer[1031]) );
  CFD1QXL \buffer_reg[1030]  ( .D(n4230), .CP(clk), .Q(buffer[1030]) );
  CFD1QXL \buffer_reg[1029]  ( .D(n4229), .CP(clk), .Q(buffer[1029]) );
  CFD1QXL \buffer_reg[1028]  ( .D(n4228), .CP(clk), .Q(buffer[1028]) );
  CFD1QXL \buffer_reg[1027]  ( .D(n4227), .CP(clk), .Q(buffer[1027]) );
  CFD1QXL \buffer_reg[1026]  ( .D(n4226), .CP(clk), .Q(buffer[1026]) );
  CFD1QXL \buffer_reg[1024]  ( .D(n4224), .CP(clk), .Q(buffer[1024]) );
  CFD1QXL \buffer_reg[780]  ( .D(n3980), .CP(clk), .Q(buffer[780]) );
  CFD1QXL \buffer_reg[769]  ( .D(n3969), .CP(clk), .Q(buffer[769]) );
  CFD1QXL \buffer_reg[522]  ( .D(n3722), .CP(clk), .Q(buffer[522]) );
  CFD1QXL \buffer_reg[520]  ( .D(n3720), .CP(clk), .Q(buffer[520]) );
  CFD1QXL \buffer_reg[518]  ( .D(n3718), .CP(clk), .Q(buffer[518]) );
  CFD1QXL \buffer_reg[516]  ( .D(n3716), .CP(clk), .Q(buffer[516]) );
  CFD1QXL \buffer_reg[514]  ( .D(n3714), .CP(clk), .Q(buffer[514]) );
  CFD1QXL \buffer_reg[512]  ( .D(n3712), .CP(clk), .Q(buffer[512]) );
  CFD1QXL \buffer_reg[525]  ( .D(n3725), .CP(clk), .Q(buffer[525]) );
  CFD1QXL \buffer_reg[521]  ( .D(n3721), .CP(clk), .Q(buffer[521]) );
  CFD1QXL \buffer_reg[519]  ( .D(n3719), .CP(clk), .Q(buffer[519]) );
  CFD1QXL \buffer_reg[517]  ( .D(n3717), .CP(clk), .Q(buffer[517]) );
  CFD1QXL \buffer_reg[515]  ( .D(n3715), .CP(clk), .Q(buffer[515]) );
  CFD1QXL \buffer_reg[513]  ( .D(n3713), .CP(clk), .Q(buffer[513]) );
  CFD1QXL \buffer_reg[266]  ( .D(n3466), .CP(clk), .Q(buffer[266]) );
  CFD1QXL \buffer_reg[264]  ( .D(n3464), .CP(clk), .Q(buffer[264]) );
  CFD1QXL \buffer_reg[262]  ( .D(n3462), .CP(clk), .Q(buffer[262]) );
  CFD1QXL \buffer_reg[260]  ( .D(n3460), .CP(clk), .Q(buffer[260]) );
  CFD1QXL \buffer_reg[258]  ( .D(n3458), .CP(clk), .Q(buffer[258]) );
  CFD1QXL \buffer_reg[256]  ( .D(n3456), .CP(clk), .Q(buffer[256]) );
  CFD1QXL \buffer_reg[269]  ( .D(n3469), .CP(clk), .Q(buffer[269]) );
  CFD1QXL \buffer_reg[265]  ( .D(n3465), .CP(clk), .Q(buffer[265]) );
  CFD1QXL \buffer_reg[263]  ( .D(n3463), .CP(clk), .Q(buffer[263]) );
  CFD1QXL \buffer_reg[261]  ( .D(n3461), .CP(clk), .Q(buffer[261]) );
  CFD1QXL \buffer_reg[259]  ( .D(n3459), .CP(clk), .Q(buffer[259]) );
  CFD1QXL \buffer_reg[257]  ( .D(n3457), .CP(clk), .Q(buffer[257]) );
  CFD1QXL \buffer_reg[781]  ( .D(n3981), .CP(clk), .Q(buffer[781]) );
  CFD1QXL \buffer_reg[777]  ( .D(n3977), .CP(clk), .Q(buffer[777]) );
  CFD1QXL \buffer_reg[775]  ( .D(n3975), .CP(clk), .Q(buffer[775]) );
  CFD1QXL \buffer_reg[773]  ( .D(n3973), .CP(clk), .Q(buffer[773]) );
  CFD1QXL \buffer_reg[771]  ( .D(n3971), .CP(clk), .Q(buffer[771]) );
  CFD1QXL \buffer_reg[778]  ( .D(n3978), .CP(clk), .Q(buffer[778]) );
  CFD1QXL \buffer_reg[776]  ( .D(n3976), .CP(clk), .Q(buffer[776]) );
  CFD1QXL \buffer_reg[774]  ( .D(n3974), .CP(clk), .Q(buffer[774]) );
  CFD1QXL \buffer_reg[772]  ( .D(n3972), .CP(clk), .Q(buffer[772]) );
  CFD1QXL \buffer_reg[770]  ( .D(n3970), .CP(clk), .Q(buffer[770]) );
  CFD1QXL \buffer_reg[768]  ( .D(n3968), .CP(clk), .Q(buffer[768]) );
  CFD1QXL \rd_ptr_reg[1]  ( .D(n3198), .CP(clk), .Q(rd_ptr[1]) );
  CFD1QXL \rd_ptr_reg[2]  ( .D(n3197), .CP(clk), .Q(rd_ptr[2]) );
  CFD2QXL \wrt_ptr_reg[0]  ( .D(n3168), .CP(clk), .CD(n7173), .Q(wrt_ptr[0])
         );
  CFD1QXL \rd_ptr_reg[3]  ( .D(n3196), .CP(clk), .Q(rd_ptr[3]) );
  CFD1QXL \rd_ptr_reg[4]  ( .D(n3195), .CP(clk), .Q(rd_ptr[4]) );
  CFD2QXL \wrt_ptr_reg[4]  ( .D(n3164), .CP(clk), .CD(n7173), .Q(wrt_ptr[4])
         );
  CFD2QXL \wrt_ptr_reg[2]  ( .D(n3166), .CP(clk), .CD(n7173), .Q(wrt_ptr[2])
         );
  CFD2QXL \wrt_ptr_reg[1]  ( .D(n3167), .CP(clk), .CD(n7173), .Q(wrt_ptr[1])
         );
  CFD2QXL \wrt_ptr_reg[3]  ( .D(n3165), .CP(clk), .CD(n7173), .Q(wrt_ptr[3])
         );
  CFD1QXL \buffer_reg[129]  ( .D(n3329), .CP(clk), .Q(buffer[129]) );
  CFD1QXL \buffer_reg[137]  ( .D(n3337), .CP(clk), .Q(buffer[137]) );
  CFD1QXL \rd_ptr_reg[5]  ( .D(n3194), .CP(clk), .Q(rd_ptr[5]) );
  CFD1QXL \rd_ptr_reg[0]  ( .D(n3199), .CP(clk), .Q(rd_ptr[0]) );
  CFD1QXL \rd_ptr_reg[6]  ( .D(n3193), .CP(clk), .Q(rd_ptr[6]) );
  CFD1QXL \lenout_stg_1_reg[3]  ( .D(N121), .CP(clk), .Q(lenout_stg_1[3]) );
  CFD1QXL \lenout_stg_1_reg[2]  ( .D(N120), .CP(clk), .Q(lenout_stg_1[2]) );
  CFD1QXL \lenout_stg_1_reg[1]  ( .D(N119), .CP(clk), .Q(lenout_stg_1[1]) );
  CFD1QXL \lenout_stg_1_reg[0]  ( .D(N118), .CP(clk), .Q(lenout_stg_1[0]) );
  CFD1QXL pushout_stg_1_reg ( .D(n6165), .CP(clk), .Q(pushout_stg_1) );
  CFD2QXL pushout_stg_2_reg ( .D(n4252), .CP(clk), .CD(n7173), .Q(pushout) );
  CFD2QXL \dataout_stg_2_reg[14]  ( .D(n4251), .CP(clk), .CD(n7173), .Q(
        dataout[14]) );
  CFD2QXL \dataout_stg_2_reg[13]  ( .D(n4250), .CP(clk), .CD(n7173), .Q(
        dataout[13]) );
  CFD2QXL \dataout_stg_2_reg[12]  ( .D(n4249), .CP(clk), .CD(n7173), .Q(
        dataout[12]) );
  CFD2QXL \dataout_stg_2_reg[11]  ( .D(n4248), .CP(clk), .CD(n7173), .Q(
        dataout[11]) );
  CFD2QXL \dataout_stg_2_reg[10]  ( .D(n4247), .CP(clk), .CD(n7173), .Q(
        dataout[10]) );
  CFD2QXL \dataout_stg_2_reg[9]  ( .D(n4246), .CP(clk), .CD(n7173), .Q(
        dataout[9]) );
  CFD2QXL \dataout_stg_2_reg[8]  ( .D(n4245), .CP(clk), .CD(n7173), .Q(
        dataout[8]) );
  CFD2QXL \dataout_stg_2_reg[7]  ( .D(n4244), .CP(clk), .CD(n7173), .Q(
        dataout[7]) );
  CFD2QXL \dataout_stg_2_reg[6]  ( .D(n6141), .CP(clk), .CD(n7173), .Q(
        dataout[6]) );
  CFD2QXL \dataout_stg_2_reg[5]  ( .D(n4292), .CP(clk), .CD(n7173), .Q(
        dataout[5]) );
  CFD2QXL \dataout_stg_2_reg[4]  ( .D(n4290), .CP(clk), .CD(n7173), .Q(
        dataout[4]) );
  CFD2QXL \dataout_stg_2_reg[3]  ( .D(n4288), .CP(clk), .CD(n7173), .Q(
        dataout[3]) );
  CFD2QXL \dataout_stg_2_reg[2]  ( .D(n4286), .CP(clk), .CD(n7173), .Q(
        dataout[2]) );
  CFD2QXL \dataout_stg_2_reg[1]  ( .D(n4284), .CP(clk), .CD(n7173), .Q(
        dataout[1]) );
  CFD2QXL \dataout_stg_2_reg[0]  ( .D(n4281), .CP(clk), .CD(n7173), .Q(
        dataout[0]) );
  CFD1XL \buffer_reg[779]  ( .D(n6109), .CP(clk), .Q(n7504), .QN(n3170) );
  CFD1XL \buffer_reg[523]  ( .D(n6103), .CP(clk), .Q(n7760), .QN(n3171) );
  CFD1XL \buffer_reg[267]  ( .D(n6101), .CP(clk), .Q(n8016), .QN(n3172) );
  CFD1XL \buffer_reg[1035]  ( .D(n6097), .CP(clk), .QN(n3169) );
  CFD1XL \buffer_reg[1013]  ( .D(n6095), .CP(clk), .QN(n7262) );
  CFD1XL \buffer_reg[1012]  ( .D(n6087), .CP(clk), .QN(n7264) );
  CFD1XL \buffer_reg[1011]  ( .D(n6085), .CP(clk), .QN(n7266) );
  CFD1XL \buffer_reg[1010]  ( .D(n6079), .CP(clk), .QN(n7267) );
  CFD1XL \buffer_reg[949]  ( .D(n6075), .CP(clk), .QN(n7334) );
  CFD1XL \buffer_reg[948]  ( .D(n6073), .CP(clk), .QN(n7335) );
  CFD1XL \buffer_reg[947]  ( .D(n6071), .CP(clk), .QN(n7336) );
  CFD1XL \buffer_reg[946]  ( .D(n6069), .CP(clk), .QN(n7337) );
  CFD1XL \buffer_reg[885]  ( .D(n6067), .CP(clk), .QN(n7398) );
  CFD1XL \buffer_reg[884]  ( .D(n6065), .CP(clk), .QN(n7399) );
  CFD1XL \buffer_reg[883]  ( .D(n6063), .CP(clk), .QN(n7400) );
  CFD1XL \buffer_reg[882]  ( .D(n6061), .CP(clk), .QN(n7401) );
  CFD1XL \buffer_reg[821]  ( .D(n6059), .CP(clk), .QN(n7462) );
  CFD1XL \buffer_reg[820]  ( .D(n6057), .CP(clk), .QN(n7463) );
  CFD1XL \buffer_reg[819]  ( .D(n6055), .CP(clk), .QN(n7464) );
  CFD1XL \buffer_reg[818]  ( .D(n6053), .CP(clk), .QN(n7465) );
  CFD1XL \buffer_reg[981]  ( .D(n6051), .CP(clk), .QN(n7302) );
  CFD1XL \buffer_reg[980]  ( .D(n6049), .CP(clk), .QN(n7303) );
  CFD1XL \buffer_reg[979]  ( .D(n6047), .CP(clk), .QN(n7304) );
  CFD1XL \buffer_reg[978]  ( .D(n6045), .CP(clk), .QN(n7305) );
  CFD1XL \buffer_reg[917]  ( .D(n6043), .CP(clk), .QN(n7366) );
  CFD1XL \buffer_reg[916]  ( .D(n6037), .CP(clk), .QN(n7367) );
  CFD1XL \buffer_reg[915]  ( .D(n6035), .CP(clk), .QN(n7368) );
  CFD1XL \buffer_reg[914]  ( .D(n6033), .CP(clk), .QN(n7369) );
  CFD1XL \buffer_reg[853]  ( .D(n6031), .CP(clk), .QN(n7430) );
  CFD1XL \buffer_reg[852]  ( .D(n6029), .CP(clk), .QN(n7431) );
  CFD1XL \buffer_reg[851]  ( .D(n6027), .CP(clk), .QN(n7432) );
  CFD1XL \buffer_reg[850]  ( .D(n6025), .CP(clk), .QN(n7433) );
  CFD1XL \buffer_reg[789]  ( .D(n6023), .CP(clk), .QN(n7494) );
  CFD1XL \buffer_reg[788]  ( .D(n6021), .CP(clk), .QN(n7495) );
  CFD1XL \buffer_reg[787]  ( .D(n6017), .CP(clk), .QN(n7496) );
  CFD1XL \buffer_reg[786]  ( .D(n6015), .CP(clk), .QN(n7497) );
  CFD1XL \buffer_reg[1009]  ( .D(n6011), .CP(clk), .QN(n7269) );
  CFD1XL \buffer_reg[1008]  ( .D(n6009), .CP(clk), .QN(n7271) );
  CFD1XL \buffer_reg[1005]  ( .D(n6007), .CP(clk), .QN(n7275) );
  CFD1XL \buffer_reg[1004]  ( .D(n6005), .CP(clk), .QN(n7276) );
  CFD1XL \buffer_reg[945]  ( .D(n6003), .CP(clk), .QN(n7338) );
  CFD1XL \buffer_reg[944]  ( .D(n5999), .CP(clk), .QN(n7339) );
  CFD1XL \buffer_reg[941]  ( .D(n5997), .CP(clk), .QN(n7342) );
  CFD1XL \buffer_reg[940]  ( .D(n5995), .CP(clk), .QN(n7343) );
  CFD1XL \buffer_reg[881]  ( .D(n5993), .CP(clk), .QN(n7402) );
  CFD1XL \buffer_reg[880]  ( .D(n5991), .CP(clk), .QN(n7403) );
  CFD1XL \buffer_reg[877]  ( .D(n5989), .CP(clk), .QN(n7406) );
  CFD1XL \buffer_reg[876]  ( .D(n5987), .CP(clk), .QN(n7407) );
  CFD1XL \buffer_reg[817]  ( .D(n5985), .CP(clk), .QN(n7466) );
  CFD1XL \buffer_reg[816]  ( .D(n5983), .CP(clk), .QN(n7467) );
  CFD1XL \buffer_reg[813]  ( .D(n5981), .CP(clk), .QN(n7470) );
  CFD1XL \buffer_reg[812]  ( .D(n5979), .CP(clk), .QN(n7471) );
  CFD1XL \buffer_reg[977]  ( .D(n5952), .CP(clk), .QN(n7306) );
  CFD1XL \buffer_reg[976]  ( .D(n5950), .CP(clk), .QN(n7307) );
  CFD1XL \buffer_reg[973]  ( .D(n5948), .CP(clk), .QN(n7310) );
  CFD1XL \buffer_reg[972]  ( .D(n5946), .CP(clk), .QN(n7311) );
  CFD1XL \buffer_reg[913]  ( .D(n5942), .CP(clk), .QN(n7370) );
  CFD1XL \buffer_reg[912]  ( .D(n5938), .CP(clk), .QN(n7371) );
  CFD1XL \buffer_reg[849]  ( .D(n5936), .CP(clk), .QN(n7434) );
  CFD1XL \buffer_reg[848]  ( .D(n5934), .CP(clk), .QN(n7435) );
  CFD1XL \buffer_reg[845]  ( .D(n5932), .CP(clk), .QN(n7438) );
  CFD1XL \buffer_reg[844]  ( .D(n5930), .CP(clk), .QN(n7439) );
  CFD1XL \buffer_reg[785]  ( .D(n5928), .CP(clk), .QN(n7498) );
  CFD1XL \buffer_reg[784]  ( .D(n5926), .CP(clk), .QN(n7499) );
  CFD1XL \buffer_reg[1023]  ( .D(n5924), .CP(clk), .QN(n7248) );
  CFD1XL \buffer_reg[1022]  ( .D(n5922), .CP(clk), .QN(n7251) );
  CFD1XL \buffer_reg[1021]  ( .D(n5920), .CP(clk), .QN(n7253) );
  CFD1XL \buffer_reg[1020]  ( .D(n5918), .CP(clk), .QN(n7254) );
  CFD1XL \buffer_reg[1019]  ( .D(n5916), .CP(clk), .QN(n7255) );
  CFD1XL \buffer_reg[1018]  ( .D(n5914), .CP(clk), .QN(n7256) );
  CFD1XL \buffer_reg[1017]  ( .D(n5910), .CP(clk), .QN(n7257) );
  CFD1XL \buffer_reg[1016]  ( .D(n5908), .CP(clk), .QN(n7259) );
  CFD1XL \buffer_reg[1015]  ( .D(n5906), .CP(clk), .QN(n7260) );
  CFD1XL \buffer_reg[1014]  ( .D(n5904), .CP(clk), .QN(n7261) );
  CFD1XL \buffer_reg[1007]  ( .D(n5902), .CP(clk), .Q(n2867), .QN(n7272) );
  CFD1XL \buffer_reg[1006]  ( .D(n5900), .CP(clk), .Q(n2404), .QN(n7273) );
  CFD1XL \buffer_reg[1003]  ( .D(n5894), .CP(clk), .QN(n7278) );
  CFD1XL \buffer_reg[1002]  ( .D(n5888), .CP(clk), .QN(n7280) );
  CFD1XL \buffer_reg[1001]  ( .D(n5886), .CP(clk), .QN(n7282) );
  CFD1XL \buffer_reg[1000]  ( .D(n5884), .CP(clk), .QN(n7283) );
  CFD1XL \buffer_reg[999]  ( .D(n5882), .CP(clk), .QN(n7284) );
  CFD1XL \buffer_reg[998]  ( .D(n5878), .CP(clk), .QN(n7285) );
  CFD1XL \buffer_reg[997]  ( .D(n5874), .CP(clk), .QN(n7286) );
  CFD1XL \buffer_reg[996]  ( .D(n5872), .CP(clk), .QN(n7287) );
  CFD1XL \buffer_reg[995]  ( .D(n5870), .CP(clk), .QN(n7288) );
  CFD1XL \buffer_reg[994]  ( .D(n5868), .CP(clk), .QN(n7289) );
  CFD1XL \buffer_reg[993]  ( .D(n5862), .CP(clk), .QN(n7290) );
  CFD1XL \buffer_reg[992]  ( .D(n5858), .CP(clk), .QN(n7291) );
  CFD1XL \buffer_reg[959]  ( .D(n5852), .CP(clk), .QN(n7324) );
  CFD1XL \buffer_reg[958]  ( .D(n5850), .CP(clk), .QN(n7325) );
  CFD1XL \buffer_reg[957]  ( .D(n5846), .CP(clk), .QN(n7326) );
  CFD1XL \buffer_reg[956]  ( .D(n5842), .CP(clk), .QN(n7327) );
  CFD1XL \buffer_reg[955]  ( .D(n5840), .CP(clk), .QN(n7328) );
  CFD1XL \buffer_reg[954]  ( .D(n5838), .CP(clk), .QN(n7329) );
  CFD1XL \buffer_reg[953]  ( .D(n5836), .CP(clk), .QN(n7330) );
  CFD1XL \buffer_reg[952]  ( .D(n5830), .CP(clk), .QN(n7331) );
  CFD1XL \buffer_reg[951]  ( .D(n5826), .CP(clk), .QN(n7332) );
  CFD1XL \buffer_reg[950]  ( .D(n5824), .CP(clk), .QN(n7333) );
  CFD1XL \buffer_reg[943]  ( .D(n5822), .CP(clk), .QN(n7340) );
  CFD1XL \buffer_reg[942]  ( .D(n5820), .CP(clk), .QN(n7341) );
  CFD1XL \buffer_reg[939]  ( .D(n5818), .CP(clk), .QN(n7344) );
  CFD1XL \buffer_reg[938]  ( .D(n5814), .CP(clk), .QN(n7345) );
  CFD1XL \buffer_reg[937]  ( .D(n5810), .CP(clk), .QN(n7346) );
  CFD1XL \buffer_reg[936]  ( .D(n5808), .CP(clk), .QN(n7347) );
  CFD1XL \buffer_reg[935]  ( .D(n5806), .CP(clk), .QN(n7348) );
  CFD1XL \buffer_reg[934]  ( .D(n5804), .CP(clk), .QN(n7349) );
  CFD1XL \buffer_reg[933]  ( .D(n5798), .CP(clk), .QN(n7350) );
  CFD1XL \buffer_reg[932]  ( .D(n5794), .CP(clk), .QN(n7351) );
  CFD1XL \buffer_reg[931]  ( .D(n5788), .CP(clk), .QN(n7352) );
  CFD1XL \buffer_reg[930]  ( .D(n5786), .CP(clk), .QN(n7353) );
  CFD1XL \buffer_reg[929]  ( .D(n5782), .CP(clk), .QN(n7354) );
  CFD1XL \buffer_reg[928]  ( .D(n5780), .CP(clk), .QN(n7355) );
  CFD1XL \buffer_reg[895]  ( .D(n5778), .CP(clk), .QN(n7388) );
  CFD1XL \buffer_reg[894]  ( .D(n5776), .CP(clk), .QN(n7389) );
  CFD1XL \buffer_reg[893]  ( .D(n5774), .CP(clk), .QN(n7390) );
  CFD1XL \buffer_reg[892]  ( .D(n5772), .CP(clk), .QN(n7391) );
  CFD1XL \buffer_reg[891]  ( .D(n5766), .CP(clk), .QN(n7392) );
  CFD1XL \buffer_reg[890]  ( .D(n5762), .CP(clk), .QN(n7393) );
  CFD1XL \buffer_reg[889]  ( .D(n5760), .CP(clk), .QN(n7394) );
  CFD1XL \buffer_reg[888]  ( .D(n5758), .CP(clk), .QN(n7395) );
  CFD1XL \buffer_reg[887]  ( .D(n5756), .CP(clk), .QN(n7396) );
  CFD1XL \buffer_reg[886]  ( .D(n5754), .CP(clk), .QN(n7397) );
  CFD1XL \buffer_reg[879]  ( .D(n5750), .CP(clk), .QN(n7404) );
  CFD1XL \buffer_reg[878]  ( .D(n5746), .CP(clk), .QN(n7405) );
  CFD1XL \buffer_reg[875]  ( .D(n5744), .CP(clk), .QN(n7408) );
  CFD1XL \buffer_reg[874]  ( .D(n5742), .CP(clk), .QN(n7409) );
  CFD1XL \buffer_reg[873]  ( .D(n5740), .CP(clk), .QN(n7410) );
  CFD1XL \buffer_reg[872]  ( .D(n5738), .CP(clk), .QN(n7411) );
  CFD1XL \buffer_reg[871]  ( .D(n5736), .CP(clk), .QN(n7412) );
  CFD1XL \buffer_reg[870]  ( .D(n5734), .CP(clk), .QN(n7413) );
  CFD1XL \buffer_reg[869]  ( .D(n5732), .CP(clk), .QN(n7414) );
  CFD1XL \buffer_reg[868]  ( .D(n5730), .CP(clk), .QN(n7415) );
  CFD1XL \buffer_reg[867]  ( .D(n5696), .CP(clk), .QN(n7416) );
  CFD1XL \buffer_reg[866]  ( .D(n5694), .CP(clk), .QN(n7417) );
  CFD1XL \buffer_reg[865]  ( .D(n5692), .CP(clk), .QN(n7418) );
  CFD1XL \buffer_reg[864]  ( .D(n5690), .CP(clk), .QN(n7419) );
  CFD1XL \buffer_reg[831]  ( .D(n5688), .CP(clk), .QN(n7452) );
  CFD1XL \buffer_reg[830]  ( .D(n5686), .CP(clk), .QN(n7453) );
  CFD1XL \buffer_reg[829]  ( .D(n5684), .CP(clk), .QN(n7454) );
  CFD1XL \buffer_reg[828]  ( .D(n5682), .CP(clk), .QN(n7455) );
  CFD1XL \buffer_reg[827]  ( .D(n5680), .CP(clk), .QN(n7456) );
  CFD1XL \buffer_reg[826]  ( .D(n5678), .CP(clk), .QN(n7457) );
  CFD1XL \buffer_reg[825]  ( .D(n5676), .CP(clk), .QN(n7458) );
  CFD1XL \buffer_reg[824]  ( .D(n5674), .CP(clk), .QN(n7459) );
  CFD1XL \buffer_reg[823]  ( .D(n5672), .CP(clk), .QN(n7460) );
  CFD1XL \buffer_reg[822]  ( .D(n5670), .CP(clk), .QN(n7461) );
  CFD1XL \buffer_reg[815]  ( .D(n5668), .CP(clk), .QN(n7468) );
  CFD1XL \buffer_reg[814]  ( .D(n5666), .CP(clk), .QN(n7469) );
  CFD1XL \buffer_reg[811]  ( .D(n5664), .CP(clk), .QN(n7472) );
  CFD1XL \buffer_reg[810]  ( .D(n5662), .CP(clk), .QN(n7473) );
  CFD1XL \buffer_reg[809]  ( .D(n5660), .CP(clk), .QN(n7474) );
  CFD1XL \buffer_reg[808]  ( .D(n5658), .CP(clk), .QN(n7475) );
  CFD1XL \buffer_reg[807]  ( .D(n5656), .CP(clk), .QN(n7476) );
  CFD1XL \buffer_reg[806]  ( .D(n5654), .CP(clk), .QN(n7477) );
  CFD1XL \buffer_reg[805]  ( .D(n5652), .CP(clk), .QN(n7478) );
  CFD1XL \buffer_reg[804]  ( .D(n5650), .CP(clk), .QN(n7479) );
  CFD1XL \buffer_reg[803]  ( .D(n5648), .CP(clk), .QN(n7480) );
  CFD1XL \buffer_reg[802]  ( .D(n5646), .CP(clk), .QN(n7481) );
  CFD1XL \buffer_reg[801]  ( .D(n5644), .CP(clk), .QN(n7482) );
  CFD1XL \buffer_reg[800]  ( .D(n5640), .CP(clk), .QN(n7483) );
  CFD1XL \buffer_reg[991]  ( .D(n5638), .CP(clk), .QN(n7292) );
  CFD1XL \buffer_reg[990]  ( .D(n5634), .CP(clk), .QN(n7293) );
  CFD1XL \buffer_reg[989]  ( .D(n5632), .CP(clk), .QN(n7294) );
  CFD1XL \buffer_reg[988]  ( .D(n5630), .CP(clk), .QN(n7295) );
  CFD1XL \buffer_reg[987]  ( .D(n5628), .CP(clk), .QN(n7296) );
  CFD1XL \buffer_reg[986]  ( .D(n5626), .CP(clk), .QN(n7297) );
  CFD1XL \buffer_reg[985]  ( .D(n5622), .CP(clk), .QN(n7298) );
  CFD1XL \buffer_reg[984]  ( .D(n5620), .CP(clk), .QN(n7299) );
  CFD1XL \buffer_reg[983]  ( .D(n5618), .CP(clk), .QN(n7300) );
  CFD1XL \buffer_reg[982]  ( .D(n5616), .CP(clk), .QN(n7301) );
  CFD1XL \buffer_reg[975]  ( .D(n5614), .CP(clk), .QN(n7308) );
  CFD1XL \buffer_reg[974]  ( .D(n5612), .CP(clk), .QN(n7309) );
  CFD1XL \buffer_reg[971]  ( .D(n5610), .CP(clk), .QN(n7312) );
  CFD1XL \buffer_reg[970]  ( .D(n5608), .CP(clk), .QN(n7313) );
  CFD1XL \buffer_reg[969]  ( .D(n5606), .CP(clk), .QN(n7314) );
  CFD1XL \buffer_reg[968]  ( .D(n5604), .CP(clk), .QN(n7315) );
  CFD1XL \buffer_reg[967]  ( .D(n5602), .CP(clk), .QN(n7316) );
  CFD1XL \buffer_reg[966]  ( .D(n5596), .CP(clk), .QN(n7317) );
  CFD1XL \buffer_reg[965]  ( .D(n5594), .CP(clk), .QN(n7318) );
  CFD1XL \buffer_reg[964]  ( .D(n5592), .CP(clk), .QN(n7319) );
  CFD1XL \buffer_reg[963]  ( .D(n5590), .CP(clk), .QN(n7320) );
  CFD1XL \buffer_reg[962]  ( .D(n5586), .CP(clk), .QN(n7321) );
  CFD1XL \buffer_reg[961]  ( .D(n5584), .CP(clk), .QN(n7322) );
  CFD1XL \buffer_reg[960]  ( .D(n5582), .CP(clk), .QN(n7323) );
  CFD1XL \buffer_reg[927]  ( .D(n5580), .CP(clk), .QN(n7356) );
  CFD1XL \buffer_reg[926]  ( .D(n5574), .CP(clk), .QN(n7357) );
  CFD1XL \buffer_reg[925]  ( .D(n5570), .CP(clk), .QN(n7358) );
  CFD1XL \buffer_reg[924]  ( .D(n5568), .CP(clk), .QN(n7359) );
  CFD1XL \buffer_reg[923]  ( .D(n5566), .CP(clk), .QN(n7360) );
  CFD1XL \buffer_reg[922]  ( .D(n5564), .CP(clk), .QN(n7361) );
  CFD1XL \buffer_reg[921]  ( .D(n5562), .CP(clk), .QN(n7362) );
  CFD1XL \buffer_reg[920]  ( .D(n5560), .CP(clk), .QN(n7363) );
  CFD1XL \buffer_reg[919]  ( .D(n5558), .CP(clk), .QN(n7364) );
  CFD1XL \buffer_reg[918]  ( .D(n5556), .CP(clk), .QN(n7365) );
  CFD1XL \buffer_reg[911]  ( .D(n5554), .CP(clk), .Q(n2851), .QN(n7372) );
  CFD1XL \buffer_reg[910]  ( .D(n5552), .CP(clk), .Q(n2388), .QN(n7373) );
  CFD1XL \buffer_reg[863]  ( .D(n5550), .CP(clk), .QN(n7420) );
  CFD1XL \buffer_reg[862]  ( .D(n5548), .CP(clk), .QN(n7421) );
  CFD1XL \buffer_reg[861]  ( .D(n5546), .CP(clk), .QN(n7422) );
  CFD1XL \buffer_reg[860]  ( .D(n5544), .CP(clk), .QN(n7423) );
  CFD1XL \buffer_reg[859]  ( .D(n5542), .CP(clk), .QN(n7424) );
  CFD1XL \buffer_reg[858]  ( .D(n5540), .CP(clk), .QN(n7425) );
  CFD1XL \buffer_reg[857]  ( .D(n5538), .CP(clk), .QN(n7426) );
  CFD1XL \buffer_reg[856]  ( .D(n5532), .CP(clk), .QN(n7427) );
  CFD1XL \buffer_reg[855]  ( .D(n5530), .CP(clk), .QN(n7428) );
  CFD1XL \buffer_reg[854]  ( .D(n5528), .CP(clk), .QN(n7429) );
  CFD1XL \buffer_reg[847]  ( .D(n5526), .CP(clk), .QN(n7436) );
  CFD1XL \buffer_reg[846]  ( .D(n5525), .CP(clk), .QN(n7437) );
  CFD1XL \buffer_reg[843]  ( .D(n5523), .CP(clk), .QN(n7440) );
  CFD1XL \buffer_reg[842]  ( .D(n5521), .CP(clk), .QN(n7441) );
  CFD1XL \buffer_reg[841]  ( .D(n5519), .CP(clk), .QN(n7442) );
  CFD1XL \buffer_reg[840]  ( .D(n5517), .CP(clk), .QN(n7443) );
  CFD1XL \buffer_reg[839]  ( .D(n5513), .CP(clk), .QN(n7444) );
  CFD1XL \buffer_reg[838]  ( .D(n5511), .CP(clk), .QN(n7445) );
  CFD1XL \buffer_reg[837]  ( .D(n5507), .CP(clk), .QN(n7446) );
  CFD1XL \buffer_reg[836]  ( .D(n5505), .CP(clk), .QN(n7447) );
  CFD1XL \buffer_reg[835]  ( .D(n5503), .CP(clk), .QN(n7448) );
  CFD1XL \buffer_reg[834]  ( .D(n5501), .CP(clk), .QN(n7449) );
  CFD1XL \buffer_reg[833]  ( .D(n5499), .CP(clk), .QN(n7450) );
  CFD1XL \buffer_reg[832]  ( .D(n5495), .CP(clk), .QN(n7451) );
  CFD1XL \buffer_reg[799]  ( .D(n5493), .CP(clk), .QN(n7484) );
  CFD1XL \buffer_reg[798]  ( .D(n5491), .CP(clk), .QN(n7485) );
  CFD1XL \buffer_reg[797]  ( .D(n5489), .CP(clk), .QN(n7486) );
  CFD1XL \buffer_reg[796]  ( .D(n5487), .CP(clk), .QN(n7487) );
  CFD1XL \buffer_reg[795]  ( .D(n5485), .CP(clk), .QN(n7488) );
  CFD1XL \buffer_reg[794]  ( .D(n5483), .CP(clk), .QN(n7489) );
  CFD1XL \buffer_reg[793]  ( .D(n5481), .CP(clk), .QN(n7490) );
  CFD1XL \buffer_reg[792]  ( .D(n5479), .CP(clk), .QN(n7491) );
  CFD1XL \buffer_reg[791]  ( .D(n5477), .CP(clk), .QN(n7492) );
  CFD1XL \buffer_reg[790]  ( .D(n5475), .CP(clk), .QN(n7493) );
  CFD1XL \buffer_reg[783]  ( .D(n5473), .CP(clk), .Q(n2847), .QN(n7500) );
  CFD1XL \buffer_reg[782]  ( .D(n5471), .CP(clk), .Q(n2384), .QN(n7501) );
  CFD1XL \buffer_reg[565]  ( .D(n5469), .CP(clk), .QN(n7718) );
  CFD1XL \buffer_reg[564]  ( .D(n5467), .CP(clk), .QN(n7719) );
  CFD1XL \buffer_reg[563]  ( .D(n5463), .CP(clk), .QN(n7720) );
  CFD1XL \buffer_reg[562]  ( .D(n5459), .CP(clk), .QN(n7721) );
  CFD1XL \buffer_reg[533]  ( .D(n5457), .CP(clk), .QN(n7750) );
  CFD1XL \buffer_reg[532]  ( .D(n5455), .CP(clk), .QN(n7751) );
  CFD1XL \buffer_reg[531]  ( .D(n5453), .CP(clk), .QN(n7752) );
  CFD1XL \buffer_reg[530]  ( .D(n5451), .CP(clk), .QN(n7753) );
  CFD1XL \buffer_reg[561]  ( .D(n5449), .CP(clk), .QN(n7722) );
  CFD1XL \buffer_reg[560]  ( .D(n5447), .CP(clk), .QN(n7723) );
  CFD1XL \buffer_reg[557]  ( .D(n5445), .CP(clk), .QN(n7726) );
  CFD1XL \buffer_reg[556]  ( .D(n5443), .CP(clk), .QN(n7727) );
  CFD1XL \buffer_reg[529]  ( .D(n5441), .CP(clk), .QN(n7754) );
  CFD1XL \buffer_reg[528]  ( .D(n5439), .CP(clk), .QN(n7755) );
  CFD1XL \buffer_reg[524]  ( .D(n5438), .CP(clk), .QN(n7759) );
  CFD1XL \buffer_reg[575]  ( .D(n5436), .CP(clk), .QN(n7708) );
  CFD1XL \buffer_reg[574]  ( .D(n5432), .CP(clk), .QN(n7709) );
  CFD1XL \buffer_reg[573]  ( .D(n5430), .CP(clk), .QN(n7710) );
  CFD1XL \buffer_reg[572]  ( .D(n5428), .CP(clk), .QN(n7711) );
  CFD1XL \buffer_reg[571]  ( .D(n5426), .CP(clk), .QN(n7712) );
  CFD1XL \buffer_reg[570]  ( .D(n5424), .CP(clk), .QN(n7713) );
  CFD1XL \buffer_reg[569]  ( .D(n5422), .CP(clk), .QN(n7714) );
  CFD1XL \buffer_reg[568]  ( .D(n5416), .CP(clk), .QN(n7715) );
  CFD1XL \buffer_reg[567]  ( .D(n5410), .CP(clk), .QN(n7716) );
  CFD1XL \buffer_reg[566]  ( .D(n5408), .CP(clk), .QN(n7717) );
  CFD1XL \buffer_reg[559]  ( .D(n5406), .CP(clk), .QN(n7724) );
  CFD1XL \buffer_reg[558]  ( .D(n5404), .CP(clk), .QN(n7725) );
  CFD1XL \buffer_reg[555]  ( .D(n5400), .CP(clk), .QN(n7728) );
  CFD1XL \buffer_reg[554]  ( .D(n5396), .CP(clk), .QN(n7729) );
  CFD1XL \buffer_reg[553]  ( .D(n5394), .CP(clk), .QN(n7730) );
  CFD1XL \buffer_reg[552]  ( .D(n5392), .CP(clk), .QN(n7731) );
  CFD1XL \buffer_reg[551]  ( .D(n5390), .CP(clk), .QN(n7732) );
  CFD1XL \buffer_reg[550]  ( .D(n5384), .CP(clk), .QN(n7733) );
  CFD1XL \buffer_reg[549]  ( .D(n5380), .CP(clk), .QN(n7734) );
  CFD1XL \buffer_reg[548]  ( .D(n5374), .CP(clk), .QN(n7735) );
  CFD1XL \buffer_reg[547]  ( .D(n5372), .CP(clk), .QN(n7736) );
  CFD1XL \buffer_reg[546]  ( .D(n5368), .CP(clk), .QN(n7737) );
  CFD1XL \buffer_reg[545]  ( .D(n5364), .CP(clk), .QN(n7738) );
  CFD1XL \buffer_reg[544]  ( .D(n5362), .CP(clk), .QN(n7739) );
  CFD1XL \buffer_reg[543]  ( .D(n5360), .CP(clk), .QN(n7740) );
  CFD1XL \buffer_reg[542]  ( .D(n5358), .CP(clk), .QN(n7741) );
  CFD1XL \buffer_reg[541]  ( .D(n5352), .CP(clk), .QN(n7742) );
  CFD1XL \buffer_reg[540]  ( .D(n5348), .CP(clk), .QN(n7743) );
  CFD1XL \buffer_reg[539]  ( .D(n5346), .CP(clk), .QN(n7744) );
  CFD1XL \buffer_reg[538]  ( .D(n5344), .CP(clk), .QN(n7745) );
  CFD1XL \buffer_reg[537]  ( .D(n5342), .CP(clk), .QN(n7746) );
  CFD1XL \buffer_reg[536]  ( .D(n5340), .CP(clk), .QN(n7747) );
  CFD1XL \buffer_reg[535]  ( .D(n5336), .CP(clk), .QN(n7748) );
  CFD1XL \buffer_reg[534]  ( .D(n5332), .CP(clk), .QN(n7749) );
  CFD1XL \buffer_reg[527]  ( .D(n5330), .CP(clk), .Q(n2846), .QN(n7756) );
  CFD1XL \buffer_reg[526]  ( .D(n5328), .CP(clk), .Q(n2383), .QN(n7757) );
  CFD1XL \buffer_reg[373]  ( .D(n5326), .CP(clk), .QN(n7910) );
  CFD1XL \buffer_reg[372]  ( .D(n5320), .CP(clk), .QN(n7911) );
  CFD1XL \buffer_reg[371]  ( .D(n5316), .CP(clk), .QN(n7912) );
  CFD1XL \buffer_reg[370]  ( .D(n5310), .CP(clk), .QN(n7913) );
  CFD1XL \buffer_reg[309]  ( .D(n5308), .CP(clk), .QN(n7974) );
  CFD1XL \buffer_reg[308]  ( .D(n5304), .CP(clk), .QN(n7975) );
  CFD1XL \buffer_reg[307]  ( .D(n5302), .CP(clk), .QN(n7976) );
  CFD1XL \buffer_reg[306]  ( .D(n5300), .CP(clk), .QN(n7977) );
  CFD1XL \buffer_reg[369]  ( .D(n5298), .CP(clk), .QN(n7914) );
  CFD1XL \buffer_reg[368]  ( .D(n5296), .CP(clk), .QN(n7915) );
  CFD1XL \buffer_reg[365]  ( .D(n5294), .CP(clk), .QN(n7918) );
  CFD1XL \buffer_reg[364]  ( .D(n5288), .CP(clk), .QN(n7919) );
  CFD1XL \buffer_reg[305]  ( .D(n5284), .CP(clk), .QN(n7978) );
  CFD1XL \buffer_reg[304]  ( .D(n5282), .CP(clk), .QN(n7979) );
  CFD1XL \buffer_reg[301]  ( .D(n5280), .CP(clk), .QN(n7982) );
  CFD1XL \buffer_reg[300]  ( .D(n5278), .CP(clk), .QN(n7983) );
  CFD1XL \buffer_reg[383]  ( .D(n5276), .CP(clk), .QN(n7900) );
  CFD1XL \buffer_reg[382]  ( .D(n5272), .CP(clk), .QN(n7901) );
  CFD1XL \buffer_reg[381]  ( .D(n5268), .CP(clk), .QN(n7902) );
  CFD1XL \buffer_reg[380]  ( .D(n5266), .CP(clk), .QN(n7903) );
  CFD1XL \buffer_reg[379]  ( .D(n5264), .CP(clk), .QN(n7904) );
  CFD1XL \buffer_reg[378]  ( .D(n5262), .CP(clk), .QN(n7905) );
  CFD1XL \buffer_reg[377]  ( .D(n5260), .CP(clk), .QN(n7906) );
  CFD1XL \buffer_reg[376]  ( .D(n5258), .CP(clk), .QN(n7907) );
  CFD1XL \buffer_reg[375]  ( .D(n5256), .CP(clk), .QN(n7908) );
  CFD1XL \buffer_reg[374]  ( .D(n5254), .CP(clk), .QN(n7909) );
  CFD1XL \buffer_reg[367]  ( .D(n5252), .CP(clk), .QN(n7916) );
  CFD1XL \buffer_reg[366]  ( .D(n5244), .CP(clk), .QN(n7917) );
  CFD1XL \buffer_reg[363]  ( .D(n5218), .CP(clk), .QN(n7920) );
  CFD1XL \buffer_reg[362]  ( .D(n5216), .CP(clk), .QN(n7921) );
  CFD1XL \buffer_reg[361]  ( .D(n5214), .CP(clk), .QN(n7922) );
  CFD1XL \buffer_reg[360]  ( .D(n5212), .CP(clk), .QN(n7923) );
  CFD1XL \buffer_reg[359]  ( .D(n5210), .CP(clk), .QN(n7924) );
  CFD1XL \buffer_reg[358]  ( .D(n5208), .CP(clk), .QN(n7925) );
  CFD1XL \buffer_reg[357]  ( .D(n5206), .CP(clk), .QN(n7926) );
  CFD1XL \buffer_reg[356]  ( .D(n5204), .CP(clk), .QN(n7927) );
  CFD1XL \buffer_reg[355]  ( .D(n5202), .CP(clk), .QN(n7928) );
  CFD1XL \buffer_reg[354]  ( .D(n5200), .CP(clk), .QN(n7929) );
  CFD1XL \buffer_reg[353]  ( .D(n5198), .CP(clk), .QN(n7930) );
  CFD1XL \buffer_reg[352]  ( .D(n5196), .CP(clk), .QN(n7931) );
  CFD1XL \buffer_reg[319]  ( .D(n5194), .CP(clk), .QN(n7964) );
  CFD1XL \buffer_reg[318]  ( .D(n5192), .CP(clk), .QN(n7965) );
  CFD1XL \buffer_reg[317]  ( .D(n5190), .CP(clk), .QN(n7966) );
  CFD1XL \buffer_reg[316]  ( .D(n5188), .CP(clk), .QN(n7967) );
  CFD1XL \buffer_reg[315]  ( .D(n5186), .CP(clk), .QN(n7968) );
  CFD1XL \buffer_reg[314]  ( .D(n5184), .CP(clk), .QN(n7969) );
  CFD1XL \buffer_reg[313]  ( .D(n5182), .CP(clk), .QN(n7970) );
  CFD1XL \buffer_reg[312]  ( .D(n5180), .CP(clk), .QN(n7971) );
  CFD1XL \buffer_reg[311]  ( .D(n5178), .CP(clk), .QN(n7972) );
  CFD1XL \buffer_reg[310]  ( .D(n5176), .CP(clk), .QN(n7973) );
  CFD1XL \buffer_reg[303]  ( .D(n5174), .CP(clk), .QN(n7980) );
  CFD1XL \buffer_reg[302]  ( .D(n5172), .CP(clk), .QN(n7981) );
  CFD1XL \buffer_reg[299]  ( .D(n5170), .CP(clk), .QN(n7984) );
  CFD1XL \buffer_reg[298]  ( .D(n5168), .CP(clk), .QN(n7985) );
  CFD1XL \buffer_reg[297]  ( .D(n5166), .CP(clk), .QN(n7986) );
  CFD1XL \buffer_reg[296]  ( .D(n5160), .CP(clk), .QN(n7987) );
  CFD1XL \buffer_reg[295]  ( .D(n5156), .CP(clk), .QN(n7988) );
  CFD1XL \buffer_reg[294]  ( .D(n5154), .CP(clk), .QN(n7989) );
  CFD1XL \buffer_reg[293]  ( .D(n5152), .CP(clk), .QN(n7990) );
  CFD1XL \buffer_reg[292]  ( .D(n5150), .CP(clk), .QN(n7991) );
  CFD1XL \buffer_reg[291]  ( .D(n5148), .CP(clk), .QN(n7992) );
  CFD1XL \buffer_reg[290]  ( .D(n5146), .CP(clk), .QN(n7993) );
  CFD1XL \buffer_reg[289]  ( .D(n5144), .CP(clk), .QN(n7994) );
  CFD1XL \buffer_reg[288]  ( .D(n5142), .CP(clk), .QN(n7995) );
  CFD1XL \buffer_reg[53]  ( .D(n5140), .CP(clk), .QN(n8230) );
  CFD1XL \buffer_reg[52]  ( .D(n5138), .CP(clk), .QN(n8231) );
  CFD1XL \buffer_reg[51]  ( .D(n5136), .CP(clk), .QN(n8232) );
  CFD1XL \buffer_reg[50]  ( .D(n5134), .CP(clk), .QN(n8233) );
  CFD1XL \buffer_reg[49]  ( .D(n5132), .CP(clk), .QN(n8234) );
  CFD1XL \buffer_reg[48]  ( .D(n5130), .CP(clk), .QN(n8235) );
  CFD1XL \buffer_reg[45]  ( .D(n5128), .CP(clk), .QN(n8238) );
  CFD1XL \buffer_reg[44]  ( .D(n5126), .CP(clk), .QN(n8239) );
  CFD1XL \buffer_reg[63]  ( .D(n5124), .CP(clk), .QN(n8220) );
  CFD1XL \buffer_reg[62]  ( .D(n5118), .CP(clk), .QN(n8221) );
  CFD1XL \buffer_reg[61]  ( .D(n5116), .CP(clk), .QN(n8222) );
  CFD1XL \buffer_reg[60]  ( .D(n5114), .CP(clk), .QN(n8223) );
  CFD1XL \buffer_reg[59]  ( .D(n5112), .CP(clk), .QN(n8224) );
  CFD1XL \buffer_reg[58]  ( .D(n5110), .CP(clk), .QN(n8225) );
  CFD1XL \buffer_reg[57]  ( .D(n5108), .CP(clk), .QN(n8226) );
  CFD1XL \buffer_reg[56]  ( .D(n5106), .CP(clk), .QN(n8227) );
  CFD1XL \buffer_reg[55]  ( .D(n5104), .CP(clk), .QN(n8228) );
  CFD1XL \buffer_reg[54]  ( .D(n5102), .CP(clk), .QN(n8229) );
  CFD1XL \buffer_reg[47]  ( .D(n5096), .CP(clk), .QN(n8236) );
  CFD1XL \buffer_reg[46]  ( .D(n5092), .CP(clk), .QN(n8237) );
  CFD1XL \buffer_reg[43]  ( .D(n5090), .CP(clk), .QN(n8240) );
  CFD1XL \buffer_reg[42]  ( .D(n5088), .CP(clk), .QN(n8241) );
  CFD1XL \buffer_reg[41]  ( .D(n5086), .CP(clk), .QN(n8242) );
  CFD1XL \buffer_reg[40]  ( .D(n5084), .CP(clk), .QN(n8243) );
  CFD1XL \buffer_reg[39]  ( .D(n5082), .CP(clk), .QN(n8244) );
  CFD1XL \buffer_reg[38]  ( .D(n5080), .CP(clk), .QN(n8245) );
  CFD1XL \buffer_reg[37]  ( .D(n5078), .CP(clk), .QN(n8246) );
  CFD1XL \buffer_reg[36]  ( .D(n5076), .CP(clk), .QN(n8247) );
  CFD1XL \buffer_reg[35]  ( .D(n5074), .CP(clk), .QN(n8248) );
  CFD1XL \buffer_reg[34]  ( .D(n5072), .CP(clk), .QN(n8249) );
  CFD1XL \buffer_reg[33]  ( .D(n5070), .CP(clk), .QN(n8250) );
  CFD1XL \buffer_reg[32]  ( .D(n5068), .CP(clk), .QN(n8251) );
  CFD1XL \buffer_reg[405]  ( .D(n5066), .CP(clk), .QN(n7878) );
  CFD1XL \buffer_reg[404]  ( .D(n5064), .CP(clk), .QN(n7879) );
  CFD1XL \buffer_reg[403]  ( .D(n5062), .CP(clk), .QN(n7880) );
  CFD1XL \buffer_reg[402]  ( .D(n5060), .CP(clk), .QN(n7881) );
  CFD1XL \buffer_reg[341]  ( .D(n5058), .CP(clk), .QN(n7942) );
  CFD1XL \buffer_reg[340]  ( .D(n5056), .CP(clk), .QN(n7943) );
  CFD1XL \buffer_reg[339]  ( .D(n5054), .CP(clk), .QN(n7944) );
  CFD1XL \buffer_reg[338]  ( .D(n5052), .CP(clk), .QN(n7945) );
  CFD1XL \buffer_reg[277]  ( .D(n5050), .CP(clk), .QN(n8006) );
  CFD1XL \buffer_reg[276]  ( .D(n5048), .CP(clk), .QN(n8007) );
  CFD1XL \buffer_reg[275]  ( .D(n5046), .CP(clk), .QN(n8008) );
  CFD1XL \buffer_reg[274]  ( .D(n5044), .CP(clk), .QN(n8009) );
  CFD1XL \buffer_reg[401]  ( .D(n5042), .CP(clk), .QN(n7882) );
  CFD1XL \buffer_reg[400]  ( .D(n5040), .CP(clk), .QN(n7883) );
  CFD1XL \buffer_reg[337]  ( .D(n5038), .CP(clk), .QN(n7946) );
  CFD1XL \buffer_reg[336]  ( .D(n5032), .CP(clk), .QN(n7947) );
  CFD1XL \buffer_reg[333]  ( .D(n5028), .CP(clk), .QN(n7950) );
  CFD1XL \buffer_reg[332]  ( .D(n5026), .CP(clk), .QN(n7951) );
  CFD1XL \buffer_reg[273]  ( .D(n5024), .CP(clk), .QN(n8010) );
  CFD1XL \buffer_reg[272]  ( .D(n5022), .CP(clk), .QN(n8011) );
  CFD1XL \buffer_reg[268]  ( .D(n5020), .CP(clk), .Q(n3162), .QN(n8015) );
  CFD1XL \buffer_reg[501]  ( .D(n5018), .CP(clk), .QN(n7782) );
  CFD1XL \buffer_reg[500]  ( .D(n5016), .CP(clk), .QN(n7783) );
  CFD1XL \buffer_reg[499]  ( .D(n5014), .CP(clk), .QN(n7784) );
  CFD1XL \buffer_reg[498]  ( .D(n5012), .CP(clk), .QN(n7785) );
  CFD1XL \buffer_reg[437]  ( .D(n5010), .CP(clk), .QN(n7846) );
  CFD1XL \buffer_reg[436]  ( .D(n5008), .CP(clk), .QN(n7847) );
  CFD1XL \buffer_reg[435]  ( .D(n5006), .CP(clk), .QN(n7848) );
  CFD1XL \buffer_reg[434]  ( .D(n5004), .CP(clk), .QN(n7849) );
  CFD1XL \buffer_reg[415]  ( .D(n5002), .CP(clk), .QN(n7868) );
  CFD1XL \buffer_reg[414]  ( .D(n5000), .CP(clk), .QN(n7869) );
  CFD1XL \buffer_reg[413]  ( .D(n4998), .CP(clk), .QN(n7870) );
  CFD1XL \buffer_reg[412]  ( .D(n4996), .CP(clk), .QN(n7871) );
  CFD1XL \buffer_reg[411]  ( .D(n4994), .CP(clk), .QN(n7872) );
  CFD1XL \buffer_reg[410]  ( .D(n4992), .CP(clk), .QN(n7873) );
  CFD1XL \buffer_reg[409]  ( .D(n4962), .CP(clk), .QN(n7874) );
  CFD1XL \buffer_reg[408]  ( .D(n4960), .CP(clk), .QN(n7875) );
  CFD1XL \buffer_reg[407]  ( .D(n4958), .CP(clk), .QN(n7876) );
  CFD1XL \buffer_reg[406]  ( .D(n4956), .CP(clk), .QN(n7877) );
  CFD1XL \buffer_reg[399]  ( .D(n4952), .CP(clk), .QN(n7884) );
  CFD1XL \buffer_reg[398]  ( .D(n4948), .CP(clk), .QN(n7885) );
  CFD1XL \buffer_reg[351]  ( .D(n4946), .CP(clk), .QN(n7932) );
  CFD1XL \buffer_reg[350]  ( .D(n4944), .CP(clk), .QN(n7933) );
  CFD1XL \buffer_reg[349]  ( .D(n4942), .CP(clk), .QN(n7934) );
  CFD1XL \buffer_reg[348]  ( .D(n4940), .CP(clk), .QN(n7935) );
  CFD1XL \buffer_reg[347]  ( .D(n4938), .CP(clk), .QN(n7936) );
  CFD1XL \buffer_reg[346]  ( .D(n4936), .CP(clk), .QN(n7937) );
  CFD1XL \buffer_reg[345]  ( .D(n4932), .CP(clk), .QN(n7938) );
  CFD1XL \buffer_reg[344]  ( .D(n4930), .CP(clk), .QN(n7939) );
  CFD1XL \buffer_reg[343]  ( .D(n4928), .CP(clk), .QN(n7940) );
  CFD1XL \buffer_reg[342]  ( .D(n4926), .CP(clk), .QN(n7941) );
  CFD1XL \buffer_reg[335]  ( .D(n4924), .CP(clk), .QN(n7948) );
  CFD1XL \buffer_reg[334]  ( .D(n4922), .CP(clk), .QN(n7949) );
  CFD1XL \buffer_reg[331]  ( .D(n4920), .CP(clk), .QN(n7952) );
  CFD1XL \buffer_reg[330]  ( .D(n4918), .CP(clk), .QN(n7953) );
  CFD1XL \buffer_reg[329]  ( .D(n4916), .CP(clk), .QN(n7954) );
  CFD1XL \buffer_reg[328]  ( .D(n4914), .CP(clk), .QN(n7955) );
  CFD1XL \buffer_reg[327]  ( .D(n4912), .CP(clk), .QN(n7956) );
  CFD1XL \buffer_reg[326]  ( .D(n4904), .CP(clk), .QN(n7957) );
  CFD1XL \buffer_reg[325]  ( .D(n4898), .CP(clk), .QN(n7958) );
  CFD1XL \buffer_reg[324]  ( .D(n4896), .CP(clk), .QN(n7959) );
  CFD1XL \buffer_reg[323]  ( .D(n4894), .CP(clk), .QN(n7960) );
  CFD1XL \buffer_reg[322]  ( .D(n4888), .CP(clk), .QN(n7961) );
  CFD1XL \buffer_reg[321]  ( .D(n4884), .CP(clk), .QN(n7962) );
  CFD1XL \buffer_reg[320]  ( .D(n4882), .CP(clk), .QN(n7963) );
  CFD1XL \buffer_reg[287]  ( .D(n4880), .CP(clk), .QN(n7996) );
  CFD1XL \buffer_reg[286]  ( .D(n4878), .CP(clk), .QN(n7997) );
  CFD1XL \buffer_reg[285]  ( .D(n4872), .CP(clk), .QN(n7998) );
  CFD1XL \buffer_reg[284]  ( .D(n4868), .CP(clk), .QN(n7999) );
  CFD1XL \buffer_reg[283]  ( .D(n4862), .CP(clk), .QN(n8000) );
  CFD1XL \buffer_reg[282]  ( .D(n4860), .CP(clk), .QN(n8001) );
  CFD1XL \buffer_reg[281]  ( .D(n4856), .CP(clk), .QN(n8002) );
  CFD1XL \buffer_reg[280]  ( .D(n4852), .CP(clk), .QN(n8003) );
  CFD1XL \buffer_reg[279]  ( .D(n4850), .CP(clk), .QN(n8004) );
  CFD1XL \buffer_reg[278]  ( .D(n4848), .CP(clk), .QN(n8005) );
  CFD1XL \buffer_reg[271]  ( .D(n4846), .CP(clk), .QN(n8012) );
  CFD1XL \buffer_reg[270]  ( .D(n4840), .CP(clk), .QN(n8013) );
  CFD1XL \buffer_reg[497]  ( .D(n4836), .CP(clk), .QN(n7786) );
  CFD1XL \buffer_reg[496]  ( .D(n4834), .CP(clk), .QN(n7787) );
  CFD1XL \buffer_reg[493]  ( .D(n4832), .CP(clk), .QN(n7790) );
  CFD1XL \buffer_reg[492]  ( .D(n4830), .CP(clk), .QN(n7791) );
  CFD1XL \buffer_reg[433]  ( .D(n4828), .CP(clk), .QN(n7850) );
  CFD1XL \buffer_reg[432]  ( .D(n4824), .CP(clk), .QN(n7851) );
  CFD1XL \buffer_reg[429]  ( .D(n4820), .CP(clk), .QN(n7854) );
  CFD1XL \buffer_reg[428]  ( .D(n4818), .CP(clk), .QN(n7855) );
  CFD1XL \buffer_reg[511]  ( .D(n4816), .CP(clk), .QN(n7772) );
  CFD1XL \buffer_reg[510]  ( .D(n4814), .CP(clk), .QN(n7773) );
  CFD1XL \buffer_reg[509]  ( .D(n4808), .CP(clk), .QN(n7774) );
  CFD1XL \buffer_reg[508]  ( .D(n4804), .CP(clk), .QN(n7775) );
  CFD1XL \buffer_reg[507]  ( .D(n4798), .CP(clk), .QN(n7776) );
  CFD1XL \buffer_reg[506]  ( .D(n4796), .CP(clk), .QN(n7777) );
  CFD1XL \buffer_reg[505]  ( .D(n4794), .CP(clk), .QN(n7778) );
  CFD1XL \buffer_reg[504]  ( .D(n4792), .CP(clk), .QN(n7779) );
  CFD1XL \buffer_reg[503]  ( .D(n4790), .CP(clk), .QN(n7780) );
  CFD1XL \buffer_reg[502]  ( .D(n4788), .CP(clk), .QN(n7781) );
  CFD1XL \buffer_reg[495]  ( .D(n4786), .CP(clk), .QN(n7788) );
  CFD1XL \buffer_reg[494]  ( .D(n4784), .CP(clk), .QN(n7789) );
  CFD1XL \buffer_reg[491]  ( .D(n4782), .CP(clk), .QN(n7792) );
  CFD1XL \buffer_reg[490]  ( .D(n4776), .CP(clk), .QN(n7793) );
  CFD1XL \buffer_reg[489]  ( .D(n4770), .CP(clk), .QN(n7794) );
  CFD1XL \buffer_reg[488]  ( .D(n4768), .CP(clk), .QN(n7795) );
  CFD1XL \buffer_reg[487]  ( .D(n4766), .CP(clk), .QN(n7796) );
  CFD1XL \buffer_reg[486]  ( .D(n4764), .CP(clk), .QN(n7797) );
  CFD1XL \buffer_reg[485]  ( .D(n4760), .CP(clk), .QN(n7798) );
  CFD1XL \buffer_reg[484]  ( .D(n4756), .CP(clk), .QN(n7799) );
  CFD1XL \buffer_reg[483]  ( .D(n4754), .CP(clk), .QN(n7800) );
  CFD1XL \buffer_reg[482]  ( .D(n4752), .CP(clk), .QN(n7801) );
  CFD1XL \buffer_reg[481]  ( .D(n4750), .CP(clk), .QN(n7802) );
  CFD1XL \buffer_reg[480]  ( .D(n4748), .CP(clk), .QN(n7803) );
  CFD1XL \buffer_reg[447]  ( .D(n4746), .CP(clk), .QN(n7836) );
  CFD1XL \buffer_reg[446]  ( .D(n4744), .CP(clk), .QN(n7837) );
  CFD1XL \buffer_reg[445]  ( .D(n4740), .CP(clk), .QN(n7838) );
  CFD1XL \buffer_reg[444]  ( .D(n4738), .CP(clk), .QN(n7839) );
  CFD1XL \buffer_reg[443]  ( .D(n4736), .CP(clk), .QN(n7840) );
  CFD1XL \buffer_reg[442]  ( .D(n4706), .CP(clk), .QN(n7841) );
  CFD1XL \buffer_reg[441]  ( .D(n4704), .CP(clk), .QN(n7842) );
  CFD1XL \buffer_reg[440]  ( .D(n4702), .CP(clk), .QN(n7843) );
  CFD1XL \buffer_reg[439]  ( .D(n4700), .CP(clk), .QN(n7844) );
  CFD1XL \buffer_reg[438]  ( .D(n4698), .CP(clk), .QN(n7845) );
  CFD1XL \buffer_reg[431]  ( .D(n4696), .CP(clk), .QN(n7852) );
  CFD1XL \buffer_reg[430]  ( .D(n4694), .CP(clk), .QN(n7853) );
  CFD1XL \buffer_reg[427]  ( .D(n4692), .CP(clk), .QN(n7856) );
  CFD1XL \buffer_reg[426]  ( .D(n4690), .CP(clk), .QN(n7857) );
  CFD1XL \buffer_reg[425]  ( .D(n4688), .CP(clk), .QN(n7858) );
  CFD1XL \buffer_reg[424]  ( .D(n4686), .CP(clk), .QN(n7859) );
  CFD1XL \buffer_reg[423]  ( .D(n4684), .CP(clk), .QN(n7860) );
  CFD1XL \buffer_reg[422]  ( .D(n4682), .CP(clk), .QN(n7861) );
  CFD1XL \buffer_reg[421]  ( .D(n4680), .CP(clk), .QN(n7862) );
  CFD1XL \buffer_reg[420]  ( .D(n4678), .CP(clk), .QN(n7863) );
  CFD1XL \buffer_reg[419]  ( .D(n4676), .CP(clk), .QN(n7864) );
  CFD1XL \buffer_reg[418]  ( .D(n4670), .CP(clk), .QN(n7865) );
  CFD1XL \buffer_reg[417]  ( .D(n4668), .CP(clk), .QN(n7866) );
  CFD1XL \buffer_reg[416]  ( .D(n4666), .CP(clk), .QN(n7867) );
  CFD1XL \buffer_reg[469]  ( .D(n4664), .CP(clk), .QN(n7814) );
  CFD1XL \buffer_reg[468]  ( .D(n4662), .CP(clk), .QN(n7815) );
  CFD1XL \buffer_reg[467]  ( .D(n4660), .CP(clk), .QN(n7816) );
  CFD1XL \buffer_reg[466]  ( .D(n4658), .CP(clk), .QN(n7817) );
  CFD1XL \buffer_reg[465]  ( .D(n4656), .CP(clk), .QN(n7818) );
  CFD1XL \buffer_reg[464]  ( .D(n4654), .CP(clk), .QN(n7819) );
  CFD1XL \buffer_reg[461]  ( .D(n4650), .CP(clk), .QN(n7822) );
  CFD1XL \buffer_reg[460]  ( .D(n4648), .CP(clk), .QN(n7823) );
  CFD1XL \buffer_reg[479]  ( .D(n4646), .CP(clk), .QN(n7804) );
  CFD1XL \buffer_reg[478]  ( .D(n4644), .CP(clk), .QN(n7805) );
  CFD1XL \buffer_reg[477]  ( .D(n4642), .CP(clk), .QN(n7806) );
  CFD1XL \buffer_reg[476]  ( .D(n4640), .CP(clk), .QN(n7807) );
  CFD1XL \buffer_reg[475]  ( .D(n4638), .CP(clk), .QN(n7808) );
  CFD1XL \buffer_reg[474]  ( .D(n4636), .CP(clk), .QN(n7809) );
  CFD1XL \buffer_reg[473]  ( .D(n4634), .CP(clk), .QN(n7810) );
  CFD1XL \buffer_reg[472]  ( .D(n4632), .CP(clk), .QN(n7811) );
  CFD1XL \buffer_reg[471]  ( .D(n4630), .CP(clk), .QN(n7812) );
  CFD1XL \buffer_reg[470]  ( .D(n4628), .CP(clk), .QN(n7813) );
  CFD1XL \buffer_reg[463]  ( .D(n4626), .CP(clk), .QN(n7820) );
  CFD1XL \buffer_reg[462]  ( .D(n4624), .CP(clk), .QN(n7821) );
  CFD1XL \buffer_reg[459]  ( .D(n4622), .CP(clk), .QN(n7824) );
  CFD1XL \buffer_reg[458]  ( .D(n4620), .CP(clk), .QN(n7825) );
  CFD1XL \buffer_reg[457]  ( .D(n4618), .CP(clk), .QN(n7826) );
  CFD1XL \buffer_reg[456]  ( .D(n4616), .CP(clk), .QN(n7827) );
  CFD1XL \buffer_reg[455]  ( .D(n4614), .CP(clk), .QN(n7828) );
  CFD1XL \buffer_reg[454]  ( .D(n4612), .CP(clk), .QN(n7829) );
  CFD1XL \buffer_reg[453]  ( .D(n4610), .CP(clk), .QN(n7830) );
  CFD1XL \buffer_reg[452]  ( .D(n4608), .CP(clk), .QN(n7831) );
  CFD1XL \buffer_reg[451]  ( .D(n4606), .CP(clk), .QN(n7832) );
  CFD1XL \buffer_reg[450]  ( .D(n4604), .CP(clk), .QN(n7833) );
  CFD1XL \buffer_reg[449]  ( .D(n4602), .CP(clk), .QN(n7834) );
  CFD1XL \buffer_reg[448]  ( .D(n4600), .CP(clk), .QN(n7835) );
  CFD1XL \buffer_reg[693]  ( .D(n4598), .CP(clk), .QN(n7590) );
  CFD1XL \buffer_reg[692]  ( .D(n4596), .CP(clk), .QN(n7591) );
  CFD1XL \buffer_reg[691]  ( .D(n4594), .CP(clk), .QN(n7592) );
  CFD1XL \buffer_reg[690]  ( .D(n4592), .CP(clk), .QN(n7593) );
  CFD1XL \buffer_reg[661]  ( .D(n4590), .CP(clk), .QN(n7622) );
  CFD1XL \buffer_reg[660]  ( .D(n4588), .CP(clk), .QN(n7623) );
  CFD1XL \buffer_reg[659]  ( .D(n4586), .CP(clk), .QN(n7624) );
  CFD1XL \buffer_reg[658]  ( .D(n4584), .CP(clk), .QN(n7625) );
  CFD1XL \buffer_reg[689]  ( .D(n4582), .CP(clk), .QN(n7594) );
  CFD1XL \buffer_reg[688]  ( .D(n4580), .CP(clk), .QN(n7595) );
  CFD1XL \buffer_reg[685]  ( .D(n4578), .CP(clk), .QN(n7598) );
  CFD1XL \buffer_reg[684]  ( .D(n4576), .CP(clk), .QN(n7599) );
  CFD1XL \buffer_reg[657]  ( .D(n4574), .CP(clk), .QN(n7626) );
  CFD1XL \buffer_reg[656]  ( .D(n4572), .CP(clk), .QN(n7627) );
  CFD1XL \buffer_reg[757]  ( .D(n4570), .CP(clk), .QN(n7526) );
  CFD1XL \buffer_reg[756]  ( .D(n4568), .CP(clk), .QN(n7527) );
  CFD1XL \buffer_reg[755]  ( .D(n4566), .CP(clk), .QN(n7528) );
  CFD1XL \buffer_reg[754]  ( .D(n4564), .CP(clk), .QN(n7529) );
  CFD1XL \buffer_reg[725]  ( .D(n4562), .CP(clk), .QN(n7558) );
  CFD1XL \buffer_reg[724]  ( .D(n4560), .CP(clk), .QN(n7559) );
  CFD1XL \buffer_reg[723]  ( .D(n4558), .CP(clk), .QN(n7560) );
  CFD1XL \buffer_reg[722]  ( .D(n4556), .CP(clk), .QN(n7561) );
  CFD1XL \buffer_reg[629]  ( .D(n4554), .CP(clk), .QN(n7654) );
  CFD1XL \buffer_reg[628]  ( .D(n4552), .CP(clk), .QN(n7655) );
  CFD1XL \buffer_reg[627]  ( .D(n4550), .CP(clk), .QN(n7656) );
  CFD1XL \buffer_reg[626]  ( .D(n4548), .CP(clk), .QN(n7657) );
  CFD1XL \buffer_reg[597]  ( .D(n4546), .CP(clk), .QN(n7686) );
  CFD1XL \buffer_reg[596]  ( .D(n4544), .CP(clk), .QN(n7687) );
  CFD1XL \buffer_reg[595]  ( .D(n4542), .CP(clk), .QN(n7688) );
  CFD1XL \buffer_reg[594]  ( .D(n4540), .CP(clk), .QN(n7689) );
  CFD1XL \buffer_reg[753]  ( .D(n4538), .CP(clk), .QN(n7530) );
  CFD1XL \buffer_reg[752]  ( .D(n4536), .CP(clk), .QN(n7531) );
  CFD1XL \buffer_reg[749]  ( .D(n4534), .CP(clk), .QN(n7534) );
  CFD1XL \buffer_reg[748]  ( .D(n4532), .CP(clk), .QN(n7535) );
  CFD1XL \buffer_reg[721]  ( .D(n4530), .CP(clk), .QN(n7562) );
  CFD1XL \buffer_reg[720]  ( .D(n4528), .CP(clk), .QN(n7563) );
  CFD1XL \buffer_reg[717]  ( .D(n4526), .CP(clk), .QN(n7566) );
  CFD1XL \buffer_reg[716]  ( .D(n4524), .CP(clk), .QN(n7567) );
  CFD1XL \buffer_reg[625]  ( .D(n4522), .CP(clk), .QN(n7658) );
  CFD1XL \buffer_reg[624]  ( .D(n4520), .CP(clk), .QN(n7659) );
  CFD1XL \buffer_reg[621]  ( .D(n4518), .CP(clk), .QN(n7662) );
  CFD1XL \buffer_reg[620]  ( .D(n4516), .CP(clk), .QN(n7663) );
  CFD1XL \buffer_reg[593]  ( .D(n4514), .CP(clk), .QN(n7690) );
  CFD1XL \buffer_reg[592]  ( .D(n4512), .CP(clk), .QN(n7691) );
  CFD1XL \buffer_reg[589]  ( .D(n4510), .CP(clk), .QN(n7694) );
  CFD1XL \buffer_reg[588]  ( .D(n4508), .CP(clk), .QN(n7695) );
  CFD1XL \buffer_reg[703]  ( .D(n4506), .CP(clk), .QN(n7580) );
  CFD1XL \buffer_reg[702]  ( .D(n4504), .CP(clk), .QN(n7581) );
  CFD1XL \buffer_reg[701]  ( .D(n4476), .CP(clk), .QN(n7582) );
  CFD1XL \buffer_reg[700]  ( .D(n4474), .CP(clk), .QN(n7583) );
  CFD1XL \buffer_reg[699]  ( .D(n4472), .CP(clk), .QN(n7584) );
  CFD1XL \buffer_reg[698]  ( .D(n4470), .CP(clk), .QN(n7585) );
  CFD1XL \buffer_reg[697]  ( .D(n4468), .CP(clk), .QN(n7586) );
  CFD1XL \buffer_reg[696]  ( .D(n4466), .CP(clk), .QN(n7587) );
  CFD1XL \buffer_reg[695]  ( .D(n4464), .CP(clk), .QN(n7588) );
  CFD1XL \buffer_reg[694]  ( .D(n4462), .CP(clk), .QN(n7589) );
  CFD1XL \buffer_reg[687]  ( .D(n4460), .CP(clk), .QN(n7596) );
  CFD1XL \buffer_reg[686]  ( .D(n4458), .CP(clk), .QN(n7597) );
  CFD1XL \buffer_reg[683]  ( .D(n4456), .CP(clk), .QN(n7600) );
  CFD1XL \buffer_reg[682]  ( .D(n4454), .CP(clk), .QN(n7601) );
  CFD1XL \buffer_reg[681]  ( .D(n4452), .CP(clk), .QN(n7602) );
  CFD1XL \buffer_reg[680]  ( .D(n4450), .CP(clk), .QN(n7603) );
  CFD1XL \buffer_reg[679]  ( .D(n4448), .CP(clk), .QN(n7604) );
  CFD1XL \buffer_reg[678]  ( .D(n4446), .CP(clk), .QN(n7605) );
  CFD1XL \buffer_reg[677]  ( .D(n4444), .CP(clk), .QN(n7606) );
  CFD1XL \buffer_reg[676]  ( .D(n4442), .CP(clk), .QN(n7607) );
  CFD1XL \buffer_reg[675]  ( .D(n4440), .CP(clk), .QN(n7608) );
  CFD1XL \buffer_reg[674]  ( .D(n4438), .CP(clk), .QN(n7609) );
  CFD1XL \buffer_reg[673]  ( .D(n4436), .CP(clk), .QN(n7610) );
  CFD1XL \buffer_reg[672]  ( .D(n4434), .CP(clk), .QN(n7611) );
  CFD1XL \buffer_reg[671]  ( .D(n4432), .CP(clk), .QN(n7612) );
  CFD1XL \buffer_reg[670]  ( .D(n4430), .CP(clk), .QN(n7613) );
  CFD1XL \buffer_reg[669]  ( .D(n4428), .CP(clk), .QN(n7614) );
  CFD1XL \buffer_reg[668]  ( .D(n4426), .CP(clk), .QN(n7615) );
  CFD1XL \buffer_reg[667]  ( .D(n4424), .CP(clk), .QN(n7616) );
  CFD1XL \buffer_reg[666]  ( .D(n4422), .CP(clk), .QN(n7617) );
  CFD1XL \buffer_reg[665]  ( .D(n4420), .CP(clk), .QN(n7618) );
  CFD1XL \buffer_reg[664]  ( .D(n4418), .CP(clk), .QN(n7619) );
  CFD1XL \buffer_reg[663]  ( .D(n4416), .CP(clk), .QN(n7620) );
  CFD1XL \buffer_reg[662]  ( .D(n4414), .CP(clk), .QN(n7621) );
  CFD1XL \buffer_reg[655]  ( .D(n4412), .CP(clk), .Q(n2850), .QN(n7628) );
  CFD1XL \buffer_reg[654]  ( .D(n4410), .CP(clk), .Q(n2387), .QN(n7629) );
  CFD1XL \buffer_reg[767]  ( .D(n4408), .CP(clk), .QN(n7516) );
  CFD1XL \buffer_reg[766]  ( .D(n4406), .CP(clk), .QN(n7517) );
  CFD1XL \buffer_reg[765]  ( .D(n4404), .CP(clk), .QN(n7518) );
  CFD1XL \buffer_reg[764]  ( .D(n4402), .CP(clk), .QN(n7519) );
  CFD1XL \buffer_reg[763]  ( .D(n4400), .CP(clk), .QN(n7520) );
  CFD1XL \buffer_reg[762]  ( .D(n4398), .CP(clk), .QN(n7521) );
  CFD1XL \buffer_reg[761]  ( .D(n4396), .CP(clk), .QN(n7522) );
  CFD1XL \buffer_reg[760]  ( .D(n4394), .CP(clk), .QN(n7523) );
  CFD1XL \buffer_reg[759]  ( .D(n4392), .CP(clk), .QN(n7524) );
  CFD1XL \buffer_reg[758]  ( .D(n4390), .CP(clk), .QN(n7525) );
  CFD1XL \buffer_reg[751]  ( .D(n4388), .CP(clk), .QN(n7532) );
  CFD1XL \buffer_reg[750]  ( .D(n4386), .CP(clk), .QN(n7533) );
  CFD1XL \buffer_reg[747]  ( .D(n4384), .CP(clk), .QN(n7536) );
  CFD1XL \buffer_reg[746]  ( .D(n4382), .CP(clk), .QN(n7537) );
  CFD1XL \buffer_reg[745]  ( .D(n4380), .CP(clk), .QN(n7538) );
  CFD1XL \buffer_reg[744]  ( .D(n4378), .CP(clk), .QN(n7539) );
  CFD1XL \buffer_reg[743]  ( .D(n4376), .CP(clk), .QN(n7540) );
  CFD1XL \buffer_reg[742]  ( .D(n4374), .CP(clk), .QN(n7541) );
  CFD1XL \buffer_reg[741]  ( .D(n4372), .CP(clk), .QN(n7542) );
  CFD1XL \buffer_reg[740]  ( .D(n4370), .CP(clk), .QN(n7543) );
  CFD1XL \buffer_reg[739]  ( .D(n4368), .CP(clk), .QN(n7544) );
  CFD1XL \buffer_reg[738]  ( .D(n4366), .CP(clk), .QN(n7545) );
  CFD1XL \buffer_reg[737]  ( .D(n4364), .CP(clk), .QN(n7546) );
  CFD1XL \buffer_reg[736]  ( .D(n4362), .CP(clk), .QN(n7547) );
  CFD1XL \buffer_reg[735]  ( .D(n4360), .CP(clk), .QN(n7548) );
  CFD1XL \buffer_reg[734]  ( .D(n4358), .CP(clk), .QN(n7549) );
  CFD1XL \buffer_reg[733]  ( .D(n4356), .CP(clk), .QN(n7550) );
  CFD1XL \buffer_reg[732]  ( .D(n4354), .CP(clk), .QN(n7551) );
  CFD1XL \buffer_reg[731]  ( .D(n4352), .CP(clk), .QN(n7552) );
  CFD1XL \buffer_reg[730]  ( .D(n4350), .CP(clk), .QN(n7553) );
  CFD1XL \buffer_reg[729]  ( .D(n4348), .CP(clk), .QN(n7554) );
  CFD1XL \buffer_reg[728]  ( .D(n4346), .CP(clk), .QN(n7555) );
  CFD1XL \buffer_reg[727]  ( .D(n4344), .CP(clk), .QN(n7556) );
  CFD1XL \buffer_reg[726]  ( .D(n4342), .CP(clk), .QN(n7557) );
  CFD1XL \buffer_reg[719]  ( .D(n4340), .CP(clk), .QN(n7564) );
  CFD1XL \buffer_reg[718]  ( .D(n4338), .CP(clk), .QN(n7565) );
  CFD1XL \buffer_reg[715]  ( .D(n4336), .CP(clk), .QN(n7568) );
  CFD1XL \buffer_reg[714]  ( .D(n4334), .CP(clk), .QN(n7569) );
  CFD1XL \buffer_reg[713]  ( .D(n4332), .CP(clk), .QN(n7570) );
  CFD1XL \buffer_reg[712]  ( .D(n4330), .CP(clk), .QN(n7571) );
  CFD1XL \buffer_reg[711]  ( .D(n4328), .CP(clk), .QN(n7572) );
  CFD1XL \buffer_reg[710]  ( .D(n4326), .CP(clk), .QN(n7573) );
  CFD1XL \buffer_reg[709]  ( .D(n4318), .CP(clk), .QN(n7574) );
  CFD1XL \buffer_reg[708]  ( .D(n4990), .CP(clk), .QN(n7575) );
  CFD1XL \buffer_reg[707]  ( .D(n4986), .CP(clk), .QN(n7576) );
  CFD1XL \buffer_reg[706]  ( .D(n4984), .CP(clk), .QN(n7577) );
  CFD1XL \buffer_reg[705]  ( .D(n4980), .CP(clk), .QN(n7578) );
  CFD1XL \buffer_reg[704]  ( .D(n4978), .CP(clk), .QN(n7579) );
  CFD1XL \buffer_reg[639]  ( .D(n4976), .CP(clk), .QN(n7644) );
  CFD1XL \buffer_reg[638]  ( .D(n4974), .CP(clk), .QN(n7645) );
  CFD1XL \buffer_reg[637]  ( .D(n4972), .CP(clk), .QN(n7646) );
  CFD1XL \buffer_reg[636]  ( .D(n4970), .CP(clk), .QN(n7647) );
  CFD1XL \buffer_reg[635]  ( .D(n4968), .CP(clk), .QN(n7648) );
  CFD1XL \buffer_reg[634]  ( .D(n4966), .CP(clk), .QN(n7649) );
  CFD1XL \buffer_reg[633]  ( .D(n4964), .CP(clk), .QN(n7650) );
  CFD1XL \buffer_reg[632]  ( .D(n4498), .CP(clk), .QN(n7651) );
  CFD1XL \buffer_reg[631]  ( .D(n4496), .CP(clk), .QN(n7652) );
  CFD1XL \buffer_reg[630]  ( .D(n4494), .CP(clk), .QN(n7653) );
  CFD1XL \buffer_reg[623]  ( .D(n4492), .CP(clk), .QN(n7660) );
  CFD1XL \buffer_reg[622]  ( .D(n4490), .CP(clk), .QN(n7661) );
  CFD1XL \buffer_reg[619]  ( .D(n4488), .CP(clk), .QN(n7664) );
  CFD1XL \buffer_reg[618]  ( .D(n4486), .CP(clk), .QN(n7665) );
  CFD1XL \buffer_reg[617]  ( .D(n4484), .CP(clk), .QN(n7666) );
  CFD1XL \buffer_reg[616]  ( .D(n4482), .CP(clk), .QN(n7667) );
  CFD1XL \buffer_reg[615]  ( .D(n4480), .CP(clk), .QN(n7668) );
  CFD1XL \buffer_reg[614]  ( .D(n4478), .CP(clk), .QN(n7669) );
  CFD1XL \buffer_reg[613]  ( .D(n6117), .CP(clk), .QN(n7670) );
  CFD1XL \buffer_reg[612]  ( .D(n4982), .CP(clk), .QN(n7671) );
  CFD1XL \buffer_reg[611]  ( .D(n4500), .CP(clk), .QN(n7672) );
  CFD1XL \buffer_reg[610]  ( .D(n4988), .CP(clk), .QN(n7673) );
  CFD1XL \buffer_reg[609]  ( .D(n4312), .CP(clk), .QN(n7674) );
  CFD1XL \buffer_reg[608]  ( .D(n4310), .CP(clk), .QN(n7675) );
  CFD1XL \buffer_reg[607]  ( .D(n5977), .CP(clk), .QN(n7676) );
  CFD1XL \buffer_reg[606]  ( .D(n5975), .CP(clk), .QN(n7677) );
  CFD1XL \buffer_reg[605]  ( .D(n5973), .CP(clk), .QN(n7678) );
  CFD1XL \buffer_reg[604]  ( .D(n5971), .CP(clk), .QN(n7679) );
  CFD1XL \buffer_reg[603]  ( .D(n5969), .CP(clk), .QN(n7680) );
  CFD1XL \buffer_reg[602]  ( .D(n5967), .CP(clk), .QN(n7681) );
  CFD1XL \buffer_reg[601]  ( .D(n5965), .CP(clk), .QN(n7682) );
  CFD1XL \buffer_reg[600]  ( .D(n5963), .CP(clk), .QN(n7683) );
  CFD1XL \buffer_reg[599]  ( .D(n5961), .CP(clk), .QN(n7684) );
  CFD1XL \buffer_reg[598]  ( .D(n5959), .CP(clk), .QN(n7685) );
  CFD1XL \buffer_reg[591]  ( .D(n5957), .CP(clk), .QN(n7692) );
  CFD1XL \buffer_reg[590]  ( .D(n5956), .CP(clk), .QN(n7693) );
  CFD1XL \buffer_reg[587]  ( .D(n5954), .CP(clk), .QN(n7696) );
  CFD1XL \buffer_reg[586]  ( .D(n6135), .CP(clk), .QN(n7697) );
  CFD1XL \buffer_reg[585]  ( .D(n6133), .CP(clk), .QN(n7698) );
  CFD1XL \buffer_reg[584]  ( .D(n6131), .CP(clk), .QN(n7699) );
  CFD1XL \buffer_reg[583]  ( .D(n6129), .CP(clk), .QN(n7700) );
  CFD1XL \buffer_reg[582]  ( .D(n6127), .CP(clk), .QN(n7701) );
  CFD1XL \buffer_reg[581]  ( .D(n6125), .CP(clk), .QN(n7702) );
  CFD1XL \buffer_reg[580]  ( .D(n6123), .CP(clk), .QN(n7703) );
  CFD1XL \buffer_reg[579]  ( .D(n6121), .CP(clk), .QN(n7704) );
  CFD1XL \buffer_reg[578]  ( .D(n6119), .CP(clk), .QN(n7705) );
  CFD1XL \buffer_reg[577]  ( .D(n6115), .CP(clk), .QN(n7706) );
  CFD1XL \buffer_reg[576]  ( .D(n4502), .CP(clk), .QN(n7707) );
  CFD1XL \buffer_reg[181]  ( .D(n5728), .CP(clk), .QN(n8102) );
  CFD1XL \buffer_reg[180]  ( .D(n5726), .CP(clk), .QN(n8103) );
  CFD1XL \buffer_reg[179]  ( .D(n4674), .CP(clk), .QN(n8104) );
  CFD1XL \buffer_reg[178]  ( .D(n4672), .CP(clk), .QN(n8105) );
  CFD1XL \buffer_reg[149]  ( .D(n5722), .CP(clk), .QN(n8134) );
  CFD1XL \buffer_reg[148]  ( .D(n6113), .CP(clk), .QN(n8135) );
  CFD1XL \buffer_reg[147]  ( .D(n6111), .CP(clk), .QN(n8136) );
  CFD1XL \buffer_reg[146]  ( .D(n5250), .CP(clk), .QN(n8137) );
  CFD1XL \buffer_reg[177]  ( .D(n5248), .CP(clk), .QN(n8106) );
  CFD1XL \buffer_reg[176]  ( .D(n4324), .CP(clk), .QN(n8107) );
  CFD1XL \buffer_reg[173]  ( .D(n4322), .CP(clk), .QN(n8110) );
  CFD1XL \buffer_reg[172]  ( .D(n4320), .CP(clk), .QN(n8111) );
  CFD1XL \buffer_reg[145]  ( .D(n4316), .CP(clk), .QN(n8138) );
  CFD1XL \buffer_reg[144]  ( .D(n4314), .CP(clk), .QN(n8139) );
  CFD1XL \buffer_reg[245]  ( .D(n4308), .CP(clk), .QN(n8038) );
  CFD1XL \buffer_reg[244]  ( .D(n4306), .CP(clk), .QN(n8039) );
  CFD1XL \buffer_reg[243]  ( .D(n4304), .CP(clk), .QN(n8040) );
  CFD1XL \buffer_reg[242]  ( .D(n4302), .CP(clk), .QN(n8041) );
  CFD1XL \buffer_reg[213]  ( .D(n4300), .CP(clk), .QN(n8070) );
  CFD1XL \buffer_reg[212]  ( .D(n4298), .CP(clk), .QN(n8071) );
  CFD1XL \buffer_reg[211]  ( .D(n4296), .CP(clk), .QN(n8072) );
  CFD1XL \buffer_reg[210]  ( .D(n4294), .CP(clk), .QN(n8073) );
  CFD1XL \buffer_reg[117]  ( .D(n5700), .CP(clk), .QN(n8166) );
  CFD1XL \buffer_reg[116]  ( .D(n5242), .CP(clk), .QN(n8167) );
  CFD1XL \buffer_reg[115]  ( .D(n4730), .CP(clk), .QN(n8168) );
  CFD1XL \buffer_reg[114]  ( .D(n6137), .CP(clk), .QN(n8169) );
  CFD1XL \buffer_reg[85]  ( .D(n4732), .CP(clk), .QN(n8198) );
  CFD1XL \buffer_reg[84]  ( .D(n5240), .CP(clk), .QN(n8199) );
  CFD1XL \buffer_reg[83]  ( .D(n5236), .CP(clk), .QN(n8200) );
  CFD1XL \buffer_reg[82]  ( .D(n5232), .CP(clk), .QN(n8201) );
  CFD1XL \buffer_reg[241]  ( .D(n5228), .CP(clk), .QN(n8042) );
  CFD1XL \buffer_reg[240]  ( .D(n5224), .CP(clk), .QN(n8043) );
  CFD1XL \buffer_reg[237]  ( .D(n5220), .CP(clk), .QN(n8046) );
  CFD1XL \buffer_reg[236]  ( .D(n5246), .CP(clk), .QN(n8047) );
  CFD1XL \buffer_reg[209]  ( .D(n5238), .CP(clk), .QN(n8074) );
  CFD1XL \buffer_reg[208]  ( .D(n5234), .CP(clk), .QN(n8075) );
  CFD1XL \buffer_reg[205]  ( .D(n5230), .CP(clk), .QN(n8078) );
  CFD1XL \buffer_reg[204]  ( .D(n5226), .CP(clk), .QN(n8079) );
  CFD1XL \buffer_reg[113]  ( .D(n5222), .CP(clk), .QN(n8170) );
  CFD1XL \buffer_reg[112]  ( .D(n4728), .CP(clk), .QN(n8171) );
  CFD1XL \buffer_reg[109]  ( .D(n4724), .CP(clk), .QN(n8174) );
  CFD1XL \buffer_reg[108]  ( .D(n4720), .CP(clk), .QN(n8175) );
  CFD1XL \buffer_reg[81]  ( .D(n4716), .CP(clk), .QN(n8202) );
  CFD1XL \buffer_reg[80]  ( .D(n4712), .CP(clk), .QN(n8203) );
  CFD1XL \buffer_reg[77]  ( .D(n4708), .CP(clk), .QN(n8206) );
  CFD1XL \buffer_reg[76]  ( .D(n4734), .CP(clk), .QN(n8207) );
  CFD1XL \buffer_reg[6]  ( .D(n4726), .CP(clk), .Q(n2453), .QN(n8277) );
  CFD1XL \buffer_reg[5]  ( .D(n4722), .CP(clk), .Q(n3030), .QN(n8278) );
  CFD1XL \buffer_reg[4]  ( .D(n4718), .CP(clk), .Q(n2624), .QN(n8279) );
  CFD1XL \buffer_reg[3]  ( .D(n4714), .CP(clk), .Q(n2755), .QN(n8280) );
  CFD1XL \buffer_reg[2]  ( .D(n4710), .CP(clk), .Q(n2567), .QN(n8281) );
  CFD1XL \buffer_reg[1]  ( .D(n5724), .CP(clk), .Q(n3136), .QN(n8282) );
  CFD1XL \buffer_reg[0]  ( .D(n5716), .CP(clk), .Q(n2235), .QN(n8283) );
  CFD1XL \buffer_reg[191]  ( .D(n5712), .CP(clk), .QN(n8092) );
  CFD1XL \buffer_reg[190]  ( .D(n5708), .CP(clk), .QN(n8093) );
  CFD1XL \buffer_reg[189]  ( .D(n5704), .CP(clk), .QN(n8094) );
  CFD1XL \buffer_reg[188]  ( .D(n5718), .CP(clk), .QN(n8095) );
  CFD1XL \buffer_reg[187]  ( .D(n5714), .CP(clk), .QN(n8096) );
  CFD1XL \buffer_reg[186]  ( .D(n5710), .CP(clk), .QN(n8097) );
  CFD1XL \buffer_reg[185]  ( .D(n5706), .CP(clk), .QN(n8098) );
  CFD1XL \buffer_reg[184]  ( .D(n5702), .CP(clk), .QN(n8099) );
  CFD1XL \buffer_reg[183]  ( .D(n5698), .CP(clk), .QN(n8100) );
  CFD1XL \buffer_reg[182]  ( .D(n5720), .CP(clk), .QN(n8101) );
  CFD1XL \buffer_reg[175]  ( .D(n4276), .CP(clk), .QN(n8108) );
  CFD1XL \buffer_reg[174]  ( .D(n4274), .CP(clk), .QN(n8109) );
  CFD1XL \buffer_reg[171]  ( .D(n6147), .CP(clk), .QN(n8112) );
  CFD1XL \buffer_reg[170]  ( .D(n4272), .CP(clk), .QN(n8113) );
  CFD1XL \buffer_reg[169]  ( .D(n4270), .CP(clk), .QN(n8114) );
  CFD1XL \buffer_reg[168]  ( .D(n6139), .CP(clk), .QN(n8115) );
  CFD1XL \buffer_reg[167]  ( .D(n6143), .CP(clk), .QN(n8116) );
  CFD1XL \buffer_reg[166]  ( .D(n6145), .CP(clk), .QN(n8117) );
  CFD1XL \buffer_reg[165]  ( .D(n4278), .CP(clk), .QN(n8118) );
  CFD1XL \buffer_reg[164]  ( .D(n6107), .CP(clk), .QN(n8119) );
  CFD1XL \buffer_reg[163]  ( .D(n6105), .CP(clk), .QN(n8120) );
  CFD1XL \buffer_reg[162]  ( .D(n6099), .CP(clk), .QN(n8121) );
  CFD1XL \buffer_reg[161]  ( .D(n6093), .CP(clk), .QN(n8122) );
  CFD1XL \buffer_reg[160]  ( .D(n6091), .CP(clk), .QN(n8123) );
  CFD1XL \buffer_reg[159]  ( .D(n6089), .CP(clk), .QN(n8124) );
  CFD1XL \buffer_reg[158]  ( .D(n6083), .CP(clk), .QN(n8125) );
  CFD1XL \buffer_reg[157]  ( .D(n6081), .CP(clk), .QN(n8126) );
  CFD1XL \buffer_reg[156]  ( .D(n6077), .CP(clk), .QN(n8127) );
  CFD1XL \buffer_reg[155]  ( .D(n6041), .CP(clk), .QN(n8128) );
  CFD1XL \buffer_reg[154]  ( .D(n6039), .CP(clk), .QN(n8129) );
  CFD1XL \buffer_reg[153]  ( .D(n6019), .CP(clk), .QN(n8130) );
  CFD1XL \buffer_reg[152]  ( .D(n6013), .CP(clk), .QN(n8131) );
  CFD1XL \buffer_reg[151]  ( .D(n6001), .CP(clk), .QN(n8132) );
  CFD1XL \buffer_reg[150]  ( .D(n5944), .CP(clk), .QN(n8133) );
  CFD1XL \buffer_reg[143]  ( .D(n5940), .CP(clk), .Q(n2848), .QN(n8140) );
  CFD1XL \buffer_reg[142]  ( .D(n5912), .CP(clk), .Q(n2385), .QN(n8141) );
  CFD1XL \buffer_reg[255]  ( .D(n5898), .CP(clk), .QN(n8028) );
  CFD1XL \buffer_reg[254]  ( .D(n5896), .CP(clk), .QN(n8029) );
  CFD1XL \buffer_reg[253]  ( .D(n5892), .CP(clk), .QN(n8030) );
  CFD1XL \buffer_reg[252]  ( .D(n5890), .CP(clk), .QN(n8031) );
  CFD1XL \buffer_reg[251]  ( .D(n5880), .CP(clk), .QN(n8032) );
  CFD1XL \buffer_reg[250]  ( .D(n5876), .CP(clk), .QN(n8033) );
  CFD1XL \buffer_reg[249]  ( .D(n5866), .CP(clk), .QN(n8034) );
  CFD1XL \buffer_reg[248]  ( .D(n5864), .CP(clk), .QN(n8035) );
  CFD1XL \buffer_reg[247]  ( .D(n5860), .CP(clk), .QN(n8036) );
  CFD1XL \buffer_reg[246]  ( .D(n5856), .CP(clk), .QN(n8037) );
  CFD1XL \buffer_reg[239]  ( .D(n5854), .CP(clk), .Q(n2864), .QN(n8044) );
  CFD1XL \buffer_reg[238]  ( .D(n5848), .CP(clk), .Q(n2401), .QN(n8045) );
  CFD1XL \buffer_reg[235]  ( .D(n5844), .CP(clk), .QN(n8048) );
  CFD1XL \buffer_reg[234]  ( .D(n5834), .CP(clk), .QN(n8049) );
  CFD1XL \buffer_reg[233]  ( .D(n5832), .CP(clk), .QN(n8050) );
  CFD1XL \buffer_reg[232]  ( .D(n5828), .CP(clk), .QN(n8051) );
  CFD1XL \buffer_reg[231]  ( .D(n5816), .CP(clk), .QN(n8052) );
  CFD1XL \buffer_reg[230]  ( .D(n5812), .CP(clk), .QN(n8053) );
  CFD1XL \buffer_reg[229]  ( .D(n5802), .CP(clk), .QN(n8054) );
  CFD1XL \buffer_reg[228]  ( .D(n5800), .CP(clk), .QN(n8055) );
  CFD1XL \buffer_reg[227]  ( .D(n5796), .CP(clk), .QN(n8056) );
  CFD1XL \buffer_reg[226]  ( .D(n5792), .CP(clk), .QN(n8057) );
  CFD1XL \buffer_reg[225]  ( .D(n5790), .CP(clk), .QN(n8058) );
  CFD1XL \buffer_reg[224]  ( .D(n5784), .CP(clk), .QN(n8059) );
  CFD1XL \buffer_reg[223]  ( .D(n5770), .CP(clk), .QN(n8060) );
  CFD1XL \buffer_reg[222]  ( .D(n5768), .CP(clk), .QN(n8061) );
  CFD1XL \buffer_reg[221]  ( .D(n5764), .CP(clk), .QN(n8062) );
  CFD1XL \buffer_reg[220]  ( .D(n5752), .CP(clk), .QN(n8063) );
  CFD1XL \buffer_reg[219]  ( .D(n5748), .CP(clk), .QN(n8064) );
  CFD1XL \buffer_reg[218]  ( .D(n5642), .CP(clk), .QN(n8065) );
  CFD1XL \buffer_reg[217]  ( .D(n5636), .CP(clk), .QN(n8066) );
  CFD1XL \buffer_reg[216]  ( .D(n5624), .CP(clk), .QN(n8067) );
  CFD1XL \buffer_reg[215]  ( .D(n5600), .CP(clk), .QN(n8068) );
  CFD1XL \buffer_reg[214]  ( .D(n5598), .CP(clk), .QN(n8069) );
  CFD1XL \buffer_reg[207]  ( .D(n5588), .CP(clk), .QN(n8076) );
  CFD1XL \buffer_reg[206]  ( .D(n5578), .CP(clk), .QN(n8077) );
  CFD1XL \buffer_reg[203]  ( .D(n5576), .CP(clk), .QN(n8080) );
  CFD1XL \buffer_reg[202]  ( .D(n5572), .CP(clk), .QN(n8081) );
  CFD1XL \buffer_reg[201]  ( .D(n5536), .CP(clk), .QN(n8082) );
  CFD1XL \buffer_reg[200]  ( .D(n5534), .CP(clk), .QN(n8083) );
  CFD1XL \buffer_reg[199]  ( .D(n5515), .CP(clk), .QN(n8084) );
  CFD1XL \buffer_reg[198]  ( .D(n5509), .CP(clk), .QN(n8085) );
  CFD1XL \buffer_reg[197]  ( .D(n5497), .CP(clk), .QN(n8086) );
  CFD1XL \buffer_reg[196]  ( .D(n5465), .CP(clk), .QN(n8087) );
  CFD1XL \buffer_reg[195]  ( .D(n5461), .CP(clk), .QN(n8088) );
  CFD1XL \buffer_reg[194]  ( .D(n5434), .CP(clk), .QN(n8089) );
  CFD1XL \buffer_reg[193]  ( .D(n5420), .CP(clk), .QN(n8090) );
  CFD1XL \buffer_reg[192]  ( .D(n5418), .CP(clk), .QN(n8091) );
  CFD1XL \buffer_reg[127]  ( .D(n5414), .CP(clk), .QN(n8156) );
  CFD1XL \buffer_reg[126]  ( .D(n5412), .CP(clk), .QN(n8157) );
  CFD1XL \buffer_reg[125]  ( .D(n5402), .CP(clk), .QN(n8158) );
  CFD1XL \buffer_reg[124]  ( .D(n5398), .CP(clk), .QN(n8159) );
  CFD1XL \buffer_reg[123]  ( .D(n5388), .CP(clk), .QN(n8160) );
  CFD1XL \buffer_reg[122]  ( .D(n5386), .CP(clk), .QN(n8161) );
  CFD1XL \buffer_reg[121]  ( .D(n5382), .CP(clk), .QN(n8162) );
  CFD1XL \buffer_reg[120]  ( .D(n5378), .CP(clk), .QN(n8163) );
  CFD1XL \buffer_reg[119]  ( .D(n5376), .CP(clk), .QN(n8164) );
  CFD1XL \buffer_reg[118]  ( .D(n5370), .CP(clk), .QN(n8165) );
  CFD1XL \buffer_reg[111]  ( .D(n5366), .CP(clk), .QN(n8172) );
  CFD1XL \buffer_reg[110]  ( .D(n5356), .CP(clk), .QN(n8173) );
  CFD1XL \buffer_reg[107]  ( .D(n5354), .CP(clk), .QN(n8176) );
  CFD1XL \buffer_reg[106]  ( .D(n5350), .CP(clk), .QN(n8177) );
  CFD1XL \buffer_reg[105]  ( .D(n5338), .CP(clk), .QN(n8178) );
  CFD1XL \buffer_reg[104]  ( .D(n5334), .CP(clk), .QN(n8179) );
  CFD1XL \buffer_reg[103]  ( .D(n5324), .CP(clk), .QN(n8180) );
  CFD1XL \buffer_reg[102]  ( .D(n5322), .CP(clk), .QN(n8181) );
  CFD1XL \buffer_reg[101]  ( .D(n5318), .CP(clk), .QN(n8182) );
  CFD1XL \buffer_reg[100]  ( .D(n5314), .CP(clk), .QN(n8183) );
  CFD1XL \buffer_reg[99]  ( .D(n5312), .CP(clk), .QN(n8184) );
  CFD1XL \buffer_reg[98]  ( .D(n5306), .CP(clk), .QN(n8185) );
  CFD1XL \buffer_reg[97]  ( .D(n5292), .CP(clk), .QN(n8186) );
  CFD1XL \buffer_reg[96]  ( .D(n5290), .CP(clk), .QN(n8187) );
  CFD1XL \buffer_reg[95]  ( .D(n5286), .CP(clk), .QN(n8188) );
  CFD1XL \buffer_reg[94]  ( .D(n5274), .CP(clk), .QN(n8189) );
  CFD1XL \buffer_reg[93]  ( .D(n5270), .CP(clk), .QN(n8190) );
  CFD1XL \buffer_reg[92]  ( .D(n5164), .CP(clk), .QN(n8191) );
  CFD1XL \buffer_reg[91]  ( .D(n5162), .CP(clk), .QN(n8192) );
  CFD1XL \buffer_reg[90]  ( .D(n5158), .CP(clk), .QN(n8193) );
  CFD1XL \buffer_reg[89]  ( .D(n5122), .CP(clk), .QN(n8194) );
  CFD1XL \buffer_reg[88]  ( .D(n5120), .CP(clk), .QN(n8195) );
  CFD1XL \buffer_reg[87]  ( .D(n5100), .CP(clk), .QN(n8196) );
  CFD1XL \buffer_reg[86]  ( .D(n5098), .CP(clk), .QN(n8197) );
  CFD1XL \buffer_reg[79]  ( .D(n5094), .CP(clk), .QN(n8204) );
  CFD1XL \buffer_reg[78]  ( .D(n5036), .CP(clk), .QN(n8205) );
  CFD1XL \buffer_reg[75]  ( .D(n5034), .CP(clk), .QN(n8208) );
  CFD1XL \buffer_reg[74]  ( .D(n5030), .CP(clk), .QN(n8209) );
  CFD1XL \buffer_reg[73]  ( .D(n4954), .CP(clk), .QN(n8210) );
  CFD1XL \buffer_reg[72]  ( .D(n4950), .CP(clk), .QN(n8211) );
  CFD1XL \buffer_reg[71]  ( .D(n4934), .CP(clk), .QN(n8212) );
  CFD1XL \buffer_reg[70]  ( .D(n4910), .CP(clk), .QN(n8213) );
  CFD1XL \buffer_reg[69]  ( .D(n4908), .CP(clk), .QN(n8214) );
  CFD1XL \buffer_reg[68]  ( .D(n4906), .CP(clk), .QN(n8215) );
  CFD1XL \buffer_reg[67]  ( .D(n4902), .CP(clk), .QN(n8216) );
  CFD1XL \buffer_reg[66]  ( .D(n4900), .CP(clk), .QN(n8217) );
  CFD1XL \buffer_reg[65]  ( .D(n4892), .CP(clk), .QN(n8218) );
  CFD1XL \buffer_reg[64]  ( .D(n4890), .CP(clk), .QN(n8219) );
  CFD1XL \buffer_reg[1036]  ( .D(n4886), .CP(clk), .QN(n7225) );
  CFD1XL \buffer_reg[31]  ( .D(n4876), .CP(clk), .QN(n8252) );
  CFD1XL \buffer_reg[30]  ( .D(n4874), .CP(clk), .QN(n8253) );
  CFD1XL \buffer_reg[29]  ( .D(n4870), .CP(clk), .QN(n8254) );
  CFD1XL \buffer_reg[28]  ( .D(n4866), .CP(clk), .QN(n8255) );
  CFD1XL \buffer_reg[27]  ( .D(n4864), .CP(clk), .QN(n8256) );
  CFD1XL \buffer_reg[26]  ( .D(n4858), .CP(clk), .QN(n8257) );
  CFD1XL \buffer_reg[25]  ( .D(n4854), .CP(clk), .QN(n8258) );
  CFD1XL \buffer_reg[24]  ( .D(n4844), .CP(clk), .QN(n8259) );
  CFD1XL \buffer_reg[23]  ( .D(n4842), .CP(clk), .QN(n8260) );
  CFD1XL \buffer_reg[22]  ( .D(n4838), .CP(clk), .QN(n8261) );
  CFD1XL \buffer_reg[21]  ( .D(n4826), .CP(clk), .QN(n8262) );
  CFD1XL \buffer_reg[20]  ( .D(n4822), .CP(clk), .QN(n8263) );
  CFD1XL \buffer_reg[19]  ( .D(n4812), .CP(clk), .QN(n8264) );
  CFD1XL \buffer_reg[18]  ( .D(n4810), .CP(clk), .QN(n8265) );
  CFD1XL \buffer_reg[17]  ( .D(n4806), .CP(clk), .QN(n8266) );
  CFD1XL \buffer_reg[16]  ( .D(n4802), .CP(clk), .QN(n8267) );
  CFD1XL \buffer_reg[15]  ( .D(n4800), .CP(clk), .Q(n2844), .QN(n8268) );
  CFD1XL \buffer_reg[14]  ( .D(n4780), .CP(clk), .Q(n2381), .QN(n8269) );
  CFD1XL \buffer_reg[13]  ( .D(n4778), .CP(clk), .Q(n2965), .QN(n8270) );
  CFD1XL \buffer_reg[12]  ( .D(n4774), .CP(clk), .QN(n8271) );
  CFD1XL \buffer_reg[11]  ( .D(n4772), .CP(clk), .Q(n2714), .QN(n8272) );
  CFD1XL \buffer_reg[10]  ( .D(n4762), .CP(clk), .Q(n2502), .QN(n8273) );
  CFD1XL \buffer_reg[9]  ( .D(n4758), .CP(clk), .Q(n3047), .QN(n8274) );
  CFD1XL \buffer_reg[8]  ( .D(n4742), .CP(clk), .Q(n2292), .QN(n8275) );
  CFD1XL \buffer_reg[7]  ( .D(n4652), .CP(clk), .Q(n2916), .QN(n8276) );
  CFD1QXL \rd_ptr_reg[7]  ( .D(n4283), .CP(clk), .Q(rd_ptr[7]) );
  CFD1QXL \rd_ptr_reg[9]  ( .D(n4280), .CP(clk), .Q(rd_ptr[9]) );
  CFD1QX1 \rd_ptr_reg[8]  ( .D(n4238), .CP(clk), .Q(rd_ptr[8]) );
  CAOR2XL U3310 ( .A(N16598), .B(n6164), .C(n7092), .D(rd_ptr[8]), .Z(n3191)
         );
  CNIVX1 U3311 ( .A(n3191), .Z(n4238) );
  CNIVX1 U3312 ( .A(rd_ptr[7]), .Z(n4239) );
  CAOR2XL U3313 ( .A(N16599), .B(n3173), .C(n4), .D(rd_ptr[9]), .Z(n3190) );
  CENXL U3314 ( .A(rd_ptr[9]), .B(n6159), .Z(N16599) );
  CNR2IXL U3315 ( .B(rd_ptr[9]), .A(n8311), .Z(n388) );
  CNR2X1 U3316 ( .A(rd_ptr[8]), .B(rd_ptr[9]), .Z(n387) );
  CIVX2 U3317 ( .A(n4239), .Z(n8310) );
  CNR3XL U3318 ( .A(n911), .B(n908), .C(n6157), .Z(n907) );
  CND2IX1 U3319 ( .B(n382), .A(n8310), .Z(n84) );
  CNIVX2 U3320 ( .A(n388), .Z(n7093) );
  COND1XL U3321 ( .A(n7247), .B(n8293), .C(n790), .Z(n289) );
  COND1XL U3322 ( .A(rd_ptr[3]), .B(n355), .C(n356), .Z(n226) );
  CND3XL U3323 ( .A(n6151), .B(n6152), .C(n6153), .Z(n6154) );
  CIVX2 U3324 ( .A(n4242), .Z(n7124) );
  CAN2X1 U3325 ( .A(n7093), .B(n4239), .Z(n4240) );
  CAN2X1 U3326 ( .A(n386), .B(n8310), .Z(n4241) );
  CAN2X1 U3327 ( .A(n387), .B(n4239), .Z(n4242) );
  CNIVXL U3328 ( .A(n284), .Z(n4243) );
  CNIVX1 U3329 ( .A(n4262), .Z(n4244) );
  CNIVX1 U3330 ( .A(n4268), .Z(n4245) );
  CNIVX1 U3331 ( .A(n4269), .Z(n4246) );
  CNIVX1 U3332 ( .A(n4263), .Z(n4247) );
  CNIVX1 U3333 ( .A(n4265), .Z(n4248) );
  CNIVX1 U3334 ( .A(n4266), .Z(n4249) );
  CNIVX1 U3335 ( .A(n4264), .Z(n4250) );
  CNIVX1 U3336 ( .A(n4267), .Z(n4251) );
  CIVDXL U3337 ( .A(pushout_stg_1), .Z1(n4253) );
  CNIVX1 U3338 ( .A(n4253), .Z(n4252) );
  CAOR2X4 U3339 ( .A(n6165), .B(n6160), .C(lenout[0]), .D(n2234), .Z(N118) );
  CAOR2X4 U3340 ( .A(n3173), .B(n6161), .C(lenout[1]), .D(n2234), .Z(N119) );
  CAOR2X4 U3341 ( .A(n3173), .B(n6162), .C(lenout[2]), .D(n2234), .Z(N120) );
  CAOR2X4 U3342 ( .A(n6165), .B(n6163), .C(lenout[3]), .D(n2234), .Z(N121) );
  CIVX3 U3343 ( .A(buffer[137]), .Z(n8146) );
  CIVX3 U3344 ( .A(buffer[129]), .Z(n8154) );
  CIVX3 U3345 ( .A(buffer[257]), .Z(n8026) );
  CIVX3 U3346 ( .A(buffer[259]), .Z(n8024) );
  CIVX3 U3347 ( .A(buffer[261]), .Z(n8022) );
  CIVX3 U3348 ( .A(buffer[263]), .Z(n8020) );
  CIVX3 U3349 ( .A(buffer[265]), .Z(n8018) );
  CIVX3 U3350 ( .A(buffer[269]), .Z(n8014) );
  CIVX3 U3351 ( .A(buffer[256]), .Z(n8027) );
  CIVX3 U3352 ( .A(buffer[258]), .Z(n8025) );
  CIVX3 U3353 ( .A(buffer[260]), .Z(n8023) );
  CIVX3 U3354 ( .A(buffer[262]), .Z(n8021) );
  CIVX3 U3355 ( .A(buffer[266]), .Z(n8017) );
  CIVX3 U3356 ( .A(buffer[513]), .Z(n7770) );
  CIVX3 U3357 ( .A(buffer[512]), .Z(n7771) );
  CIVX3 U3358 ( .A(buffer[514]), .Z(n7769) );
  CIVX3 U3359 ( .A(buffer[516]), .Z(n7767) );
  CIVX3 U3360 ( .A(buffer[780]), .Z(n7503) );
  CIVX3 U3361 ( .A(buffer[1024]), .Z(n7243) );
  CIVX3 U3362 ( .A(buffer[1026]), .Z(n7239) );
  CIVX3 U3363 ( .A(buffer[1027]), .Z(n7238) );
  CIVX3 U3364 ( .A(buffer[1028]), .Z(n7236) );
  CIVX3 U3365 ( .A(buffer[1029]), .Z(n7235) );
  CIVX3 U3366 ( .A(buffer[1030]), .Z(n7234) );
  CIVX3 U3367 ( .A(buffer[1031]), .Z(n7232) );
  CIVX3 U3368 ( .A(buffer[1032]), .Z(n7231) );
  CIVX3 U3369 ( .A(buffer[1033]), .Z(n7229) );
  CIVX3 U3370 ( .A(buffer[1034]), .Z(n7228) );
  CIVX3 U3371 ( .A(buffer[896]), .Z(n7387) );
  CIVX3 U3372 ( .A(buffer[897]), .Z(n7386) );
  CIVX3 U3373 ( .A(buffer[898]), .Z(n7385) );
  CIVX3 U3374 ( .A(buffer[899]), .Z(n7384) );
  CIVX3 U3375 ( .A(buffer[900]), .Z(n7383) );
  CIVX3 U3376 ( .A(buffer[901]), .Z(n7382) );
  CIVX3 U3377 ( .A(buffer[902]), .Z(n7381) );
  CIVX3 U3378 ( .A(buffer[903]), .Z(n7380) );
  CIVX3 U3379 ( .A(buffer[904]), .Z(n7379) );
  CIVX3 U3380 ( .A(buffer[905]), .Z(n7378) );
  CIVX3 U3381 ( .A(buffer[906]), .Z(n7377) );
  CIVX3 U3382 ( .A(buffer[907]), .Z(n7376) );
  CIVX3 U3383 ( .A(buffer[909]), .Z(n7374) );
  CIVX3 U3384 ( .A(buffer[393]), .Z(n7890) );
  CIVX3 U3385 ( .A(buffer[1025]), .Z(n7242) );
  CIVX3 U3386 ( .A(buffer[128]), .Z(n8155) );
  CIVX3 U3387 ( .A(buffer[130]), .Z(n8153) );
  CIVX3 U3388 ( .A(buffer[131]), .Z(n8152) );
  CIVX3 U3389 ( .A(buffer[132]), .Z(n8151) );
  CIVX3 U3390 ( .A(buffer[133]), .Z(n8150) );
  CIVX3 U3391 ( .A(buffer[134]), .Z(n8149) );
  CIVX3 U3392 ( .A(buffer[135]), .Z(n8148) );
  CIVX3 U3393 ( .A(buffer[136]), .Z(n8147) );
  CIVX3 U3394 ( .A(buffer[138]), .Z(n8145) );
  CIVX3 U3395 ( .A(buffer[139]), .Z(n8144) );
  CIVX3 U3396 ( .A(buffer[141]), .Z(n8142) );
  CIVX3 U3397 ( .A(buffer[384]), .Z(n7899) );
  CIVX3 U3398 ( .A(buffer[385]), .Z(n7898) );
  CIVX3 U3399 ( .A(buffer[386]), .Z(n7897) );
  CIVX3 U3400 ( .A(buffer[387]), .Z(n7896) );
  CIVX3 U3401 ( .A(buffer[388]), .Z(n7895) );
  CIVX3 U3402 ( .A(buffer[389]), .Z(n7894) );
  CIVX3 U3403 ( .A(buffer[390]), .Z(n7893) );
  CIVX3 U3404 ( .A(buffer[391]), .Z(n7892) );
  CIVX3 U3405 ( .A(buffer[392]), .Z(n7891) );
  CIVX3 U3406 ( .A(buffer[394]), .Z(n7889) );
  CIVX3 U3407 ( .A(buffer[395]), .Z(n7888) );
  CIVX3 U3408 ( .A(buffer[397]), .Z(n7886) );
  CIVX3 U3409 ( .A(buffer[140]), .Z(n8143) );
  COND2XL U3410 ( .A(n7643), .B(n6510), .C(n7206), .D(n6501), .Z(n3840) );
  CIVX3 U3411 ( .A(buffer[640]), .Z(n7643) );
  COND2XL U3412 ( .A(n7642), .B(n6511), .C(n7205), .D(n6502), .Z(n3841) );
  CIVX3 U3413 ( .A(buffer[641]), .Z(n7642) );
  COND2XL U3414 ( .A(n7641), .B(n6512), .C(n7204), .D(n6501), .Z(n3842) );
  CIVX3 U3415 ( .A(buffer[642]), .Z(n7641) );
  COND2XL U3416 ( .A(n7640), .B(n6513), .C(n7203), .D(n6502), .Z(n3843) );
  CIVX3 U3417 ( .A(buffer[643]), .Z(n7640) );
  COND2XL U3418 ( .A(n7639), .B(n6514), .C(n7202), .D(n6503), .Z(n3844) );
  CIVX3 U3419 ( .A(buffer[644]), .Z(n7639) );
  COND2XL U3420 ( .A(n7638), .B(n6515), .C(n7201), .D(n6501), .Z(n3845) );
  CIVX3 U3421 ( .A(buffer[645]), .Z(n7638) );
  COND2XL U3422 ( .A(n7637), .B(n6517), .C(n7200), .D(n6503), .Z(n3846) );
  CIVX3 U3423 ( .A(buffer[646]), .Z(n7637) );
  COND2XL U3424 ( .A(n7636), .B(n6518), .C(n7199), .D(n6504), .Z(n3847) );
  CIVX3 U3425 ( .A(buffer[647]), .Z(n7636) );
  COND2XL U3426 ( .A(n7635), .B(n6519), .C(n7198), .D(n6504), .Z(n3848) );
  CIVX3 U3427 ( .A(buffer[648]), .Z(n7635) );
  COND2XL U3428 ( .A(n7634), .B(n6520), .C(n7197), .D(n6505), .Z(n3849) );
  CIVX3 U3429 ( .A(buffer[649]), .Z(n7634) );
  COND2XL U3430 ( .A(n7633), .B(n6521), .C(n7196), .D(n6506), .Z(n3850) );
  CIVX3 U3431 ( .A(buffer[650]), .Z(n7633) );
  COND2XL U3432 ( .A(n7632), .B(n6522), .C(n7195), .D(n6502), .Z(n3851) );
  CIVX3 U3433 ( .A(buffer[651]), .Z(n7632) );
  CIVX3 U3434 ( .A(buffer[652]), .Z(n7631) );
  COND2XL U3435 ( .A(n7630), .B(n6525), .C(n7193), .D(n6506), .Z(n3853) );
  CIVX3 U3436 ( .A(buffer[653]), .Z(n7630) );
  CIVX3 U3437 ( .A(buffer[908]), .Z(n7375) );
  CIVDXL U3438 ( .A(lenout_stg_1[0]), .Z1(n4255) );
  CNIVX1 U3439 ( .A(n4255), .Z(n4254) );
  CIVDXL U3440 ( .A(lenout_stg_1[1]), .Z1(n4257) );
  CNIVX1 U3441 ( .A(n4257), .Z(n4256) );
  CIVDXL U3442 ( .A(lenout_stg_1[2]), .Z1(n4259) );
  CNIVX1 U3443 ( .A(n4259), .Z(n4258) );
  CIVDXL U3444 ( .A(lenout_stg_1[3]), .Z1(n4261) );
  CNIVX1 U3445 ( .A(n4261), .Z(n4260) );
  CIVX3 U3446 ( .A(buffer[1037]), .Z(n7223) );
  CNIVX1 U3447 ( .A(dataout_stg_1[7]), .Z(n4262) );
  CNIVX1 U3448 ( .A(dataout_stg_1[10]), .Z(n4263) );
  CNIVX1 U3449 ( .A(dataout_stg_1[13]), .Z(n4264) );
  CNIVX1 U3450 ( .A(dataout_stg_1[11]), .Z(n4265) );
  CAOR2X2 U3451 ( .A(n4265), .B(n7091), .C(n7211), .D(n130), .Z(n3178) );
  CNIVX1 U3452 ( .A(dataout_stg_1[12]), .Z(n4266) );
  CAOR2X2 U3453 ( .A(n4266), .B(n7092), .C(n7211), .D(n96), .Z(n3177) );
  CNIVX1 U3454 ( .A(dataout_stg_1[14]), .Z(n4267) );
  CNIVX1 U3455 ( .A(dataout_stg_1[8]), .Z(n4268) );
  CNIVX1 U3456 ( .A(dataout_stg_1[9]), .Z(n4269) );
  CNIVX1 U3457 ( .A(n4271), .Z(n4270) );
  CNIVX1 U3458 ( .A(n3369), .Z(n4271) );
  CNIVX1 U3459 ( .A(n4273), .Z(n4272) );
  CNIVX1 U3460 ( .A(n3370), .Z(n4273) );
  CNIVX1 U3461 ( .A(n4275), .Z(n4274) );
  CNIVX1 U3462 ( .A(n3374), .Z(n4275) );
  CNIVX1 U3463 ( .A(n4277), .Z(n4276) );
  CNIVX1 U3464 ( .A(n3375), .Z(n4277) );
  CNIVX1 U3465 ( .A(n4279), .Z(n4278) );
  CNIVX1 U3466 ( .A(n3365), .Z(n4279) );
  CNIVX1 U3467 ( .A(n3190), .Z(n4280) );
  CNIVX1 U3468 ( .A(n4282), .Z(n4281) );
  CNIVX1 U3469 ( .A(dataout_stg_1[0]), .Z(n4282) );
  CNIVX1 U3470 ( .A(n3192), .Z(n4283) );
  CNIVX1 U3471 ( .A(n4285), .Z(n4284) );
  CNIVX1 U3472 ( .A(dataout_stg_1[1]), .Z(n4285) );
  CNIVX1 U3473 ( .A(n4287), .Z(n4286) );
  CNIVX1 U3474 ( .A(dataout_stg_1[2]), .Z(n4287) );
  CNIVX1 U3475 ( .A(n4289), .Z(n4288) );
  CNIVX1 U3476 ( .A(dataout_stg_1[3]), .Z(n4289) );
  CNIVX1 U3477 ( .A(n4291), .Z(n4290) );
  CNIVX1 U3478 ( .A(dataout_stg_1[4]), .Z(n4291) );
  CNIVX1 U3479 ( .A(n4293), .Z(n4292) );
  CNIVX1 U3480 ( .A(dataout_stg_1[5]), .Z(n4293) );
  CNIVX1 U3481 ( .A(n4295), .Z(n4294) );
  CNIVX1 U3482 ( .A(n3410), .Z(n4295) );
  CNIVX1 U3483 ( .A(n4297), .Z(n4296) );
  CNIVX1 U3484 ( .A(n3411), .Z(n4297) );
  CNIVX1 U3485 ( .A(n4299), .Z(n4298) );
  CNIVX1 U3486 ( .A(n3412), .Z(n4299) );
  CNIVX1 U3487 ( .A(n4301), .Z(n4300) );
  CNIVX1 U3488 ( .A(n3413), .Z(n4301) );
  CNIVX1 U3489 ( .A(n4303), .Z(n4302) );
  CNIVX1 U3490 ( .A(n3442), .Z(n4303) );
  CNIVX1 U3491 ( .A(n4305), .Z(n4304) );
  CNIVX1 U3492 ( .A(n3443), .Z(n4305) );
  CNIVX1 U3493 ( .A(n4307), .Z(n4306) );
  CNIVX1 U3494 ( .A(n3444), .Z(n4307) );
  CNIVX1 U3495 ( .A(n4309), .Z(n4308) );
  CNIVX1 U3496 ( .A(n3445), .Z(n4309) );
  CNIVX1 U3497 ( .A(n4311), .Z(n4310) );
  CNIVX1 U3498 ( .A(n3808), .Z(n4311) );
  CNIVX1 U3499 ( .A(n4313), .Z(n4312) );
  CNIVX1 U3500 ( .A(n3809), .Z(n4313) );
  CNIVX1 U3501 ( .A(n4315), .Z(n4314) );
  CNIVX1 U3502 ( .A(n3344), .Z(n4315) );
  CNIVX1 U3503 ( .A(n4317), .Z(n4316) );
  CNIVX1 U3504 ( .A(n3345), .Z(n4317) );
  CNIVX1 U3505 ( .A(n4319), .Z(n4318) );
  CNIVX1 U3506 ( .A(n3909), .Z(n4319) );
  CNIVX1 U3507 ( .A(n4321), .Z(n4320) );
  CNIVX1 U3508 ( .A(n3372), .Z(n4321) );
  CNIVX1 U3509 ( .A(n4323), .Z(n4322) );
  CNIVX1 U3510 ( .A(n3373), .Z(n4323) );
  CNIVX1 U3511 ( .A(n4325), .Z(n4324) );
  CNIVX1 U3512 ( .A(n3376), .Z(n4325) );
  CNIVX1 U3513 ( .A(n4327), .Z(n4326) );
  CNIVX1 U3514 ( .A(n3910), .Z(n4327) );
  CNIVX1 U3515 ( .A(n4329), .Z(n4328) );
  CNIVX1 U3516 ( .A(n3911), .Z(n4329) );
  CNIVX1 U3517 ( .A(n4331), .Z(n4330) );
  CNIVX1 U3518 ( .A(n3912), .Z(n4331) );
  CNIVX1 U3519 ( .A(n4333), .Z(n4332) );
  CNIVX1 U3520 ( .A(n3913), .Z(n4333) );
  CNIVX1 U3521 ( .A(n4335), .Z(n4334) );
  CNIVX1 U3522 ( .A(n3914), .Z(n4335) );
  CNIVX1 U3523 ( .A(n4337), .Z(n4336) );
  CNIVX1 U3524 ( .A(n3915), .Z(n4337) );
  CNIVX1 U3525 ( .A(n4339), .Z(n4338) );
  CNIVX1 U3526 ( .A(n3918), .Z(n4339) );
  CNIVX1 U3527 ( .A(n4341), .Z(n4340) );
  CNIVX1 U3528 ( .A(n3919), .Z(n4341) );
  CNIVX1 U3529 ( .A(n4343), .Z(n4342) );
  CNIVX1 U3530 ( .A(n3926), .Z(n4343) );
  CNIVX1 U3531 ( .A(n4345), .Z(n4344) );
  CNIVX1 U3532 ( .A(n3927), .Z(n4345) );
  CNIVX1 U3533 ( .A(n4347), .Z(n4346) );
  CNIVX1 U3534 ( .A(n3928), .Z(n4347) );
  CNIVX1 U3535 ( .A(n4349), .Z(n4348) );
  CNIVX1 U3536 ( .A(n3929), .Z(n4349) );
  CNIVX1 U3537 ( .A(n4351), .Z(n4350) );
  CNIVX1 U3538 ( .A(n3930), .Z(n4351) );
  CNIVX1 U3539 ( .A(n4353), .Z(n4352) );
  CNIVX1 U3540 ( .A(n3931), .Z(n4353) );
  CNIVX1 U3541 ( .A(n4355), .Z(n4354) );
  CNIVX1 U3542 ( .A(n3932), .Z(n4355) );
  CNIVX1 U3543 ( .A(n4357), .Z(n4356) );
  CNIVX1 U3544 ( .A(n3933), .Z(n4357) );
  CNIVX1 U3545 ( .A(n4359), .Z(n4358) );
  CNIVX1 U3546 ( .A(n3934), .Z(n4359) );
  CNIVX1 U3547 ( .A(n4361), .Z(n4360) );
  CNIVX1 U3548 ( .A(n3935), .Z(n4361) );
  CNIVX1 U3549 ( .A(n4363), .Z(n4362) );
  CNIVX1 U3550 ( .A(n3936), .Z(n4363) );
  CNIVX1 U3551 ( .A(n4365), .Z(n4364) );
  CNIVX1 U3552 ( .A(n3937), .Z(n4365) );
  CNIVX1 U3553 ( .A(n4367), .Z(n4366) );
  CNIVX1 U3554 ( .A(n3938), .Z(n4367) );
  CNIVX1 U3555 ( .A(n4369), .Z(n4368) );
  CNIVX1 U3556 ( .A(n3939), .Z(n4369) );
  CNIVX1 U3557 ( .A(n4371), .Z(n4370) );
  CNIVX1 U3558 ( .A(n3940), .Z(n4371) );
  CNIVX1 U3559 ( .A(n4373), .Z(n4372) );
  CNIVX1 U3560 ( .A(n3941), .Z(n4373) );
  CNIVX1 U3561 ( .A(n4375), .Z(n4374) );
  CNIVX1 U3562 ( .A(n3942), .Z(n4375) );
  CNIVX1 U3563 ( .A(n4377), .Z(n4376) );
  CNIVX1 U3564 ( .A(n3943), .Z(n4377) );
  CNIVX1 U3565 ( .A(n4379), .Z(n4378) );
  CNIVX1 U3566 ( .A(n3944), .Z(n4379) );
  CNIVX1 U3567 ( .A(n4381), .Z(n4380) );
  CNIVX1 U3568 ( .A(n3945), .Z(n4381) );
  CNIVX1 U3569 ( .A(n4383), .Z(n4382) );
  CNIVX1 U3570 ( .A(n3946), .Z(n4383) );
  CNIVX1 U3571 ( .A(n4385), .Z(n4384) );
  CNIVX1 U3572 ( .A(n3947), .Z(n4385) );
  CNIVX1 U3573 ( .A(n4387), .Z(n4386) );
  CNIVX1 U3574 ( .A(n3950), .Z(n4387) );
  CNIVX1 U3575 ( .A(n4389), .Z(n4388) );
  CNIVX1 U3576 ( .A(n3951), .Z(n4389) );
  CNIVX1 U3577 ( .A(n4391), .Z(n4390) );
  CNIVX1 U3578 ( .A(n3958), .Z(n4391) );
  CNIVX1 U3579 ( .A(n4393), .Z(n4392) );
  CNIVX1 U3580 ( .A(n3959), .Z(n4393) );
  CNIVX1 U3581 ( .A(n4395), .Z(n4394) );
  CNIVX1 U3582 ( .A(n3960), .Z(n4395) );
  CNIVX1 U3583 ( .A(n4397), .Z(n4396) );
  CNIVX1 U3584 ( .A(n3961), .Z(n4397) );
  CNIVX1 U3585 ( .A(n4399), .Z(n4398) );
  CNIVX1 U3586 ( .A(n3962), .Z(n4399) );
  CNIVX1 U3587 ( .A(n4401), .Z(n4400) );
  CNIVX1 U3588 ( .A(n3963), .Z(n4401) );
  CNIVX1 U3589 ( .A(n4403), .Z(n4402) );
  CNIVX1 U3590 ( .A(n3964), .Z(n4403) );
  CNIVX1 U3591 ( .A(n4405), .Z(n4404) );
  CNIVX1 U3592 ( .A(n3965), .Z(n4405) );
  CNIVX1 U3593 ( .A(n4407), .Z(n4406) );
  CNIVX1 U3594 ( .A(n3966), .Z(n4407) );
  CNIVX1 U3595 ( .A(n4409), .Z(n4408) );
  CNIVX1 U3596 ( .A(n3967), .Z(n4409) );
  CNIVX1 U3597 ( .A(n4411), .Z(n4410) );
  CNIVX1 U3598 ( .A(n3854), .Z(n4411) );
  CNIVX1 U3599 ( .A(n4413), .Z(n4412) );
  CNIVX1 U3600 ( .A(n3855), .Z(n4413) );
  CNIVX1 U3601 ( .A(n4415), .Z(n4414) );
  CNIVX1 U3602 ( .A(n3862), .Z(n4415) );
  CNIVX1 U3603 ( .A(n4417), .Z(n4416) );
  CNIVX1 U3604 ( .A(n3863), .Z(n4417) );
  CNIVX1 U3605 ( .A(n4419), .Z(n4418) );
  CNIVX1 U3606 ( .A(n3864), .Z(n4419) );
  CNIVX1 U3607 ( .A(n4421), .Z(n4420) );
  CNIVX1 U3608 ( .A(n3865), .Z(n4421) );
  CNIVX1 U3609 ( .A(n4423), .Z(n4422) );
  CNIVX1 U3610 ( .A(n3866), .Z(n4423) );
  CNIVX1 U3611 ( .A(n4425), .Z(n4424) );
  CNIVX1 U3612 ( .A(n3867), .Z(n4425) );
  CNIVX1 U3613 ( .A(n4427), .Z(n4426) );
  CNIVX1 U3614 ( .A(n3868), .Z(n4427) );
  CNIVX1 U3615 ( .A(n4429), .Z(n4428) );
  CNIVX1 U3616 ( .A(n3869), .Z(n4429) );
  CNIVX1 U3617 ( .A(n4431), .Z(n4430) );
  CNIVX1 U3618 ( .A(n3870), .Z(n4431) );
  CNIVX1 U3619 ( .A(n4433), .Z(n4432) );
  CNIVX1 U3620 ( .A(n3871), .Z(n4433) );
  CNIVX1 U3621 ( .A(n4435), .Z(n4434) );
  CNIVX1 U3622 ( .A(n3872), .Z(n4435) );
  CNIVX1 U3623 ( .A(n4437), .Z(n4436) );
  CNIVX1 U3624 ( .A(n3873), .Z(n4437) );
  CNIVX1 U3625 ( .A(n4439), .Z(n4438) );
  CNIVX1 U3626 ( .A(n3874), .Z(n4439) );
  CNIVX1 U3627 ( .A(n4441), .Z(n4440) );
  CNIVX1 U3628 ( .A(n3875), .Z(n4441) );
  CNIVX1 U3629 ( .A(n4443), .Z(n4442) );
  CNIVX1 U3630 ( .A(n3876), .Z(n4443) );
  CNIVX1 U3631 ( .A(n4445), .Z(n4444) );
  CNIVX1 U3632 ( .A(n3877), .Z(n4445) );
  CNIVX1 U3633 ( .A(n4447), .Z(n4446) );
  CNIVX1 U3634 ( .A(n3878), .Z(n4447) );
  CNIVX1 U3635 ( .A(n4449), .Z(n4448) );
  CNIVX1 U3636 ( .A(n3879), .Z(n4449) );
  CNIVX1 U3637 ( .A(n4451), .Z(n4450) );
  CNIVX1 U3638 ( .A(n3880), .Z(n4451) );
  CNIVX1 U3639 ( .A(n4453), .Z(n4452) );
  CNIVX1 U3640 ( .A(n3881), .Z(n4453) );
  CNIVX1 U3641 ( .A(n4455), .Z(n4454) );
  CNIVX1 U3642 ( .A(n3882), .Z(n4455) );
  CNIVX1 U3643 ( .A(n4457), .Z(n4456) );
  CNIVX1 U3644 ( .A(n3883), .Z(n4457) );
  CNIVX1 U3645 ( .A(n4459), .Z(n4458) );
  CNIVX1 U3646 ( .A(n3886), .Z(n4459) );
  CNIVX1 U3647 ( .A(n4461), .Z(n4460) );
  CNIVX1 U3648 ( .A(n3887), .Z(n4461) );
  CNIVX1 U3649 ( .A(n4463), .Z(n4462) );
  CNIVX1 U3650 ( .A(n3894), .Z(n4463) );
  CNIVX1 U3651 ( .A(n4465), .Z(n4464) );
  CNIVX1 U3652 ( .A(n3895), .Z(n4465) );
  CNIVX1 U3653 ( .A(n4467), .Z(n4466) );
  CNIVX1 U3654 ( .A(n3896), .Z(n4467) );
  CNIVX1 U3655 ( .A(n4469), .Z(n4468) );
  CNIVX1 U3656 ( .A(n3897), .Z(n4469) );
  CNIVX1 U3657 ( .A(n4471), .Z(n4470) );
  CNIVX1 U3658 ( .A(n3898), .Z(n4471) );
  CNIVX1 U3659 ( .A(n4473), .Z(n4472) );
  CNIVX1 U3660 ( .A(n3899), .Z(n4473) );
  CNIVX1 U3661 ( .A(n4475), .Z(n4474) );
  CNIVX1 U3662 ( .A(n3900), .Z(n4475) );
  CNIVX1 U3663 ( .A(n4477), .Z(n4476) );
  CNIVX1 U3664 ( .A(n3901), .Z(n4477) );
  CNIVX1 U3665 ( .A(n4479), .Z(n4478) );
  CNIVX1 U3666 ( .A(n3814), .Z(n4479) );
  CNIVX1 U3667 ( .A(n4481), .Z(n4480) );
  CNIVX1 U3668 ( .A(n3815), .Z(n4481) );
  CNIVX1 U3669 ( .A(n4483), .Z(n4482) );
  CNIVX1 U3670 ( .A(n3816), .Z(n4483) );
  CNIVX1 U3671 ( .A(n4485), .Z(n4484) );
  CNIVX1 U3672 ( .A(n3817), .Z(n4485) );
  CNIVX1 U3673 ( .A(n4487), .Z(n4486) );
  CNIVX1 U3674 ( .A(n3818), .Z(n4487) );
  CNIVX1 U3675 ( .A(n4489), .Z(n4488) );
  CNIVX1 U3676 ( .A(n3819), .Z(n4489) );
  CNIVX1 U3677 ( .A(n4491), .Z(n4490) );
  CNIVX1 U3678 ( .A(n3822), .Z(n4491) );
  CNIVX1 U3679 ( .A(n4493), .Z(n4492) );
  CNIVX1 U3680 ( .A(n3823), .Z(n4493) );
  CNIVX1 U3681 ( .A(n4495), .Z(n4494) );
  CNIVX1 U3682 ( .A(n3830), .Z(n4495) );
  CNIVX1 U3683 ( .A(n4497), .Z(n4496) );
  CNIVX1 U3684 ( .A(n3831), .Z(n4497) );
  CNIVX1 U3685 ( .A(n4499), .Z(n4498) );
  CNIVX1 U3686 ( .A(n3832), .Z(n4499) );
  CNIVX1 U3687 ( .A(n4501), .Z(n4500) );
  CNIVX1 U3688 ( .A(n3811), .Z(n4501) );
  CNIVX1 U3689 ( .A(n4503), .Z(n4502) );
  CNIVX1 U3690 ( .A(n3776), .Z(n4503) );
  CNIVX1 U3691 ( .A(n4505), .Z(n4504) );
  CNIVX1 U3692 ( .A(n3902), .Z(n4505) );
  CNIVX1 U3693 ( .A(n4507), .Z(n4506) );
  CNIVX1 U3694 ( .A(n3903), .Z(n4507) );
  CNIVX1 U3695 ( .A(n4509), .Z(n4508) );
  CNIVX1 U3696 ( .A(n3788), .Z(n4509) );
  CNIVX1 U3697 ( .A(n4511), .Z(n4510) );
  CNIVX1 U3698 ( .A(n3789), .Z(n4511) );
  CNIVX1 U3699 ( .A(n4513), .Z(n4512) );
  CNIVX1 U3700 ( .A(n3792), .Z(n4513) );
  CNIVX1 U3701 ( .A(n4515), .Z(n4514) );
  CNIVX1 U3702 ( .A(n3793), .Z(n4515) );
  CNIVX1 U3703 ( .A(n4517), .Z(n4516) );
  CNIVX1 U3704 ( .A(n3820), .Z(n4517) );
  CNIVX1 U3705 ( .A(n4519), .Z(n4518) );
  CNIVX1 U3706 ( .A(n3821), .Z(n4519) );
  CNIVX1 U3707 ( .A(n4521), .Z(n4520) );
  CNIVX1 U3708 ( .A(n3824), .Z(n4521) );
  CNIVX1 U3709 ( .A(n4523), .Z(n4522) );
  CNIVX1 U3710 ( .A(n3825), .Z(n4523) );
  CNIVX1 U3711 ( .A(n4525), .Z(n4524) );
  CNIVX1 U3712 ( .A(n3916), .Z(n4525) );
  CNIVX1 U3713 ( .A(n4527), .Z(n4526) );
  CNIVX1 U3714 ( .A(n3917), .Z(n4527) );
  CNIVX1 U3715 ( .A(n4529), .Z(n4528) );
  CNIVX1 U3716 ( .A(n3920), .Z(n4529) );
  CNIVX1 U3717 ( .A(n4531), .Z(n4530) );
  CNIVX1 U3718 ( .A(n3921), .Z(n4531) );
  CNIVX1 U3719 ( .A(n4533), .Z(n4532) );
  CNIVX1 U3720 ( .A(n3948), .Z(n4533) );
  CNIVX1 U3721 ( .A(n4535), .Z(n4534) );
  CNIVX1 U3722 ( .A(n3949), .Z(n4535) );
  CNIVX1 U3723 ( .A(n4537), .Z(n4536) );
  CNIVX1 U3724 ( .A(n3952), .Z(n4537) );
  CNIVX1 U3725 ( .A(n4539), .Z(n4538) );
  CNIVX1 U3726 ( .A(n3953), .Z(n4539) );
  CNIVX1 U3727 ( .A(n4541), .Z(n4540) );
  CNIVX1 U3728 ( .A(n3794), .Z(n4541) );
  CNIVX1 U3729 ( .A(n4543), .Z(n4542) );
  CNIVX1 U3730 ( .A(n3795), .Z(n4543) );
  CNIVX1 U3731 ( .A(n4545), .Z(n4544) );
  CNIVX1 U3732 ( .A(n3796), .Z(n4545) );
  CNIVX1 U3733 ( .A(n4547), .Z(n4546) );
  CNIVX1 U3734 ( .A(n3797), .Z(n4547) );
  CNIVX1 U3735 ( .A(n4549), .Z(n4548) );
  CNIVX1 U3736 ( .A(n3826), .Z(n4549) );
  CNIVX1 U3737 ( .A(n4551), .Z(n4550) );
  CNIVX1 U3738 ( .A(n3827), .Z(n4551) );
  CNIVX1 U3739 ( .A(n4553), .Z(n4552) );
  CNIVX1 U3740 ( .A(n3828), .Z(n4553) );
  CNIVX1 U3741 ( .A(n4555), .Z(n4554) );
  CNIVX1 U3742 ( .A(n3829), .Z(n4555) );
  CNIVX1 U3743 ( .A(n4557), .Z(n4556) );
  CNIVX1 U3744 ( .A(n3922), .Z(n4557) );
  CNIVX1 U3745 ( .A(n4559), .Z(n4558) );
  CNIVX1 U3746 ( .A(n3923), .Z(n4559) );
  CNIVX1 U3747 ( .A(n4561), .Z(n4560) );
  CNIVX1 U3748 ( .A(n3924), .Z(n4561) );
  CNIVX1 U3749 ( .A(n4563), .Z(n4562) );
  CNIVX1 U3750 ( .A(n3925), .Z(n4563) );
  CNIVX1 U3751 ( .A(n4565), .Z(n4564) );
  CNIVX1 U3752 ( .A(n3954), .Z(n4565) );
  CNIVX1 U3753 ( .A(n4567), .Z(n4566) );
  CNIVX1 U3754 ( .A(n3955), .Z(n4567) );
  CNIVX1 U3755 ( .A(n4569), .Z(n4568) );
  CNIVX1 U3756 ( .A(n3956), .Z(n4569) );
  CNIVX1 U3757 ( .A(n4571), .Z(n4570) );
  CNIVX1 U3758 ( .A(n3957), .Z(n4571) );
  CNIVX1 U3759 ( .A(n4573), .Z(n4572) );
  CNIVX1 U3760 ( .A(n3856), .Z(n4573) );
  CNIVX1 U3761 ( .A(n4575), .Z(n4574) );
  CNIVX1 U3762 ( .A(n3857), .Z(n4575) );
  CNIVX1 U3763 ( .A(n4577), .Z(n4576) );
  CNIVX1 U3764 ( .A(n3884), .Z(n4577) );
  CNIVX1 U3765 ( .A(n4579), .Z(n4578) );
  CNIVX1 U3766 ( .A(n3885), .Z(n4579) );
  CNIVX1 U3767 ( .A(n4581), .Z(n4580) );
  CNIVX1 U3768 ( .A(n3888), .Z(n4581) );
  CNIVX1 U3769 ( .A(n4583), .Z(n4582) );
  CNIVX1 U3770 ( .A(n3889), .Z(n4583) );
  CNIVX1 U3771 ( .A(n4585), .Z(n4584) );
  CNIVX1 U3772 ( .A(n3858), .Z(n4585) );
  CNIVX1 U3773 ( .A(n4587), .Z(n4586) );
  CNIVX1 U3774 ( .A(n3859), .Z(n4587) );
  CNIVX1 U3775 ( .A(n4589), .Z(n4588) );
  CNIVX1 U3776 ( .A(n3860), .Z(n4589) );
  CNIVX1 U3777 ( .A(n4591), .Z(n4590) );
  CNIVX1 U3778 ( .A(n3861), .Z(n4591) );
  CNIVX1 U3779 ( .A(n4593), .Z(n4592) );
  CNIVX1 U3780 ( .A(n3890), .Z(n4593) );
  CNIVX1 U3781 ( .A(n4595), .Z(n4594) );
  CNIVX1 U3782 ( .A(n3891), .Z(n4595) );
  CNIVX1 U3783 ( .A(n4597), .Z(n4596) );
  CNIVX1 U3784 ( .A(n3892), .Z(n4597) );
  CNIVX1 U3785 ( .A(n4599), .Z(n4598) );
  CNIVX1 U3786 ( .A(n3893), .Z(n4599) );
  CNIVX1 U3787 ( .A(n4601), .Z(n4600) );
  CNIVX1 U3788 ( .A(n3648), .Z(n4601) );
  CNIVX1 U3789 ( .A(n4603), .Z(n4602) );
  CNIVX1 U3790 ( .A(n3649), .Z(n4603) );
  CNIVX1 U3791 ( .A(n4605), .Z(n4604) );
  CNIVX1 U3792 ( .A(n3650), .Z(n4605) );
  CNIVX1 U3793 ( .A(n4607), .Z(n4606) );
  CNIVX1 U3794 ( .A(n3651), .Z(n4607) );
  CNIVX1 U3795 ( .A(n4609), .Z(n4608) );
  CNIVX1 U3796 ( .A(n3652), .Z(n4609) );
  CNIVX1 U3797 ( .A(n4611), .Z(n4610) );
  CNIVX1 U3798 ( .A(n3653), .Z(n4611) );
  CNIVX1 U3799 ( .A(n4613), .Z(n4612) );
  CNIVX1 U3800 ( .A(n3654), .Z(n4613) );
  CNIVX1 U3801 ( .A(n4615), .Z(n4614) );
  CNIVX1 U3802 ( .A(n3655), .Z(n4615) );
  CNIVX1 U3803 ( .A(n4617), .Z(n4616) );
  CNIVX1 U3804 ( .A(n3656), .Z(n4617) );
  CNIVX1 U3805 ( .A(n4619), .Z(n4618) );
  CNIVX1 U3806 ( .A(n3657), .Z(n4619) );
  CNIVX1 U3807 ( .A(n4621), .Z(n4620) );
  CNIVX1 U3808 ( .A(n3658), .Z(n4621) );
  CNIVX1 U3809 ( .A(n4623), .Z(n4622) );
  CNIVX1 U3810 ( .A(n3659), .Z(n4623) );
  CNIVX1 U3811 ( .A(n4625), .Z(n4624) );
  CNIVX1 U3812 ( .A(n3662), .Z(n4625) );
  CNIVX1 U3813 ( .A(n4627), .Z(n4626) );
  CNIVX1 U3814 ( .A(n3663), .Z(n4627) );
  CNIVX1 U3815 ( .A(n4629), .Z(n4628) );
  CNIVX1 U3816 ( .A(n3670), .Z(n4629) );
  CNIVX1 U3817 ( .A(n4631), .Z(n4630) );
  CNIVX1 U3818 ( .A(n3671), .Z(n4631) );
  CNIVX1 U3819 ( .A(n4633), .Z(n4632) );
  CNIVX1 U3820 ( .A(n3672), .Z(n4633) );
  CNIVX1 U3821 ( .A(n4635), .Z(n4634) );
  CNIVX1 U3822 ( .A(n3673), .Z(n4635) );
  CNIVX1 U3823 ( .A(n4637), .Z(n4636) );
  CNIVX1 U3824 ( .A(n3674), .Z(n4637) );
  CNIVX1 U3825 ( .A(n4639), .Z(n4638) );
  CNIVX1 U3826 ( .A(n3675), .Z(n4639) );
  CNIVX1 U3827 ( .A(n4641), .Z(n4640) );
  CNIVX1 U3828 ( .A(n3676), .Z(n4641) );
  CNIVX1 U3829 ( .A(n4643), .Z(n4642) );
  CNIVX1 U3830 ( .A(n3677), .Z(n4643) );
  CNIVX1 U3831 ( .A(n4645), .Z(n4644) );
  CNIVX1 U3832 ( .A(n3678), .Z(n4645) );
  CNIVX1 U3833 ( .A(n4647), .Z(n4646) );
  CNIVX1 U3834 ( .A(n3679), .Z(n4647) );
  CNIVX1 U3835 ( .A(n4649), .Z(n4648) );
  CNIVX1 U3836 ( .A(n3660), .Z(n4649) );
  CNIVX1 U3837 ( .A(n4651), .Z(n4650) );
  CNIVX1 U3838 ( .A(n3661), .Z(n4651) );
  CNIVX1 U3839 ( .A(n4653), .Z(n4652) );
  CNIVX1 U3840 ( .A(n3207), .Z(n4653) );
  CNIVX1 U3841 ( .A(n4655), .Z(n4654) );
  CNIVX1 U3842 ( .A(n3664), .Z(n4655) );
  CNIVX1 U3843 ( .A(n4657), .Z(n4656) );
  CNIVX1 U3844 ( .A(n3665), .Z(n4657) );
  CNIVX1 U3845 ( .A(n4659), .Z(n4658) );
  CNIVX1 U3846 ( .A(n3666), .Z(n4659) );
  CNIVX1 U3847 ( .A(n4661), .Z(n4660) );
  CNIVX1 U3848 ( .A(n3667), .Z(n4661) );
  CNIVX1 U3849 ( .A(n4663), .Z(n4662) );
  CNIVX1 U3850 ( .A(n3668), .Z(n4663) );
  CNIVX1 U3851 ( .A(n4665), .Z(n4664) );
  CNIVX1 U3852 ( .A(n3669), .Z(n4665) );
  CNIVX1 U3853 ( .A(n4667), .Z(n4666) );
  CNIVX1 U3854 ( .A(n3616), .Z(n4667) );
  CNIVX1 U3855 ( .A(n4669), .Z(n4668) );
  CNIVX1 U3856 ( .A(n3617), .Z(n4669) );
  CNIVX1 U3857 ( .A(n4671), .Z(n4670) );
  CNIVX1 U3858 ( .A(n3618), .Z(n4671) );
  CNIVX1 U3859 ( .A(n4673), .Z(n4672) );
  CNIVX1 U3860 ( .A(n3378), .Z(n4673) );
  CNIVX1 U3861 ( .A(n4675), .Z(n4674) );
  CNIVX1 U3862 ( .A(n3379), .Z(n4675) );
  CNIVX1 U3863 ( .A(n4677), .Z(n4676) );
  CNIVX1 U3864 ( .A(n3619), .Z(n4677) );
  CNIVX1 U3865 ( .A(n4679), .Z(n4678) );
  CNIVX1 U3866 ( .A(n3620), .Z(n4679) );
  CNIVX1 U3867 ( .A(n4681), .Z(n4680) );
  CNIVX1 U3868 ( .A(n3621), .Z(n4681) );
  CNIVX1 U3869 ( .A(n4683), .Z(n4682) );
  CNIVX1 U3870 ( .A(n3622), .Z(n4683) );
  CNIVX1 U3871 ( .A(n4685), .Z(n4684) );
  CNIVX1 U3872 ( .A(n3623), .Z(n4685) );
  CNIVX1 U3873 ( .A(n4687), .Z(n4686) );
  CNIVX1 U3874 ( .A(n3624), .Z(n4687) );
  CNIVX1 U3875 ( .A(n4689), .Z(n4688) );
  CNIVX1 U3876 ( .A(n3625), .Z(n4689) );
  CNIVX1 U3877 ( .A(n4691), .Z(n4690) );
  CNIVX1 U3878 ( .A(n3626), .Z(n4691) );
  CNIVX1 U3879 ( .A(n4693), .Z(n4692) );
  CNIVX1 U3880 ( .A(n3627), .Z(n4693) );
  CNIVX1 U3881 ( .A(n4695), .Z(n4694) );
  CNIVX1 U3882 ( .A(n3630), .Z(n4695) );
  CNIVX1 U3883 ( .A(n4697), .Z(n4696) );
  CNIVX1 U3884 ( .A(n3631), .Z(n4697) );
  CNIVX1 U3885 ( .A(n4699), .Z(n4698) );
  CNIVX1 U3886 ( .A(n3638), .Z(n4699) );
  CNIVX1 U3887 ( .A(n4701), .Z(n4700) );
  CNIVX1 U3888 ( .A(n3639), .Z(n4701) );
  CNIVX1 U3889 ( .A(n4703), .Z(n4702) );
  CNIVX1 U3890 ( .A(n3640), .Z(n4703) );
  CNIVX1 U3891 ( .A(n4705), .Z(n4704) );
  CNIVX1 U3892 ( .A(n3641), .Z(n4705) );
  CNIVX1 U3893 ( .A(n4707), .Z(n4706) );
  CNIVX1 U3894 ( .A(n3642), .Z(n4707) );
  CNIVX1 U3895 ( .A(n4709), .Z(n4708) );
  CNIVX1 U3896 ( .A(n3277), .Z(n4709) );
  CNIVX1 U3897 ( .A(n4711), .Z(n4710) );
  CNIVX1 U3898 ( .A(n3202), .Z(n4711) );
  CNIVX1 U3899 ( .A(n4713), .Z(n4712) );
  CNIVX1 U3900 ( .A(n3280), .Z(n4713) );
  CNIVX1 U3901 ( .A(n4715), .Z(n4714) );
  CNIVX1 U3902 ( .A(n3203), .Z(n4715) );
  CNIVX1 U3903 ( .A(n4717), .Z(n4716) );
  CNIVX1 U3904 ( .A(n3281), .Z(n4717) );
  CNIVX1 U3905 ( .A(n4719), .Z(n4718) );
  CNIVX1 U3906 ( .A(n3204), .Z(n4719) );
  CNIVX1 U3907 ( .A(n4721), .Z(n4720) );
  CNIVX1 U3908 ( .A(n3308), .Z(n4721) );
  CNIVX1 U3909 ( .A(n4723), .Z(n4722) );
  CNIVX1 U3910 ( .A(n3205), .Z(n4723) );
  CNIVX1 U3911 ( .A(n4725), .Z(n4724) );
  CNIVX1 U3912 ( .A(n3309), .Z(n4725) );
  CNIVX1 U3913 ( .A(n4727), .Z(n4726) );
  CNIVX1 U3914 ( .A(n3206), .Z(n4727) );
  CNIVX1 U3915 ( .A(n4729), .Z(n4728) );
  CNIVX1 U3916 ( .A(n3312), .Z(n4729) );
  CNIVX1 U3917 ( .A(n4731), .Z(n4730) );
  CNIVX1 U3918 ( .A(n3315), .Z(n4731) );
  CNIVX1 U3919 ( .A(n4733), .Z(n4732) );
  CNIVX1 U3920 ( .A(n3285), .Z(n4733) );
  CNIVX1 U3921 ( .A(n4735), .Z(n4734) );
  CNIVX1 U3922 ( .A(n3276), .Z(n4735) );
  CNIVX1 U3923 ( .A(n4737), .Z(n4736) );
  CNIVX1 U3924 ( .A(n3643), .Z(n4737) );
  CNIVX1 U3925 ( .A(n4739), .Z(n4738) );
  CNIVX1 U3926 ( .A(n3644), .Z(n4739) );
  CNIVX1 U3927 ( .A(n4741), .Z(n4740) );
  CNIVX1 U3928 ( .A(n3645), .Z(n4741) );
  CNIVX1 U3929 ( .A(n4743), .Z(n4742) );
  CNIVX1 U3930 ( .A(n3208), .Z(n4743) );
  CNIVX1 U3931 ( .A(n4745), .Z(n4744) );
  CNIVX1 U3932 ( .A(n3646), .Z(n4745) );
  CNIVX1 U3933 ( .A(n4747), .Z(n4746) );
  CNIVX1 U3934 ( .A(n3647), .Z(n4747) );
  CNIVX1 U3935 ( .A(n4749), .Z(n4748) );
  CNIVX1 U3936 ( .A(n3680), .Z(n4749) );
  CNIVX1 U3937 ( .A(n4751), .Z(n4750) );
  CNIVX1 U3938 ( .A(n3681), .Z(n4751) );
  CNIVX1 U3939 ( .A(n4753), .Z(n4752) );
  CNIVX1 U3940 ( .A(n3682), .Z(n4753) );
  CNIVX1 U3941 ( .A(n4755), .Z(n4754) );
  CNIVX1 U3942 ( .A(n3683), .Z(n4755) );
  CNIVX1 U3943 ( .A(n4757), .Z(n4756) );
  CNIVX1 U3944 ( .A(n3684), .Z(n4757) );
  CNIVX1 U3945 ( .A(n4759), .Z(n4758) );
  CNIVX1 U3946 ( .A(n3209), .Z(n4759) );
  CNIVX1 U3947 ( .A(n4761), .Z(n4760) );
  CNIVX1 U3948 ( .A(n3685), .Z(n4761) );
  CNIVX1 U3949 ( .A(n4763), .Z(n4762) );
  CNIVX1 U3950 ( .A(n3210), .Z(n4763) );
  CNIVX1 U3951 ( .A(n4765), .Z(n4764) );
  CNIVX1 U3952 ( .A(n3686), .Z(n4765) );
  CNIVX1 U3953 ( .A(n4767), .Z(n4766) );
  CNIVX1 U3954 ( .A(n3687), .Z(n4767) );
  CNIVX1 U3955 ( .A(n4769), .Z(n4768) );
  CNIVX1 U3956 ( .A(n3688), .Z(n4769) );
  CNIVX1 U3957 ( .A(n4771), .Z(n4770) );
  CNIVX1 U3958 ( .A(n3689), .Z(n4771) );
  CNIVX1 U3959 ( .A(n4773), .Z(n4772) );
  CNIVX1 U3960 ( .A(n3211), .Z(n4773) );
  CNIVX1 U3961 ( .A(n4775), .Z(n4774) );
  CNIVX1 U3962 ( .A(n3212), .Z(n4775) );
  CNIVX1 U3963 ( .A(n4777), .Z(n4776) );
  CNIVX1 U3964 ( .A(n3690), .Z(n4777) );
  CNIVX1 U3965 ( .A(n4779), .Z(n4778) );
  CNIVX1 U3966 ( .A(n3213), .Z(n4779) );
  CNIVX1 U3967 ( .A(n4781), .Z(n4780) );
  CNIVX1 U3968 ( .A(n3214), .Z(n4781) );
  CNIVX1 U3969 ( .A(n4783), .Z(n4782) );
  CNIVX1 U3970 ( .A(n3691), .Z(n4783) );
  CNIVX1 U3971 ( .A(n4785), .Z(n4784) );
  CNIVX1 U3972 ( .A(n3694), .Z(n4785) );
  CNIVX1 U3973 ( .A(n4787), .Z(n4786) );
  CNIVX1 U3974 ( .A(n3695), .Z(n4787) );
  CNIVX1 U3975 ( .A(n4789), .Z(n4788) );
  CNIVX1 U3976 ( .A(n3702), .Z(n4789) );
  CNIVX1 U3977 ( .A(n4791), .Z(n4790) );
  CNIVX1 U3978 ( .A(n3703), .Z(n4791) );
  CNIVX1 U3979 ( .A(n4793), .Z(n4792) );
  CNIVX1 U3980 ( .A(n3704), .Z(n4793) );
  CNIVX1 U3981 ( .A(n4795), .Z(n4794) );
  CNIVX1 U3982 ( .A(n3705), .Z(n4795) );
  CNIVX1 U3983 ( .A(n4797), .Z(n4796) );
  CNIVX1 U3984 ( .A(n3706), .Z(n4797) );
  CNIVX1 U3985 ( .A(n4799), .Z(n4798) );
  CNIVX1 U3986 ( .A(n3707), .Z(n4799) );
  CNIVX1 U3987 ( .A(n4801), .Z(n4800) );
  CNIVX1 U3988 ( .A(n3215), .Z(n4801) );
  CNIVX1 U3989 ( .A(n4803), .Z(n4802) );
  CNIVX1 U3990 ( .A(n3216), .Z(n4803) );
  CNIVX1 U3991 ( .A(n4805), .Z(n4804) );
  CNIVX1 U3992 ( .A(n3708), .Z(n4805) );
  CNIVX1 U3993 ( .A(n4807), .Z(n4806) );
  CNIVX1 U3994 ( .A(n3217), .Z(n4807) );
  CNIVX1 U3995 ( .A(n4809), .Z(n4808) );
  CNIVX1 U3996 ( .A(n3709), .Z(n4809) );
  CNIVX1 U3997 ( .A(n4811), .Z(n4810) );
  CNIVX1 U3998 ( .A(n3218), .Z(n4811) );
  CNIVX1 U3999 ( .A(n4813), .Z(n4812) );
  CNIVX1 U4000 ( .A(n3219), .Z(n4813) );
  CNIVX1 U4001 ( .A(n4815), .Z(n4814) );
  CNIVX1 U4002 ( .A(n3710), .Z(n4815) );
  CNIVX1 U4003 ( .A(n4817), .Z(n4816) );
  CNIVX1 U4004 ( .A(n3711), .Z(n4817) );
  CNIVX1 U4005 ( .A(n4819), .Z(n4818) );
  CNIVX1 U4006 ( .A(n3628), .Z(n4819) );
  CNIVX1 U4007 ( .A(n4821), .Z(n4820) );
  CNIVX1 U4008 ( .A(n3629), .Z(n4821) );
  CNIVX1 U4009 ( .A(n4823), .Z(n4822) );
  CNIVX1 U4010 ( .A(n3220), .Z(n4823) );
  CNIVX1 U4011 ( .A(n4825), .Z(n4824) );
  CNIVX1 U4012 ( .A(n3632), .Z(n4825) );
  CNIVX1 U4013 ( .A(n4827), .Z(n4826) );
  CNIVX1 U4014 ( .A(n3221), .Z(n4827) );
  CNIVX1 U4015 ( .A(n4829), .Z(n4828) );
  CNIVX1 U4016 ( .A(n3633), .Z(n4829) );
  CNIVX1 U4017 ( .A(n4831), .Z(n4830) );
  CNIVX1 U4018 ( .A(n3692), .Z(n4831) );
  CNIVX1 U4019 ( .A(n4833), .Z(n4832) );
  CNIVX1 U4020 ( .A(n3693), .Z(n4833) );
  CNIVX1 U4021 ( .A(n4835), .Z(n4834) );
  CNIVX1 U4022 ( .A(n3696), .Z(n4835) );
  CNIVX1 U4023 ( .A(n4837), .Z(n4836) );
  CNIVX1 U4024 ( .A(n3697), .Z(n4837) );
  CNIVX1 U4025 ( .A(n4839), .Z(n4838) );
  CNIVX1 U4026 ( .A(n3222), .Z(n4839) );
  CNIVX1 U4027 ( .A(n4841), .Z(n4840) );
  CNIVX1 U4028 ( .A(n3470), .Z(n4841) );
  CNIVX1 U4029 ( .A(n4843), .Z(n4842) );
  CNIVX1 U4030 ( .A(n3223), .Z(n4843) );
  CNIVX1 U4031 ( .A(n4845), .Z(n4844) );
  CNIVX1 U4032 ( .A(n3224), .Z(n4845) );
  CNIVX1 U4033 ( .A(n4847), .Z(n4846) );
  CNIVX1 U4034 ( .A(n3471), .Z(n4847) );
  CNIVX1 U4035 ( .A(n4849), .Z(n4848) );
  CNIVX1 U4036 ( .A(n3478), .Z(n4849) );
  CNIVX1 U4037 ( .A(n4851), .Z(n4850) );
  CNIVX1 U4038 ( .A(n3479), .Z(n4851) );
  CNIVX1 U4039 ( .A(n4853), .Z(n4852) );
  CNIVX1 U4040 ( .A(n3480), .Z(n4853) );
  CNIVX1 U4041 ( .A(n4855), .Z(n4854) );
  CNIVX1 U4042 ( .A(n3225), .Z(n4855) );
  CNIVX1 U4043 ( .A(n4857), .Z(n4856) );
  CNIVX1 U4044 ( .A(n3481), .Z(n4857) );
  CNIVX1 U4045 ( .A(n4859), .Z(n4858) );
  CNIVX1 U4046 ( .A(n3226), .Z(n4859) );
  CNIVX1 U4047 ( .A(n4861), .Z(n4860) );
  CNIVX1 U4048 ( .A(n3482), .Z(n4861) );
  CNIVX1 U4049 ( .A(n4863), .Z(n4862) );
  CNIVX1 U4050 ( .A(n3483), .Z(n4863) );
  CNIVX1 U4051 ( .A(n4865), .Z(n4864) );
  CNIVX1 U4052 ( .A(n3227), .Z(n4865) );
  CNIVX1 U4053 ( .A(n4867), .Z(n4866) );
  CNIVX1 U4054 ( .A(n3228), .Z(n4867) );
  CNIVX1 U4055 ( .A(n4869), .Z(n4868) );
  CNIVX1 U4056 ( .A(n3484), .Z(n4869) );
  CNIVX1 U4057 ( .A(n4871), .Z(n4870) );
  CNIVX1 U4058 ( .A(n3229), .Z(n4871) );
  CNIVX1 U4059 ( .A(n4873), .Z(n4872) );
  CNIVX1 U4060 ( .A(n3485), .Z(n4873) );
  CNIVX1 U4061 ( .A(n4875), .Z(n4874) );
  CNIVX1 U4062 ( .A(n3230), .Z(n4875) );
  CNIVX1 U4063 ( .A(n4877), .Z(n4876) );
  CNIVX1 U4064 ( .A(n3231), .Z(n4877) );
  CNIVX1 U4065 ( .A(n4879), .Z(n4878) );
  CNIVX1 U4066 ( .A(n3486), .Z(n4879) );
  CNIVX1 U4067 ( .A(n4881), .Z(n4880) );
  CNIVX1 U4068 ( .A(n3487), .Z(n4881) );
  CNIVX1 U4069 ( .A(n4883), .Z(n4882) );
  CNIVX1 U4070 ( .A(n3520), .Z(n4883) );
  CNIVX1 U4071 ( .A(n4885), .Z(n4884) );
  CNIVX1 U4072 ( .A(n3521), .Z(n4885) );
  CNIVX1 U4073 ( .A(n4887), .Z(n4886) );
  CNIVX1 U4074 ( .A(n4236), .Z(n4887) );
  CNIVX1 U4075 ( .A(n4889), .Z(n4888) );
  CNIVX1 U4076 ( .A(n3522), .Z(n4889) );
  CNIVX1 U4077 ( .A(n4891), .Z(n4890) );
  CNIVX1 U4078 ( .A(n3264), .Z(n4891) );
  CNIVX1 U4079 ( .A(n4893), .Z(n4892) );
  CNIVX1 U4080 ( .A(n3265), .Z(n4893) );
  CNIVX1 U4081 ( .A(n4895), .Z(n4894) );
  CNIVX1 U4082 ( .A(n3523), .Z(n4895) );
  CNIVX1 U4083 ( .A(n4897), .Z(n4896) );
  CNIVX1 U4084 ( .A(n3524), .Z(n4897) );
  CNIVX1 U4085 ( .A(n4899), .Z(n4898) );
  CNIVX1 U4086 ( .A(n3525), .Z(n4899) );
  CNIVX1 U4087 ( .A(n4901), .Z(n4900) );
  CNIVX1 U4088 ( .A(n3266), .Z(n4901) );
  CNIVX1 U4089 ( .A(n4903), .Z(n4902) );
  CNIVX1 U4090 ( .A(n3267), .Z(n4903) );
  CNIVX1 U4091 ( .A(n4905), .Z(n4904) );
  CNIVX1 U4092 ( .A(n3526), .Z(n4905) );
  CNIVX1 U4093 ( .A(n4907), .Z(n4906) );
  CNIVX1 U4094 ( .A(n3268), .Z(n4907) );
  CNIVX1 U4095 ( .A(n4909), .Z(n4908) );
  CNIVX1 U4096 ( .A(n3269), .Z(n4909) );
  CNIVX1 U4097 ( .A(n4911), .Z(n4910) );
  CNIVX1 U4098 ( .A(n3270), .Z(n4911) );
  CNIVX1 U4099 ( .A(n4913), .Z(n4912) );
  CNIVX1 U4100 ( .A(n3527), .Z(n4913) );
  CNIVX1 U4101 ( .A(n4915), .Z(n4914) );
  CNIVX1 U4102 ( .A(n3528), .Z(n4915) );
  CNIVX1 U4103 ( .A(n4917), .Z(n4916) );
  CNIVX1 U4104 ( .A(n3529), .Z(n4917) );
  CNIVX1 U4105 ( .A(n4919), .Z(n4918) );
  CNIVX1 U4106 ( .A(n3530), .Z(n4919) );
  CNIVX1 U4107 ( .A(n4921), .Z(n4920) );
  CNIVX1 U4108 ( .A(n3531), .Z(n4921) );
  CNIVX1 U4109 ( .A(n4923), .Z(n4922) );
  CNIVX1 U4110 ( .A(n3534), .Z(n4923) );
  CNIVX1 U4111 ( .A(n4925), .Z(n4924) );
  CNIVX1 U4112 ( .A(n3535), .Z(n4925) );
  CNIVX1 U4113 ( .A(n4927), .Z(n4926) );
  CNIVX1 U4114 ( .A(n3542), .Z(n4927) );
  CNIVX1 U4115 ( .A(n4929), .Z(n4928) );
  CNIVX1 U4116 ( .A(n3543), .Z(n4929) );
  CNIVX1 U4117 ( .A(n4931), .Z(n4930) );
  CNIVX1 U4118 ( .A(n3544), .Z(n4931) );
  CNIVX1 U4119 ( .A(n4933), .Z(n4932) );
  CNIVX1 U4120 ( .A(n3545), .Z(n4933) );
  CNIVX1 U4121 ( .A(n4935), .Z(n4934) );
  CNIVX1 U4122 ( .A(n3271), .Z(n4935) );
  CNIVX1 U4123 ( .A(n4937), .Z(n4936) );
  CNIVX1 U4124 ( .A(n3546), .Z(n4937) );
  CNIVX1 U4125 ( .A(n4939), .Z(n4938) );
  CNIVX1 U4126 ( .A(n3547), .Z(n4939) );
  CNIVX1 U4127 ( .A(n4941), .Z(n4940) );
  CNIVX1 U4128 ( .A(n3548), .Z(n4941) );
  CNIVX1 U4129 ( .A(n4943), .Z(n4942) );
  CNIVX1 U4130 ( .A(n3549), .Z(n4943) );
  CNIVX1 U4131 ( .A(n4945), .Z(n4944) );
  CNIVX1 U4132 ( .A(n3550), .Z(n4945) );
  CNIVX1 U4133 ( .A(n4947), .Z(n4946) );
  CNIVX1 U4134 ( .A(n3551), .Z(n4947) );
  CNIVX1 U4135 ( .A(n4949), .Z(n4948) );
  CNIVX1 U4136 ( .A(n3598), .Z(n4949) );
  CNIVX1 U4137 ( .A(n4951), .Z(n4950) );
  CNIVX1 U4138 ( .A(n3272), .Z(n4951) );
  CNIVX1 U4139 ( .A(n4953), .Z(n4952) );
  CNIVX1 U4140 ( .A(n3599), .Z(n4953) );
  CNIVX1 U4141 ( .A(n4955), .Z(n4954) );
  CNIVX1 U4142 ( .A(n3273), .Z(n4955) );
  CNIVX1 U4143 ( .A(n4957), .Z(n4956) );
  CNIVX1 U4144 ( .A(n3606), .Z(n4957) );
  CNIVX1 U4145 ( .A(n4959), .Z(n4958) );
  CNIVX1 U4146 ( .A(n3607), .Z(n4959) );
  CNIVX1 U4147 ( .A(n4961), .Z(n4960) );
  CNIVX1 U4148 ( .A(n3608), .Z(n4961) );
  CNIVX1 U4149 ( .A(n4963), .Z(n4962) );
  CNIVX1 U4150 ( .A(n3609), .Z(n4963) );
  CNIVX1 U4151 ( .A(n4965), .Z(n4964) );
  CNIVX1 U4152 ( .A(n3833), .Z(n4965) );
  CNIVX1 U4153 ( .A(n4967), .Z(n4966) );
  CNIVX1 U4154 ( .A(n3834), .Z(n4967) );
  CNIVX1 U4155 ( .A(n4969), .Z(n4968) );
  CNIVX1 U4156 ( .A(n3835), .Z(n4969) );
  CNIVX1 U4157 ( .A(n4971), .Z(n4970) );
  CNIVX1 U4158 ( .A(n3836), .Z(n4971) );
  CNIVX1 U4159 ( .A(n4973), .Z(n4972) );
  CNIVX1 U4160 ( .A(n3837), .Z(n4973) );
  CNIVX1 U4161 ( .A(n4975), .Z(n4974) );
  CNIVX1 U4162 ( .A(n3838), .Z(n4975) );
  CNIVX1 U4163 ( .A(n4977), .Z(n4976) );
  CNIVX1 U4164 ( .A(n3839), .Z(n4977) );
  CNIVX1 U4165 ( .A(n4979), .Z(n4978) );
  CNIVX1 U4166 ( .A(n3904), .Z(n4979) );
  CNIVX1 U4167 ( .A(n4981), .Z(n4980) );
  CNIVX1 U4168 ( .A(n3905), .Z(n4981) );
  CNIVX1 U4169 ( .A(n4983), .Z(n4982) );
  CNIVX1 U4170 ( .A(n3812), .Z(n4983) );
  CNIVX1 U4171 ( .A(n4985), .Z(n4984) );
  CNIVX1 U4172 ( .A(n3906), .Z(n4985) );
  CNIVX1 U4173 ( .A(n4987), .Z(n4986) );
  CNIVX1 U4174 ( .A(n3907), .Z(n4987) );
  CNIVX1 U4175 ( .A(n4989), .Z(n4988) );
  CNIVX1 U4176 ( .A(n3810), .Z(n4989) );
  CNIVX1 U4177 ( .A(n4991), .Z(n4990) );
  CNIVX1 U4178 ( .A(n3908), .Z(n4991) );
  CNIVX1 U4179 ( .A(n4993), .Z(n4992) );
  CNIVX1 U4180 ( .A(n3610), .Z(n4993) );
  CNIVX1 U4181 ( .A(n4995), .Z(n4994) );
  CNIVX1 U4182 ( .A(n3611), .Z(n4995) );
  CNIVX1 U4183 ( .A(n4997), .Z(n4996) );
  CNIVX1 U4184 ( .A(n3612), .Z(n4997) );
  CNIVX1 U4185 ( .A(n4999), .Z(n4998) );
  CNIVX1 U4186 ( .A(n3613), .Z(n4999) );
  CNIVX1 U4187 ( .A(n5001), .Z(n5000) );
  CNIVX1 U4188 ( .A(n3614), .Z(n5001) );
  CNIVX1 U4189 ( .A(n5003), .Z(n5002) );
  CNIVX1 U4190 ( .A(n3615), .Z(n5003) );
  CNIVX1 U4191 ( .A(n5005), .Z(n5004) );
  CNIVX1 U4192 ( .A(n3634), .Z(n5005) );
  CNIVX1 U4193 ( .A(n5007), .Z(n5006) );
  CNIVX1 U4194 ( .A(n3635), .Z(n5007) );
  CNIVX1 U4195 ( .A(n5009), .Z(n5008) );
  CNIVX1 U4196 ( .A(n3636), .Z(n5009) );
  CNIVX1 U4197 ( .A(n5011), .Z(n5010) );
  CNIVX1 U4198 ( .A(n3637), .Z(n5011) );
  CNIVX1 U4199 ( .A(n5013), .Z(n5012) );
  CNIVX1 U4200 ( .A(n3698), .Z(n5013) );
  CNIVX1 U4201 ( .A(n5015), .Z(n5014) );
  CNIVX1 U4202 ( .A(n3699), .Z(n5015) );
  CNIVX1 U4203 ( .A(n5017), .Z(n5016) );
  CNIVX1 U4204 ( .A(n3700), .Z(n5017) );
  CNIVX1 U4205 ( .A(n5019), .Z(n5018) );
  CNIVX1 U4206 ( .A(n3701), .Z(n5019) );
  CNIVX1 U4207 ( .A(n5021), .Z(n5020) );
  CNIVX1 U4208 ( .A(n3468), .Z(n5021) );
  CNIVX1 U4209 ( .A(n5023), .Z(n5022) );
  CNIVX1 U4210 ( .A(n3472), .Z(n5023) );
  CNIVX1 U4211 ( .A(n5025), .Z(n5024) );
  CNIVX1 U4212 ( .A(n3473), .Z(n5025) );
  CNIVX1 U4213 ( .A(n5027), .Z(n5026) );
  CNIVX1 U4214 ( .A(n3532), .Z(n5027) );
  CNIVX1 U4215 ( .A(n5029), .Z(n5028) );
  CNIVX1 U4216 ( .A(n3533), .Z(n5029) );
  CNIVX1 U4217 ( .A(n5031), .Z(n5030) );
  CNIVX1 U4218 ( .A(n3274), .Z(n5031) );
  CNIVX1 U4219 ( .A(n5033), .Z(n5032) );
  CNIVX1 U4220 ( .A(n3536), .Z(n5033) );
  CNIVX1 U4221 ( .A(n5035), .Z(n5034) );
  CNIVX1 U4222 ( .A(n3275), .Z(n5035) );
  CNIVX1 U4223 ( .A(n5037), .Z(n5036) );
  CNIVX1 U4224 ( .A(n3278), .Z(n5037) );
  CNIVX1 U4225 ( .A(n5039), .Z(n5038) );
  CNIVX1 U4226 ( .A(n3537), .Z(n5039) );
  CNIVX1 U4227 ( .A(n5041), .Z(n5040) );
  CNIVX1 U4228 ( .A(n3600), .Z(n5041) );
  CNIVX1 U4229 ( .A(n5043), .Z(n5042) );
  CNIVX1 U4230 ( .A(n3601), .Z(n5043) );
  CNIVX1 U4231 ( .A(n5045), .Z(n5044) );
  CNIVX1 U4232 ( .A(n3474), .Z(n5045) );
  CNIVX1 U4233 ( .A(n5047), .Z(n5046) );
  CNIVX1 U4234 ( .A(n3475), .Z(n5047) );
  CNIVX1 U4235 ( .A(n5049), .Z(n5048) );
  CNIVX1 U4236 ( .A(n3476), .Z(n5049) );
  CNIVX1 U4237 ( .A(n5051), .Z(n5050) );
  CNIVX1 U4238 ( .A(n3477), .Z(n5051) );
  CNIVX1 U4239 ( .A(n5053), .Z(n5052) );
  CNIVX1 U4240 ( .A(n3538), .Z(n5053) );
  CNIVX1 U4241 ( .A(n5055), .Z(n5054) );
  CNIVX1 U4242 ( .A(n3539), .Z(n5055) );
  CNIVX1 U4243 ( .A(n5057), .Z(n5056) );
  CNIVX1 U4244 ( .A(n3540), .Z(n5057) );
  CNIVX1 U4245 ( .A(n5059), .Z(n5058) );
  CNIVX1 U4246 ( .A(n3541), .Z(n5059) );
  CNIVX1 U4247 ( .A(n5061), .Z(n5060) );
  CNIVX1 U4248 ( .A(n3602), .Z(n5061) );
  CNIVX1 U4249 ( .A(n5063), .Z(n5062) );
  CNIVX1 U4250 ( .A(n3603), .Z(n5063) );
  CNIVX1 U4251 ( .A(n5065), .Z(n5064) );
  CNIVX1 U4252 ( .A(n3604), .Z(n5065) );
  CNIVX1 U4253 ( .A(n5067), .Z(n5066) );
  CNIVX1 U4254 ( .A(n3605), .Z(n5067) );
  CNIVX1 U4255 ( .A(n5069), .Z(n5068) );
  CNIVX1 U4256 ( .A(n3232), .Z(n5069) );
  CNIVX1 U4257 ( .A(n5071), .Z(n5070) );
  CNIVX1 U4258 ( .A(n3233), .Z(n5071) );
  CNIVX1 U4259 ( .A(n5073), .Z(n5072) );
  CNIVX1 U4260 ( .A(n3234), .Z(n5073) );
  CNIVX1 U4261 ( .A(n5075), .Z(n5074) );
  CNIVX1 U4262 ( .A(n3235), .Z(n5075) );
  CNIVX1 U4263 ( .A(n5077), .Z(n5076) );
  CNIVX1 U4264 ( .A(n3236), .Z(n5077) );
  CNIVX1 U4265 ( .A(n5079), .Z(n5078) );
  CNIVX1 U4266 ( .A(n3237), .Z(n5079) );
  CNIVX1 U4267 ( .A(n5081), .Z(n5080) );
  CNIVX1 U4268 ( .A(n3238), .Z(n5081) );
  CNIVX1 U4269 ( .A(n5083), .Z(n5082) );
  CNIVX1 U4270 ( .A(n3239), .Z(n5083) );
  CNIVX1 U4271 ( .A(n5085), .Z(n5084) );
  CNIVX1 U4272 ( .A(n3240), .Z(n5085) );
  CNIVX1 U4273 ( .A(n5087), .Z(n5086) );
  CNIVX1 U4274 ( .A(n3241), .Z(n5087) );
  CNIVX1 U4275 ( .A(n5089), .Z(n5088) );
  CNIVX1 U4276 ( .A(n3242), .Z(n5089) );
  CNIVX1 U4277 ( .A(n5091), .Z(n5090) );
  CNIVX1 U4278 ( .A(n3243), .Z(n5091) );
  CNIVX1 U4279 ( .A(n5093), .Z(n5092) );
  CNIVX1 U4280 ( .A(n3246), .Z(n5093) );
  CNIVX1 U4281 ( .A(n5095), .Z(n5094) );
  CNIVX1 U4282 ( .A(n3279), .Z(n5095) );
  CNIVX1 U4283 ( .A(n5097), .Z(n5096) );
  CNIVX1 U4284 ( .A(n3247), .Z(n5097) );
  CNIVX1 U4285 ( .A(n5099), .Z(n5098) );
  CNIVX1 U4286 ( .A(n3286), .Z(n5099) );
  CNIVX1 U4287 ( .A(n5101), .Z(n5100) );
  CNIVX1 U4288 ( .A(n3287), .Z(n5101) );
  CNIVX1 U4289 ( .A(n5103), .Z(n5102) );
  CNIVX1 U4290 ( .A(n3254), .Z(n5103) );
  CNIVX1 U4291 ( .A(n5105), .Z(n5104) );
  CNIVX1 U4292 ( .A(n3255), .Z(n5105) );
  CNIVX1 U4293 ( .A(n5107), .Z(n5106) );
  CNIVX1 U4294 ( .A(n3256), .Z(n5107) );
  CNIVX1 U4295 ( .A(n5109), .Z(n5108) );
  CNIVX1 U4296 ( .A(n3257), .Z(n5109) );
  CNIVX1 U4297 ( .A(n5111), .Z(n5110) );
  CNIVX1 U4298 ( .A(n3258), .Z(n5111) );
  CNIVX1 U4299 ( .A(n5113), .Z(n5112) );
  CNIVX1 U4300 ( .A(n3259), .Z(n5113) );
  CNIVX1 U4301 ( .A(n5115), .Z(n5114) );
  CNIVX1 U4302 ( .A(n3260), .Z(n5115) );
  CNIVX1 U4303 ( .A(n5117), .Z(n5116) );
  CNIVX1 U4304 ( .A(n3261), .Z(n5117) );
  CNIVX1 U4305 ( .A(n5119), .Z(n5118) );
  CNIVX1 U4306 ( .A(n3262), .Z(n5119) );
  CNIVX1 U4307 ( .A(n5121), .Z(n5120) );
  CNIVX1 U4308 ( .A(n3288), .Z(n5121) );
  CNIVX1 U4309 ( .A(n5123), .Z(n5122) );
  CNIVX1 U4310 ( .A(n3289), .Z(n5123) );
  CNIVX1 U4311 ( .A(n5125), .Z(n5124) );
  CNIVX1 U4312 ( .A(n3263), .Z(n5125) );
  CNIVX1 U4313 ( .A(n5127), .Z(n5126) );
  CNIVX1 U4314 ( .A(n3244), .Z(n5127) );
  CNIVX1 U4315 ( .A(n5129), .Z(n5128) );
  CNIVX1 U4316 ( .A(n3245), .Z(n5129) );
  CNIVX1 U4317 ( .A(n5131), .Z(n5130) );
  CNIVX1 U4318 ( .A(n3248), .Z(n5131) );
  CNIVX1 U4319 ( .A(n5133), .Z(n5132) );
  CNIVX1 U4320 ( .A(n3249), .Z(n5133) );
  CNIVX1 U4321 ( .A(n5135), .Z(n5134) );
  CNIVX1 U4322 ( .A(n3250), .Z(n5135) );
  CNIVX1 U4323 ( .A(n5137), .Z(n5136) );
  CNIVX1 U4324 ( .A(n3251), .Z(n5137) );
  CNIVX1 U4325 ( .A(n5139), .Z(n5138) );
  CNIVX1 U4326 ( .A(n3252), .Z(n5139) );
  CNIVX1 U4327 ( .A(n5141), .Z(n5140) );
  CNIVX1 U4328 ( .A(n3253), .Z(n5141) );
  CNIVX1 U4329 ( .A(n5143), .Z(n5142) );
  CNIVX1 U4330 ( .A(n3488), .Z(n5143) );
  CNIVX1 U4331 ( .A(n5145), .Z(n5144) );
  CNIVX1 U4332 ( .A(n3489), .Z(n5145) );
  CNIVX1 U4333 ( .A(n5147), .Z(n5146) );
  CNIVX1 U4334 ( .A(n3490), .Z(n5147) );
  CNIVX1 U4335 ( .A(n5149), .Z(n5148) );
  CNIVX1 U4336 ( .A(n3491), .Z(n5149) );
  CNIVX1 U4337 ( .A(n5151), .Z(n5150) );
  CNIVX1 U4338 ( .A(n3492), .Z(n5151) );
  CNIVX1 U4339 ( .A(n5153), .Z(n5152) );
  CNIVX1 U4340 ( .A(n3493), .Z(n5153) );
  CNIVX1 U4341 ( .A(n5155), .Z(n5154) );
  CNIVX1 U4342 ( .A(n3494), .Z(n5155) );
  CNIVX1 U4343 ( .A(n5157), .Z(n5156) );
  CNIVX1 U4344 ( .A(n3495), .Z(n5157) );
  CNIVX1 U4345 ( .A(n5159), .Z(n5158) );
  CNIVX1 U4346 ( .A(n3290), .Z(n5159) );
  CNIVX1 U4347 ( .A(n5161), .Z(n5160) );
  CNIVX1 U4348 ( .A(n3496), .Z(n5161) );
  CNIVX1 U4349 ( .A(n5163), .Z(n5162) );
  CNIVX1 U4350 ( .A(n3291), .Z(n5163) );
  CNIVX1 U4351 ( .A(n5165), .Z(n5164) );
  CNIVX1 U4352 ( .A(n3292), .Z(n5165) );
  CNIVX1 U4353 ( .A(n5167), .Z(n5166) );
  CNIVX1 U4354 ( .A(n3497), .Z(n5167) );
  CNIVX1 U4355 ( .A(n5169), .Z(n5168) );
  CNIVX1 U4356 ( .A(n3498), .Z(n5169) );
  CNIVX1 U4357 ( .A(n5171), .Z(n5170) );
  CNIVX1 U4358 ( .A(n3499), .Z(n5171) );
  CNIVX1 U4359 ( .A(n5173), .Z(n5172) );
  CNIVX1 U4360 ( .A(n3502), .Z(n5173) );
  CNIVX1 U4361 ( .A(n5175), .Z(n5174) );
  CNIVX1 U4362 ( .A(n3503), .Z(n5175) );
  CNIVX1 U4363 ( .A(n5177), .Z(n5176) );
  CNIVX1 U4364 ( .A(n3510), .Z(n5177) );
  CNIVX1 U4365 ( .A(n5179), .Z(n5178) );
  CNIVX1 U4366 ( .A(n3511), .Z(n5179) );
  CNIVX1 U4367 ( .A(n5181), .Z(n5180) );
  CNIVX1 U4368 ( .A(n3512), .Z(n5181) );
  CNIVX1 U4369 ( .A(n5183), .Z(n5182) );
  CNIVX1 U4370 ( .A(n3513), .Z(n5183) );
  CNIVX1 U4371 ( .A(n5185), .Z(n5184) );
  CNIVX1 U4372 ( .A(n3514), .Z(n5185) );
  CNIVX1 U4373 ( .A(n5187), .Z(n5186) );
  CNIVX1 U4374 ( .A(n3515), .Z(n5187) );
  CNIVX1 U4375 ( .A(n5189), .Z(n5188) );
  CNIVX1 U4376 ( .A(n3516), .Z(n5189) );
  CNIVX1 U4377 ( .A(n5191), .Z(n5190) );
  CNIVX1 U4378 ( .A(n3517), .Z(n5191) );
  CNIVX1 U4379 ( .A(n5193), .Z(n5192) );
  CNIVX1 U4380 ( .A(n3518), .Z(n5193) );
  CNIVX1 U4381 ( .A(n5195), .Z(n5194) );
  CNIVX1 U4382 ( .A(n3519), .Z(n5195) );
  CNIVX1 U4383 ( .A(n5197), .Z(n5196) );
  CNIVX1 U4384 ( .A(n3552), .Z(n5197) );
  CNIVX1 U4385 ( .A(n5199), .Z(n5198) );
  CNIVX1 U4386 ( .A(n3553), .Z(n5199) );
  CNIVX1 U4387 ( .A(n5201), .Z(n5200) );
  CNIVX1 U4388 ( .A(n3554), .Z(n5201) );
  CNIVX1 U4389 ( .A(n5203), .Z(n5202) );
  CNIVX1 U4390 ( .A(n3555), .Z(n5203) );
  CNIVX1 U4391 ( .A(n5205), .Z(n5204) );
  CNIVX1 U4392 ( .A(n3556), .Z(n5205) );
  CNIVX1 U4393 ( .A(n5207), .Z(n5206) );
  CNIVX1 U4394 ( .A(n3557), .Z(n5207) );
  CNIVX1 U4395 ( .A(n5209), .Z(n5208) );
  CNIVX1 U4396 ( .A(n3558), .Z(n5209) );
  CNIVX1 U4397 ( .A(n5211), .Z(n5210) );
  CNIVX1 U4398 ( .A(n3559), .Z(n5211) );
  CNIVX1 U4399 ( .A(n5213), .Z(n5212) );
  CNIVX1 U4400 ( .A(n3560), .Z(n5213) );
  CNIVX1 U4401 ( .A(n5215), .Z(n5214) );
  CNIVX1 U4402 ( .A(n3561), .Z(n5215) );
  CNIVX1 U4403 ( .A(n5217), .Z(n5216) );
  CNIVX1 U4404 ( .A(n3562), .Z(n5217) );
  CNIVX1 U4405 ( .A(n5219), .Z(n5218) );
  CNIVX1 U4406 ( .A(n3563), .Z(n5219) );
  CNIVX1 U4407 ( .A(n5221), .Z(n5220) );
  CNIVX1 U4408 ( .A(n3437), .Z(n5221) );
  CNIVX1 U4409 ( .A(n5223), .Z(n5222) );
  CNIVX1 U4410 ( .A(n3313), .Z(n5223) );
  CNIVX1 U4411 ( .A(n5225), .Z(n5224) );
  CNIVX1 U4412 ( .A(n3440), .Z(n5225) );
  CNIVX1 U4413 ( .A(n5227), .Z(n5226) );
  CNIVX1 U4414 ( .A(n3404), .Z(n5227) );
  CNIVX1 U4415 ( .A(n5229), .Z(n5228) );
  CNIVX1 U4416 ( .A(n3441), .Z(n5229) );
  CNIVX1 U4417 ( .A(n5231), .Z(n5230) );
  CNIVX1 U4418 ( .A(n3405), .Z(n5231) );
  CNIVX1 U4419 ( .A(n5233), .Z(n5232) );
  CNIVX1 U4420 ( .A(n3282), .Z(n5233) );
  CNIVX1 U4421 ( .A(n5235), .Z(n5234) );
  CNIVX1 U4422 ( .A(n3408), .Z(n5235) );
  CNIVX1 U4423 ( .A(n5237), .Z(n5236) );
  CNIVX1 U4424 ( .A(n3283), .Z(n5237) );
  CNIVX1 U4425 ( .A(n5239), .Z(n5238) );
  CNIVX1 U4426 ( .A(n3409), .Z(n5239) );
  CNIVX1 U4427 ( .A(n5241), .Z(n5240) );
  CNIVX1 U4428 ( .A(n3284), .Z(n5241) );
  CNIVX1 U4429 ( .A(n5243), .Z(n5242) );
  CNIVX1 U4430 ( .A(n3316), .Z(n5243) );
  CNIVX1 U4431 ( .A(n5245), .Z(n5244) );
  CNIVX1 U4432 ( .A(n3566), .Z(n5245) );
  CNIVX1 U4433 ( .A(n5247), .Z(n5246) );
  CNIVX1 U4434 ( .A(n3436), .Z(n5247) );
  CNIVX1 U4435 ( .A(n5249), .Z(n5248) );
  CNIVX1 U4436 ( .A(n3377), .Z(n5249) );
  CNIVX1 U4437 ( .A(n5251), .Z(n5250) );
  CNIVX1 U4438 ( .A(n3346), .Z(n5251) );
  CNIVX1 U4439 ( .A(n5253), .Z(n5252) );
  CNIVX1 U4440 ( .A(n3567), .Z(n5253) );
  CNIVX1 U4441 ( .A(n5255), .Z(n5254) );
  CNIVX1 U4442 ( .A(n3574), .Z(n5255) );
  CNIVX1 U4443 ( .A(n5257), .Z(n5256) );
  CNIVX1 U4444 ( .A(n3575), .Z(n5257) );
  CNIVX1 U4445 ( .A(n5259), .Z(n5258) );
  CNIVX1 U4446 ( .A(n3576), .Z(n5259) );
  CNIVX1 U4447 ( .A(n5261), .Z(n5260) );
  CNIVX1 U4448 ( .A(n3577), .Z(n5261) );
  CNIVX1 U4449 ( .A(n5263), .Z(n5262) );
  CNIVX1 U4450 ( .A(n3578), .Z(n5263) );
  CNIVX1 U4451 ( .A(n5265), .Z(n5264) );
  CNIVX1 U4452 ( .A(n3579), .Z(n5265) );
  CNIVX1 U4453 ( .A(n5267), .Z(n5266) );
  CNIVX1 U4454 ( .A(n3580), .Z(n5267) );
  CNIVX1 U4455 ( .A(n5269), .Z(n5268) );
  CNIVX1 U4456 ( .A(n3581), .Z(n5269) );
  CNIVX1 U4457 ( .A(n5271), .Z(n5270) );
  CNIVX1 U4458 ( .A(n3293), .Z(n5271) );
  CNIVX1 U4459 ( .A(n5273), .Z(n5272) );
  CNIVX1 U4460 ( .A(n3582), .Z(n5273) );
  CNIVX1 U4461 ( .A(n5275), .Z(n5274) );
  CNIVX1 U4462 ( .A(n3294), .Z(n5275) );
  CNIVX1 U4463 ( .A(n5277), .Z(n5276) );
  CNIVX1 U4464 ( .A(n3583), .Z(n5277) );
  CNIVX1 U4465 ( .A(n5279), .Z(n5278) );
  CNIVX1 U4466 ( .A(n3500), .Z(n5279) );
  CNIVX1 U4467 ( .A(n5281), .Z(n5280) );
  CNIVX1 U4468 ( .A(n3501), .Z(n5281) );
  CNIVX1 U4469 ( .A(n5283), .Z(n5282) );
  CNIVX1 U4470 ( .A(n3504), .Z(n5283) );
  CNIVX1 U4471 ( .A(n5285), .Z(n5284) );
  CNIVX1 U4472 ( .A(n3505), .Z(n5285) );
  CNIVX1 U4473 ( .A(n5287), .Z(n5286) );
  CNIVX1 U4474 ( .A(n3295), .Z(n5287) );
  CNIVX1 U4475 ( .A(n5289), .Z(n5288) );
  CNIVX1 U4476 ( .A(n3564), .Z(n5289) );
  CNIVX1 U4477 ( .A(n5291), .Z(n5290) );
  CNIVX1 U4478 ( .A(n3296), .Z(n5291) );
  CNIVX1 U4479 ( .A(n5293), .Z(n5292) );
  CNIVX1 U4480 ( .A(n3297), .Z(n5293) );
  CNIVX1 U4481 ( .A(n5295), .Z(n5294) );
  CNIVX1 U4482 ( .A(n3565), .Z(n5295) );
  CNIVX1 U4483 ( .A(n5297), .Z(n5296) );
  CNIVX1 U4484 ( .A(n3568), .Z(n5297) );
  CNIVX1 U4485 ( .A(n5299), .Z(n5298) );
  CNIVX1 U4486 ( .A(n3569), .Z(n5299) );
  CNIVX1 U4487 ( .A(n5301), .Z(n5300) );
  CNIVX1 U4488 ( .A(n3506), .Z(n5301) );
  CNIVX1 U4489 ( .A(n5303), .Z(n5302) );
  CNIVX1 U4490 ( .A(n3507), .Z(n5303) );
  CNIVX1 U4491 ( .A(n5305), .Z(n5304) );
  CNIVX1 U4492 ( .A(n3508), .Z(n5305) );
  CNIVX1 U4493 ( .A(n5307), .Z(n5306) );
  CNIVX1 U4494 ( .A(n3298), .Z(n5307) );
  CNIVX1 U4495 ( .A(n5309), .Z(n5308) );
  CNIVX1 U4496 ( .A(n3509), .Z(n5309) );
  CNIVX1 U4497 ( .A(n5311), .Z(n5310) );
  CNIVX1 U4498 ( .A(n3570), .Z(n5311) );
  CNIVX1 U4499 ( .A(n5313), .Z(n5312) );
  CNIVX1 U4500 ( .A(n3299), .Z(n5313) );
  CNIVX1 U4501 ( .A(n5315), .Z(n5314) );
  CNIVX1 U4502 ( .A(n3300), .Z(n5315) );
  CNIVX1 U4503 ( .A(n5317), .Z(n5316) );
  CNIVX1 U4504 ( .A(n3571), .Z(n5317) );
  CNIVX1 U4505 ( .A(n5319), .Z(n5318) );
  CNIVX1 U4506 ( .A(n3301), .Z(n5319) );
  CNIVX1 U4507 ( .A(n5321), .Z(n5320) );
  CNIVX1 U4508 ( .A(n3572), .Z(n5321) );
  CNIVX1 U4509 ( .A(n5323), .Z(n5322) );
  CNIVX1 U4510 ( .A(n3302), .Z(n5323) );
  CNIVX1 U4511 ( .A(n5325), .Z(n5324) );
  CNIVX1 U4512 ( .A(n3303), .Z(n5325) );
  CNIVX1 U4513 ( .A(n5327), .Z(n5326) );
  CNIVX1 U4514 ( .A(n3573), .Z(n5327) );
  CNIVX1 U4515 ( .A(n5329), .Z(n5328) );
  CNIVX1 U4516 ( .A(n3726), .Z(n5329) );
  CNIVX1 U4517 ( .A(n5331), .Z(n5330) );
  CNIVX1 U4518 ( .A(n3727), .Z(n5331) );
  CNIVX1 U4519 ( .A(n5333), .Z(n5332) );
  CNIVX1 U4520 ( .A(n3734), .Z(n5333) );
  CNIVX1 U4521 ( .A(n5335), .Z(n5334) );
  CNIVX1 U4522 ( .A(n3304), .Z(n5335) );
  CNIVX1 U4523 ( .A(n5337), .Z(n5336) );
  CNIVX1 U4524 ( .A(n3735), .Z(n5337) );
  CNIVX1 U4525 ( .A(n5339), .Z(n5338) );
  CNIVX1 U4526 ( .A(n3305), .Z(n5339) );
  CNIVX1 U4527 ( .A(n5341), .Z(n5340) );
  CNIVX1 U4528 ( .A(n3736), .Z(n5341) );
  CNIVX1 U4529 ( .A(n5343), .Z(n5342) );
  CNIVX1 U4530 ( .A(n3737), .Z(n5343) );
  CNIVX1 U4531 ( .A(n5345), .Z(n5344) );
  CNIVX1 U4532 ( .A(n3738), .Z(n5345) );
  CNIVX1 U4533 ( .A(n5347), .Z(n5346) );
  CNIVX1 U4534 ( .A(n3739), .Z(n5347) );
  CNIVX1 U4535 ( .A(n5349), .Z(n5348) );
  CNIVX1 U4536 ( .A(n3740), .Z(n5349) );
  CNIVX1 U4537 ( .A(n5351), .Z(n5350) );
  CNIVX1 U4538 ( .A(n3306), .Z(n5351) );
  CNIVX1 U4539 ( .A(n5353), .Z(n5352) );
  CNIVX1 U4540 ( .A(n3741), .Z(n5353) );
  CNIVX1 U4541 ( .A(n5355), .Z(n5354) );
  CNIVX1 U4542 ( .A(n3307), .Z(n5355) );
  CNIVX1 U4543 ( .A(n5357), .Z(n5356) );
  CNIVX1 U4544 ( .A(n3310), .Z(n5357) );
  CNIVX1 U4545 ( .A(n5359), .Z(n5358) );
  CNIVX1 U4546 ( .A(n3742), .Z(n5359) );
  CNIVX1 U4547 ( .A(n5361), .Z(n5360) );
  CNIVX1 U4548 ( .A(n3743), .Z(n5361) );
  CNIVX1 U4549 ( .A(n5363), .Z(n5362) );
  CNIVX1 U4550 ( .A(n3744), .Z(n5363) );
  CNIVX1 U4551 ( .A(n5365), .Z(n5364) );
  CNIVX1 U4552 ( .A(n3745), .Z(n5365) );
  CNIVX1 U4553 ( .A(n5367), .Z(n5366) );
  CNIVX1 U4554 ( .A(n3311), .Z(n5367) );
  CNIVX1 U4555 ( .A(n5369), .Z(n5368) );
  CNIVX1 U4556 ( .A(n3746), .Z(n5369) );
  CNIVX1 U4557 ( .A(n5371), .Z(n5370) );
  CNIVX1 U4558 ( .A(n3318), .Z(n5371) );
  CNIVX1 U4559 ( .A(n5373), .Z(n5372) );
  CNIVX1 U4560 ( .A(n3747), .Z(n5373) );
  CNIVX1 U4561 ( .A(n5375), .Z(n5374) );
  CNIVX1 U4562 ( .A(n3748), .Z(n5375) );
  CNIVX1 U4563 ( .A(n5377), .Z(n5376) );
  CNIVX1 U4564 ( .A(n3319), .Z(n5377) );
  CNIVX1 U4565 ( .A(n5379), .Z(n5378) );
  CNIVX1 U4566 ( .A(n3320), .Z(n5379) );
  CNIVX1 U4567 ( .A(n5381), .Z(n5380) );
  CNIVX1 U4568 ( .A(n3749), .Z(n5381) );
  CNIVX1 U4569 ( .A(n5383), .Z(n5382) );
  CNIVX1 U4570 ( .A(n3321), .Z(n5383) );
  CNIVX1 U4571 ( .A(n5385), .Z(n5384) );
  CNIVX1 U4572 ( .A(n3750), .Z(n5385) );
  CNIVX1 U4573 ( .A(n5387), .Z(n5386) );
  CNIVX1 U4574 ( .A(n3322), .Z(n5387) );
  CNIVX1 U4575 ( .A(n5389), .Z(n5388) );
  CNIVX1 U4576 ( .A(n3323), .Z(n5389) );
  CNIVX1 U4577 ( .A(n5391), .Z(n5390) );
  CNIVX1 U4578 ( .A(n3751), .Z(n5391) );
  CNIVX1 U4579 ( .A(n5393), .Z(n5392) );
  CNIVX1 U4580 ( .A(n3752), .Z(n5393) );
  CNIVX1 U4581 ( .A(n5395), .Z(n5394) );
  CNIVX1 U4582 ( .A(n3753), .Z(n5395) );
  CNIVX1 U4583 ( .A(n5397), .Z(n5396) );
  CNIVX1 U4584 ( .A(n3754), .Z(n5397) );
  CNIVX1 U4585 ( .A(n5399), .Z(n5398) );
  CNIVX1 U4586 ( .A(n3324), .Z(n5399) );
  CNIVX1 U4587 ( .A(n5401), .Z(n5400) );
  CNIVX1 U4588 ( .A(n3755), .Z(n5401) );
  CNIVX1 U4589 ( .A(n5403), .Z(n5402) );
  CNIVX1 U4590 ( .A(n3325), .Z(n5403) );
  CNIVX1 U4591 ( .A(n5405), .Z(n5404) );
  CNIVX1 U4592 ( .A(n3758), .Z(n5405) );
  CNIVX1 U4593 ( .A(n5407), .Z(n5406) );
  CNIVX1 U4594 ( .A(n3759), .Z(n5407) );
  CNIVX1 U4595 ( .A(n5409), .Z(n5408) );
  CNIVX1 U4596 ( .A(n3766), .Z(n5409) );
  CNIVX1 U4597 ( .A(n5411), .Z(n5410) );
  CNIVX1 U4598 ( .A(n3767), .Z(n5411) );
  CNIVX1 U4599 ( .A(n5413), .Z(n5412) );
  CNIVX1 U4600 ( .A(n3326), .Z(n5413) );
  CNIVX1 U4601 ( .A(n5415), .Z(n5414) );
  CNIVX1 U4602 ( .A(n3327), .Z(n5415) );
  CNIVX1 U4603 ( .A(n5417), .Z(n5416) );
  CNIVX1 U4604 ( .A(n3768), .Z(n5417) );
  CNIVX1 U4605 ( .A(n5419), .Z(n5418) );
  CNIVX1 U4606 ( .A(n3392), .Z(n5419) );
  CNIVX1 U4607 ( .A(n5421), .Z(n5420) );
  CNIVX1 U4608 ( .A(n3393), .Z(n5421) );
  CNIVX1 U4609 ( .A(n5423), .Z(n5422) );
  CNIVX1 U4610 ( .A(n3769), .Z(n5423) );
  CNIVX1 U4611 ( .A(n5425), .Z(n5424) );
  CNIVX1 U4612 ( .A(n3770), .Z(n5425) );
  CNIVX1 U4613 ( .A(n5427), .Z(n5426) );
  CNIVX1 U4614 ( .A(n3771), .Z(n5427) );
  CNIVX1 U4615 ( .A(n5429), .Z(n5428) );
  CNIVX1 U4616 ( .A(n3772), .Z(n5429) );
  CNIVX1 U4617 ( .A(n5431), .Z(n5430) );
  CNIVX1 U4618 ( .A(n3773), .Z(n5431) );
  CNIVX1 U4619 ( .A(n5433), .Z(n5432) );
  CNIVX1 U4620 ( .A(n3774), .Z(n5433) );
  CNIVX1 U4621 ( .A(n5435), .Z(n5434) );
  CNIVX1 U4622 ( .A(n3394), .Z(n5435) );
  CNIVX1 U4623 ( .A(n5437), .Z(n5436) );
  CNIVX1 U4624 ( .A(n3775), .Z(n5437) );
  CNIVX1 U4625 ( .A(n3724), .Z(n5438) );
  CNIVX1 U4626 ( .A(n5440), .Z(n5439) );
  CNIVX1 U4627 ( .A(n3728), .Z(n5440) );
  CNIVX1 U4628 ( .A(n5442), .Z(n5441) );
  CNIVX1 U4629 ( .A(n3729), .Z(n5442) );
  CNIVX1 U4630 ( .A(n5444), .Z(n5443) );
  CNIVX1 U4631 ( .A(n3756), .Z(n5444) );
  CNIVX1 U4632 ( .A(n5446), .Z(n5445) );
  CNIVX1 U4633 ( .A(n3757), .Z(n5446) );
  CNIVX1 U4634 ( .A(n5448), .Z(n5447) );
  CNIVX1 U4635 ( .A(n3760), .Z(n5448) );
  CNIVX1 U4636 ( .A(n5450), .Z(n5449) );
  CNIVX1 U4637 ( .A(n3761), .Z(n5450) );
  CNIVX1 U4638 ( .A(n5452), .Z(n5451) );
  CNIVX1 U4639 ( .A(n3730), .Z(n5452) );
  CNIVX1 U4640 ( .A(n5454), .Z(n5453) );
  CNIVX1 U4641 ( .A(n3731), .Z(n5454) );
  CNIVX1 U4642 ( .A(n5456), .Z(n5455) );
  CNIVX1 U4643 ( .A(n3732), .Z(n5456) );
  CNIVX1 U4644 ( .A(n5458), .Z(n5457) );
  CNIVX1 U4645 ( .A(n3733), .Z(n5458) );
  CNIVX1 U4646 ( .A(n5460), .Z(n5459) );
  CNIVX1 U4647 ( .A(n3762), .Z(n5460) );
  CNIVX1 U4648 ( .A(n5462), .Z(n5461) );
  CNIVX1 U4649 ( .A(n3395), .Z(n5462) );
  CNIVX1 U4650 ( .A(n5464), .Z(n5463) );
  CNIVX1 U4651 ( .A(n3763), .Z(n5464) );
  CNIVX1 U4652 ( .A(n5466), .Z(n5465) );
  CNIVX1 U4653 ( .A(n3396), .Z(n5466) );
  CNIVX1 U4654 ( .A(n5468), .Z(n5467) );
  CNIVX1 U4655 ( .A(n3764), .Z(n5468) );
  CNIVX1 U4656 ( .A(n5470), .Z(n5469) );
  CNIVX1 U4657 ( .A(n3765), .Z(n5470) );
  CNIVX1 U4658 ( .A(n5472), .Z(n5471) );
  CNIVX1 U4659 ( .A(n3982), .Z(n5472) );
  CNIVX1 U4660 ( .A(n5474), .Z(n5473) );
  CNIVX1 U4661 ( .A(n3983), .Z(n5474) );
  CNIVX1 U4662 ( .A(n5476), .Z(n5475) );
  CNIVX1 U4663 ( .A(n3990), .Z(n5476) );
  CNIVX1 U4664 ( .A(n5478), .Z(n5477) );
  CNIVX1 U4665 ( .A(n3991), .Z(n5478) );
  CNIVX1 U4666 ( .A(n5480), .Z(n5479) );
  CNIVX1 U4667 ( .A(n3992), .Z(n5480) );
  CNIVX1 U4668 ( .A(n5482), .Z(n5481) );
  CNIVX1 U4669 ( .A(n3993), .Z(n5482) );
  CNIVX1 U4670 ( .A(n5484), .Z(n5483) );
  CNIVX1 U4671 ( .A(n3994), .Z(n5484) );
  CNIVX1 U4672 ( .A(n5486), .Z(n5485) );
  CNIVX1 U4673 ( .A(n3995), .Z(n5486) );
  CNIVX1 U4674 ( .A(n5488), .Z(n5487) );
  CNIVX1 U4675 ( .A(n3996), .Z(n5488) );
  CNIVX1 U4676 ( .A(n5490), .Z(n5489) );
  CNIVX1 U4677 ( .A(n3997), .Z(n5490) );
  CNIVX1 U4678 ( .A(n5492), .Z(n5491) );
  CNIVX1 U4679 ( .A(n3998), .Z(n5492) );
  CNIVX1 U4680 ( .A(n5494), .Z(n5493) );
  CNIVX1 U4681 ( .A(n3999), .Z(n5494) );
  CNIVX1 U4682 ( .A(n5496), .Z(n5495) );
  CNIVX1 U4683 ( .A(n4032), .Z(n5496) );
  CNIVX1 U4684 ( .A(n5498), .Z(n5497) );
  CNIVX1 U4685 ( .A(n3397), .Z(n5498) );
  CNIVX1 U4686 ( .A(n5500), .Z(n5499) );
  CNIVX1 U4687 ( .A(n4033), .Z(n5500) );
  CNIVX1 U4688 ( .A(n5502), .Z(n5501) );
  CNIVX1 U4689 ( .A(n4034), .Z(n5502) );
  CNIVX1 U4690 ( .A(n5504), .Z(n5503) );
  CNIVX1 U4691 ( .A(n4035), .Z(n5504) );
  CNIVX1 U4692 ( .A(n5506), .Z(n5505) );
  CNIVX1 U4693 ( .A(n4036), .Z(n5506) );
  CNIVX1 U4694 ( .A(n5508), .Z(n5507) );
  CNIVX1 U4695 ( .A(n4037), .Z(n5508) );
  CNIVX1 U4696 ( .A(n5510), .Z(n5509) );
  CNIVX1 U4697 ( .A(n3398), .Z(n5510) );
  CNIVX1 U4698 ( .A(n5512), .Z(n5511) );
  CNIVX1 U4699 ( .A(n4038), .Z(n5512) );
  CNIVX1 U4700 ( .A(n5514), .Z(n5513) );
  CNIVX1 U4701 ( .A(n4039), .Z(n5514) );
  CNIVX1 U4702 ( .A(n5516), .Z(n5515) );
  CNIVX1 U4703 ( .A(n3399), .Z(n5516) );
  CNIVX1 U4704 ( .A(n5518), .Z(n5517) );
  CNIVX1 U4705 ( .A(n4040), .Z(n5518) );
  CNIVX1 U4706 ( .A(n5520), .Z(n5519) );
  CNIVX1 U4707 ( .A(n4041), .Z(n5520) );
  CNIVX1 U4708 ( .A(n5522), .Z(n5521) );
  CNIVX1 U4709 ( .A(n4042), .Z(n5522) );
  CNIVX1 U4710 ( .A(n5524), .Z(n5523) );
  CNIVX1 U4711 ( .A(n4043), .Z(n5524) );
  CNIVX1 U4712 ( .A(n4046), .Z(n5525) );
  CNIVX1 U4713 ( .A(n5527), .Z(n5526) );
  CNIVX1 U4714 ( .A(n4047), .Z(n5527) );
  CNIVX1 U4715 ( .A(n5529), .Z(n5528) );
  CNIVX1 U4716 ( .A(n4054), .Z(n5529) );
  CNIVX1 U4717 ( .A(n5531), .Z(n5530) );
  CNIVX1 U4718 ( .A(n4055), .Z(n5531) );
  CNIVX1 U4719 ( .A(n5533), .Z(n5532) );
  CNIVX1 U4720 ( .A(n4056), .Z(n5533) );
  CNIVX1 U4721 ( .A(n5535), .Z(n5534) );
  CNIVX1 U4722 ( .A(n3400), .Z(n5535) );
  CNIVX1 U4723 ( .A(n5537), .Z(n5536) );
  CNIVX1 U4724 ( .A(n3401), .Z(n5537) );
  CNIVX1 U4725 ( .A(n5539), .Z(n5538) );
  CNIVX1 U4726 ( .A(n4057), .Z(n5539) );
  CNIVX1 U4727 ( .A(n5541), .Z(n5540) );
  CNIVX1 U4728 ( .A(n4058), .Z(n5541) );
  CNIVX1 U4729 ( .A(n5543), .Z(n5542) );
  CNIVX1 U4730 ( .A(n4059), .Z(n5543) );
  CNIVX1 U4731 ( .A(n5545), .Z(n5544) );
  CNIVX1 U4732 ( .A(n4060), .Z(n5545) );
  CNIVX1 U4733 ( .A(n5547), .Z(n5546) );
  CNIVX1 U4734 ( .A(n4061), .Z(n5547) );
  CNIVX1 U4735 ( .A(n5549), .Z(n5548) );
  CNIVX1 U4736 ( .A(n4062), .Z(n5549) );
  CNIVX1 U4737 ( .A(n5551), .Z(n5550) );
  CNIVX1 U4738 ( .A(n4063), .Z(n5551) );
  CNIVX1 U4739 ( .A(n5553), .Z(n5552) );
  CNIVX1 U4740 ( .A(n4110), .Z(n5553) );
  CNIVX1 U4741 ( .A(n5555), .Z(n5554) );
  CNIVX1 U4742 ( .A(n4111), .Z(n5555) );
  CNIVX1 U4743 ( .A(n5557), .Z(n5556) );
  CNIVX1 U4744 ( .A(n4118), .Z(n5557) );
  CNIVX1 U4745 ( .A(n5559), .Z(n5558) );
  CNIVX1 U4746 ( .A(n4119), .Z(n5559) );
  CNIVX1 U4747 ( .A(n5561), .Z(n5560) );
  CNIVX1 U4748 ( .A(n4120), .Z(n5561) );
  CNIVX1 U4749 ( .A(n5563), .Z(n5562) );
  CNIVX1 U4750 ( .A(n4121), .Z(n5563) );
  CNIVX1 U4751 ( .A(n5565), .Z(n5564) );
  CNIVX1 U4752 ( .A(n4122), .Z(n5565) );
  CNIVX1 U4753 ( .A(n5567), .Z(n5566) );
  CNIVX1 U4754 ( .A(n4123), .Z(n5567) );
  CNIVX1 U4755 ( .A(n5569), .Z(n5568) );
  CNIVX1 U4756 ( .A(n4124), .Z(n5569) );
  CNIVX1 U4757 ( .A(n5571), .Z(n5570) );
  CNIVX1 U4758 ( .A(n4125), .Z(n5571) );
  CNIVX1 U4759 ( .A(n5573), .Z(n5572) );
  CNIVX1 U4760 ( .A(n3402), .Z(n5573) );
  CNIVX1 U4761 ( .A(n5575), .Z(n5574) );
  CNIVX1 U4762 ( .A(n4126), .Z(n5575) );
  CNIVX1 U4763 ( .A(n5577), .Z(n5576) );
  CNIVX1 U4764 ( .A(n3403), .Z(n5577) );
  CNIVX1 U4765 ( .A(n5579), .Z(n5578) );
  CNIVX1 U4766 ( .A(n3406), .Z(n5579) );
  CNIVX1 U4767 ( .A(n5581), .Z(n5580) );
  CNIVX1 U4768 ( .A(n4127), .Z(n5581) );
  CNIVX1 U4769 ( .A(n5583), .Z(n5582) );
  CNIVX1 U4770 ( .A(n4160), .Z(n5583) );
  CNIVX1 U4771 ( .A(n5585), .Z(n5584) );
  CNIVX1 U4772 ( .A(n4161), .Z(n5585) );
  CNIVX1 U4773 ( .A(n5587), .Z(n5586) );
  CNIVX1 U4774 ( .A(n4162), .Z(n5587) );
  CNIVX1 U4775 ( .A(n5589), .Z(n5588) );
  CNIVX1 U4776 ( .A(n3407), .Z(n5589) );
  CNIVX1 U4777 ( .A(n5591), .Z(n5590) );
  CNIVX1 U4778 ( .A(n4163), .Z(n5591) );
  CNIVX1 U4779 ( .A(n5593), .Z(n5592) );
  CNIVX1 U4780 ( .A(n4164), .Z(n5593) );
  CNIVX1 U4781 ( .A(n5595), .Z(n5594) );
  CNIVX1 U4782 ( .A(n4165), .Z(n5595) );
  CNIVX1 U4783 ( .A(n5597), .Z(n5596) );
  CNIVX1 U4784 ( .A(n4166), .Z(n5597) );
  CNIVX1 U4785 ( .A(n5599), .Z(n5598) );
  CNIVX1 U4786 ( .A(n3414), .Z(n5599) );
  CNIVX1 U4787 ( .A(n5601), .Z(n5600) );
  CNIVX1 U4788 ( .A(n3415), .Z(n5601) );
  CNIVX1 U4789 ( .A(n5603), .Z(n5602) );
  CNIVX1 U4790 ( .A(n4167), .Z(n5603) );
  CNIVX1 U4791 ( .A(n5605), .Z(n5604) );
  CNIVX1 U4792 ( .A(n4168), .Z(n5605) );
  CNIVX1 U4793 ( .A(n5607), .Z(n5606) );
  CNIVX1 U4794 ( .A(n4169), .Z(n5607) );
  CNIVX1 U4795 ( .A(n5609), .Z(n5608) );
  CNIVX1 U4796 ( .A(n4170), .Z(n5609) );
  CNIVX1 U4797 ( .A(n5611), .Z(n5610) );
  CNIVX1 U4798 ( .A(n4171), .Z(n5611) );
  CNIVX1 U4799 ( .A(n5613), .Z(n5612) );
  CNIVX1 U4800 ( .A(n4174), .Z(n5613) );
  CNIVX1 U4801 ( .A(n5615), .Z(n5614) );
  CNIVX1 U4802 ( .A(n4175), .Z(n5615) );
  CNIVX1 U4803 ( .A(n5617), .Z(n5616) );
  CNIVX1 U4804 ( .A(n4182), .Z(n5617) );
  CNIVX1 U4805 ( .A(n5619), .Z(n5618) );
  CNIVX1 U4806 ( .A(n4183), .Z(n5619) );
  CNIVX1 U4807 ( .A(n5621), .Z(n5620) );
  CNIVX1 U4808 ( .A(n4184), .Z(n5621) );
  CNIVX1 U4809 ( .A(n5623), .Z(n5622) );
  CNIVX1 U4810 ( .A(n4185), .Z(n5623) );
  CNIVX1 U4811 ( .A(n5625), .Z(n5624) );
  CNIVX1 U4812 ( .A(n3416), .Z(n5625) );
  CNIVX1 U4813 ( .A(n5627), .Z(n5626) );
  CNIVX1 U4814 ( .A(n4186), .Z(n5627) );
  CNIVX1 U4815 ( .A(n5629), .Z(n5628) );
  CNIVX1 U4816 ( .A(n4187), .Z(n5629) );
  CNIVX1 U4817 ( .A(n5631), .Z(n5630) );
  CNIVX1 U4818 ( .A(n4188), .Z(n5631) );
  CNIVX1 U4819 ( .A(n5633), .Z(n5632) );
  CNIVX1 U4820 ( .A(n4189), .Z(n5633) );
  CNIVX1 U4821 ( .A(n5635), .Z(n5634) );
  CNIVX1 U4822 ( .A(n4190), .Z(n5635) );
  CNIVX1 U4823 ( .A(n5637), .Z(n5636) );
  CNIVX1 U4824 ( .A(n3417), .Z(n5637) );
  CNIVX1 U4825 ( .A(n5639), .Z(n5638) );
  CNIVX1 U4826 ( .A(n4191), .Z(n5639) );
  CNIVX1 U4827 ( .A(n5641), .Z(n5640) );
  CNIVX1 U4828 ( .A(n4000), .Z(n5641) );
  CNIVX1 U4829 ( .A(n5643), .Z(n5642) );
  CNIVX1 U4830 ( .A(n3418), .Z(n5643) );
  CNIVX1 U4831 ( .A(n5645), .Z(n5644) );
  CNIVX1 U4832 ( .A(n4001), .Z(n5645) );
  CNIVX1 U4833 ( .A(n5647), .Z(n5646) );
  CNIVX1 U4834 ( .A(n4002), .Z(n5647) );
  CNIVX1 U4835 ( .A(n5649), .Z(n5648) );
  CNIVX1 U4836 ( .A(n4003), .Z(n5649) );
  CNIVX1 U4837 ( .A(n5651), .Z(n5650) );
  CNIVX1 U4838 ( .A(n4004), .Z(n5651) );
  CNIVX1 U4839 ( .A(n5653), .Z(n5652) );
  CNIVX1 U4840 ( .A(n4005), .Z(n5653) );
  CNIVX1 U4841 ( .A(n5655), .Z(n5654) );
  CNIVX1 U4842 ( .A(n4006), .Z(n5655) );
  CNIVX1 U4843 ( .A(n5657), .Z(n5656) );
  CNIVX1 U4844 ( .A(n4007), .Z(n5657) );
  CNIVX1 U4845 ( .A(n5659), .Z(n5658) );
  CNIVX1 U4846 ( .A(n4008), .Z(n5659) );
  CNIVX1 U4847 ( .A(n5661), .Z(n5660) );
  CNIVX1 U4848 ( .A(n4009), .Z(n5661) );
  CNIVX1 U4849 ( .A(n5663), .Z(n5662) );
  CNIVX1 U4850 ( .A(n4010), .Z(n5663) );
  CNIVX1 U4851 ( .A(n5665), .Z(n5664) );
  CNIVX1 U4852 ( .A(n4011), .Z(n5665) );
  CNIVX1 U4853 ( .A(n5667), .Z(n5666) );
  CNIVX1 U4854 ( .A(n4014), .Z(n5667) );
  CNIVX1 U4855 ( .A(n5669), .Z(n5668) );
  CNIVX1 U4856 ( .A(n4015), .Z(n5669) );
  CNIVX1 U4857 ( .A(n5671), .Z(n5670) );
  CNIVX1 U4858 ( .A(n4022), .Z(n5671) );
  CNIVX1 U4859 ( .A(n5673), .Z(n5672) );
  CNIVX1 U4860 ( .A(n4023), .Z(n5673) );
  CNIVX1 U4861 ( .A(n5675), .Z(n5674) );
  CNIVX1 U4862 ( .A(n4024), .Z(n5675) );
  CNIVX1 U4863 ( .A(n5677), .Z(n5676) );
  CNIVX1 U4864 ( .A(n4025), .Z(n5677) );
  CNIVX1 U4865 ( .A(n5679), .Z(n5678) );
  CNIVX1 U4866 ( .A(n4026), .Z(n5679) );
  CNIVX1 U4867 ( .A(n5681), .Z(n5680) );
  CNIVX1 U4868 ( .A(n4027), .Z(n5681) );
  CNIVX1 U4869 ( .A(n5683), .Z(n5682) );
  CNIVX1 U4870 ( .A(n4028), .Z(n5683) );
  CNIVX1 U4871 ( .A(n5685), .Z(n5684) );
  CNIVX1 U4872 ( .A(n4029), .Z(n5685) );
  CNIVX1 U4873 ( .A(n5687), .Z(n5686) );
  CNIVX1 U4874 ( .A(n4030), .Z(n5687) );
  CNIVX1 U4875 ( .A(n5689), .Z(n5688) );
  CNIVX1 U4876 ( .A(n4031), .Z(n5689) );
  CNIVX1 U4877 ( .A(n5691), .Z(n5690) );
  CNIVX1 U4878 ( .A(n4064), .Z(n5691) );
  CNIVX1 U4879 ( .A(n5693), .Z(n5692) );
  CNIVX1 U4880 ( .A(n4065), .Z(n5693) );
  CNIVX1 U4881 ( .A(n5695), .Z(n5694) );
  CNIVX1 U4882 ( .A(n4066), .Z(n5695) );
  CNIVX1 U4883 ( .A(n5697), .Z(n5696) );
  CNIVX1 U4884 ( .A(n4067), .Z(n5697) );
  CNIVX1 U4885 ( .A(n5699), .Z(n5698) );
  CNIVX1 U4886 ( .A(n3383), .Z(n5699) );
  CNIVX1 U4887 ( .A(n5701), .Z(n5700) );
  CNIVX1 U4888 ( .A(n3317), .Z(n5701) );
  CNIVX1 U4889 ( .A(n5703), .Z(n5702) );
  CNIVX1 U4890 ( .A(n3384), .Z(n5703) );
  CNIVX1 U4891 ( .A(n5705), .Z(n5704) );
  CNIVX1 U4892 ( .A(n3389), .Z(n5705) );
  CNIVX1 U4893 ( .A(n5707), .Z(n5706) );
  CNIVX1 U4894 ( .A(n3385), .Z(n5707) );
  CNIVX1 U4895 ( .A(n5709), .Z(n5708) );
  CNIVX1 U4896 ( .A(n3390), .Z(n5709) );
  CNIVX1 U4897 ( .A(n5711), .Z(n5710) );
  CNIVX1 U4898 ( .A(n3386), .Z(n5711) );
  CNIVX1 U4899 ( .A(n5713), .Z(n5712) );
  CNIVX1 U4900 ( .A(n3391), .Z(n5713) );
  CNIVX1 U4901 ( .A(n5715), .Z(n5714) );
  CNIVX1 U4902 ( .A(n3387), .Z(n5715) );
  CNIVX1 U4903 ( .A(n5717), .Z(n5716) );
  CNIVX1 U4904 ( .A(n3200), .Z(n5717) );
  CNIVX1 U4905 ( .A(n5719), .Z(n5718) );
  CNIVX1 U4906 ( .A(n3388), .Z(n5719) );
  CNIVX1 U4907 ( .A(n5721), .Z(n5720) );
  CNIVX1 U4908 ( .A(n3382), .Z(n5721) );
  CNIVX1 U4909 ( .A(n5723), .Z(n5722) );
  CNIVX1 U4910 ( .A(n3349), .Z(n5723) );
  CNIVX1 U4911 ( .A(n5725), .Z(n5724) );
  CNIVX1 U4912 ( .A(n3201), .Z(n5725) );
  CNIVX1 U4913 ( .A(n5727), .Z(n5726) );
  CNIVX1 U4914 ( .A(n3380), .Z(n5727) );
  CNIVX1 U4915 ( .A(n5729), .Z(n5728) );
  CNIVX1 U4916 ( .A(n3381), .Z(n5729) );
  CNIVX1 U4917 ( .A(n5731), .Z(n5730) );
  CNIVX1 U4918 ( .A(n4068), .Z(n5731) );
  CNIVX1 U4919 ( .A(n5733), .Z(n5732) );
  CNIVX1 U4920 ( .A(n4069), .Z(n5733) );
  CNIVX1 U4921 ( .A(n5735), .Z(n5734) );
  CNIVX1 U4922 ( .A(n4070), .Z(n5735) );
  CNIVX1 U4923 ( .A(n5737), .Z(n5736) );
  CNIVX1 U4924 ( .A(n4071), .Z(n5737) );
  CNIVX1 U4925 ( .A(n5739), .Z(n5738) );
  CNIVX1 U4926 ( .A(n4072), .Z(n5739) );
  CNIVX1 U4927 ( .A(n5741), .Z(n5740) );
  CNIVX1 U4928 ( .A(n4073), .Z(n5741) );
  CNIVX1 U4929 ( .A(n5743), .Z(n5742) );
  CNIVX1 U4930 ( .A(n4074), .Z(n5743) );
  CNIVX1 U4931 ( .A(n5745), .Z(n5744) );
  CNIVX1 U4932 ( .A(n4075), .Z(n5745) );
  CNIVX1 U4933 ( .A(n5747), .Z(n5746) );
  CNIVX1 U4934 ( .A(n4078), .Z(n5747) );
  CNIVX1 U4935 ( .A(n5749), .Z(n5748) );
  CNIVX1 U4936 ( .A(n3419), .Z(n5749) );
  CNIVX1 U4937 ( .A(n5751), .Z(n5750) );
  CNIVX1 U4938 ( .A(n4079), .Z(n5751) );
  CNIVX1 U4939 ( .A(n5753), .Z(n5752) );
  CNIVX1 U4940 ( .A(n3420), .Z(n5753) );
  CNIVX1 U4941 ( .A(n5755), .Z(n5754) );
  CNIVX1 U4942 ( .A(n4086), .Z(n5755) );
  CNIVX1 U4943 ( .A(n5757), .Z(n5756) );
  CNIVX1 U4944 ( .A(n4087), .Z(n5757) );
  CNIVX1 U4945 ( .A(n5759), .Z(n5758) );
  CNIVX1 U4946 ( .A(n4088), .Z(n5759) );
  CNIVX1 U4947 ( .A(n5761), .Z(n5760) );
  CNIVX1 U4948 ( .A(n4089), .Z(n5761) );
  CNIVX1 U4949 ( .A(n5763), .Z(n5762) );
  CNIVX1 U4950 ( .A(n4090), .Z(n5763) );
  CNIVX1 U4951 ( .A(n5765), .Z(n5764) );
  CNIVX1 U4952 ( .A(n3421), .Z(n5765) );
  CNIVX1 U4953 ( .A(n5767), .Z(n5766) );
  CNIVX1 U4954 ( .A(n4091), .Z(n5767) );
  CNIVX1 U4955 ( .A(n5769), .Z(n5768) );
  CNIVX1 U4956 ( .A(n3422), .Z(n5769) );
  CNIVX1 U4957 ( .A(n5771), .Z(n5770) );
  CNIVX1 U4958 ( .A(n3423), .Z(n5771) );
  CNIVX1 U4959 ( .A(n5773), .Z(n5772) );
  CNIVX1 U4960 ( .A(n4092), .Z(n5773) );
  CNIVX1 U4961 ( .A(n5775), .Z(n5774) );
  CNIVX1 U4962 ( .A(n4093), .Z(n5775) );
  CNIVX1 U4963 ( .A(n5777), .Z(n5776) );
  CNIVX1 U4964 ( .A(n4094), .Z(n5777) );
  CNIVX1 U4965 ( .A(n5779), .Z(n5778) );
  CNIVX1 U4966 ( .A(n4095), .Z(n5779) );
  CNIVX1 U4967 ( .A(n5781), .Z(n5780) );
  CNIVX1 U4968 ( .A(n4128), .Z(n5781) );
  CNIVX1 U4969 ( .A(n5783), .Z(n5782) );
  CNIVX1 U4970 ( .A(n4129), .Z(n5783) );
  CNIVX1 U4971 ( .A(n5785), .Z(n5784) );
  CNIVX1 U4972 ( .A(n3424), .Z(n5785) );
  CNIVX1 U4973 ( .A(n5787), .Z(n5786) );
  CNIVX1 U4974 ( .A(n4130), .Z(n5787) );
  CNIVX1 U4975 ( .A(n5789), .Z(n5788) );
  CNIVX1 U4976 ( .A(n4131), .Z(n5789) );
  CNIVX1 U4977 ( .A(n5791), .Z(n5790) );
  CNIVX1 U4978 ( .A(n3425), .Z(n5791) );
  CNIVX1 U4979 ( .A(n5793), .Z(n5792) );
  CNIVX1 U4980 ( .A(n3426), .Z(n5793) );
  CNIVX1 U4981 ( .A(n5795), .Z(n5794) );
  CNIVX1 U4982 ( .A(n4132), .Z(n5795) );
  CNIVX1 U4983 ( .A(n5797), .Z(n5796) );
  CNIVX1 U4984 ( .A(n3427), .Z(n5797) );
  CNIVX1 U4985 ( .A(n5799), .Z(n5798) );
  CNIVX1 U4986 ( .A(n4133), .Z(n5799) );
  CNIVX1 U4987 ( .A(n5801), .Z(n5800) );
  CNIVX1 U4988 ( .A(n3428), .Z(n5801) );
  CNIVX1 U4989 ( .A(n5803), .Z(n5802) );
  CNIVX1 U4990 ( .A(n3429), .Z(n5803) );
  CNIVX1 U4991 ( .A(n5805), .Z(n5804) );
  CNIVX1 U4992 ( .A(n4134), .Z(n5805) );
  CNIVX1 U4993 ( .A(n5807), .Z(n5806) );
  CNIVX1 U4994 ( .A(n4135), .Z(n5807) );
  CNIVX1 U4995 ( .A(n5809), .Z(n5808) );
  CNIVX1 U4996 ( .A(n4136), .Z(n5809) );
  CNIVX1 U4997 ( .A(n5811), .Z(n5810) );
  CNIVX1 U4998 ( .A(n4137), .Z(n5811) );
  CNIVX1 U4999 ( .A(n5813), .Z(n5812) );
  CNIVX1 U5000 ( .A(n3430), .Z(n5813) );
  CNIVX1 U5001 ( .A(n5815), .Z(n5814) );
  CNIVX1 U5002 ( .A(n4138), .Z(n5815) );
  CNIVX1 U5003 ( .A(n5817), .Z(n5816) );
  CNIVX1 U5004 ( .A(n3431), .Z(n5817) );
  CNIVX1 U5005 ( .A(n5819), .Z(n5818) );
  CNIVX1 U5006 ( .A(n4139), .Z(n5819) );
  CNIVX1 U5007 ( .A(n5821), .Z(n5820) );
  CNIVX1 U5008 ( .A(n4142), .Z(n5821) );
  CNIVX1 U5009 ( .A(n5823), .Z(n5822) );
  CNIVX1 U5010 ( .A(n4143), .Z(n5823) );
  CNIVX1 U5011 ( .A(n5825), .Z(n5824) );
  CNIVX1 U5012 ( .A(n4150), .Z(n5825) );
  CNIVX1 U5013 ( .A(n5827), .Z(n5826) );
  CNIVX1 U5014 ( .A(n4151), .Z(n5827) );
  CNIVX1 U5015 ( .A(n5829), .Z(n5828) );
  CNIVX1 U5016 ( .A(n3432), .Z(n5829) );
  CNIVX1 U5017 ( .A(n5831), .Z(n5830) );
  CNIVX1 U5018 ( .A(n4152), .Z(n5831) );
  CNIVX1 U5019 ( .A(n5833), .Z(n5832) );
  CNIVX1 U5020 ( .A(n3433), .Z(n5833) );
  CNIVX1 U5021 ( .A(n5835), .Z(n5834) );
  CNIVX1 U5022 ( .A(n3434), .Z(n5835) );
  CNIVX1 U5023 ( .A(n5837), .Z(n5836) );
  CNIVX1 U5024 ( .A(n4153), .Z(n5837) );
  CNIVX1 U5025 ( .A(n5839), .Z(n5838) );
  CNIVX1 U5026 ( .A(n4154), .Z(n5839) );
  CNIVX1 U5027 ( .A(n5841), .Z(n5840) );
  CNIVX1 U5028 ( .A(n4155), .Z(n5841) );
  CNIVX1 U5029 ( .A(n5843), .Z(n5842) );
  CNIVX1 U5030 ( .A(n4156), .Z(n5843) );
  CNIVX1 U5031 ( .A(n5845), .Z(n5844) );
  CNIVX1 U5032 ( .A(n3435), .Z(n5845) );
  CNIVX1 U5033 ( .A(n5847), .Z(n5846) );
  CNIVX1 U5034 ( .A(n4157), .Z(n5847) );
  CNIVX1 U5035 ( .A(n5849), .Z(n5848) );
  CNIVX1 U5036 ( .A(n3438), .Z(n5849) );
  CNIVX1 U5037 ( .A(n5851), .Z(n5850) );
  CNIVX1 U5038 ( .A(n4158), .Z(n5851) );
  CNIVX1 U5039 ( .A(n5853), .Z(n5852) );
  CNIVX1 U5040 ( .A(n4159), .Z(n5853) );
  CNIVX1 U5041 ( .A(n5855), .Z(n5854) );
  CNIVX1 U5042 ( .A(n3439), .Z(n5855) );
  CNIVX1 U5043 ( .A(n5857), .Z(n5856) );
  CNIVX1 U5044 ( .A(n3446), .Z(n5857) );
  CNIVX1 U5045 ( .A(n5859), .Z(n5858) );
  CNIVX1 U5046 ( .A(n4192), .Z(n5859) );
  CNIVX1 U5047 ( .A(n5861), .Z(n5860) );
  CNIVX1 U5048 ( .A(n3447), .Z(n5861) );
  CNIVX1 U5049 ( .A(n5863), .Z(n5862) );
  CNIVX1 U5050 ( .A(n4193), .Z(n5863) );
  CNIVX1 U5051 ( .A(n5865), .Z(n5864) );
  CNIVX1 U5052 ( .A(n3448), .Z(n5865) );
  CNIVX1 U5053 ( .A(n5867), .Z(n5866) );
  CNIVX1 U5054 ( .A(n3449), .Z(n5867) );
  CNIVX1 U5055 ( .A(n5869), .Z(n5868) );
  CNIVX1 U5056 ( .A(n4194), .Z(n5869) );
  CNIVX1 U5057 ( .A(n5871), .Z(n5870) );
  CNIVX1 U5058 ( .A(n4195), .Z(n5871) );
  CNIVX1 U5059 ( .A(n5873), .Z(n5872) );
  CNIVX1 U5060 ( .A(n4196), .Z(n5873) );
  CNIVX1 U5061 ( .A(n5875), .Z(n5874) );
  CNIVX1 U5062 ( .A(n4197), .Z(n5875) );
  CNIVX1 U5063 ( .A(n5877), .Z(n5876) );
  CNIVX1 U5064 ( .A(n3450), .Z(n5877) );
  CNIVX1 U5065 ( .A(n5879), .Z(n5878) );
  CNIVX1 U5066 ( .A(n4198), .Z(n5879) );
  CNIVX1 U5067 ( .A(n5881), .Z(n5880) );
  CNIVX1 U5068 ( .A(n3451), .Z(n5881) );
  CNIVX1 U5069 ( .A(n5883), .Z(n5882) );
  CNIVX1 U5070 ( .A(n4199), .Z(n5883) );
  CNIVX1 U5071 ( .A(n5885), .Z(n5884) );
  CNIVX1 U5072 ( .A(n4200), .Z(n5885) );
  CNIVX1 U5073 ( .A(n5887), .Z(n5886) );
  CNIVX1 U5074 ( .A(n4201), .Z(n5887) );
  CNIVX1 U5075 ( .A(n5889), .Z(n5888) );
  CNIVX1 U5076 ( .A(n4202), .Z(n5889) );
  CNIVX1 U5077 ( .A(n5891), .Z(n5890) );
  CNIVX1 U5078 ( .A(n3452), .Z(n5891) );
  CNIVX1 U5079 ( .A(n5893), .Z(n5892) );
  CNIVX1 U5080 ( .A(n3453), .Z(n5893) );
  CNIVX1 U5081 ( .A(n5895), .Z(n5894) );
  CNIVX1 U5082 ( .A(n4203), .Z(n5895) );
  CNIVX1 U5083 ( .A(n5897), .Z(n5896) );
  CNIVX1 U5084 ( .A(n3454), .Z(n5897) );
  CNIVX1 U5085 ( .A(n5899), .Z(n5898) );
  CNIVX1 U5086 ( .A(n3455), .Z(n5899) );
  CNIVX1 U5087 ( .A(n5901), .Z(n5900) );
  CNIVX1 U5088 ( .A(n4206), .Z(n5901) );
  CNIVX1 U5089 ( .A(n5903), .Z(n5902) );
  CNIVX1 U5090 ( .A(n4207), .Z(n5903) );
  CNIVX1 U5091 ( .A(n5905), .Z(n5904) );
  CNIVX1 U5092 ( .A(n4214), .Z(n5905) );
  CNIVX1 U5093 ( .A(n5907), .Z(n5906) );
  CNIVX1 U5094 ( .A(n4215), .Z(n5907) );
  CNIVX1 U5095 ( .A(n5909), .Z(n5908) );
  CNIVX1 U5096 ( .A(n4216), .Z(n5909) );
  CNIVX1 U5097 ( .A(n5911), .Z(n5910) );
  CNIVX1 U5098 ( .A(n4217), .Z(n5911) );
  CNIVX1 U5099 ( .A(n5913), .Z(n5912) );
  CNIVX1 U5100 ( .A(n3342), .Z(n5913) );
  CNIVX1 U5101 ( .A(n5915), .Z(n5914) );
  CNIVX1 U5102 ( .A(n4218), .Z(n5915) );
  CNIVX1 U5103 ( .A(n5917), .Z(n5916) );
  CNIVX1 U5104 ( .A(n4219), .Z(n5917) );
  CNIVX1 U5105 ( .A(n5919), .Z(n5918) );
  CNIVX1 U5106 ( .A(n4220), .Z(n5919) );
  CNIVX1 U5107 ( .A(n5921), .Z(n5920) );
  CNIVX1 U5108 ( .A(n4221), .Z(n5921) );
  CNIVX1 U5109 ( .A(n5923), .Z(n5922) );
  CNIVX1 U5110 ( .A(n4222), .Z(n5923) );
  CNIVX1 U5111 ( .A(n5925), .Z(n5924) );
  CNIVX1 U5112 ( .A(n4223), .Z(n5925) );
  CNIVX1 U5113 ( .A(n5927), .Z(n5926) );
  CNIVX1 U5114 ( .A(n3984), .Z(n5927) );
  CNIVX1 U5115 ( .A(n5929), .Z(n5928) );
  CNIVX1 U5116 ( .A(n3985), .Z(n5929) );
  CNIVX1 U5117 ( .A(n5931), .Z(n5930) );
  CNIVX1 U5118 ( .A(n4044), .Z(n5931) );
  CNIVX1 U5119 ( .A(n5933), .Z(n5932) );
  CNIVX1 U5120 ( .A(n4045), .Z(n5933) );
  CNIVX1 U5121 ( .A(n5935), .Z(n5934) );
  CNIVX1 U5122 ( .A(n4048), .Z(n5935) );
  CNIVX1 U5123 ( .A(n5937), .Z(n5936) );
  CNIVX1 U5124 ( .A(n4049), .Z(n5937) );
  CNIVX1 U5125 ( .A(n5939), .Z(n5938) );
  CNIVX1 U5126 ( .A(n4112), .Z(n5939) );
  CNIVX1 U5127 ( .A(n5941), .Z(n5940) );
  CNIVX1 U5128 ( .A(n3343), .Z(n5941) );
  CNIVX1 U5129 ( .A(n5943), .Z(n5942) );
  CNIVX1 U5130 ( .A(n4113), .Z(n5943) );
  CNIVX1 U5131 ( .A(n5945), .Z(n5944) );
  CNIVX1 U5132 ( .A(n3350), .Z(n5945) );
  CNIVX1 U5133 ( .A(n5947), .Z(n5946) );
  CNIVX1 U5134 ( .A(n4172), .Z(n5947) );
  CNIVX1 U5135 ( .A(n5949), .Z(n5948) );
  CNIVX1 U5136 ( .A(n4173), .Z(n5949) );
  CNIVX1 U5137 ( .A(n5951), .Z(n5950) );
  CNIVX1 U5138 ( .A(n4176), .Z(n5951) );
  CNIVX1 U5139 ( .A(n5953), .Z(n5952) );
  CNIVX1 U5140 ( .A(n4177), .Z(n5953) );
  CNIVX1 U5141 ( .A(n5955), .Z(n5954) );
  CNIVX1 U5142 ( .A(n3787), .Z(n5955) );
  CNIVX1 U5143 ( .A(n3790), .Z(n5956) );
  CNIVX1 U5144 ( .A(n5958), .Z(n5957) );
  CNIVX1 U5145 ( .A(n3791), .Z(n5958) );
  CNIVX1 U5146 ( .A(n5960), .Z(n5959) );
  CNIVX1 U5147 ( .A(n3798), .Z(n5960) );
  CNIVX1 U5148 ( .A(n5962), .Z(n5961) );
  CNIVX1 U5149 ( .A(n3799), .Z(n5962) );
  CNIVX1 U5150 ( .A(n5964), .Z(n5963) );
  CNIVX1 U5151 ( .A(n3800), .Z(n5964) );
  CNIVX1 U5152 ( .A(n5966), .Z(n5965) );
  CNIVX1 U5153 ( .A(n3801), .Z(n5966) );
  CNIVX1 U5154 ( .A(n5968), .Z(n5967) );
  CNIVX1 U5155 ( .A(n3802), .Z(n5968) );
  CNIVX1 U5156 ( .A(n5970), .Z(n5969) );
  CNIVX1 U5157 ( .A(n3803), .Z(n5970) );
  CNIVX1 U5158 ( .A(n5972), .Z(n5971) );
  CNIVX1 U5159 ( .A(n3804), .Z(n5972) );
  CNIVX1 U5160 ( .A(n5974), .Z(n5973) );
  CNIVX1 U5161 ( .A(n3805), .Z(n5974) );
  CNIVX1 U5162 ( .A(n5976), .Z(n5975) );
  CNIVX1 U5163 ( .A(n3806), .Z(n5976) );
  CNIVX1 U5164 ( .A(n5978), .Z(n5977) );
  CNIVX1 U5165 ( .A(n3807), .Z(n5978) );
  CNIVX1 U5166 ( .A(n5980), .Z(n5979) );
  CNIVX1 U5167 ( .A(n4012), .Z(n5980) );
  CNIVX1 U5168 ( .A(n5982), .Z(n5981) );
  CNIVX1 U5169 ( .A(n4013), .Z(n5982) );
  CNIVX1 U5170 ( .A(n5984), .Z(n5983) );
  CNIVX1 U5171 ( .A(n4016), .Z(n5984) );
  CNIVX1 U5172 ( .A(n5986), .Z(n5985) );
  CNIVX1 U5173 ( .A(n4017), .Z(n5986) );
  CNIVX1 U5174 ( .A(n5988), .Z(n5987) );
  CNIVX1 U5175 ( .A(n4076), .Z(n5988) );
  CNIVX1 U5176 ( .A(n5990), .Z(n5989) );
  CNIVX1 U5177 ( .A(n4077), .Z(n5990) );
  CNIVX1 U5178 ( .A(n5992), .Z(n5991) );
  CNIVX1 U5179 ( .A(n4080), .Z(n5992) );
  CNIVX1 U5180 ( .A(n5994), .Z(n5993) );
  CNIVX1 U5181 ( .A(n4081), .Z(n5994) );
  CNIVX1 U5182 ( .A(n5996), .Z(n5995) );
  CNIVX1 U5183 ( .A(n4140), .Z(n5996) );
  CNIVX1 U5184 ( .A(n5998), .Z(n5997) );
  CNIVX1 U5185 ( .A(n4141), .Z(n5998) );
  CNIVX1 U5186 ( .A(n6000), .Z(n5999) );
  CNIVX1 U5187 ( .A(n4144), .Z(n6000) );
  CNIVX1 U5188 ( .A(n6002), .Z(n6001) );
  CNIVX1 U5189 ( .A(n3351), .Z(n6002) );
  CNIVX1 U5190 ( .A(n6004), .Z(n6003) );
  CNIVX1 U5191 ( .A(n4145), .Z(n6004) );
  CNIVX1 U5192 ( .A(n6006), .Z(n6005) );
  CNIVX1 U5193 ( .A(n4204), .Z(n6006) );
  CNIVX1 U5194 ( .A(n6008), .Z(n6007) );
  CNIVX1 U5195 ( .A(n4205), .Z(n6008) );
  CNIVX1 U5196 ( .A(n6010), .Z(n6009) );
  CNIVX1 U5197 ( .A(n4208), .Z(n6010) );
  CNIVX1 U5198 ( .A(n6012), .Z(n6011) );
  CNIVX1 U5199 ( .A(n4209), .Z(n6012) );
  CNIVX1 U5200 ( .A(n6014), .Z(n6013) );
  CNIVX1 U5201 ( .A(n3352), .Z(n6014) );
  CNIVX1 U5202 ( .A(n6016), .Z(n6015) );
  CNIVX1 U5203 ( .A(n3986), .Z(n6016) );
  CNIVX1 U5204 ( .A(n6018), .Z(n6017) );
  CNIVX1 U5205 ( .A(n3987), .Z(n6018) );
  CNIVX1 U5206 ( .A(n6020), .Z(n6019) );
  CNIVX1 U5207 ( .A(n3353), .Z(n6020) );
  CNIVX1 U5208 ( .A(n6022), .Z(n6021) );
  CNIVX1 U5209 ( .A(n3988), .Z(n6022) );
  CNIVX1 U5210 ( .A(n6024), .Z(n6023) );
  CNIVX1 U5211 ( .A(n3989), .Z(n6024) );
  CNIVX1 U5212 ( .A(n6026), .Z(n6025) );
  CNIVX1 U5213 ( .A(n4050), .Z(n6026) );
  CNIVX1 U5214 ( .A(n6028), .Z(n6027) );
  CNIVX1 U5215 ( .A(n4051), .Z(n6028) );
  CNIVX1 U5216 ( .A(n6030), .Z(n6029) );
  CNIVX1 U5217 ( .A(n4052), .Z(n6030) );
  CNIVX1 U5218 ( .A(n6032), .Z(n6031) );
  CNIVX1 U5219 ( .A(n4053), .Z(n6032) );
  CNIVX1 U5220 ( .A(n6034), .Z(n6033) );
  CNIVX1 U5221 ( .A(n4114), .Z(n6034) );
  CNIVX1 U5222 ( .A(n6036), .Z(n6035) );
  CNIVX1 U5223 ( .A(n4115), .Z(n6036) );
  CNIVX1 U5224 ( .A(n6038), .Z(n6037) );
  CNIVX1 U5225 ( .A(n4116), .Z(n6038) );
  CNIVX1 U5226 ( .A(n6040), .Z(n6039) );
  CNIVX1 U5227 ( .A(n3354), .Z(n6040) );
  CNIVX1 U5228 ( .A(n6042), .Z(n6041) );
  CNIVX1 U5229 ( .A(n3355), .Z(n6042) );
  CNIVX1 U5230 ( .A(n6044), .Z(n6043) );
  CNIVX1 U5231 ( .A(n4117), .Z(n6044) );
  CNIVX1 U5232 ( .A(n6046), .Z(n6045) );
  CNIVX1 U5233 ( .A(n4178), .Z(n6046) );
  CNIVX1 U5234 ( .A(n6048), .Z(n6047) );
  CNIVX1 U5235 ( .A(n4179), .Z(n6048) );
  CNIVX1 U5236 ( .A(n6050), .Z(n6049) );
  CNIVX1 U5237 ( .A(n4180), .Z(n6050) );
  CNIVX1 U5238 ( .A(n6052), .Z(n6051) );
  CNIVX1 U5239 ( .A(n4181), .Z(n6052) );
  CNIVX1 U5240 ( .A(n6054), .Z(n6053) );
  CNIVX1 U5241 ( .A(n4018), .Z(n6054) );
  CNIVX1 U5242 ( .A(n6056), .Z(n6055) );
  CNIVX1 U5243 ( .A(n4019), .Z(n6056) );
  CNIVX1 U5244 ( .A(n6058), .Z(n6057) );
  CNIVX1 U5245 ( .A(n4020), .Z(n6058) );
  CNIVX1 U5246 ( .A(n6060), .Z(n6059) );
  CNIVX1 U5247 ( .A(n4021), .Z(n6060) );
  CNIVX1 U5248 ( .A(n6062), .Z(n6061) );
  CNIVX1 U5249 ( .A(n4082), .Z(n6062) );
  CNIVX1 U5250 ( .A(n6064), .Z(n6063) );
  CNIVX1 U5251 ( .A(n4083), .Z(n6064) );
  CNIVX1 U5252 ( .A(n6066), .Z(n6065) );
  CNIVX1 U5253 ( .A(n4084), .Z(n6066) );
  CNIVX1 U5254 ( .A(n6068), .Z(n6067) );
  CNIVX1 U5255 ( .A(n4085), .Z(n6068) );
  CNIVX1 U5256 ( .A(n6070), .Z(n6069) );
  CNIVX1 U5257 ( .A(n4146), .Z(n6070) );
  CNIVX1 U5258 ( .A(n6072), .Z(n6071) );
  CNIVX1 U5259 ( .A(n4147), .Z(n6072) );
  CNIVX1 U5260 ( .A(n6074), .Z(n6073) );
  CNIVX1 U5261 ( .A(n4148), .Z(n6074) );
  CNIVX1 U5262 ( .A(n6076), .Z(n6075) );
  CNIVX1 U5263 ( .A(n4149), .Z(n6076) );
  CNIVX1 U5264 ( .A(n6078), .Z(n6077) );
  CNIVX1 U5265 ( .A(n3356), .Z(n6078) );
  CNIVX1 U5266 ( .A(n6080), .Z(n6079) );
  CNIVX1 U5267 ( .A(n4210), .Z(n6080) );
  CNIVX1 U5268 ( .A(n6082), .Z(n6081) );
  CNIVX1 U5269 ( .A(n3357), .Z(n6082) );
  CNIVX1 U5270 ( .A(n6084), .Z(n6083) );
  CNIVX1 U5271 ( .A(n3358), .Z(n6084) );
  CNIVX1 U5272 ( .A(n6086), .Z(n6085) );
  CNIVX1 U5273 ( .A(n4211), .Z(n6086) );
  CNIVX1 U5274 ( .A(n6088), .Z(n6087) );
  CNIVX1 U5275 ( .A(n4212), .Z(n6088) );
  CNIVX1 U5276 ( .A(n6090), .Z(n6089) );
  CNIVX1 U5277 ( .A(n3359), .Z(n6090) );
  CNIVX1 U5278 ( .A(n6092), .Z(n6091) );
  CNIVX1 U5279 ( .A(n3360), .Z(n6092) );
  CNIVX1 U5280 ( .A(n6094), .Z(n6093) );
  CNIVX1 U5281 ( .A(n3361), .Z(n6094) );
  CNIVX1 U5282 ( .A(n6096), .Z(n6095) );
  CNIVX1 U5283 ( .A(n4213), .Z(n6096) );
  CNIVX1 U5284 ( .A(n6098), .Z(n6097) );
  CNIVX1 U5285 ( .A(n4235), .Z(n6098) );
  CNIVX1 U5286 ( .A(n6100), .Z(n6099) );
  CNIVX1 U5287 ( .A(n3362), .Z(n6100) );
  CNIVX1 U5288 ( .A(n6102), .Z(n6101) );
  CNIVX1 U5289 ( .A(n3467), .Z(n6102) );
  CNIVX1 U5290 ( .A(n6104), .Z(n6103) );
  CNIVX1 U5291 ( .A(n3723), .Z(n6104) );
  CNIVX1 U5292 ( .A(n6106), .Z(n6105) );
  CNIVX1 U5293 ( .A(n3363), .Z(n6106) );
  CNIVX1 U5294 ( .A(n6108), .Z(n6107) );
  CNIVX1 U5295 ( .A(n3364), .Z(n6108) );
  CNIVX1 U5296 ( .A(n6110), .Z(n6109) );
  CNIVX1 U5297 ( .A(n3979), .Z(n6110) );
  CNIVX1 U5298 ( .A(n6112), .Z(n6111) );
  CNIVX1 U5299 ( .A(n3347), .Z(n6112) );
  CNIVX1 U5300 ( .A(n6114), .Z(n6113) );
  CNIVX1 U5301 ( .A(n3348), .Z(n6114) );
  CNIVX1 U5302 ( .A(n6116), .Z(n6115) );
  CNIVX1 U5303 ( .A(n3777), .Z(n6116) );
  CNIVX1 U5304 ( .A(n6118), .Z(n6117) );
  CNIVX1 U5305 ( .A(n3813), .Z(n6118) );
  CNIVX1 U5306 ( .A(n6120), .Z(n6119) );
  CNIVX1 U5307 ( .A(n3778), .Z(n6120) );
  CNIVX1 U5308 ( .A(n6122), .Z(n6121) );
  CNIVX1 U5309 ( .A(n3779), .Z(n6122) );
  CNIVX1 U5310 ( .A(n6124), .Z(n6123) );
  CNIVX1 U5311 ( .A(n3780), .Z(n6124) );
  CNIVX1 U5312 ( .A(n6126), .Z(n6125) );
  CNIVX1 U5313 ( .A(n3781), .Z(n6126) );
  CNIVX1 U5314 ( .A(n6128), .Z(n6127) );
  CNIVX1 U5315 ( .A(n3782), .Z(n6128) );
  CNIVX1 U5316 ( .A(n6130), .Z(n6129) );
  CNIVX1 U5317 ( .A(n3783), .Z(n6130) );
  CNIVX1 U5318 ( .A(n6132), .Z(n6131) );
  CNIVX1 U5319 ( .A(n3784), .Z(n6132) );
  CNIVX1 U5320 ( .A(n6134), .Z(n6133) );
  CNIVX1 U5321 ( .A(n3785), .Z(n6134) );
  CNIVX1 U5322 ( .A(n6136), .Z(n6135) );
  CNIVX1 U5323 ( .A(n3786), .Z(n6136) );
  CNIVX1 U5324 ( .A(n6138), .Z(n6137) );
  CNIVX1 U5325 ( .A(n3314), .Z(n6138) );
  CNIVX1 U5326 ( .A(n6140), .Z(n6139) );
  CNIVX1 U5327 ( .A(n3368), .Z(n6140) );
  CNIVX1 U5328 ( .A(n6142), .Z(n6141) );
  CNIVX1 U5329 ( .A(dataout_stg_1[6]), .Z(n6142) );
  CNIVX1 U5330 ( .A(n6144), .Z(n6143) );
  CNIVX1 U5331 ( .A(n3367), .Z(n6144) );
  CNIVX1 U5332 ( .A(n6146), .Z(n6145) );
  CNIVX1 U5333 ( .A(n3366), .Z(n6146) );
  CNIVX1 U5334 ( .A(n6148), .Z(n6147) );
  CNIVX1 U5335 ( .A(n3371), .Z(n6148) );
  CANR1XL U5336 ( .A(n8303), .B(n904), .C(n905), .Z(n903) );
  CAN4X1 U5337 ( .A(n591), .B(n592), .C(n593), .D(n594), .Z(n590) );
  CIVX1 U5338 ( .A(rd_ptr[8]), .Z(n8311) );
  CANR2X1 U5339 ( .A(n7096), .B(buffer[515]), .C(n8301), .D(n298), .Z(n592) );
  COND2X2 U5340 ( .A(n7140), .B(n7693), .C(n7139), .D(n7437), .Z(n1922) );
  COND2X1 U5341 ( .A(n906), .B(n76), .C(n907), .D(n35), .Z(n905) );
  COND1XL U5342 ( .A(n8287), .B(n6155), .C(n287), .Z(n284) );
  CIVX1 U5343 ( .A(n258), .Z(n7213) );
  COND1XL U5344 ( .A(n8307), .B(n7789), .C(n1911), .Z(n1906) );
  COND1XL U5345 ( .A(n8296), .B(n187), .C(n1302), .Z(n355) );
  CAN2XL U5346 ( .A(n284), .B(n6163), .Z(n285) );
  CNR2XL U5347 ( .A(n8311), .B(rd_ptr[9]), .Z(n6149) );
  CANR2X1 U5348 ( .A(n7237), .B(n8285), .C(n60), .D(n8286), .Z(n104) );
  CANR2X1 U5349 ( .A(n8301), .B(n278), .C(n8303), .D(n279), .Z(n1403) );
  CNIVXL U5350 ( .A(n84), .Z(n7146) );
  CNIVX8 U5351 ( .A(n86), .Z(n7139) );
  COND4CX1 U5352 ( .A(n7216), .B(n178), .C(n349), .D(n351), .Z(n343) );
  COND2XL U5353 ( .A(n7136), .B(n7790), .C(n7130), .D(n8046), .Z(n1185) );
  COND2XL U5354 ( .A(n7136), .B(n7854), .C(n7130), .D(n8110), .Z(n1173) );
  COND2XL U5355 ( .A(n7113), .B(n7986), .C(n7168), .D(n8242), .Z(n510) );
  CANR2XL U5356 ( .A(n8288), .B(n48), .C(n8286), .D(n17), .Z(n109) );
  COND2X1 U5357 ( .A(n7141), .B(n7733), .C(n7139), .D(n7477), .Z(n1824) );
  CND2XL U5358 ( .A(n8288), .B(n17), .Z(n153) );
  CANR2XL U5359 ( .A(n8286), .B(n207), .C(n8285), .D(n288), .Z(n287) );
  COND2XL U5360 ( .A(n7136), .B(n7798), .C(n7131), .D(n8054), .Z(n1010) );
  COND2XL U5361 ( .A(n7136), .B(n7862), .C(n7131), .D(n8118), .Z(n1022) );
  COND2XL U5362 ( .A(n7135), .B(n7867), .C(n7129), .D(n8123), .Z(n1226) );
  COND2XL U5363 ( .A(n7122), .B(n7987), .C(n7164), .D(n8243), .Z(n1323) );
  COND2XL U5364 ( .A(n7136), .B(n7830), .C(n7131), .D(n8086), .Z(n1034) );
  COND2XL U5365 ( .A(n7120), .B(n7923), .C(n7164), .D(n8179), .Z(n1335) );
  COND2XL U5366 ( .A(n7112), .B(n7971), .C(n7164), .D(n8227), .Z(n1351) );
  COND2XL U5367 ( .A(n7112), .B(n7939), .C(n7164), .D(n8195), .Z(n1377) );
  COND2XL U5368 ( .A(n7112), .B(n7907), .C(n7163), .D(n8163), .Z(n1389) );
  CND4XL U5369 ( .A(n1606), .B(n1607), .C(n1608), .D(n1609), .Z(n1605) );
  COR2X1 U5370 ( .A(n330), .B(n8287), .Z(n372) );
  CNR2XL U5371 ( .A(n8311), .B(rd_ptr[9]), .Z(n386) );
  COR3X1 U5372 ( .A(n8), .B(n7233), .C(n172), .Z(n6150) );
  CND2X1 U5373 ( .A(n6150), .B(n173), .Z(n170) );
  CIVXL U5374 ( .A(n199), .Z(n7233) );
  CND2X1 U5375 ( .A(n6154), .B(n306), .Z(n301) );
  CIVX2 U5376 ( .A(n7216), .Z(n6151) );
  CIVX2 U5377 ( .A(n7241), .Z(n6152) );
  CIVX2 U5378 ( .A(n7219), .Z(n6153) );
  CIVXL U5379 ( .A(n301), .Z(n7214) );
  COND2XL U5380 ( .A(rd_ptr[2]), .B(n289), .C(n8290), .D(n155), .Z(n6155) );
  COND2XL U5381 ( .A(n7136), .B(n7868), .C(n7125), .D(n8124), .Z(n962) );
  COND2XL U5382 ( .A(n7136), .B(n7772), .C(n7129), .D(n8028), .Z(n988) );
  COND2XL U5383 ( .A(n7136), .B(n7836), .C(n7126), .D(n8092), .Z(n950) );
  COND2XL U5384 ( .A(n7136), .B(n7804), .C(n7127), .D(n8060), .Z(n976) );
  COND2XL U5385 ( .A(n7137), .B(n7780), .C(n7129), .D(n8036), .Z(n880) );
  COND2XL U5386 ( .A(n7137), .B(n7812), .C(n7127), .D(n8068), .Z(n868) );
  CNIVXL U5387 ( .A(n8309), .Z(n7098) );
  CNIVXL U5388 ( .A(n8309), .Z(n7103) );
  CNIVXL U5389 ( .A(n8309), .Z(n7102) );
  CNIVXL U5390 ( .A(n8309), .Z(n7105) );
  CNIVXL U5391 ( .A(n8309), .Z(n7104) );
  CNIVXL U5392 ( .A(n8309), .Z(n7099) );
  CNIVXL U5393 ( .A(n8309), .Z(n7107) );
  CNR2XL U5394 ( .A(n33), .B(n7161), .Z(n381) );
  CNR2XL U5395 ( .A(n33), .B(n7139), .Z(n390) );
  CNIVXL U5396 ( .A(n84), .Z(n7148) );
  CNIVXL U5397 ( .A(n84), .Z(n7147) );
  CNIVXL U5398 ( .A(n84), .Z(n7143) );
  CNIVXL U5399 ( .A(n84), .Z(n7144) );
  CNIVXL U5400 ( .A(n84), .Z(n7145) );
  CNIVXL U5401 ( .A(n84), .Z(n7141) );
  CNIVXL U5402 ( .A(n84), .Z(n7142) );
  CNIVXL U5403 ( .A(n80), .Z(n7168) );
  CANR2XL U5404 ( .A(n8301), .B(n195), .C(n8298), .D(n197), .Z(n188) );
  CANR2XL U5405 ( .A(n8301), .B(n325), .C(n8303), .D(n326), .Z(n1606) );
  CANR2XL U5406 ( .A(n8303), .B(n218), .C(n8298), .D(n219), .Z(n212) );
  CANR2XL U5407 ( .A(n8306), .B(n299), .C(n8303), .D(n300), .Z(n591) );
  CANR2XL U5408 ( .A(n8306), .B(n341), .C(n8303), .D(n342), .Z(n376) );
  CNIVXL U5409 ( .A(n84), .Z(n7149) );
  CANR2XL U5410 ( .A(n8291), .B(n114), .C(n8295), .D(n115), .Z(n113) );
  COND2XL U5411 ( .A(n7148), .B(n7666), .C(n7139), .D(n7410), .Z(n523) );
  COND2XL U5412 ( .A(n7144), .B(n7662), .C(n7139), .D(n7406), .Z(n1184) );
  COND2XL U5413 ( .A(n7133), .B(n7793), .C(n7124), .D(n8049), .Z(n1791) );
  COND2XL U5414 ( .A(n7148), .B(n7730), .C(n7139), .D(n7474), .Z(n511) );
  COND2XL U5415 ( .A(n7144), .B(n7726), .C(n7139), .D(n7470), .Z(n1172) );
  COND2XL U5416 ( .A(n7133), .B(n7857), .C(n7124), .D(n8113), .Z(n1779) );
  CNIVXL U5417 ( .A(n396), .Z(n7138) );
  CANR2XL U5418 ( .A(n266), .B(n8285), .C(n198), .D(n8286), .Z(n265) );
  COND3XL U5419 ( .A(n156), .B(n69), .C(n157), .D(n158), .Z(n17) );
  CANR2XL U5420 ( .A(n8291), .B(n159), .C(n8295), .D(n160), .Z(n158) );
  COND11XL U5421 ( .A(n161), .B(n162), .C(n163), .D(n8294), .Z(n157) );
  CND2XL U5422 ( .A(n132), .B(n104), .Z(n101) );
  CND2XL U5423 ( .A(n8285), .B(n129), .Z(n108) );
  CND2XL U5424 ( .A(n8285), .B(n198), .Z(n180) );
  COND2XL U5425 ( .A(n7151), .B(n7275), .C(n7102), .D(n7534), .Z(n1186) );
  COND2XL U5426 ( .A(n7154), .B(n7346), .C(n7098), .D(n7602), .Z(n513) );
  COND2XL U5427 ( .A(n7155), .B(n7342), .C(n7102), .D(n7598), .Z(n1174) );
  COND2XL U5428 ( .A(n7150), .B(n7280), .C(n7106), .D(n7537), .Z(n1792) );
  COND2XL U5429 ( .A(n7151), .B(n7345), .C(n7106), .D(n7601), .Z(n1780) );
  COND2XL U5430 ( .A(n7147), .B(n7728), .C(n7139), .D(n7472), .Z(n703) );
  COND2XL U5431 ( .A(n142), .B(n33), .C(n143), .D(n35), .Z(n141) );
  COND2XL U5432 ( .A(n164), .B(n33), .C(n165), .D(n35), .Z(n163) );
  COND2XL U5433 ( .A(n7138), .B(n7794), .C(n7128), .D(n8050), .Z(n524) );
  COND2XL U5434 ( .A(n1198), .B(n16), .C(n7249), .D(n21), .Z(n1196) );
  CANR3XL U5435 ( .A(n8292), .B(n23), .C(n24), .D(n25), .Z(n20) );
  COND2XL U5436 ( .A(n7137), .B(n7792), .C(n7130), .D(n8048), .Z(n713) );
  COND2XL U5437 ( .A(n7137), .B(n7856), .C(n7130), .D(n8112), .Z(n701) );
  COND2XL U5438 ( .A(n7159), .B(n7278), .C(n7099), .D(n7536), .Z(n712) );
  COND2XL U5439 ( .A(n7153), .B(n7276), .C(n7104), .D(n7535), .Z(n1537) );
  COND2XL U5440 ( .A(n7115), .B(n7980), .C(n7166), .D(n8236), .Z(n926) );
  COND2XL U5441 ( .A(n7123), .B(n7988), .C(n7166), .D(n8244), .Z(n811) );
  COND2XL U5442 ( .A(n7123), .B(n7956), .C(n7166), .D(n8212), .Z(n823) );
  COND2XL U5443 ( .A(n7123), .B(n7924), .C(n7166), .D(n8180), .Z(n799) );
  COND2XL U5444 ( .A(n7123), .B(n7940), .C(n7166), .D(n8196), .Z(n865) );
  COND2XL U5445 ( .A(n7123), .B(n7972), .C(n7166), .D(n8228), .Z(n839) );
  COND2XL U5446 ( .A(n7112), .B(n7968), .C(n7166), .D(n8224), .Z(n752) );
  COND2XL U5447 ( .A(n7112), .B(n7936), .C(n7166), .D(n8192), .Z(n766) );
  COND2XL U5448 ( .A(n7112), .B(n7904), .C(n7166), .D(n8160), .Z(n778) );
  COND2XL U5449 ( .A(n7123), .B(n7909), .C(n7161), .D(n8165), .Z(n1889) );
  COND2XL U5450 ( .A(n7123), .B(n8005), .C(n7161), .D(n8261), .Z(n1863) );
  COND2XL U5451 ( .A(n7115), .B(n7964), .C(n7166), .D(n8220), .Z(n947) );
  COND2XL U5452 ( .A(n7115), .B(n7996), .C(n7166), .D(n8252), .Z(n959) );
  COND2XL U5453 ( .A(n7120), .B(n7908), .C(n7166), .D(n8164), .Z(n877) );
  COND2XL U5454 ( .A(n7123), .B(n8004), .C(n7166), .D(n8260), .Z(n851) );
  COND2XL U5455 ( .A(n7140), .B(n7725), .C(n7139), .D(n7469), .Z(n1938) );
  COND2XL U5456 ( .A(n7147), .B(n7648), .C(n7139), .D(n7392), .Z(n779) );
  COND2XL U5457 ( .A(n7149), .B(n7674), .C(n7139), .D(n7418), .Z(n422) );
  COND2XL U5458 ( .A(n7147), .B(n7752), .C(n7139), .D(n7496), .Z(n651) );
  COND2XL U5459 ( .A(n7148), .B(n7650), .C(n7139), .D(n7394), .Z(n577) );
  COND2XL U5460 ( .A(n7146), .B(n7748), .C(n7139), .D(n7492), .Z(n852) );
  COND2XL U5461 ( .A(n7149), .B(n7754), .C(n7139), .D(n7498), .Z(n450) );
  COND2XL U5462 ( .A(n7140), .B(n7677), .C(n7139), .D(n7421), .Z(n1982) );
  COND2XL U5463 ( .A(n7140), .B(n7709), .C(n7139), .D(n7453), .Z(n1956) );
  COND2XL U5464 ( .A(n7140), .B(n7741), .C(n7139), .D(n7485), .Z(n1968) );
  COND2XL U5465 ( .A(n7140), .B(n7749), .C(n7139), .D(n7493), .Z(n1864) );
  COND2XL U5466 ( .A(n7144), .B(n7645), .C(n7139), .D(n7389), .Z(n1994) );
  COND2XL U5467 ( .A(n7144), .B(n7755), .C(n7139), .D(n7499), .Z(n1265) );
  COND2XL U5468 ( .A(n7143), .B(n7747), .C(n7139), .D(n7491), .Z(n1364) );
  COND2XL U5469 ( .A(n7145), .B(n7734), .C(n7139), .D(n7478), .Z(n1020) );
  COND2XL U5470 ( .A(n7137), .B(n7844), .C(n7132), .D(n8100), .Z(n842) );
  COND2XL U5471 ( .A(n7146), .B(n7716), .C(n7139), .D(n7460), .Z(n840) );
  COND2XL U5472 ( .A(n7150), .B(n7349), .C(n7106), .D(n7605), .Z(n1825) );
  COND2XL U5473 ( .A(n7150), .B(n7317), .C(n7106), .D(n7573), .Z(n1837) );
  COND2XL U5474 ( .A(n7150), .B(n7301), .C(n7106), .D(n7557), .Z(n1879) );
  COND2XL U5475 ( .A(n7150), .B(n7333), .C(n7106), .D(n7589), .Z(n1853) );
  COND2XL U5476 ( .A(n7150), .B(n7365), .C(n7106), .D(n7621), .Z(n1865) );
  COND2XL U5477 ( .A(n7151), .B(n7297), .C(n7105), .D(n7553), .Z(n1735) );
  COND2XL U5478 ( .A(n7151), .B(n7256), .C(n7105), .D(n7521), .Z(n1747) );
  COND2XL U5479 ( .A(n7151), .B(n7329), .C(n7105), .D(n7585), .Z(n1709) );
  COND2XL U5480 ( .A(n7151), .B(n7361), .C(n7105), .D(n7617), .Z(n1721) );
  COND2XL U5481 ( .A(n7152), .B(n7305), .C(n7105), .D(n7561), .Z(n1681) );
  COND2XL U5482 ( .A(n7151), .B(n7267), .C(n7105), .D(n7529), .Z(n1693) );
  COND2XL U5483 ( .A(n7152), .B(n7337), .C(n7105), .D(n7593), .Z(n1655) );
  COND2XL U5484 ( .A(n7152), .B(n7369), .C(n7105), .D(n7625), .Z(n1667) );
  COND2XL U5485 ( .A(n7152), .B(n7254), .C(n7104), .D(n7519), .Z(n1593) );
  COND2XL U5486 ( .A(n7160), .B(n7322), .C(n7098), .D(n7578), .Z(n394) );
  COND2XL U5487 ( .A(n7137), .B(n7872), .C(n7131), .D(n8128), .Z(n743) );
  COND2XL U5488 ( .A(n7159), .B(n7360), .C(n7100), .D(n7616), .Z(n742) );
  COND2XL U5489 ( .A(n7147), .B(n7744), .C(n7139), .D(n7488), .Z(n741) );
  COND2XL U5490 ( .A(n7160), .B(n7338), .C(n7098), .D(n7594), .Z(n439) );
  COND2XL U5491 ( .A(n7160), .B(n7306), .C(n7098), .D(n7562), .Z(n465) );
  COND2XL U5492 ( .A(n7160), .B(n7315), .C(n7103), .D(n7571), .Z(n1313) );
  COND2XL U5493 ( .A(n7150), .B(n7310), .C(n7102), .D(n7566), .Z(n1160) );
  COND2XL U5494 ( .A(n7155), .B(n7339), .C(n7102), .D(n7595), .Z(n1254) );
  COND2XL U5495 ( .A(n7155), .B(n7307), .C(n7103), .D(n7563), .Z(n1280) );
  COND2XL U5496 ( .A(n7159), .B(n7331), .C(n7103), .D(n7587), .Z(n1353) );
  COND2XL U5497 ( .A(n7154), .B(n7299), .C(n7103), .D(n7555), .Z(n1379) );
  COND2XL U5498 ( .A(n7138), .B(n7864), .C(n7124), .D(n8120), .Z(n612) );
  COND2XL U5499 ( .A(n7155), .B(n7371), .C(n7102), .D(n7627), .Z(n1266) );
  COND2XL U5500 ( .A(n7155), .B(n7271), .C(n7103), .D(n7531), .Z(n1292) );
  COND2XL U5501 ( .A(n7152), .B(n7326), .C(n7102), .D(n7582), .Z(n1103) );
  COND2XL U5502 ( .A(n7159), .B(n7294), .C(n7102), .D(n7550), .Z(n1129) );
  COND2XL U5503 ( .A(n7143), .B(n7719), .C(n7139), .D(n7463), .Z(n1451) );
  COND2XL U5504 ( .A(n7154), .B(n7335), .C(n7104), .D(n7591), .Z(n1452) );
  COND2XL U5505 ( .A(n7143), .B(n7687), .C(n7139), .D(n7431), .Z(n1477) );
  COND2XL U5506 ( .A(n7154), .B(n7303), .C(n7104), .D(n7559), .Z(n1478) );
  COND2XL U5507 ( .A(n7152), .B(n7363), .C(n7103), .D(n7619), .Z(n1365) );
  COND2XL U5508 ( .A(n7151), .B(n7313), .C(n7105), .D(n7569), .Z(n1766) );
  COND2XL U5509 ( .A(n7152), .B(n7353), .C(n7105), .D(n7609), .Z(n1627) );
  COND2XL U5510 ( .A(n7137), .B(n7800), .C(n7124), .D(n8056), .Z(n624) );
  COND2XL U5511 ( .A(n7155), .B(n7259), .C(n7103), .D(n7523), .Z(n1391) );
  COND2XL U5512 ( .A(n7150), .B(n7358), .C(n7102), .D(n7614), .Z(n1115) );
  COND2XL U5513 ( .A(n7151), .B(n7253), .C(n7102), .D(n7518), .Z(n1141) );
  COND2XL U5514 ( .A(n7152), .B(n7321), .C(n7105), .D(n7577), .Z(n1639) );
  COND2XL U5515 ( .A(n7150), .B(n7285), .C(n7106), .D(n7541), .Z(n1813) );
  COND2XL U5516 ( .A(n7160), .B(n7370), .C(n7098), .D(n7626), .Z(n451) );
  COND2XL U5517 ( .A(n7154), .B(n7269), .C(n7098), .D(n7530), .Z(n477) );
  COND2XL U5518 ( .A(n7154), .B(n7264), .C(n7104), .D(n7527), .Z(n1490) );
  COND2XL U5519 ( .A(n7157), .B(n7292), .C(n7101), .D(n7548), .Z(n975) );
  COND2XL U5520 ( .A(n7157), .B(n7248), .C(n7101), .D(n7516), .Z(n987) );
  COND2XL U5521 ( .A(n7156), .B(n7366), .C(n7101), .D(n7622), .Z(n1061) );
  COND2XL U5522 ( .A(n7153), .B(n7327), .C(n7104), .D(n7583), .Z(n1567) );
  COND2XL U5523 ( .A(n7137), .B(n7816), .C(n7127), .D(n8072), .Z(n667) );
  COND2XL U5524 ( .A(n7137), .B(n7784), .C(n7125), .D(n8040), .Z(n679) );
  COND2XL U5525 ( .A(n7137), .B(n7848), .C(n7127), .D(n8104), .Z(n641) );
  COND2XL U5526 ( .A(n7137), .B(n7880), .C(n7128), .D(n8136), .Z(n653) );
  COND2XL U5527 ( .A(n7137), .B(n7776), .C(n7132), .D(n8032), .Z(n781) );
  COND2XL U5528 ( .A(n7138), .B(n7778), .C(n7128), .D(n8034), .Z(n579) );
  COND2XL U5529 ( .A(n7160), .B(n7354), .C(n7098), .D(n7610), .Z(n412) );
  COND2XL U5530 ( .A(n7159), .B(n7347), .C(n7103), .D(n7603), .Z(n1326) );
  COND2XL U5531 ( .A(n7154), .B(n7283), .C(n7103), .D(n7539), .Z(n1338) );
  COND2XL U5532 ( .A(n7138), .B(n7832), .C(n7131), .D(n8088), .Z(n601) );
  COND2XL U5533 ( .A(n7137), .B(n7876), .C(n7132), .D(n8132), .Z(n854) );
  COND2XL U5534 ( .A(n7138), .B(n7882), .C(n7126), .D(n8138), .Z(n452) );
  COND2XL U5535 ( .A(n7133), .B(n7877), .C(n7124), .D(n8133), .Z(n1866) );
  CANR2XL U5536 ( .A(n8289), .B(n129), .C(n8285), .D(n155), .Z(n154) );
  CANR2XL U5537 ( .A(n8292), .B(n44), .C(n8291), .D(n249), .Z(n248) );
  CANR2XL U5538 ( .A(n8292), .B(n184), .C(n8291), .D(n185), .Z(n183) );
  COND2XL U5539 ( .A(n7146), .B(n7660), .C(n7139), .D(n7404), .Z(n921) );
  COND2XL U5540 ( .A(n7115), .B(n7916), .C(n7166), .D(n8172), .Z(n920) );
  CANR2XL U5541 ( .A(n8289), .B(n198), .C(n8285), .D(n226), .Z(n225) );
  COND3XL U5542 ( .A(n179), .B(n19), .C(n224), .D(n225), .Z(n202) );
  COND2XL U5543 ( .A(n7123), .B(n7989), .C(n7161), .D(n8245), .Z(n1823) );
  COND2XL U5544 ( .A(n7133), .B(n7861), .C(n7124), .D(n8117), .Z(n1826) );
  COND2XL U5545 ( .A(n7133), .B(n7797), .C(n7124), .D(n8053), .Z(n1814) );
  COND2XL U5546 ( .A(n7144), .B(n7699), .C(n7139), .D(n7443), .Z(n1312) );
  COND2XL U5547 ( .A(n7112), .B(n7962), .C(n7161), .D(n8218), .Z(n392) );
  COND2XL U5548 ( .A(n7160), .B(n7320), .C(n7099), .D(n7576), .Z(n600) );
  COND2XL U5549 ( .A(n7148), .B(n7736), .C(n7139), .D(n7480), .Z(n611) );
  COND2XL U5550 ( .A(n7159), .B(n7352), .C(n7099), .D(n7608), .Z(n613) );
  COND2XL U5551 ( .A(n7149), .B(n7738), .C(n7139), .D(n7482), .Z(n410) );
  COND2XL U5552 ( .A(n7138), .B(n7866), .C(n7124), .D(n8122), .Z(n411) );
  COND2XL U5553 ( .A(n7143), .B(n7735), .C(n7139), .D(n7479), .Z(n1423) );
  COND2XL U5554 ( .A(n7154), .B(n7351), .C(n7103), .D(n7607), .Z(n1424) );
  COND2XL U5555 ( .A(n7143), .B(n7731), .C(n7139), .D(n7475), .Z(n1324) );
  COND2XL U5556 ( .A(n7155), .B(n7355), .C(n7102), .D(n7611), .Z(n1227) );
  COND2XL U5557 ( .A(n7137), .B(n7860), .C(n7132), .D(n8116), .Z(n814) );
  COND2XL U5558 ( .A(n7146), .B(n7732), .C(n7139), .D(n7476), .Z(n812) );
  COND2XL U5559 ( .A(n7144), .B(n7707), .C(n7139), .D(n7451), .Z(n1213) );
  COND2XL U5560 ( .A(n7155), .B(n7291), .C(n7102), .D(n7547), .Z(n1239) );
  COND2XL U5561 ( .A(n7144), .B(n7675), .C(n7139), .D(n7419), .Z(n1237) );
  COND2XL U5562 ( .A(n7123), .B(n7957), .C(n7161), .D(n8213), .Z(n1835) );
  COND2XL U5563 ( .A(n7140), .B(n7701), .C(n7139), .D(n7445), .Z(n1836) );
  COND2XL U5564 ( .A(n7133), .B(n7829), .C(n7124), .D(n8085), .Z(n1838) );
  COND2XL U5565 ( .A(n7148), .B(n7672), .C(n7139), .D(n7416), .Z(n623) );
  COND2XL U5566 ( .A(n7154), .B(n7288), .C(n7099), .D(n7544), .Z(n625) );
  COND2XL U5567 ( .A(n7160), .B(n7290), .C(n7098), .D(n7546), .Z(n424) );
  COND2XL U5568 ( .A(n7138), .B(n7802), .C(n7132), .D(n8058), .Z(n423) );
  COND2XL U5569 ( .A(n7143), .B(n7703), .C(n7139), .D(n7447), .Z(n1435) );
  COND2XL U5570 ( .A(n7154), .B(n7319), .C(n7103), .D(n7575), .Z(n1436) );
  COND2XL U5571 ( .A(n7145), .B(n7702), .C(n7139), .D(n7446), .Z(n1032) );
  COND2XL U5572 ( .A(n7143), .B(n7667), .C(n7139), .D(n7411), .Z(n1336) );
  COND2XL U5573 ( .A(n7137), .B(n7828), .C(n7132), .D(n8084), .Z(n826) );
  COND2XL U5574 ( .A(n7146), .B(n7700), .C(n7139), .D(n7444), .Z(n824) );
  COND2XL U5575 ( .A(n7133), .B(n7825), .C(n7125), .D(n8081), .Z(n1767) );
  COND2XL U5576 ( .A(n7154), .B(n7314), .C(n7098), .D(n7570), .Z(n499) );
  COND2XL U5577 ( .A(n7138), .B(n7826), .C(n7131), .D(n8082), .Z(n500) );
  COND2XL U5578 ( .A(n7148), .B(n7698), .C(n7139), .D(n7442), .Z(n498) );
  COND2XL U5579 ( .A(n7144), .B(n7694), .C(n7139), .D(n7438), .Z(n1159) );
  COND2XL U5580 ( .A(n7137), .B(n7796), .C(n7132), .D(n8052), .Z(n802) );
  COND2XL U5581 ( .A(n7147), .B(n7668), .C(n7139), .D(n7412), .Z(n800) );
  COND2XL U5582 ( .A(n7137), .B(n7824), .C(n7129), .D(n8080), .Z(n727) );
  COND2XL U5583 ( .A(n7147), .B(n7696), .C(n7139), .D(n7440), .Z(n725) );
  COND2XL U5584 ( .A(n7145), .B(n7670), .C(n7139), .D(n7414), .Z(n1008) );
  COND2XL U5585 ( .A(n7149), .B(n7722), .C(n7139), .D(n7466), .Z(n438) );
  COND2XL U5586 ( .A(n7138), .B(n7850), .C(n7131), .D(n8106), .Z(n440) );
  COND2XL U5587 ( .A(n7148), .B(n7690), .C(n7139), .D(n7434), .Z(n464) );
  COND2XL U5588 ( .A(n7138), .B(n7818), .C(n7131), .D(n8074), .Z(n466) );
  COND2XL U5589 ( .A(n7146), .B(n7684), .C(n7139), .D(n7428), .Z(n866) );
  COND2XL U5590 ( .A(n7158), .B(n7300), .C(n7100), .D(n7556), .Z(n867) );
  COND2XL U5591 ( .A(n7156), .B(n7334), .C(n7101), .D(n7590), .Z(n1049) );
  COND2XL U5592 ( .A(n7145), .B(n7718), .C(n7139), .D(n7462), .Z(n1048) );
  COND2XL U5593 ( .A(n7156), .B(n7302), .C(n7101), .D(n7558), .Z(n1075) );
  COND2XL U5594 ( .A(n7145), .B(n7686), .C(n7139), .D(n7430), .Z(n1074) );
  COND2XL U5595 ( .A(n7123), .B(n7941), .C(n7161), .D(n8197), .Z(n1877) );
  COND2XL U5596 ( .A(n7140), .B(n7685), .C(n7139), .D(n7429), .Z(n1878) );
  COND2XL U5597 ( .A(n7133), .B(n7813), .C(n7124), .D(n8069), .Z(n1880) );
  COND2XL U5598 ( .A(n7123), .B(n7973), .C(n7161), .D(n8229), .Z(n1851) );
  COND2XL U5599 ( .A(n7140), .B(n7717), .C(n7139), .D(n7461), .Z(n1852) );
  COND2XL U5600 ( .A(n7133), .B(n7845), .C(n7124), .D(n8101), .Z(n1854) );
  COND2XL U5601 ( .A(n7137), .B(n7808), .C(n7132), .D(n8064), .Z(n769) );
  COND2XL U5602 ( .A(n7159), .B(n7296), .C(n7100), .D(n7552), .Z(n768) );
  COND2XL U5603 ( .A(n7147), .B(n7680), .C(n7139), .D(n7424), .Z(n767) );
  COND2XL U5604 ( .A(n7147), .B(n7720), .C(n7139), .D(n7464), .Z(n639) );
  COND2XL U5605 ( .A(n7147), .B(n7688), .C(n7139), .D(n7432), .Z(n665) );
  COND2XL U5606 ( .A(n7154), .B(n7304), .C(n7099), .D(n7560), .Z(n666) );
  COND2XL U5607 ( .A(n7138), .B(n7842), .C(n7128), .D(n8098), .Z(n541) );
  COND2XL U5608 ( .A(n7148), .B(n7714), .C(n7139), .D(n7458), .Z(n539) );
  COND2XL U5609 ( .A(n7151), .B(n7330), .C(n7098), .D(n7586), .Z(n540) );
  COND2XL U5610 ( .A(n7144), .B(n7723), .C(n7139), .D(n7467), .Z(n1253) );
  COND2XL U5611 ( .A(n7144), .B(n7691), .C(n7139), .D(n7435), .Z(n1279) );
  COND2XL U5612 ( .A(n7143), .B(n7715), .C(n7139), .D(n7459), .Z(n1352) );
  COND2XL U5613 ( .A(n7143), .B(n7683), .C(n7139), .D(n7427), .Z(n1378) );
  COND2XL U5614 ( .A(n7138), .B(n7810), .C(n7128), .D(n8066), .Z(n567) );
  COND2XL U5615 ( .A(n7150), .B(n7298), .C(n7099), .D(n7554), .Z(n566) );
  COND2XL U5616 ( .A(n7148), .B(n7682), .C(n7139), .D(n7426), .Z(n565) );
  COND2XL U5617 ( .A(n7145), .B(n7710), .C(n7139), .D(n7454), .Z(n1102) );
  COND2XL U5618 ( .A(n7145), .B(n7678), .C(n7139), .D(n7422), .Z(n1128) );
  COND2XL U5619 ( .A(n7157), .B(n7324), .C(n7101), .D(n7580), .Z(n949) );
  COND2XL U5620 ( .A(n7146), .B(n7708), .C(n7139), .D(n7452), .Z(n948) );
  COND2XL U5621 ( .A(n7146), .B(n7676), .C(n7139), .D(n7420), .Z(n974) );
  COND2XL U5622 ( .A(n7140), .B(n7653), .C(n7139), .D(n7397), .Z(n1890) );
  COND2XL U5623 ( .A(n7137), .B(n7840), .C(n7132), .D(n8096), .Z(n755) );
  COND2XL U5624 ( .A(n7159), .B(n7328), .C(n7100), .D(n7584), .Z(n754) );
  COND2XL U5625 ( .A(n7147), .B(n7712), .C(n7139), .D(n7456), .Z(n753) );
  COND2XL U5626 ( .A(n7147), .B(n7656), .C(n7139), .D(n7400), .Z(n677) );
  COND2XL U5627 ( .A(n7159), .B(n7266), .C(n7099), .D(n7528), .Z(n678) );
  COND2XL U5628 ( .A(n7138), .B(n7874), .C(n7126), .D(n8130), .Z(n553) );
  COND2XL U5629 ( .A(n7148), .B(n7746), .C(n7139), .D(n7490), .Z(n551) );
  COND2XL U5630 ( .A(n7152), .B(n7362), .C(n7098), .D(n7618), .Z(n552) );
  COND2XL U5631 ( .A(n7144), .B(n7659), .C(n7139), .D(n7403), .Z(n1291) );
  COND2XL U5632 ( .A(n7143), .B(n7651), .C(n7139), .D(n7395), .Z(n1390) );
  COND2XL U5633 ( .A(n7145), .B(n7646), .C(n7139), .D(n7390), .Z(n1140) );
  COND2XL U5634 ( .A(n7143), .B(n7751), .C(n7139), .D(n7495), .Z(n1463) );
  COND2XL U5635 ( .A(n7154), .B(n7367), .C(n7104), .D(n7623), .Z(n1464) );
  COND2XL U5636 ( .A(n7148), .B(n7658), .C(n7139), .D(n7402), .Z(n476) );
  COND2XL U5637 ( .A(n7138), .B(n7786), .C(n7124), .D(n8042), .Z(n478) );
  COND2XL U5638 ( .A(n7157), .B(n7356), .C(n7101), .D(n7612), .Z(n961) );
  COND2XL U5639 ( .A(n7146), .B(n7740), .C(n7139), .D(n7484), .Z(n960) );
  COND2XL U5640 ( .A(n7145), .B(n7644), .C(n7139), .D(n7388), .Z(n986) );
  COND2XL U5641 ( .A(n7146), .B(n7652), .C(n7139), .D(n7396), .Z(n878) );
  COND2XL U5642 ( .A(n7157), .B(n7260), .C(n7100), .D(n7524), .Z(n879) );
  COND2XL U5643 ( .A(n7156), .B(n7262), .C(n7101), .D(n7526), .Z(n1087) );
  COND2XL U5644 ( .A(n7145), .B(n7654), .C(n7139), .D(n7398), .Z(n1086) );
  COND2XL U5645 ( .A(n32), .B(n33), .C(n34), .D(n35), .Z(n31) );
  COND2XL U5646 ( .A(n7140), .B(n7661), .C(n7139), .D(n7405), .Z(n1932) );
  CNR2XL U5647 ( .A(n1931), .B(n1932), .Z(n1917) );
  CANR2XL U5648 ( .A(n8295), .B(n318), .C(n8294), .D(n138), .Z(n1603) );
  CND2XL U5649 ( .A(buffer[902]), .B(n7093), .Z(n1808) );
  CND2XL U5650 ( .A(buffer[897]), .B(n7093), .Z(n384) );
  CND2XL U5651 ( .A(buffer[899]), .B(n7093), .Z(n596) );
  CND2XL U5652 ( .A(buffer[898]), .B(n7093), .Z(n1611) );
  CND2XL U5653 ( .A(buffer[900]), .B(n7093), .Z(n1408) );
  CND2XL U5654 ( .A(buffer[896]), .B(n7093), .Z(n1210) );
  CND2XL U5655 ( .A(buffer[904]), .B(n7093), .Z(n1309) );
  CND2XL U5656 ( .A(buffer[906]), .B(n7093), .Z(n1762) );
  CND2XL U5657 ( .A(buffer[909]), .B(n7093), .Z(n1156) );
  CND2XL U5658 ( .A(buffer[903]), .B(n7093), .Z(n797) );
  CND2XL U5659 ( .A(buffer[907]), .B(n7093), .Z(n694) );
  CND2XL U5660 ( .A(buffer[901]), .B(n7093), .Z(n1005) );
  COND2XL U5661 ( .A(n7159), .B(n7344), .C(n7099), .D(n7600), .Z(n700) );
  CND2XL U5662 ( .A(buffer[905]), .B(n7093), .Z(n495) );
  CANR2XL U5663 ( .A(buffer[393]), .B(n6149), .C(buffer[137]), .D(n387), .Z(
        n496) );
  COND2XL U5664 ( .A(n7161), .B(n8143), .C(n7160), .D(n7225), .Z(n79) );
  COND2XL U5665 ( .A(n7140), .B(n7631), .C(n7139), .D(n7375), .Z(n78) );
  COND2XL U5666 ( .A(n64), .B(n65), .C(n7263), .D(n67), .Z(n62) );
  CANR2XL U5667 ( .A(buffer[518]), .B(n40), .C(buffer[262]), .D(n7097), .Z(
        n234) );
  COND4CXL U5668 ( .A(n332), .B(rd_ptr[3]), .C(n374), .D(n8285), .Z(n373) );
  CANR2XL U5669 ( .A(buffer[520]), .B(n40), .C(buffer[264]), .D(n7097), .Z(
        n191) );
  CANR2XL U5670 ( .A(buffer[521]), .B(n40), .C(buffer[265]), .D(n7097), .Z(
        n169) );
  CANR2XL U5671 ( .A(n3162), .B(n8297), .C(buffer[780]), .D(n7095), .Z(n1519)
         );
  CANR2XL U5672 ( .A(n8297), .B(buffer[263]), .C(n7095), .D(buffer[775]), .Z(
        n794) );
  CANR2XL U5673 ( .A(buffer[260]), .B(n8297), .C(buffer[772]), .D(n7095), .Z(
        n1405) );
  CANR2XL U5674 ( .A(buffer[262]), .B(n8297), .C(buffer[774]), .D(n7095), .Z(
        n1805) );
  CANR2XL U5675 ( .A(n8297), .B(buffer[261]), .C(n7095), .D(buffer[773]), .Z(
        n1002) );
  CANR2XL U5676 ( .A(buffer[258]), .B(n8297), .C(buffer[770]), .D(n7095), .Z(
        n1608) );
  COND3XL U5677 ( .A(n7133), .B(n7884), .C(n940), .D(n941), .Z(n938) );
  COND3XL U5678 ( .A(n7133), .B(n7885), .C(n1951), .D(n1952), .Z(n1949) );
  CANR2XL U5679 ( .A(buffer[514]), .B(n7096), .C(n8306), .D(n324), .Z(n1607)
         );
  CANR2XL U5680 ( .A(buffer[516]), .B(n7096), .C(n8306), .D(n277), .Z(n1404)
         );
  COND2XL U5681 ( .A(rd_ptr[2]), .B(n289), .C(n8290), .D(n155), .Z(n245) );
  CANR2XL U5682 ( .A(buffer[525]), .B(n40), .C(buffer[269]), .D(n7097), .Z(n27) );
  CANR2XL U5683 ( .A(n8297), .B(buffer[259]), .C(n7095), .D(buffer[771]), .Z(
        n593) );
  CANR2XL U5684 ( .A(n7096), .B(buffer[513]), .C(n8301), .D(n340), .Z(n377) );
  CANR2XL U5685 ( .A(buffer[512]), .B(n7096), .C(n8301), .D(n363), .Z(n1206)
         );
  CANR2XL U5686 ( .A(buffer[514]), .B(n40), .C(buffer[258]), .D(n7097), .Z(
        n322) );
  CANR2XL U5687 ( .A(n2847), .B(n7095), .C(n2846), .D(n7096), .Z(n899) );
  CANR2XL U5688 ( .A(n2384), .B(n7095), .C(n2383), .D(n7096), .Z(n1911) );
  CIVX1 U5689 ( .A(n239), .Z(n7208) );
  CANR2XL U5690 ( .A(buffer[512]), .B(n40), .C(buffer[256]), .D(n7097), .Z(
        n360) );
  CANR2XL U5691 ( .A(n8297), .B(buffer[269]), .C(n7095), .D(buffer[781]), .Z(
        n1153) );
  CANR2XL U5692 ( .A(buffer[517]), .B(n40), .C(buffer[261]), .D(n7097), .Z(
        n253) );
  CANR2XL U5693 ( .A(n8303), .B(n256), .C(n8298), .D(n257), .Z(n250) );
  COND3XL U5694 ( .A(n8), .B(n221), .C(n222), .D(n223), .Z(n3182) );
  COND3XL U5695 ( .A(n8), .B(n149), .C(n150), .D(n151), .Z(n3179) );
  CANR2XL U5696 ( .A(buffer[519]), .B(n40), .C(buffer[263]), .D(n7097), .Z(
        n215) );
  CANR2XL U5697 ( .A(buffer[516]), .B(n40), .C(buffer[260]), .D(n7097), .Z(
        n275) );
  CANR2XL U5698 ( .A(buffer[513]), .B(n40), .C(buffer[257]), .D(n7097), .Z(
        n338) );
  CANR2XL U5699 ( .A(buffer[515]), .B(n40), .C(buffer[259]), .D(n7097), .Z(
        n296) );
  CANR2XL U5700 ( .A(buffer[522]), .B(n40), .C(buffer[266]), .D(n7097), .Z(
        n147) );
  CANR2XL U5701 ( .A(n8297), .B(buffer[257]), .C(n7095), .D(buffer[769]), .Z(
        n378) );
  COND2XL U5702 ( .A(n7268), .B(n69), .C(n375), .D(n67), .Z(n374) );
  CANR2XL U5703 ( .A(n8306), .B(n362), .C(n8303), .D(n364), .Z(n1205) );
  CANR2XL U5704 ( .A(buffer[256]), .B(n8297), .C(buffer[768]), .D(n7095), .Z(
        n1207) );
  CANR2XL U5705 ( .A(n8297), .B(buffer[265]), .C(n7095), .D(buffer[777]), .Z(
        n491) );
  CANR2XL U5706 ( .A(n8297), .B(n8016), .C(n7095), .D(n7504), .Z(n691) );
  COND2XL U5707 ( .A(n8307), .B(n7759), .C(n75), .D(n76), .Z(n72) );
  COND2XL U5708 ( .A(n68), .B(n69), .C(n70), .D(n29), .Z(n61) );
  CND2XL U5709 ( .A(\add_121/carry [8]), .B(rd_ptr[8]), .Z(n6159) );
  CND2XL U5710 ( .A(n344), .B(n345), .Z(n3188) );
  CANR2XL U5711 ( .A(n7171), .B(n343), .C(n4285), .D(n7092), .Z(n344) );
  CANR2XL U5712 ( .A(buffer[266]), .B(n8297), .C(buffer[778]), .D(n7095), .Z(
        n1759) );
  COND3XL U5713 ( .A(n239), .B(n8), .C(n240), .D(n241), .Z(n3183) );
  CIVX1 U5714 ( .A(n49), .Z(n7224) );
  CNR3XL U5715 ( .A(wrt_ptr[2]), .B(wrt_ptr[3]), .C(n7221), .Z(n2061) );
  CNR3XL U5716 ( .A(wrt_ptr[1]), .B(wrt_ptr[3]), .C(n7222), .Z(n2082) );
  CNR3XL U5717 ( .A(n7222), .B(wrt_ptr[3]), .C(n7221), .Z(n2087) );
  CNR3XL U5718 ( .A(wrt_ptr[2]), .B(wrt_ptr[3]), .C(wrt_ptr[1]), .Z(n2058) );
  CNR3X1 U5719 ( .A(wrt_ptr[0]), .B(wrt_ptr[4]), .C(n7174), .Z(n2062) );
  CNR3X1 U5720 ( .A(n7174), .B(wrt_ptr[4]), .C(n7220), .Z(n2057) );
  CIVX3 U5721 ( .A(rst), .Z(n7173) );
  CNR2X2 U5722 ( .A(n909), .B(n910), .Z(n6156) );
  CIVX1 U5723 ( .A(n6156), .Z(n6157) );
  COND2XL U5724 ( .A(n7146), .B(n7692), .C(n7139), .D(n7436), .Z(n911) );
  CDLY1XL U5725 ( .A(n382), .Z(n6158) );
  CIVX2 U5726 ( .A(n900), .Z(n8297) );
  CNIVX1 U5727 ( .A(n8309), .Z(n7101) );
  CND2X1 U5728 ( .A(n8298), .B(n4241), .Z(n900) );
  CNIVX1 U5729 ( .A(n8309), .Z(n7100) );
  CIVX2 U5730 ( .A(n120), .Z(n8304) );
  CIVX2 U5731 ( .A(n92), .Z(n8305) );
  CNIVX1 U5732 ( .A(n8309), .Z(n7106) );
  CNR2X1 U5733 ( .A(n7211), .B(n174), .Z(n172) );
  CNIVX1 U5734 ( .A(n80), .Z(n7166) );
  CNIVX1 U5735 ( .A(n84), .Z(n7140) );
  CIVX2 U5736 ( .A(n33), .Z(n8298) );
  CNIVX1 U5737 ( .A(n2007), .Z(n7111) );
  CND2X1 U5738 ( .A(n1248), .B(n1249), .Z(n185) );
  CANR2X1 U5739 ( .A(n8298), .B(n1250), .C(n8303), .D(n1251), .Z(n1249) );
  CANR2X1 U5740 ( .A(n8306), .B(n1276), .C(n8301), .D(n1277), .Z(n1248) );
  CND2X1 U5741 ( .A(n835), .B(n836), .Z(n211) );
  CANR2X1 U5742 ( .A(n8298), .B(n837), .C(n8303), .D(n838), .Z(n836) );
  CANR2X1 U5743 ( .A(n8306), .B(n863), .C(n8301), .D(n864), .Z(n835) );
  CANR2X1 U5744 ( .A(n8301), .B(n237), .C(n8303), .D(n238), .Z(n1803) );
  CANR2X1 U5745 ( .A(n8301), .B(n218), .C(n8303), .D(n219), .Z(n792) );
  CANR2X1 U5746 ( .A(n8306), .B(n195), .C(n8303), .D(n197), .Z(n1303) );
  CANR2X1 U5747 ( .A(n8301), .B(n256), .C(n8303), .D(n257), .Z(n1000) );
  CANR2X1 U5748 ( .A(n8303), .B(n237), .C(n8298), .D(n238), .Z(n231) );
  CNIVX1 U5749 ( .A(n2008), .Z(n6169) );
  CND2X1 U5750 ( .A(n4240), .B(n8306), .Z(n120) );
  CANR2X1 U5751 ( .A(n8301), .B(n299), .C(n8298), .D(n300), .Z(n293) );
  CANR2X1 U5752 ( .A(n8303), .B(n278), .C(n8298), .D(n279), .Z(n272) );
  CND2X1 U5753 ( .A(n1703), .B(n1704), .Z(n138) );
  CANR2X1 U5754 ( .A(n8298), .B(n1705), .C(n8303), .D(n1706), .Z(n1704) );
  CANR2X1 U5755 ( .A(n8306), .B(n1731), .C(n8301), .D(n1732), .Z(n1703) );
  CND2X1 U5756 ( .A(n1649), .B(n1650), .Z(n137) );
  CANR2X1 U5757 ( .A(n8298), .B(n1651), .C(n8303), .D(n1652), .Z(n1650) );
  CANR2X1 U5758 ( .A(n8306), .B(n1677), .C(n8301), .D(n1678), .Z(n1649) );
  CNIVX1 U5759 ( .A(n391), .Z(n7096) );
  CNR2X1 U5760 ( .A(n33), .B(n7149), .Z(n391) );
  CND2X1 U5761 ( .A(n1097), .B(n1098), .Z(n44) );
  CANR2X1 U5762 ( .A(n8298), .B(n1099), .C(n8303), .D(n1100), .Z(n1098) );
  CANR2X1 U5763 ( .A(n8306), .B(n1125), .C(n8301), .D(n1126), .Z(n1097) );
  CND2X1 U5764 ( .A(n1043), .B(n1044), .Z(n46) );
  CANR2X1 U5765 ( .A(n8298), .B(n1045), .C(n8303), .D(n1046), .Z(n1044) );
  CANR2X1 U5766 ( .A(n8306), .B(n1071), .C(n8301), .D(n1072), .Z(n1043) );
  CAN2X1 U5767 ( .A(n1549), .B(n1550), .Z(n64) );
  CANR2X1 U5768 ( .A(n8303), .B(n1551), .C(n8298), .D(n1552), .Z(n1550) );
  CANR2X1 U5769 ( .A(n8306), .B(n1577), .C(n8301), .D(n1578), .Z(n1549) );
  CND2X1 U5770 ( .A(n1847), .B(n1848), .Z(n230) );
  CANR2X1 U5771 ( .A(n8298), .B(n1849), .C(n8303), .D(n1850), .Z(n1848) );
  CANR2X1 U5772 ( .A(n8306), .B(n1875), .C(n8301), .D(n1876), .Z(n1847) );
  CND2X1 U5773 ( .A(n1347), .B(n1348), .Z(n187) );
  CANR2X1 U5774 ( .A(n8298), .B(n1349), .C(n8303), .D(n1350), .Z(n1348) );
  CANR2X1 U5775 ( .A(n8306), .B(n1375), .C(n8301), .D(n1376), .Z(n1347) );
  CND2X1 U5776 ( .A(n433), .B(n434), .Z(n159) );
  CANR2X1 U5777 ( .A(n8298), .B(n435), .C(n8303), .D(n436), .Z(n434) );
  CANR2X1 U5778 ( .A(n8306), .B(n461), .C(n8301), .D(n462), .Z(n433) );
  CND2X1 U5779 ( .A(n634), .B(n635), .Z(n114) );
  CANR2X1 U5780 ( .A(n8298), .B(n636), .C(n8303), .D(n637), .Z(n635) );
  CANR2X1 U5781 ( .A(n8306), .B(n662), .C(n8301), .D(n663), .Z(n634) );
  CNIVX1 U5782 ( .A(n80), .Z(n7165) );
  CNIVX1 U5783 ( .A(n80), .Z(n7162) );
  CNIVX1 U5784 ( .A(n80), .Z(n7164) );
  CNIVX1 U5785 ( .A(n390), .Z(n7095) );
  CNIVX1 U5786 ( .A(n381), .Z(n7094) );
  CNIVX1 U5787 ( .A(n80), .Z(n7161) );
  CND2X1 U5788 ( .A(n152), .B(n175), .Z(n149) );
  CND2X1 U5789 ( .A(n736), .B(n737), .Z(n115) );
  CANR2X1 U5790 ( .A(n8306), .B(n764), .C(n8301), .D(n765), .Z(n736) );
  CANR2X1 U5791 ( .A(n8303), .B(n738), .C(n8298), .D(n739), .Z(n737) );
  CNIVX1 U5792 ( .A(n80), .Z(n7167) );
  CND2X1 U5793 ( .A(n534), .B(n535), .Z(n160) );
  CANR2X1 U5794 ( .A(n8306), .B(n562), .C(n8301), .D(n563), .Z(n534) );
  CANR2X1 U5795 ( .A(n8298), .B(n536), .C(n8303), .D(n537), .Z(n535) );
  CNIVX1 U5796 ( .A(n80), .Z(n7163) );
  CND2X1 U5797 ( .A(n1446), .B(n1447), .Z(n271) );
  CANR2X1 U5798 ( .A(n8306), .B(n1474), .C(n8301), .D(n1475), .Z(n1446) );
  CANR2X1 U5799 ( .A(n8298), .B(n1448), .C(n8303), .D(n1449), .Z(n1447) );
  COND1XL U5800 ( .A(n7210), .B(n178), .C(n10), .Z(n152) );
  CNR2X1 U5801 ( .A(n7210), .B(n7217), .Z(n174) );
  CNIVX1 U5802 ( .A(n2008), .Z(n6166) );
  CNIVX1 U5803 ( .A(n2008), .Z(n6167) );
  CNIVX1 U5804 ( .A(n2008), .Z(n6168) );
  CND2X1 U5805 ( .A(n7216), .B(n7210), .Z(n310) );
  CIVX2 U5806 ( .A(n14), .Z(n8285) );
  CNIVX1 U5807 ( .A(n2132), .Z(n6706) );
  CNIVX1 U5808 ( .A(n2134), .Z(n6679) );
  CNIVX1 U5809 ( .A(n2137), .Z(n6652) );
  CNIVX1 U5810 ( .A(n2132), .Z(n6704) );
  CNIVX1 U5811 ( .A(n2132), .Z(n6705) );
  CNIVX1 U5812 ( .A(n2134), .Z(n6677) );
  CNIVX1 U5813 ( .A(n2134), .Z(n6678) );
  CNIVX1 U5814 ( .A(n2137), .Z(n6650) );
  CNIVX1 U5815 ( .A(n2137), .Z(n6651) );
  COND1XL U5816 ( .A(n7219), .B(n7210), .C(n172), .Z(n203) );
  CNIVX1 U5817 ( .A(n2132), .Z(n6707) );
  CNIVX1 U5818 ( .A(n2134), .Z(n6680) );
  CNIVX1 U5819 ( .A(n2137), .Z(n6653) );
  CNIVX1 U5820 ( .A(n2056), .Z(n7066) );
  CNIVX1 U5821 ( .A(n2060), .Z(n7036) );
  CNIVX1 U5822 ( .A(n2064), .Z(n7006) );
  CNIVX1 U5823 ( .A(n2067), .Z(n6976) );
  CNIVX1 U5824 ( .A(n2084), .Z(n6946) );
  CNIVX1 U5825 ( .A(n2086), .Z(n6916) );
  CNIVX1 U5826 ( .A(n2089), .Z(n6886) );
  CNIVX1 U5827 ( .A(n2094), .Z(n6856) );
  CNIVX1 U5828 ( .A(n2109), .Z(n6826) );
  CNIVX1 U5829 ( .A(n2111), .Z(n6796) );
  CNIVX1 U5830 ( .A(n2114), .Z(n6766) );
  CNIVX1 U5831 ( .A(n2117), .Z(n6736) );
  CNIVX1 U5832 ( .A(n2141), .Z(n6625) );
  CNIVX1 U5833 ( .A(n2157), .Z(n6595) );
  CNIVX1 U5834 ( .A(n2160), .Z(n6565) );
  CNIVX1 U5835 ( .A(n2162), .Z(n6535) );
  CNIVX1 U5836 ( .A(n2165), .Z(n6505) );
  CNIVX1 U5837 ( .A(n2169), .Z(n6475) );
  CNIVX1 U5838 ( .A(n2172), .Z(n6445) );
  CNIVX1 U5839 ( .A(n2174), .Z(n6415) );
  CNIVX1 U5840 ( .A(n2177), .Z(n6385) );
  CNIVX1 U5841 ( .A(n2192), .Z(n6355) );
  CNIVX1 U5842 ( .A(n2194), .Z(n6325) );
  CNIVX1 U5843 ( .A(n2196), .Z(n6295) );
  CNIVX1 U5844 ( .A(n2199), .Z(n6265) );
  CNIVX1 U5845 ( .A(n2215), .Z(n6235) );
  CNIVX1 U5846 ( .A(n2217), .Z(n6205) );
  CNIVX1 U5847 ( .A(n2219), .Z(n6175) );
  CNIVX1 U5848 ( .A(n2056), .Z(n7065) );
  CNIVX1 U5849 ( .A(n2060), .Z(n7035) );
  CNIVX1 U5850 ( .A(n2064), .Z(n7005) );
  CNIVX1 U5851 ( .A(n2067), .Z(n6975) );
  CNIVX1 U5852 ( .A(n2084), .Z(n6945) );
  CNIVX1 U5853 ( .A(n2086), .Z(n6915) );
  CNIVX1 U5854 ( .A(n2089), .Z(n6885) );
  CNIVX1 U5855 ( .A(n2094), .Z(n6855) );
  CNIVX1 U5856 ( .A(n2109), .Z(n6825) );
  CNIVX1 U5857 ( .A(n2111), .Z(n6795) );
  CNIVX1 U5858 ( .A(n2114), .Z(n6765) );
  CNIVX1 U5859 ( .A(n2117), .Z(n6735) );
  CNIVX1 U5860 ( .A(n2141), .Z(n6624) );
  CNIVX1 U5861 ( .A(n2157), .Z(n6594) );
  CNIVX1 U5862 ( .A(n2160), .Z(n6564) );
  CNIVX1 U5863 ( .A(n2162), .Z(n6534) );
  CNIVX1 U5864 ( .A(n2165), .Z(n6504) );
  CNIVX1 U5865 ( .A(n2169), .Z(n6474) );
  CNIVX1 U5866 ( .A(n2172), .Z(n6444) );
  CNIVX1 U5867 ( .A(n2174), .Z(n6414) );
  CNIVX1 U5868 ( .A(n2177), .Z(n6384) );
  CNIVX1 U5869 ( .A(n2192), .Z(n6354) );
  CNIVX1 U5870 ( .A(n2194), .Z(n6324) );
  CNIVX1 U5871 ( .A(n2196), .Z(n6294) );
  CNIVX1 U5872 ( .A(n2199), .Z(n6264) );
  CNIVX1 U5873 ( .A(n2215), .Z(n6234) );
  CNIVX1 U5874 ( .A(n2217), .Z(n6204) );
  CNIVX1 U5875 ( .A(n2219), .Z(n6174) );
  CNIVX1 U5876 ( .A(n7061), .Z(n7062) );
  CNIVX1 U5877 ( .A(n7061), .Z(n7063) );
  CNIVX1 U5878 ( .A(n7061), .Z(n7064) );
  CNIVX1 U5879 ( .A(n7031), .Z(n7032) );
  CNIVX1 U5880 ( .A(n7031), .Z(n7033) );
  CNIVX1 U5881 ( .A(n7031), .Z(n7034) );
  CNIVX1 U5882 ( .A(n7001), .Z(n7002) );
  CNIVX1 U5883 ( .A(n7001), .Z(n7003) );
  CNIVX1 U5884 ( .A(n7001), .Z(n7004) );
  CNIVX1 U5885 ( .A(n6971), .Z(n6972) );
  CNIVX1 U5886 ( .A(n6971), .Z(n6973) );
  CNIVX1 U5887 ( .A(n6971), .Z(n6974) );
  CNIVX1 U5888 ( .A(n6941), .Z(n6942) );
  CNIVX1 U5889 ( .A(n6941), .Z(n6943) );
  CNIVX1 U5890 ( .A(n6941), .Z(n6944) );
  CNIVX1 U5891 ( .A(n6911), .Z(n6912) );
  CNIVX1 U5892 ( .A(n6911), .Z(n6913) );
  CNIVX1 U5893 ( .A(n6911), .Z(n6914) );
  CNIVX1 U5894 ( .A(n6881), .Z(n6882) );
  CNIVX1 U5895 ( .A(n6881), .Z(n6883) );
  CNIVX1 U5896 ( .A(n6881), .Z(n6884) );
  CNIVX1 U5897 ( .A(n6851), .Z(n6852) );
  CNIVX1 U5898 ( .A(n6851), .Z(n6853) );
  CNIVX1 U5899 ( .A(n6851), .Z(n6854) );
  CNIVX1 U5900 ( .A(n6821), .Z(n6822) );
  CNIVX1 U5901 ( .A(n6821), .Z(n6823) );
  CNIVX1 U5902 ( .A(n6821), .Z(n6824) );
  CNIVX1 U5903 ( .A(n6791), .Z(n6792) );
  CNIVX1 U5904 ( .A(n6791), .Z(n6793) );
  CNIVX1 U5905 ( .A(n6791), .Z(n6794) );
  CNIVX1 U5906 ( .A(n6761), .Z(n6762) );
  CNIVX1 U5907 ( .A(n6761), .Z(n6763) );
  CNIVX1 U5908 ( .A(n6761), .Z(n6764) );
  CNIVX1 U5909 ( .A(n6731), .Z(n6732) );
  CNIVX1 U5910 ( .A(n6731), .Z(n6733) );
  CNIVX1 U5911 ( .A(n6731), .Z(n6734) );
  CNIVX1 U5912 ( .A(n6620), .Z(n6621) );
  CNIVX1 U5913 ( .A(n6620), .Z(n6622) );
  CNIVX1 U5914 ( .A(n6620), .Z(n6623) );
  CNIVX1 U5915 ( .A(n6590), .Z(n6591) );
  CNIVX1 U5916 ( .A(n6590), .Z(n6592) );
  CNIVX1 U5917 ( .A(n6590), .Z(n6593) );
  CNIVX1 U5918 ( .A(n6560), .Z(n6561) );
  CNIVX1 U5919 ( .A(n6560), .Z(n6562) );
  CNIVX1 U5920 ( .A(n6560), .Z(n6563) );
  CNIVX1 U5921 ( .A(n6530), .Z(n6531) );
  CNIVX1 U5922 ( .A(n6530), .Z(n6532) );
  CNIVX1 U5923 ( .A(n6530), .Z(n6533) );
  CNIVX1 U5924 ( .A(n6500), .Z(n6501) );
  CNIVX1 U5925 ( .A(n6500), .Z(n6502) );
  CNIVX1 U5926 ( .A(n6500), .Z(n6503) );
  CNIVX1 U5927 ( .A(n6470), .Z(n6471) );
  CNIVX1 U5928 ( .A(n6470), .Z(n6472) );
  CNIVX1 U5929 ( .A(n6470), .Z(n6473) );
  CNIVX1 U5930 ( .A(n6440), .Z(n6441) );
  CNIVX1 U5931 ( .A(n6440), .Z(n6442) );
  CNIVX1 U5932 ( .A(n6440), .Z(n6443) );
  CNIVX1 U5933 ( .A(n6410), .Z(n6411) );
  CNIVX1 U5934 ( .A(n6410), .Z(n6412) );
  CNIVX1 U5935 ( .A(n6410), .Z(n6413) );
  CNIVX1 U5936 ( .A(n6380), .Z(n6381) );
  CNIVX1 U5937 ( .A(n6380), .Z(n6382) );
  CNIVX1 U5938 ( .A(n6380), .Z(n6383) );
  CNIVX1 U5939 ( .A(n6350), .Z(n6351) );
  CNIVX1 U5940 ( .A(n6350), .Z(n6352) );
  CNIVX1 U5941 ( .A(n6350), .Z(n6353) );
  CNIVX1 U5942 ( .A(n6320), .Z(n6321) );
  CNIVX1 U5943 ( .A(n6320), .Z(n6322) );
  CNIVX1 U5944 ( .A(n6320), .Z(n6323) );
  CNIVX1 U5945 ( .A(n6290), .Z(n6291) );
  CNIVX1 U5946 ( .A(n6290), .Z(n6292) );
  CNIVX1 U5947 ( .A(n6290), .Z(n6293) );
  CNIVX1 U5948 ( .A(n6260), .Z(n6261) );
  CNIVX1 U5949 ( .A(n6260), .Z(n6262) );
  CNIVX1 U5950 ( .A(n6260), .Z(n6263) );
  CNIVX1 U5951 ( .A(n6230), .Z(n6231) );
  CNIVX1 U5952 ( .A(n6230), .Z(n6232) );
  CNIVX1 U5953 ( .A(n6230), .Z(n6233) );
  CNIVX1 U5954 ( .A(n6200), .Z(n6201) );
  CNIVX1 U5955 ( .A(n6200), .Z(n6202) );
  CNIVX1 U5956 ( .A(n6200), .Z(n6203) );
  CNIVX1 U5957 ( .A(n6170), .Z(n6171) );
  CNIVX1 U5958 ( .A(n6170), .Z(n6172) );
  CNIVX1 U5959 ( .A(n6170), .Z(n6173) );
  CIVX2 U5960 ( .A(n67), .Z(n8291) );
  CNIVX1 U5961 ( .A(n2056), .Z(n7067) );
  CNIVX1 U5962 ( .A(n2060), .Z(n7037) );
  CNIVX1 U5963 ( .A(n2064), .Z(n7007) );
  CNIVX1 U5964 ( .A(n2067), .Z(n6977) );
  CNIVX1 U5965 ( .A(n2084), .Z(n6947) );
  CNIVX1 U5966 ( .A(n2086), .Z(n6917) );
  CNIVX1 U5967 ( .A(n2089), .Z(n6887) );
  CNIVX1 U5968 ( .A(n2094), .Z(n6857) );
  CNIVX1 U5969 ( .A(n2109), .Z(n6827) );
  CNIVX1 U5970 ( .A(n2111), .Z(n6797) );
  CNIVX1 U5971 ( .A(n2114), .Z(n6767) );
  CNIVX1 U5972 ( .A(n2117), .Z(n6737) );
  CNIVX1 U5973 ( .A(n2141), .Z(n6626) );
  CNIVX1 U5974 ( .A(n2157), .Z(n6596) );
  CNIVX1 U5975 ( .A(n2160), .Z(n6566) );
  CNIVX1 U5976 ( .A(n2162), .Z(n6536) );
  CNIVX1 U5977 ( .A(n2165), .Z(n6506) );
  CNIVX1 U5978 ( .A(n2169), .Z(n6476) );
  CNIVX1 U5979 ( .A(n2172), .Z(n6446) );
  CNIVX1 U5980 ( .A(n2174), .Z(n6416) );
  CNIVX1 U5981 ( .A(n2177), .Z(n6386) );
  CNIVX1 U5982 ( .A(n2192), .Z(n6356) );
  CNIVX1 U5983 ( .A(n2194), .Z(n6326) );
  CNIVX1 U5984 ( .A(n2196), .Z(n6296) );
  CNIVX1 U5985 ( .A(n2199), .Z(n6266) );
  CNIVX1 U5986 ( .A(n2215), .Z(n6236) );
  CNIVX1 U5987 ( .A(n2217), .Z(n6206) );
  CNIVX1 U5988 ( .A(n2219), .Z(n6176) );
  CNIVX1 U5989 ( .A(n2007), .Z(n7110) );
  CNIVX1 U5990 ( .A(n2007), .Z(n7109) );
  CNIVX1 U5991 ( .A(n2007), .Z(n7108) );
  COND11X1 U5992 ( .A(n116), .B(n117), .C(n118), .D(n8294), .Z(n112) );
  CND2X1 U5993 ( .A(n8308), .B(n8302), .Z(n33) );
  CNR2X1 U5994 ( .A(n76), .B(n7138), .Z(n40) );
  CNR2X1 U5995 ( .A(n33), .B(n8310), .Z(n380) );
  CNR4X1 U5996 ( .A(n510), .B(n511), .C(n512), .D(n513), .Z(n164) );
  COND2X1 U5997 ( .A(n7138), .B(n7858), .C(n7132), .D(n8114), .Z(n512) );
  CNR4X1 U5998 ( .A(n1171), .B(n1172), .C(n1173), .D(n1174), .Z(n32) );
  COND2X1 U5999 ( .A(n7117), .B(n7982), .C(n7165), .D(n8238), .Z(n1171) );
  CNR4X1 U6000 ( .A(n1777), .B(n1778), .C(n1779), .D(n1780), .Z(n142) );
  COND2X1 U6001 ( .A(n7141), .B(n7729), .C(n7139), .D(n7473), .Z(n1778) );
  COND2X1 U6002 ( .A(n7122), .B(n7985), .C(n7162), .D(n8241), .Z(n1777) );
  CNR4X1 U6003 ( .A(n522), .B(n523), .C(n524), .D(n525), .Z(n165) );
  COND2X1 U6004 ( .A(n7113), .B(n7922), .C(n7168), .D(n8178), .Z(n522) );
  COND2X1 U6005 ( .A(n7154), .B(n7282), .C(n7098), .D(n7538), .Z(n525) );
  CNR4X1 U6006 ( .A(n1183), .B(n1184), .C(n1185), .D(n1186), .Z(n34) );
  COND2X1 U6007 ( .A(n7117), .B(n7918), .C(n7164), .D(n8174), .Z(n1183) );
  CNR4X1 U6008 ( .A(n1789), .B(n1790), .C(n1791), .D(n1792), .Z(n143) );
  COND2X1 U6009 ( .A(n7141), .B(n7665), .C(n7139), .D(n7409), .Z(n1790) );
  COND2X1 U6010 ( .A(n7122), .B(n7921), .C(n7162), .D(n8177), .Z(n1789) );
  CNR4X1 U6011 ( .A(n1919), .B(n1920), .C(n1921), .D(n1922), .Z(n1918) );
  CANR11X1 U6012 ( .A(n7218), .B(n262), .C(n6162), .D(n263), .Z(n239) );
  CANR1XL U6013 ( .A(n264), .B(n265), .C(n7210), .Z(n263) );
  CANR2X1 U6014 ( .A(n6163), .B(n307), .C(n308), .D(n6162), .Z(n306) );
  CANR4CX1 U6015 ( .A(n8287), .B(n267), .C(n7244), .D(n7217), .Z(n308) );
  COND2X1 U6016 ( .A(n7147), .B(n7664), .C(n7139), .D(n7408), .Z(n715) );
  COND2X1 U6017 ( .A(n7142), .B(n7663), .C(n7139), .D(n7407), .Z(n1540) );
  COND2X1 U6018 ( .A(n7117), .B(n7920), .C(n7167), .D(n8176), .Z(n714) );
  COND2X1 U6019 ( .A(n7113), .B(n7984), .C(n7167), .D(n8240), .Z(n702) );
  COND2X1 U6020 ( .A(n7134), .B(n7823), .C(n7127), .D(n8079), .Z(n1506) );
  COND2X1 U6021 ( .A(n7120), .B(n7919), .C(n7163), .D(n8175), .Z(n1539) );
  COND2X1 U6022 ( .A(n7120), .B(n7983), .C(n7163), .D(n8239), .Z(n1527) );
  CNR4X1 U6023 ( .A(n1504), .B(n1505), .C(n1506), .D(n1507), .Z(n94) );
  COND2X1 U6024 ( .A(n7142), .B(n7695), .C(n7139), .D(n7439), .Z(n1505) );
  COND2X1 U6025 ( .A(n7120), .B(n7951), .C(n7163), .D(n8207), .Z(n1504) );
  COND2X1 U6026 ( .A(n7134), .B(n7791), .C(n7127), .D(n8047), .Z(n1538) );
  COND2X1 U6027 ( .A(n7134), .B(n7855), .C(n7127), .D(n8111), .Z(n1526) );
  COND2X1 U6028 ( .A(n7226), .B(n19), .C(n20), .D(n21), .Z(n11) );
  CANR11X1 U6029 ( .A(n26), .B(n27), .C(n28), .D(n29), .Z(n25) );
  CANR1X1 U6030 ( .A(n8293), .B(n269), .C(n270), .Z(n179) );
  COND2X1 U6031 ( .A(n29), .B(n68), .C(n65), .D(n7263), .Z(n270) );
  CND2X1 U6032 ( .A(n8286), .B(n129), .Z(n205) );
  COND3X1 U6033 ( .A(n179), .B(n16), .C(n180), .D(n181), .Z(n175) );
  CANR2X1 U6034 ( .A(n8288), .B(n60), .C(n8286), .D(n105), .Z(n181) );
  CANR2X1 U6035 ( .A(n226), .B(n8289), .C(n7237), .D(n8288), .Z(n264) );
  CANR11X1 U6036 ( .A(n6162), .B(n4243), .C(n6161), .D(n285), .Z(n258) );
  CIVX2 U6037 ( .A(n76), .Z(n8306) );
  CIVX2 U6038 ( .A(n93), .Z(n8303) );
  COND11X1 U6039 ( .A(n1905), .B(n1906), .C(n1907), .D(n8296), .Z(n1904) );
  COND1XL U6040 ( .A(n92), .B(n7533), .C(n1909), .Z(n1907) );
  COND11X1 U6041 ( .A(n893), .B(n894), .C(n895), .D(n8296), .Z(n892) );
  COND1XL U6042 ( .A(n92), .B(n7532), .C(n897), .Z(n895) );
  COND1XL U6043 ( .A(n8307), .B(n7788), .C(n899), .Z(n894) );
  CIVX2 U6044 ( .A(n35), .Z(n8301) );
  COND1XL U6045 ( .A(n1520), .B(n1521), .C(n8298), .Z(n1518) );
  COND2X1 U6046 ( .A(n7134), .B(n7887), .C(n7127), .D(n8143), .Z(n1521) );
  CANR2X1 U6047 ( .A(n39), .B(n361), .C(n8301), .D(n362), .Z(n358) );
  CANR2X1 U6048 ( .A(n39), .B(n235), .C(n8301), .D(n236), .Z(n232) );
  COND2X1 U6049 ( .A(n76), .B(n34), .C(n93), .D(n32), .Z(n1170) );
  COND2X1 U6050 ( .A(n76), .B(n143), .C(n93), .D(n142), .Z(n1776) );
  CND2X1 U6051 ( .A(n168), .B(n169), .Z(n161) );
  CND2X1 U6052 ( .A(n316), .B(n317), .Z(n198) );
  CANR2X1 U6053 ( .A(n8292), .B(n138), .C(n8291), .D(n318), .Z(n317) );
  CANR2X1 U6054 ( .A(n8294), .B(n148), .C(n8295), .D(n137), .Z(n316) );
  COND2X1 U6055 ( .A(n7115), .B(n8000), .C(n7167), .D(n8256), .Z(n740) );
  COND2X1 U6056 ( .A(n7112), .B(n7952), .C(n7167), .D(n8208), .Z(n724) );
  COND2X1 U6057 ( .A(n7116), .B(n7942), .C(n7165), .D(n8198), .Z(n1073) );
  COND2X1 U6058 ( .A(n7116), .B(n7974), .C(n7165), .D(n8230), .Z(n1047) );
  COND2X1 U6059 ( .A(n7113), .B(n7954), .C(n7168), .D(n8210), .Z(n497) );
  COND2X1 U6060 ( .A(n7113), .B(n7970), .C(n7167), .D(n8226), .Z(n538) );
  COND2X1 U6061 ( .A(n7113), .B(n8002), .C(n7167), .D(n8258), .Z(n550) );
  COND2X1 U6062 ( .A(n7113), .B(n7938), .C(n7167), .D(n8194), .Z(n564) );
  COND2X1 U6063 ( .A(n7113), .B(n7906), .C(n7167), .D(n8162), .Z(n576) );
  COND2X1 U6064 ( .A(n7118), .B(n8011), .C(n7164), .D(n8267), .Z(n1264) );
  COND2X1 U6065 ( .A(n7117), .B(n7998), .C(n7165), .D(n8254), .Z(n1113) );
  COND2X1 U6066 ( .A(n7116), .B(n7926), .C(n7165), .D(n8182), .Z(n1007) );
  COND2X1 U6067 ( .A(n7118), .B(n7931), .C(n7164), .D(n8187), .Z(n1236) );
  COND2X1 U6068 ( .A(n7118), .B(n7995), .C(n7164), .D(n8251), .Z(n1224) );
  COND2X1 U6069 ( .A(n7120), .B(n7935), .C(n7163), .D(n8191), .Z(n1579) );
  COND2X1 U6070 ( .A(n7120), .B(n7999), .C(n7163), .D(n8255), .Z(n1553) );
  COND2X1 U6071 ( .A(n7120), .B(n7967), .C(n7163), .D(n8223), .Z(n1565) );
  COND2X1 U6072 ( .A(n7116), .B(n7990), .C(n7165), .D(n8246), .Z(n1019) );
  COND2X1 U6073 ( .A(n7116), .B(n7958), .C(n7165), .D(n8214), .Z(n1031) );
  COND2X1 U6074 ( .A(n7112), .B(n8010), .C(n7168), .D(n8266), .Z(n449) );
  COND2X1 U6075 ( .A(n7116), .B(n7910), .C(n7165), .D(n8166), .Z(n1085) );
  COND2X1 U6076 ( .A(n7116), .B(n8006), .C(n7165), .D(n8262), .Z(n1059) );
  COND2X1 U6077 ( .A(n7122), .B(n8001), .C(n7162), .D(n8257), .Z(n1719) );
  COND2X1 U6078 ( .A(n7112), .B(n8003), .C(n7164), .D(n8259), .Z(n1363) );
  COND2X1 U6079 ( .A(n7121), .B(n8009), .C(n7162), .D(n8265), .Z(n1665) );
  COND2X1 U6080 ( .A(n7146), .B(n7724), .C(n7139), .D(n7468), .Z(n927) );
  COND2X1 U6081 ( .A(n7142), .B(n7655), .C(n7139), .D(n7399), .Z(n1489) );
  COND2X1 U6082 ( .A(n7145), .B(n7750), .C(n7139), .D(n7494), .Z(n1060) );
  COND2X1 U6083 ( .A(n7145), .B(n7742), .C(n7139), .D(n7486), .Z(n1114) );
  COND2X1 U6084 ( .A(n7141), .B(n7745), .C(n7139), .D(n7489), .Z(n1720) );
  COND2X1 U6085 ( .A(n7141), .B(n7753), .C(n7139), .D(n7497), .Z(n1666) );
  COND2X1 U6086 ( .A(n7142), .B(n7711), .C(n7139), .D(n7455), .Z(n1566) );
  COND2X1 U6087 ( .A(n7157), .B(n7340), .C(n7101), .D(n7596), .Z(n928) );
  COND2X1 U6088 ( .A(n7152), .B(n7289), .C(n7105), .D(n7545), .Z(n1615) );
  CND2X1 U6089 ( .A(n7173), .B(n6169), .Z(n2007) );
  COND2X1 U6090 ( .A(n7135), .B(n7863), .C(n7128), .D(n8119), .Z(n1425) );
  COND2X1 U6091 ( .A(n7135), .B(n7831), .C(n7128), .D(n8087), .Z(n1437) );
  COND2X1 U6092 ( .A(n7135), .B(n7847), .C(n7127), .D(n8103), .Z(n1453) );
  COND2X1 U6093 ( .A(n7135), .B(n7879), .C(n7127), .D(n8135), .Z(n1465) );
  COND2X1 U6094 ( .A(n7135), .B(n7815), .C(n7127), .D(n8071), .Z(n1479) );
  COND2X1 U6095 ( .A(n7134), .B(n7783), .C(n7127), .D(n8039), .Z(n1491) );
  COND2X1 U6096 ( .A(n7135), .B(n7799), .C(n7128), .D(n8055), .Z(n1413) );
  COND2X1 U6097 ( .A(n7135), .B(n7773), .C(n7130), .D(n8029), .Z(n1996) );
  COND2X1 U6098 ( .A(n7136), .B(n7878), .C(n7131), .D(n8134), .Z(n1062) );
  COND2X1 U6099 ( .A(n7135), .B(n7883), .C(n7129), .D(n8139), .Z(n1267) );
  COND2X1 U6100 ( .A(n7136), .B(n7870), .C(n7130), .D(n8126), .Z(n1116) );
  COND2X1 U6101 ( .A(n7134), .B(n7873), .C(n7125), .D(n8129), .Z(n1722) );
  COND2X1 U6102 ( .A(n7135), .B(n7875), .C(n7128), .D(n8131), .Z(n1366) );
  COND2X1 U6103 ( .A(n7134), .B(n7881), .C(n7125), .D(n8137), .Z(n1668) );
  COND2X1 U6104 ( .A(n7134), .B(n7839), .C(n7126), .D(n8095), .Z(n1568) );
  CND2X1 U6105 ( .A(n182), .B(n183), .Z(n60) );
  CANR2X1 U6106 ( .A(n8294), .B(n186), .C(n8295), .D(n187), .Z(n182) );
  CND4X1 U6107 ( .A(n188), .B(n189), .C(n190), .D(n191), .Z(n186) );
  CANR1XL U6108 ( .A(n8303), .B(n1915), .C(n1916), .Z(n1914) );
  COND2XL U6109 ( .A(n1917), .B(n76), .C(n1918), .D(n35), .Z(n1916) );
  COND2X1 U6110 ( .A(n7141), .B(n7669), .C(n7139), .D(n7413), .Z(n1812) );
  COND2X1 U6111 ( .A(n7123), .B(n7925), .C(n7162), .D(n8181), .Z(n1811) );
  COND2X1 U6112 ( .A(n7112), .B(n7994), .C(n7168), .D(n8250), .Z(n409) );
  COND2X1 U6113 ( .A(n7135), .B(n7859), .C(n7129), .D(n8115), .Z(n1325) );
  COND2X1 U6114 ( .A(n7144), .B(n7739), .C(n7139), .D(n7483), .Z(n1225) );
  COND2X1 U6115 ( .A(n7142), .B(n7737), .C(n7139), .D(n7481), .Z(n1626) );
  COND2X1 U6116 ( .A(n7134), .B(n7865), .C(n7126), .D(n8121), .Z(n1628) );
  COND2X1 U6117 ( .A(n7121), .B(n7993), .C(n7162), .D(n8249), .Z(n1625) );
  COND2X1 U6118 ( .A(n7136), .B(n7835), .C(n7130), .D(n8091), .Z(n1215) );
  COND2X1 U6119 ( .A(n7118), .B(n7963), .C(n7164), .D(n8219), .Z(n1212) );
  COND2X1 U6120 ( .A(n7135), .B(n7803), .C(n7129), .D(n8059), .Z(n1238) );
  COND2X1 U6121 ( .A(n7112), .B(n7930), .C(n7168), .D(n8186), .Z(n421) );
  COND2X1 U6122 ( .A(n7135), .B(n7795), .C(n7128), .D(n8051), .Z(n1337) );
  COND2X1 U6123 ( .A(n7142), .B(n7705), .C(n7139), .D(n7449), .Z(n1638) );
  COND2X1 U6124 ( .A(n7134), .B(n7833), .C(n7126), .D(n8089), .Z(n1640) );
  COND2X1 U6125 ( .A(n7121), .B(n7961), .C(n7162), .D(n8217), .Z(n1637) );
  COND3X1 U6126 ( .A(n7240), .B(n69), .C(n135), .D(n136), .Z(n107) );
  CANR2X1 U6127 ( .A(n8291), .B(n137), .C(n8295), .D(n138), .Z(n136) );
  COND11X1 U6128 ( .A(n139), .B(n140), .C(n141), .D(n8294), .Z(n135) );
  CND2X1 U6129 ( .A(n247), .B(n248), .Z(n129) );
  CANR2X1 U6130 ( .A(n8294), .B(n23), .C(n8295), .D(n46), .Z(n247) );
  COND2X1 U6131 ( .A(n7149), .B(n7706), .C(n7139), .D(n7450), .Z(n393) );
  COND2X1 U6132 ( .A(n7148), .B(n7704), .C(n7139), .D(n7448), .Z(n599) );
  COND2X1 U6133 ( .A(n7142), .B(n7673), .C(n7139), .D(n7417), .Z(n1614) );
  COND2X1 U6134 ( .A(n7134), .B(n7801), .C(n7126), .D(n8057), .Z(n1616) );
  COND2X1 U6135 ( .A(n7121), .B(n7929), .C(n7162), .D(n8185), .Z(n1613) );
  COND2X1 U6136 ( .A(n7154), .B(n7287), .C(n7103), .D(n7543), .Z(n1412) );
  COND2X1 U6137 ( .A(n7143), .B(n7671), .C(n7139), .D(n7415), .Z(n1411) );
  COND2X1 U6138 ( .A(n7135), .B(n7827), .C(n7129), .D(n8083), .Z(n1314) );
  COND2X1 U6139 ( .A(n7121), .B(n7955), .C(n7164), .D(n8211), .Z(n1311) );
  COND2X1 U6140 ( .A(n7141), .B(n7697), .C(n7139), .D(n7441), .Z(n1765) );
  COND2X1 U6141 ( .A(n7122), .B(n7953), .C(n7162), .D(n8209), .Z(n1764) );
  COND2X1 U6142 ( .A(n7136), .B(n7822), .C(n7130), .D(n8078), .Z(n1161) );
  COND2X1 U6143 ( .A(n7117), .B(n7950), .C(n7165), .D(n8206), .Z(n1158) );
  CNIVX1 U6144 ( .A(n396), .Z(n7135) );
  CNIVX1 U6145 ( .A(n396), .Z(n7134) );
  COND2X1 U6146 ( .A(n7112), .B(n7946), .C(n7168), .D(n8202), .Z(n463) );
  COND2X1 U6147 ( .A(n7112), .B(n7978), .C(n7168), .D(n8234), .Z(n437) );
  COND2X1 U6148 ( .A(n7136), .B(n7814), .C(n7131), .D(n8070), .Z(n1076) );
  COND2X1 U6149 ( .A(n7136), .B(n7846), .C(n7131), .D(n8102), .Z(n1050) );
  COND2X1 U6150 ( .A(n7135), .B(n7819), .C(n7129), .D(n8075), .Z(n1281) );
  COND2X1 U6151 ( .A(n7118), .B(n7947), .C(n7164), .D(n8203), .Z(n1278) );
  COND2X1 U6152 ( .A(n7135), .B(n7851), .C(n7129), .D(n8107), .Z(n1255) );
  COND2X1 U6153 ( .A(n7118), .B(n7979), .C(n7164), .D(n8235), .Z(n1252) );
  COND2X1 U6154 ( .A(n7136), .B(n7806), .C(n7130), .D(n8062), .Z(n1130) );
  COND2X1 U6155 ( .A(n7117), .B(n7934), .C(n7165), .D(n8190), .Z(n1127) );
  COND2X1 U6156 ( .A(n7136), .B(n7838), .C(n7131), .D(n8094), .Z(n1104) );
  COND2X1 U6157 ( .A(n7117), .B(n7966), .C(n7165), .D(n8222), .Z(n1101) );
  COND2X1 U6158 ( .A(n7141), .B(n7681), .C(n7139), .D(n7425), .Z(n1734) );
  COND2X1 U6159 ( .A(n7134), .B(n7809), .C(n7125), .D(n8065), .Z(n1736) );
  COND2X1 U6160 ( .A(n7122), .B(n7937), .C(n7162), .D(n8193), .Z(n1733) );
  COND2X1 U6161 ( .A(n7141), .B(n7713), .C(n7139), .D(n7457), .Z(n1708) );
  COND2X1 U6162 ( .A(n7134), .B(n7841), .C(n7125), .D(n8097), .Z(n1710) );
  COND2X1 U6163 ( .A(n7122), .B(n7969), .C(n7162), .D(n8225), .Z(n1707) );
  COND2X1 U6164 ( .A(n7135), .B(n7811), .C(n7128), .D(n8067), .Z(n1380) );
  COND2X1 U6165 ( .A(n7135), .B(n7843), .C(n7128), .D(n8099), .Z(n1354) );
  COND2X1 U6166 ( .A(n7141), .B(n7689), .C(n7139), .D(n7433), .Z(n1680) );
  COND2X1 U6167 ( .A(n7134), .B(n7817), .C(n7125), .D(n8073), .Z(n1682) );
  COND2X1 U6168 ( .A(n7121), .B(n7945), .C(n7162), .D(n8201), .Z(n1679) );
  COND2X1 U6169 ( .A(n7142), .B(n7721), .C(n7139), .D(n7465), .Z(n1654) );
  COND2X1 U6170 ( .A(n7134), .B(n7849), .C(n7126), .D(n8105), .Z(n1656) );
  COND2X1 U6171 ( .A(n7121), .B(n7977), .C(n7162), .D(n8233), .Z(n1653) );
  COND2X1 U6172 ( .A(n7142), .B(n7679), .C(n7139), .D(n7423), .Z(n1580) );
  COND2X1 U6173 ( .A(n7134), .B(n7807), .C(n7126), .D(n8063), .Z(n1582) );
  COND2X1 U6174 ( .A(n7142), .B(n7743), .C(n7139), .D(n7487), .Z(n1554) );
  COND2X1 U6175 ( .A(n7134), .B(n7871), .C(n7126), .D(n8127), .Z(n1556) );
  COND2X1 U6176 ( .A(n7115), .B(n7932), .C(n7165), .D(n8188), .Z(n973) );
  COND2X1 U6177 ( .A(n7135), .B(n7787), .C(n7129), .D(n8043), .Z(n1293) );
  COND2X1 U6178 ( .A(n7118), .B(n7915), .C(n7164), .D(n8171), .Z(n1290) );
  COND2X1 U6179 ( .A(n7136), .B(n7774), .C(n7130), .D(n8030), .Z(n1142) );
  COND2X1 U6180 ( .A(n7117), .B(n7902), .C(n7165), .D(n8158), .Z(n1139) );
  COND2X1 U6181 ( .A(n7141), .B(n7649), .C(n7139), .D(n7393), .Z(n1746) );
  COND2X1 U6182 ( .A(n7134), .B(n7777), .C(n7125), .D(n8033), .Z(n1748) );
  COND2X1 U6183 ( .A(n7122), .B(n7905), .C(n7162), .D(n8161), .Z(n1745) );
  COND2X1 U6184 ( .A(n7135), .B(n7779), .C(n7128), .D(n8035), .Z(n1392) );
  COND2X1 U6185 ( .A(n7141), .B(n7657), .C(n7139), .D(n7401), .Z(n1692) );
  COND2X1 U6186 ( .A(n7134), .B(n7785), .C(n7125), .D(n8041), .Z(n1694) );
  COND2X1 U6187 ( .A(n7121), .B(n7913), .C(n7162), .D(n8169), .Z(n1691) );
  COND2X1 U6188 ( .A(n7142), .B(n7647), .C(n7139), .D(n7391), .Z(n1592) );
  COND2X1 U6189 ( .A(n7134), .B(n7775), .C(n7126), .D(n8031), .Z(n1594) );
  COND2X1 U6190 ( .A(n7120), .B(n7903), .C(n7163), .D(n8159), .Z(n1591) );
  COND2X1 U6191 ( .A(n7115), .B(n7900), .C(n7165), .D(n8156), .Z(n985) );
  COND2X1 U6192 ( .A(n7112), .B(n7914), .C(n7168), .D(n8170), .Z(n475) );
  COND2X1 U6193 ( .A(n7136), .B(n7782), .C(n7131), .D(n8038), .Z(n1088) );
  CND2X1 U6194 ( .A(n6163), .B(n243), .Z(n221) );
  CNIVX1 U6195 ( .A(n396), .Z(n7137) );
  CNR2X1 U6196 ( .A(n30), .B(n31), .Z(n28) );
  CNIVX1 U6197 ( .A(n396), .Z(n7136) );
  CNIVX1 U6198 ( .A(n396), .Z(n7133) );
  CND2X1 U6199 ( .A(n997), .B(n998), .Z(n288) );
  CANR2X1 U6200 ( .A(n8292), .B(n46), .C(n8291), .D(n999), .Z(n998) );
  CANR2X1 U6201 ( .A(n8295), .B(n249), .C(n8294), .D(n44), .Z(n997) );
  CND4X1 U6202 ( .A(n1000), .B(n1001), .C(n1002), .D(n1003), .Z(n999) );
  COND2X1 U6203 ( .A(n314), .B(n14), .C(n7245), .D(n19), .Z(n313) );
  CND2X1 U6204 ( .A(n310), .B(n370), .Z(n348) );
  CAN2X1 U6205 ( .A(n1603), .B(n1604), .Z(n1198) );
  CANR2X1 U6206 ( .A(n8292), .B(n137), .C(n8291), .D(n1605), .Z(n1604) );
  CND2X1 U6207 ( .A(n312), .B(n7244), .Z(n307) );
  CANR2X1 U6208 ( .A(n8288), .B(n198), .C(n8289), .D(n266), .Z(n312) );
  CANR2X1 U6209 ( .A(n8298), .B(n1953), .C(n8303), .D(n1954), .Z(n1903) );
  CANR2X1 U6210 ( .A(n8306), .B(n1979), .C(n8301), .D(n1980), .Z(n1902) );
  CNR2X1 U6211 ( .A(n920), .B(n921), .Z(n906) );
  CND2X1 U6212 ( .A(n2058), .B(n2062), .Z(n2008) );
  CNIVX1 U6213 ( .A(n41), .Z(n7097) );
  CANR2X1 U6214 ( .A(n8306), .B(n971), .C(n8301), .D(n972), .Z(n890) );
  CANR2X1 U6215 ( .A(n8298), .B(n945), .C(n8303), .D(n946), .Z(n891) );
  CAN2X1 U6216 ( .A(n167), .B(n380), .Z(n493) );
  CAN2X1 U6217 ( .A(n192), .B(n380), .Z(n1307) );
  COND2X1 U6218 ( .A(n76), .B(n165), .C(n93), .D(n164), .Z(n509) );
  CND2X1 U6219 ( .A(n8293), .B(n8296), .Z(n67) );
  CND2X1 U6220 ( .A(n6165), .B(n8284), .Z(n8) );
  COND2X1 U6221 ( .A(n8271), .B(n7110), .C(n6168), .D(n7194), .Z(n3212) );
  COND2X1 U6222 ( .A(n8267), .B(n7110), .C(n6166), .D(n7190), .Z(n3216) );
  COND2X1 U6223 ( .A(n8266), .B(n7110), .C(n6167), .D(n7189), .Z(n3217) );
  COND2X1 U6224 ( .A(n8265), .B(n7110), .C(n6166), .D(n7188), .Z(n3218) );
  COND2X1 U6225 ( .A(n8264), .B(n7110), .C(n6166), .D(n7187), .Z(n3219) );
  COND2X1 U6226 ( .A(n8263), .B(n7109), .C(n6168), .D(n7186), .Z(n3220) );
  COND2X1 U6227 ( .A(n8262), .B(n7109), .C(n6169), .D(n7185), .Z(n3221) );
  COND2X1 U6228 ( .A(n8261), .B(n7109), .C(n6167), .D(n7184), .Z(n3222) );
  COND2X1 U6229 ( .A(n8260), .B(n7109), .C(n6167), .D(n7183), .Z(n3223) );
  COND2X1 U6230 ( .A(n8259), .B(n7109), .C(n6166), .D(n7182), .Z(n3224) );
  COND2X1 U6231 ( .A(n8258), .B(n7109), .C(n6167), .D(n7181), .Z(n3225) );
  COND2X1 U6232 ( .A(n8257), .B(n7109), .C(n6168), .D(n7180), .Z(n3226) );
  COND2X1 U6233 ( .A(n8256), .B(n7109), .C(n6168), .D(n7179), .Z(n3227) );
  COND2X1 U6234 ( .A(n8255), .B(n7109), .C(n6168), .D(n7178), .Z(n3228) );
  COND2X1 U6235 ( .A(n8254), .B(n7109), .C(n6169), .D(n7177), .Z(n3229) );
  COND2X1 U6236 ( .A(n8253), .B(n7109), .C(n6169), .D(n7176), .Z(n3230) );
  COND2X1 U6237 ( .A(n8252), .B(n7109), .C(n6169), .D(n7175), .Z(n3231) );
  COND2X1 U6238 ( .A(n8251), .B(n7071), .C(n7206), .D(n7062), .Z(n3232) );
  COND2X1 U6239 ( .A(n8250), .B(n7072), .C(n7205), .D(n7063), .Z(n3233) );
  COND2X1 U6240 ( .A(n8249), .B(n7073), .C(n7204), .D(n7062), .Z(n3234) );
  COND2X1 U6241 ( .A(n8248), .B(n7074), .C(n7203), .D(n7063), .Z(n3235) );
  COND2X1 U6242 ( .A(n8247), .B(n7075), .C(n7202), .D(n7064), .Z(n3236) );
  COND2X1 U6243 ( .A(n8246), .B(n7076), .C(n7201), .D(n7062), .Z(n3237) );
  COND2X1 U6244 ( .A(n8245), .B(n7078), .C(n7200), .D(n7064), .Z(n3238) );
  COND2X1 U6245 ( .A(n8244), .B(n7079), .C(n7199), .D(n7065), .Z(n3239) );
  COND2X1 U6246 ( .A(n8243), .B(n7080), .C(n7198), .D(n7065), .Z(n3240) );
  COND2X1 U6247 ( .A(n8242), .B(n7081), .C(n7197), .D(n7066), .Z(n3241) );
  COND2X1 U6248 ( .A(n8241), .B(n7082), .C(n7196), .D(n7067), .Z(n3242) );
  COND2X1 U6249 ( .A(n8240), .B(n7083), .C(n7195), .D(n7063), .Z(n3243) );
  COND2X1 U6250 ( .A(n8239), .B(n7085), .C(n7194), .D(n7066), .Z(n3244) );
  COND2X1 U6251 ( .A(n8238), .B(n7086), .C(n7193), .D(n7067), .Z(n3245) );
  COND2X1 U6252 ( .A(n8237), .B(n7082), .C(n7192), .D(n7062), .Z(n3246) );
  COND2X1 U6253 ( .A(n8236), .B(n7083), .C(n7191), .D(n7063), .Z(n3247) );
  COND2X1 U6254 ( .A(n8235), .B(n7085), .C(n7190), .D(n7064), .Z(n3248) );
  COND2X1 U6255 ( .A(n8234), .B(n7086), .C(n7189), .D(n7064), .Z(n3249) );
  COND2X1 U6256 ( .A(n8233), .B(n7087), .C(n7188), .D(n7062), .Z(n3250) );
  COND2X1 U6257 ( .A(n8232), .B(n7088), .C(n7187), .D(n7063), .Z(n3251) );
  COND2X1 U6258 ( .A(n8231), .B(n7089), .C(n7186), .D(n7065), .Z(n3252) );
  COND2X1 U6259 ( .A(n8230), .B(n7090), .C(n7185), .D(n7066), .Z(n3253) );
  COND2X1 U6260 ( .A(n8229), .B(n7071), .C(n7184), .D(n7067), .Z(n3254) );
  COND2X1 U6261 ( .A(n8228), .B(n7072), .C(n7183), .D(n7065), .Z(n3255) );
  COND2X1 U6262 ( .A(n8227), .B(n7073), .C(n7182), .D(n7064), .Z(n3256) );
  COND2X1 U6263 ( .A(n8226), .B(n7074), .C(n7181), .D(n7065), .Z(n3257) );
  COND2X1 U6264 ( .A(n8225), .B(n7075), .C(n7180), .D(n7062), .Z(n3258) );
  COND2X1 U6265 ( .A(n8224), .B(n7076), .C(n7179), .D(n7063), .Z(n3259) );
  COND2X1 U6266 ( .A(n8223), .B(n7078), .C(n7178), .D(n7064), .Z(n3260) );
  COND2X1 U6267 ( .A(n8222), .B(n7079), .C(n7177), .D(n7066), .Z(n3261) );
  COND2X1 U6268 ( .A(n8221), .B(n7080), .C(n7176), .D(n7066), .Z(n3262) );
  COND2X1 U6269 ( .A(n8220), .B(n7081), .C(n7175), .D(n7067), .Z(n3263) );
  COND2X1 U6270 ( .A(n8219), .B(n7041), .C(n7206), .D(n7032), .Z(n3264) );
  COND2X1 U6271 ( .A(n8218), .B(n7042), .C(n7205), .D(n7033), .Z(n3265) );
  COND2X1 U6272 ( .A(n8217), .B(n7043), .C(n7204), .D(n7032), .Z(n3266) );
  COND2X1 U6273 ( .A(n8216), .B(n7044), .C(n7203), .D(n7033), .Z(n3267) );
  COND2X1 U6274 ( .A(n8215), .B(n7045), .C(n7202), .D(n7034), .Z(n3268) );
  COND2X1 U6275 ( .A(n8214), .B(n7046), .C(n7201), .D(n7032), .Z(n3269) );
  COND2X1 U6276 ( .A(n8213), .B(n7048), .C(n7200), .D(n7034), .Z(n3270) );
  COND2X1 U6277 ( .A(n8212), .B(n7049), .C(n7199), .D(n7035), .Z(n3271) );
  COND2X1 U6278 ( .A(n8211), .B(n7050), .C(n7198), .D(n7035), .Z(n3272) );
  COND2X1 U6279 ( .A(n8210), .B(n7051), .C(n7197), .D(n7036), .Z(n3273) );
  COND2X1 U6280 ( .A(n8209), .B(n7052), .C(n7196), .D(n7037), .Z(n3274) );
  COND2X1 U6281 ( .A(n8208), .B(n7053), .C(n7195), .D(n7033), .Z(n3275) );
  COND2X1 U6282 ( .A(n8207), .B(n7055), .C(n7194), .D(n7036), .Z(n3276) );
  COND2X1 U6283 ( .A(n8206), .B(n7056), .C(n7193), .D(n7037), .Z(n3277) );
  COND2X1 U6284 ( .A(n8205), .B(n7052), .C(n7192), .D(n7032), .Z(n3278) );
  COND2X1 U6285 ( .A(n8204), .B(n7053), .C(n7191), .D(n7033), .Z(n3279) );
  COND2X1 U6286 ( .A(n8203), .B(n7055), .C(n7190), .D(n7034), .Z(n3280) );
  COND2X1 U6287 ( .A(n8202), .B(n7056), .C(n7189), .D(n7034), .Z(n3281) );
  COND2X1 U6288 ( .A(n8201), .B(n7057), .C(n7188), .D(n7032), .Z(n3282) );
  COND2X1 U6289 ( .A(n8200), .B(n7058), .C(n7187), .D(n7033), .Z(n3283) );
  COND2X1 U6290 ( .A(n8199), .B(n7059), .C(n7186), .D(n7035), .Z(n3284) );
  COND2X1 U6291 ( .A(n8198), .B(n7060), .C(n7185), .D(n7036), .Z(n3285) );
  COND2X1 U6292 ( .A(n8197), .B(n7041), .C(n7184), .D(n7037), .Z(n3286) );
  COND2X1 U6293 ( .A(n8196), .B(n7042), .C(n7183), .D(n7035), .Z(n3287) );
  COND2X1 U6294 ( .A(n8195), .B(n7043), .C(n7182), .D(n7034), .Z(n3288) );
  COND2X1 U6295 ( .A(n8194), .B(n7044), .C(n7181), .D(n7035), .Z(n3289) );
  COND2X1 U6296 ( .A(n8193), .B(n7045), .C(n7180), .D(n7032), .Z(n3290) );
  COND2X1 U6297 ( .A(n8192), .B(n7046), .C(n7179), .D(n7033), .Z(n3291) );
  COND2X1 U6298 ( .A(n8191), .B(n7048), .C(n7178), .D(n7034), .Z(n3292) );
  COND2X1 U6299 ( .A(n8190), .B(n7049), .C(n7177), .D(n7036), .Z(n3293) );
  COND2X1 U6300 ( .A(n8189), .B(n7050), .C(n7176), .D(n7036), .Z(n3294) );
  COND2X1 U6301 ( .A(n8188), .B(n7051), .C(n7175), .D(n7037), .Z(n3295) );
  COND2X1 U6302 ( .A(n8187), .B(n7011), .C(n7206), .D(n7002), .Z(n3296) );
  COND2X1 U6303 ( .A(n8186), .B(n7012), .C(n7205), .D(n7003), .Z(n3297) );
  COND2X1 U6304 ( .A(n8185), .B(n7013), .C(n7204), .D(n7002), .Z(n3298) );
  COND2X1 U6305 ( .A(n8184), .B(n7014), .C(n7203), .D(n7003), .Z(n3299) );
  COND2X1 U6306 ( .A(n8183), .B(n7015), .C(n7202), .D(n7004), .Z(n3300) );
  COND2X1 U6307 ( .A(n8182), .B(n7016), .C(n7201), .D(n7002), .Z(n3301) );
  COND2X1 U6308 ( .A(n8181), .B(n7018), .C(n7200), .D(n7004), .Z(n3302) );
  COND2X1 U6309 ( .A(n8180), .B(n7019), .C(n7199), .D(n7005), .Z(n3303) );
  COND2X1 U6310 ( .A(n8179), .B(n7020), .C(n7198), .D(n7005), .Z(n3304) );
  COND2X1 U6311 ( .A(n8178), .B(n7021), .C(n7197), .D(n7006), .Z(n3305) );
  COND2X1 U6312 ( .A(n8177), .B(n7022), .C(n7196), .D(n7007), .Z(n3306) );
  COND2X1 U6313 ( .A(n8176), .B(n7023), .C(n7195), .D(n7003), .Z(n3307) );
  COND2X1 U6314 ( .A(n8175), .B(n7025), .C(n7194), .D(n7006), .Z(n3308) );
  COND2X1 U6315 ( .A(n8174), .B(n7026), .C(n7193), .D(n7007), .Z(n3309) );
  COND2X1 U6316 ( .A(n8173), .B(n7022), .C(n7192), .D(n7002), .Z(n3310) );
  COND2X1 U6317 ( .A(n8172), .B(n7023), .C(n7191), .D(n7003), .Z(n3311) );
  COND2X1 U6318 ( .A(n8171), .B(n7025), .C(n7190), .D(n7004), .Z(n3312) );
  COND2X1 U6319 ( .A(n8170), .B(n7026), .C(n7189), .D(n7004), .Z(n3313) );
  COND2X1 U6320 ( .A(n8169), .B(n7027), .C(n7188), .D(n7002), .Z(n3314) );
  COND2X1 U6321 ( .A(n8168), .B(n7028), .C(n7187), .D(n7003), .Z(n3315) );
  COND2X1 U6322 ( .A(n8167), .B(n7029), .C(n7186), .D(n7005), .Z(n3316) );
  COND2X1 U6323 ( .A(n8166), .B(n7030), .C(n7185), .D(n7006), .Z(n3317) );
  COND2X1 U6324 ( .A(n8165), .B(n7011), .C(n7184), .D(n7007), .Z(n3318) );
  COND2X1 U6325 ( .A(n8164), .B(n7012), .C(n7183), .D(n7005), .Z(n3319) );
  COND2X1 U6326 ( .A(n8163), .B(n7013), .C(n7182), .D(n7004), .Z(n3320) );
  COND2X1 U6327 ( .A(n8162), .B(n7014), .C(n7181), .D(n7005), .Z(n3321) );
  COND2X1 U6328 ( .A(n8161), .B(n7015), .C(n7180), .D(n7002), .Z(n3322) );
  COND2X1 U6329 ( .A(n8160), .B(n7016), .C(n7179), .D(n7003), .Z(n3323) );
  COND2X1 U6330 ( .A(n8159), .B(n7018), .C(n7178), .D(n7004), .Z(n3324) );
  COND2X1 U6331 ( .A(n8158), .B(n7019), .C(n7177), .D(n7006), .Z(n3325) );
  COND2X1 U6332 ( .A(n8157), .B(n7020), .C(n7176), .D(n7006), .Z(n3326) );
  COND2X1 U6333 ( .A(n8156), .B(n7021), .C(n7175), .D(n7007), .Z(n3327) );
  COND2X1 U6334 ( .A(n8139), .B(n6995), .C(n7190), .D(n6974), .Z(n3344) );
  COND2X1 U6335 ( .A(n8138), .B(n6996), .C(n7189), .D(n6974), .Z(n3345) );
  COND2X1 U6336 ( .A(n8137), .B(n6997), .C(n7188), .D(n6972), .Z(n3346) );
  COND2X1 U6337 ( .A(n8136), .B(n6998), .C(n7187), .D(n6973), .Z(n3347) );
  COND2X1 U6338 ( .A(n8135), .B(n6999), .C(n7186), .D(n6975), .Z(n3348) );
  COND2X1 U6339 ( .A(n8134), .B(n7000), .C(n7185), .D(n6976), .Z(n3349) );
  COND2X1 U6340 ( .A(n8133), .B(n6981), .C(n7184), .D(n6977), .Z(n3350) );
  COND2X1 U6341 ( .A(n8132), .B(n6982), .C(n7183), .D(n6975), .Z(n3351) );
  COND2X1 U6342 ( .A(n8131), .B(n6983), .C(n7182), .D(n6974), .Z(n3352) );
  COND2X1 U6343 ( .A(n8130), .B(n6984), .C(n7181), .D(n6975), .Z(n3353) );
  COND2X1 U6344 ( .A(n8129), .B(n6985), .C(n7180), .D(n6972), .Z(n3354) );
  COND2X1 U6345 ( .A(n8128), .B(n6986), .C(n7179), .D(n6973), .Z(n3355) );
  COND2X1 U6346 ( .A(n8127), .B(n6988), .C(n7178), .D(n6974), .Z(n3356) );
  COND2X1 U6347 ( .A(n8126), .B(n6989), .C(n7177), .D(n6976), .Z(n3357) );
  COND2X1 U6348 ( .A(n8125), .B(n6990), .C(n7176), .D(n6976), .Z(n3358) );
  COND2X1 U6349 ( .A(n8124), .B(n6991), .C(n7175), .D(n6977), .Z(n3359) );
  COND2X1 U6350 ( .A(n8123), .B(n6951), .C(n7206), .D(n6942), .Z(n3360) );
  COND2X1 U6351 ( .A(n8122), .B(n6952), .C(n7205), .D(n6943), .Z(n3361) );
  COND2X1 U6352 ( .A(n8121), .B(n6953), .C(n7204), .D(n6942), .Z(n3362) );
  COND2X1 U6353 ( .A(n8120), .B(n6954), .C(n7203), .D(n6943), .Z(n3363) );
  COND2X1 U6354 ( .A(n8119), .B(n6955), .C(n7202), .D(n6944), .Z(n3364) );
  COND2X1 U6355 ( .A(n8118), .B(n6956), .C(n7201), .D(n6942), .Z(n3365) );
  COND2X1 U6356 ( .A(n8117), .B(n6958), .C(n7200), .D(n6944), .Z(n3366) );
  COND2X1 U6357 ( .A(n8116), .B(n6959), .C(n7199), .D(n6945), .Z(n3367) );
  COND2X1 U6358 ( .A(n8115), .B(n6960), .C(n7198), .D(n6945), .Z(n3368) );
  COND2X1 U6359 ( .A(n8114), .B(n6961), .C(n7197), .D(n6946), .Z(n3369) );
  COND2X1 U6360 ( .A(n8113), .B(n6962), .C(n7196), .D(n6947), .Z(n3370) );
  COND2X1 U6361 ( .A(n8112), .B(n6963), .C(n7195), .D(n6943), .Z(n3371) );
  COND2X1 U6362 ( .A(n8111), .B(n6965), .C(n7194), .D(n6946), .Z(n3372) );
  COND2X1 U6363 ( .A(n8110), .B(n6966), .C(n7193), .D(n6947), .Z(n3373) );
  COND2X1 U6364 ( .A(n8109), .B(n6962), .C(n7192), .D(n6942), .Z(n3374) );
  COND2X1 U6365 ( .A(n8108), .B(n6963), .C(n7191), .D(n6943), .Z(n3375) );
  COND2X1 U6366 ( .A(n8107), .B(n6965), .C(n7190), .D(n6944), .Z(n3376) );
  COND2X1 U6367 ( .A(n8106), .B(n6966), .C(n7189), .D(n6944), .Z(n3377) );
  COND2X1 U6368 ( .A(n8105), .B(n6967), .C(n7188), .D(n6942), .Z(n3378) );
  COND2X1 U6369 ( .A(n8104), .B(n6968), .C(n7187), .D(n6943), .Z(n3379) );
  COND2X1 U6370 ( .A(n8103), .B(n6969), .C(n7186), .D(n6945), .Z(n3380) );
  COND2X1 U6371 ( .A(n8102), .B(n6970), .C(n7185), .D(n6946), .Z(n3381) );
  COND2X1 U6372 ( .A(n8101), .B(n6951), .C(n7184), .D(n6947), .Z(n3382) );
  COND2X1 U6373 ( .A(n8100), .B(n6952), .C(n7183), .D(n6945), .Z(n3383) );
  COND2X1 U6374 ( .A(n8099), .B(n6953), .C(n7182), .D(n6944), .Z(n3384) );
  COND2X1 U6375 ( .A(n8098), .B(n6954), .C(n7181), .D(n6945), .Z(n3385) );
  COND2X1 U6376 ( .A(n8097), .B(n6955), .C(n7180), .D(n6942), .Z(n3386) );
  COND2X1 U6377 ( .A(n8096), .B(n6956), .C(n7179), .D(n6943), .Z(n3387) );
  COND2X1 U6378 ( .A(n8095), .B(n6958), .C(n7178), .D(n6944), .Z(n3388) );
  COND2X1 U6379 ( .A(n8094), .B(n6959), .C(n7177), .D(n6946), .Z(n3389) );
  COND2X1 U6380 ( .A(n8093), .B(n6960), .C(n7176), .D(n6946), .Z(n3390) );
  COND2X1 U6381 ( .A(n8092), .B(n6961), .C(n7175), .D(n6947), .Z(n3391) );
  COND2X1 U6382 ( .A(n8091), .B(n6921), .C(n7206), .D(n6912), .Z(n3392) );
  COND2X1 U6383 ( .A(n8090), .B(n6922), .C(n7205), .D(n6913), .Z(n3393) );
  COND2X1 U6384 ( .A(n8089), .B(n6923), .C(n7204), .D(n6912), .Z(n3394) );
  COND2X1 U6385 ( .A(n8088), .B(n6924), .C(n7203), .D(n6913), .Z(n3395) );
  COND2X1 U6386 ( .A(n8087), .B(n6925), .C(n7202), .D(n6914), .Z(n3396) );
  COND2X1 U6387 ( .A(n8086), .B(n6926), .C(n7201), .D(n6912), .Z(n3397) );
  COND2X1 U6388 ( .A(n8085), .B(n6928), .C(n7200), .D(n6914), .Z(n3398) );
  COND2X1 U6389 ( .A(n8084), .B(n6929), .C(n7199), .D(n6915), .Z(n3399) );
  COND2X1 U6390 ( .A(n8083), .B(n6930), .C(n7198), .D(n6915), .Z(n3400) );
  COND2X1 U6391 ( .A(n8082), .B(n6931), .C(n7197), .D(n6916), .Z(n3401) );
  COND2X1 U6392 ( .A(n8081), .B(n6932), .C(n7196), .D(n6917), .Z(n3402) );
  COND2X1 U6393 ( .A(n8080), .B(n6933), .C(n7195), .D(n6913), .Z(n3403) );
  COND2X1 U6394 ( .A(n8079), .B(n6935), .C(n7194), .D(n6916), .Z(n3404) );
  COND2X1 U6395 ( .A(n8078), .B(n6936), .C(n7193), .D(n6917), .Z(n3405) );
  COND2X1 U6396 ( .A(n8077), .B(n6932), .C(n7192), .D(n6912), .Z(n3406) );
  COND2X1 U6397 ( .A(n8076), .B(n6933), .C(n7191), .D(n6913), .Z(n3407) );
  COND2X1 U6398 ( .A(n8075), .B(n6935), .C(n7190), .D(n6914), .Z(n3408) );
  COND2X1 U6399 ( .A(n8074), .B(n6936), .C(n7189), .D(n6914), .Z(n3409) );
  COND2X1 U6400 ( .A(n8073), .B(n6937), .C(n7188), .D(n6912), .Z(n3410) );
  COND2X1 U6401 ( .A(n8072), .B(n6938), .C(n7187), .D(n6913), .Z(n3411) );
  COND2X1 U6402 ( .A(n8071), .B(n6939), .C(n7186), .D(n6915), .Z(n3412) );
  COND2X1 U6403 ( .A(n8070), .B(n6940), .C(n7185), .D(n6916), .Z(n3413) );
  COND2X1 U6404 ( .A(n8069), .B(n6921), .C(n7184), .D(n6917), .Z(n3414) );
  COND2X1 U6405 ( .A(n8068), .B(n6922), .C(n7183), .D(n6915), .Z(n3415) );
  COND2X1 U6406 ( .A(n8067), .B(n6923), .C(n7182), .D(n6914), .Z(n3416) );
  COND2X1 U6407 ( .A(n8066), .B(n6924), .C(n7181), .D(n6915), .Z(n3417) );
  COND2X1 U6408 ( .A(n8065), .B(n6925), .C(n7180), .D(n6912), .Z(n3418) );
  COND2X1 U6409 ( .A(n8064), .B(n6926), .C(n7179), .D(n6913), .Z(n3419) );
  COND2X1 U6410 ( .A(n8063), .B(n6928), .C(n7178), .D(n6914), .Z(n3420) );
  COND2X1 U6411 ( .A(n8062), .B(n6929), .C(n7177), .D(n6916), .Z(n3421) );
  COND2X1 U6412 ( .A(n8061), .B(n6930), .C(n7176), .D(n6916), .Z(n3422) );
  COND2X1 U6413 ( .A(n8060), .B(n6931), .C(n7175), .D(n6917), .Z(n3423) );
  COND2X1 U6414 ( .A(n8059), .B(n6891), .C(n7206), .D(n6882), .Z(n3424) );
  COND2X1 U6415 ( .A(n8058), .B(n6892), .C(n7205), .D(n6883), .Z(n3425) );
  COND2X1 U6416 ( .A(n8057), .B(n6893), .C(n7204), .D(n6882), .Z(n3426) );
  COND2X1 U6417 ( .A(n8056), .B(n6894), .C(n7203), .D(n6883), .Z(n3427) );
  COND2X1 U6418 ( .A(n8055), .B(n6895), .C(n7202), .D(n6884), .Z(n3428) );
  COND2X1 U6419 ( .A(n8054), .B(n6896), .C(n7201), .D(n6882), .Z(n3429) );
  COND2X1 U6420 ( .A(n8053), .B(n6898), .C(n7200), .D(n6884), .Z(n3430) );
  COND2X1 U6421 ( .A(n8052), .B(n6899), .C(n7199), .D(n6885), .Z(n3431) );
  COND2X1 U6422 ( .A(n8051), .B(n6900), .C(n7198), .D(n6885), .Z(n3432) );
  COND2X1 U6423 ( .A(n8050), .B(n6901), .C(n7197), .D(n6886), .Z(n3433) );
  COND2X1 U6424 ( .A(n8049), .B(n6902), .C(n7196), .D(n6887), .Z(n3434) );
  COND2X1 U6425 ( .A(n8048), .B(n6903), .C(n7195), .D(n6883), .Z(n3435) );
  COND2X1 U6426 ( .A(n8047), .B(n6905), .C(n7194), .D(n6886), .Z(n3436) );
  COND2X1 U6427 ( .A(n8046), .B(n6906), .C(n7193), .D(n6887), .Z(n3437) );
  COND2X1 U6428 ( .A(n8043), .B(n6905), .C(n7190), .D(n6884), .Z(n3440) );
  COND2X1 U6429 ( .A(n8042), .B(n6906), .C(n7189), .D(n6884), .Z(n3441) );
  COND2X1 U6430 ( .A(n8041), .B(n6907), .C(n7188), .D(n6882), .Z(n3442) );
  COND2X1 U6431 ( .A(n8040), .B(n6908), .C(n7187), .D(n6883), .Z(n3443) );
  COND2X1 U6432 ( .A(n8039), .B(n6909), .C(n7186), .D(n6885), .Z(n3444) );
  COND2X1 U6433 ( .A(n8038), .B(n6910), .C(n7185), .D(n6886), .Z(n3445) );
  COND2X1 U6434 ( .A(n8037), .B(n6891), .C(n7184), .D(n6887), .Z(n3446) );
  COND2X1 U6435 ( .A(n8036), .B(n6892), .C(n7183), .D(n6885), .Z(n3447) );
  COND2X1 U6436 ( .A(n8035), .B(n6893), .C(n7182), .D(n6884), .Z(n3448) );
  COND2X1 U6437 ( .A(n8034), .B(n6894), .C(n7181), .D(n6885), .Z(n3449) );
  COND2X1 U6438 ( .A(n8033), .B(n6895), .C(n7180), .D(n6882), .Z(n3450) );
  COND2X1 U6439 ( .A(n8032), .B(n6896), .C(n7179), .D(n6883), .Z(n3451) );
  COND2X1 U6440 ( .A(n8031), .B(n6898), .C(n7178), .D(n6884), .Z(n3452) );
  COND2X1 U6441 ( .A(n8030), .B(n6899), .C(n7177), .D(n6886), .Z(n3453) );
  COND2X1 U6442 ( .A(n8029), .B(n6900), .C(n7176), .D(n6886), .Z(n3454) );
  COND2X1 U6443 ( .A(n8028), .B(n6901), .C(n7175), .D(n6887), .Z(n3455) );
  COND2X1 U6444 ( .A(n8013), .B(n6872), .C(n7192), .D(n6852), .Z(n3470) );
  COND2X1 U6445 ( .A(n8012), .B(n6873), .C(n7191), .D(n6853), .Z(n3471) );
  COND2X1 U6446 ( .A(n8011), .B(n6875), .C(n7190), .D(n6854), .Z(n3472) );
  COND2X1 U6447 ( .A(n8010), .B(n6876), .C(n7189), .D(n6854), .Z(n3473) );
  COND2X1 U6448 ( .A(n8009), .B(n6877), .C(n7188), .D(n6852), .Z(n3474) );
  COND2X1 U6449 ( .A(n8008), .B(n6878), .C(n7187), .D(n6853), .Z(n3475) );
  COND2X1 U6450 ( .A(n8007), .B(n6879), .C(n7186), .D(n6855), .Z(n3476) );
  COND2X1 U6451 ( .A(n8006), .B(n6880), .C(n7185), .D(n6856), .Z(n3477) );
  COND2X1 U6452 ( .A(n8005), .B(n6861), .C(n7184), .D(n6857), .Z(n3478) );
  COND2X1 U6453 ( .A(n8004), .B(n6862), .C(n7183), .D(n6855), .Z(n3479) );
  COND2X1 U6454 ( .A(n8003), .B(n6863), .C(n7182), .D(n6854), .Z(n3480) );
  COND2X1 U6455 ( .A(n8002), .B(n6864), .C(n7181), .D(n6855), .Z(n3481) );
  COND2X1 U6456 ( .A(n8001), .B(n6865), .C(n7180), .D(n6852), .Z(n3482) );
  COND2X1 U6457 ( .A(n8000), .B(n6866), .C(n7179), .D(n6853), .Z(n3483) );
  COND2X1 U6458 ( .A(n7999), .B(n6868), .C(n7178), .D(n6854), .Z(n3484) );
  COND2X1 U6459 ( .A(n7998), .B(n6869), .C(n7177), .D(n6856), .Z(n3485) );
  COND2X1 U6460 ( .A(n7997), .B(n6870), .C(n7176), .D(n6856), .Z(n3486) );
  COND2X1 U6461 ( .A(n7996), .B(n6871), .C(n7175), .D(n6857), .Z(n3487) );
  COND2X1 U6462 ( .A(n7995), .B(n6831), .C(n7206), .D(n6822), .Z(n3488) );
  COND2X1 U6463 ( .A(n7994), .B(n6832), .C(n7205), .D(n6823), .Z(n3489) );
  COND2X1 U6464 ( .A(n7993), .B(n6833), .C(n7204), .D(n6822), .Z(n3490) );
  COND2X1 U6465 ( .A(n7992), .B(n6834), .C(n7203), .D(n6823), .Z(n3491) );
  COND2X1 U6466 ( .A(n7991), .B(n6835), .C(n7202), .D(n6824), .Z(n3492) );
  COND2X1 U6467 ( .A(n7990), .B(n6836), .C(n7201), .D(n6822), .Z(n3493) );
  COND2X1 U6468 ( .A(n7989), .B(n6838), .C(n7200), .D(n6824), .Z(n3494) );
  COND2X1 U6469 ( .A(n7988), .B(n6839), .C(n7199), .D(n6825), .Z(n3495) );
  COND2X1 U6470 ( .A(n7987), .B(n6840), .C(n7198), .D(n6825), .Z(n3496) );
  COND2X1 U6471 ( .A(n7986), .B(n6841), .C(n7197), .D(n6826), .Z(n3497) );
  COND2X1 U6472 ( .A(n7985), .B(n6842), .C(n7196), .D(n6827), .Z(n3498) );
  COND2X1 U6473 ( .A(n7984), .B(n6843), .C(n7195), .D(n6823), .Z(n3499) );
  COND2X1 U6474 ( .A(n7983), .B(n6845), .C(n7194), .D(n6826), .Z(n3500) );
  COND2X1 U6475 ( .A(n7982), .B(n6846), .C(n7193), .D(n6827), .Z(n3501) );
  COND2X1 U6476 ( .A(n7981), .B(n6842), .C(n7192), .D(n6822), .Z(n3502) );
  COND2X1 U6477 ( .A(n7980), .B(n6843), .C(n7191), .D(n6823), .Z(n3503) );
  COND2X1 U6478 ( .A(n7979), .B(n6845), .C(n7190), .D(n6824), .Z(n3504) );
  COND2X1 U6479 ( .A(n7978), .B(n6846), .C(n7189), .D(n6824), .Z(n3505) );
  COND2X1 U6480 ( .A(n7977), .B(n6847), .C(n7188), .D(n6822), .Z(n3506) );
  COND2X1 U6481 ( .A(n7976), .B(n6848), .C(n7187), .D(n6823), .Z(n3507) );
  COND2X1 U6482 ( .A(n7975), .B(n6849), .C(n7186), .D(n6825), .Z(n3508) );
  COND2X1 U6483 ( .A(n7974), .B(n6850), .C(n7185), .D(n6826), .Z(n3509) );
  COND2X1 U6484 ( .A(n7973), .B(n6831), .C(n7184), .D(n6827), .Z(n3510) );
  COND2X1 U6485 ( .A(n7972), .B(n6832), .C(n7183), .D(n6825), .Z(n3511) );
  COND2X1 U6486 ( .A(n7971), .B(n6833), .C(n7182), .D(n6824), .Z(n3512) );
  COND2X1 U6487 ( .A(n7970), .B(n6834), .C(n7181), .D(n6825), .Z(n3513) );
  COND2X1 U6488 ( .A(n7969), .B(n6835), .C(n7180), .D(n6822), .Z(n3514) );
  COND2X1 U6489 ( .A(n7968), .B(n6836), .C(n7179), .D(n6823), .Z(n3515) );
  COND2X1 U6490 ( .A(n7967), .B(n6838), .C(n7178), .D(n6824), .Z(n3516) );
  COND2X1 U6491 ( .A(n7966), .B(n6839), .C(n7177), .D(n6826), .Z(n3517) );
  COND2X1 U6492 ( .A(n7965), .B(n6840), .C(n7176), .D(n6826), .Z(n3518) );
  COND2X1 U6493 ( .A(n7964), .B(n6841), .C(n7175), .D(n6827), .Z(n3519) );
  COND2X1 U6494 ( .A(n7963), .B(n6801), .C(n7206), .D(n6792), .Z(n3520) );
  COND2X1 U6495 ( .A(n7962), .B(n6802), .C(n7205), .D(n6793), .Z(n3521) );
  COND2X1 U6496 ( .A(n7961), .B(n6803), .C(n7204), .D(n6792), .Z(n3522) );
  COND2X1 U6497 ( .A(n7960), .B(n6804), .C(n7203), .D(n6793), .Z(n3523) );
  COND2X1 U6498 ( .A(n7959), .B(n6805), .C(n7202), .D(n6794), .Z(n3524) );
  COND2X1 U6499 ( .A(n7958), .B(n6806), .C(n7201), .D(n6792), .Z(n3525) );
  COND2X1 U6500 ( .A(n7957), .B(n6808), .C(n7200), .D(n6794), .Z(n3526) );
  COND2X1 U6501 ( .A(n7956), .B(n6809), .C(n7199), .D(n6795), .Z(n3527) );
  COND2X1 U6502 ( .A(n7955), .B(n6810), .C(n7198), .D(n6795), .Z(n3528) );
  COND2X1 U6503 ( .A(n7954), .B(n6811), .C(n7197), .D(n6796), .Z(n3529) );
  COND2X1 U6504 ( .A(n7953), .B(n6812), .C(n7196), .D(n6797), .Z(n3530) );
  COND2X1 U6505 ( .A(n7952), .B(n6813), .C(n7195), .D(n6793), .Z(n3531) );
  COND2X1 U6506 ( .A(n7951), .B(n6815), .C(n7194), .D(n6796), .Z(n3532) );
  COND2X1 U6507 ( .A(n7950), .B(n6816), .C(n7193), .D(n6797), .Z(n3533) );
  COND2X1 U6508 ( .A(n7949), .B(n6812), .C(n7192), .D(n6792), .Z(n3534) );
  COND2X1 U6509 ( .A(n7948), .B(n6813), .C(n7191), .D(n6793), .Z(n3535) );
  COND2X1 U6510 ( .A(n7947), .B(n6815), .C(n7190), .D(n6794), .Z(n3536) );
  COND2X1 U6511 ( .A(n7946), .B(n6816), .C(n7189), .D(n6794), .Z(n3537) );
  COND2X1 U6512 ( .A(n7945), .B(n6817), .C(n7188), .D(n6792), .Z(n3538) );
  COND2X1 U6513 ( .A(n7944), .B(n6818), .C(n7187), .D(n6793), .Z(n3539) );
  COND2X1 U6514 ( .A(n7943), .B(n6819), .C(n7186), .D(n6795), .Z(n3540) );
  COND2X1 U6515 ( .A(n7942), .B(n6820), .C(n7185), .D(n6796), .Z(n3541) );
  COND2X1 U6516 ( .A(n7941), .B(n6801), .C(n7184), .D(n6797), .Z(n3542) );
  COND2X1 U6517 ( .A(n7940), .B(n6802), .C(n7183), .D(n6795), .Z(n3543) );
  COND2X1 U6518 ( .A(n7939), .B(n6803), .C(n7182), .D(n6794), .Z(n3544) );
  COND2X1 U6519 ( .A(n7938), .B(n6804), .C(n7181), .D(n6795), .Z(n3545) );
  COND2X1 U6520 ( .A(n7937), .B(n6805), .C(n7180), .D(n6792), .Z(n3546) );
  COND2X1 U6521 ( .A(n7936), .B(n6806), .C(n7179), .D(n6793), .Z(n3547) );
  COND2X1 U6522 ( .A(n7935), .B(n6808), .C(n7178), .D(n6794), .Z(n3548) );
  COND2X1 U6523 ( .A(n7934), .B(n6809), .C(n7177), .D(n6796), .Z(n3549) );
  COND2X1 U6524 ( .A(n7933), .B(n6810), .C(n7176), .D(n6796), .Z(n3550) );
  COND2X1 U6525 ( .A(n7932), .B(n6811), .C(n7175), .D(n6797), .Z(n3551) );
  COND2X1 U6526 ( .A(n7931), .B(n6771), .C(n7206), .D(n6762), .Z(n3552) );
  COND2X1 U6527 ( .A(n7930), .B(n6772), .C(n7205), .D(n6763), .Z(n3553) );
  COND2X1 U6528 ( .A(n7929), .B(n6773), .C(n7204), .D(n6762), .Z(n3554) );
  COND2X1 U6529 ( .A(n7928), .B(n6774), .C(n7203), .D(n6763), .Z(n3555) );
  COND2X1 U6530 ( .A(n7927), .B(n6775), .C(n7202), .D(n6764), .Z(n3556) );
  COND2X1 U6531 ( .A(n7926), .B(n6776), .C(n7201), .D(n6762), .Z(n3557) );
  COND2X1 U6532 ( .A(n7925), .B(n6778), .C(n7200), .D(n6764), .Z(n3558) );
  COND2X1 U6533 ( .A(n7924), .B(n6779), .C(n7199), .D(n6765), .Z(n3559) );
  COND2X1 U6534 ( .A(n7923), .B(n6780), .C(n7198), .D(n6765), .Z(n3560) );
  COND2X1 U6535 ( .A(n7922), .B(n6781), .C(n7197), .D(n6766), .Z(n3561) );
  COND2X1 U6536 ( .A(n7921), .B(n6782), .C(n7196), .D(n6767), .Z(n3562) );
  COND2X1 U6537 ( .A(n7920), .B(n6783), .C(n7195), .D(n6763), .Z(n3563) );
  COND2X1 U6538 ( .A(n7919), .B(n6785), .C(n7194), .D(n6766), .Z(n3564) );
  COND2X1 U6539 ( .A(n7918), .B(n6786), .C(n7193), .D(n6767), .Z(n3565) );
  COND2X1 U6540 ( .A(n7917), .B(n6782), .C(n7192), .D(n6762), .Z(n3566) );
  COND2X1 U6541 ( .A(n7916), .B(n6783), .C(n7191), .D(n6763), .Z(n3567) );
  COND2X1 U6542 ( .A(n7915), .B(n6785), .C(n7190), .D(n6764), .Z(n3568) );
  COND2X1 U6543 ( .A(n7914), .B(n6786), .C(n7189), .D(n6764), .Z(n3569) );
  COND2X1 U6544 ( .A(n7913), .B(n6787), .C(n7188), .D(n6762), .Z(n3570) );
  COND2X1 U6545 ( .A(n7912), .B(n6788), .C(n7187), .D(n6763), .Z(n3571) );
  COND2X1 U6546 ( .A(n7911), .B(n6789), .C(n7186), .D(n6765), .Z(n3572) );
  COND2X1 U6547 ( .A(n7910), .B(n6790), .C(n7185), .D(n6766), .Z(n3573) );
  COND2X1 U6548 ( .A(n7909), .B(n6771), .C(n7184), .D(n6767), .Z(n3574) );
  COND2X1 U6549 ( .A(n7908), .B(n6772), .C(n7183), .D(n6765), .Z(n3575) );
  COND2X1 U6550 ( .A(n7907), .B(n6773), .C(n7182), .D(n6764), .Z(n3576) );
  COND2X1 U6551 ( .A(n7906), .B(n6774), .C(n7181), .D(n6765), .Z(n3577) );
  COND2X1 U6552 ( .A(n7905), .B(n6775), .C(n7180), .D(n6762), .Z(n3578) );
  COND2X1 U6553 ( .A(n7904), .B(n6776), .C(n7179), .D(n6763), .Z(n3579) );
  COND2X1 U6554 ( .A(n7903), .B(n6778), .C(n7178), .D(n6764), .Z(n3580) );
  COND2X1 U6555 ( .A(n7902), .B(n6779), .C(n7177), .D(n6766), .Z(n3581) );
  COND2X1 U6556 ( .A(n7901), .B(n6780), .C(n7176), .D(n6766), .Z(n3582) );
  COND2X1 U6557 ( .A(n7900), .B(n6781), .C(n7175), .D(n6767), .Z(n3583) );
  COND2X1 U6558 ( .A(n7885), .B(n6752), .C(n7192), .D(n6732), .Z(n3598) );
  COND2X1 U6559 ( .A(n7884), .B(n6753), .C(n7191), .D(n6733), .Z(n3599) );
  COND2X1 U6560 ( .A(n7883), .B(n6755), .C(n7190), .D(n6734), .Z(n3600) );
  COND2X1 U6561 ( .A(n7882), .B(n6756), .C(n7189), .D(n6734), .Z(n3601) );
  COND2X1 U6562 ( .A(n7881), .B(n6757), .C(n7188), .D(n6732), .Z(n3602) );
  COND2X1 U6563 ( .A(n7880), .B(n6758), .C(n7187), .D(n6733), .Z(n3603) );
  COND2X1 U6564 ( .A(n7879), .B(n6759), .C(n7186), .D(n6735), .Z(n3604) );
  COND2X1 U6565 ( .A(n7878), .B(n6760), .C(n7185), .D(n6736), .Z(n3605) );
  COND2X1 U6566 ( .A(n7877), .B(n6741), .C(n7184), .D(n6737), .Z(n3606) );
  COND2X1 U6567 ( .A(n7876), .B(n6742), .C(n7183), .D(n6735), .Z(n3607) );
  COND2X1 U6568 ( .A(n7875), .B(n6743), .C(n7182), .D(n6734), .Z(n3608) );
  COND2X1 U6569 ( .A(n7874), .B(n6744), .C(n7181), .D(n6735), .Z(n3609) );
  COND2X1 U6570 ( .A(n7873), .B(n6745), .C(n7180), .D(n6732), .Z(n3610) );
  COND2X1 U6571 ( .A(n7872), .B(n6746), .C(n7179), .D(n6733), .Z(n3611) );
  COND2X1 U6572 ( .A(n7871), .B(n6748), .C(n7178), .D(n6734), .Z(n3612) );
  COND2X1 U6573 ( .A(n7870), .B(n6749), .C(n7177), .D(n6736), .Z(n3613) );
  COND2X1 U6574 ( .A(n7869), .B(n6750), .C(n7176), .D(n6736), .Z(n3614) );
  COND2X1 U6575 ( .A(n7868), .B(n6751), .C(n7175), .D(n6737), .Z(n3615) );
  COND2X1 U6576 ( .A(n7867), .B(n6711), .C(n7206), .D(n6704), .Z(n3616) );
  COND2X1 U6577 ( .A(n7866), .B(n6712), .C(n7205), .D(n6705), .Z(n3617) );
  COND2X1 U6578 ( .A(n7865), .B(n6713), .C(n7204), .D(n6706), .Z(n3618) );
  COND2X1 U6579 ( .A(n7864), .B(n6714), .C(n7203), .D(n6707), .Z(n3619) );
  COND2X1 U6580 ( .A(n7863), .B(n6715), .C(n7202), .D(n6707), .Z(n3620) );
  COND2X1 U6581 ( .A(n7862), .B(n6716), .C(n7201), .D(n6704), .Z(n3621) );
  COND2X1 U6582 ( .A(n7861), .B(n6718), .C(n7200), .D(n6705), .Z(n3622) );
  COND2X1 U6583 ( .A(n7860), .B(n6719), .C(n7199), .D(n6704), .Z(n3623) );
  COND2X1 U6584 ( .A(n7859), .B(n6720), .C(n7198), .D(n6706), .Z(n3624) );
  COND2X1 U6585 ( .A(n7858), .B(n6721), .C(n7197), .D(n6707), .Z(n3625) );
  COND2X1 U6586 ( .A(n7857), .B(n6722), .C(n7196), .D(n6704), .Z(n3626) );
  COND2X1 U6587 ( .A(n7856), .B(n6723), .C(n7195), .D(n6705), .Z(n3627) );
  COND2X1 U6588 ( .A(n7855), .B(n6725), .C(n7194), .D(n6705), .Z(n3628) );
  COND2X1 U6589 ( .A(n7854), .B(n6726), .C(n7193), .D(n6706), .Z(n3629) );
  COND2X1 U6590 ( .A(n7853), .B(n6722), .C(n7192), .D(n6707), .Z(n3630) );
  COND2X1 U6591 ( .A(n7852), .B(n6723), .C(n7191), .D(n6706), .Z(n3631) );
  COND2X1 U6592 ( .A(n7851), .B(n6725), .C(n7190), .D(n6704), .Z(n3632) );
  COND2X1 U6593 ( .A(n7850), .B(n6726), .C(n7189), .D(n6705), .Z(n3633) );
  COND2X1 U6594 ( .A(n7849), .B(n6727), .C(n7188), .D(n6706), .Z(n3634) );
  COND2X1 U6595 ( .A(n7848), .B(n6728), .C(n7187), .D(n6707), .Z(n3635) );
  COND2X1 U6596 ( .A(n7847), .B(n6729), .C(n7186), .D(n6707), .Z(n3636) );
  COND2X1 U6597 ( .A(n7846), .B(n6730), .C(n7185), .D(n6704), .Z(n3637) );
  COND2X1 U6598 ( .A(n7845), .B(n6711), .C(n7184), .D(n6705), .Z(n3638) );
  COND2X1 U6599 ( .A(n7844), .B(n6712), .C(n7183), .D(n6704), .Z(n3639) );
  COND2X1 U6600 ( .A(n7843), .B(n6713), .C(n7182), .D(n6706), .Z(n3640) );
  COND2X1 U6601 ( .A(n7842), .B(n6714), .C(n7181), .D(n6707), .Z(n3641) );
  COND2X1 U6602 ( .A(n7841), .B(n6715), .C(n7180), .D(n6704), .Z(n3642) );
  COND2X1 U6603 ( .A(n7840), .B(n6716), .C(n7179), .D(n6705), .Z(n3643) );
  COND2X1 U6604 ( .A(n7839), .B(n6718), .C(n7178), .D(n6705), .Z(n3644) );
  COND2X1 U6605 ( .A(n7838), .B(n6719), .C(n7177), .D(n6706), .Z(n3645) );
  COND2X1 U6606 ( .A(n7837), .B(n6720), .C(n7176), .D(n6707), .Z(n3646) );
  COND2X1 U6607 ( .A(n7836), .B(n6721), .C(n7175), .D(n6706), .Z(n3647) );
  COND2X1 U6608 ( .A(n7835), .B(n6684), .C(n7206), .D(n6677), .Z(n3648) );
  COND2X1 U6609 ( .A(n7834), .B(n6685), .C(n7205), .D(n6678), .Z(n3649) );
  COND2X1 U6610 ( .A(n7833), .B(n6686), .C(n7204), .D(n6679), .Z(n3650) );
  COND2X1 U6611 ( .A(n7832), .B(n6687), .C(n7203), .D(n6680), .Z(n3651) );
  COND2X1 U6612 ( .A(n7831), .B(n6688), .C(n7202), .D(n6680), .Z(n3652) );
  COND2X1 U6613 ( .A(n7830), .B(n6689), .C(n7201), .D(n6677), .Z(n3653) );
  COND2X1 U6614 ( .A(n7829), .B(n6691), .C(n7200), .D(n6678), .Z(n3654) );
  COND2X1 U6615 ( .A(n7828), .B(n6692), .C(n7199), .D(n6677), .Z(n3655) );
  COND2X1 U6616 ( .A(n7827), .B(n6693), .C(n7198), .D(n6679), .Z(n3656) );
  COND2X1 U6617 ( .A(n7826), .B(n6694), .C(n7197), .D(n6680), .Z(n3657) );
  COND2X1 U6618 ( .A(n7825), .B(n6695), .C(n7196), .D(n6677), .Z(n3658) );
  COND2X1 U6619 ( .A(n7824), .B(n6696), .C(n7195), .D(n6678), .Z(n3659) );
  COND2X1 U6620 ( .A(n7823), .B(n6698), .C(n7194), .D(n6678), .Z(n3660) );
  COND2X1 U6621 ( .A(n7822), .B(n6699), .C(n7193), .D(n6679), .Z(n3661) );
  COND2X1 U6622 ( .A(n7821), .B(n6695), .C(n7192), .D(n6680), .Z(n3662) );
  COND2X1 U6623 ( .A(n7820), .B(n6696), .C(n7191), .D(n6679), .Z(n3663) );
  COND2X1 U6624 ( .A(n7819), .B(n6698), .C(n7190), .D(n6677), .Z(n3664) );
  COND2X1 U6625 ( .A(n7818), .B(n6699), .C(n7189), .D(n6678), .Z(n3665) );
  COND2X1 U6626 ( .A(n7817), .B(n6700), .C(n7188), .D(n6679), .Z(n3666) );
  COND2X1 U6627 ( .A(n7816), .B(n6701), .C(n7187), .D(n6680), .Z(n3667) );
  COND2X1 U6628 ( .A(n7815), .B(n6702), .C(n7186), .D(n6680), .Z(n3668) );
  COND2X1 U6629 ( .A(n7814), .B(n6703), .C(n7185), .D(n6677), .Z(n3669) );
  COND2X1 U6630 ( .A(n7813), .B(n6684), .C(n7184), .D(n6678), .Z(n3670) );
  COND2X1 U6631 ( .A(n7812), .B(n6685), .C(n7183), .D(n6677), .Z(n3671) );
  COND2X1 U6632 ( .A(n7811), .B(n6686), .C(n7182), .D(n6679), .Z(n3672) );
  COND2X1 U6633 ( .A(n7810), .B(n6687), .C(n7181), .D(n6680), .Z(n3673) );
  COND2X1 U6634 ( .A(n7809), .B(n6688), .C(n7180), .D(n6677), .Z(n3674) );
  COND2X1 U6635 ( .A(n7808), .B(n6689), .C(n7179), .D(n6678), .Z(n3675) );
  COND2X1 U6636 ( .A(n7807), .B(n6691), .C(n7178), .D(n6678), .Z(n3676) );
  COND2X1 U6637 ( .A(n7806), .B(n6692), .C(n7177), .D(n6679), .Z(n3677) );
  COND2X1 U6638 ( .A(n7805), .B(n6693), .C(n7176), .D(n6680), .Z(n3678) );
  COND2X1 U6639 ( .A(n7804), .B(n6694), .C(n7175), .D(n6679), .Z(n3679) );
  COND2X1 U6640 ( .A(n7803), .B(n6657), .C(n7206), .D(n6650), .Z(n3680) );
  COND2X1 U6641 ( .A(n7802), .B(n6658), .C(n7205), .D(n6651), .Z(n3681) );
  COND2X1 U6642 ( .A(n7801), .B(n6659), .C(n7204), .D(n6652), .Z(n3682) );
  COND2X1 U6643 ( .A(n7800), .B(n6660), .C(n7203), .D(n6653), .Z(n3683) );
  COND2X1 U6644 ( .A(n7799), .B(n6661), .C(n7202), .D(n6653), .Z(n3684) );
  COND2X1 U6645 ( .A(n7798), .B(n6662), .C(n7201), .D(n6650), .Z(n3685) );
  COND2X1 U6646 ( .A(n7797), .B(n6664), .C(n7200), .D(n6651), .Z(n3686) );
  COND2X1 U6647 ( .A(n7796), .B(n6665), .C(n7199), .D(n6650), .Z(n3687) );
  COND2X1 U6648 ( .A(n7795), .B(n6666), .C(n7198), .D(n6652), .Z(n3688) );
  COND2X1 U6649 ( .A(n7794), .B(n6667), .C(n7197), .D(n6653), .Z(n3689) );
  COND2X1 U6650 ( .A(n7793), .B(n6668), .C(n7196), .D(n6650), .Z(n3690) );
  COND2X1 U6651 ( .A(n7792), .B(n6669), .C(n7195), .D(n6651), .Z(n3691) );
  COND2X1 U6652 ( .A(n7791), .B(n6671), .C(n7194), .D(n6651), .Z(n3692) );
  COND2X1 U6653 ( .A(n7790), .B(n6672), .C(n7193), .D(n6652), .Z(n3693) );
  COND2X1 U6654 ( .A(n7789), .B(n6668), .C(n7192), .D(n6653), .Z(n3694) );
  COND2X1 U6655 ( .A(n7788), .B(n6669), .C(n7191), .D(n6652), .Z(n3695) );
  COND2X1 U6656 ( .A(n7787), .B(n6671), .C(n7190), .D(n6650), .Z(n3696) );
  COND2X1 U6657 ( .A(n7786), .B(n6672), .C(n7189), .D(n6651), .Z(n3697) );
  COND2X1 U6658 ( .A(n7785), .B(n6673), .C(n7188), .D(n6652), .Z(n3698) );
  COND2X1 U6659 ( .A(n7784), .B(n6674), .C(n7187), .D(n6653), .Z(n3699) );
  COND2X1 U6660 ( .A(n7783), .B(n6675), .C(n7186), .D(n6653), .Z(n3700) );
  COND2X1 U6661 ( .A(n7782), .B(n6676), .C(n7185), .D(n6650), .Z(n3701) );
  COND2X1 U6662 ( .A(n7781), .B(n6657), .C(n7184), .D(n6651), .Z(n3702) );
  COND2X1 U6663 ( .A(n7780), .B(n6658), .C(n7183), .D(n6650), .Z(n3703) );
  COND2X1 U6664 ( .A(n7779), .B(n6659), .C(n7182), .D(n6652), .Z(n3704) );
  COND2X1 U6665 ( .A(n7778), .B(n6660), .C(n7181), .D(n6653), .Z(n3705) );
  COND2X1 U6666 ( .A(n7777), .B(n6661), .C(n7180), .D(n6650), .Z(n3706) );
  COND2X1 U6667 ( .A(n7776), .B(n6662), .C(n7179), .D(n6651), .Z(n3707) );
  COND2X1 U6668 ( .A(n7775), .B(n6664), .C(n7178), .D(n6651), .Z(n3708) );
  COND2X1 U6669 ( .A(n7774), .B(n6665), .C(n7177), .D(n6652), .Z(n3709) );
  COND2X1 U6670 ( .A(n7773), .B(n6666), .C(n7176), .D(n6653), .Z(n3710) );
  COND2X1 U6671 ( .A(n7772), .B(n6667), .C(n7175), .D(n6652), .Z(n3711) );
  COND2X1 U6672 ( .A(n7759), .B(n6644), .C(n7194), .D(n6625), .Z(n3724) );
  COND2X1 U6673 ( .A(n7755), .B(n6644), .C(n7190), .D(n6623), .Z(n3728) );
  COND2X1 U6674 ( .A(n7754), .B(n6645), .C(n7189), .D(n6623), .Z(n3729) );
  COND2X1 U6675 ( .A(n7753), .B(n6646), .C(n7188), .D(n6621), .Z(n3730) );
  COND2X1 U6676 ( .A(n7752), .B(n6647), .C(n7187), .D(n6622), .Z(n3731) );
  COND2X1 U6677 ( .A(n7751), .B(n6648), .C(n7186), .D(n6624), .Z(n3732) );
  COND2X1 U6678 ( .A(n7750), .B(n6649), .C(n7185), .D(n6625), .Z(n3733) );
  COND2X1 U6679 ( .A(n7749), .B(n6630), .C(n7184), .D(n6626), .Z(n3734) );
  COND2X1 U6680 ( .A(n7748), .B(n6631), .C(n7183), .D(n6624), .Z(n3735) );
  COND2X1 U6681 ( .A(n7747), .B(n6632), .C(n7182), .D(n6623), .Z(n3736) );
  COND2X1 U6682 ( .A(n7746), .B(n6633), .C(n7181), .D(n6624), .Z(n3737) );
  COND2X1 U6683 ( .A(n7745), .B(n6634), .C(n7180), .D(n6621), .Z(n3738) );
  COND2X1 U6684 ( .A(n7744), .B(n6635), .C(n7179), .D(n6622), .Z(n3739) );
  COND2X1 U6685 ( .A(n7743), .B(n6637), .C(n7178), .D(n6623), .Z(n3740) );
  COND2X1 U6686 ( .A(n7742), .B(n6638), .C(n7177), .D(n6625), .Z(n3741) );
  COND2X1 U6687 ( .A(n7741), .B(n6639), .C(n7176), .D(n6625), .Z(n3742) );
  COND2X1 U6688 ( .A(n7740), .B(n6640), .C(n7175), .D(n6626), .Z(n3743) );
  COND2X1 U6689 ( .A(n7739), .B(n6600), .C(n7206), .D(n6591), .Z(n3744) );
  COND2X1 U6690 ( .A(n7738), .B(n6601), .C(n7205), .D(n6592), .Z(n3745) );
  COND2X1 U6691 ( .A(n7737), .B(n6602), .C(n7204), .D(n6591), .Z(n3746) );
  COND2X1 U6692 ( .A(n7736), .B(n6603), .C(n7203), .D(n6592), .Z(n3747) );
  COND2X1 U6693 ( .A(n7735), .B(n6604), .C(n7202), .D(n6593), .Z(n3748) );
  COND2X1 U6694 ( .A(n7734), .B(n6605), .C(n7201), .D(n6591), .Z(n3749) );
  COND2X1 U6695 ( .A(n7733), .B(n6607), .C(n7200), .D(n6593), .Z(n3750) );
  COND2X1 U6696 ( .A(n7732), .B(n6608), .C(n7199), .D(n6594), .Z(n3751) );
  COND2X1 U6697 ( .A(n7731), .B(n6609), .C(n7198), .D(n6594), .Z(n3752) );
  COND2X1 U6698 ( .A(n7730), .B(n6610), .C(n7197), .D(n6595), .Z(n3753) );
  COND2X1 U6699 ( .A(n7729), .B(n6611), .C(n7196), .D(n6596), .Z(n3754) );
  COND2X1 U6700 ( .A(n7728), .B(n6612), .C(n7195), .D(n6592), .Z(n3755) );
  COND2X1 U6701 ( .A(n7727), .B(n6614), .C(n7194), .D(n6595), .Z(n3756) );
  COND2X1 U6702 ( .A(n7726), .B(n6615), .C(n7193), .D(n6596), .Z(n3757) );
  COND2X1 U6703 ( .A(n7725), .B(n6611), .C(n7192), .D(n6591), .Z(n3758) );
  COND2X1 U6704 ( .A(n7724), .B(n6612), .C(n7191), .D(n6592), .Z(n3759) );
  COND2X1 U6705 ( .A(n7723), .B(n6614), .C(n7190), .D(n6593), .Z(n3760) );
  COND2X1 U6706 ( .A(n7722), .B(n6615), .C(n7189), .D(n6593), .Z(n3761) );
  COND2X1 U6707 ( .A(n7721), .B(n6616), .C(n7188), .D(n6591), .Z(n3762) );
  COND2X1 U6708 ( .A(n7720), .B(n6617), .C(n7187), .D(n6592), .Z(n3763) );
  COND2X1 U6709 ( .A(n7719), .B(n6618), .C(n7186), .D(n6594), .Z(n3764) );
  COND2X1 U6710 ( .A(n7718), .B(n6619), .C(n7185), .D(n6595), .Z(n3765) );
  COND2X1 U6711 ( .A(n7717), .B(n6600), .C(n7184), .D(n6596), .Z(n3766) );
  COND2X1 U6712 ( .A(n7716), .B(n6601), .C(n7183), .D(n6594), .Z(n3767) );
  COND2X1 U6713 ( .A(n7715), .B(n6602), .C(n7182), .D(n6593), .Z(n3768) );
  COND2X1 U6714 ( .A(n7714), .B(n6603), .C(n7181), .D(n6594), .Z(n3769) );
  COND2X1 U6715 ( .A(n7713), .B(n6604), .C(n7180), .D(n6591), .Z(n3770) );
  COND2X1 U6716 ( .A(n7712), .B(n6605), .C(n7179), .D(n6592), .Z(n3771) );
  COND2X1 U6717 ( .A(n7711), .B(n6607), .C(n7178), .D(n6593), .Z(n3772) );
  COND2X1 U6718 ( .A(n7710), .B(n6608), .C(n7177), .D(n6595), .Z(n3773) );
  COND2X1 U6719 ( .A(n7709), .B(n6609), .C(n7176), .D(n6595), .Z(n3774) );
  COND2X1 U6720 ( .A(n7708), .B(n6610), .C(n7175), .D(n6596), .Z(n3775) );
  COND2X1 U6721 ( .A(n7707), .B(n6570), .C(n7206), .D(n6561), .Z(n3776) );
  COND2X1 U6722 ( .A(n7706), .B(n6571), .C(n7205), .D(n6562), .Z(n3777) );
  COND2X1 U6723 ( .A(n7705), .B(n6572), .C(n7204), .D(n6561), .Z(n3778) );
  COND2X1 U6724 ( .A(n7704), .B(n6573), .C(n7203), .D(n6562), .Z(n3779) );
  COND2X1 U6725 ( .A(n7703), .B(n6574), .C(n7202), .D(n6563), .Z(n3780) );
  COND2X1 U6726 ( .A(n7702), .B(n6575), .C(n7201), .D(n6561), .Z(n3781) );
  COND2X1 U6727 ( .A(n7701), .B(n6577), .C(n7200), .D(n6563), .Z(n3782) );
  COND2X1 U6728 ( .A(n7700), .B(n6578), .C(n7199), .D(n6564), .Z(n3783) );
  COND2X1 U6729 ( .A(n7699), .B(n6579), .C(n7198), .D(n6564), .Z(n3784) );
  COND2X1 U6730 ( .A(n7698), .B(n6580), .C(n7197), .D(n6565), .Z(n3785) );
  COND2X1 U6731 ( .A(n7697), .B(n6581), .C(n7196), .D(n6566), .Z(n3786) );
  COND2X1 U6732 ( .A(n7696), .B(n6582), .C(n7195), .D(n6562), .Z(n3787) );
  COND2X1 U6733 ( .A(n7695), .B(n6584), .C(n7194), .D(n6565), .Z(n3788) );
  COND2X1 U6734 ( .A(n7694), .B(n6585), .C(n7193), .D(n6566), .Z(n3789) );
  COND2X1 U6735 ( .A(n7693), .B(n6581), .C(n7192), .D(n6561), .Z(n3790) );
  COND2X1 U6736 ( .A(n7692), .B(n6582), .C(n7191), .D(n6562), .Z(n3791) );
  COND2X1 U6737 ( .A(n7691), .B(n6584), .C(n7190), .D(n6563), .Z(n3792) );
  COND2X1 U6738 ( .A(n7690), .B(n6585), .C(n7189), .D(n6563), .Z(n3793) );
  COND2X1 U6739 ( .A(n7689), .B(n6586), .C(n7188), .D(n6561), .Z(n3794) );
  COND2X1 U6740 ( .A(n7688), .B(n6587), .C(n7187), .D(n6562), .Z(n3795) );
  COND2X1 U6741 ( .A(n7687), .B(n6588), .C(n7186), .D(n6564), .Z(n3796) );
  COND2X1 U6742 ( .A(n7686), .B(n6589), .C(n7185), .D(n6565), .Z(n3797) );
  COND2X1 U6743 ( .A(n7685), .B(n6570), .C(n7184), .D(n6566), .Z(n3798) );
  COND2X1 U6744 ( .A(n7684), .B(n6571), .C(n7183), .D(n6564), .Z(n3799) );
  COND2X1 U6745 ( .A(n7683), .B(n6572), .C(n7182), .D(n6563), .Z(n3800) );
  COND2X1 U6746 ( .A(n7682), .B(n6573), .C(n7181), .D(n6564), .Z(n3801) );
  COND2X1 U6747 ( .A(n7681), .B(n6574), .C(n7180), .D(n6561), .Z(n3802) );
  COND2X1 U6748 ( .A(n7680), .B(n6575), .C(n7179), .D(n6562), .Z(n3803) );
  COND2X1 U6749 ( .A(n7679), .B(n6577), .C(n7178), .D(n6563), .Z(n3804) );
  COND2X1 U6750 ( .A(n7678), .B(n6578), .C(n7177), .D(n6565), .Z(n3805) );
  COND2X1 U6751 ( .A(n7677), .B(n6579), .C(n7176), .D(n6565), .Z(n3806) );
  COND2X1 U6752 ( .A(n7676), .B(n6580), .C(n7175), .D(n6566), .Z(n3807) );
  COND2X1 U6753 ( .A(n7675), .B(n6540), .C(n7206), .D(n6531), .Z(n3808) );
  COND2X1 U6754 ( .A(n7674), .B(n6541), .C(n7205), .D(n6532), .Z(n3809) );
  COND2X1 U6755 ( .A(n7673), .B(n6542), .C(n7204), .D(n6531), .Z(n3810) );
  COND2X1 U6756 ( .A(n7672), .B(n6543), .C(n7203), .D(n6532), .Z(n3811) );
  COND2X1 U6757 ( .A(n7671), .B(n6544), .C(n7202), .D(n6533), .Z(n3812) );
  COND2X1 U6758 ( .A(n7670), .B(n6545), .C(n7201), .D(n6531), .Z(n3813) );
  COND2X1 U6759 ( .A(n7669), .B(n6547), .C(n7200), .D(n6533), .Z(n3814) );
  COND2X1 U6760 ( .A(n7668), .B(n6548), .C(n7199), .D(n6534), .Z(n3815) );
  COND2X1 U6761 ( .A(n7667), .B(n6549), .C(n7198), .D(n6534), .Z(n3816) );
  COND2X1 U6762 ( .A(n7666), .B(n6550), .C(n7197), .D(n6535), .Z(n3817) );
  COND2X1 U6763 ( .A(n7665), .B(n6551), .C(n7196), .D(n6536), .Z(n3818) );
  COND2X1 U6764 ( .A(n7664), .B(n6552), .C(n7195), .D(n6532), .Z(n3819) );
  COND2X1 U6765 ( .A(n7663), .B(n6554), .C(n7194), .D(n6535), .Z(n3820) );
  COND2X1 U6766 ( .A(n7662), .B(n6555), .C(n7193), .D(n6536), .Z(n3821) );
  COND2X1 U6767 ( .A(n7661), .B(n6551), .C(n7192), .D(n6531), .Z(n3822) );
  COND2X1 U6768 ( .A(n7660), .B(n6552), .C(n7191), .D(n6532), .Z(n3823) );
  COND2X1 U6769 ( .A(n7659), .B(n6554), .C(n7190), .D(n6533), .Z(n3824) );
  COND2X1 U6770 ( .A(n7658), .B(n6555), .C(n7189), .D(n6533), .Z(n3825) );
  COND2X1 U6771 ( .A(n7657), .B(n6556), .C(n7188), .D(n6531), .Z(n3826) );
  COND2X1 U6772 ( .A(n7656), .B(n6557), .C(n7187), .D(n6532), .Z(n3827) );
  COND2X1 U6773 ( .A(n7655), .B(n6558), .C(n7186), .D(n6534), .Z(n3828) );
  COND2X1 U6774 ( .A(n7654), .B(n6559), .C(n7185), .D(n6535), .Z(n3829) );
  COND2X1 U6775 ( .A(n7653), .B(n6540), .C(n7184), .D(n6536), .Z(n3830) );
  COND2X1 U6776 ( .A(n7652), .B(n6541), .C(n7183), .D(n6534), .Z(n3831) );
  COND2X1 U6777 ( .A(n7651), .B(n6542), .C(n7182), .D(n6533), .Z(n3832) );
  COND2X1 U6778 ( .A(n7650), .B(n6543), .C(n7181), .D(n6534), .Z(n3833) );
  COND2X1 U6779 ( .A(n7649), .B(n6544), .C(n7180), .D(n6531), .Z(n3834) );
  COND2X1 U6780 ( .A(n7648), .B(n6545), .C(n7179), .D(n6532), .Z(n3835) );
  COND2X1 U6781 ( .A(n7647), .B(n6547), .C(n7178), .D(n6533), .Z(n3836) );
  COND2X1 U6782 ( .A(n7646), .B(n6548), .C(n7177), .D(n6535), .Z(n3837) );
  COND2X1 U6783 ( .A(n7645), .B(n6549), .C(n7176), .D(n6535), .Z(n3838) );
  COND2X1 U6784 ( .A(n7644), .B(n6550), .C(n7175), .D(n6536), .Z(n3839) );
  COND2X1 U6785 ( .A(n7627), .B(n6524), .C(n7190), .D(n6503), .Z(n3856) );
  COND2X1 U6786 ( .A(n7626), .B(n6525), .C(n7189), .D(n6503), .Z(n3857) );
  COND2X1 U6787 ( .A(n7625), .B(n6526), .C(n7188), .D(n6501), .Z(n3858) );
  COND2X1 U6788 ( .A(n7624), .B(n6527), .C(n7187), .D(n6502), .Z(n3859) );
  COND2X1 U6789 ( .A(n7623), .B(n6528), .C(n7186), .D(n6504), .Z(n3860) );
  COND2X1 U6790 ( .A(n7622), .B(n6529), .C(n7185), .D(n6505), .Z(n3861) );
  COND2X1 U6791 ( .A(n7621), .B(n6510), .C(n7184), .D(n6506), .Z(n3862) );
  COND2X1 U6792 ( .A(n7620), .B(n6511), .C(n7183), .D(n6504), .Z(n3863) );
  COND2X1 U6793 ( .A(n7619), .B(n6512), .C(n7182), .D(n6503), .Z(n3864) );
  COND2X1 U6794 ( .A(n7618), .B(n6513), .C(n7181), .D(n6504), .Z(n3865) );
  COND2X1 U6795 ( .A(n7617), .B(n6514), .C(n7180), .D(n6501), .Z(n3866) );
  COND2X1 U6796 ( .A(n7616), .B(n6515), .C(n7179), .D(n6502), .Z(n3867) );
  COND2X1 U6797 ( .A(n7615), .B(n6517), .C(n7178), .D(n6503), .Z(n3868) );
  COND2X1 U6798 ( .A(n7614), .B(n6518), .C(n7177), .D(n6505), .Z(n3869) );
  COND2X1 U6799 ( .A(n7613), .B(n6519), .C(n7176), .D(n6505), .Z(n3870) );
  COND2X1 U6800 ( .A(n7612), .B(n6520), .C(n7175), .D(n6506), .Z(n3871) );
  COND2X1 U6801 ( .A(n7611), .B(n6480), .C(n7206), .D(n6471), .Z(n3872) );
  COND2X1 U6802 ( .A(n7610), .B(n6481), .C(n7205), .D(n6472), .Z(n3873) );
  COND2X1 U6803 ( .A(n7609), .B(n6482), .C(n7204), .D(n6471), .Z(n3874) );
  COND2X1 U6804 ( .A(n7608), .B(n6483), .C(n7203), .D(n6472), .Z(n3875) );
  COND2X1 U6805 ( .A(n7607), .B(n6484), .C(n7202), .D(n6473), .Z(n3876) );
  COND2X1 U6806 ( .A(n7606), .B(n6485), .C(n7201), .D(n6471), .Z(n3877) );
  COND2X1 U6807 ( .A(n7605), .B(n6487), .C(n7200), .D(n6473), .Z(n3878) );
  COND2X1 U6808 ( .A(n7604), .B(n6488), .C(n7199), .D(n6474), .Z(n3879) );
  COND2X1 U6809 ( .A(n7603), .B(n6489), .C(n7198), .D(n6474), .Z(n3880) );
  COND2X1 U6810 ( .A(n7602), .B(n6490), .C(n7197), .D(n6475), .Z(n3881) );
  COND2X1 U6811 ( .A(n7601), .B(n6491), .C(n7196), .D(n6476), .Z(n3882) );
  COND2X1 U6812 ( .A(n7600), .B(n6492), .C(n7195), .D(n6472), .Z(n3883) );
  COND2X1 U6813 ( .A(n7599), .B(n6494), .C(n7194), .D(n6475), .Z(n3884) );
  COND2X1 U6814 ( .A(n7598), .B(n6495), .C(n7193), .D(n6476), .Z(n3885) );
  COND2X1 U6815 ( .A(n7597), .B(n6491), .C(n7192), .D(n6471), .Z(n3886) );
  COND2X1 U6816 ( .A(n7596), .B(n6492), .C(n7191), .D(n6472), .Z(n3887) );
  COND2X1 U6817 ( .A(n7595), .B(n6494), .C(n7190), .D(n6473), .Z(n3888) );
  COND2X1 U6818 ( .A(n7594), .B(n6495), .C(n7189), .D(n6473), .Z(n3889) );
  COND2X1 U6819 ( .A(n7593), .B(n6496), .C(n7188), .D(n6471), .Z(n3890) );
  COND2X1 U6820 ( .A(n7592), .B(n6497), .C(n7187), .D(n6472), .Z(n3891) );
  COND2X1 U6821 ( .A(n7591), .B(n6498), .C(n7186), .D(n6474), .Z(n3892) );
  COND2X1 U6822 ( .A(n7590), .B(n6499), .C(n7185), .D(n6475), .Z(n3893) );
  COND2X1 U6823 ( .A(n7589), .B(n6480), .C(n7184), .D(n6476), .Z(n3894) );
  COND2X1 U6824 ( .A(n7588), .B(n6481), .C(n7183), .D(n6474), .Z(n3895) );
  COND2X1 U6825 ( .A(n7587), .B(n6482), .C(n7182), .D(n6473), .Z(n3896) );
  COND2X1 U6826 ( .A(n7586), .B(n6483), .C(n7181), .D(n6474), .Z(n3897) );
  COND2X1 U6827 ( .A(n7585), .B(n6484), .C(n7180), .D(n6471), .Z(n3898) );
  COND2X1 U6828 ( .A(n7584), .B(n6485), .C(n7179), .D(n6472), .Z(n3899) );
  COND2X1 U6829 ( .A(n7583), .B(n6487), .C(n7178), .D(n6473), .Z(n3900) );
  COND2X1 U6830 ( .A(n7582), .B(n6488), .C(n7177), .D(n6475), .Z(n3901) );
  COND2X1 U6831 ( .A(n7581), .B(n6489), .C(n7176), .D(n6475), .Z(n3902) );
  COND2X1 U6832 ( .A(n7580), .B(n6490), .C(n7175), .D(n6476), .Z(n3903) );
  COND2X1 U6833 ( .A(n7579), .B(n6450), .C(n7206), .D(n6441), .Z(n3904) );
  COND2X1 U6834 ( .A(n7578), .B(n6451), .C(n7205), .D(n6442), .Z(n3905) );
  COND2X1 U6835 ( .A(n7577), .B(n6452), .C(n7204), .D(n6441), .Z(n3906) );
  COND2X1 U6836 ( .A(n7576), .B(n6453), .C(n7203), .D(n6442), .Z(n3907) );
  COND2X1 U6837 ( .A(n7575), .B(n6454), .C(n7202), .D(n6443), .Z(n3908) );
  COND2X1 U6838 ( .A(n7574), .B(n6455), .C(n7201), .D(n6441), .Z(n3909) );
  COND2X1 U6839 ( .A(n7573), .B(n6457), .C(n7200), .D(n6443), .Z(n3910) );
  COND2X1 U6840 ( .A(n7572), .B(n6458), .C(n7199), .D(n6444), .Z(n3911) );
  COND2X1 U6841 ( .A(n7571), .B(n6459), .C(n7198), .D(n6444), .Z(n3912) );
  COND2X1 U6842 ( .A(n7570), .B(n6460), .C(n7197), .D(n6445), .Z(n3913) );
  COND2X1 U6843 ( .A(n7569), .B(n6461), .C(n7196), .D(n6446), .Z(n3914) );
  COND2X1 U6844 ( .A(n7568), .B(n6462), .C(n7195), .D(n6442), .Z(n3915) );
  COND2X1 U6845 ( .A(n7567), .B(n6464), .C(n7194), .D(n6445), .Z(n3916) );
  COND2X1 U6846 ( .A(n7566), .B(n6465), .C(n7193), .D(n6446), .Z(n3917) );
  COND2X1 U6847 ( .A(n7565), .B(n6461), .C(n7192), .D(n6441), .Z(n3918) );
  COND2X1 U6848 ( .A(n7564), .B(n6462), .C(n7191), .D(n6442), .Z(n3919) );
  COND2X1 U6849 ( .A(n7563), .B(n6464), .C(n7190), .D(n6443), .Z(n3920) );
  COND2X1 U6850 ( .A(n7562), .B(n6465), .C(n7189), .D(n6443), .Z(n3921) );
  COND2X1 U6851 ( .A(n7561), .B(n6466), .C(n7188), .D(n6441), .Z(n3922) );
  COND2X1 U6852 ( .A(n7560), .B(n6467), .C(n7187), .D(n6442), .Z(n3923) );
  COND2X1 U6853 ( .A(n7559), .B(n6468), .C(n7186), .D(n6444), .Z(n3924) );
  COND2X1 U6854 ( .A(n7558), .B(n6469), .C(n7185), .D(n6445), .Z(n3925) );
  COND2X1 U6855 ( .A(n7557), .B(n6450), .C(n7184), .D(n6446), .Z(n3926) );
  COND2X1 U6856 ( .A(n7556), .B(n6451), .C(n7183), .D(n6444), .Z(n3927) );
  COND2X1 U6857 ( .A(n7555), .B(n6452), .C(n7182), .D(n6443), .Z(n3928) );
  COND2X1 U6858 ( .A(n7554), .B(n6453), .C(n7181), .D(n6444), .Z(n3929) );
  COND2X1 U6859 ( .A(n7553), .B(n6454), .C(n7180), .D(n6441), .Z(n3930) );
  COND2X1 U6860 ( .A(n7552), .B(n6455), .C(n7179), .D(n6442), .Z(n3931) );
  COND2X1 U6861 ( .A(n7551), .B(n6457), .C(n7178), .D(n6443), .Z(n3932) );
  COND2X1 U6862 ( .A(n7550), .B(n6458), .C(n7177), .D(n6445), .Z(n3933) );
  COND2X1 U6863 ( .A(n7549), .B(n6459), .C(n7176), .D(n6445), .Z(n3934) );
  COND2X1 U6864 ( .A(n7548), .B(n6460), .C(n7175), .D(n6446), .Z(n3935) );
  COND2X1 U6865 ( .A(n7547), .B(n6420), .C(n7206), .D(n6411), .Z(n3936) );
  COND2X1 U6866 ( .A(n7546), .B(n6421), .C(n7205), .D(n6412), .Z(n3937) );
  COND2X1 U6867 ( .A(n7545), .B(n6422), .C(n7204), .D(n6411), .Z(n3938) );
  COND2X1 U6868 ( .A(n7544), .B(n6423), .C(n7203), .D(n6412), .Z(n3939) );
  COND2X1 U6869 ( .A(n7543), .B(n6424), .C(n7202), .D(n6413), .Z(n3940) );
  COND2X1 U6870 ( .A(n7542), .B(n6425), .C(n7201), .D(n6411), .Z(n3941) );
  COND2X1 U6871 ( .A(n7541), .B(n6427), .C(n7200), .D(n6413), .Z(n3942) );
  COND2X1 U6872 ( .A(n7540), .B(n6428), .C(n7199), .D(n6414), .Z(n3943) );
  COND2X1 U6873 ( .A(n7539), .B(n6429), .C(n7198), .D(n6414), .Z(n3944) );
  COND2X1 U6874 ( .A(n7538), .B(n6430), .C(n7197), .D(n6415), .Z(n3945) );
  COND2X1 U6875 ( .A(n7537), .B(n6431), .C(n7196), .D(n6416), .Z(n3946) );
  COND2X1 U6876 ( .A(n7536), .B(n6432), .C(n7195), .D(n6412), .Z(n3947) );
  COND2X1 U6877 ( .A(n7535), .B(n6434), .C(n7194), .D(n6415), .Z(n3948) );
  COND2X1 U6878 ( .A(n7534), .B(n6435), .C(n7193), .D(n6416), .Z(n3949) );
  COND2X1 U6879 ( .A(n7533), .B(n6431), .C(n7192), .D(n6411), .Z(n3950) );
  COND2X1 U6880 ( .A(n7532), .B(n6432), .C(n7191), .D(n6412), .Z(n3951) );
  COND2X1 U6881 ( .A(n7531), .B(n6434), .C(n7190), .D(n6413), .Z(n3952) );
  COND2X1 U6882 ( .A(n7530), .B(n6435), .C(n7189), .D(n6413), .Z(n3953) );
  COND2X1 U6883 ( .A(n7529), .B(n6436), .C(n7188), .D(n6411), .Z(n3954) );
  COND2X1 U6884 ( .A(n7528), .B(n6437), .C(n7187), .D(n6412), .Z(n3955) );
  COND2X1 U6885 ( .A(n7527), .B(n6438), .C(n7186), .D(n6414), .Z(n3956) );
  COND2X1 U6886 ( .A(n7526), .B(n6439), .C(n7185), .D(n6415), .Z(n3957) );
  COND2X1 U6887 ( .A(n7525), .B(n6420), .C(n7184), .D(n6416), .Z(n3958) );
  COND2X1 U6888 ( .A(n7524), .B(n6421), .C(n7183), .D(n6414), .Z(n3959) );
  COND2X1 U6889 ( .A(n7523), .B(n6422), .C(n7182), .D(n6413), .Z(n3960) );
  COND2X1 U6890 ( .A(n7522), .B(n6423), .C(n7181), .D(n6414), .Z(n3961) );
  COND2X1 U6891 ( .A(n7521), .B(n6424), .C(n7180), .D(n6411), .Z(n3962) );
  COND2X1 U6892 ( .A(n7520), .B(n6425), .C(n7179), .D(n6412), .Z(n3963) );
  COND2X1 U6893 ( .A(n7519), .B(n6427), .C(n7178), .D(n6413), .Z(n3964) );
  COND2X1 U6894 ( .A(n7518), .B(n6428), .C(n7177), .D(n6415), .Z(n3965) );
  COND2X1 U6895 ( .A(n7517), .B(n6429), .C(n7176), .D(n6415), .Z(n3966) );
  COND2X1 U6896 ( .A(n7516), .B(n6430), .C(n7175), .D(n6416), .Z(n3967) );
  COND2X1 U6897 ( .A(n7499), .B(n6404), .C(n7190), .D(n6383), .Z(n3984) );
  COND2X1 U6898 ( .A(n7498), .B(n6405), .C(n7189), .D(n6383), .Z(n3985) );
  COND2X1 U6899 ( .A(n7497), .B(n6406), .C(n7188), .D(n6381), .Z(n3986) );
  COND2X1 U6900 ( .A(n7496), .B(n6407), .C(n7187), .D(n6382), .Z(n3987) );
  COND2X1 U6901 ( .A(n7495), .B(n6408), .C(n7186), .D(n6384), .Z(n3988) );
  COND2X1 U6902 ( .A(n7494), .B(n6409), .C(n7185), .D(n6385), .Z(n3989) );
  COND2X1 U6903 ( .A(n7493), .B(n6390), .C(n7184), .D(n6386), .Z(n3990) );
  COND2X1 U6904 ( .A(n7492), .B(n6391), .C(n7183), .D(n6384), .Z(n3991) );
  COND2X1 U6905 ( .A(n7491), .B(n6392), .C(n7182), .D(n6383), .Z(n3992) );
  COND2X1 U6906 ( .A(n7490), .B(n6393), .C(n7181), .D(n6384), .Z(n3993) );
  COND2X1 U6907 ( .A(n7489), .B(n6394), .C(n7180), .D(n6381), .Z(n3994) );
  COND2X1 U6908 ( .A(n7488), .B(n6395), .C(n7179), .D(n6382), .Z(n3995) );
  COND2X1 U6909 ( .A(n7487), .B(n6397), .C(n7178), .D(n6383), .Z(n3996) );
  COND2X1 U6910 ( .A(n7486), .B(n6398), .C(n7177), .D(n6385), .Z(n3997) );
  COND2X1 U6911 ( .A(n7485), .B(n6399), .C(n7176), .D(n6385), .Z(n3998) );
  COND2X1 U6912 ( .A(n7484), .B(n6400), .C(n7175), .D(n6386), .Z(n3999) );
  COND2X1 U6913 ( .A(n7483), .B(n6360), .C(n7206), .D(n6351), .Z(n4000) );
  COND2X1 U6914 ( .A(n7482), .B(n6361), .C(n7205), .D(n6352), .Z(n4001) );
  COND2X1 U6915 ( .A(n7481), .B(n6362), .C(n7204), .D(n6351), .Z(n4002) );
  COND2X1 U6916 ( .A(n7480), .B(n6363), .C(n7203), .D(n6352), .Z(n4003) );
  COND2X1 U6917 ( .A(n7479), .B(n6364), .C(n7202), .D(n6353), .Z(n4004) );
  COND2X1 U6918 ( .A(n7478), .B(n6365), .C(n7201), .D(n6351), .Z(n4005) );
  COND2X1 U6919 ( .A(n7477), .B(n6367), .C(n7200), .D(n6353), .Z(n4006) );
  COND2X1 U6920 ( .A(n7476), .B(n6368), .C(n7199), .D(n6354), .Z(n4007) );
  COND2X1 U6921 ( .A(n7475), .B(n6369), .C(n7198), .D(n6354), .Z(n4008) );
  COND2X1 U6922 ( .A(n7474), .B(n6370), .C(n7197), .D(n6355), .Z(n4009) );
  COND2X1 U6923 ( .A(n7473), .B(n6371), .C(n7196), .D(n6356), .Z(n4010) );
  COND2X1 U6924 ( .A(n7472), .B(n6372), .C(n7195), .D(n6352), .Z(n4011) );
  COND2X1 U6925 ( .A(n7471), .B(n6374), .C(n7194), .D(n6355), .Z(n4012) );
  COND2X1 U6926 ( .A(n7470), .B(n6375), .C(n7193), .D(n6356), .Z(n4013) );
  COND2X1 U6927 ( .A(n7469), .B(n6371), .C(n7192), .D(n6351), .Z(n4014) );
  COND2X1 U6928 ( .A(n7468), .B(n6372), .C(n7191), .D(n6352), .Z(n4015) );
  COND2X1 U6929 ( .A(n7467), .B(n6374), .C(n7190), .D(n6353), .Z(n4016) );
  COND2X1 U6930 ( .A(n7466), .B(n6375), .C(n7189), .D(n6353), .Z(n4017) );
  COND2X1 U6931 ( .A(n7465), .B(n6376), .C(n7188), .D(n6351), .Z(n4018) );
  COND2X1 U6932 ( .A(n7464), .B(n6377), .C(n7187), .D(n6352), .Z(n4019) );
  COND2X1 U6933 ( .A(n7463), .B(n6378), .C(n7186), .D(n6354), .Z(n4020) );
  COND2X1 U6934 ( .A(n7462), .B(n6379), .C(n7185), .D(n6355), .Z(n4021) );
  COND2X1 U6935 ( .A(n7461), .B(n6360), .C(n7184), .D(n6356), .Z(n4022) );
  COND2X1 U6936 ( .A(n7460), .B(n6361), .C(n7183), .D(n6354), .Z(n4023) );
  COND2X1 U6937 ( .A(n7459), .B(n6362), .C(n7182), .D(n6353), .Z(n4024) );
  COND2X1 U6938 ( .A(n7458), .B(n6363), .C(n7181), .D(n6354), .Z(n4025) );
  COND2X1 U6939 ( .A(n7457), .B(n6364), .C(n7180), .D(n6351), .Z(n4026) );
  COND2X1 U6940 ( .A(n7456), .B(n6365), .C(n7179), .D(n6352), .Z(n4027) );
  COND2X1 U6941 ( .A(n7455), .B(n6367), .C(n7178), .D(n6353), .Z(n4028) );
  COND2X1 U6942 ( .A(n7454), .B(n6368), .C(n7177), .D(n6355), .Z(n4029) );
  COND2X1 U6943 ( .A(n7453), .B(n6369), .C(n7176), .D(n6355), .Z(n4030) );
  COND2X1 U6944 ( .A(n7452), .B(n6370), .C(n7175), .D(n6356), .Z(n4031) );
  COND2X1 U6945 ( .A(n7451), .B(n6330), .C(n7206), .D(n6321), .Z(n4032) );
  COND2X1 U6946 ( .A(n7450), .B(n6331), .C(n7205), .D(n6322), .Z(n4033) );
  COND2X1 U6947 ( .A(n7449), .B(n6332), .C(n7204), .D(n6321), .Z(n4034) );
  COND2X1 U6948 ( .A(n7448), .B(n6333), .C(n7203), .D(n6322), .Z(n4035) );
  COND2X1 U6949 ( .A(n7447), .B(n6334), .C(n7202), .D(n6323), .Z(n4036) );
  COND2X1 U6950 ( .A(n7446), .B(n6335), .C(n7201), .D(n6321), .Z(n4037) );
  COND2X1 U6951 ( .A(n7445), .B(n6337), .C(n7200), .D(n6323), .Z(n4038) );
  COND2X1 U6952 ( .A(n7444), .B(n6338), .C(n7199), .D(n6324), .Z(n4039) );
  COND2X1 U6953 ( .A(n7443), .B(n6339), .C(n7198), .D(n6324), .Z(n4040) );
  COND2X1 U6954 ( .A(n7442), .B(n6340), .C(n7197), .D(n6325), .Z(n4041) );
  COND2X1 U6955 ( .A(n7441), .B(n6341), .C(n7196), .D(n6326), .Z(n4042) );
  COND2X1 U6956 ( .A(n7440), .B(n6342), .C(n7195), .D(n6322), .Z(n4043) );
  COND2X1 U6957 ( .A(n7439), .B(n6344), .C(n7194), .D(n6325), .Z(n4044) );
  COND2X1 U6958 ( .A(n7438), .B(n6345), .C(n7193), .D(n6326), .Z(n4045) );
  COND2X1 U6959 ( .A(n7437), .B(n6341), .C(n7192), .D(n6321), .Z(n4046) );
  COND2X1 U6960 ( .A(n7436), .B(n6342), .C(n7191), .D(n6322), .Z(n4047) );
  COND2X1 U6961 ( .A(n7435), .B(n6344), .C(n7190), .D(n6323), .Z(n4048) );
  COND2X1 U6962 ( .A(n7434), .B(n6345), .C(n7189), .D(n6323), .Z(n4049) );
  COND2X1 U6963 ( .A(n7433), .B(n6346), .C(n7188), .D(n6321), .Z(n4050) );
  COND2X1 U6964 ( .A(n7432), .B(n6347), .C(n7187), .D(n6322), .Z(n4051) );
  COND2X1 U6965 ( .A(n7431), .B(n6348), .C(n7186), .D(n6324), .Z(n4052) );
  COND2X1 U6966 ( .A(n7430), .B(n6349), .C(n7185), .D(n6325), .Z(n4053) );
  COND2X1 U6967 ( .A(n7429), .B(n6330), .C(n7184), .D(n6326), .Z(n4054) );
  COND2X1 U6968 ( .A(n7428), .B(n6331), .C(n7183), .D(n6324), .Z(n4055) );
  COND2X1 U6969 ( .A(n7427), .B(n6332), .C(n7182), .D(n6323), .Z(n4056) );
  COND2X1 U6970 ( .A(n7426), .B(n6333), .C(n7181), .D(n6324), .Z(n4057) );
  COND2X1 U6971 ( .A(n7425), .B(n6334), .C(n7180), .D(n6321), .Z(n4058) );
  COND2X1 U6972 ( .A(n7424), .B(n6335), .C(n7179), .D(n6322), .Z(n4059) );
  COND2X1 U6973 ( .A(n7423), .B(n6337), .C(n7178), .D(n6323), .Z(n4060) );
  COND2X1 U6974 ( .A(n7422), .B(n6338), .C(n7177), .D(n6325), .Z(n4061) );
  COND2X1 U6975 ( .A(n7421), .B(n6339), .C(n7176), .D(n6325), .Z(n4062) );
  COND2X1 U6976 ( .A(n7420), .B(n6340), .C(n7175), .D(n6326), .Z(n4063) );
  COND2X1 U6977 ( .A(n7419), .B(n6300), .C(n7206), .D(n6291), .Z(n4064) );
  COND2X1 U6978 ( .A(n7418), .B(n6301), .C(n7205), .D(n6292), .Z(n4065) );
  COND2X1 U6979 ( .A(n7417), .B(n6302), .C(n7204), .D(n6291), .Z(n4066) );
  COND2X1 U6980 ( .A(n7416), .B(n6303), .C(n7203), .D(n6292), .Z(n4067) );
  COND2X1 U6981 ( .A(n7415), .B(n6304), .C(n7202), .D(n6293), .Z(n4068) );
  COND2X1 U6982 ( .A(n7414), .B(n6305), .C(n7201), .D(n6291), .Z(n4069) );
  COND2X1 U6983 ( .A(n7413), .B(n6307), .C(n7200), .D(n6293), .Z(n4070) );
  COND2X1 U6984 ( .A(n7412), .B(n6308), .C(n7199), .D(n6294), .Z(n4071) );
  COND2X1 U6985 ( .A(n7411), .B(n6309), .C(n7198), .D(n6294), .Z(n4072) );
  COND2X1 U6986 ( .A(n7410), .B(n6310), .C(n7197), .D(n6295), .Z(n4073) );
  COND2X1 U6987 ( .A(n7409), .B(n6311), .C(n7196), .D(n6296), .Z(n4074) );
  COND2X1 U6988 ( .A(n7408), .B(n6312), .C(n7195), .D(n6292), .Z(n4075) );
  COND2X1 U6989 ( .A(n7407), .B(n6314), .C(n7194), .D(n6295), .Z(n4076) );
  COND2X1 U6990 ( .A(n7406), .B(n6315), .C(n7193), .D(n6296), .Z(n4077) );
  COND2X1 U6991 ( .A(n7405), .B(n6311), .C(n7192), .D(n6291), .Z(n4078) );
  COND2X1 U6992 ( .A(n7404), .B(n6312), .C(n7191), .D(n6292), .Z(n4079) );
  COND2X1 U6993 ( .A(n7403), .B(n6314), .C(n7190), .D(n6293), .Z(n4080) );
  COND2X1 U6994 ( .A(n7402), .B(n6315), .C(n7189), .D(n6293), .Z(n4081) );
  COND2X1 U6995 ( .A(n7401), .B(n6316), .C(n7188), .D(n6291), .Z(n4082) );
  COND2X1 U6996 ( .A(n7400), .B(n6317), .C(n7187), .D(n6292), .Z(n4083) );
  COND2X1 U6997 ( .A(n7399), .B(n6318), .C(n7186), .D(n6294), .Z(n4084) );
  COND2X1 U6998 ( .A(n7398), .B(n6319), .C(n7185), .D(n6295), .Z(n4085) );
  COND2X1 U6999 ( .A(n7397), .B(n6300), .C(n7184), .D(n6296), .Z(n4086) );
  COND2X1 U7000 ( .A(n7396), .B(n6301), .C(n7183), .D(n6294), .Z(n4087) );
  COND2X1 U7001 ( .A(n7395), .B(n6302), .C(n7182), .D(n6293), .Z(n4088) );
  COND2X1 U7002 ( .A(n7394), .B(n6303), .C(n7181), .D(n6294), .Z(n4089) );
  COND2X1 U7003 ( .A(n7393), .B(n6304), .C(n7180), .D(n6291), .Z(n4090) );
  COND2X1 U7004 ( .A(n7392), .B(n6305), .C(n7179), .D(n6292), .Z(n4091) );
  COND2X1 U7005 ( .A(n7391), .B(n6307), .C(n7178), .D(n6293), .Z(n4092) );
  COND2X1 U7006 ( .A(n7390), .B(n6308), .C(n7177), .D(n6295), .Z(n4093) );
  COND2X1 U7007 ( .A(n7389), .B(n6309), .C(n7176), .D(n6295), .Z(n4094) );
  COND2X1 U7008 ( .A(n7388), .B(n6310), .C(n7175), .D(n6296), .Z(n4095) );
  COND2X1 U7009 ( .A(n7371), .B(n6284), .C(n7190), .D(n6263), .Z(n4112) );
  COND2X1 U7010 ( .A(n7370), .B(n6285), .C(n7189), .D(n6263), .Z(n4113) );
  COND2X1 U7011 ( .A(n7369), .B(n6286), .C(n7188), .D(n6261), .Z(n4114) );
  COND2X1 U7012 ( .A(n7368), .B(n6287), .C(n7187), .D(n6262), .Z(n4115) );
  COND2X1 U7013 ( .A(n7367), .B(n6288), .C(n7186), .D(n6264), .Z(n4116) );
  COND2X1 U7014 ( .A(n7366), .B(n6289), .C(n7185), .D(n6265), .Z(n4117) );
  COND2X1 U7015 ( .A(n7365), .B(n6270), .C(n7184), .D(n6266), .Z(n4118) );
  COND2X1 U7016 ( .A(n7364), .B(n6271), .C(n7183), .D(n6264), .Z(n4119) );
  COND2X1 U7017 ( .A(n7363), .B(n6272), .C(n7182), .D(n6263), .Z(n4120) );
  COND2X1 U7018 ( .A(n7362), .B(n6273), .C(n7181), .D(n6264), .Z(n4121) );
  COND2X1 U7019 ( .A(n7361), .B(n6274), .C(n7180), .D(n6261), .Z(n4122) );
  COND2X1 U7020 ( .A(n7360), .B(n6275), .C(n7179), .D(n6262), .Z(n4123) );
  COND2X1 U7021 ( .A(n7359), .B(n6277), .C(n7178), .D(n6263), .Z(n4124) );
  COND2X1 U7022 ( .A(n7358), .B(n6278), .C(n7177), .D(n6265), .Z(n4125) );
  COND2X1 U7023 ( .A(n7357), .B(n6279), .C(n7176), .D(n6265), .Z(n4126) );
  COND2X1 U7024 ( .A(n7356), .B(n6280), .C(n7175), .D(n6266), .Z(n4127) );
  COND2X1 U7025 ( .A(n7355), .B(n6240), .C(n7206), .D(n6231), .Z(n4128) );
  COND2X1 U7026 ( .A(n7354), .B(n6241), .C(n7205), .D(n6232), .Z(n4129) );
  COND2X1 U7027 ( .A(n7353), .B(n6242), .C(n7204), .D(n6231), .Z(n4130) );
  COND2X1 U7028 ( .A(n7352), .B(n6243), .C(n7203), .D(n6232), .Z(n4131) );
  COND2X1 U7029 ( .A(n7351), .B(n6244), .C(n7202), .D(n6233), .Z(n4132) );
  COND2X1 U7030 ( .A(n7350), .B(n6245), .C(n7201), .D(n6231), .Z(n4133) );
  COND2X1 U7031 ( .A(n7349), .B(n6247), .C(n7200), .D(n6233), .Z(n4134) );
  COND2X1 U7032 ( .A(n7348), .B(n6248), .C(n7199), .D(n6234), .Z(n4135) );
  COND2X1 U7033 ( .A(n7347), .B(n6249), .C(n7198), .D(n6234), .Z(n4136) );
  COND2X1 U7034 ( .A(n7346), .B(n6250), .C(n7197), .D(n6235), .Z(n4137) );
  COND2X1 U7035 ( .A(n7345), .B(n6251), .C(n7196), .D(n6236), .Z(n4138) );
  COND2X1 U7036 ( .A(n7344), .B(n6252), .C(n7195), .D(n6232), .Z(n4139) );
  COND2X1 U7037 ( .A(n7343), .B(n6254), .C(n7194), .D(n6235), .Z(n4140) );
  COND2X1 U7038 ( .A(n7342), .B(n6255), .C(n7193), .D(n6236), .Z(n4141) );
  COND2X1 U7039 ( .A(n7341), .B(n6251), .C(n7192), .D(n6231), .Z(n4142) );
  COND2X1 U7040 ( .A(n7340), .B(n6252), .C(n7191), .D(n6232), .Z(n4143) );
  COND2X1 U7041 ( .A(n7339), .B(n6254), .C(n7190), .D(n6233), .Z(n4144) );
  COND2X1 U7042 ( .A(n7338), .B(n6255), .C(n7189), .D(n6233), .Z(n4145) );
  COND2X1 U7043 ( .A(n7337), .B(n6256), .C(n7188), .D(n6231), .Z(n4146) );
  COND2X1 U7044 ( .A(n7336), .B(n6257), .C(n7187), .D(n6232), .Z(n4147) );
  COND2X1 U7045 ( .A(n7335), .B(n6258), .C(n7186), .D(n6234), .Z(n4148) );
  COND2X1 U7046 ( .A(n7334), .B(n6259), .C(n7185), .D(n6235), .Z(n4149) );
  COND2X1 U7047 ( .A(n7333), .B(n6240), .C(n7184), .D(n6236), .Z(n4150) );
  COND2X1 U7048 ( .A(n7332), .B(n6241), .C(n7183), .D(n6234), .Z(n4151) );
  COND2X1 U7049 ( .A(n7331), .B(n6242), .C(n7182), .D(n6233), .Z(n4152) );
  COND2X1 U7050 ( .A(n7330), .B(n6243), .C(n7181), .D(n6234), .Z(n4153) );
  COND2X1 U7051 ( .A(n7329), .B(n6244), .C(n7180), .D(n6231), .Z(n4154) );
  COND2X1 U7052 ( .A(n7328), .B(n6245), .C(n7179), .D(n6232), .Z(n4155) );
  COND2X1 U7053 ( .A(n7327), .B(n6247), .C(n7178), .D(n6233), .Z(n4156) );
  COND2X1 U7054 ( .A(n7326), .B(n6248), .C(n7177), .D(n6235), .Z(n4157) );
  COND2X1 U7055 ( .A(n7325), .B(n6249), .C(n7176), .D(n6235), .Z(n4158) );
  COND2X1 U7056 ( .A(n7324), .B(n6250), .C(n7175), .D(n6236), .Z(n4159) );
  COND2X1 U7057 ( .A(n7323), .B(n6210), .C(n7206), .D(n6201), .Z(n4160) );
  COND2X1 U7058 ( .A(n7322), .B(n6211), .C(n7205), .D(n6202), .Z(n4161) );
  COND2X1 U7059 ( .A(n7321), .B(n6212), .C(n7204), .D(n6201), .Z(n4162) );
  COND2X1 U7060 ( .A(n7320), .B(n6213), .C(n7203), .D(n6202), .Z(n4163) );
  COND2X1 U7061 ( .A(n7319), .B(n6214), .C(n7202), .D(n6203), .Z(n4164) );
  COND2X1 U7062 ( .A(n7318), .B(n6215), .C(n7201), .D(n6201), .Z(n4165) );
  COND2X1 U7063 ( .A(n7317), .B(n6217), .C(n7200), .D(n6203), .Z(n4166) );
  COND2X1 U7064 ( .A(n7316), .B(n6218), .C(n7199), .D(n6204), .Z(n4167) );
  COND2X1 U7065 ( .A(n7315), .B(n6219), .C(n7198), .D(n6204), .Z(n4168) );
  COND2X1 U7066 ( .A(n7314), .B(n6220), .C(n7197), .D(n6205), .Z(n4169) );
  COND2X1 U7067 ( .A(n7313), .B(n6221), .C(n7196), .D(n6206), .Z(n4170) );
  COND2X1 U7068 ( .A(n7312), .B(n6222), .C(n7195), .D(n6202), .Z(n4171) );
  COND2X1 U7069 ( .A(n7311), .B(n6224), .C(n7194), .D(n6205), .Z(n4172) );
  COND2X1 U7070 ( .A(n7310), .B(n6225), .C(n7193), .D(n6206), .Z(n4173) );
  COND2X1 U7071 ( .A(n7309), .B(n6221), .C(n7192), .D(n6201), .Z(n4174) );
  COND2X1 U7072 ( .A(n7308), .B(n6222), .C(n7191), .D(n6202), .Z(n4175) );
  COND2X1 U7073 ( .A(n7307), .B(n6224), .C(n7190), .D(n6203), .Z(n4176) );
  COND2X1 U7074 ( .A(n7306), .B(n6225), .C(n7189), .D(n6203), .Z(n4177) );
  COND2X1 U7075 ( .A(n7305), .B(n6226), .C(n7188), .D(n6201), .Z(n4178) );
  COND2X1 U7076 ( .A(n7304), .B(n6227), .C(n7187), .D(n6202), .Z(n4179) );
  COND2X1 U7077 ( .A(n7303), .B(n6228), .C(n7186), .D(n6204), .Z(n4180) );
  COND2X1 U7078 ( .A(n7302), .B(n6229), .C(n7185), .D(n6205), .Z(n4181) );
  COND2X1 U7079 ( .A(n7301), .B(n6210), .C(n7184), .D(n6206), .Z(n4182) );
  COND2X1 U7080 ( .A(n7300), .B(n6211), .C(n7183), .D(n6204), .Z(n4183) );
  COND2X1 U7081 ( .A(n7299), .B(n6212), .C(n7182), .D(n6203), .Z(n4184) );
  COND2X1 U7082 ( .A(n7298), .B(n6213), .C(n7181), .D(n6204), .Z(n4185) );
  COND2X1 U7083 ( .A(n7297), .B(n6214), .C(n7180), .D(n6201), .Z(n4186) );
  COND2X1 U7084 ( .A(n7296), .B(n6215), .C(n7179), .D(n6202), .Z(n4187) );
  COND2X1 U7085 ( .A(n7295), .B(n6217), .C(n7178), .D(n6203), .Z(n4188) );
  COND2X1 U7086 ( .A(n7294), .B(n6218), .C(n7177), .D(n6205), .Z(n4189) );
  COND2X1 U7087 ( .A(n7293), .B(n6219), .C(n7176), .D(n6205), .Z(n4190) );
  COND2X1 U7088 ( .A(n7292), .B(n6220), .C(n7175), .D(n6206), .Z(n4191) );
  COND2X1 U7089 ( .A(n7291), .B(n6180), .C(n7206), .D(n6171), .Z(n4192) );
  COND2X1 U7090 ( .A(n7290), .B(n6181), .C(n7205), .D(n6172), .Z(n4193) );
  COND2X1 U7091 ( .A(n7289), .B(n6182), .C(n7204), .D(n6171), .Z(n4194) );
  COND2X1 U7092 ( .A(n7288), .B(n6183), .C(n7203), .D(n6172), .Z(n4195) );
  COND2X1 U7093 ( .A(n7287), .B(n6184), .C(n7202), .D(n6173), .Z(n4196) );
  COND2X1 U7094 ( .A(n7286), .B(n6185), .C(n7201), .D(n6171), .Z(n4197) );
  COND2X1 U7095 ( .A(n7285), .B(n6187), .C(n7200), .D(n6173), .Z(n4198) );
  COND2X1 U7096 ( .A(n7284), .B(n6188), .C(n7199), .D(n6174), .Z(n4199) );
  COND2X1 U7097 ( .A(n7283), .B(n6189), .C(n7198), .D(n6174), .Z(n4200) );
  COND2X1 U7098 ( .A(n7282), .B(n6190), .C(n7197), .D(n6175), .Z(n4201) );
  COND2X1 U7099 ( .A(n7280), .B(n6191), .C(n7196), .D(n6176), .Z(n4202) );
  COND2X1 U7100 ( .A(n7278), .B(n6192), .C(n7195), .D(n6172), .Z(n4203) );
  COND2X1 U7101 ( .A(n7276), .B(n6194), .C(n7194), .D(n6175), .Z(n4204) );
  COND2X1 U7102 ( .A(n7275), .B(n6195), .C(n7193), .D(n6176), .Z(n4205) );
  COND2X1 U7103 ( .A(n7271), .B(n6194), .C(n7190), .D(n6173), .Z(n4208) );
  COND2X1 U7104 ( .A(n7269), .B(n6195), .C(n7189), .D(n6173), .Z(n4209) );
  COND2X1 U7105 ( .A(n7267), .B(n6196), .C(n7188), .D(n6171), .Z(n4210) );
  COND2X1 U7106 ( .A(n7266), .B(n6197), .C(n7187), .D(n6172), .Z(n4211) );
  COND2X1 U7107 ( .A(n7264), .B(n6198), .C(n7186), .D(n6174), .Z(n4212) );
  COND2X1 U7108 ( .A(n7262), .B(n6199), .C(n7185), .D(n6175), .Z(n4213) );
  COND2X1 U7109 ( .A(n7261), .B(n6180), .C(n7184), .D(n6176), .Z(n4214) );
  COND2X1 U7110 ( .A(n7260), .B(n6181), .C(n7183), .D(n6174), .Z(n4215) );
  COND2X1 U7111 ( .A(n7259), .B(n6182), .C(n7182), .D(n6173), .Z(n4216) );
  COND2X1 U7112 ( .A(n7257), .B(n6183), .C(n7181), .D(n6174), .Z(n4217) );
  COND2X1 U7113 ( .A(n7256), .B(n6184), .C(n7180), .D(n6171), .Z(n4218) );
  COND2X1 U7114 ( .A(n7255), .B(n6185), .C(n7179), .D(n6172), .Z(n4219) );
  COND2X1 U7115 ( .A(n7254), .B(n6187), .C(n7178), .D(n6173), .Z(n4220) );
  COND2X1 U7116 ( .A(n7253), .B(n6188), .C(n7177), .D(n6175), .Z(n4221) );
  COND2X1 U7117 ( .A(n7251), .B(n6189), .C(n7176), .D(n6175), .Z(n4222) );
  COND2X1 U7118 ( .A(n7248), .B(n6190), .C(n7175), .D(n6176), .Z(n4223) );
  COND2X1 U7119 ( .A(n7225), .B(n7108), .C(n6168), .D(n7194), .Z(n4236) );
  COND2X1 U7120 ( .A(n8143), .B(n6995), .C(n7194), .D(n6976), .Z(n3340) );
  COND2X1 U7121 ( .A(n7887), .B(n6755), .C(n7194), .D(n6736), .Z(n3596) );
  COND2X1 U7122 ( .A(n7631), .B(n6524), .C(n7194), .D(n6505), .Z(n3852) );
  COND2X1 U7123 ( .A(n7503), .B(n6404), .C(n7194), .D(n6385), .Z(n3980) );
  COND2X1 U7124 ( .A(n7375), .B(n6284), .C(n7194), .D(n6265), .Z(n4108) );
  CNR2X1 U7125 ( .A(n6161), .B(n6160), .Z(n99) );
  CIVX2 U7126 ( .A(n97), .Z(n7171) );
  CND2X1 U7127 ( .A(n8290), .B(n8287), .Z(n14) );
  CND2X1 U7128 ( .A(n6161), .B(n6160), .Z(n178) );
  CND2X1 U7129 ( .A(n6163), .B(n6162), .Z(n10) );
  CIVX2 U7130 ( .A(n65), .Z(n8295) );
  CIVX2 U7131 ( .A(n29), .Z(n8294) );
  CND2X1 U7132 ( .A(n2057), .B(n2058), .Z(n2056) );
  CND2X1 U7133 ( .A(n2057), .B(n2058), .Z(n7061) );
  CND2X1 U7134 ( .A(n2061), .B(n2062), .Z(n2060) );
  CND2X1 U7135 ( .A(n2061), .B(n2062), .Z(n7031) );
  CND2X1 U7136 ( .A(n2061), .B(n2057), .Z(n2064) );
  CND2X1 U7137 ( .A(n2061), .B(n2057), .Z(n7001) );
  CND2X1 U7138 ( .A(n2082), .B(n2062), .Z(n2067) );
  CND2X1 U7139 ( .A(n2082), .B(n2062), .Z(n6971) );
  CND2X1 U7140 ( .A(n2082), .B(n2057), .Z(n2084) );
  CND2X1 U7141 ( .A(n2082), .B(n2057), .Z(n6941) );
  CND2X1 U7142 ( .A(n2087), .B(n2062), .Z(n2086) );
  CND2X1 U7143 ( .A(n2087), .B(n2062), .Z(n6911) );
  CND2X1 U7144 ( .A(n2087), .B(n2057), .Z(n2089) );
  CND2X1 U7145 ( .A(n2087), .B(n2057), .Z(n6881) );
  CND2X1 U7146 ( .A(n2107), .B(n2062), .Z(n2094) );
  CND2X1 U7147 ( .A(n2107), .B(n2062), .Z(n6851) );
  CND2X1 U7148 ( .A(n2107), .B(n2057), .Z(n2109) );
  CND2X1 U7149 ( .A(n2107), .B(n2057), .Z(n6821) );
  CND2X1 U7150 ( .A(n2112), .B(n2062), .Z(n2111) );
  CND2X1 U7151 ( .A(n2112), .B(n2062), .Z(n6791) );
  CND2X1 U7152 ( .A(n2112), .B(n2057), .Z(n2114) );
  CND2X1 U7153 ( .A(n2112), .B(n2057), .Z(n6761) );
  CND2X1 U7154 ( .A(n2130), .B(n2062), .Z(n2117) );
  CND2X1 U7155 ( .A(n2130), .B(n2062), .Z(n6731) );
  CND2X1 U7156 ( .A(n2155), .B(n2058), .Z(n2141) );
  CND2X1 U7157 ( .A(n2155), .B(n2058), .Z(n6620) );
  CND2X1 U7158 ( .A(n2158), .B(n2058), .Z(n2157) );
  CND2X1 U7159 ( .A(n2158), .B(n2058), .Z(n6590) );
  CND2X1 U7160 ( .A(n2155), .B(n2061), .Z(n2160) );
  CND2X1 U7161 ( .A(n2155), .B(n2061), .Z(n6560) );
  CND2X1 U7162 ( .A(n2158), .B(n2061), .Z(n2162) );
  CND2X1 U7163 ( .A(n2158), .B(n2061), .Z(n6530) );
  CND2X1 U7164 ( .A(n2155), .B(n2082), .Z(n2165) );
  CND2X1 U7165 ( .A(n2155), .B(n2082), .Z(n6500) );
  CND2X1 U7166 ( .A(n2158), .B(n2082), .Z(n2169) );
  CND2X1 U7167 ( .A(n2158), .B(n2082), .Z(n6470) );
  CND2X1 U7168 ( .A(n2155), .B(n2087), .Z(n2172) );
  CND2X1 U7169 ( .A(n2155), .B(n2087), .Z(n6440) );
  CND2X1 U7170 ( .A(n2158), .B(n2087), .Z(n2174) );
  CND2X1 U7171 ( .A(n2158), .B(n2087), .Z(n6410) );
  CND2X1 U7172 ( .A(n2155), .B(n2107), .Z(n2177) );
  CND2X1 U7173 ( .A(n2155), .B(n2107), .Z(n6380) );
  CND2X1 U7174 ( .A(n2158), .B(n2107), .Z(n2192) );
  CND2X1 U7175 ( .A(n2158), .B(n2107), .Z(n6350) );
  CND2X1 U7176 ( .A(n2155), .B(n2112), .Z(n2194) );
  CND2X1 U7177 ( .A(n2155), .B(n2112), .Z(n6320) );
  CND2X1 U7178 ( .A(n2158), .B(n2112), .Z(n2196) );
  CND2X1 U7179 ( .A(n2158), .B(n2112), .Z(n6290) );
  CND2X1 U7180 ( .A(n2155), .B(n2130), .Z(n2199) );
  CND2X1 U7181 ( .A(n2155), .B(n2130), .Z(n6260) );
  CND2X1 U7182 ( .A(n2158), .B(n2130), .Z(n2215) );
  CND2X1 U7183 ( .A(n2158), .B(n2130), .Z(n6230) );
  CND2X1 U7184 ( .A(n2155), .B(n2135), .Z(n2217) );
  CND2X1 U7185 ( .A(n2155), .B(n2135), .Z(n6200) );
  CND2X1 U7186 ( .A(n2158), .B(n2135), .Z(n2219) );
  CND2X1 U7187 ( .A(n2158), .B(n2135), .Z(n6170) );
  CIVX2 U7188 ( .A(n21), .Z(n8288) );
  CND2X1 U7189 ( .A(n7173), .B(n7067), .Z(n2055) );
  CND2X1 U7190 ( .A(n7173), .B(n7037), .Z(n2059) );
  CND2X1 U7191 ( .A(n7173), .B(n7007), .Z(n2063) );
  CND2X1 U7192 ( .A(n7173), .B(n6977), .Z(n2066) );
  CND2X1 U7193 ( .A(n7173), .B(n6947), .Z(n2083) );
  CND2X1 U7194 ( .A(n7173), .B(n6917), .Z(n2085) );
  CND2X1 U7195 ( .A(n7173), .B(n6887), .Z(n2088) );
  CND2X1 U7196 ( .A(n7173), .B(n6857), .Z(n2093) );
  CND2X1 U7197 ( .A(n7173), .B(n6827), .Z(n2108) );
  CND2X1 U7198 ( .A(n7173), .B(n6797), .Z(n2110) );
  CND2X1 U7199 ( .A(n7173), .B(n6767), .Z(n2113) );
  CND2X1 U7200 ( .A(n7173), .B(n6737), .Z(n2116) );
  CND2X1 U7201 ( .A(n7173), .B(n6706), .Z(n2131) );
  CND2X1 U7202 ( .A(n7173), .B(n6679), .Z(n2133) );
  CND2X1 U7203 ( .A(n7173), .B(n6652), .Z(n2136) );
  CND2X1 U7204 ( .A(n7173), .B(n6626), .Z(n2140) );
  CND2X1 U7205 ( .A(n7173), .B(n6596), .Z(n2156) );
  CND2X1 U7206 ( .A(n7173), .B(n6566), .Z(n2159) );
  CND2X1 U7207 ( .A(n7173), .B(n6536), .Z(n2161) );
  CND2X1 U7208 ( .A(n7173), .B(n6506), .Z(n2164) );
  CND2X1 U7209 ( .A(n7173), .B(n6476), .Z(n2168) );
  CND2X1 U7210 ( .A(n7173), .B(n6446), .Z(n2171) );
  CND2X1 U7211 ( .A(n7173), .B(n6416), .Z(n2173) );
  CND2X1 U7212 ( .A(n7173), .B(n6386), .Z(n2176) );
  CND2X1 U7213 ( .A(n7173), .B(n6356), .Z(n2191) );
  CND2X1 U7214 ( .A(n7173), .B(n6326), .Z(n2193) );
  CND2X1 U7215 ( .A(n7173), .B(n6296), .Z(n2195) );
  CND2X1 U7216 ( .A(n7173), .B(n6266), .Z(n2198) );
  CND2X1 U7217 ( .A(n7173), .B(n6236), .Z(n2214) );
  CND2X1 U7218 ( .A(n7173), .B(n6206), .Z(n2216) );
  CND2X1 U7219 ( .A(n7173), .B(n6176), .Z(n2218) );
  CIVX2 U7220 ( .A(n69), .Z(n8292) );
  CND2X1 U7221 ( .A(n2130), .B(n2057), .Z(n2132) );
  CND2X1 U7222 ( .A(n2135), .B(n2062), .Z(n2134) );
  CND2X1 U7223 ( .A(n2135), .B(n2057), .Z(n2137) );
  CND2X1 U7224 ( .A(n7173), .B(n7066), .Z(n7068) );
  CND2X1 U7225 ( .A(n7173), .B(n7065), .Z(n7069) );
  CND2X1 U7226 ( .A(n7173), .B(n7036), .Z(n7038) );
  CND2X1 U7227 ( .A(n7173), .B(n7035), .Z(n7039) );
  CND2X1 U7228 ( .A(n7173), .B(n7006), .Z(n7008) );
  CND2X1 U7229 ( .A(n7173), .B(n7005), .Z(n7009) );
  CND2X1 U7230 ( .A(n7173), .B(n6976), .Z(n6978) );
  CND2X1 U7231 ( .A(n7173), .B(n6975), .Z(n6979) );
  CND2X1 U7232 ( .A(n7173), .B(n6946), .Z(n6948) );
  CND2X1 U7233 ( .A(n7173), .B(n6945), .Z(n6949) );
  CND2X1 U7234 ( .A(n7173), .B(n6916), .Z(n6918) );
  CND2X1 U7235 ( .A(n7173), .B(n6915), .Z(n6919) );
  CND2X1 U7236 ( .A(n7173), .B(n6886), .Z(n6888) );
  CND2X1 U7237 ( .A(n7173), .B(n6885), .Z(n6889) );
  CND2X1 U7238 ( .A(n7173), .B(n6856), .Z(n6858) );
  CND2X1 U7239 ( .A(n7173), .B(n6855), .Z(n6859) );
  CND2X1 U7240 ( .A(n7173), .B(n6826), .Z(n6828) );
  CND2X1 U7241 ( .A(n7173), .B(n6825), .Z(n6829) );
  CND2X1 U7242 ( .A(n7173), .B(n6796), .Z(n6798) );
  CND2X1 U7243 ( .A(n7173), .B(n6795), .Z(n6799) );
  CND2X1 U7244 ( .A(n7173), .B(n6766), .Z(n6768) );
  CND2X1 U7245 ( .A(n7173), .B(n6765), .Z(n6769) );
  CND2X1 U7246 ( .A(n7173), .B(n6736), .Z(n6738) );
  CND2X1 U7247 ( .A(n7173), .B(n6735), .Z(n6739) );
  CND2X1 U7248 ( .A(n7173), .B(n6705), .Z(n6708) );
  CND2X1 U7249 ( .A(n7173), .B(n6704), .Z(n6709) );
  CND2X1 U7250 ( .A(n7173), .B(n6678), .Z(n6681) );
  CND2X1 U7251 ( .A(n7173), .B(n6677), .Z(n6682) );
  CND2X1 U7252 ( .A(n7173), .B(n6651), .Z(n6654) );
  CND2X1 U7253 ( .A(n7173), .B(n6650), .Z(n6655) );
  CND2X1 U7254 ( .A(n7173), .B(n6625), .Z(n6627) );
  CND2X1 U7255 ( .A(n7173), .B(n6624), .Z(n6628) );
  CND2X1 U7256 ( .A(n7173), .B(n6595), .Z(n6597) );
  CND2X1 U7257 ( .A(n7173), .B(n6594), .Z(n6598) );
  CND2X1 U7258 ( .A(n7173), .B(n6565), .Z(n6567) );
  CND2X1 U7259 ( .A(n7173), .B(n6564), .Z(n6568) );
  CND2X1 U7260 ( .A(n7173), .B(n6535), .Z(n6537) );
  CND2X1 U7261 ( .A(n7173), .B(n6534), .Z(n6538) );
  CND2X1 U7262 ( .A(n7173), .B(n6505), .Z(n6507) );
  CND2X1 U7263 ( .A(n7173), .B(n6504), .Z(n6508) );
  CND2X1 U7264 ( .A(n7173), .B(n6475), .Z(n6477) );
  CND2X1 U7265 ( .A(n7173), .B(n6474), .Z(n6478) );
  CND2X1 U7266 ( .A(n7173), .B(n6445), .Z(n6447) );
  CND2X1 U7267 ( .A(n7173), .B(n6444), .Z(n6448) );
  CND2X1 U7268 ( .A(n7173), .B(n6415), .Z(n6417) );
  CND2X1 U7269 ( .A(n7173), .B(n6414), .Z(n6418) );
  CND2X1 U7270 ( .A(n7173), .B(n6385), .Z(n6387) );
  CND2X1 U7271 ( .A(n7173), .B(n6384), .Z(n6388) );
  CND2X1 U7272 ( .A(n7173), .B(n6355), .Z(n6357) );
  CND2X1 U7273 ( .A(n7173), .B(n6354), .Z(n6358) );
  CND2X1 U7274 ( .A(n7173), .B(n6325), .Z(n6327) );
  CND2X1 U7275 ( .A(n7173), .B(n6324), .Z(n6328) );
  CND2X1 U7276 ( .A(n7173), .B(n6295), .Z(n6297) );
  CND2X1 U7277 ( .A(n7173), .B(n6294), .Z(n6298) );
  CND2X1 U7278 ( .A(n7173), .B(n6265), .Z(n6267) );
  CND2X1 U7279 ( .A(n7173), .B(n6264), .Z(n6268) );
  CND2X1 U7280 ( .A(n7173), .B(n6235), .Z(n6237) );
  CND2X1 U7281 ( .A(n7173), .B(n6234), .Z(n6238) );
  CND2X1 U7282 ( .A(n7173), .B(n6205), .Z(n6207) );
  CND2X1 U7283 ( .A(n7173), .B(n6204), .Z(n6208) );
  CND2X1 U7284 ( .A(n7173), .B(n6175), .Z(n6177) );
  CND2X1 U7285 ( .A(n7173), .B(n6174), .Z(n6178) );
  CIVX2 U7286 ( .A(n16), .Z(n8289) );
  CND2X1 U7287 ( .A(n7171), .B(n6162), .Z(n286) );
  CANR2X1 U7288 ( .A(n7258), .B(rd_ptr[3]), .C(n1202), .D(n8293), .Z(n1200) );
  COND2X1 U7289 ( .A(n7270), .B(n8296), .C(rd_ptr[4]), .D(n1204), .Z(n1202) );
  CND2X1 U7290 ( .A(rd_ptr[6]), .B(n8302), .Z(n35) );
  COND1XL U7291 ( .A(rd_ptr[1]), .B(n352), .C(n354), .Z(n349) );
  COND1XL U7292 ( .A(n61), .B(n62), .C(n8288), .Z(n57) );
  CND2X1 U7293 ( .A(n8289), .B(n60), .Z(n58) );
  CND2X1 U7294 ( .A(rd_ptr[5]), .B(n8308), .Z(n93) );
  COND2X1 U7295 ( .A(n64), .B(n8296), .C(rd_ptr[4]), .D(n1500), .Z(n269) );
  CANR3X1 U7296 ( .A(rd_ptr[5]), .B(n89), .C(n1501), .D(n1502), .Z(n1500) );
  COND3X1 U7297 ( .A(n8299), .B(n8271), .C(n1518), .D(n1519), .Z(n1501) );
  COND1XL U7298 ( .A(rd_ptr[1]), .B(n245), .C(n246), .Z(n243) );
  COND1X1 U7299 ( .A(n7250), .B(n8293), .C(n1801), .Z(n266) );
  CANR2X1 U7300 ( .A(n8292), .B(n230), .C(n8291), .D(n1802), .Z(n1801) );
  CND4X1 U7301 ( .A(n1803), .B(n1804), .C(n1805), .D(n1806), .Z(n1802) );
  CANR2X1 U7302 ( .A(n380), .B(n235), .C(n2453), .D(n7094), .Z(n1806) );
  CANR2X1 U7303 ( .A(n380), .B(n339), .C(n3136), .D(n7094), .Z(n379) );
  COND2X1 U7304 ( .A(n697), .B(n8308), .C(rd_ptr[6]), .D(n699), .Z(n127) );
  CNR4X1 U7305 ( .A(n700), .B(n701), .C(n702), .D(n703), .Z(n699) );
  CNR4X1 U7306 ( .A(n712), .B(n713), .C(n714), .D(n715), .Z(n697) );
  COND1X1 U7307 ( .A(rd_ptr[3]), .B(n7250), .C(n228), .Z(n105) );
  CANR2X1 U7308 ( .A(n8294), .B(n229), .C(n8295), .D(n230), .Z(n228) );
  CND4X1 U7309 ( .A(n231), .B(n232), .C(n233), .D(n234), .Z(n229) );
  COND1XL U7310 ( .A(rd_ptr[1]), .B(n330), .C(n331), .Z(n311) );
  CANR3X1 U7311 ( .A(buffer[396]), .B(n4241), .C(n78), .D(n79), .Z(n75) );
  CANR2X1 U7312 ( .A(n8295), .B(n185), .C(n8294), .D(n184), .Z(n356) );
  CANR2X1 U7313 ( .A(n7171), .B(n7208), .C(dataout_stg_1[5]), .D(n7092), .Z(
        n260) );
  COND2X1 U7314 ( .A(rd_ptr[2]), .B(n266), .C(n8290), .D(n198), .Z(n267) );
  COND2X1 U7315 ( .A(n1523), .B(n8308), .C(rd_ptr[6]), .D(n1524), .Z(n89) );
  CNR4X1 U7316 ( .A(n1525), .B(n1526), .C(n1527), .D(n1528), .Z(n1524) );
  CNR4X1 U7317 ( .A(n1537), .B(n1538), .C(n1539), .D(n1540), .Z(n1523) );
  COND2X1 U7318 ( .A(n7142), .B(n7727), .C(n7139), .D(n7471), .Z(n1528) );
  CANR2X1 U7319 ( .A(n289), .B(rd_ptr[2]), .C(n8290), .D(n588), .Z(n330) );
  COND2X1 U7320 ( .A(n7265), .B(n69), .C(n590), .D(n67), .Z(n589) );
  CND2X1 U7321 ( .A(rd_ptr[6]), .B(rd_ptr[5]), .Z(n76) );
  COND2X1 U7322 ( .A(n7249), .B(n8290), .C(rd_ptr[2]), .D(n1198), .Z(n352) );
  CANR2X1 U7323 ( .A(n2864), .B(n7097), .C(n2867), .D(n8304), .Z(n897) );
  CANR2X1 U7324 ( .A(n2401), .B(n7097), .C(n2404), .D(n8304), .Z(n1909) );
  CANR1X1 U7325 ( .A(n269), .B(rd_ptr[3]), .C(n1401), .Z(n314) );
  CND4X1 U7326 ( .A(n1403), .B(n1404), .C(n1405), .D(n1406), .Z(n1402) );
  CANR2X1 U7327 ( .A(n380), .B(n276), .C(n2624), .D(n7094), .Z(n1406) );
  CANR2X1 U7328 ( .A(n380), .B(n254), .C(n3030), .D(n7094), .Z(n1003) );
  CANR2X1 U7329 ( .A(n380), .B(n323), .C(n2567), .D(n7094), .Z(n1609) );
  CANR3X1 U7330 ( .A(n3162), .B(n7097), .C(n71), .D(n72), .Z(n70) );
  CANR2X1 U7331 ( .A(buffer[1030]), .B(n8304), .C(buffer[774]), .D(n8305), .Z(
        n233) );
  CANR2X1 U7332 ( .A(buffer[1032]), .B(n8304), .C(buffer[776]), .D(n8305), .Z(
        n190) );
  CANR2X1 U7333 ( .A(buffer[1031]), .B(n8304), .C(buffer[775]), .D(n8305), .Z(
        n214) );
  COND2X1 U7334 ( .A(n3170), .B(n92), .C(n3169), .D(n120), .Z(n118) );
  CANR2X1 U7335 ( .A(buffer[1033]), .B(n8304), .C(buffer[777]), .D(n8305), .Z(
        n168) );
  CND2X1 U7336 ( .A(n146), .B(n147), .Z(n139) );
  CANR2X1 U7337 ( .A(buffer[1034]), .B(n8304), .C(buffer[778]), .D(n8305), .Z(
        n146) );
  CANR2X1 U7338 ( .A(buffer[518]), .B(n7096), .C(n8306), .D(n236), .Z(n1804)
         );
  CANR2X1 U7339 ( .A(n7096), .B(buffer[519]), .C(n8306), .D(n217), .Z(n793) );
  CANR2X1 U7340 ( .A(n7096), .B(buffer[521]), .C(n8301), .D(n166), .Z(n490) );
  CANR2X1 U7341 ( .A(buffer[520]), .B(n7096), .C(n8301), .D(n193), .Z(n1304)
         );
  CANR2X1 U7342 ( .A(n7096), .B(buffer[525]), .C(n8301), .D(n36), .Z(n1152) );
  CANR2X1 U7343 ( .A(n7096), .B(buffer[517]), .C(n8306), .D(n255), .Z(n1001)
         );
  CANR2X1 U7344 ( .A(buffer[522]), .B(n7096), .C(n8301), .D(n144), .Z(n1758)
         );
  COND1XL U7345 ( .A(rd_ptr[1]), .B(n267), .C(n264), .Z(n262) );
  CANR2X1 U7346 ( .A(buffer[1037]), .B(n8304), .C(buffer[781]), .D(n8305), .Z(
        n26) );
  COND11X1 U7347 ( .A(n10), .B(n50), .C(n7217), .D(n52), .Z(n3176) );
  CND2X1 U7348 ( .A(n4264), .B(n7091), .Z(n52) );
  CANR2X1 U7349 ( .A(n7172), .B(n54), .C(n7171), .D(n49), .Z(n50) );
  CANR2X1 U7350 ( .A(n8292), .B(n211), .C(n8291), .D(n791), .Z(n790) );
  CND4X1 U7351 ( .A(n792), .B(n793), .C(n794), .D(n795), .Z(n791) );
  CANR2X1 U7352 ( .A(n380), .B(n216), .C(n2916), .D(n7094), .Z(n795) );
  CND4X1 U7353 ( .A(n1303), .B(n1304), .C(n1305), .D(n1306), .Z(n1302) );
  CANR3X1 U7354 ( .A(n2292), .B(n7094), .C(rd_ptr[4]), .D(n1307), .Z(n1306) );
  CANR2X1 U7355 ( .A(buffer[264]), .B(n8297), .C(buffer[776]), .D(n7095), .Z(
        n1305) );
  COND2X1 U7356 ( .A(n8283), .B(n7111), .C(n6166), .D(n7206), .Z(n3200) );
  COND2X1 U7357 ( .A(n8282), .B(n7111), .C(n6167), .D(n7205), .Z(n3201) );
  COND2X1 U7358 ( .A(n8281), .B(n7111), .C(n6166), .D(n7204), .Z(n3202) );
  COND2X1 U7359 ( .A(n8280), .B(n7111), .C(n6166), .D(n7203), .Z(n3203) );
  COND2X1 U7360 ( .A(n8279), .B(n7111), .C(n6168), .D(n7202), .Z(n3204) );
  COND2X1 U7361 ( .A(n8278), .B(n7111), .C(n6169), .D(n7201), .Z(n3205) );
  COND2X1 U7362 ( .A(n8277), .B(n7111), .C(n6167), .D(n7200), .Z(n3206) );
  CANR2X1 U7363 ( .A(n8298), .B(n938), .C(n2844), .D(n7094), .Z(n902) );
  CND2X1 U7364 ( .A(n2848), .B(n4242), .Z(n940) );
  CANR2X1 U7365 ( .A(n8298), .B(n1949), .C(n2381), .D(n7094), .Z(n1913) );
  CANR2X1 U7366 ( .A(n380), .B(n297), .C(n2755), .D(n7094), .Z(n594) );
  CANR2X1 U7367 ( .A(buffer[1028]), .B(n8304), .C(buffer[772]), .D(n8305), .Z(
        n274) );
  CND4X1 U7368 ( .A(n7281), .B(n490), .C(n491), .D(n492), .Z(n488) );
  CANR3X1 U7369 ( .A(n3047), .B(n7094), .C(rd_ptr[4]), .D(n493), .Z(n492) );
  CANR2X1 U7370 ( .A(n7171), .B(n369), .C(dataout_stg_1[0]), .D(n4), .Z(n368)
         );
  COND1XL U7371 ( .A(n7246), .B(n99), .C(n348), .Z(n369) );
  COND1XL U7372 ( .A(n6161), .B(n310), .C(n8284), .Z(n365) );
  COND3X1 U7373 ( .A(n1195), .B(n1196), .C(n6160), .D(n7172), .Z(n367) );
  CND3XL U7374 ( .A(n310), .B(n311), .C(n7172), .Z(n303) );
  CANR2X1 U7375 ( .A(n7171), .B(n301), .C(dataout_stg_1[3]), .D(n7091), .Z(
        n304) );
  CND3XL U7376 ( .A(n6160), .B(n4243), .C(n7170), .Z(n281) );
  CANR2X1 U7377 ( .A(n7171), .B(n7213), .C(dataout_stg_1[4]), .D(n4), .Z(n282)
         );
  CND4X1 U7378 ( .A(n357), .B(n358), .C(n359), .D(n360), .Z(n184) );
  CANR2X1 U7379 ( .A(buffer[1024]), .B(n8304), .C(buffer[768]), .D(n8305), .Z(
        n359) );
  CANR2X1 U7380 ( .A(n8303), .B(n363), .C(n8298), .D(n364), .Z(n357) );
  CND4X1 U7381 ( .A(n7279), .B(n1758), .C(n1759), .D(n1760), .Z(n318) );
  CANR2X1 U7382 ( .A(n380), .B(n145), .C(n2502), .D(n7094), .Z(n1760) );
  CND4X1 U7383 ( .A(n7274), .B(n1152), .C(n1153), .D(n1154), .Z(n249) );
  CANR2X1 U7384 ( .A(n380), .B(n38), .C(n2965), .D(n7094), .Z(n1154) );
  CND4X1 U7385 ( .A(n250), .B(n251), .C(n252), .D(n253), .Z(n23) );
  CANR2X1 U7386 ( .A(buffer[1029]), .B(n8304), .C(buffer[773]), .D(n8305), .Z(
        n252) );
  CND4X1 U7387 ( .A(n319), .B(n320), .C(n321), .D(n322), .Z(n148) );
  CANR2X1 U7388 ( .A(buffer[1026]), .B(n8304), .C(buffer[770]), .D(n8305), .Z(
        n321) );
  CANR2X1 U7389 ( .A(n8303), .B(n325), .C(n8298), .D(n326), .Z(n319) );
  COND1XL U7390 ( .A(rd_ptr[5]), .B(n7277), .C(n124), .Z(n116) );
  COND3X1 U7391 ( .A(n7215), .B(n8), .C(n328), .D(n329), .Z(n3187) );
  CND2X1 U7392 ( .A(n4287), .B(n7091), .Z(n329) );
  COND3X1 U7393 ( .A(n7218), .B(n310), .C(n311), .D(n7171), .Z(n328) );
  CND3XL U7394 ( .A(n7218), .B(n243), .C(n7170), .Z(n240) );
  CANR2X1 U7395 ( .A(n7212), .B(n7171), .C(dataout_stg_1[6]), .D(n7091), .Z(
        n241) );
  CND2X1 U7396 ( .A(n4262), .B(n4), .Z(n223) );
  CND3XL U7397 ( .A(n6163), .B(n202), .C(n7171), .Z(n222) );
  CND2X1 U7398 ( .A(n4263), .B(n7092), .Z(n151) );
  CND3XL U7399 ( .A(n152), .B(n131), .C(n7171), .Z(n150) );
  CANR2X1 U7400 ( .A(n8294), .B(n210), .C(n8295), .D(n211), .Z(n209) );
  CND4X1 U7401 ( .A(n212), .B(n213), .C(n214), .D(n215), .Z(n210) );
  CAN4X1 U7402 ( .A(n335), .B(n336), .C(n337), .D(n338), .Z(n156) );
  CANR2X1 U7403 ( .A(n8301), .B(n341), .C(n8298), .D(n342), .Z(n335) );
  CANR2X1 U7404 ( .A(n380), .B(n361), .C(n2235), .D(n7094), .Z(n1208) );
  CANR2X1 U7405 ( .A(buffer[1027]), .B(n8304), .C(buffer[771]), .D(n8305), .Z(
        n295) );
  CANR2X1 U7406 ( .A(n380), .B(n125), .C(n2714), .D(n7094), .Z(n692) );
  CNIVX1 U7407 ( .A(reqlen[0]), .Z(n6160) );
  CNIVX1 U7408 ( .A(reqlen[2]), .Z(n6162) );
  CNIVX1 U7409 ( .A(reqlen[1]), .Z(n6161) );
  COND11X1 U7410 ( .A(n97), .B(n7227), .C(n99), .D(n100), .Z(n96) );
  COND4CX1 U7411 ( .A(n6160), .B(n101), .C(n102), .D(n7172), .Z(n100) );
  COND3X1 U7412 ( .A(n11), .B(n12), .C(n6164), .D(rd_ptr[0]), .Z(n9) );
  CANR11X1 U7413 ( .A(n7172), .B(n202), .C(n203), .D(n204), .Z(n201) );
  COND4CX1 U7414 ( .A(n174), .B(n175), .C(n7207), .D(n7171), .Z(n173) );
  CND2X1 U7415 ( .A(rd_ptr[5]), .B(n127), .Z(n690) );
  CANR2X1 U7416 ( .A(n6161), .B(n346), .C(n7209), .D(n7172), .Z(n345) );
  CND2X1 U7417 ( .A(rd_ptr[4]), .B(n8293), .Z(n69) );
  CNR2X1 U7418 ( .A(n6164), .B(rst), .Z(n7092) );
  CNR2X1 U7419 ( .A(n6165), .B(rst), .Z(n7091) );
  CND2X1 U7420 ( .A(rd_ptr[4]), .B(rd_ptr[3]), .Z(n29) );
  CND2X1 U7421 ( .A(rd_ptr[1]), .B(n8290), .Z(n16) );
  CND2X1 U7422 ( .A(rd_ptr[3]), .B(n8296), .Z(n65) );
  CND2X1 U7423 ( .A(rd_ptr[2]), .B(rd_ptr[1]), .Z(n21) );
  CND2X1 U7424 ( .A(rd_ptr[2]), .B(n8287), .Z(n19) );
  CND2X1 U7425 ( .A(rd_ptr[0]), .B(n6164), .Z(n97) );
  CAN2X1 U7426 ( .A(reqin), .B(n7173), .Z(n6164) );
  COND2X1 U7427 ( .A(n8276), .B(n7110), .C(n6167), .D(n7199), .Z(n3207) );
  COND2X1 U7428 ( .A(n8275), .B(n7110), .C(n6166), .D(n7198), .Z(n3208) );
  COND2X1 U7429 ( .A(n8274), .B(n7110), .C(n6167), .D(n7197), .Z(n3209) );
  COND2X1 U7430 ( .A(n8273), .B(n7110), .C(n6168), .D(n7196), .Z(n3210) );
  COND2X1 U7431 ( .A(n8272), .B(n7110), .C(n6168), .D(n7195), .Z(n3211) );
  COND2X1 U7432 ( .A(n8270), .B(n7110), .C(n6169), .D(n7193), .Z(n3213) );
  COND2X1 U7433 ( .A(n8269), .B(n7110), .C(n6169), .D(n7192), .Z(n3214) );
  COND2X1 U7434 ( .A(n8268), .B(n7110), .C(n6169), .D(n7191), .Z(n3215) );
  COND2X1 U7435 ( .A(n8141), .B(n6992), .C(n7192), .D(n6972), .Z(n3342) );
  COND2X1 U7436 ( .A(n8140), .B(n6993), .C(n7191), .D(n6973), .Z(n3343) );
  COND2X1 U7437 ( .A(n8045), .B(n6902), .C(n7192), .D(n6882), .Z(n3438) );
  COND2X1 U7438 ( .A(n8044), .B(n6903), .C(n7191), .D(n6883), .Z(n3439) );
  COND2X1 U7439 ( .A(n3172), .B(n6873), .C(n7195), .D(n6853), .Z(n3467) );
  COND2X1 U7440 ( .A(n8015), .B(n6875), .C(n7194), .D(n6856), .Z(n3468) );
  COND2X1 U7441 ( .A(n3171), .B(n6642), .C(n7195), .D(n6622), .Z(n3723) );
  COND2X1 U7442 ( .A(n7757), .B(n6641), .C(n7192), .D(n6621), .Z(n3726) );
  COND2X1 U7443 ( .A(n7756), .B(n6642), .C(n7191), .D(n6622), .Z(n3727) );
  COND2X1 U7444 ( .A(n7629), .B(n6521), .C(n7192), .D(n6501), .Z(n3854) );
  COND2X1 U7445 ( .A(n7628), .B(n6522), .C(n7191), .D(n6502), .Z(n3855) );
  COND2X1 U7446 ( .A(n3170), .B(n6402), .C(n7195), .D(n6382), .Z(n3979) );
  COND2X1 U7447 ( .A(n7501), .B(n6401), .C(n7192), .D(n6381), .Z(n3982) );
  COND2X1 U7448 ( .A(n7500), .B(n6402), .C(n7191), .D(n6382), .Z(n3983) );
  COND2X1 U7449 ( .A(n7373), .B(n6281), .C(n7192), .D(n6261), .Z(n4110) );
  COND2X1 U7450 ( .A(n7372), .B(n6282), .C(n7191), .D(n6262), .Z(n4111) );
  COND2X1 U7451 ( .A(n7273), .B(n6191), .C(n7192), .D(n6171), .Z(n4206) );
  COND2X1 U7452 ( .A(n7272), .B(n6192), .C(n7191), .D(n6172), .Z(n4207) );
  COND2X1 U7453 ( .A(n3169), .B(n7108), .C(n6168), .D(n7195), .Z(n4235) );
  COND2X1 U7454 ( .A(n8155), .B(n6981), .C(n7206), .D(n6972), .Z(n3328) );
  COND2X1 U7455 ( .A(n8154), .B(n6982), .C(n7205), .D(n6973), .Z(n3329) );
  COND2X1 U7456 ( .A(n8153), .B(n6983), .C(n7204), .D(n6972), .Z(n3330) );
  COND2X1 U7457 ( .A(n8152), .B(n6984), .C(n7203), .D(n6973), .Z(n3331) );
  COND2X1 U7458 ( .A(n8151), .B(n6985), .C(n7202), .D(n6974), .Z(n3332) );
  COND2X1 U7459 ( .A(n8150), .B(n6986), .C(n7201), .D(n6972), .Z(n3333) );
  COND2X1 U7460 ( .A(n8149), .B(n6988), .C(n7200), .D(n6974), .Z(n3334) );
  COND2X1 U7461 ( .A(n8148), .B(n6989), .C(n7199), .D(n6975), .Z(n3335) );
  COND2X1 U7462 ( .A(n8147), .B(n6990), .C(n7198), .D(n6975), .Z(n3336) );
  COND2X1 U7463 ( .A(n8146), .B(n6991), .C(n7197), .D(n6976), .Z(n3337) );
  COND2X1 U7464 ( .A(n8145), .B(n6992), .C(n7196), .D(n6977), .Z(n3338) );
  COND2X1 U7465 ( .A(n8144), .B(n6993), .C(n7195), .D(n6973), .Z(n3339) );
  COND2X1 U7466 ( .A(n8142), .B(n6996), .C(n7193), .D(n6977), .Z(n3341) );
  COND2X1 U7467 ( .A(n8027), .B(n6861), .C(n7206), .D(n6852), .Z(n3456) );
  COND2X1 U7468 ( .A(n8026), .B(n6862), .C(n7205), .D(n6853), .Z(n3457) );
  COND2X1 U7469 ( .A(n8025), .B(n6863), .C(n7204), .D(n6852), .Z(n3458) );
  COND2X1 U7470 ( .A(n8024), .B(n6864), .C(n7203), .D(n6853), .Z(n3459) );
  COND2X1 U7471 ( .A(n8023), .B(n6865), .C(n7202), .D(n6854), .Z(n3460) );
  COND2X1 U7472 ( .A(n8022), .B(n6866), .C(n7201), .D(n6852), .Z(n3461) );
  COND2X1 U7473 ( .A(n8021), .B(n6868), .C(n7200), .D(n6854), .Z(n3462) );
  COND2X1 U7474 ( .A(n8020), .B(n6869), .C(n7199), .D(n6855), .Z(n3463) );
  COND2X1 U7475 ( .A(n8019), .B(n6870), .C(n7198), .D(n6855), .Z(n3464) );
  COND2X1 U7476 ( .A(n8018), .B(n6871), .C(n7197), .D(n6856), .Z(n3465) );
  COND2X1 U7477 ( .A(n8017), .B(n6872), .C(n7196), .D(n6857), .Z(n3466) );
  COND2X1 U7478 ( .A(n8014), .B(n6876), .C(n7193), .D(n6857), .Z(n3469) );
  COND2X1 U7479 ( .A(n7899), .B(n6741), .C(n7206), .D(n6732), .Z(n3584) );
  COND2X1 U7480 ( .A(n7898), .B(n6742), .C(n7205), .D(n6733), .Z(n3585) );
  COND2X1 U7481 ( .A(n7897), .B(n6743), .C(n7204), .D(n6732), .Z(n3586) );
  COND2X1 U7482 ( .A(n7896), .B(n6744), .C(n7203), .D(n6733), .Z(n3587) );
  COND2X1 U7483 ( .A(n7895), .B(n6745), .C(n7202), .D(n6734), .Z(n3588) );
  COND2X1 U7484 ( .A(n7894), .B(n6746), .C(n7201), .D(n6732), .Z(n3589) );
  COND2X1 U7485 ( .A(n7893), .B(n6748), .C(n7200), .D(n6734), .Z(n3590) );
  COND2X1 U7486 ( .A(n7892), .B(n6749), .C(n7199), .D(n6735), .Z(n3591) );
  COND2X1 U7487 ( .A(n7891), .B(n6750), .C(n7198), .D(n6735), .Z(n3592) );
  COND2X1 U7488 ( .A(n7890), .B(n6751), .C(n7197), .D(n6736), .Z(n3593) );
  COND2X1 U7489 ( .A(n7889), .B(n6752), .C(n7196), .D(n6737), .Z(n3594) );
  COND2X1 U7490 ( .A(n7888), .B(n6753), .C(n7195), .D(n6733), .Z(n3595) );
  COND2X1 U7491 ( .A(n7886), .B(n6756), .C(n7193), .D(n6737), .Z(n3597) );
  COND2X1 U7492 ( .A(n7771), .B(n6630), .C(n7206), .D(n6621), .Z(n3712) );
  COND2X1 U7493 ( .A(n7770), .B(n6631), .C(n7205), .D(n6622), .Z(n3713) );
  COND2X1 U7494 ( .A(n7769), .B(n6632), .C(n7204), .D(n6621), .Z(n3714) );
  COND2X1 U7495 ( .A(n7768), .B(n6633), .C(n7203), .D(n6622), .Z(n3715) );
  COND2X1 U7496 ( .A(n7767), .B(n6634), .C(n7202), .D(n6623), .Z(n3716) );
  COND2X1 U7497 ( .A(n7766), .B(n6635), .C(n7201), .D(n6621), .Z(n3717) );
  COND2X1 U7498 ( .A(n7765), .B(n6637), .C(n7200), .D(n6623), .Z(n3718) );
  COND2X1 U7499 ( .A(n7764), .B(n6638), .C(n7199), .D(n6624), .Z(n3719) );
  COND2X1 U7500 ( .A(n7763), .B(n6639), .C(n7198), .D(n6624), .Z(n3720) );
  COND2X1 U7501 ( .A(n7762), .B(n6640), .C(n7197), .D(n6625), .Z(n3721) );
  COND2X1 U7502 ( .A(n7761), .B(n6641), .C(n7196), .D(n6626), .Z(n3722) );
  COND2X1 U7503 ( .A(n7758), .B(n6645), .C(n7193), .D(n6626), .Z(n3725) );
  COND2X1 U7504 ( .A(n7515), .B(n6390), .C(n7206), .D(n6381), .Z(n3968) );
  COND2X1 U7505 ( .A(n7514), .B(n6391), .C(n7205), .D(n6382), .Z(n3969) );
  COND2X1 U7506 ( .A(n7513), .B(n6392), .C(n7204), .D(n6381), .Z(n3970) );
  COND2X1 U7507 ( .A(n7512), .B(n6393), .C(n7203), .D(n6382), .Z(n3971) );
  COND2X1 U7508 ( .A(n7511), .B(n6394), .C(n7202), .D(n6383), .Z(n3972) );
  COND2X1 U7509 ( .A(n7510), .B(n6395), .C(n7201), .D(n6381), .Z(n3973) );
  COND2X1 U7510 ( .A(n7509), .B(n6397), .C(n7200), .D(n6383), .Z(n3974) );
  COND2X1 U7511 ( .A(n7508), .B(n6398), .C(n7199), .D(n6384), .Z(n3975) );
  COND2X1 U7512 ( .A(n7507), .B(n6399), .C(n7198), .D(n6384), .Z(n3976) );
  COND2X1 U7513 ( .A(n7506), .B(n6400), .C(n7197), .D(n6385), .Z(n3977) );
  COND2X1 U7514 ( .A(n7505), .B(n6401), .C(n7196), .D(n6386), .Z(n3978) );
  COND2X1 U7515 ( .A(n7502), .B(n6405), .C(n7193), .D(n6386), .Z(n3981) );
  COND2X1 U7516 ( .A(n7387), .B(n6270), .C(n7206), .D(n6261), .Z(n4096) );
  COND2X1 U7517 ( .A(n7386), .B(n6271), .C(n7205), .D(n6262), .Z(n4097) );
  COND2X1 U7518 ( .A(n7385), .B(n6272), .C(n7204), .D(n6261), .Z(n4098) );
  COND2X1 U7519 ( .A(n7384), .B(n6273), .C(n7203), .D(n6262), .Z(n4099) );
  COND2X1 U7520 ( .A(n7383), .B(n6274), .C(n7202), .D(n6263), .Z(n4100) );
  COND2X1 U7521 ( .A(n7382), .B(n6275), .C(n7201), .D(n6261), .Z(n4101) );
  COND2X1 U7522 ( .A(n7381), .B(n6277), .C(n7200), .D(n6263), .Z(n4102) );
  COND2X1 U7523 ( .A(n7380), .B(n6278), .C(n7199), .D(n6264), .Z(n4103) );
  COND2X1 U7524 ( .A(n7379), .B(n6279), .C(n7198), .D(n6264), .Z(n4104) );
  COND2X1 U7525 ( .A(n7378), .B(n6280), .C(n7197), .D(n6265), .Z(n4105) );
  COND2X1 U7526 ( .A(n7377), .B(n6281), .C(n7196), .D(n6266), .Z(n4106) );
  COND2X1 U7527 ( .A(n7376), .B(n6282), .C(n7195), .D(n6262), .Z(n4107) );
  COND2X1 U7528 ( .A(n7374), .B(n6285), .C(n7193), .D(n6266), .Z(n4109) );
  COND2X1 U7529 ( .A(n7243), .B(n7109), .C(n6166), .D(n7206), .Z(n4224) );
  COND2X1 U7530 ( .A(n7242), .B(n7108), .C(n6167), .D(n7205), .Z(n4225) );
  COND2X1 U7531 ( .A(n7239), .B(n7108), .C(n6166), .D(n7204), .Z(n4226) );
  COND2X1 U7532 ( .A(n7238), .B(n7108), .C(n6166), .D(n7203), .Z(n4227) );
  COND2X1 U7533 ( .A(n7236), .B(n7108), .C(n6168), .D(n7202), .Z(n4228) );
  COND2X1 U7534 ( .A(n7235), .B(n7108), .C(n6169), .D(n7201), .Z(n4229) );
  COND2X1 U7535 ( .A(n7234), .B(n7108), .C(n6167), .D(n7200), .Z(n4230) );
  COND2X1 U7536 ( .A(n7232), .B(n7108), .C(n6167), .D(n7199), .Z(n4231) );
  COND2X1 U7537 ( .A(n7231), .B(n7108), .C(n6166), .D(n7198), .Z(n4232) );
  COND2X1 U7538 ( .A(n7229), .B(n7108), .C(n6167), .D(n7197), .Z(n4233) );
  COND2X1 U7539 ( .A(n7228), .B(n7108), .C(n6168), .D(n7196), .Z(n4234) );
  COND2X1 U7540 ( .A(n7223), .B(n7108), .C(n6169), .D(n7193), .Z(n4237) );
  CAN2X1 U7541 ( .A(reqin), .B(n7173), .Z(n6165) );
  CIVX2 U7542 ( .A(rd_ptr[4]), .Z(n8296) );
  CNIVX1 U7543 ( .A(reqlen[3]), .Z(n6163) );
  CNR2X1 U7544 ( .A(n3173), .B(rst), .Z(n4) );
  CIVX2 U7545 ( .A(datain[0]), .Z(n7206) );
  CIVX2 U7546 ( .A(datain[1]), .Z(n7205) );
  CIVX2 U7547 ( .A(datain[2]), .Z(n7204) );
  CIVX2 U7548 ( .A(datain[3]), .Z(n7203) );
  CIVX2 U7549 ( .A(datain[4]), .Z(n7202) );
  CIVX2 U7550 ( .A(datain[5]), .Z(n7201) );
  CIVX2 U7551 ( .A(datain[6]), .Z(n7200) );
  CIVX2 U7552 ( .A(datain[7]), .Z(n7199) );
  CIVX2 U7553 ( .A(datain[8]), .Z(n7198) );
  CIVX2 U7554 ( .A(datain[9]), .Z(n7197) );
  CIVX2 U7555 ( .A(datain[10]), .Z(n7196) );
  CIVX2 U7556 ( .A(datain[11]), .Z(n7195) );
  CIVX2 U7557 ( .A(datain[12]), .Z(n7194) );
  CIVX2 U7558 ( .A(datain[13]), .Z(n7193) );
  CIVX2 U7559 ( .A(datain[14]), .Z(n7192) );
  CIVX2 U7560 ( .A(datain[15]), .Z(n7191) );
  CIVX2 U7561 ( .A(datain[16]), .Z(n7190) );
  CIVX2 U7562 ( .A(datain[17]), .Z(n7189) );
  CIVX2 U7563 ( .A(datain[18]), .Z(n7188) );
  CIVX2 U7564 ( .A(datain[19]), .Z(n7187) );
  CIVX2 U7565 ( .A(datain[20]), .Z(n7186) );
  CIVX2 U7566 ( .A(datain[21]), .Z(n7185) );
  CIVX2 U7567 ( .A(datain[22]), .Z(n7184) );
  CIVX2 U7568 ( .A(datain[23]), .Z(n7183) );
  CIVX2 U7569 ( .A(datain[24]), .Z(n7182) );
  CIVX2 U7570 ( .A(datain[25]), .Z(n7181) );
  CIVX2 U7571 ( .A(datain[26]), .Z(n7180) );
  CIVX2 U7572 ( .A(datain[27]), .Z(n7179) );
  CIVX2 U7573 ( .A(datain[28]), .Z(n7178) );
  CIVX2 U7574 ( .A(datain[29]), .Z(n7177) );
  CIVX2 U7575 ( .A(datain[30]), .Z(n7176) );
  CIVX2 U7576 ( .A(datain[31]), .Z(n7175) );
  CNR2X1 U7577 ( .A(reqin), .B(rst), .Z(n2234) );
  CAN2X1 U7578 ( .A(reqin), .B(n7173), .Z(n3173) );
  CANR4CX1 U7579 ( .A(n7224), .B(n8), .C(n9), .D(n10), .Z(n5) );
  COND3X1 U7580 ( .A(rd_ptr[1]), .B(n56), .C(n57), .D(n58), .Z(n49) );
  CANR4CX1 U7581 ( .A(n8287), .B(n56), .C(n104), .D(n7217), .Z(n102) );
  CND2X1 U7582 ( .A(n7093), .B(n8310), .Z(n86) );
  COND2X1 U7583 ( .A(n7156), .B(n7286), .C(n7101), .D(n7542), .Z(n1009) );
  COND2X1 U7584 ( .A(n7156), .B(n7350), .C(n7101), .D(n7606), .Z(n1021) );
  COND2X1 U7585 ( .A(n7156), .B(n7318), .C(n7101), .D(n7574), .Z(n1033) );
  CIVX2 U7586 ( .A(n4241), .Z(n7115) );
  COND2X1 U7587 ( .A(n7155), .B(n7323), .C(n7102), .D(n7579), .Z(n1214) );
  COND2X1 U7588 ( .A(n7114), .B(n8008), .C(n7167), .D(n8264), .Z(n650) );
  COND2X1 U7589 ( .A(n7114), .B(n7912), .C(n7167), .D(n8168), .Z(n676) );
  COND2X1 U7590 ( .A(n7114), .B(n7976), .C(n7167), .D(n8232), .Z(n638) );
  COND2X1 U7591 ( .A(n7114), .B(n7944), .C(n7167), .D(n8200), .Z(n664) );
  COND2X1 U7592 ( .A(n7114), .B(n7928), .C(n7167), .D(n8184), .Z(n622) );
  COND2X1 U7593 ( .A(n7114), .B(n7960), .C(n7167), .D(n8216), .Z(n598) );
  COND2X1 U7594 ( .A(n7114), .B(n7992), .C(n7167), .D(n8248), .Z(n610) );
  COND2X1 U7595 ( .A(n7136), .B(n7852), .C(n7130), .D(n8108), .Z(n929) );
  COND2X1 U7596 ( .A(n7137), .B(n7820), .C(n7124), .D(n8076), .Z(n909) );
  COND2X1 U7597 ( .A(n7157), .B(n7308), .C(n7100), .D(n7564), .Z(n908) );
  COND2XL U7598 ( .A(n7133), .B(n7869), .C(n7132), .D(n8125), .Z(n1970) );
  COND2X1 U7599 ( .A(n7133), .B(n7837), .C(n7126), .D(n8093), .Z(n1958) );
  COND2X1 U7600 ( .A(n7133), .B(n7805), .C(n7125), .D(n8061), .Z(n1984) );
  CANR2XL U7601 ( .A(buffer[397]), .B(n6149), .C(buffer[141]), .D(n387), .Z(
        n1157) );
  CND2X1 U7602 ( .A(n2385), .B(n4242), .Z(n1951) );
  CANR2XL U7603 ( .A(buffer[391]), .B(n6149), .C(buffer[135]), .D(n387), .Z(
        n798) );
  CANR2XL U7604 ( .A(buffer[394]), .B(n6149), .C(buffer[138]), .D(n387), .Z(
        n1763) );
  CANR2XL U7605 ( .A(buffer[386]), .B(n6149), .C(buffer[130]), .D(n387), .Z(
        n1612) );
  CANR2XL U7606 ( .A(buffer[389]), .B(n6149), .C(buffer[133]), .D(n387), .Z(
        n1006) );
  COND2X1 U7607 ( .A(n7133), .B(n7781), .C(n7125), .D(n8037), .Z(n1892) );
  CANR2XL U7608 ( .A(buffer[390]), .B(n6149), .C(buffer[134]), .D(n387), .Z(
        n1809) );
  CANR2XL U7609 ( .A(buffer[395]), .B(n6149), .C(buffer[139]), .D(n387), .Z(
        n695) );
  CANR2XL U7610 ( .A(buffer[392]), .B(n6149), .C(buffer[136]), .D(n387), .Z(
        n1310) );
  CNR2X1 U7611 ( .A(n7132), .B(n76), .Z(n41) );
  CANR2XL U7612 ( .A(buffer[384]), .B(n6149), .C(buffer[128]), .D(n387), .Z(
        n1211) );
  CANR2XL U7613 ( .A(buffer[387]), .B(n6149), .C(buffer[131]), .D(n387), .Z(
        n597) );
  CANR2XL U7614 ( .A(buffer[388]), .B(n6149), .C(buffer[132]), .D(n387), .Z(
        n1409) );
  COND2X1 U7615 ( .A(n7133), .B(n7853), .C(n7124), .D(n8109), .Z(n1940) );
  CANR2XL U7616 ( .A(buffer[385]), .B(n6149), .C(buffer[129]), .D(n387), .Z(
        n385) );
  COND2X1 U7617 ( .A(n7133), .B(n7834), .C(n7124), .D(n8090), .Z(n395) );
  COND2X1 U7618 ( .A(n7133), .B(n7821), .C(n7132), .D(n8077), .Z(n1920) );
  CND2X1 U7619 ( .A(n387), .B(n8310), .Z(n80) );
  COND2X1 U7620 ( .A(n29), .B(n156), .C(n65), .D(n7268), .Z(n333) );
  COND3X1 U7621 ( .A(n365), .B(n366), .C(n367), .D(n368), .Z(n3189) );
  COND2XL U7622 ( .A(n7158), .B(n7364), .C(n7100), .D(n7620), .Z(n853) );
  COND2X1 U7623 ( .A(n7158), .B(n7332), .C(n7100), .D(n7588), .Z(n841) );
  COND2X1 U7624 ( .A(n7158), .B(n7316), .C(n7100), .D(n7572), .Z(n825) );
  COND2X1 U7625 ( .A(n7158), .B(n7284), .C(n7100), .D(n7540), .Z(n801) );
  COND2X1 U7626 ( .A(n7158), .B(n7348), .C(n7100), .D(n7604), .Z(n813) );
  COND2X1 U7627 ( .A(n7158), .B(n7255), .C(n7100), .D(n7520), .Z(n780) );
  CAOR2XL U7628 ( .A(n36), .B(n8303), .C(n38), .D(n39), .Z(n30) );
  CANR2XL U7629 ( .A(n39), .B(n216), .C(n8301), .D(n217), .Z(n213) );
  CAOR2XL U7630 ( .A(n166), .B(n8303), .C(n167), .D(n39), .Z(n162) );
  CANR2XL U7631 ( .A(n39), .B(n254), .C(n8301), .D(n255), .Z(n251) );
  CANR2XL U7632 ( .A(n39), .B(n125), .C(n8303), .D(n126), .Z(n124) );
  CANR2X1 U7633 ( .A(n39), .B(n192), .C(n8303), .D(n193), .Z(n189) );
  CANR2X1 U7634 ( .A(n39), .B(n323), .C(n8301), .D(n324), .Z(n320) );
  CANR2X1 U7635 ( .A(n39), .B(n297), .C(n8303), .D(n298), .Z(n294) );
  CANR2X1 U7636 ( .A(n39), .B(n276), .C(n8301), .D(n277), .Z(n273) );
  CND2XL U7637 ( .A(rd_ptr[9]), .B(n8311), .Z(n382) );
  COND2X1 U7638 ( .A(n7115), .B(n7948), .C(n7166), .D(n8204), .Z(n910) );
  CIVX1 U7639 ( .A(n4240), .Z(n7157) );
  COND2X1 U7640 ( .A(n7159), .B(n7312), .C(n7099), .D(n7568), .Z(n726) );
  CIVX1 U7641 ( .A(n4240), .Z(n7159) );
  CAOR2XL U7642 ( .A(N16597), .B(n6165), .C(n7091), .D(n4239), .Z(n3192) );
  CND3XL U7643 ( .A(n6161), .B(n262), .C(n7170), .Z(n259) );
  CEOXL U7644 ( .A(n4239), .B(\add_121/carry [7]), .Z(N16597) );
  CAN2XL U7645 ( .A(\add_121/carry [7]), .B(n4239), .Z(\add_121/carry [8]) );
  CNR2XL U7646 ( .A(n76), .B(n4239), .Z(n39) );
  COND2XL U7647 ( .A(n7119), .B(n7911), .C(n7163), .D(n8167), .Z(n1488) );
  COND2XL U7648 ( .A(n7119), .B(n8007), .C(n7163), .D(n8263), .Z(n1462) );
  COND2X1 U7649 ( .A(n7119), .B(n7943), .C(n7163), .D(n8199), .Z(n1476) );
  COND2X1 U7650 ( .A(n7119), .B(n7975), .C(n7163), .D(n8231), .Z(n1450) );
  COND2X1 U7651 ( .A(n7119), .B(n7959), .C(n7163), .D(n8215), .Z(n1434) );
  COND2X1 U7652 ( .A(n7119), .B(n7991), .C(n7163), .D(n8247), .Z(n1422) );
  COND2X1 U7653 ( .A(n7119), .B(n7927), .C(n7163), .D(n8183), .Z(n1410) );
  CND2X1 U7654 ( .A(n4239), .B(n386), .Z(n396) );
  COND3X1 U7655 ( .A(n900), .B(n8013), .C(n1913), .D(n1914), .Z(n1905) );
  CANR2XL U7656 ( .A(n7245), .B(n8288), .C(n314), .D(n8289), .Z(n354) );
  COND2XL U7657 ( .A(n314), .B(n16), .C(n7245), .D(n21), .Z(n353) );
  COND2XL U7658 ( .A(n314), .B(n19), .C(n1200), .D(n14), .Z(n1195) );
  COND2XL U7659 ( .A(n7503), .B(n92), .C(n93), .D(n94), .Z(n90) );
  COND2X1 U7660 ( .A(n94), .B(n35), .C(n8300), .D(n7759), .Z(n1502) );
  COND2XL U7661 ( .A(n7153), .B(n7343), .C(n7104), .D(n7599), .Z(n1525) );
  COND2X1 U7662 ( .A(n7153), .B(n7375), .C(n7104), .D(n7631), .Z(n1520) );
  COND2X1 U7663 ( .A(n7153), .B(n7359), .C(n7104), .D(n7615), .Z(n1555) );
  COND2X1 U7664 ( .A(n7153), .B(n7295), .C(n7104), .D(n7551), .Z(n1581) );
  COND2X1 U7665 ( .A(n7153), .B(n7311), .C(n7104), .D(n7567), .Z(n1507) );
  CIVX1 U7666 ( .A(n370), .Z(n7246) );
  COND3X1 U7667 ( .A(n7252), .B(n19), .C(n372), .D(n373), .Z(n370) );
  CND4X1 U7668 ( .A(n689), .B(n690), .C(n691), .D(n692), .Z(n688) );
  CANR2X1 U7669 ( .A(n7096), .B(n7760), .C(n8301), .D(n126), .Z(n689) );
  CANR2X1 U7670 ( .A(n39), .B(n339), .C(n8303), .D(n340), .Z(n336) );
  CANR2X1 U7671 ( .A(buffer[1025]), .B(n8304), .C(buffer[769]), .D(n8305), .Z(
        n337) );
  CIVX1 U7672 ( .A(n4241), .Z(n7112) );
  COND3X1 U7673 ( .A(n900), .B(n8012), .C(n902), .D(n903), .Z(n893) );
  COND2XL U7674 ( .A(n7123), .B(n7997), .C(n7161), .D(n8253), .Z(n1967) );
  COND2XL U7675 ( .A(n7118), .B(n7901), .C(n7164), .D(n8157), .Z(n1993) );
  COND2XL U7676 ( .A(n7123), .B(n7965), .C(n7161), .D(n8221), .Z(n1955) );
  COND2X1 U7677 ( .A(n7118), .B(n7933), .C(n7161), .D(n8189), .Z(n1981) );
  COND2X1 U7678 ( .A(n7119), .B(n7917), .C(n7161), .D(n8173), .Z(n1931) );
  COND2X1 U7679 ( .A(n7112), .B(n7981), .C(n7161), .D(n8237), .Z(n1937) );
  COND2X1 U7680 ( .A(n7115), .B(n7949), .C(n7161), .D(n8205), .Z(n1921) );
  CIVX1 U7681 ( .A(n4240), .Z(n7160) );
  COND3X1 U7682 ( .A(n7241), .B(n286), .C(n303), .D(n304), .Z(n3186) );
  COND3XL U7683 ( .A(n111), .B(n69), .C(n112), .D(n113), .Z(n48) );
  COND2X1 U7684 ( .A(n29), .B(n111), .C(n65), .D(n7265), .Z(n291) );
  COND2XL U7685 ( .A(n7155), .B(n7257), .C(n7099), .D(n7522), .Z(n578) );
  COND2XL U7686 ( .A(n7159), .B(n7368), .C(n7099), .D(n7624), .Z(n652) );
  COND2XL U7687 ( .A(n7159), .B(n7336), .C(n7099), .D(n7592), .Z(n640) );
  COND2X1 U7688 ( .A(n13), .B(n14), .C(n7230), .D(n16), .Z(n12) );
  COND3X1 U7689 ( .A(n13), .B(n16), .C(n108), .D(n109), .Z(n54) );
  COND3X1 U7690 ( .A(n13), .B(n19), .C(n153), .D(n154), .Z(n131) );
  COND4CX1 U7691 ( .A(n890), .B(n891), .C(n8296), .D(n892), .Z(n889) );
  CIVX1 U7692 ( .A(n4240), .Z(n7154) );
  CND2XL U7693 ( .A(n8288), .B(n105), .Z(n224) );
  CANR2XL U7694 ( .A(n8288), .B(n107), .C(n8289), .D(n105), .Z(n132) );
  COND2X1 U7695 ( .A(rd_ptr[2]), .B(n105), .C(n8290), .D(n107), .Z(n56) );
  COND4CX1 U7696 ( .A(n1902), .B(n1903), .C(n8296), .D(n1904), .Z(n1901) );
  COND2XL U7697 ( .A(n7151), .B(n7357), .C(n7107), .D(n7613), .Z(n1969) );
  COND2XL U7698 ( .A(n7150), .B(n7251), .C(n7107), .D(n7517), .Z(n1995) );
  COND2XL U7699 ( .A(n7153), .B(n7325), .C(n7106), .D(n7581), .Z(n1957) );
  COND2XL U7700 ( .A(n7159), .B(n7293), .C(n7107), .D(n7549), .Z(n1983) );
  COND2XL U7701 ( .A(n7154), .B(n7261), .C(n7106), .D(n7525), .Z(n1891) );
  COND2X1 U7702 ( .A(n7157), .B(n7341), .C(n7106), .D(n7597), .Z(n1939) );
  COND2X1 U7703 ( .A(n7160), .B(n7309), .C(n7106), .D(n7565), .Z(n1919) );
  CND2XL U7704 ( .A(n942), .B(n8306), .Z(n92) );
  CANR2XL U7705 ( .A(n2850), .B(n942), .C(n2851), .D(n4240), .Z(n941) );
  CANR2XL U7706 ( .A(n2387), .B(n942), .C(n2388), .D(n4240), .Z(n1952) );
  COND4CXL U7707 ( .A(rd_ptr[1]), .B(n352), .C(n1195), .D(n3173), .Z(n366) );
  COND2X1 U7708 ( .A(n97), .B(n349), .C(n7246), .D(n8), .Z(n346) );
  COND4CX1 U7709 ( .A(n352), .B(n8287), .C(n353), .D(n6163), .Z(n351) );
  CANR2XL U7710 ( .A(n8288), .B(n207), .C(n8289), .D(n288), .Z(n331) );
  CAN3X1 U7711 ( .A(n203), .B(n199), .C(n7171), .Z(n204) );
  CANR2XL U7712 ( .A(n8288), .B(n129), .C(n8289), .D(n207), .Z(n246) );
  COND3X1 U7713 ( .A(n13), .B(n21), .C(n205), .D(n206), .Z(n199) );
  CANR2X1 U7714 ( .A(n8289), .B(n155), .C(n8285), .D(n207), .Z(n206) );
  COND3XL U7715 ( .A(n258), .B(n8), .C(n259), .D(n260), .Z(n3184) );
  COND3X1 U7716 ( .A(n7214), .B(n8), .C(n281), .D(n282), .Z(n3185) );
  COND3XL U7717 ( .A(n6158), .B(n7641), .C(n1611), .D(n1612), .Z(n323) );
  COND3XL U7718 ( .A(n6158), .B(n7633), .C(n1762), .D(n1763), .Z(n145) );
  COND3XL U7719 ( .A(n6158), .B(n7637), .C(n1808), .D(n1809), .Z(n235) );
  COND3XL U7720 ( .A(n6158), .B(n7630), .C(n1156), .D(n1157), .Z(n38) );
  COND3XL U7721 ( .A(n6158), .B(n7638), .C(n1005), .D(n1006), .Z(n254) );
  COND3XL U7722 ( .A(n6158), .B(n7636), .C(n797), .D(n798), .Z(n216) );
  COND3XL U7723 ( .A(n6158), .B(n7643), .C(n1210), .D(n1211), .Z(n361) );
  COND3XL U7724 ( .A(n6158), .B(n7632), .C(n694), .D(n695), .Z(n125) );
  COND3XL U7725 ( .A(n6158), .B(n7635), .C(n1309), .D(n1310), .Z(n192) );
  COND3XL U7726 ( .A(n6158), .B(n7639), .C(n1408), .D(n1409), .Z(n276) );
  COND3XL U7727 ( .A(n6158), .B(n7640), .C(n596), .D(n597), .Z(n297) );
  COND3XL U7728 ( .A(n6158), .B(n7642), .C(n384), .D(n385), .Z(n339) );
  COND3XL U7729 ( .A(n6158), .B(n7634), .C(n495), .D(n496), .Z(n167) );
  CNR2XL U7730 ( .A(n382), .B(n8310), .Z(n942) );
  CIVX1 U7731 ( .A(n6177), .Z(n6179) );
  CIVX1 U7732 ( .A(n6179), .Z(n6180) );
  CIVX1 U7733 ( .A(n6179), .Z(n6181) );
  CIVX1 U7734 ( .A(n6186), .Z(n6182) );
  CIVX1 U7735 ( .A(n6179), .Z(n6183) );
  CIVX1 U7736 ( .A(n6179), .Z(n6184) );
  CIVX1 U7737 ( .A(n6179), .Z(n6185) );
  CIVX1 U7738 ( .A(n6178), .Z(n6186) );
  CIVX1 U7739 ( .A(n6186), .Z(n6187) );
  CIVX1 U7740 ( .A(n6186), .Z(n6188) );
  CIVX1 U7741 ( .A(n6186), .Z(n6189) );
  CIVX1 U7742 ( .A(n6186), .Z(n6190) );
  CIVX1 U7743 ( .A(n6193), .Z(n6191) );
  CIVX1 U7744 ( .A(n6193), .Z(n6192) );
  CIVX1 U7745 ( .A(n2218), .Z(n6193) );
  CIVX1 U7746 ( .A(n6193), .Z(n6194) );
  CIVX1 U7747 ( .A(n6193), .Z(n6195) );
  CIVX1 U7748 ( .A(n6193), .Z(n6196) );
  CIVX1 U7749 ( .A(n6193), .Z(n6197) );
  CIVX1 U7750 ( .A(n6179), .Z(n6198) );
  CIVX1 U7751 ( .A(n6193), .Z(n6199) );
  CIVX1 U7752 ( .A(n6207), .Z(n6209) );
  CIVX1 U7753 ( .A(n6209), .Z(n6210) );
  CIVX1 U7754 ( .A(n6209), .Z(n6211) );
  CIVX1 U7755 ( .A(n6216), .Z(n6212) );
  CIVX1 U7756 ( .A(n6209), .Z(n6213) );
  CIVX1 U7757 ( .A(n6209), .Z(n6214) );
  CIVX1 U7758 ( .A(n6209), .Z(n6215) );
  CIVX1 U7759 ( .A(n6208), .Z(n6216) );
  CIVX1 U7760 ( .A(n6216), .Z(n6217) );
  CIVX1 U7761 ( .A(n6216), .Z(n6218) );
  CIVX1 U7762 ( .A(n6223), .Z(n6219) );
  CIVX1 U7763 ( .A(n6223), .Z(n6220) );
  CIVX1 U7764 ( .A(n6216), .Z(n6221) );
  CIVX1 U7765 ( .A(n6216), .Z(n6222) );
  CIVX1 U7766 ( .A(n2216), .Z(n6223) );
  CIVX1 U7767 ( .A(n6223), .Z(n6224) );
  CIVX1 U7768 ( .A(n6223), .Z(n6225) );
  CIVX1 U7769 ( .A(n6223), .Z(n6226) );
  CIVX1 U7770 ( .A(n6223), .Z(n6227) );
  CIVX1 U7771 ( .A(n6209), .Z(n6228) );
  CIVX1 U7772 ( .A(n6223), .Z(n6229) );
  CIVX1 U7773 ( .A(n6237), .Z(n6239) );
  CIVX1 U7774 ( .A(n6239), .Z(n6240) );
  CIVX1 U7775 ( .A(n6239), .Z(n6241) );
  CIVX1 U7776 ( .A(n6246), .Z(n6242) );
  CIVX1 U7777 ( .A(n6239), .Z(n6243) );
  CIVX1 U7778 ( .A(n6239), .Z(n6244) );
  CIVX1 U7779 ( .A(n6239), .Z(n6245) );
  CIVX1 U7780 ( .A(n6238), .Z(n6246) );
  CIVX1 U7781 ( .A(n6246), .Z(n6247) );
  CIVX1 U7782 ( .A(n6246), .Z(n6248) );
  CIVX1 U7783 ( .A(n6253), .Z(n6249) );
  CIVX1 U7784 ( .A(n6253), .Z(n6250) );
  CIVX1 U7785 ( .A(n6246), .Z(n6251) );
  CIVX1 U7786 ( .A(n6246), .Z(n6252) );
  CIVX1 U7787 ( .A(n2214), .Z(n6253) );
  CIVX1 U7788 ( .A(n6253), .Z(n6254) );
  CIVX1 U7789 ( .A(n6253), .Z(n6255) );
  CIVX1 U7790 ( .A(n6253), .Z(n6256) );
  CIVX1 U7791 ( .A(n6253), .Z(n6257) );
  CIVX1 U7792 ( .A(n6239), .Z(n6258) );
  CIVX1 U7793 ( .A(n6253), .Z(n6259) );
  CIVX1 U7794 ( .A(n6267), .Z(n6269) );
  CIVX1 U7795 ( .A(n6269), .Z(n6270) );
  CIVX1 U7796 ( .A(n6269), .Z(n6271) );
  CIVX1 U7797 ( .A(n6276), .Z(n6272) );
  CIVX1 U7798 ( .A(n6269), .Z(n6273) );
  CIVX1 U7799 ( .A(n6269), .Z(n6274) );
  CIVX1 U7800 ( .A(n6269), .Z(n6275) );
  CIVX1 U7801 ( .A(n6268), .Z(n6276) );
  CIVX1 U7802 ( .A(n6276), .Z(n6277) );
  CIVX1 U7803 ( .A(n6276), .Z(n6278) );
  CIVX1 U7804 ( .A(n6276), .Z(n6279) );
  CIVX1 U7805 ( .A(n6276), .Z(n6280) );
  CIVX1 U7806 ( .A(n6283), .Z(n6281) );
  CIVX1 U7807 ( .A(n6283), .Z(n6282) );
  CIVX1 U7808 ( .A(n2198), .Z(n6283) );
  CIVX1 U7809 ( .A(n6283), .Z(n6284) );
  CIVX1 U7810 ( .A(n6283), .Z(n6285) );
  CIVX1 U7811 ( .A(n6283), .Z(n6286) );
  CIVX1 U7812 ( .A(n6283), .Z(n6287) );
  CIVX1 U7813 ( .A(n6269), .Z(n6288) );
  CIVX1 U7814 ( .A(n6283), .Z(n6289) );
  CIVX1 U7815 ( .A(n6297), .Z(n6299) );
  CIVX1 U7816 ( .A(n6299), .Z(n6300) );
  CIVX1 U7817 ( .A(n6299), .Z(n6301) );
  CIVX1 U7818 ( .A(n6306), .Z(n6302) );
  CIVX1 U7819 ( .A(n6299), .Z(n6303) );
  CIVX1 U7820 ( .A(n6299), .Z(n6304) );
  CIVX1 U7821 ( .A(n6299), .Z(n6305) );
  CIVX1 U7822 ( .A(n6298), .Z(n6306) );
  CIVX1 U7823 ( .A(n6306), .Z(n6307) );
  CIVX1 U7824 ( .A(n6306), .Z(n6308) );
  CIVX1 U7825 ( .A(n6313), .Z(n6309) );
  CIVX1 U7826 ( .A(n6313), .Z(n6310) );
  CIVX1 U7827 ( .A(n6306), .Z(n6311) );
  CIVX1 U7828 ( .A(n6306), .Z(n6312) );
  CIVX1 U7829 ( .A(n2195), .Z(n6313) );
  CIVX1 U7830 ( .A(n6313), .Z(n6314) );
  CIVX1 U7831 ( .A(n6313), .Z(n6315) );
  CIVX1 U7832 ( .A(n6313), .Z(n6316) );
  CIVX1 U7833 ( .A(n6313), .Z(n6317) );
  CIVX1 U7834 ( .A(n6299), .Z(n6318) );
  CIVX1 U7835 ( .A(n6313), .Z(n6319) );
  CIVX1 U7836 ( .A(n6327), .Z(n6329) );
  CIVX1 U7837 ( .A(n6329), .Z(n6330) );
  CIVX1 U7838 ( .A(n6329), .Z(n6331) );
  CIVX1 U7839 ( .A(n6336), .Z(n6332) );
  CIVX1 U7840 ( .A(n6329), .Z(n6333) );
  CIVX1 U7841 ( .A(n6329), .Z(n6334) );
  CIVX1 U7842 ( .A(n6329), .Z(n6335) );
  CIVX1 U7843 ( .A(n6328), .Z(n6336) );
  CIVX1 U7844 ( .A(n6336), .Z(n6337) );
  CIVX1 U7845 ( .A(n6336), .Z(n6338) );
  CIVX1 U7846 ( .A(n6343), .Z(n6339) );
  CIVX1 U7847 ( .A(n6343), .Z(n6340) );
  CIVX1 U7848 ( .A(n6336), .Z(n6341) );
  CIVX1 U7849 ( .A(n6336), .Z(n6342) );
  CIVX1 U7850 ( .A(n2193), .Z(n6343) );
  CIVX1 U7851 ( .A(n6343), .Z(n6344) );
  CIVX1 U7852 ( .A(n6343), .Z(n6345) );
  CIVX1 U7853 ( .A(n6343), .Z(n6346) );
  CIVX1 U7854 ( .A(n6343), .Z(n6347) );
  CIVX1 U7855 ( .A(n6329), .Z(n6348) );
  CIVX1 U7856 ( .A(n6343), .Z(n6349) );
  CIVX1 U7857 ( .A(n6357), .Z(n6359) );
  CIVX1 U7858 ( .A(n6359), .Z(n6360) );
  CIVX1 U7859 ( .A(n6359), .Z(n6361) );
  CIVX1 U7860 ( .A(n6366), .Z(n6362) );
  CIVX1 U7861 ( .A(n6359), .Z(n6363) );
  CIVX1 U7862 ( .A(n6359), .Z(n6364) );
  CIVX1 U7863 ( .A(n6359), .Z(n6365) );
  CIVX1 U7864 ( .A(n6358), .Z(n6366) );
  CIVX1 U7865 ( .A(n6366), .Z(n6367) );
  CIVX1 U7866 ( .A(n6366), .Z(n6368) );
  CIVX1 U7867 ( .A(n6373), .Z(n6369) );
  CIVX1 U7868 ( .A(n6373), .Z(n6370) );
  CIVX1 U7869 ( .A(n6366), .Z(n6371) );
  CIVX1 U7870 ( .A(n6366), .Z(n6372) );
  CIVX1 U7871 ( .A(n2191), .Z(n6373) );
  CIVX1 U7872 ( .A(n6373), .Z(n6374) );
  CIVX1 U7873 ( .A(n6373), .Z(n6375) );
  CIVX1 U7874 ( .A(n6373), .Z(n6376) );
  CIVX1 U7875 ( .A(n6373), .Z(n6377) );
  CIVX1 U7876 ( .A(n6359), .Z(n6378) );
  CIVX1 U7877 ( .A(n6373), .Z(n6379) );
  CIVX1 U7878 ( .A(n6387), .Z(n6389) );
  CIVX1 U7879 ( .A(n6389), .Z(n6390) );
  CIVX1 U7880 ( .A(n6389), .Z(n6391) );
  CIVX1 U7881 ( .A(n6396), .Z(n6392) );
  CIVX1 U7882 ( .A(n6389), .Z(n6393) );
  CIVX1 U7883 ( .A(n6389), .Z(n6394) );
  CIVX1 U7884 ( .A(n6389), .Z(n6395) );
  CIVX1 U7885 ( .A(n6388), .Z(n6396) );
  CIVX1 U7886 ( .A(n6396), .Z(n6397) );
  CIVX1 U7887 ( .A(n6396), .Z(n6398) );
  CIVX1 U7888 ( .A(n6396), .Z(n6399) );
  CIVX1 U7889 ( .A(n6396), .Z(n6400) );
  CIVX1 U7890 ( .A(n6403), .Z(n6401) );
  CIVX1 U7891 ( .A(n6403), .Z(n6402) );
  CIVX1 U7892 ( .A(n2176), .Z(n6403) );
  CIVX1 U7893 ( .A(n6403), .Z(n6404) );
  CIVX1 U7894 ( .A(n6403), .Z(n6405) );
  CIVX1 U7895 ( .A(n6403), .Z(n6406) );
  CIVX1 U7896 ( .A(n6403), .Z(n6407) );
  CIVX1 U7897 ( .A(n6389), .Z(n6408) );
  CIVX1 U7898 ( .A(n6403), .Z(n6409) );
  CIVX1 U7899 ( .A(n6417), .Z(n6419) );
  CIVX1 U7900 ( .A(n6419), .Z(n6420) );
  CIVX1 U7901 ( .A(n6419), .Z(n6421) );
  CIVX1 U7902 ( .A(n6426), .Z(n6422) );
  CIVX1 U7903 ( .A(n6419), .Z(n6423) );
  CIVX1 U7904 ( .A(n6419), .Z(n6424) );
  CIVX1 U7905 ( .A(n6419), .Z(n6425) );
  CIVX1 U7906 ( .A(n6418), .Z(n6426) );
  CIVX1 U7907 ( .A(n6426), .Z(n6427) );
  CIVX1 U7908 ( .A(n6426), .Z(n6428) );
  CIVX1 U7909 ( .A(n6433), .Z(n6429) );
  CIVX1 U7910 ( .A(n6433), .Z(n6430) );
  CIVX1 U7911 ( .A(n6426), .Z(n6431) );
  CIVX1 U7912 ( .A(n6426), .Z(n6432) );
  CIVX1 U7913 ( .A(n2173), .Z(n6433) );
  CIVX1 U7914 ( .A(n6433), .Z(n6434) );
  CIVX1 U7915 ( .A(n6433), .Z(n6435) );
  CIVX1 U7916 ( .A(n6433), .Z(n6436) );
  CIVX1 U7917 ( .A(n6433), .Z(n6437) );
  CIVX1 U7918 ( .A(n6419), .Z(n6438) );
  CIVX1 U7919 ( .A(n6433), .Z(n6439) );
  CIVX1 U7920 ( .A(n6447), .Z(n6449) );
  CIVX1 U7921 ( .A(n6449), .Z(n6450) );
  CIVX1 U7922 ( .A(n6449), .Z(n6451) );
  CIVX1 U7923 ( .A(n6456), .Z(n6452) );
  CIVX1 U7924 ( .A(n6449), .Z(n6453) );
  CIVX1 U7925 ( .A(n6449), .Z(n6454) );
  CIVX1 U7926 ( .A(n6449), .Z(n6455) );
  CIVX1 U7927 ( .A(n6448), .Z(n6456) );
  CIVX1 U7928 ( .A(n6456), .Z(n6457) );
  CIVX1 U7929 ( .A(n6456), .Z(n6458) );
  CIVX1 U7930 ( .A(n6463), .Z(n6459) );
  CIVX1 U7931 ( .A(n6463), .Z(n6460) );
  CIVX1 U7932 ( .A(n6456), .Z(n6461) );
  CIVX1 U7933 ( .A(n6456), .Z(n6462) );
  CIVX1 U7934 ( .A(n2171), .Z(n6463) );
  CIVX1 U7935 ( .A(n6463), .Z(n6464) );
  CIVX1 U7936 ( .A(n6463), .Z(n6465) );
  CIVX1 U7937 ( .A(n6463), .Z(n6466) );
  CIVX1 U7938 ( .A(n6463), .Z(n6467) );
  CIVX1 U7939 ( .A(n6449), .Z(n6468) );
  CIVX1 U7940 ( .A(n6463), .Z(n6469) );
  CIVX1 U7941 ( .A(n6477), .Z(n6479) );
  CIVX1 U7942 ( .A(n6479), .Z(n6480) );
  CIVX1 U7943 ( .A(n6479), .Z(n6481) );
  CIVX1 U7944 ( .A(n6486), .Z(n6482) );
  CIVX1 U7945 ( .A(n6479), .Z(n6483) );
  CIVX1 U7946 ( .A(n6479), .Z(n6484) );
  CIVX1 U7947 ( .A(n6479), .Z(n6485) );
  CIVX1 U7948 ( .A(n6478), .Z(n6486) );
  CIVX1 U7949 ( .A(n6486), .Z(n6487) );
  CIVX1 U7950 ( .A(n6486), .Z(n6488) );
  CIVX1 U7951 ( .A(n6493), .Z(n6489) );
  CIVX1 U7952 ( .A(n6493), .Z(n6490) );
  CIVX1 U7953 ( .A(n6486), .Z(n6491) );
  CIVX1 U7954 ( .A(n6486), .Z(n6492) );
  CIVX1 U7955 ( .A(n2168), .Z(n6493) );
  CIVX1 U7956 ( .A(n6493), .Z(n6494) );
  CIVX1 U7957 ( .A(n6493), .Z(n6495) );
  CIVX1 U7958 ( .A(n6493), .Z(n6496) );
  CIVX1 U7959 ( .A(n6493), .Z(n6497) );
  CIVX1 U7960 ( .A(n6479), .Z(n6498) );
  CIVX1 U7961 ( .A(n6493), .Z(n6499) );
  CIVX1 U7962 ( .A(n6507), .Z(n6509) );
  CIVX1 U7963 ( .A(n6509), .Z(n6510) );
  CIVX1 U7964 ( .A(n6509), .Z(n6511) );
  CIVX1 U7965 ( .A(n6523), .Z(n6512) );
  CIVX1 U7966 ( .A(n6509), .Z(n6513) );
  CIVX1 U7967 ( .A(n6509), .Z(n6514) );
  CIVX1 U7968 ( .A(n6509), .Z(n6515) );
  CIVX1 U7969 ( .A(n6508), .Z(n6516) );
  CIVX1 U7970 ( .A(n6516), .Z(n6517) );
  CIVX1 U7971 ( .A(n6516), .Z(n6518) );
  CIVX1 U7972 ( .A(n6516), .Z(n6519) );
  CIVX1 U7973 ( .A(n6516), .Z(n6520) );
  CIVX1 U7974 ( .A(n6516), .Z(n6521) );
  CIVX1 U7975 ( .A(n6523), .Z(n6522) );
  CIVX1 U7976 ( .A(n2164), .Z(n6523) );
  CIVX1 U7977 ( .A(n6523), .Z(n6524) );
  CIVX1 U7978 ( .A(n6523), .Z(n6525) );
  CIVX1 U7979 ( .A(n6523), .Z(n6526) );
  CIVX1 U7980 ( .A(n6523), .Z(n6527) );
  CIVX1 U7981 ( .A(n6523), .Z(n6528) );
  CIVX1 U7982 ( .A(n6516), .Z(n6529) );
  CIVX1 U7983 ( .A(n6537), .Z(n6539) );
  CIVX1 U7984 ( .A(n6539), .Z(n6540) );
  CIVX1 U7985 ( .A(n6539), .Z(n6541) );
  CIVX1 U7986 ( .A(n6546), .Z(n6542) );
  CIVX1 U7987 ( .A(n6539), .Z(n6543) );
  CIVX1 U7988 ( .A(n6539), .Z(n6544) );
  CIVX1 U7989 ( .A(n6539), .Z(n6545) );
  CIVX1 U7990 ( .A(n6538), .Z(n6546) );
  CIVX1 U7991 ( .A(n6546), .Z(n6547) );
  CIVX1 U7992 ( .A(n6546), .Z(n6548) );
  CIVX1 U7993 ( .A(n6553), .Z(n6549) );
  CIVX1 U7994 ( .A(n6553), .Z(n6550) );
  CIVX1 U7995 ( .A(n6546), .Z(n6551) );
  CIVX1 U7996 ( .A(n6546), .Z(n6552) );
  CIVX1 U7997 ( .A(n2161), .Z(n6553) );
  CIVX1 U7998 ( .A(n6553), .Z(n6554) );
  CIVX1 U7999 ( .A(n6553), .Z(n6555) );
  CIVX1 U8000 ( .A(n6553), .Z(n6556) );
  CIVX1 U8001 ( .A(n6553), .Z(n6557) );
  CIVX1 U8002 ( .A(n6539), .Z(n6558) );
  CIVX1 U8003 ( .A(n6553), .Z(n6559) );
  CIVX1 U8004 ( .A(n6567), .Z(n6569) );
  CIVX1 U8005 ( .A(n6569), .Z(n6570) );
  CIVX1 U8006 ( .A(n6569), .Z(n6571) );
  CIVX1 U8007 ( .A(n6576), .Z(n6572) );
  CIVX1 U8008 ( .A(n6569), .Z(n6573) );
  CIVX1 U8009 ( .A(n6569), .Z(n6574) );
  CIVX1 U8010 ( .A(n6569), .Z(n6575) );
  CIVX1 U8011 ( .A(n6568), .Z(n6576) );
  CIVX1 U8012 ( .A(n6576), .Z(n6577) );
  CIVX1 U8013 ( .A(n6576), .Z(n6578) );
  CIVX1 U8014 ( .A(n6583), .Z(n6579) );
  CIVX1 U8015 ( .A(n6583), .Z(n6580) );
  CIVX1 U8016 ( .A(n6576), .Z(n6581) );
  CIVX1 U8017 ( .A(n6576), .Z(n6582) );
  CIVX1 U8018 ( .A(n2159), .Z(n6583) );
  CIVX1 U8019 ( .A(n6583), .Z(n6584) );
  CIVX1 U8020 ( .A(n6583), .Z(n6585) );
  CIVX1 U8021 ( .A(n6583), .Z(n6586) );
  CIVX1 U8022 ( .A(n6583), .Z(n6587) );
  CIVX1 U8023 ( .A(n6569), .Z(n6588) );
  CIVX1 U8024 ( .A(n6583), .Z(n6589) );
  CIVX1 U8025 ( .A(n6597), .Z(n6599) );
  CIVX1 U8026 ( .A(n6599), .Z(n6600) );
  CIVX1 U8027 ( .A(n6599), .Z(n6601) );
  CIVX1 U8028 ( .A(n6599), .Z(n6602) );
  CIVX1 U8029 ( .A(n6599), .Z(n6603) );
  CIVX1 U8030 ( .A(n6599), .Z(n6604) );
  CIVX1 U8031 ( .A(n6599), .Z(n6605) );
  CIVX1 U8032 ( .A(n6598), .Z(n6606) );
  CIVX1 U8033 ( .A(n6606), .Z(n6607) );
  CIVX1 U8034 ( .A(n6606), .Z(n6608) );
  CIVX1 U8035 ( .A(n6606), .Z(n6609) );
  CIVX1 U8036 ( .A(n6606), .Z(n6610) );
  CIVX1 U8037 ( .A(n6606), .Z(n6611) );
  CIVX1 U8038 ( .A(n6606), .Z(n6612) );
  CIVX1 U8039 ( .A(n2156), .Z(n6613) );
  CIVX1 U8040 ( .A(n6613), .Z(n6614) );
  CIVX1 U8041 ( .A(n6613), .Z(n6615) );
  CIVX1 U8042 ( .A(n6613), .Z(n6616) );
  CIVX1 U8043 ( .A(n6613), .Z(n6617) );
  CIVX1 U8044 ( .A(n6613), .Z(n6618) );
  CIVX1 U8045 ( .A(n6613), .Z(n6619) );
  CIVX1 U8046 ( .A(n6627), .Z(n6629) );
  CIVX1 U8047 ( .A(n6629), .Z(n6630) );
  CIVX1 U8048 ( .A(n6629), .Z(n6631) );
  CIVX1 U8049 ( .A(n6629), .Z(n6632) );
  CIVX1 U8050 ( .A(n6629), .Z(n6633) );
  CIVX1 U8051 ( .A(n6629), .Z(n6634) );
  CIVX1 U8052 ( .A(n6629), .Z(n6635) );
  CIVX1 U8053 ( .A(n6628), .Z(n6636) );
  CIVX1 U8054 ( .A(n6636), .Z(n6637) );
  CIVX1 U8055 ( .A(n6636), .Z(n6638) );
  CIVX1 U8056 ( .A(n6636), .Z(n6639) );
  CIVX1 U8057 ( .A(n6636), .Z(n6640) );
  CIVX1 U8058 ( .A(n6636), .Z(n6641) );
  CIVX1 U8059 ( .A(n6636), .Z(n6642) );
  CIVX1 U8060 ( .A(n2140), .Z(n6643) );
  CIVX1 U8061 ( .A(n6643), .Z(n6644) );
  CIVX1 U8062 ( .A(n6643), .Z(n6645) );
  CIVX1 U8063 ( .A(n6643), .Z(n6646) );
  CIVX1 U8064 ( .A(n6643), .Z(n6647) );
  CIVX1 U8065 ( .A(n6643), .Z(n6648) );
  CIVX1 U8066 ( .A(n6643), .Z(n6649) );
  CIVX1 U8067 ( .A(n6654), .Z(n6656) );
  CIVX1 U8068 ( .A(n6656), .Z(n6657) );
  CIVX1 U8069 ( .A(n6656), .Z(n6658) );
  CIVX1 U8070 ( .A(n6656), .Z(n6659) );
  CIVX1 U8071 ( .A(n6656), .Z(n6660) );
  CIVX1 U8072 ( .A(n6656), .Z(n6661) );
  CIVX1 U8073 ( .A(n6656), .Z(n6662) );
  CIVX1 U8074 ( .A(n6655), .Z(n6663) );
  CIVX1 U8075 ( .A(n6663), .Z(n6664) );
  CIVX1 U8076 ( .A(n6663), .Z(n6665) );
  CIVX1 U8077 ( .A(n6663), .Z(n6666) );
  CIVX1 U8078 ( .A(n6663), .Z(n6667) );
  CIVX1 U8079 ( .A(n6663), .Z(n6668) );
  CIVX1 U8080 ( .A(n6663), .Z(n6669) );
  CIVX1 U8081 ( .A(n2136), .Z(n6670) );
  CIVX1 U8082 ( .A(n6670), .Z(n6671) );
  CIVX1 U8083 ( .A(n6670), .Z(n6672) );
  CIVX1 U8084 ( .A(n6670), .Z(n6673) );
  CIVX1 U8085 ( .A(n6670), .Z(n6674) );
  CIVX1 U8086 ( .A(n6670), .Z(n6675) );
  CIVX1 U8087 ( .A(n6670), .Z(n6676) );
  CIVX1 U8088 ( .A(n6681), .Z(n6683) );
  CIVX1 U8089 ( .A(n6683), .Z(n6684) );
  CIVX1 U8090 ( .A(n6683), .Z(n6685) );
  CIVX1 U8091 ( .A(n6683), .Z(n6686) );
  CIVX1 U8092 ( .A(n6683), .Z(n6687) );
  CIVX1 U8093 ( .A(n6683), .Z(n6688) );
  CIVX1 U8094 ( .A(n6683), .Z(n6689) );
  CIVX1 U8095 ( .A(n6682), .Z(n6690) );
  CIVX1 U8096 ( .A(n6690), .Z(n6691) );
  CIVX1 U8097 ( .A(n6690), .Z(n6692) );
  CIVX1 U8098 ( .A(n6690), .Z(n6693) );
  CIVX1 U8099 ( .A(n6690), .Z(n6694) );
  CIVX1 U8100 ( .A(n6690), .Z(n6695) );
  CIVX1 U8101 ( .A(n6690), .Z(n6696) );
  CIVX1 U8102 ( .A(n2133), .Z(n6697) );
  CIVX1 U8103 ( .A(n6697), .Z(n6698) );
  CIVX1 U8104 ( .A(n6697), .Z(n6699) );
  CIVX1 U8105 ( .A(n6697), .Z(n6700) );
  CIVX1 U8106 ( .A(n6697), .Z(n6701) );
  CIVX1 U8107 ( .A(n6697), .Z(n6702) );
  CIVX1 U8108 ( .A(n6697), .Z(n6703) );
  CIVX1 U8109 ( .A(n6708), .Z(n6710) );
  CIVX1 U8110 ( .A(n6710), .Z(n6711) );
  CIVX1 U8111 ( .A(n6710), .Z(n6712) );
  CIVX1 U8112 ( .A(n6710), .Z(n6713) );
  CIVX1 U8113 ( .A(n6710), .Z(n6714) );
  CIVX1 U8114 ( .A(n6710), .Z(n6715) );
  CIVX1 U8115 ( .A(n6710), .Z(n6716) );
  CIVX1 U8116 ( .A(n6709), .Z(n6717) );
  CIVX1 U8117 ( .A(n6717), .Z(n6718) );
  CIVX1 U8118 ( .A(n6717), .Z(n6719) );
  CIVX1 U8119 ( .A(n6717), .Z(n6720) );
  CIVX1 U8120 ( .A(n6717), .Z(n6721) );
  CIVX1 U8121 ( .A(n6717), .Z(n6722) );
  CIVX1 U8122 ( .A(n6717), .Z(n6723) );
  CIVX1 U8123 ( .A(n2131), .Z(n6724) );
  CIVX1 U8124 ( .A(n6724), .Z(n6725) );
  CIVX1 U8125 ( .A(n6724), .Z(n6726) );
  CIVX1 U8126 ( .A(n6724), .Z(n6727) );
  CIVX1 U8127 ( .A(n6724), .Z(n6728) );
  CIVX1 U8128 ( .A(n6724), .Z(n6729) );
  CIVX1 U8129 ( .A(n6724), .Z(n6730) );
  CIVX1 U8130 ( .A(n6738), .Z(n6740) );
  CIVX1 U8131 ( .A(n6740), .Z(n6741) );
  CIVX1 U8132 ( .A(n6740), .Z(n6742) );
  CIVX1 U8133 ( .A(n6747), .Z(n6743) );
  CIVX1 U8134 ( .A(n6740), .Z(n6744) );
  CIVX1 U8135 ( .A(n6740), .Z(n6745) );
  CIVX1 U8136 ( .A(n6740), .Z(n6746) );
  CIVX1 U8137 ( .A(n6739), .Z(n6747) );
  CIVX1 U8138 ( .A(n6747), .Z(n6748) );
  CIVX1 U8139 ( .A(n6747), .Z(n6749) );
  CIVX1 U8140 ( .A(n6747), .Z(n6750) );
  CIVX1 U8141 ( .A(n6747), .Z(n6751) );
  CIVX1 U8142 ( .A(n6754), .Z(n6752) );
  CIVX1 U8143 ( .A(n6754), .Z(n6753) );
  CIVX1 U8144 ( .A(n2116), .Z(n6754) );
  CIVX1 U8145 ( .A(n6754), .Z(n6755) );
  CIVX1 U8146 ( .A(n6754), .Z(n6756) );
  CIVX1 U8147 ( .A(n6754), .Z(n6757) );
  CIVX1 U8148 ( .A(n6754), .Z(n6758) );
  CIVX1 U8149 ( .A(n6740), .Z(n6759) );
  CIVX1 U8150 ( .A(n6754), .Z(n6760) );
  CIVX1 U8151 ( .A(n6768), .Z(n6770) );
  CIVX1 U8152 ( .A(n6770), .Z(n6771) );
  CIVX1 U8153 ( .A(n6770), .Z(n6772) );
  CIVX1 U8154 ( .A(n6777), .Z(n6773) );
  CIVX1 U8155 ( .A(n6770), .Z(n6774) );
  CIVX1 U8156 ( .A(n6770), .Z(n6775) );
  CIVX1 U8157 ( .A(n6770), .Z(n6776) );
  CIVX1 U8158 ( .A(n6769), .Z(n6777) );
  CIVX1 U8159 ( .A(n6777), .Z(n6778) );
  CIVX1 U8160 ( .A(n6777), .Z(n6779) );
  CIVX1 U8161 ( .A(n6784), .Z(n6780) );
  CIVX1 U8162 ( .A(n6784), .Z(n6781) );
  CIVX1 U8163 ( .A(n6777), .Z(n6782) );
  CIVX1 U8164 ( .A(n6777), .Z(n6783) );
  CIVX1 U8165 ( .A(n2113), .Z(n6784) );
  CIVX1 U8166 ( .A(n6784), .Z(n6785) );
  CIVX1 U8167 ( .A(n6784), .Z(n6786) );
  CIVX1 U8168 ( .A(n6784), .Z(n6787) );
  CIVX1 U8169 ( .A(n6784), .Z(n6788) );
  CIVX1 U8170 ( .A(n6770), .Z(n6789) );
  CIVX1 U8171 ( .A(n6784), .Z(n6790) );
  CIVX1 U8172 ( .A(n6798), .Z(n6800) );
  CIVX1 U8173 ( .A(n6800), .Z(n6801) );
  CIVX1 U8174 ( .A(n6800), .Z(n6802) );
  CIVX1 U8175 ( .A(n6807), .Z(n6803) );
  CIVX1 U8176 ( .A(n6800), .Z(n6804) );
  CIVX1 U8177 ( .A(n6800), .Z(n6805) );
  CIVX1 U8178 ( .A(n6800), .Z(n6806) );
  CIVX1 U8179 ( .A(n6799), .Z(n6807) );
  CIVX1 U8180 ( .A(n6807), .Z(n6808) );
  CIVX1 U8181 ( .A(n6807), .Z(n6809) );
  CIVX1 U8182 ( .A(n6814), .Z(n6810) );
  CIVX1 U8183 ( .A(n6814), .Z(n6811) );
  CIVX1 U8184 ( .A(n6807), .Z(n6812) );
  CIVX1 U8185 ( .A(n6807), .Z(n6813) );
  CIVX1 U8186 ( .A(n2110), .Z(n6814) );
  CIVX1 U8187 ( .A(n6814), .Z(n6815) );
  CIVX1 U8188 ( .A(n6814), .Z(n6816) );
  CIVX1 U8189 ( .A(n6814), .Z(n6817) );
  CIVX1 U8190 ( .A(n6814), .Z(n6818) );
  CIVX1 U8191 ( .A(n6800), .Z(n6819) );
  CIVX1 U8192 ( .A(n6814), .Z(n6820) );
  CIVX1 U8193 ( .A(n6828), .Z(n6830) );
  CIVX1 U8194 ( .A(n6830), .Z(n6831) );
  CIVX1 U8195 ( .A(n6830), .Z(n6832) );
  CIVX1 U8196 ( .A(n6837), .Z(n6833) );
  CIVX1 U8197 ( .A(n6830), .Z(n6834) );
  CIVX1 U8198 ( .A(n6830), .Z(n6835) );
  CIVX1 U8199 ( .A(n6830), .Z(n6836) );
  CIVX1 U8200 ( .A(n6829), .Z(n6837) );
  CIVX1 U8201 ( .A(n6837), .Z(n6838) );
  CIVX1 U8202 ( .A(n6837), .Z(n6839) );
  CIVX1 U8203 ( .A(n6844), .Z(n6840) );
  CIVX1 U8204 ( .A(n6844), .Z(n6841) );
  CIVX1 U8205 ( .A(n6837), .Z(n6842) );
  CIVX1 U8206 ( .A(n6837), .Z(n6843) );
  CIVX1 U8207 ( .A(n2108), .Z(n6844) );
  CIVX1 U8208 ( .A(n6844), .Z(n6845) );
  CIVX1 U8209 ( .A(n6844), .Z(n6846) );
  CIVX1 U8210 ( .A(n6844), .Z(n6847) );
  CIVX1 U8211 ( .A(n6844), .Z(n6848) );
  CIVX1 U8212 ( .A(n6830), .Z(n6849) );
  CIVX1 U8213 ( .A(n6844), .Z(n6850) );
  CIVX1 U8214 ( .A(n6858), .Z(n6860) );
  CIVX1 U8215 ( .A(n6860), .Z(n6861) );
  CIVX1 U8216 ( .A(n6860), .Z(n6862) );
  CIVX1 U8217 ( .A(n6867), .Z(n6863) );
  CIVX1 U8218 ( .A(n6860), .Z(n6864) );
  CIVX1 U8219 ( .A(n6860), .Z(n6865) );
  CIVX1 U8220 ( .A(n6860), .Z(n6866) );
  CIVX1 U8221 ( .A(n6859), .Z(n6867) );
  CIVX1 U8222 ( .A(n6867), .Z(n6868) );
  CIVX1 U8223 ( .A(n6867), .Z(n6869) );
  CIVX1 U8224 ( .A(n6867), .Z(n6870) );
  CIVX1 U8225 ( .A(n6867), .Z(n6871) );
  CIVX1 U8226 ( .A(n6874), .Z(n6872) );
  CIVX1 U8227 ( .A(n6874), .Z(n6873) );
  CIVX1 U8228 ( .A(n2093), .Z(n6874) );
  CIVX1 U8229 ( .A(n6874), .Z(n6875) );
  CIVX1 U8230 ( .A(n6874), .Z(n6876) );
  CIVX1 U8231 ( .A(n6874), .Z(n6877) );
  CIVX1 U8232 ( .A(n6874), .Z(n6878) );
  CIVX1 U8233 ( .A(n6860), .Z(n6879) );
  CIVX1 U8234 ( .A(n6874), .Z(n6880) );
  CIVX1 U8235 ( .A(n6888), .Z(n6890) );
  CIVX1 U8236 ( .A(n6890), .Z(n6891) );
  CIVX1 U8237 ( .A(n6890), .Z(n6892) );
  CIVX1 U8238 ( .A(n6897), .Z(n6893) );
  CIVX1 U8239 ( .A(n6890), .Z(n6894) );
  CIVX1 U8240 ( .A(n6890), .Z(n6895) );
  CIVX1 U8241 ( .A(n6890), .Z(n6896) );
  CIVX1 U8242 ( .A(n6889), .Z(n6897) );
  CIVX1 U8243 ( .A(n6897), .Z(n6898) );
  CIVX1 U8244 ( .A(n6897), .Z(n6899) );
  CIVX1 U8245 ( .A(n6897), .Z(n6900) );
  CIVX1 U8246 ( .A(n6897), .Z(n6901) );
  CIVX1 U8247 ( .A(n6904), .Z(n6902) );
  CIVX1 U8248 ( .A(n6904), .Z(n6903) );
  CIVX1 U8249 ( .A(n2088), .Z(n6904) );
  CIVX1 U8250 ( .A(n6904), .Z(n6905) );
  CIVX1 U8251 ( .A(n6904), .Z(n6906) );
  CIVX1 U8252 ( .A(n6904), .Z(n6907) );
  CIVX1 U8253 ( .A(n6904), .Z(n6908) );
  CIVX1 U8254 ( .A(n6890), .Z(n6909) );
  CIVX1 U8255 ( .A(n6904), .Z(n6910) );
  CIVX1 U8256 ( .A(n6918), .Z(n6920) );
  CIVX1 U8257 ( .A(n6920), .Z(n6921) );
  CIVX1 U8258 ( .A(n6920), .Z(n6922) );
  CIVX1 U8259 ( .A(n6927), .Z(n6923) );
  CIVX1 U8260 ( .A(n6920), .Z(n6924) );
  CIVX1 U8261 ( .A(n6920), .Z(n6925) );
  CIVX1 U8262 ( .A(n6920), .Z(n6926) );
  CIVX1 U8263 ( .A(n6919), .Z(n6927) );
  CIVX1 U8264 ( .A(n6927), .Z(n6928) );
  CIVX1 U8265 ( .A(n6927), .Z(n6929) );
  CIVX1 U8266 ( .A(n6934), .Z(n6930) );
  CIVX1 U8267 ( .A(n6934), .Z(n6931) );
  CIVX1 U8268 ( .A(n6927), .Z(n6932) );
  CIVX1 U8269 ( .A(n6927), .Z(n6933) );
  CIVX1 U8270 ( .A(n2085), .Z(n6934) );
  CIVX1 U8271 ( .A(n6934), .Z(n6935) );
  CIVX1 U8272 ( .A(n6934), .Z(n6936) );
  CIVX1 U8273 ( .A(n6934), .Z(n6937) );
  CIVX1 U8274 ( .A(n6934), .Z(n6938) );
  CIVX1 U8275 ( .A(n6920), .Z(n6939) );
  CIVX1 U8276 ( .A(n6934), .Z(n6940) );
  CIVX1 U8277 ( .A(n6948), .Z(n6950) );
  CIVX1 U8278 ( .A(n6950), .Z(n6951) );
  CIVX1 U8279 ( .A(n6950), .Z(n6952) );
  CIVX1 U8280 ( .A(n6957), .Z(n6953) );
  CIVX1 U8281 ( .A(n6950), .Z(n6954) );
  CIVX1 U8282 ( .A(n6950), .Z(n6955) );
  CIVX1 U8283 ( .A(n6950), .Z(n6956) );
  CIVX1 U8284 ( .A(n6949), .Z(n6957) );
  CIVX1 U8285 ( .A(n6957), .Z(n6958) );
  CIVX1 U8286 ( .A(n6957), .Z(n6959) );
  CIVX1 U8287 ( .A(n6964), .Z(n6960) );
  CIVX1 U8288 ( .A(n6964), .Z(n6961) );
  CIVX1 U8289 ( .A(n6957), .Z(n6962) );
  CIVX1 U8290 ( .A(n6957), .Z(n6963) );
  CIVX1 U8291 ( .A(n2083), .Z(n6964) );
  CIVX1 U8292 ( .A(n6964), .Z(n6965) );
  CIVX1 U8293 ( .A(n6964), .Z(n6966) );
  CIVX1 U8294 ( .A(n6964), .Z(n6967) );
  CIVX1 U8295 ( .A(n6964), .Z(n6968) );
  CIVX1 U8296 ( .A(n6950), .Z(n6969) );
  CIVX1 U8297 ( .A(n6964), .Z(n6970) );
  CIVX1 U8298 ( .A(n6978), .Z(n6980) );
  CIVX1 U8299 ( .A(n6980), .Z(n6981) );
  CIVX1 U8300 ( .A(n6980), .Z(n6982) );
  CIVX1 U8301 ( .A(n6987), .Z(n6983) );
  CIVX1 U8302 ( .A(n6980), .Z(n6984) );
  CIVX1 U8303 ( .A(n6980), .Z(n6985) );
  CIVX1 U8304 ( .A(n6980), .Z(n6986) );
  CIVX1 U8305 ( .A(n6979), .Z(n6987) );
  CIVX1 U8306 ( .A(n6987), .Z(n6988) );
  CIVX1 U8307 ( .A(n6987), .Z(n6989) );
  CIVX1 U8308 ( .A(n6987), .Z(n6990) );
  CIVX1 U8309 ( .A(n6987), .Z(n6991) );
  CIVX1 U8310 ( .A(n6994), .Z(n6992) );
  CIVX1 U8311 ( .A(n6994), .Z(n6993) );
  CIVX1 U8312 ( .A(n2066), .Z(n6994) );
  CIVX1 U8313 ( .A(n6994), .Z(n6995) );
  CIVX1 U8314 ( .A(n6994), .Z(n6996) );
  CIVX1 U8315 ( .A(n6994), .Z(n6997) );
  CIVX1 U8316 ( .A(n6994), .Z(n6998) );
  CIVX1 U8317 ( .A(n6980), .Z(n6999) );
  CIVX1 U8318 ( .A(n6994), .Z(n7000) );
  CIVX1 U8319 ( .A(n7008), .Z(n7010) );
  CIVX1 U8320 ( .A(n7010), .Z(n7011) );
  CIVX1 U8321 ( .A(n7010), .Z(n7012) );
  CIVX1 U8322 ( .A(n7017), .Z(n7013) );
  CIVX1 U8323 ( .A(n7010), .Z(n7014) );
  CIVX1 U8324 ( .A(n7010), .Z(n7015) );
  CIVX1 U8325 ( .A(n7010), .Z(n7016) );
  CIVX1 U8326 ( .A(n7009), .Z(n7017) );
  CIVX1 U8327 ( .A(n7017), .Z(n7018) );
  CIVX1 U8328 ( .A(n7017), .Z(n7019) );
  CIVX1 U8329 ( .A(n7024), .Z(n7020) );
  CIVX1 U8330 ( .A(n7024), .Z(n7021) );
  CIVX1 U8331 ( .A(n7017), .Z(n7022) );
  CIVX1 U8332 ( .A(n7017), .Z(n7023) );
  CIVX1 U8333 ( .A(n2063), .Z(n7024) );
  CIVX1 U8334 ( .A(n7024), .Z(n7025) );
  CIVX1 U8335 ( .A(n7024), .Z(n7026) );
  CIVX1 U8336 ( .A(n7024), .Z(n7027) );
  CIVX1 U8337 ( .A(n7024), .Z(n7028) );
  CIVX1 U8338 ( .A(n7010), .Z(n7029) );
  CIVX1 U8339 ( .A(n7024), .Z(n7030) );
  CIVX1 U8340 ( .A(n7038), .Z(n7040) );
  CIVX1 U8341 ( .A(n7040), .Z(n7041) );
  CIVX1 U8342 ( .A(n7040), .Z(n7042) );
  CIVX1 U8343 ( .A(n7047), .Z(n7043) );
  CIVX1 U8344 ( .A(n7040), .Z(n7044) );
  CIVX1 U8345 ( .A(n7040), .Z(n7045) );
  CIVX1 U8346 ( .A(n7040), .Z(n7046) );
  CIVX1 U8347 ( .A(n7039), .Z(n7047) );
  CIVX1 U8348 ( .A(n7047), .Z(n7048) );
  CIVX1 U8349 ( .A(n7047), .Z(n7049) );
  CIVX1 U8350 ( .A(n7054), .Z(n7050) );
  CIVX1 U8351 ( .A(n7054), .Z(n7051) );
  CIVX1 U8352 ( .A(n7047), .Z(n7052) );
  CIVX1 U8353 ( .A(n7047), .Z(n7053) );
  CIVX1 U8354 ( .A(n2059), .Z(n7054) );
  CIVX1 U8355 ( .A(n7054), .Z(n7055) );
  CIVX1 U8356 ( .A(n7054), .Z(n7056) );
  CIVX1 U8357 ( .A(n7054), .Z(n7057) );
  CIVX1 U8358 ( .A(n7054), .Z(n7058) );
  CIVX1 U8359 ( .A(n7040), .Z(n7059) );
  CIVX1 U8360 ( .A(n7054), .Z(n7060) );
  CIVX1 U8361 ( .A(n7068), .Z(n7070) );
  CIVX1 U8362 ( .A(n7070), .Z(n7071) );
  CIVX1 U8363 ( .A(n7070), .Z(n7072) );
  CIVX1 U8364 ( .A(n7077), .Z(n7073) );
  CIVX1 U8365 ( .A(n7070), .Z(n7074) );
  CIVX1 U8366 ( .A(n7070), .Z(n7075) );
  CIVX1 U8367 ( .A(n7070), .Z(n7076) );
  CIVX1 U8368 ( .A(n7069), .Z(n7077) );
  CIVX1 U8369 ( .A(n7077), .Z(n7078) );
  CIVX1 U8370 ( .A(n7077), .Z(n7079) );
  CIVX1 U8371 ( .A(n7084), .Z(n7080) );
  CIVX1 U8372 ( .A(n7084), .Z(n7081) );
  CIVX1 U8373 ( .A(n7077), .Z(n7082) );
  CIVX1 U8374 ( .A(n7077), .Z(n7083) );
  CIVX1 U8375 ( .A(n2055), .Z(n7084) );
  CIVX1 U8376 ( .A(n7084), .Z(n7085) );
  CIVX1 U8377 ( .A(n7084), .Z(n7086) );
  CIVX1 U8378 ( .A(n7084), .Z(n7087) );
  CIVX1 U8379 ( .A(n7084), .Z(n7088) );
  CIVX1 U8380 ( .A(n7070), .Z(n7089) );
  CIVX1 U8381 ( .A(n7084), .Z(n7090) );
  CIVXL U8382 ( .A(n4241), .Z(n7113) );
  CIVXL U8383 ( .A(n4241), .Z(n7114) );
  CIVXL U8384 ( .A(n4241), .Z(n7116) );
  CIVXL U8385 ( .A(n4241), .Z(n7117) );
  CIVXL U8386 ( .A(n4241), .Z(n7118) );
  CIVXL U8387 ( .A(n4241), .Z(n7119) );
  CIVXL U8388 ( .A(n4241), .Z(n7120) );
  CIVXL U8389 ( .A(n4241), .Z(n7121) );
  CIVXL U8390 ( .A(n4241), .Z(n7122) );
  CIVXL U8391 ( .A(n4241), .Z(n7123) );
  CIVXL U8392 ( .A(n4242), .Z(n7125) );
  CIVXL U8393 ( .A(n4242), .Z(n7126) );
  CIVXL U8394 ( .A(n4242), .Z(n7127) );
  CIVXL U8395 ( .A(n4242), .Z(n7128) );
  CIVXL U8396 ( .A(n4242), .Z(n7129) );
  CIVXL U8397 ( .A(n4242), .Z(n7130) );
  CIVXL U8398 ( .A(n4242), .Z(n7131) );
  CIVXL U8399 ( .A(n4242), .Z(n7132) );
  CIVXL U8400 ( .A(n4240), .Z(n7150) );
  CIVXL U8401 ( .A(n4240), .Z(n7151) );
  CIVXL U8402 ( .A(n4240), .Z(n7152) );
  CIVXL U8403 ( .A(n4240), .Z(n7153) );
  CIVXL U8404 ( .A(n4240), .Z(n7155) );
  CIVXL U8405 ( .A(n4240), .Z(n7156) );
  CIVXL U8406 ( .A(n4240), .Z(n7158) );
  CEOX1 U8407 ( .A(rd_ptr[8]), .B(\add_121/carry [8]), .Z(N16598) );
  CAN2X1 U8408 ( .A(\add_121/carry [6]), .B(rd_ptr[6]), .Z(\add_121/carry [7])
         );
  CEOX1 U8409 ( .A(rd_ptr[6]), .B(\add_121/carry [6]), .Z(N16596) );
  CAN2X1 U8410 ( .A(\add_121/carry [5]), .B(rd_ptr[5]), .Z(\add_121/carry [6])
         );
  CEOX1 U8411 ( .A(rd_ptr[5]), .B(\add_121/carry [5]), .Z(N16595) );
  CAN2X1 U8412 ( .A(\add_121/carry [4]), .B(rd_ptr[4]), .Z(\add_121/carry [5])
         );
  CEOX1 U8413 ( .A(rd_ptr[4]), .B(\add_121/carry [4]), .Z(N16594) );
  CAN2X1 U8414 ( .A(rd_ptr[0]), .B(n6160), .Z(\add_121/carry [1]) );
  CEOX1 U8415 ( .A(n6160), .B(rd_ptr[0]), .Z(N16590) );
  CEOX1 U8416 ( .A(\add_44/carry [4]), .B(wrt_ptr[4]), .Z(N114) );
  CIVX2 U8417 ( .A(n201), .Z(n7169) );
  CIVX2 U8418 ( .A(n286), .Z(n7170) );
  CIVX2 U8419 ( .A(n8), .Z(n7172) );
  CIVX2 U8420 ( .A(pushin), .Z(n7174) );
  CIVX2 U8421 ( .A(n149), .Z(n7207) );
  CIVX2 U8422 ( .A(n348), .Z(n7209) );
  CIVX2 U8423 ( .A(n6163), .Z(n7210) );
  CIVX2 U8424 ( .A(n10), .Z(n7211) );
  CIVX2 U8425 ( .A(n221), .Z(n7212) );
  CIVX2 U8426 ( .A(n343), .Z(n7215) );
  CIVX2 U8427 ( .A(n6162), .Z(n7216) );
  CIVX2 U8428 ( .A(n6161), .Z(n7217) );
  CIVX2 U8429 ( .A(n178), .Z(n7218) );
  CIVX2 U8430 ( .A(n6160), .Z(n7219) );
  CIVX2 U8431 ( .A(wrt_ptr[0]), .Z(n7220) );
  CIVX2 U8432 ( .A(wrt_ptr[1]), .Z(n7221) );
  CIVX2 U8433 ( .A(wrt_ptr[2]), .Z(n7222) );
  CIVX2 U8434 ( .A(n48), .Z(n7226) );
  CIVX2 U8435 ( .A(n54), .Z(n7227) );
  CIVX2 U8436 ( .A(n17), .Z(n7230) );
  CIVX2 U8437 ( .A(n179), .Z(n7237) );
  CIVX2 U8438 ( .A(n148), .Z(n7240) );
  CIVX2 U8439 ( .A(n307), .Z(n7241) );
  CIVX2 U8440 ( .A(n313), .Z(n7244) );
  CIVX2 U8441 ( .A(n226), .Z(n7245) );
  CIVX2 U8442 ( .A(n889), .Z(n7247) );
  CIVX2 U8443 ( .A(n266), .Z(n7249) );
  CIVX2 U8444 ( .A(n1901), .Z(n7250) );
  CIVX2 U8445 ( .A(n288), .Z(n7252) );
  CIVX2 U8446 ( .A(n355), .Z(n7258) );
  CIVX2 U8447 ( .A(n271), .Z(n7263) );
  CIVX2 U8448 ( .A(n114), .Z(n7265) );
  CIVX2 U8449 ( .A(n159), .Z(n7268) );
  CIVX2 U8450 ( .A(n185), .Z(n7270) );
  CIVX2 U8451 ( .A(n1170), .Z(n7274) );
  CIVX2 U8452 ( .A(n127), .Z(n7277) );
  CIVX2 U8453 ( .A(n1776), .Z(n7279) );
  CIVX2 U8454 ( .A(n509), .Z(n7281) );
  CIVX2 U8455 ( .A(buffer[781]), .Z(n7502) );
  CIVX2 U8456 ( .A(buffer[778]), .Z(n7505) );
  CIVX2 U8457 ( .A(buffer[777]), .Z(n7506) );
  CIVX2 U8458 ( .A(buffer[776]), .Z(n7507) );
  CIVX2 U8459 ( .A(buffer[775]), .Z(n7508) );
  CIVX2 U8460 ( .A(buffer[774]), .Z(n7509) );
  CIVX2 U8461 ( .A(buffer[773]), .Z(n7510) );
  CIVX2 U8462 ( .A(buffer[772]), .Z(n7511) );
  CIVX2 U8463 ( .A(buffer[771]), .Z(n7512) );
  CIVX2 U8464 ( .A(buffer[770]), .Z(n7513) );
  CIVX2 U8465 ( .A(buffer[769]), .Z(n7514) );
  CIVX2 U8466 ( .A(buffer[768]), .Z(n7515) );
  CIVX2 U8467 ( .A(buffer[525]), .Z(n7758) );
  CIVX2 U8468 ( .A(buffer[522]), .Z(n7761) );
  CIVX2 U8469 ( .A(buffer[521]), .Z(n7762) );
  CIVX2 U8470 ( .A(buffer[520]), .Z(n7763) );
  CIVX2 U8471 ( .A(buffer[519]), .Z(n7764) );
  CIVX2 U8472 ( .A(buffer[518]), .Z(n7765) );
  CIVX2 U8473 ( .A(buffer[517]), .Z(n7766) );
  CIVX2 U8474 ( .A(buffer[515]), .Z(n7768) );
  CIVX2 U8475 ( .A(buffer[396]), .Z(n7887) );
  CIVX2 U8476 ( .A(buffer[264]), .Z(n8019) );
  CIVX2 U8477 ( .A(rd_ptr[0]), .Z(n8284) );
  CIVX2 U8478 ( .A(n19), .Z(n8286) );
  CIVX2 U8479 ( .A(rd_ptr[1]), .Z(n8287) );
  CIVX2 U8480 ( .A(rd_ptr[2]), .Z(n8290) );
  CIVX2 U8481 ( .A(rd_ptr[3]), .Z(n8293) );
  CIVX2 U8482 ( .A(n7094), .Z(n8299) );
  CIVX2 U8483 ( .A(n7096), .Z(n8300) );
  CIVX2 U8484 ( .A(rd_ptr[5]), .Z(n8302) );
  CIVX2 U8485 ( .A(n40), .Z(n8307) );
  CIVX2 U8486 ( .A(rd_ptr[6]), .Z(n8308) );
  CIVX2 U8487 ( .A(n942), .Z(n8309) );
endmodule

