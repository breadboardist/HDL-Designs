module();

endmodule
