module FLMultiplier	();

endmodule
