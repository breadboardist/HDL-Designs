
module sqrt64 ( clk, rdy, reset, x, acc );
  input [63:0] x;
  output [31:0] acc;
  input clk, reset;
  output rdy;
  wire   n2689, N130, N131, N132, N133, N134, n297, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688;
  wire   [4:0] bitl;
  wire   [63:0] acc2;

  CFD2QX1 \acc_reg[9]  ( .D(n2666), .CP(clk), .CD(n2613), .Q(acc[9]) );
  CFD2QX1 \acc_reg[25]  ( .D(n2665), .CP(clk), .CD(n2613), .Q(acc[25]) );
  CFD2QX1 \acc_reg[1]  ( .D(n2685), .CP(clk), .CD(n2613), .Q(acc[1]) );
  CFD2QX1 \acc_reg[17]  ( .D(n2664), .CP(clk), .CD(n2613), .Q(acc[17]) );
  CFD2QX1 \acc_reg[23]  ( .D(n2674), .CP(clk), .CD(n2613), .Q(acc[23]) );
  CFD2QX1 \acc_reg[15]  ( .D(n2670), .CP(clk), .CD(n2613), .Q(acc[15]) );
  CFD2QX1 \acc_reg[29]  ( .D(n2677), .CP(clk), .CD(n2613), .Q(acc[29]) );
  CFD2QX1 \acc_reg[21]  ( .D(n2673), .CP(clk), .CD(n2613), .Q(acc[21]) );
  CFD2QX1 \acc_reg[13]  ( .D(n2669), .CP(clk), .CD(n2613), .Q(acc[13]) );
  CFD2QX1 \acc_reg[3]  ( .D(n2684), .CP(clk), .CD(n2613), .Q(acc[3]) );
  CFD2QX1 \acc_reg[27]  ( .D(n2663), .CP(clk), .CD(n2613), .Q(acc[27]) );
  CFD2QX1 \acc_reg[19]  ( .D(n2662), .CP(clk), .CD(n2613), .Q(acc[19]) );
  CFD2QX1 \acc_reg[11]  ( .D(n2661), .CP(clk), .CD(n2613), .Q(acc[11]) );
  CFD2QX1 \acc_reg[6]  ( .D(n2680), .CP(clk), .CD(n2613), .Q(acc[6]) );
  CFD2QX1 \acc_reg[30]  ( .D(n2676), .CP(clk), .CD(n2613), .Q(acc[30]) );
  CFD2QX1 \acc_reg[22]  ( .D(n2672), .CP(clk), .CD(n2613), .Q(acc[22]) );
  CFD2QX1 \acc_reg[14]  ( .D(n2668), .CP(clk), .CD(n2613), .Q(acc[14]) );
  CFD2QX1 \acc_reg[4]  ( .D(n2679), .CP(clk), .CD(n2613), .Q(acc[4]) );
  CFD2QX1 \acc_reg[28]  ( .D(n2675), .CP(clk), .CD(n2613), .Q(acc[28]) );
  CFD2QX1 \acc_reg[20]  ( .D(n2671), .CP(clk), .CD(n2613), .Q(acc[20]) );
  CFD2QX1 \acc_reg[12]  ( .D(n2667), .CP(clk), .CD(n2613), .Q(acc[12]) );
  CFD2QX1 \acc_reg[26]  ( .D(n2660), .CP(clk), .CD(n2613), .Q(acc[26]) );
  CFD2QX1 \acc_reg[18]  ( .D(n2659), .CP(clk), .CD(n2613), .Q(acc[18]) );
  CFD2QX1 \acc_reg[24]  ( .D(n2687), .CP(clk), .CD(n2613), .Q(acc[24]) );
  CFD4QX4 \bitl_reg[4]  ( .D(N133), .CP(clk), .SD(n2613), .Q(bitl[4]) );
  CFD4QX4 \bitl_reg[2]  ( .D(N131), .CP(clk), .SD(n2613), .Q(bitl[2]) );
  CFD4QX4 \bitl_reg[3]  ( .D(N132), .CP(clk), .SD(n2613), .Q(bitl[3]) );
  CFD4QX4 \bitl_reg[0]  ( .D(n452), .CP(clk), .SD(n2613), .Q(bitl[0]) );
  CFD2QX4 \acc_reg[2]  ( .D(n2683), .CP(clk), .CD(n2613), .Q(acc[2]) );
  CFD2QX4 \acc_reg[0]  ( .D(n297), .CP(clk), .CD(n2613), .Q(acc[0]) );
  CFD4QX4 \bitl_reg[1]  ( .D(N130), .CP(clk), .SD(n2613), .Q(bitl[1]) );
  CFD2QX1 \acc_reg[10]  ( .D(n2658), .CP(clk), .CD(n2613), .Q(acc[10]) );
  CFD2QX1 \acc_reg[8]  ( .D(n2688), .CP(clk), .CD(n2613), .Q(acc[8]) );
  CFD2QX1 \acc_reg[5]  ( .D(n2681), .CP(clk), .CD(n2613), .Q(acc[5]) );
  CFD2QX1 \acc_reg[7]  ( .D(n2682), .CP(clk), .CD(n2613), .Q(acc[7]) );
  CFD2XL \acc2_reg[54]  ( .D(n383), .CP(clk), .CD(n2613), .Q(acc2[54]), .QN(
        n2624) );
  CFD2XL \acc2_reg[30]  ( .D(n359), .CP(clk), .CD(n2613), .Q(acc2[30]), .QN(
        n2591) );
  CFD2XL \acc2_reg[37]  ( .D(n366), .CP(clk), .CD(n2613), .Q(acc2[37]), .QN(
        n2598) );
  CFD2XL \acc2_reg[41]  ( .D(n370), .CP(clk), .CD(n2613), .Q(acc2[41]), .QN(
        n2634) );
  CFD2XL \acc2_reg[46]  ( .D(n375), .CP(clk), .CD(n2613), .Q(acc2[46]), .QN(
        n2630) );
  CFD2XL \acc2_reg[33]  ( .D(n362), .CP(clk), .CD(n2613), .Q(acc2[33]), .QN(
        n2609) );
  CFD2XL \acc2_reg[40]  ( .D(n369), .CP(clk), .CD(n2613), .Q(acc2[40]), .QN(
        n2635) );
  CFD2XL \acc2_reg[16]  ( .D(n345), .CP(clk), .CD(n2613), .Q(acc2[16]), .QN(
        n2646) );
  CFD2XL \acc2_reg[49]  ( .D(n378), .CP(clk), .CD(n2613), .Q(acc2[49]), .QN(
        n2602) );
  CFD2XL \acc2_reg[22]  ( .D(n351), .CP(clk), .CD(n2613), .Q(acc2[22]), .QN(
        n2643) );
  CFD2XL \acc2_reg[24]  ( .D(n353), .CP(clk), .CD(n2613), .Q(acc2[24]), .QN(
        n2595) );
  CFD2XL \acc2_reg[15]  ( .D(n344), .CP(clk), .CD(n2613), .Q(acc2[15]), .QN(
        n2647) );
  CFD2XL \acc2_reg[13]  ( .D(n342), .CP(clk), .CD(n2613), .Q(acc2[13]), .QN(
        n2648) );
  CFD2XL \acc2_reg[34]  ( .D(n363), .CP(clk), .CD(n2613), .Q(acc2[34]), .QN(
        n2639) );
  CFD2XL \acc2_reg[10]  ( .D(n339), .CP(clk), .CD(n2613), .Q(acc2[10]), .QN(
        n2650) );
  CFD2XL \acc2_reg[28]  ( .D(n357), .CP(clk), .CD(n2613), .Q(acc2[28]), .QN(
        n2596) );
  CFD2XL \acc2_reg[45]  ( .D(n374), .CP(clk), .CD(n2613), .Q(acc2[45]), .QN(
        n2593) );
  CFD2XL \acc2_reg[58]  ( .D(n387), .CP(clk), .CD(n2613), .Q(acc2[58]), .QN(
        n2620) );
  CFD2XL \acc2_reg[32]  ( .D(n361), .CP(clk), .CD(n2613), .Q(acc2[32]), .QN(
        n2640) );
  CFD2XL \acc2_reg[1]  ( .D(n330), .CP(clk), .CD(n2613), .Q(acc2[1]), .QN(
        n2655) );
  CFD2XL \acc2_reg[19]  ( .D(n348), .CP(clk), .CD(n2613), .Q(acc2[19]), .QN(
        n2608) );
  CFD2XL \acc2_reg[7]  ( .D(n336), .CP(clk), .CD(n2613), .Q(acc2[7]), .QN(
        n2651) );
  CFD2XL \acc2_reg[36]  ( .D(n365), .CP(clk), .CD(n2613), .Q(acc2[36]), .QN(
        n2637) );
  CFD2XL \acc2_reg[20]  ( .D(n349), .CP(clk), .CD(n2613), .Q(acc2[20]), .QN(
        n2594) );
  CFD2XL \acc2_reg[0]  ( .D(n329), .CP(clk), .CD(n2613), .Q(acc2[0]), .QN(
        n2656) );
  CFD2XL \acc2_reg[21]  ( .D(n350), .CP(clk), .CD(n2613), .Q(acc2[21]), .QN(
        n2644) );
  CFD2XL \acc2_reg[31]  ( .D(n360), .CP(clk), .CD(n2613), .Q(acc2[31]), .QN(
        n2600) );
  CFD2XL \acc2_reg[47]  ( .D(n376), .CP(clk), .CD(n2613), .Q(acc2[47]), .QN(
        n2629) );
  CFD2XL \acc2_reg[53]  ( .D(n382), .CP(clk), .CD(n2613), .Q(acc2[53]), .QN(
        n2597) );
  CFD2XL \acc2_reg[4]  ( .D(n333), .CP(clk), .CD(n2613), .Q(acc2[4]), .QN(
        n2610) );
  CFD2XL \acc2_reg[3]  ( .D(n332), .CP(clk), .CD(n2613), .Q(acc2[3]), .QN(
        n2653) );
  CFD2XL \acc2_reg[43]  ( .D(n372), .CP(clk), .CD(n2613), .Q(acc2[43]), .QN(
        n2632) );
  CFD2XL \acc2_reg[55]  ( .D(n384), .CP(clk), .CD(n2613), .Q(acc2[55]), .QN(
        n2623) );
  CFD2XL \acc2_reg[50]  ( .D(n379), .CP(clk), .CD(n2613), .Q(acc2[50]), .QN(
        n2627) );
  CFD2XL \acc2_reg[2]  ( .D(n331), .CP(clk), .CD(n2613), .Q(acc2[2]), .QN(
        n2654) );
  CFD2XL \acc2_reg[5]  ( .D(n334), .CP(clk), .CD(n2613), .Q(acc2[5]), .QN(
        n2605) );
  CFD2XL \acc2_reg[44]  ( .D(n373), .CP(clk), .CD(n2613), .Q(acc2[44]), .QN(
        n2631) );
  CFD2XL \acc2_reg[48]  ( .D(n377), .CP(clk), .CD(n2613), .Q(acc2[48]), .QN(
        n2628) );
  CFD2XL \acc2_reg[57]  ( .D(n386), .CP(clk), .CD(n2613), .Q(acc2[57]), .QN(
        n2621) );
  CFD2XL \acc2_reg[9]  ( .D(n338), .CP(clk), .CD(n2613), .Q(acc2[9]), .QN(
        n2612) );
  CFD2XL \acc2_reg[56]  ( .D(n385), .CP(clk), .CD(n2613), .Q(acc2[56]), .QN(
        n2622) );
  CFD2XL \acc2_reg[59]  ( .D(n388), .CP(clk), .CD(n2613), .Q(acc2[59]), .QN(
        n2619) );
  CFD2XL \acc2_reg[52]  ( .D(n381), .CP(clk), .CD(n2613), .Q(acc2[52]), .QN(
        n2625) );
  CFD2XL \acc2_reg[61]  ( .D(n390), .CP(clk), .CD(n2613), .Q(acc2[61]), .QN(
        n2617) );
  CFD2XL \acc2_reg[60]  ( .D(n389), .CP(clk), .CD(n2613), .Q(acc2[60]), .QN(
        n2618) );
  CFD2XL \acc2_reg[51]  ( .D(n380), .CP(clk), .CD(n2613), .Q(acc2[51]), .QN(
        n2626) );
  CFD2XL \acc2_reg[14]  ( .D(n343), .CP(clk), .CD(n2613), .Q(acc2[14]), .QN(
        n2592) );
  CFD2XL \acc2_reg[62]  ( .D(n391), .CP(clk), .CD(n2613), .Q(acc2[62]), .QN(
        n2616) );
  CFD2XL \acc2_reg[23]  ( .D(n352), .CP(clk), .CD(n2613), .Q(acc2[23]), .QN(
        n2604) );
  CFD2XL \acc2_reg[63]  ( .D(n392), .CP(clk), .CD(n2613), .Q(acc2[63]), .QN(
        n2615) );
  CFD2XL \acc2_reg[11]  ( .D(n340), .CP(clk), .CD(n2613), .Q(acc2[11]), .QN(
        n2649) );
  CFD2XL \acc2_reg[12]  ( .D(n341), .CP(clk), .CD(n2613), .Q(acc2[12]), .QN(
        n2611) );
  CFD2XL \acc2_reg[17]  ( .D(n346), .CP(clk), .CD(n2613), .Q(acc2[17]), .QN(
        n2599) );
  CFD2XL \acc2_reg[25]  ( .D(n354), .CP(clk), .CD(n2613), .Q(acc2[25]), .QN(
        n2607) );
  CFD2XL \acc2_reg[26]  ( .D(n355), .CP(clk), .CD(n2613), .Q(acc2[26]), .QN(
        n2642) );
  CFD2XL \acc2_reg[27]  ( .D(n356), .CP(clk), .CD(n2613), .Q(acc2[27]), .QN(
        n2603) );
  CFD2XL \acc2_reg[38]  ( .D(n367), .CP(clk), .CD(n2613), .Q(acc2[38]), .QN(
        n2636) );
  CFD2XL \acc2_reg[39]  ( .D(n368), .CP(clk), .CD(n2613), .Q(acc2[39]), .QN(
        n2606) );
  CFD2XL \acc2_reg[42]  ( .D(n371), .CP(clk), .CD(n2613), .Q(acc2[42]), .QN(
        n2633) );
  CFD2XL \acc2_reg[8]  ( .D(n337), .CP(clk), .CD(n2613), .Q(acc2[8]), .QN(
        n2601) );
  CFD2XL \acc2_reg[6]  ( .D(n335), .CP(clk), .CD(n2613), .Q(acc2[6]), .QN(
        n2652) );
  CFD2XL \acc2_reg[35]  ( .D(n364), .CP(clk), .CD(n2613), .Q(acc2[35]), .QN(
        n2638) );
  CFD2XL \acc2_reg[18]  ( .D(n347), .CP(clk), .CD(n2613), .Q(acc2[18]), .QN(
        n2645) );
  CFD2XL \acc2_reg[29]  ( .D(n358), .CP(clk), .CD(n2613), .Q(acc2[29]), .QN(
        n2641) );
  CFD2QX2 \acc_reg[16]  ( .D(n2686), .CP(clk), .CD(n2613), .Q(acc[16]) );
  CFD2QX1 \bitl_reg[5]  ( .D(N134), .CP(clk), .CD(n2613), .Q(n2689) );
  CFD2X2 \acc_reg[31]  ( .D(n2678), .CP(clk), .CD(n2613), .Q(acc[31]), .QN(
        n2614) );
  CND2X2 U491 ( .A(n393), .B(n1316), .Z(n1359) );
  CNR2X2 U492 ( .A(n393), .B(n1316), .Z(n1351) );
  CENX2 U493 ( .A(n1308), .B(n1307), .Z(n393) );
  CND2X1 U494 ( .A(n2558), .B(x[40]), .Z(n1550) );
  CND2X2 U495 ( .A(n2067), .B(n2087), .Z(n1401) );
  CND2X2 U496 ( .A(n396), .B(n394), .Z(n1427) );
  CND2X2 U497 ( .A(n1962), .B(n395), .Z(n394) );
  CIVX2 U498 ( .A(n1425), .Z(n395) );
  CND2X2 U499 ( .A(n1426), .B(n1425), .Z(n396) );
  CND2X4 U500 ( .A(n2063), .B(n2449), .Z(n1039) );
  CND4X2 U501 ( .A(n398), .B(n397), .C(n399), .D(n2305), .Z(n2528) );
  CND2X4 U502 ( .A(n2528), .B(x[51]), .Z(n2349) );
  CIVX2 U503 ( .A(n2579), .Z(n2348) );
  CND2X2 U504 ( .A(n400), .B(n2349), .Z(n2354) );
  CND2X2 U505 ( .A(n2299), .B(n2303), .Z(n397) );
  CND3X2 U506 ( .A(n2319), .B(n2302), .C(n2298), .Z(n398) );
  CND2X2 U507 ( .A(n2303), .B(n2304), .Z(n399) );
  CND2X2 U508 ( .A(n2579), .B(x[50]), .Z(n400) );
  CENX2 U509 ( .A(n564), .B(n563), .Z(n2579) );
  CND2X4 U510 ( .A(n402), .B(n401), .Z(n1017) );
  CND2X2 U511 ( .A(n787), .B(acc[6]), .Z(n401) );
  CND2X2 U512 ( .A(n1201), .B(acc[7]), .Z(n402) );
  CIVX2 U513 ( .A(n1332), .Z(n815) );
  CIVX3 U514 ( .A(n403), .Z(n818) );
  CND2X2 U515 ( .A(n1017), .B(n1332), .Z(n403) );
  CND2X4 U516 ( .A(n404), .B(n816), .Z(n1085) );
  CIVX4 U517 ( .A(n1017), .Z(n404) );
  CIVX2 U518 ( .A(n405), .Z(n1903) );
  COND1X2 U519 ( .A(n405), .B(n1900), .C(n1901), .Z(n1885) );
  CND2XL U520 ( .A(n1905), .B(n405), .Z(n1899) );
  CND2X4 U521 ( .A(n1141), .B(n1140), .Z(n405) );
  CND4X4 U522 ( .A(n1090), .B(n1089), .C(n1087), .D(n1088), .Z(n406) );
  CND2X1 U523 ( .A(n406), .B(n2087), .Z(n464) );
  CND2X2 U524 ( .A(n406), .B(n2080), .Z(n1281) );
  CND2X2 U525 ( .A(n406), .B(n1420), .Z(n1095) );
  CNR2X2 U526 ( .A(n2119), .B(n2120), .Z(n2293) );
  CND2X2 U527 ( .A(n408), .B(n407), .Z(n2120) );
  CND2X2 U528 ( .A(n2032), .B(acc2[50]), .Z(n407) );
  CND2X2 U529 ( .A(n2033), .B(n409), .Z(n408) );
  CND2IX1 U530 ( .B(n2032), .A(n410), .Z(n409) );
  CIVX2 U531 ( .A(acc2[50]), .Z(n410) );
  CIVX2 U532 ( .A(n411), .Z(n2117) );
  CNR2X2 U533 ( .A(n2293), .B(n2292), .Z(n2126) );
  CNR2IX2 U534 ( .B(n411), .A(n2118), .Z(n2292) );
  CENX2 U535 ( .A(n2024), .B(n2033), .Z(n2118) );
  CND2X2 U536 ( .A(n2042), .B(acc2[49]), .Z(n411) );
  CND2X2 U537 ( .A(n2030), .B(n2031), .Z(n2042) );
  CIVX3 U538 ( .A(n412), .Z(n414) );
  CND2X4 U539 ( .A(n847), .B(n758), .Z(n412) );
  CND2X4 U540 ( .A(n2053), .B(n2080), .Z(n847) );
  CND2X4 U541 ( .A(n2052), .B(n2449), .Z(n848) );
  CND2X4 U542 ( .A(n415), .B(n413), .Z(n1147) );
  CND2X2 U543 ( .A(n414), .B(n848), .Z(n413) );
  CIVX3 U544 ( .A(n416), .Z(n415) );
  CANR1X2 U545 ( .A(n847), .B(n848), .C(n758), .Z(n416) );
  CNR2X4 U546 ( .A(n1351), .B(n1348), .Z(n1441) );
  CIVDX3 U547 ( .A(n1808), .Z0(n1114), .Z1(n1812) );
  CIVX2 U548 ( .A(n417), .Z(n1467) );
  CND2X2 U549 ( .A(n1434), .B(acc2[41]), .Z(n417) );
  CNR2X4 U550 ( .A(n1464), .B(n1465), .Z(n1544) );
  CENX2 U551 ( .A(n418), .B(n1434), .Z(n1465) );
  CIVX2 U552 ( .A(acc2[41]), .Z(n418) );
  CND2X2 U553 ( .A(n2011), .B(n2087), .Z(n1336) );
  CND2X2 U554 ( .A(n988), .B(n1981), .Z(n708) );
  CNIVX4 U555 ( .A(n1440), .Z(n419) );
  CND2X2 U556 ( .A(n2334), .B(n2355), .Z(n2335) );
  CIVX16 U557 ( .A(n641), .Z(n862) );
  CND2X2 U558 ( .A(n2052), .B(n2080), .Z(n1429) );
  CIVX4 U559 ( .A(n2121), .Z(n2128) );
  COND1X4 U560 ( .A(n1312), .B(n1311), .C(n1310), .Z(n1313) );
  CND2X4 U561 ( .A(n1285), .B(n1284), .Z(n1310) );
  CND2X4 U562 ( .A(n2523), .B(x[62]), .Z(n2180) );
  CND2X2 U563 ( .A(n2083), .B(n2087), .Z(n1409) );
  COND1X2 U564 ( .A(n2293), .B(n2306), .C(n2294), .Z(n2121) );
  CNR2X4 U565 ( .A(n1285), .B(n1284), .Z(n1311) );
  CIVX4 U566 ( .A(n1043), .Z(n1047) );
  CND2X2 U567 ( .A(n1196), .B(n1981), .Z(n778) );
  CIVX4 U568 ( .A(n420), .Z(n1295) );
  CNR2X2 U569 ( .A(n1398), .B(n1288), .Z(n420) );
  CND2X2 U570 ( .A(n1275), .B(n1967), .Z(n1278) );
  CND3X4 U571 ( .A(n1278), .B(n1277), .C(n1276), .Z(n1983) );
  CND2X2 U572 ( .A(n1963), .B(n2087), .Z(n1484) );
  CND3X4 U573 ( .A(n1484), .B(n1483), .C(n1482), .Z(n492) );
  CENX2 U574 ( .A(n662), .B(n1165), .Z(n697) );
  COND1X4 U575 ( .A(n660), .B(n661), .C(n659), .Z(n1165) );
  CND2X1 U576 ( .A(n641), .B(acc[1]), .Z(n716) );
  CNIVX4 U577 ( .A(n2074), .Z(n421) );
  CIVX2 U578 ( .A(n422), .Z(n2123) );
  CND2X2 U579 ( .A(n423), .B(acc2[47]), .Z(n422) );
  CENX2 U580 ( .A(n424), .B(n423), .Z(n1505) );
  CND3X2 U581 ( .A(n1504), .B(n1502), .C(n1503), .Z(n423) );
  CIVX2 U582 ( .A(acc2[47]), .Z(n424) );
  CIVX4 U583 ( .A(n1170), .Z(n1183) );
  CND2X4 U584 ( .A(n2501), .B(acc[30]), .Z(n672) );
  CND4X4 U585 ( .A(n622), .B(n621), .C(n620), .D(n619), .Z(n1061) );
  CIVX8 U586 ( .A(n1061), .Z(n834) );
  CND2X4 U587 ( .A(n1095), .B(n1094), .Z(n1108) );
  CND2X4 U588 ( .A(n2067), .B(n1420), .Z(n954) );
  CND2X4 U589 ( .A(n954), .B(n2601), .Z(n957) );
  CND2X2 U590 ( .A(n464), .B(n425), .Z(n2005) );
  CIVX2 U591 ( .A(n426), .Z(n425) );
  CND2X2 U592 ( .A(n462), .B(n463), .Z(n426) );
  CIVX2 U593 ( .A(n427), .Z(n2154) );
  CND2X2 U594 ( .A(n428), .B(acc2[59]), .Z(n427) );
  CENX2 U595 ( .A(n432), .B(n428), .Z(n2151) );
  CND3X2 U596 ( .A(n2055), .B(n2054), .C(n429), .Z(n428) );
  CND2X2 U597 ( .A(n431), .B(n430), .Z(n429) );
  CIVX2 U598 ( .A(n2056), .Z(n430) );
  CIVX2 U599 ( .A(n2057), .Z(n431) );
  CIVX2 U600 ( .A(acc2[59]), .Z(n432) );
  CND2X2 U601 ( .A(n1193), .B(n1332), .Z(n1194) );
  CIVX4 U602 ( .A(n1018), .Z(n721) );
  COAN1X2 U603 ( .A(n1048), .B(n2070), .C(n1401), .Z(n1403) );
  CIVX4 U604 ( .A(n433), .Z(n1171) );
  CND2X1 U605 ( .A(n629), .B(bitl[1]), .Z(n433) );
  CND3X2 U606 ( .A(n1410), .B(n1409), .C(n1411), .Z(n1434) );
  CENX4 U607 ( .A(n2599), .B(n1034), .Z(n437) );
  CND2X4 U608 ( .A(n1029), .B(n1030), .Z(n1034) );
  CND2X2 U609 ( .A(n991), .B(n1221), .Z(n712) );
  CND3X4 U610 ( .A(n690), .B(n548), .C(n549), .Z(n991) );
  CNIVX1 U611 ( .A(n2292), .Z(n434) );
  CIVX3 U612 ( .A(n1021), .Z(n741) );
  CND2X4 U613 ( .A(n1402), .B(n1403), .Z(n1413) );
  COND1X4 U614 ( .A(acc2[40]), .B(n1413), .C(n1412), .Z(n1406) );
  CND2X4 U615 ( .A(n2273), .B(n2366), .Z(n2356) );
  CND2X4 U616 ( .A(n2576), .B(x[55]), .Z(n2366) );
  CND3X4 U617 ( .A(n945), .B(n944), .C(n946), .Z(n2092) );
  CIVX2 U618 ( .A(n435), .Z(n2000) );
  CND3X2 U619 ( .A(n1999), .B(n2091), .C(n1998), .Z(n435) );
  CNR2IX4 U620 ( .B(n1332), .A(n834), .Z(n700) );
  CNR2IX2 U621 ( .B(acc[10]), .A(n1220), .Z(n767) );
  CNR2X4 U622 ( .A(n1148), .B(n595), .Z(n1867) );
  CND3X4 U623 ( .A(n1996), .B(n1995), .C(n1997), .Z(n1272) );
  CNIVX1 U624 ( .A(n1613), .Z(n436) );
  CND2X4 U625 ( .A(n1201), .B(acc[12]), .Z(n768) );
  CND2X2 U626 ( .A(n1111), .B(n1112), .Z(n1806) );
  CND2X2 U627 ( .A(n1054), .B(n1055), .Z(n1111) );
  CND2X2 U628 ( .A(n1121), .B(n437), .Z(n1653) );
  CAN2X1 U629 ( .A(n1550), .B(n1549), .Z(n534) );
  CND2X2 U630 ( .A(n438), .B(n2355), .Z(n2376) );
  COND1X2 U631 ( .A(n2354), .B(n2353), .C(n2352), .Z(n438) );
  CND2X2 U632 ( .A(n641), .B(acc[27]), .Z(n671) );
  CND2X4 U633 ( .A(n672), .B(n671), .Z(n673) );
  CND4X4 U634 ( .A(n994), .B(n993), .C(n439), .D(n992), .Z(n1989) );
  CND2X2 U635 ( .A(n988), .B(n1332), .Z(n439) );
  CNIVX4 U636 ( .A(n2589), .Z(n440) );
  CND2X4 U637 ( .A(n713), .B(n441), .Z(n1096) );
  CND2X2 U638 ( .A(n2011), .B(n2080), .Z(n441) );
  CND2X2 U639 ( .A(n2475), .B(acc[8]), .Z(n681) );
  CND3X4 U640 ( .A(n683), .B(n682), .C(n681), .Z(n989) );
  CND2X2 U641 ( .A(n442), .B(n1435), .Z(n1391) );
  CND3X2 U642 ( .A(n1388), .B(n1386), .C(n443), .Z(n442) );
  CNR2X2 U643 ( .A(n444), .B(acc2[44]), .Z(n443) );
  CIVX2 U644 ( .A(n1387), .Z(n444) );
  CND2X2 U645 ( .A(n1268), .B(n1267), .Z(n1384) );
  CIVX4 U646 ( .A(n2057), .Z(n445) );
  CND2X2 U647 ( .A(n445), .B(n2449), .Z(n1430) );
  CANR1X2 U648 ( .A(n1346), .B(n1904), .C(n1345), .Z(n1347) );
  CIVX3 U649 ( .A(n2026), .Z(n2056) );
  CND2X1 U650 ( .A(n2026), .B(n1998), .Z(n2437) );
  CNR2IX4 U651 ( .B(bitl[4]), .A(rdy), .Z(n2026) );
  CNIVX3 U652 ( .A(n1840), .Z(n1846) );
  COND1X4 U653 ( .A(n986), .B(n985), .C(n984), .Z(n446) );
  CANR1X4 U654 ( .A(n1752), .B(n1693), .C(n1692), .Z(n986) );
  COND1X2 U655 ( .A(n986), .B(n985), .C(n984), .Z(n1646) );
  CND3X4 U656 ( .A(n744), .B(n743), .C(n742), .Z(n2082) );
  CND2X4 U657 ( .A(n2082), .B(n2449), .Z(n745) );
  CND2X2 U658 ( .A(n2088), .B(n2449), .Z(n802) );
  CNIVX2 U659 ( .A(n2330), .Z(n447) );
  CIVX4 U660 ( .A(n1015), .Z(n819) );
  CIVDX2 U661 ( .A(n1867), .Z0(n1862), .Z1(n1871) );
  CAN2XL U662 ( .A(n1431), .B(acc2[42]), .Z(n1424) );
  CIVX4 U663 ( .A(n536), .Z(n2583) );
  CANR11X2 U664 ( .A(n1997), .B(n1996), .C(n1995), .D(n2056), .Z(n2001) );
  CND2X4 U665 ( .A(n752), .B(n751), .Z(n1142) );
  CND2X2 U666 ( .A(n2209), .B(n2319), .Z(n2214) );
  CAOR1X1 U667 ( .A(n2287), .B(n2319), .C(n2286), .Z(n2288) );
  CNIVX1 U668 ( .A(n2101), .Z(n448) );
  CNR2X4 U669 ( .A(n2000), .B(n2001), .Z(n572) );
  CNR2IX4 U670 ( .B(x[29]), .A(n1929), .Z(n1933) );
  CNR2X1 U671 ( .A(n1492), .B(n1495), .Z(n1493) );
  CND2XL U672 ( .A(n1492), .B(n1491), .Z(n1489) );
  CNIVX1 U673 ( .A(n2555), .Z(n449) );
  CIVDX2 U674 ( .A(n1809), .Z0(n451), .Z1(n450) );
  CND3X4 U675 ( .A(n1109), .B(n1134), .C(n1600), .Z(n1137) );
  CNR2X2 U676 ( .A(n1524), .B(n1523), .Z(n1583) );
  CND2IXL U677 ( .B(n1647), .A(n446), .Z(n1648) );
  CNIVX1 U678 ( .A(n791), .Z(n452) );
  CNIVX1 U679 ( .A(n2614), .Z(n453) );
  CNIVX1 U680 ( .A(n2469), .Z(n454) );
  CND2X2 U681 ( .A(n1110), .B(n455), .Z(n1808) );
  CNR2X2 U682 ( .A(n455), .B(n1110), .Z(n1809) );
  CENX2 U683 ( .A(n1053), .B(n1045), .Z(n455) );
  CIVX3 U684 ( .A(n456), .Z(n1778) );
  CNR2X2 U685 ( .A(n912), .B(n911), .Z(n456) );
  CND2X2 U686 ( .A(n459), .B(n457), .Z(n911) );
  CIVX2 U687 ( .A(n458), .Z(n457) );
  CNR2X2 U688 ( .A(n902), .B(n2610), .Z(n458) );
  CND2X2 U689 ( .A(n904), .B(n903), .Z(n459) );
  CENX2 U690 ( .A(n2605), .B(n917), .Z(n912) );
  CND2X2 U691 ( .A(n908), .B(n907), .Z(n917) );
  CND2X2 U692 ( .A(n551), .B(n550), .Z(n1986) );
  CANR11X2 U693 ( .A(n461), .B(n550), .C(n551), .D(n460), .Z(n2133) );
  CNR2X2 U694 ( .A(n1985), .B(acc2[52]), .Z(n460) );
  CND2X2 U695 ( .A(n1985), .B(acc2[52]), .Z(n461) );
  CND2X2 U696 ( .A(n2133), .B(n2134), .Z(n2275) );
  CENX2 U697 ( .A(n2597), .B(n2005), .Z(n2134) );
  CND2X2 U698 ( .A(n1984), .B(n2091), .Z(n462) );
  CND2X2 U699 ( .A(n1983), .B(n2080), .Z(n463) );
  CND3X2 U700 ( .A(n467), .B(n466), .C(n465), .Z(n469) );
  CND2X2 U701 ( .A(n2590), .B(acc[31]), .Z(n465) );
  CND2X1 U702 ( .A(n787), .B(acc[29]), .Z(n466) );
  CND2X2 U703 ( .A(n1201), .B(acc[30]), .Z(n467) );
  CND2X1 U704 ( .A(n2047), .B(n588), .Z(n1400) );
  CNR2X4 U705 ( .A(n469), .B(n468), .Z(n2047) );
  CNR2X4 U706 ( .A(n2003), .B(n2447), .Z(n468) );
  CIVX2 U707 ( .A(n1031), .Z(n1037) );
  CND2IX2 U708 ( .B(n1031), .A(acc2[16]), .Z(n1033) );
  CND2X2 U709 ( .A(n470), .B(n1036), .Z(n1032) );
  CND2X2 U710 ( .A(n1031), .B(n471), .Z(n470) );
  CIVX2 U711 ( .A(acc2[16]), .Z(n471) );
  CNIVX4 U712 ( .A(n2011), .Z(n472) );
  CND2X4 U713 ( .A(n2011), .B(n478), .Z(n477) );
  CND2X4 U714 ( .A(n712), .B(n711), .Z(n2011) );
  CANR11X2 U715 ( .A(n711), .B(n476), .C(n712), .D(n473), .Z(n480) );
  CIVX2 U716 ( .A(n474), .Z(n473) );
  CND2X2 U717 ( .A(n475), .B(n476), .Z(n474) );
  CIVX2 U718 ( .A(n1420), .Z(n475) );
  CIVX2 U719 ( .A(n481), .Z(n476) );
  CND2X2 U720 ( .A(n472), .B(n1420), .Z(n931) );
  CND2X2 U721 ( .A(n935), .B(n934), .Z(n1741) );
  CND2X2 U722 ( .A(n480), .B(n477), .Z(n934) );
  CIVX2 U723 ( .A(n479), .Z(n478) );
  CND2X2 U724 ( .A(n1420), .B(n481), .Z(n479) );
  CIVX2 U725 ( .A(acc2[7]), .Z(n481) );
  CND2X2 U726 ( .A(n923), .B(n924), .Z(n928) );
  CANR1X2 U727 ( .A(n923), .B(n483), .C(n482), .Z(n935) );
  CNR2X2 U728 ( .A(n927), .B(acc2[6]), .Z(n482) );
  CIVX2 U729 ( .A(n484), .Z(n483) );
  CND2X2 U730 ( .A(n485), .B(n924), .Z(n484) );
  CND2X2 U731 ( .A(n927), .B(acc2[6]), .Z(n485) );
  CIVX2 U732 ( .A(n486), .Z(n2144) );
  CND2X2 U733 ( .A(n487), .B(acc2[55]), .Z(n486) );
  CENX2 U734 ( .A(n488), .B(n487), .Z(n2138) );
  CND2X2 U735 ( .A(n2013), .B(n2014), .Z(n487) );
  CIVX2 U736 ( .A(acc2[55]), .Z(n488) );
  CNR2X4 U737 ( .A(n1488), .B(n1487), .Z(n1972) );
  CENX2 U738 ( .A(n1485), .B(n492), .Z(n1488) );
  CNR2X2 U739 ( .A(n1505), .B(n1506), .Z(n2112) );
  CND2X2 U740 ( .A(n490), .B(n489), .Z(n1506) );
  CND2X2 U741 ( .A(n1500), .B(acc2[46]), .Z(n489) );
  CND2X2 U742 ( .A(n492), .B(n491), .Z(n490) );
  COR2X1 U743 ( .A(acc2[46]), .B(n1500), .Z(n491) );
  CNR2X2 U744 ( .A(n2112), .B(n1972), .Z(n2108) );
  CND2IX1 U745 ( .B(n2566), .A(n1915), .Z(n1916) );
  CENX2 U746 ( .A(n493), .B(n1898), .Z(n2566) );
  CIVX2 U747 ( .A(n1899), .Z(n493) );
  CND3X2 U748 ( .A(n497), .B(n496), .C(n494), .Z(n1368) );
  CIVX2 U749 ( .A(n1370), .Z(n494) );
  CNR2IX2 U750 ( .B(x[37]), .A(n1371), .Z(n1370) );
  CENX2 U751 ( .A(n495), .B(n1357), .Z(n1371) );
  CIVX2 U752 ( .A(n1358), .Z(n495) );
  CIVX2 U753 ( .A(n1372), .Z(n496) );
  CNR2IX2 U754 ( .B(x[38]), .A(n1376), .Z(n1372) );
  CENX2 U755 ( .A(n1326), .B(n1325), .Z(n1376) );
  CIVX2 U756 ( .A(n1377), .Z(n497) );
  CNR2IX2 U757 ( .B(x[39]), .A(n1378), .Z(n1377) );
  CENX2 U758 ( .A(n589), .B(n1347), .Z(n1378) );
  CND2X4 U759 ( .A(n499), .B(n498), .Z(n2124) );
  CND2X2 U760 ( .A(n2044), .B(acc2[48]), .Z(n498) );
  COND1X4 U761 ( .A(acc2[48]), .B(n2044), .C(n2043), .Z(n499) );
  COND1X4 U762 ( .A(n503), .B(n501), .C(n500), .Z(n2044) );
  CND2X1 U763 ( .A(n2040), .B(n2087), .Z(n500) );
  CND3X1 U764 ( .A(n2039), .B(n2038), .C(n502), .Z(n501) );
  CIVX4 U765 ( .A(n2056), .Z(n502) );
  CND2X1 U766 ( .A(n2037), .B(n2036), .Z(n503) );
  CND2X2 U767 ( .A(n505), .B(n504), .Z(n507) );
  CIVX2 U768 ( .A(n508), .Z(n504) );
  CND2X2 U769 ( .A(n2214), .B(n2213), .Z(n505) );
  CND2X4 U770 ( .A(n507), .B(n506), .Z(n2508) );
  CND3X2 U771 ( .A(n2214), .B(n2213), .C(n508), .Z(n506) );
  CIVX4 U772 ( .A(n2215), .Z(n508) );
  CND3X4 U773 ( .A(n2390), .B(n2389), .C(n2388), .Z(n2393) );
  CND2X4 U774 ( .A(n2508), .B(x[59]), .Z(n2388) );
  CIVX2 U775 ( .A(n2565), .Z(n2360) );
  CND2X4 U776 ( .A(n2565), .B(x[53]), .Z(n2358) );
  CENX4 U777 ( .A(n541), .B(n509), .Z(n2565) );
  CND2X4 U778 ( .A(n511), .B(n510), .Z(n509) );
  CIVX1 U779 ( .A(n2280), .Z(n510) );
  CND2X1 U780 ( .A(n2281), .B(n2319), .Z(n511) );
  CND2X2 U781 ( .A(n512), .B(n1826), .Z(n1828) );
  CNR2X2 U782 ( .A(n1822), .B(n1815), .Z(n1826) );
  CNR2IX2 U783 ( .B(x[15]), .A(n2541), .Z(n1822) );
  CND2X2 U784 ( .A(n518), .B(n513), .Z(n512) );
  COND1X2 U785 ( .A(n517), .B(n516), .C(n514), .Z(n513) );
  CNR2X2 U786 ( .A(n1819), .B(n1803), .Z(n514) );
  CNR2IX2 U787 ( .B(x[12]), .A(n2518), .Z(n1803) );
  CENX2 U788 ( .A(n515), .B(n1739), .Z(n2518) );
  CIVX2 U789 ( .A(n1740), .Z(n515) );
  CANR1X2 U790 ( .A(n1718), .B(n1719), .C(n520), .Z(n516) );
  CND2X2 U791 ( .A(n1725), .B(n1724), .Z(n517) );
  CND3X2 U792 ( .A(n1804), .B(n1805), .C(n519), .Z(n518) );
  CNR2X2 U793 ( .A(n1819), .B(n520), .Z(n519) );
  CND2X2 U794 ( .A(n1705), .B(n1722), .Z(n520) );
  CNR2IX2 U795 ( .B(x[13]), .A(n1816), .Z(n1819) );
  CENX2 U796 ( .A(n521), .B(n1732), .Z(n1816) );
  CIVX2 U797 ( .A(n1733), .Z(n521) );
  COND1X1 U798 ( .A(n1476), .B(n1570), .C(n1573), .Z(n1524) );
  CENX2 U799 ( .A(n1475), .B(n1474), .Z(n1570) );
  CIVX2 U800 ( .A(n1477), .Z(n1517) );
  CIVX2 U801 ( .A(n1492), .Z(n1509) );
  COND1X2 U802 ( .A(n523), .B(n1477), .C(n522), .Z(n1492) );
  CIVX2 U803 ( .A(n2109), .Z(n522) );
  CIVX2 U804 ( .A(n1973), .Z(n523) );
  CND2X1 U805 ( .A(n1700), .B(n1698), .Z(n524) );
  CNR2X1 U806 ( .A(n1508), .B(n1972), .Z(n1511) );
  CND2XL U807 ( .A(n1645), .B(n1644), .Z(n525) );
  CND2X1 U808 ( .A(n524), .B(n1697), .Z(n526) );
  CIVX3 U809 ( .A(n2368), .Z(n2576) );
  CND2X2 U810 ( .A(n1960), .B(n2080), .Z(n879) );
  CNR2X2 U811 ( .A(n1855), .B(n1847), .Z(n1849) );
  CND2X2 U812 ( .A(n1841), .B(n1846), .Z(n1855) );
  CEOX2 U813 ( .A(n2599), .B(n1034), .Z(n527) );
  CIVX3 U814 ( .A(n1691), .Z(n973) );
  CND2IX1 U815 ( .B(acc2[14]), .A(n1047), .Z(n1052) );
  CNR2X2 U816 ( .A(n1570), .B(n1476), .Z(n1572) );
  CND2X4 U817 ( .A(n930), .B(n929), .Z(n1742) );
  CAN2X2 U818 ( .A(n1001), .B(n586), .Z(n921) );
  COND1X2 U819 ( .A(n2016), .B(n2015), .C(n2087), .Z(n2023) );
  CNR2IX1 U820 ( .B(acc[23]), .A(n610), .Z(n771) );
  CNR2X2 U821 ( .A(n610), .B(n1227), .Z(n903) );
  CND2X2 U822 ( .A(n2475), .B(acc[13]), .Z(n640) );
  CNR2X4 U823 ( .A(n1852), .B(n1837), .Z(n1156) );
  CIVDX2 U824 ( .A(n1852), .Z0(n1854), .Z1(n1847) );
  CNR2X4 U825 ( .A(n1152), .B(n1151), .Z(n1852) );
  CND2X4 U826 ( .A(n1152), .B(n1151), .Z(n1853) );
  CENX4 U827 ( .A(n873), .B(n872), .Z(n1152) );
  CNR2X2 U828 ( .A(n1169), .B(n1168), .Z(n2029) );
  CNR2X2 U829 ( .A(n2574), .B(x[43]), .Z(n1562) );
  CIVX4 U830 ( .A(n1560), .Z(n2574) );
  CENX2 U831 ( .A(n1539), .B(n1538), .Z(n1560) );
  CANR1X2 U832 ( .A(n1537), .B(n2269), .C(n1536), .Z(n1538) );
  CIVX2 U833 ( .A(n937), .Z(n528) );
  CIVX4 U834 ( .A(n1749), .Z(n937) );
  CND2X2 U835 ( .A(n967), .B(n948), .Z(n529) );
  CND2X2 U836 ( .A(n967), .B(n948), .Z(n1691) );
  CNR2X2 U837 ( .A(n1082), .B(n1982), .Z(n1103) );
  CIVX16 U838 ( .A(n1389), .Z(n1332) );
  CND2IX2 U839 ( .B(n1389), .A(n1180), .Z(n1040) );
  CIVX4 U840 ( .A(n974), .Z(n1698) );
  CEOX1 U841 ( .A(acc2[58]), .B(n2098), .Z(n530) );
  CEOX2 U842 ( .A(n530), .B(n2099), .Z(n2149) );
  CND2X1 U843 ( .A(n2099), .B(n2098), .Z(n531) );
  CND2X1 U844 ( .A(n2099), .B(acc2[58]), .Z(n532) );
  CND2X1 U845 ( .A(n2098), .B(acc2[58]), .Z(n533) );
  CND3X2 U846 ( .A(n531), .B(n532), .C(n533), .Z(n2150) );
  CND3X4 U847 ( .A(n2095), .B(n2094), .C(n2093), .Z(n2099) );
  CNR2X1 U848 ( .A(n608), .B(n2096), .Z(n2098) );
  CND2X2 U849 ( .A(n2151), .B(n2150), .Z(n2206) );
  CNR2X4 U850 ( .A(n2149), .B(n2148), .Z(n2208) );
  CNR2X2 U851 ( .A(n2208), .B(n2205), .Z(n2153) );
  CIVX4 U852 ( .A(n2208), .Z(n2217) );
  CND2X4 U853 ( .A(n979), .B(n978), .Z(n1735) );
  CENX4 U854 ( .A(n942), .B(n941), .Z(n979) );
  CNR2X4 U855 ( .A(n1454), .B(n1442), .Z(n1457) );
  CND3X2 U856 ( .A(n1583), .B(n1559), .C(n534), .Z(n1957) );
  COND1X1 U857 ( .A(n1492), .B(n1490), .C(n1489), .Z(n1499) );
  CANR1X2 U858 ( .A(n1384), .B(n1954), .C(n1383), .Z(n1585) );
  CNIVX2 U859 ( .A(n2327), .Z(n2328) );
  COR2XL U860 ( .A(n1132), .B(n1131), .Z(n535) );
  CND2X2 U861 ( .A(n2393), .B(n2392), .Z(n2394) );
  CND2IX4 U862 ( .B(n782), .A(acc[8]), .Z(n784) );
  CNR2X2 U863 ( .A(n933), .B(n932), .Z(n1744) );
  CNR2X1 U864 ( .A(n2318), .B(n2324), .Z(n579) );
  CENX4 U865 ( .A(n2332), .B(n2331), .Z(n536) );
  COND1X2 U866 ( .A(n2056), .B(n2002), .C(n1273), .Z(n537) );
  COND1X2 U867 ( .A(n2056), .B(n2002), .C(n1273), .Z(n1328) );
  CND2X4 U868 ( .A(n675), .B(n674), .Z(n1426) );
  CND2X2 U869 ( .A(n1034), .B(acc2[17]), .Z(n1118) );
  CND2X1 U870 ( .A(n1222), .B(n1967), .Z(n1223) );
  CND2X1 U871 ( .A(n1222), .B(n1221), .Z(n707) );
  COR2XL U872 ( .A(n2133), .B(n2134), .Z(n538) );
  CNR2X2 U873 ( .A(n1285), .B(n1284), .Z(n539) );
  CIVX3 U874 ( .A(n2405), .Z(n2523) );
  CND2X1 U875 ( .A(n2405), .B(n2404), .Z(n2410) );
  CND2X4 U876 ( .A(n1297), .B(n594), .Z(n902) );
  CANR1X4 U877 ( .A(n914), .B(n1778), .C(n913), .Z(n915) );
  CIVX2 U878 ( .A(n1777), .Z(n913) );
  CIVX2 U879 ( .A(n1782), .Z(n914) );
  CND3X4 U880 ( .A(n1388), .B(n1387), .C(n1386), .Z(n540) );
  CND2X4 U881 ( .A(n2045), .B(n2080), .Z(n1388) );
  CAN2X2 U882 ( .A(n538), .B(n2275), .Z(n541) );
  CIVX4 U883 ( .A(n2407), .Z(n2511) );
  CND2IX1 U884 ( .B(x[63]), .A(n2407), .Z(n2408) );
  CENX4 U885 ( .A(n846), .B(n845), .Z(n1148) );
  CND2X4 U886 ( .A(n1120), .B(n1119), .Z(n1643) );
  CNIVX1 U887 ( .A(n2508), .Z(n542) );
  CANR1X4 U888 ( .A(acc[11]), .B(n2590), .C(n642), .Z(n644) );
  CNR2X4 U889 ( .A(n862), .B(n1425), .Z(n2440) );
  CNR2X4 U890 ( .A(n966), .B(n958), .Z(n959) );
  CND2X4 U891 ( .A(n529), .B(n1707), .Z(n1699) );
  CNR2X2 U892 ( .A(n1834), .B(n1833), .Z(n1835) );
  CENX2 U893 ( .A(n565), .B(n566), .Z(n1829) );
  COND1X2 U894 ( .A(n1672), .B(n1813), .C(n1671), .Z(n565) );
  CND2IX2 U895 ( .B(n819), .A(n1981), .Z(n822) );
  CND2X4 U896 ( .A(n1587), .B(n1656), .Z(n1591) );
  CIVX3 U897 ( .A(n1591), .Z(n1612) );
  CANR1X4 U898 ( .A(n2153), .B(n2219), .C(n2152), .Z(n2183) );
  CENX4 U899 ( .A(n2202), .B(n2201), .Z(n2515) );
  CNR2X4 U900 ( .A(n1514), .B(n1479), .Z(n1973) );
  CANR1X2 U901 ( .A(n1221), .B(n1086), .C(n814), .Z(n824) );
  CND2X2 U902 ( .A(n981), .B(n980), .Z(n1727) );
  CND2X1 U903 ( .A(n2560), .B(n2341), .Z(n2342) );
  CNR2IX2 U904 ( .B(x[49]), .A(n2560), .Z(n2343) );
  CENX4 U905 ( .A(n2641), .B(n874), .Z(n1150) );
  CND2X4 U906 ( .A(n825), .B(n826), .Z(n874) );
  CND2X1 U907 ( .A(n1270), .B(n1221), .Z(n775) );
  CANR1X2 U908 ( .A(acc[21]), .B(n2590), .C(n763), .Z(n766) );
  CND2X2 U909 ( .A(n1084), .B(n1332), .Z(n1090) );
  CND2X1 U910 ( .A(n1201), .B(acc[20]), .Z(n765) );
  COR2X1 U911 ( .A(n905), .B(n1389), .Z(n1092) );
  CND2X2 U912 ( .A(n2522), .B(x[11]), .Z(n1722) );
  CND2X1 U913 ( .A(n1205), .B(n1981), .Z(n868) );
  CND2X1 U914 ( .A(n1175), .B(n1221), .Z(n1089) );
  CND2X2 U915 ( .A(n1086), .B(n1981), .Z(n1087) );
  CNR2X1 U916 ( .A(n1372), .B(n1377), .Z(n1373) );
  COND1X2 U917 ( .A(n1022), .B(n1021), .C(n1221), .Z(n1027) );
  COND1X2 U918 ( .A(n1018), .B(n1017), .C(n1981), .Z(n1019) );
  CND2X1 U919 ( .A(n970), .B(acc2[10]), .Z(n961) );
  CENX1 U920 ( .A(n2051), .B(n2059), .Z(n2155) );
  CND2X2 U921 ( .A(n1196), .B(n1332), .Z(n1076) );
  CND2X1 U922 ( .A(n1196), .B(n1967), .Z(n871) );
  CAN2X1 U923 ( .A(n2555), .B(x[31]), .Z(n1939) );
  CEOX1 U924 ( .A(n1553), .B(n1552), .Z(n1555) );
  CND2X2 U925 ( .A(n1205), .B(n1967), .Z(n1207) );
  CND2X1 U926 ( .A(n1201), .B(acc[18]), .Z(n622) );
  CAN2X1 U927 ( .A(n2020), .B(n2087), .Z(n1204) );
  CND2X2 U928 ( .A(n1193), .B(n1221), .Z(n1041) );
  COND1XL U929 ( .A(n1823), .B(n1822), .C(n1821), .Z(n1824) );
  CIVX16 U930 ( .A(n628), .Z(n1981) );
  CND2X1 U931 ( .A(n864), .B(acc[28]), .Z(n675) );
  CIVX2 U932 ( .A(n827), .Z(n830) );
  CND2X2 U933 ( .A(n1989), .B(n2080), .Z(n1229) );
  CND2X1 U934 ( .A(n1201), .B(acc[6]), .Z(n648) );
  CND2X2 U935 ( .A(n1984), .B(n2080), .Z(n1094) );
  CND2X1 U936 ( .A(n1983), .B(n2449), .Z(n1280) );
  CND2X2 U937 ( .A(n1984), .B(n2087), .Z(n1279) );
  CND2X2 U938 ( .A(n2515), .B(x[61]), .Z(n2398) );
  CNR2XL U939 ( .A(n842), .B(acc2[28]), .Z(n840) );
  CND2XL U940 ( .A(n798), .B(acc2[26]), .Z(n796) );
  CND2X1 U941 ( .A(n1275), .B(n1332), .Z(n811) );
  CND2X1 U942 ( .A(n1989), .B(n2087), .Z(n1993) );
  CND2X1 U943 ( .A(n2010), .B(n2087), .Z(n2014) );
  CNR2IX2 U944 ( .B(n1468), .A(n1469), .Z(n1529) );
  CNR2X1 U945 ( .A(n880), .B(acc2[30]), .Z(n881) );
  CND3X1 U946 ( .A(n1072), .B(n1071), .C(n996), .Z(n997) );
  CND2X1 U947 ( .A(n2088), .B(n2087), .Z(n2095) );
  COR2X1 U948 ( .A(n2029), .B(n2028), .Z(n2030) );
  CND2X2 U949 ( .A(n2010), .B(n2080), .Z(n1338) );
  CND2X1 U950 ( .A(n1413), .B(acc2[40]), .Z(n1405) );
  CNR2XL U951 ( .A(n1303), .B(acc2[36]), .Z(n1300) );
  CIVX2 U952 ( .A(bitl[1]), .Z(n617) );
  CENX2 U953 ( .A(n1012), .B(n2645), .Z(n1014) );
  CND2X1 U954 ( .A(n2269), .B(n2175), .Z(n2176) );
  CND2X1 U955 ( .A(n2059), .B(acc2[60]), .Z(n2060) );
  CND2X1 U956 ( .A(n2077), .B(acc2[56]), .Z(n2078) );
  CIVX3 U957 ( .A(n894), .Z(n895) );
  CND2IX2 U958 ( .B(n1125), .A(n1124), .Z(n1592) );
  COND1X1 U959 ( .A(n1734), .B(n577), .C(n1735), .Z(n1730) );
  CDLY1XL U960 ( .A(n1670), .Z(n1671) );
  CNR2X2 U961 ( .A(n2339), .B(n2335), .Z(n2336) );
  CNR3X2 U962 ( .A(n1956), .B(n1957), .C(n1955), .Z(n2337) );
  CANR1X1 U963 ( .A(n2196), .B(n2195), .C(n2194), .Z(n2197) );
  CND2X2 U964 ( .A(n964), .B(n963), .Z(n965) );
  CNR2X2 U965 ( .A(n895), .B(n896), .Z(n1754) );
  CAN2XL U966 ( .A(n1742), .B(n1741), .Z(n1743) );
  CIVX3 U967 ( .A(n967), .Z(n972) );
  CENX1 U968 ( .A(n2650), .B(n968), .Z(n947) );
  CND2X1 U969 ( .A(n1665), .B(n1813), .Z(n1666) );
  CENX2 U970 ( .A(n1704), .B(n1703), .Z(n2522) );
  CIVX3 U971 ( .A(n1567), .Z(n2562) );
  CENX2 U972 ( .A(n2323), .B(n2322), .Z(n2560) );
  CNR2XL U973 ( .A(n440), .B(n1961), .Z(n2586) );
  CMXI2X2 U974 ( .A0(acc[31]), .A1(acc[30]), .S(n1208), .Z(n543) );
  CNR2IX4 U975 ( .B(n1209), .A(n543), .Z(n1416) );
  CND2X1 U976 ( .A(n1297), .B(n1296), .Z(n1304) );
  CIVX1 U977 ( .A(n1304), .Z(n1298) );
  CAN2X2 U978 ( .A(n917), .B(acc2[5]), .Z(n933) );
  CNR2X1 U979 ( .A(n2237), .B(n2198), .Z(n544) );
  CND2X1 U980 ( .A(n2269), .B(n544), .Z(n2200) );
  CIVX2 U981 ( .A(n1762), .Z(n545) );
  CANR1X4 U982 ( .A(n1764), .B(n1763), .C(n545), .Z(n1756) );
  CIVXL U983 ( .A(n2584), .Z(n546) );
  CMXI2X1 U984 ( .A0(n546), .A1(n2631), .S(n2585), .Z(n373) );
  CANR2XL U985 ( .A(n1964), .B(n2087), .C(n1965), .D(n2485), .Z(n547) );
  CND2X1 U986 ( .A(n1966), .B(n547), .Z(n583) );
  CND2X2 U987 ( .A(n2475), .B(acc[4]), .Z(n548) );
  CND2X2 U988 ( .A(n1201), .B(acc[5]), .Z(n549) );
  CND2X1 U989 ( .A(n2087), .B(n1975), .Z(n550) );
  CANR2X4 U990 ( .A(n1979), .B(n2080), .C(n1978), .D(n1991), .Z(n551) );
  CNR2X1 U991 ( .A(n2237), .B(n2234), .Z(n552) );
  CND2X2 U992 ( .A(n2319), .B(n552), .Z(n2231) );
  CIVX2 U993 ( .A(n1806), .Z(n1113) );
  CIVXL U994 ( .A(n2540), .Z(n553) );
  CMXI2X1 U995 ( .A0(n553), .A1(n2651), .S(n2580), .Z(n336) );
  CIVX2 U996 ( .A(n862), .Z(n554) );
  CANR2X4 U997 ( .A(acc[24]), .B(n1201), .C(acc[22]), .D(n554), .Z(n774) );
  CND3XL U998 ( .A(n1202), .B(n1425), .C(acc[26]), .Z(n1203) );
  CND2IXL U999 ( .B(x[15]), .A(n2541), .Z(n1821) );
  CND2X1 U1000 ( .A(n1967), .B(n990), .Z(n555) );
  CND2X1 U1001 ( .A(n1332), .B(n1331), .Z(n556) );
  CND3X2 U1002 ( .A(n679), .B(n555), .C(n556), .Z(n1958) );
  CND2XL U1003 ( .A(n1961), .B(acc[0]), .Z(n557) );
  CNR2X2 U1004 ( .A(n2589), .B(n557), .Z(n718) );
  CIVXL U1005 ( .A(n940), .Z(n558) );
  CANR5CX4 U1006 ( .A(n941), .B(n2611), .C(n558), .Z(n980) );
  CND2IXL U1007 ( .B(n1253), .A(n1252), .Z(n559) );
  COND3X1 U1008 ( .A(n1362), .B(n1247), .C(n1312), .D(n559), .Z(n1248) );
  CND2X1 U1009 ( .A(n1781), .B(n1780), .Z(n560) );
  CND2X1 U1010 ( .A(n560), .B(n1782), .Z(n561) );
  CND2XL U1011 ( .A(n1777), .B(n1778), .Z(n562) );
  CENX1 U1012 ( .A(n561), .B(n562), .Z(n1790) );
  CANR1X4 U1013 ( .A(n2313), .B(n2319), .C(n2312), .Z(n563) );
  CND2XL U1014 ( .A(n2307), .B(n2306), .Z(n564) );
  CND2IXL U1015 ( .B(n1673), .A(n1674), .Z(n566) );
  CIVXL U1016 ( .A(n2572), .Z(n567) );
  CMXI2X1 U1017 ( .A0(n567), .A1(n2655), .S(n2573), .Z(n330) );
  CND2IXL U1018 ( .B(x[7]), .A(n2540), .Z(n1786) );
  CND4XL U1019 ( .A(n1201), .B(n586), .C(n1425), .D(acc[28]), .Z(n568) );
  CND4XL U1020 ( .A(n586), .B(n1425), .C(n724), .D(acc[29]), .Z(n569) );
  COND3X1 U1021 ( .A(n1961), .B(n1203), .C(n568), .D(n569), .Z(n2019) );
  CENX2 U1022 ( .A(n1931), .B(n1930), .Z(n570) );
  CND2IX2 U1023 ( .B(x[28]), .A(n570), .Z(n1932) );
  CIVXL U1024 ( .A(n2087), .Z(n571) );
  COND1X2 U1025 ( .A(n571), .B(n2002), .C(n572), .Z(n2007) );
  CAOR2X1 U1026 ( .A(n1960), .B(n2091), .C(n1962), .D(n2485), .Z(n573) );
  CANR1XL U1027 ( .A(n1958), .B(n2087), .C(n573), .Z(n574) );
  CENX1 U1028 ( .A(acc2[63]), .B(n574), .Z(n1969) );
  CND2X1 U1029 ( .A(n1072), .B(n1071), .Z(n575) );
  CND2X2 U1030 ( .A(n575), .B(acc2[19]), .Z(n1125) );
  CAN2X4 U1031 ( .A(n1096), .B(acc2[23]), .Z(n1140) );
  CND2X1 U1032 ( .A(n2283), .B(n2278), .Z(n576) );
  COND3X1 U1033 ( .A(n2317), .B(n2279), .C(n2282), .D(n576), .Z(n2280) );
  CIVX4 U1034 ( .A(n526), .Z(n577) );
  CND2XL U1035 ( .A(n1360), .B(n1353), .Z(n578) );
  COND3X1 U1036 ( .A(n1362), .B(n1354), .C(n1359), .D(n578), .Z(n1355) );
  CND2X1 U1037 ( .A(n2319), .B(n579), .Z(n2320) );
  CND2IXL U1038 ( .B(n1754), .A(n1755), .Z(n580) );
  CENX1 U1039 ( .A(n1756), .B(n580), .Z(n593) );
  CIVXL U1040 ( .A(n2541), .Z(n581) );
  CMXI2X1 U1041 ( .A0(n581), .A1(n2647), .S(n2573), .Z(n344) );
  CND2IX1 U1042 ( .B(x[6]), .A(n2563), .Z(n1788) );
  COR2X1 U1043 ( .A(n1220), .B(n2495), .Z(n625) );
  CND2IX1 U1044 ( .B(x[18]), .A(n2534), .Z(n1678) );
  CNR2IX1 U1045 ( .B(n921), .A(n1425), .Z(n919) );
  CNR2X1 U1046 ( .A(n2003), .B(n2096), .Z(n582) );
  CENX1 U1047 ( .A(n582), .B(acc2[62]), .Z(n584) );
  CENX1 U1048 ( .A(n583), .B(n584), .Z(n2159) );
  CANR5CXL U1049 ( .A(n582), .B(acc2[62]), .C(n583), .Z(n585) );
  CIVX1 U1050 ( .A(n585), .Z(n1968) );
  CNR2IX1 U1051 ( .B(n2265), .A(n2261), .Z(n2254) );
  CNR2IX1 U1052 ( .B(n1893), .A(n1890), .Z(n1887) );
  CND2IX1 U1053 ( .B(n1468), .A(n1469), .Z(n1530) );
  CNR2IX1 U1054 ( .B(n1738), .A(n1734), .Z(n1731) );
  CND2IX1 U1055 ( .B(n1972), .A(n2111), .Z(n1491) );
  CND2IX1 U1056 ( .B(n2293), .A(n2294), .Z(n2301) );
  CND2IX1 U1057 ( .B(n1544), .A(n1545), .Z(n1553) );
  COND1XL U1058 ( .A(n587), .B(acc2[0]), .C(n1761), .Z(n600) );
  CIVX8 U1059 ( .A(n636), .Z(n586) );
  CIVX16 U1060 ( .A(n1048), .Z(n1420) );
  CIVX20 U1061 ( .A(n2056), .Z(n2080) );
  CAN2X2 U1062 ( .A(n918), .B(n724), .Z(n587) );
  CIVX4 U1063 ( .A(n641), .Z(n1220) );
  CIVX12 U1064 ( .A(n613), .Z(n1425) );
  CAN2X2 U1065 ( .A(n1332), .B(n1001), .Z(n601) );
  CAN2X2 U1066 ( .A(n607), .B(n1446), .Z(n589) );
  CIVDXL U1067 ( .A(n1885), .Z0(n590), .Z1(n591) );
  CAN2X2 U1068 ( .A(n1302), .B(acc2[37]), .Z(n592) );
  CAN3X2 U1069 ( .A(n886), .B(n1180), .C(n1976), .Z(n594) );
  CAN2X2 U1070 ( .A(n849), .B(acc2[27]), .Z(n595) );
  CNIVX20 U1071 ( .A(n1420), .Z(n2449) );
  CND2X1 U1072 ( .A(n1296), .B(n1990), .Z(n596) );
  CAOR1X1 U1073 ( .A(n1587), .B(n1659), .C(n1586), .Z(n597) );
  CIVDX2 U1074 ( .A(n1865), .Z0(n1845), .Z1(n1870) );
  CIVDX2 U1075 ( .A(n1201), .Z0(n598), .Z1(n599) );
  CIVDX4 U1076 ( .A(n1202), .Z0(n2003), .Z1(n2491) );
  CIVX2 U1077 ( .A(n597), .Z(n602) );
  CAN2X1 U1078 ( .A(n1981), .B(n1420), .Z(n603) );
  COAN1X1 U1079 ( .A(n2234), .B(n2230), .C(n2235), .Z(n604) );
  CAN2X1 U1080 ( .A(n1967), .B(n1420), .Z(n605) );
  CAN2X1 U1081 ( .A(n1496), .B(n1495), .Z(n606) );
  CND3X4 U1082 ( .A(n1174), .B(n1173), .C(n1172), .Z(n1408) );
  CIVX4 U1083 ( .A(n1961), .Z(n1998) );
  CAN2X2 U1084 ( .A(n1862), .B(n1869), .Z(n1863) );
  COR2XL U1085 ( .A(n1439), .B(n1438), .Z(n607) );
  CIVDX4 U1086 ( .A(n599), .Z0(n608), .Z1(n609) );
  CIVX8 U1087 ( .A(n616), .Z(n610) );
  CNR2X4 U1088 ( .A(n2151), .B(n2150), .Z(n2205) );
  CND2X2 U1089 ( .A(n1233), .B(n1200), .Z(n1219) );
  CND2X1 U1090 ( .A(n2007), .B(acc2[54]), .Z(n2008) );
  CND2X4 U1091 ( .A(n844), .B(n843), .Z(n845) );
  CNR2X4 U1092 ( .A(n1130), .B(n1129), .Z(n1617) );
  CNR2IX2 U1093 ( .B(acc[26]), .A(n862), .Z(n863) );
  CND2X4 U1094 ( .A(n1269), .B(n2449), .Z(n1081) );
  CND2X4 U1095 ( .A(n1270), .B(n1967), .Z(n1996) );
  CIVX12 U1096 ( .A(n2422), .Z(n2472) );
  CIVX2 U1097 ( .A(n1291), .Z(n837) );
  CIVX12 U1098 ( .A(n611), .Z(n2590) );
  CIVX2 U1099 ( .A(bitl[0]), .Z(n791) );
  CNIVX12 U1100 ( .A(bitl[4]), .Z(n1980) );
  CIVX8 U1101 ( .A(n1980), .Z(n1180) );
  CNR2X4 U1102 ( .A(bitl[1]), .B(bitl[0]), .Z(n668) );
  CIVX12 U1103 ( .A(bitl[2]), .Z(n613) );
  CND2X4 U1104 ( .A(n2590), .B(n588), .Z(n2589) );
  CNIVX12 U1105 ( .A(bitl[3]), .Z(n1961) );
  CENX1 U1106 ( .A(n1180), .B(n2586), .Z(N133) );
  CNIVX4 U1107 ( .A(n2689), .Z(rdy) );
  CNR2X4 U1108 ( .A(n2689), .B(bitl[4]), .Z(n1001) );
  CIVX8 U1109 ( .A(n1001), .Z(n1048) );
  CMXI2XL U1110 ( .A0(rdy), .A1(n2449), .S(n2586), .Z(n612) );
  CND2X4 U1111 ( .A(rdy), .B(n1980), .Z(n1959) );
  CND2XL U1112 ( .A(n612), .B(n1959), .Z(N134) );
  CNIVX4 U1113 ( .A(n1404), .Z(n2074) );
  CND2X4 U1114 ( .A(bitl[1]), .B(bitl[0]), .Z(n650) );
  CND2XL U1115 ( .A(n421), .B(n2003), .Z(N130) );
  CIVX4 U1116 ( .A(reset), .Z(n2613) );
  CNIVX4 U1117 ( .A(bitl[3]), .Z(n636) );
  CIVDX4 U1118 ( .A(n613), .Z0(n614), .Z1(n588) );
  CIVX4 U1119 ( .A(n614), .Z(n615) );
  CND2X4 U1120 ( .A(n586), .B(n615), .Z(n885) );
  CAN2X4 U1121 ( .A(n1001), .B(n1221), .Z(n2471) );
  CIVX4 U1122 ( .A(bitl[0]), .Z(n629) );
  CAN2X2 U1123 ( .A(n629), .B(bitl[1]), .Z(n616) );
  CNIVX1 U1124 ( .A(n864), .Z(n2484) );
  CND2X1 U1125 ( .A(n2471), .B(n2484), .Z(n2424) );
  CIVX2 U1126 ( .A(n629), .Z(n618) );
  CND2X4 U1127 ( .A(n618), .B(n617), .Z(n782) );
  CIVX16 U1128 ( .A(n782), .Z(n1201) );
  CND2X1 U1129 ( .A(n2590), .B(acc[19]), .Z(n621) );
  CIVX8 U1130 ( .A(n650), .Z(n641) );
  CIVX2 U1131 ( .A(acc[16]), .Z(n2469) );
  COR2X2 U1132 ( .A(n862), .B(n2469), .Z(n620) );
  CND2X1 U1133 ( .A(n1171), .B(acc[17]), .Z(n619) );
  CND2X4 U1134 ( .A(n1961), .B(n1425), .Z(n1290) );
  CIVX8 U1135 ( .A(n1290), .Z(n1967) );
  CND2X1 U1136 ( .A(n834), .B(n1967), .Z(n2039) );
  CAN2X2 U1137 ( .A(n1201), .B(acc[22]), .Z(n627) );
  CIVX2 U1138 ( .A(acc[20]), .Z(n2495) );
  CND2X1 U1139 ( .A(n2590), .B(acc[23]), .Z(n624) );
  CND2X1 U1140 ( .A(n1171), .B(acc[21]), .Z(n623) );
  CND3X2 U1141 ( .A(n625), .B(n624), .C(n623), .Z(n626) );
  CNR2X4 U1142 ( .A(n626), .B(n627), .Z(n1291) );
  CND2X4 U1143 ( .A(n613), .B(n1961), .Z(n628) );
  CND2X1 U1144 ( .A(n1291), .B(n1981), .Z(n2037) );
  CND2X2 U1145 ( .A(n2039), .B(n2037), .Z(n661) );
  CAN2X4 U1146 ( .A(n629), .B(bitl[1]), .Z(n787) );
  CIVX2 U1147 ( .A(acc[28]), .Z(n2447) );
  CIVX12 U1148 ( .A(n885), .Z(n1221) );
  CND2X2 U1149 ( .A(n2047), .B(n1221), .Z(n2038) );
  CND2X1 U1150 ( .A(n1201), .B(acc[26]), .Z(n631) );
  CND2X1 U1151 ( .A(n1202), .B(acc[24]), .Z(n630) );
  CND2X2 U1152 ( .A(n631), .B(n630), .Z(n635) );
  CND2X1 U1153 ( .A(n2590), .B(acc[27]), .Z(n633) );
  CND2X1 U1154 ( .A(n1171), .B(acc[25]), .Z(n632) );
  CND2X2 U1155 ( .A(n633), .B(n632), .Z(n634) );
  CNR2X4 U1156 ( .A(n635), .B(n634), .Z(n1398) );
  CND2X4 U1157 ( .A(n586), .B(n1425), .Z(n1389) );
  CND2X1 U1158 ( .A(n1398), .B(n1332), .Z(n2036) );
  CND3X2 U1159 ( .A(n2036), .B(n2038), .C(n2449), .Z(n660) );
  CIVX8 U1160 ( .A(n610), .Z(n2475) );
  CND2X1 U1161 ( .A(n1201), .B(acc[14]), .Z(n639) );
  CNR2IX2 U1162 ( .B(acc[12]), .A(n862), .Z(n637) );
  CANR1X4 U1163 ( .A(acc[15]), .B(n2590), .C(n637), .Z(n638) );
  CND3X4 U1164 ( .A(n639), .B(n640), .C(n638), .Z(n1058) );
  CND2X2 U1165 ( .A(n1058), .B(n1221), .Z(n658) );
  CND2X1 U1166 ( .A(n1201), .B(acc[10]), .Z(n645) );
  CNR2IX2 U1167 ( .B(acc[8]), .A(n862), .Z(n642) );
  CND2X1 U1168 ( .A(n1171), .B(acc[9]), .Z(n643) );
  CND3X4 U1169 ( .A(n645), .B(n644), .C(n643), .Z(n1063) );
  CND2X4 U1170 ( .A(n1063), .B(n1332), .Z(n657) );
  CNR2IX2 U1171 ( .B(acc[4]), .A(n862), .Z(n646) );
  CANR1X2 U1172 ( .A(acc[7]), .B(n2590), .C(n646), .Z(n649) );
  CND2X1 U1173 ( .A(n1171), .B(acc[5]), .Z(n647) );
  CND3X4 U1174 ( .A(n649), .B(n648), .C(n647), .Z(n1062) );
  CND2X2 U1175 ( .A(n1062), .B(n1981), .Z(n656) );
  CND2X1 U1176 ( .A(n1171), .B(acc[1]), .Z(n652) );
  CIVX4 U1177 ( .A(n650), .Z(n1202) );
  CND2X1 U1178 ( .A(n1202), .B(acc[0]), .Z(n651) );
  CND2X2 U1179 ( .A(n652), .B(n651), .Z(n828) );
  CND2X2 U1180 ( .A(n1201), .B(acc[2]), .Z(n654) );
  CND2X2 U1181 ( .A(n2590), .B(acc[3]), .Z(n653) );
  CND2X4 U1182 ( .A(n654), .B(n653), .Z(n827) );
  COND1X2 U1183 ( .A(n828), .B(n827), .C(n1967), .Z(n655) );
  CND4X4 U1184 ( .A(n658), .B(n656), .C(n657), .D(n655), .Z(n2040) );
  CND2X2 U1185 ( .A(n2040), .B(n2080), .Z(n659) );
  CND2X4 U1186 ( .A(n1221), .B(n1980), .Z(n1977) );
  CNR2X4 U1187 ( .A(n1977), .B(n421), .Z(n1164) );
  CENX2 U1188 ( .A(acc2[32]), .B(n1164), .Z(n662) );
  CIVDX3 U1189 ( .A(n668), .Z0(n611), .Z1(n724) );
  CND2X1 U1190 ( .A(n2501), .B(acc[18]), .Z(n664) );
  CND2X1 U1191 ( .A(acc[15]), .B(n1202), .Z(n663) );
  CAN2X2 U1192 ( .A(n664), .B(n663), .Z(n667) );
  CND2X1 U1193 ( .A(n1201), .B(acc[17]), .Z(n666) );
  CND2X1 U1194 ( .A(n1171), .B(acc[16]), .Z(n665) );
  CND3X4 U1195 ( .A(n667), .B(n666), .C(n665), .Z(n990) );
  CANR2X2 U1196 ( .A(n2475), .B(acc[24]), .C(acc[23]), .D(n1202), .Z(n670) );
  CIVDX2 U1197 ( .A(n668), .Z0(n1404), .Z1(n2501) );
  CANR2X1 U1198 ( .A(n1201), .B(acc[25]), .C(n724), .D(acc[26]), .Z(n669) );
  CND2X2 U1199 ( .A(n670), .B(n669), .Z(n1331) );
  CANR1X2 U1200 ( .A(acc[29]), .B(n1201), .C(n673), .Z(n674) );
  CND2X2 U1201 ( .A(n2475), .B(acc[20]), .Z(n678) );
  CANR2X2 U1202 ( .A(n724), .B(acc[22]), .C(acc[19]), .D(n1202), .Z(n677) );
  CND2X2 U1203 ( .A(n1201), .B(acc[21]), .Z(n676) );
  CND3X4 U1204 ( .A(n678), .B(n677), .C(n676), .Z(n1222) );
  CANR2X2 U1205 ( .A(n1426), .B(n1221), .C(n1981), .D(n1222), .Z(n679) );
  CND2X2 U1206 ( .A(n1958), .B(n1420), .Z(n878) );
  CND2X1 U1207 ( .A(n1201), .B(acc[9]), .Z(n683) );
  CIVX2 U1208 ( .A(acc[7]), .Z(n2492) );
  CIVX2 U1209 ( .A(acc[10]), .Z(n2477) );
  COND2X1 U1210 ( .A(n1220), .B(n2492), .C(n2477), .D(n1404), .Z(n680) );
  CIVX2 U1211 ( .A(n680), .Z(n682) );
  CND2X2 U1212 ( .A(n989), .B(n1332), .Z(n694) );
  CANR2X2 U1213 ( .A(n724), .B(acc[14]), .C(acc[11]), .D(n1202), .Z(n686) );
  CND2X2 U1214 ( .A(n1201), .B(acc[13]), .Z(n685) );
  CND2X1 U1215 ( .A(n787), .B(acc[12]), .Z(n684) );
  CND3X2 U1216 ( .A(n686), .B(n685), .C(n684), .Z(n988) );
  CND2X2 U1217 ( .A(n988), .B(n1221), .Z(n693) );
  CND2X2 U1218 ( .A(n1201), .B(acc[1]), .Z(n689) );
  CND2X2 U1219 ( .A(n787), .B(acc[0]), .Z(n688) );
  CND2X2 U1220 ( .A(n2590), .B(acc[2]), .Z(n687) );
  CND3X4 U1221 ( .A(n689), .B(n688), .C(n687), .Z(n987) );
  CND2X2 U1222 ( .A(n987), .B(n1967), .Z(n692) );
  CANR2X2 U1223 ( .A(n2590), .B(acc[6]), .C(acc[3]), .D(n1202), .Z(n690) );
  CND2X2 U1224 ( .A(n991), .B(n1981), .Z(n691) );
  CND4X4 U1225 ( .A(n694), .B(n693), .C(n692), .D(n691), .Z(n1960) );
  CND2X2 U1226 ( .A(n878), .B(n879), .Z(n695) );
  CND2X2 U1227 ( .A(n695), .B(acc2[31]), .Z(n696) );
  CIVX2 U1228 ( .A(n696), .Z(n698) );
  CNR2X2 U1229 ( .A(n697), .B(n698), .Z(n1238) );
  CIVXL U1230 ( .A(n1238), .Z(n1185) );
  CND2X2 U1231 ( .A(n698), .B(n697), .Z(n1244) );
  CND2X1 U1232 ( .A(n1185), .B(n1244), .Z(n1163) );
  COR2X2 U1233 ( .A(n1980), .B(n1290), .Z(n1385) );
  CNR2X1 U1234 ( .A(n1385), .B(n421), .Z(n749) );
  CENX2 U1235 ( .A(acc2[24]), .B(n749), .Z(n706) );
  CNR2IX2 U1236 ( .B(n1221), .A(n1291), .Z(n699) );
  CNR2X4 U1237 ( .A(n700), .B(n699), .Z(n702) );
  CANR2X2 U1238 ( .A(n1063), .B(n1967), .C(n1981), .D(n1058), .Z(n701) );
  CND2X4 U1239 ( .A(n702), .B(n701), .Z(n2069) );
  CND2X4 U1240 ( .A(n2069), .B(n2449), .Z(n748) );
  CND2X2 U1241 ( .A(n1062), .B(n1221), .Z(n704) );
  COND1X2 U1242 ( .A(n828), .B(n827), .C(n1332), .Z(n703) );
  CND2X4 U1243 ( .A(n704), .B(n703), .Z(n2067) );
  CND2X2 U1244 ( .A(n2067), .B(n2080), .Z(n705) );
  CND2X4 U1245 ( .A(n748), .B(n705), .Z(n747) );
  CENX4 U1246 ( .A(n706), .B(n747), .Z(n1141) );
  CND2X1 U1247 ( .A(n990), .B(n1332), .Z(n710) );
  CND2X2 U1248 ( .A(n989), .B(n1967), .Z(n709) );
  CND4X4 U1249 ( .A(n710), .B(n708), .C(n709), .D(n707), .Z(n2010) );
  CND2X2 U1250 ( .A(n2010), .B(n1420), .Z(n713) );
  CND2X4 U1251 ( .A(n987), .B(n1332), .Z(n711) );
  CNR2X2 U1252 ( .A(n1141), .B(n1140), .Z(n1897) );
  CND2X2 U1253 ( .A(n1201), .B(acc[3]), .Z(n715) );
  CND2X1 U1254 ( .A(n787), .B(acc[2]), .Z(n714) );
  CND2X4 U1255 ( .A(n714), .B(n715), .Z(n1015) );
  CND2X2 U1256 ( .A(n2590), .B(acc[4]), .Z(n717) );
  CIVX2 U1257 ( .A(acc[1]), .Z(n2473) );
  CND2X4 U1258 ( .A(n717), .B(n716), .Z(n1016) );
  CIVX4 U1259 ( .A(n1016), .Z(n820) );
  CND2X4 U1260 ( .A(n819), .B(n820), .Z(n1091) );
  CANR1X4 U1261 ( .A(n1332), .B(n1091), .C(n718), .Z(n723) );
  CND2X2 U1262 ( .A(n2590), .B(acc[8]), .Z(n720) );
  CND2X1 U1263 ( .A(n1202), .B(acc[5]), .Z(n719) );
  CND2X4 U1264 ( .A(n720), .B(n719), .Z(n1018) );
  CND2X2 U1265 ( .A(n1085), .B(n1221), .Z(n722) );
  CND2X4 U1266 ( .A(n723), .B(n722), .Z(n2083) );
  CND2X2 U1267 ( .A(n2083), .B(n2080), .Z(n746) );
  CANR2X1 U1268 ( .A(n1202), .B(acc[21]), .C(acc[24]), .D(n2501), .Z(n727) );
  CND2X2 U1269 ( .A(n864), .B(acc[22]), .Z(n726) );
  CND2X1 U1270 ( .A(n1201), .B(acc[23]), .Z(n725) );
  CND3X2 U1271 ( .A(n727), .B(n726), .C(n725), .Z(n1275) );
  CANR2X2 U1272 ( .A(n2590), .B(acc[20]), .C(acc[17]), .D(n1202), .Z(n730) );
  CND2X1 U1273 ( .A(n1171), .B(acc[18]), .Z(n729) );
  CND2X2 U1274 ( .A(n1201), .B(acc[19]), .Z(n728) );
  CND3X4 U1275 ( .A(n730), .B(n729), .C(n728), .Z(n1175) );
  CANR2X2 U1276 ( .A(n1275), .B(n1221), .C(n1332), .D(n1175), .Z(n744) );
  CND2X4 U1277 ( .A(n1201), .B(acc[11]), .Z(n732) );
  CND2X2 U1278 ( .A(n787), .B(acc[10]), .Z(n731) );
  CND2X4 U1279 ( .A(n732), .B(n731), .Z(n1025) );
  CIVX4 U1280 ( .A(n1025), .Z(n736) );
  CND2X4 U1281 ( .A(n2590), .B(acc[12]), .Z(n733) );
  CIVX4 U1282 ( .A(n733), .Z(n735) );
  CIVX2 U1283 ( .A(acc[9]), .Z(n2460) );
  CNR2X1 U1284 ( .A(n1220), .B(n2460), .Z(n734) );
  CNR2X4 U1285 ( .A(n735), .B(n734), .Z(n1023) );
  CND2X4 U1286 ( .A(n736), .B(n1023), .Z(n1086) );
  CND2X1 U1287 ( .A(n1086), .B(n1967), .Z(n743) );
  CND2X2 U1288 ( .A(n1201), .B(acc[15]), .Z(n738) );
  CND2X2 U1289 ( .A(n2475), .B(acc[14]), .Z(n737) );
  CND2X2 U1290 ( .A(n738), .B(n737), .Z(n1021) );
  CIVX2 U1291 ( .A(acc[13]), .Z(n2443) );
  CND2X2 U1292 ( .A(n2590), .B(acc[16]), .Z(n739) );
  COND1X4 U1293 ( .A(n2443), .B(n2003), .C(n739), .Z(n1022) );
  CIVX2 U1294 ( .A(n1022), .Z(n740) );
  CND2X4 U1295 ( .A(n741), .B(n740), .Z(n1084) );
  CND2X2 U1296 ( .A(n1084), .B(n1981), .Z(n742) );
  CND2X4 U1297 ( .A(n745), .B(n746), .Z(n806) );
  CENX2 U1298 ( .A(n2607), .B(n806), .Z(n1143) );
  CND2X2 U1299 ( .A(n747), .B(acc2[24]), .Z(n752) );
  CND2X1 U1300 ( .A(n2595), .B(n748), .Z(n750) );
  CND2X2 U1301 ( .A(n750), .B(n749), .Z(n751) );
  CNR2X4 U1302 ( .A(n1143), .B(n1142), .Z(n1900) );
  CNR2X2 U1303 ( .A(n1897), .B(n1900), .Z(n1893) );
  CND2X1 U1304 ( .A(n989), .B(n1221), .Z(n754) );
  CANR2X2 U1305 ( .A(n991), .B(n1332), .C(n1981), .D(n987), .Z(n753) );
  CND2X2 U1306 ( .A(n754), .B(n753), .Z(n2053) );
  CANR2X2 U1307 ( .A(n1967), .B(n988), .C(n1981), .D(n990), .Z(n757) );
  CND2X1 U1308 ( .A(n1222), .B(n1332), .Z(n756) );
  CND2X1 U1309 ( .A(n1331), .B(n1221), .Z(n755) );
  CND3X4 U1310 ( .A(n757), .B(n756), .C(n755), .Z(n2052) );
  CIVX2 U1311 ( .A(n2603), .Z(n758) );
  CNR2IX2 U1312 ( .B(acc[14]), .A(n862), .Z(n759) );
  CANR1X2 U1313 ( .A(acc[17]), .B(n2590), .C(n759), .Z(n762) );
  CND2IX1 U1314 ( .B(n2469), .A(n1201), .Z(n761) );
  CND2X1 U1315 ( .A(n787), .B(acc[15]), .Z(n760) );
  CND3X4 U1316 ( .A(n762), .B(n761), .C(n760), .Z(n1196) );
  CNR2IX2 U1317 ( .B(acc[18]), .A(n862), .Z(n763) );
  CND2X1 U1318 ( .A(n1171), .B(acc[19]), .Z(n764) );
  CND3X4 U1319 ( .A(n766), .B(n765), .C(n764), .Z(n1205) );
  CND2X1 U1320 ( .A(n1205), .B(n1332), .Z(n777) );
  CANR2X4 U1321 ( .A(n2590), .B(acc[13]), .C(acc[11]), .D(n787), .Z(n770) );
  CIVX2 U1322 ( .A(n767), .Z(n769) );
  CND3X4 U1323 ( .A(n770), .B(n768), .C(n769), .Z(n1193) );
  CND2X1 U1324 ( .A(n1193), .B(n1967), .Z(n776) );
  CIVX2 U1325 ( .A(n771), .Z(n773) );
  CND2X1 U1326 ( .A(n2590), .B(acc[25]), .Z(n772) );
  CND3X4 U1327 ( .A(n774), .B(n773), .C(n772), .Z(n1270) );
  CND4X4 U1328 ( .A(n775), .B(n778), .C(n777), .D(n776), .Z(n2088) );
  CND2X4 U1329 ( .A(n1171), .B(acc[7]), .Z(n779) );
  CIVX4 U1330 ( .A(n779), .Z(n781) );
  CNR2IX2 U1331 ( .B(acc[6]), .A(n1220), .Z(n780) );
  CNR2X4 U1332 ( .A(n781), .B(n780), .Z(n785) );
  CND2X2 U1333 ( .A(n2590), .B(acc[9]), .Z(n783) );
  CND3X4 U1334 ( .A(n785), .B(n784), .C(n783), .Z(n1192) );
  CND2X2 U1335 ( .A(n1192), .B(n1221), .Z(n945) );
  CND2X2 U1336 ( .A(n1201), .B(acc[4]), .Z(n790) );
  CNR2IX4 U1337 ( .B(acc[2]), .A(n862), .Z(n786) );
  CANR1X4 U1338 ( .A(acc[5]), .B(n2590), .C(n786), .Z(n789) );
  CND2X1 U1339 ( .A(n787), .B(acc[3]), .Z(n788) );
  CND3X4 U1340 ( .A(n789), .B(n790), .C(n788), .Z(n1197) );
  CND2X2 U1341 ( .A(n1197), .B(n1332), .Z(n944) );
  CIVX3 U1342 ( .A(n791), .Z(n1208) );
  CMXI2X1 U1343 ( .A0(acc[1]), .A1(acc[0]), .S(n1208), .Z(n792) );
  CNIVX1 U1344 ( .A(bitl[1]), .Z(n1209) );
  CNR2X2 U1345 ( .A(n792), .B(n1209), .Z(n920) );
  CND2X2 U1346 ( .A(n920), .B(n588), .Z(n1006) );
  CIVX3 U1347 ( .A(n1006), .Z(n793) );
  CND2X4 U1348 ( .A(n793), .B(n1961), .Z(n946) );
  CND2X2 U1349 ( .A(n2092), .B(n2080), .Z(n801) );
  CND2X2 U1350 ( .A(n802), .B(n801), .Z(n795) );
  CNR2X2 U1351 ( .A(n1385), .B(n598), .Z(n798) );
  COR2X1 U1352 ( .A(acc2[26]), .B(n798), .Z(n794) );
  CND2X2 U1353 ( .A(n795), .B(n794), .Z(n797) );
  CND2X2 U1354 ( .A(n797), .B(n796), .Z(n1146) );
  CNR2X4 U1355 ( .A(n1147), .B(n1146), .Z(n1882) );
  CENX1 U1356 ( .A(acc2[26]), .B(n798), .Z(n799) );
  CND2IX2 U1357 ( .B(n802), .A(n799), .Z(n805) );
  CND2IX2 U1358 ( .B(n801), .A(n799), .Z(n804) );
  CIVX2 U1359 ( .A(n799), .Z(n800) );
  CND3X2 U1360 ( .A(n802), .B(n801), .C(n800), .Z(n803) );
  CND3X4 U1361 ( .A(n805), .B(n804), .C(n803), .Z(n1144) );
  CND2X2 U1362 ( .A(n806), .B(acc2[25]), .Z(n807) );
  CIVX3 U1363 ( .A(n807), .Z(n1145) );
  CNR2X4 U1364 ( .A(n1144), .B(n1145), .Z(n1890) );
  CNR2X2 U1365 ( .A(n1882), .B(n1890), .Z(n1843) );
  CND2X2 U1366 ( .A(n1893), .B(n1843), .Z(n1864) );
  CANR2X2 U1367 ( .A(n2590), .B(acc[28]), .C(acc[25]), .D(n1202), .Z(n810) );
  CND2X1 U1368 ( .A(n1171), .B(acc[26]), .Z(n809) );
  CND2X4 U1369 ( .A(n1201), .B(acc[27]), .Z(n808) );
  CND3X4 U1370 ( .A(n810), .B(n809), .C(n808), .Z(n1407) );
  CANR2X2 U1371 ( .A(n1175), .B(n1981), .C(n1221), .D(n1407), .Z(n813) );
  CND2X2 U1372 ( .A(n1084), .B(n1967), .Z(n812) );
  CND3X4 U1373 ( .A(n813), .B(n812), .C(n811), .Z(n2062) );
  CND2X2 U1374 ( .A(n2062), .B(n2449), .Z(n826) );
  CND2X2 U1375 ( .A(n2590), .B(acc[0]), .Z(n905) );
  CNR2X1 U1376 ( .A(n905), .B(n1290), .Z(n814) );
  CIVX2 U1377 ( .A(n1018), .Z(n816) );
  CNR2X2 U1378 ( .A(n721), .B(n815), .Z(n817) );
  CNR2X4 U1379 ( .A(n817), .B(n818), .Z(n823) );
  CND2IX2 U1380 ( .B(n820), .A(n1981), .Z(n821) );
  CND4X4 U1381 ( .A(n824), .B(n823), .C(n822), .D(n821), .Z(n2063) );
  CND2X2 U1382 ( .A(n2063), .B(n2080), .Z(n825) );
  CIVX2 U1383 ( .A(n828), .Z(n829) );
  CND2X4 U1384 ( .A(n830), .B(n829), .Z(n1297) );
  CND2X4 U1385 ( .A(n1297), .B(n1981), .Z(n833) );
  CND2X1 U1386 ( .A(n1062), .B(n1332), .Z(n832) );
  CND2X2 U1387 ( .A(n1063), .B(n1221), .Z(n831) );
  CND3X4 U1388 ( .A(n833), .B(n832), .C(n831), .Z(n2046) );
  CND2X2 U1389 ( .A(n2046), .B(n2080), .Z(n843) );
  CIVDX4 U1390 ( .A(n610), .Z0(n864), .Z1(n1982) );
  CNR2X1 U1391 ( .A(n1385), .B(n610), .Z(n842) );
  CND2IX1 U1392 ( .B(n2596), .A(n842), .Z(n841) );
  CIVX2 U1393 ( .A(n1981), .Z(n1288) );
  CNR2X2 U1394 ( .A(n834), .B(n1288), .Z(n836) );
  CIVX2 U1395 ( .A(n1221), .Z(n1059) );
  CNR2X2 U1396 ( .A(n1398), .B(n1059), .Z(n835) );
  CNR2X4 U1397 ( .A(n836), .B(n835), .Z(n839) );
  CANR2X4 U1398 ( .A(n837), .B(n1332), .C(n1967), .D(n1058), .Z(n838) );
  CND2X4 U1399 ( .A(n839), .B(n838), .Z(n2045) );
  CND2X4 U1400 ( .A(n2045), .B(n1420), .Z(n844) );
  CANR11X2 U1401 ( .A(n843), .B(n841), .C(n844), .D(n840), .Z(n1149) );
  CNR2X4 U1402 ( .A(n1150), .B(n1149), .Z(n1874) );
  CENX1 U1403 ( .A(acc2[28]), .B(n842), .Z(n846) );
  CND2X2 U1404 ( .A(n848), .B(n847), .Z(n849) );
  CNR2X2 U1405 ( .A(n1874), .B(n1867), .Z(n1840) );
  CNR2X2 U1406 ( .A(n1385), .B(n2003), .Z(n880) );
  CENX2 U1407 ( .A(acc2[30]), .B(n880), .Z(n873) );
  CND3X1 U1408 ( .A(n920), .B(n1961), .C(n1425), .Z(n859) );
  CND3X1 U1409 ( .A(n2440), .B(n1961), .C(acc[2]), .Z(n850) );
  CIVX2 U1410 ( .A(n850), .Z(n853) );
  CND2X4 U1411 ( .A(n1201), .B(n588), .Z(n2429) );
  CND2X1 U1412 ( .A(n1961), .B(acc[4]), .Z(n851) );
  CNR2X2 U1413 ( .A(n2429), .B(n851), .Z(n852) );
  CNR2X2 U1414 ( .A(n853), .B(n852), .Z(n857) );
  CIVX2 U1415 ( .A(acc[5]), .Z(n2445) );
  COR4X1 U1416 ( .A(n1425), .B(n2445), .C(n586), .D(n2074), .Z(n856) );
  CNR2IX1 U1417 ( .B(acc[3]), .A(n1425), .Z(n854) );
  CND3X1 U1418 ( .A(n864), .B(n854), .C(n1961), .Z(n855) );
  CND3X2 U1419 ( .A(n856), .B(n857), .C(n855), .Z(n858) );
  CNR2IX4 U1420 ( .B(n859), .A(n858), .Z(n1044) );
  CND2X4 U1421 ( .A(n1192), .B(n1332), .Z(n1042) );
  CND2X2 U1422 ( .A(n1042), .B(n1041), .Z(n860) );
  CIVX2 U1423 ( .A(n860), .Z(n861) );
  CND2X2 U1424 ( .A(n1044), .B(n861), .Z(n1963) );
  CND2X2 U1425 ( .A(n1963), .B(n2080), .Z(n883) );
  CND2X1 U1426 ( .A(n1270), .B(n1332), .Z(n870) );
  CANR1X2 U1427 ( .A(acc[29]), .B(n2590), .C(n863), .Z(n867) );
  CND2X2 U1428 ( .A(n864), .B(acc[27]), .Z(n866) );
  CND2X1 U1429 ( .A(n1201), .B(acc[28]), .Z(n865) );
  CND3X2 U1430 ( .A(n867), .B(n866), .C(n865), .Z(n1417) );
  CND2X1 U1431 ( .A(n1417), .B(n1221), .Z(n869) );
  CND4X2 U1432 ( .A(n871), .B(n870), .C(n869), .D(n868), .Z(n1964) );
  CND2X2 U1433 ( .A(n1964), .B(n2449), .Z(n882) );
  CND2X2 U1434 ( .A(n883), .B(n882), .Z(n872) );
  CND2X2 U1435 ( .A(n874), .B(acc2[29]), .Z(n875) );
  CIVX2 U1436 ( .A(n875), .Z(n1151) );
  CIVX2 U1437 ( .A(n2600), .Z(n877) );
  CND3X4 U1438 ( .A(n878), .B(n879), .C(n877), .Z(n876) );
  COND4CX4 U1439 ( .A(n879), .B(n878), .C(n877), .D(n876), .Z(n1153) );
  CND2IX1 U1440 ( .B(n2591), .A(n880), .Z(n884) );
  CANR11X2 U1441 ( .A(n884), .B(n883), .C(n882), .D(n881), .Z(n1154) );
  CNR2X4 U1442 ( .A(n1153), .B(n1154), .Z(n1837) );
  CND2X2 U1443 ( .A(n1840), .B(n1156), .Z(n1159) );
  CNR2X4 U1444 ( .A(n1864), .B(n1159), .Z(n1443) );
  CIVX2 U1445 ( .A(n1443), .Z(n1361) );
  CIVX2 U1446 ( .A(n1361), .Z(n1161) );
  CIVX4 U1447 ( .A(n885), .Z(n886) );
  CND2X4 U1448 ( .A(n886), .B(n1180), .Z(n1227) );
  CENX1 U1449 ( .A(n2610), .B(n903), .Z(n887) );
  CIVX2 U1450 ( .A(rdy), .Z(n1976) );
  CENX2 U1451 ( .A(n887), .B(n902), .Z(n910) );
  CIVX3 U1452 ( .A(n910), .Z(n889) );
  CND2X2 U1453 ( .A(n987), .B(n594), .Z(n897) );
  CNR2IX2 U1454 ( .B(acc2[3]), .A(n897), .Z(n909) );
  CIVX2 U1455 ( .A(n909), .Z(n888) );
  CND2X4 U1456 ( .A(n889), .B(n888), .Z(n1780) );
  CIVX2 U1457 ( .A(n1227), .Z(n918) );
  CND2X2 U1458 ( .A(n587), .B(acc2[0]), .Z(n1761) );
  CIVX2 U1459 ( .A(n1761), .Z(n1764) );
  CND2X2 U1460 ( .A(acc[0]), .B(n1998), .Z(n1028) );
  CNR3X2 U1461 ( .A(n1048), .B(n2589), .C(n1028), .Z(n890) );
  COR2X2 U1462 ( .A(n890), .B(acc2[1]), .Z(n1763) );
  CIVX4 U1463 ( .A(n440), .Z(n2588) );
  CIVX1 U1464 ( .A(n1028), .Z(n891) );
  CND2X2 U1465 ( .A(n891), .B(acc2[1]), .Z(n892) );
  CNR2X2 U1466 ( .A(n1048), .B(n892), .Z(n893) );
  CND2X2 U1467 ( .A(n2588), .B(n893), .Z(n1762) );
  CNR2X2 U1468 ( .A(n1006), .B(n1961), .Z(n2020) );
  CND2X2 U1469 ( .A(n2020), .B(n2449), .Z(n894) );
  CNR2X2 U1470 ( .A(n598), .B(n1227), .Z(n898) );
  CND2X2 U1471 ( .A(n896), .B(n895), .Z(n1755) );
  COND1X4 U1472 ( .A(n1756), .B(n1754), .C(n1755), .Z(n1759) );
  CENX2 U1473 ( .A(acc2[3]), .B(n897), .Z(n900) );
  CHA1X1 U1474 ( .A(acc2[2]), .B(n898), .CO(n899), .S(n896) );
  COR2X1 U1475 ( .A(n900), .B(n899), .Z(n1758) );
  CND2X2 U1476 ( .A(n1759), .B(n1758), .Z(n901) );
  CND2X1 U1477 ( .A(n900), .B(n899), .Z(n1757) );
  CND2X4 U1478 ( .A(n901), .B(n1757), .Z(n1779) );
  CND2X2 U1479 ( .A(n902), .B(n2610), .Z(n904) );
  CND2IX1 U1480 ( .B(n1092), .A(n1420), .Z(n908) );
  CNR2X2 U1481 ( .A(n1048), .B(n1059), .Z(n906) );
  CND2X2 U1482 ( .A(n1091), .B(n906), .Z(n907) );
  CND3X2 U1483 ( .A(n1780), .B(n1779), .C(n1778), .Z(n916) );
  CND2X4 U1484 ( .A(n910), .B(n909), .Z(n1782) );
  CND2X2 U1485 ( .A(n912), .B(n911), .Z(n1777) );
  CND2X4 U1486 ( .A(n916), .B(n915), .Z(n1752) );
  CND2X2 U1487 ( .A(n2491), .B(n918), .Z(n926) );
  CENX2 U1488 ( .A(n926), .B(n2652), .Z(n925) );
  CND2X2 U1489 ( .A(n919), .B(n1197), .Z(n924) );
  CND2IX1 U1490 ( .B(n588), .A(n920), .Z(n1078) );
  CIVX2 U1491 ( .A(n1078), .Z(n922) );
  CND2X2 U1492 ( .A(n922), .B(n921), .Z(n923) );
  CENX2 U1493 ( .A(n925), .B(n928), .Z(n932) );
  CIVX2 U1494 ( .A(n934), .Z(n930) );
  CIVX2 U1495 ( .A(n926), .Z(n927) );
  CIVX2 U1496 ( .A(n935), .Z(n929) );
  CND2X1 U1497 ( .A(n1750), .B(n1742), .Z(n1714) );
  CNR2X1 U1498 ( .A(n1040), .B(n421), .Z(n955) );
  CEN3X1 U1499 ( .A(acc2[8]), .B(n955), .C(n954), .Z(n939) );
  CNR2IX2 U1500 ( .B(acc2[7]), .A(n931), .Z(n938) );
  CNR2X2 U1501 ( .A(n939), .B(n938), .Z(n1710) );
  CNR2X2 U1502 ( .A(n1714), .B(n1710), .Z(n1693) );
  CND2X2 U1503 ( .A(n933), .B(n932), .Z(n1749) );
  CIVX2 U1504 ( .A(n1741), .Z(n936) );
  CANR1X4 U1505 ( .A(n1742), .B(n937), .C(n936), .Z(n1713) );
  CND2X1 U1506 ( .A(n939), .B(n938), .Z(n1711) );
  COND1X4 U1507 ( .A(n1710), .B(n1713), .C(n1711), .Z(n1692) );
  CENX2 U1508 ( .A(acc2[13]), .B(n1039), .Z(n981) );
  CND2X4 U1509 ( .A(n2046), .B(n2449), .Z(n941) );
  CNR2X1 U1510 ( .A(n1040), .B(n610), .Z(n940) );
  CNR2X4 U1511 ( .A(n981), .B(n980), .Z(n1726) );
  CENX1 U1512 ( .A(n2611), .B(n940), .Z(n942) );
  CND2X2 U1513 ( .A(n2053), .B(n1420), .Z(n960) );
  CNR2IX2 U1514 ( .B(acc2[11]), .A(n960), .Z(n978) );
  CNR2X4 U1515 ( .A(n979), .B(n978), .Z(n1734) );
  CNR2X2 U1516 ( .A(n1726), .B(n1734), .Z(n983) );
  CND2X4 U1517 ( .A(n2083), .B(n1420), .Z(n951) );
  CIVX3 U1518 ( .A(n951), .Z(n943) );
  CND2X4 U1519 ( .A(n943), .B(acc2[9]), .Z(n967) );
  CANR11X4 U1520 ( .A(n946), .B(n945), .C(n944), .D(n1048), .Z(n970) );
  CNR2X4 U1521 ( .A(n1040), .B(n598), .Z(n968) );
  CENX2 U1522 ( .A(n970), .B(n947), .Z(n948) );
  CIVX2 U1523 ( .A(n2612), .Z(n950) );
  CNR2IX2 U1524 ( .B(n1420), .A(n950), .Z(n949) );
  CND2X2 U1525 ( .A(n2083), .B(n949), .Z(n953) );
  CND2X4 U1526 ( .A(n951), .B(n950), .Z(n952) );
  CND2X4 U1527 ( .A(n953), .B(n952), .Z(n966) );
  CNIVX2 U1528 ( .A(n955), .Z(n956) );
  CND2X4 U1529 ( .A(n957), .B(n956), .Z(n964) );
  CND3X2 U1530 ( .A(n2067), .B(n1420), .C(acc2[8]), .Z(n963) );
  CND2X2 U1531 ( .A(n964), .B(n963), .Z(n958) );
  CIVX4 U1532 ( .A(n959), .Z(n1707) );
  CENX2 U1533 ( .A(n960), .B(acc2[11]), .Z(n976) );
  COND1X2 U1534 ( .A(acc2[10]), .B(n970), .C(n968), .Z(n962) );
  CND2X2 U1535 ( .A(n962), .B(n961), .Z(n975) );
  CNR2X4 U1536 ( .A(n976), .B(n975), .Z(n974) );
  CNR2X2 U1537 ( .A(n1699), .B(n974), .Z(n1738) );
  CND2X2 U1538 ( .A(n983), .B(n1738), .Z(n985) );
  CND2X4 U1539 ( .A(n966), .B(n965), .Z(n1706) );
  CENX1 U1540 ( .A(acc2[10]), .B(n968), .Z(n969) );
  CENX1 U1541 ( .A(n970), .B(n969), .Z(n971) );
  CND2X4 U1542 ( .A(n972), .B(n971), .Z(n1690) );
  COND1X4 U1543 ( .A(n1706), .B(n973), .C(n1690), .Z(n1700) );
  CND2X4 U1544 ( .A(n1700), .B(n1698), .Z(n977) );
  CND2X1 U1545 ( .A(n976), .B(n975), .Z(n1697) );
  CND2X4 U1546 ( .A(n977), .B(n1697), .Z(n1729) );
  COND1X2 U1547 ( .A(n1726), .B(n1735), .C(n1727), .Z(n982) );
  CANR1X4 U1548 ( .A(n983), .B(n1729), .C(n982), .Z(n984) );
  CNR2X2 U1549 ( .A(n2437), .B(n1425), .Z(n1068) );
  CNIVX4 U1550 ( .A(n987), .Z(n1990) );
  CND2X2 U1551 ( .A(n1068), .B(n1990), .Z(n1072) );
  CND2X2 U1552 ( .A(n989), .B(n1981), .Z(n994) );
  CND2X2 U1553 ( .A(n990), .B(n1221), .Z(n993) );
  CND2X2 U1554 ( .A(n991), .B(n1967), .Z(n992) );
  CND2X2 U1555 ( .A(n1989), .B(n2449), .Z(n1071) );
  CIVX2 U1556 ( .A(n2608), .Z(n996) );
  CANR1X2 U1557 ( .A(n1072), .B(n1071), .C(n996), .Z(n995) );
  CIVX2 U1558 ( .A(n995), .Z(n998) );
  CND2X4 U1559 ( .A(n998), .B(n997), .Z(n1123) );
  CND2X1 U1560 ( .A(n1197), .B(n605), .Z(n1000) );
  CND2X2 U1561 ( .A(n1192), .B(n603), .Z(n999) );
  CND2X2 U1562 ( .A(n1000), .B(n999), .Z(n1005) );
  CND2X2 U1563 ( .A(n1196), .B(n2471), .Z(n1003) );
  CND2X1 U1564 ( .A(n1193), .B(n601), .Z(n1002) );
  CND2X2 U1565 ( .A(n1003), .B(n1002), .Z(n1004) );
  CNR2X4 U1566 ( .A(n1005), .B(n1004), .Z(n1008) );
  COR2X1 U1567 ( .A(n2437), .B(n1006), .Z(n1007) );
  CND2X4 U1568 ( .A(n1008), .B(n1007), .Z(n1013) );
  CND2X4 U1569 ( .A(n1981), .B(n1180), .Z(n1082) );
  CNIVX4 U1570 ( .A(n1082), .Z(n1009) );
  CNR2X4 U1571 ( .A(n1009), .B(n608), .Z(n1012) );
  COND1X4 U1572 ( .A(acc2[18]), .B(n1013), .C(n1012), .Z(n1011) );
  CND2X2 U1573 ( .A(n1013), .B(acc2[18]), .Z(n1010) );
  CND2X4 U1574 ( .A(n1011), .B(n1010), .Z(n1122) );
  CNR2X4 U1575 ( .A(n1123), .B(n1122), .Z(n1638) );
  CENX4 U1576 ( .A(n1014), .B(n1013), .Z(n1117) );
  COND1X2 U1577 ( .A(n1016), .B(n1015), .C(n1967), .Z(n1020) );
  CND2X4 U1578 ( .A(n1020), .B(n1019), .Z(n1168) );
  CIVX4 U1579 ( .A(n1023), .Z(n1024) );
  COND1X4 U1580 ( .A(n1025), .B(n1024), .C(n1332), .Z(n1026) );
  CND2X4 U1581 ( .A(n1026), .B(n1027), .Z(n1169) );
  COND1X4 U1582 ( .A(n1168), .B(n1169), .C(n1420), .Z(n1030) );
  COR2X1 U1583 ( .A(n2589), .B(n1028), .Z(n1179) );
  COR2X1 U1584 ( .A(n1179), .B(n2056), .Z(n1029) );
  CND2X4 U1585 ( .A(n1118), .B(n1117), .Z(n1644) );
  CND2IX4 U1586 ( .B(n1048), .A(n2040), .Z(n1031) );
  CNR2X2 U1587 ( .A(n1082), .B(n421), .Z(n1036) );
  CND2X4 U1588 ( .A(n1033), .B(n1032), .Z(n1121) );
  CIVX2 U1589 ( .A(n1121), .Z(n1035) );
  CND2X4 U1590 ( .A(n1035), .B(n527), .Z(n1655) );
  CND2X4 U1591 ( .A(n1644), .B(n1655), .Z(n1632) );
  CNR2X4 U1592 ( .A(n1638), .B(n1632), .Z(n1587) );
  CENX2 U1593 ( .A(acc2[16]), .B(n1036), .Z(n1038) );
  CENX4 U1594 ( .A(n1038), .B(n1037), .Z(n1116) );
  CND2X4 U1595 ( .A(n1960), .B(n1420), .Z(n1046) );
  CNR2IX2 U1596 ( .B(acc2[15]), .A(n1046), .Z(n1115) );
  CNR2X4 U1597 ( .A(n1116), .B(n1115), .Z(n1673) );
  CNR2IX2 U1598 ( .B(acc2[13]), .A(n1039), .Z(n1110) );
  CNR2X1 U1599 ( .A(n1040), .B(n2003), .Z(n1050) );
  CENX1 U1600 ( .A(acc2[14]), .B(n1050), .Z(n1045) );
  CND2X2 U1601 ( .A(n1042), .B(n1041), .Z(n1043) );
  CANR1X4 U1602 ( .A(n1044), .B(n1047), .C(n1048), .Z(n1053) );
  CENX4 U1603 ( .A(acc2[15]), .B(n1046), .Z(n1112) );
  CIVX2 U1604 ( .A(n1112), .Z(n1057) );
  CND2IX1 U1605 ( .B(acc2[14]), .A(n1048), .Z(n1049) );
  CAN2X1 U1606 ( .A(n1050), .B(n1049), .Z(n1051) );
  CND2X2 U1607 ( .A(n1052), .B(n1051), .Z(n1055) );
  CND2X2 U1608 ( .A(n1053), .B(acc2[14]), .Z(n1054) );
  CIVX2 U1609 ( .A(n1111), .Z(n1056) );
  CND2X4 U1610 ( .A(n1057), .B(n1056), .Z(n1807) );
  CND2X2 U1611 ( .A(n451), .B(n1807), .Z(n1672) );
  CNR2X4 U1612 ( .A(n1673), .B(n1672), .Z(n1656) );
  CENX1 U1613 ( .A(acc2[20]), .B(n1103), .Z(n1070) );
  CND2X1 U1614 ( .A(n1058), .B(n1332), .Z(n1067) );
  CIVX2 U1615 ( .A(n1059), .Z(n1060) );
  CND2X2 U1616 ( .A(n1061), .B(n1060), .Z(n1066) );
  CND2X1 U1617 ( .A(n1062), .B(n1967), .Z(n1065) );
  CND2X2 U1618 ( .A(n1063), .B(n1981), .Z(n1064) );
  CND4X4 U1619 ( .A(n1067), .B(n1066), .C(n1065), .D(n1064), .Z(n1975) );
  CND2X2 U1620 ( .A(n1975), .B(n2449), .Z(n1102) );
  CNIVX4 U1621 ( .A(n1297), .Z(n1978) );
  CND2X1 U1622 ( .A(n1978), .B(n1068), .Z(n1069) );
  CND2X2 U1623 ( .A(n1102), .B(n1069), .Z(n1101) );
  CENX2 U1624 ( .A(n1070), .B(n1101), .Z(n1124) );
  CIVX2 U1625 ( .A(n1125), .Z(n1073) );
  CNR2X2 U1626 ( .A(n1124), .B(n1073), .Z(n1588) );
  CIVX2 U1627 ( .A(n1588), .Z(n1109) );
  CND2X2 U1628 ( .A(n1192), .B(n1967), .Z(n1077) );
  CND2X2 U1629 ( .A(n1205), .B(n1221), .Z(n1075) );
  CND2X2 U1630 ( .A(n1193), .B(n1981), .Z(n1074) );
  CND4X4 U1631 ( .A(n1077), .B(n1076), .C(n1075), .D(n1074), .Z(n1269) );
  CND2X4 U1632 ( .A(n1197), .B(n588), .Z(n1079) );
  CND2X4 U1633 ( .A(n1079), .B(n1078), .Z(n1999) );
  CND2IX1 U1634 ( .B(n2437), .A(n1999), .Z(n1080) );
  CND2X4 U1635 ( .A(n1081), .B(n1080), .Z(n1098) );
  CNR2X2 U1636 ( .A(n1082), .B(n2003), .Z(n1097) );
  CENX2 U1637 ( .A(acc2[22]), .B(n1097), .Z(n1083) );
  CENX2 U1638 ( .A(n1083), .B(n1098), .Z(n1130) );
  CND2X4 U1639 ( .A(n1085), .B(n1967), .Z(n1088) );
  CND2X4 U1640 ( .A(n1091), .B(n1221), .Z(n1093) );
  CND2X4 U1641 ( .A(n1093), .B(n1092), .Z(n1984) );
  CAN2X2 U1642 ( .A(n1108), .B(acc2[21]), .Z(n1129) );
  CENX4 U1643 ( .A(n2604), .B(n1096), .Z(n1132) );
  COND1X4 U1644 ( .A(acc2[22]), .B(n1098), .C(n1097), .Z(n1100) );
  CND2X2 U1645 ( .A(n1098), .B(acc2[22]), .Z(n1099) );
  CND2X4 U1646 ( .A(n1100), .B(n1099), .Z(n1131) );
  CNR2X4 U1647 ( .A(n1131), .B(n1132), .Z(n1607) );
  CNR2X4 U1648 ( .A(n1617), .B(n1607), .Z(n1134) );
  CND2X2 U1649 ( .A(n1101), .B(acc2[20]), .Z(n1107) );
  CIVX1 U1650 ( .A(n2594), .Z(n1105) );
  CIVX2 U1651 ( .A(n1102), .Z(n1104) );
  COND1X4 U1652 ( .A(n1105), .B(n1104), .C(n1103), .Z(n1106) );
  CND2X4 U1653 ( .A(n1107), .B(n1106), .Z(n1126) );
  CENX2 U1654 ( .A(n2644), .B(n1108), .Z(n1127) );
  CNR2X4 U1655 ( .A(n1126), .B(n1127), .Z(n1128) );
  CIVX3 U1656 ( .A(n1128), .Z(n1600) );
  CNR2X4 U1657 ( .A(n1591), .B(n1137), .Z(n1445) );
  CND2X4 U1658 ( .A(n1646), .B(n1445), .Z(n1139) );
  CANR1X4 U1659 ( .A(n1807), .B(n1114), .C(n1113), .Z(n1670) );
  CND2X2 U1660 ( .A(n1116), .B(n1115), .Z(n1674) );
  COND1X4 U1661 ( .A(n1673), .B(n1670), .C(n1674), .Z(n1659) );
  CIVX2 U1662 ( .A(n1117), .Z(n1120) );
  CIVX2 U1663 ( .A(n1118), .Z(n1119) );
  CND2X4 U1664 ( .A(n1645), .B(n1644), .Z(n1633) );
  CND2X2 U1665 ( .A(n1123), .B(n1122), .Z(n1639) );
  COND4CX4 U1666 ( .A(n1643), .B(n1633), .C(n1638), .D(n1639), .Z(n1586) );
  CANR1X2 U1667 ( .A(n1587), .B(n1659), .C(n1586), .Z(n1136) );
  CND2X2 U1668 ( .A(n1127), .B(n1126), .Z(n1596) );
  COND1X4 U1669 ( .A(n1592), .B(n1128), .C(n1596), .Z(n1613) );
  CND2X2 U1670 ( .A(n1130), .B(n1129), .Z(n1618) );
  CND2X2 U1671 ( .A(n1132), .B(n1131), .Z(n1608) );
  COND1X2 U1672 ( .A(n1618), .B(n1607), .C(n1608), .Z(n1133) );
  CANR1X2 U1673 ( .A(n1134), .B(n1613), .C(n1133), .Z(n1135) );
  COND1X2 U1674 ( .A(n1137), .B(n1136), .C(n1135), .Z(n1444) );
  CIVX2 U1675 ( .A(n1444), .Z(n1138) );
  CND2X4 U1676 ( .A(n1139), .B(n1138), .Z(n1904) );
  CND2X2 U1677 ( .A(n1143), .B(n1142), .Z(n1901) );
  CND2X2 U1678 ( .A(n1144), .B(n1145), .Z(n1891) );
  CND2X2 U1679 ( .A(n1147), .B(n1146), .Z(n1883) );
  COND1X2 U1680 ( .A(n1891), .B(n1882), .C(n1883), .Z(n1842) );
  CANR1X2 U1681 ( .A(n1843), .B(n1885), .C(n1842), .Z(n1158) );
  CND2X2 U1682 ( .A(n1148), .B(n595), .Z(n1869) );
  CND2X2 U1683 ( .A(n1150), .B(n1149), .Z(n1875) );
  COND1X2 U1684 ( .A(n1874), .B(n1869), .C(n1875), .Z(n1844) );
  CND2X2 U1685 ( .A(n1154), .B(n1153), .Z(n1838) );
  COND1X2 U1686 ( .A(n1837), .B(n1853), .C(n1838), .Z(n1155) );
  CANR1X2 U1687 ( .A(n1156), .B(n1844), .C(n1155), .Z(n1157) );
  COND1X2 U1688 ( .A(n1159), .B(n1158), .C(n1157), .Z(n1456) );
  CIVX3 U1689 ( .A(n1456), .Z(n1362) );
  CIVX2 U1690 ( .A(n1362), .Z(n1160) );
  CANR1X1 U1691 ( .A(n1161), .B(n1904), .C(n1160), .Z(n1162) );
  CEOX2 U1692 ( .A(n1163), .B(n1162), .Z(n1949) );
  CIVX2 U1693 ( .A(n1949), .Z(n2532) );
  COND1X4 U1694 ( .A(acc2[32]), .B(n1165), .C(n1164), .Z(n1167) );
  CND2X2 U1695 ( .A(n1165), .B(acc2[32]), .Z(n1166) );
  CND2X4 U1696 ( .A(n1167), .B(n1166), .Z(n1241) );
  CNR2X2 U1697 ( .A(n2029), .B(n2056), .Z(n1170) );
  CND2X2 U1698 ( .A(n1201), .B(acc[31]), .Z(n1174) );
  CND2X1 U1699 ( .A(n1171), .B(acc[30]), .Z(n1173) );
  CND2X1 U1700 ( .A(n1202), .B(acc[29]), .Z(n1172) );
  CANR2X2 U1701 ( .A(n1175), .B(n1967), .C(n1221), .D(n1408), .Z(n1178) );
  CND2X1 U1702 ( .A(n1407), .B(n1332), .Z(n1177) );
  CND2X1 U1703 ( .A(n1275), .B(n1981), .Z(n1176) );
  CND3X2 U1704 ( .A(n1178), .B(n1177), .C(n1176), .Z(n2027) );
  CIVX2 U1705 ( .A(n1179), .Z(n2025) );
  CND2X4 U1706 ( .A(n1180), .B(rdy), .Z(n2028) );
  CIVX12 U1707 ( .A(n2028), .Z(n2087) );
  CAN2X2 U1708 ( .A(n2025), .B(n2087), .Z(n1181) );
  CANR1X4 U1709 ( .A(n2449), .B(n2027), .C(n1181), .Z(n1182) );
  CND2X4 U1710 ( .A(n1183), .B(n1182), .Z(n1236) );
  CENX4 U1711 ( .A(n2609), .B(n1236), .Z(n1240) );
  CNR2X2 U1712 ( .A(n1241), .B(n1240), .Z(n1239) );
  CIVXL U1713 ( .A(n1239), .Z(n1184) );
  CND2X2 U1714 ( .A(n1240), .B(n1241), .Z(n1242) );
  CND2X1 U1715 ( .A(n1184), .B(n1242), .Z(n1190) );
  CIVX1 U1716 ( .A(n1185), .Z(n1186) );
  CNR2X1 U1717 ( .A(n1361), .B(n1186), .Z(n1188) );
  COND1X1 U1718 ( .A(n1186), .B(n1362), .C(n1244), .Z(n1187) );
  CANR1X2 U1719 ( .A(n1188), .B(n1904), .C(n1187), .Z(n1189) );
  CEOX2 U1720 ( .A(n1190), .B(n1189), .Z(n1191) );
  CNR2IX4 U1721 ( .B(x[33]), .A(n1191), .Z(n1950) );
  CNR3X1 U1722 ( .A(n2532), .B(x[32]), .C(n1950), .Z(n1262) );
  CIVX2 U1723 ( .A(n1191), .Z(n2556) );
  CNR2X1 U1724 ( .A(n2556), .B(x[33]), .Z(n1261) );
  CNR2X2 U1725 ( .A(n608), .B(n1977), .Z(n1233) );
  CND2X2 U1726 ( .A(n1192), .B(n1981), .Z(n1195) );
  CND2X4 U1727 ( .A(n1195), .B(n1194), .Z(n2015) );
  CND2X2 U1728 ( .A(n1196), .B(n1221), .Z(n1199) );
  CND2X1 U1729 ( .A(n1197), .B(n1967), .Z(n1198) );
  CND2X2 U1730 ( .A(n1199), .B(n1198), .Z(n2016) );
  COND1X4 U1731 ( .A(n2015), .B(n2016), .C(n2080), .Z(n1217) );
  CND2X2 U1732 ( .A(n1217), .B(n2639), .Z(n1200) );
  CANR1X2 U1733 ( .A(n2449), .B(n2019), .C(n1204), .Z(n1216) );
  CND2X2 U1734 ( .A(n1270), .B(n1981), .Z(n1206) );
  CND2X4 U1735 ( .A(n1206), .B(n1207), .Z(n2017) );
  CIVX4 U1736 ( .A(n2017), .Z(n1213) );
  CND2X2 U1737 ( .A(n1416), .B(n1221), .Z(n1211) );
  CND4X1 U1738 ( .A(n864), .B(n1425), .C(acc[27]), .D(n1998), .Z(n1210) );
  CND2X2 U1739 ( .A(n1211), .B(n1210), .Z(n2018) );
  CIVX3 U1740 ( .A(n2018), .Z(n1212) );
  CND2X4 U1741 ( .A(n1213), .B(n1212), .Z(n1214) );
  CND2X4 U1742 ( .A(n1214), .B(n2449), .Z(n1215) );
  CND3X4 U1743 ( .A(n1217), .B(n1215), .C(n1216), .Z(n1234) );
  CND2X2 U1744 ( .A(n1234), .B(acc2[34]), .Z(n1218) );
  CND2X4 U1745 ( .A(n1218), .B(n1219), .Z(n1285) );
  CNIVX1 U1746 ( .A(n1285), .Z(n1230) );
  CND2X2 U1747 ( .A(n1331), .B(n1981), .Z(n1226) );
  CND2X2 U1748 ( .A(n1426), .B(n1332), .Z(n1225) );
  CNR2IX2 U1749 ( .B(acc[31]), .A(n1220), .Z(n1962) );
  CND2X1 U1750 ( .A(n1962), .B(n1221), .Z(n1224) );
  CND4X4 U1751 ( .A(n1226), .B(n1223), .C(n1224), .D(n1225), .Z(n1988) );
  CND2X4 U1752 ( .A(n1988), .B(n2449), .Z(n1228) );
  CNR2X1 U1753 ( .A(n1227), .B(n1976), .Z(n1296) );
  CND3X4 U1754 ( .A(n1229), .B(n1228), .C(n596), .Z(n1309) );
  CENX4 U1755 ( .A(n2638), .B(n1309), .Z(n1284) );
  CNR2X1 U1756 ( .A(n1230), .B(n1284), .Z(n1231) );
  CIVX2 U1757 ( .A(n1231), .Z(n1232) );
  CND2X1 U1758 ( .A(n1232), .B(n1310), .Z(n1251) );
  CENX1 U1759 ( .A(acc2[34]), .B(n1233), .Z(n1235) );
  CENX2 U1760 ( .A(n1235), .B(n1234), .Z(n1246) );
  CND2X2 U1761 ( .A(n1236), .B(acc2[33]), .Z(n1237) );
  CIVX3 U1762 ( .A(n1237), .Z(n1245) );
  CNR2X4 U1763 ( .A(n1246), .B(n1245), .Z(n1286) );
  CIVX2 U1764 ( .A(n1286), .Z(n1252) );
  CNR2X4 U1765 ( .A(n1239), .B(n1238), .Z(n1287) );
  CND2X1 U1766 ( .A(n1252), .B(n1287), .Z(n1247) );
  CNR2X1 U1767 ( .A(n1361), .B(n1247), .Z(n1249) );
  CNR2X2 U1768 ( .A(n1241), .B(n1240), .Z(n1243) );
  COND1X2 U1769 ( .A(n1244), .B(n1243), .C(n1242), .Z(n1314) );
  CIVX2 U1770 ( .A(n1314), .Z(n1253) );
  CND2X4 U1771 ( .A(n1246), .B(n1245), .Z(n1312) );
  CANR1X1 U1772 ( .A(n1249), .B(n1904), .C(n1248), .Z(n1250) );
  CEOX2 U1773 ( .A(n1251), .B(n1250), .Z(n1263) );
  CNR2IX2 U1774 ( .B(x[35]), .A(n1263), .Z(n1260) );
  CND2X2 U1775 ( .A(n1252), .B(n1312), .Z(n1258) );
  CIVX2 U1776 ( .A(n1287), .Z(n1254) );
  CNR2X1 U1777 ( .A(n1361), .B(n1254), .Z(n1256) );
  COND1X1 U1778 ( .A(n1254), .B(n1362), .C(n1253), .Z(n1255) );
  CANR1X1 U1779 ( .A(n1256), .B(n1904), .C(n1255), .Z(n1257) );
  CEOX2 U1780 ( .A(n1258), .B(n1257), .Z(n1264) );
  CNR2IX1 U1781 ( .B(x[34]), .A(n1264), .Z(n1259) );
  CNR2X2 U1782 ( .A(n1260), .B(n1259), .Z(n1952) );
  COND1X1 U1783 ( .A(n1262), .B(n1261), .C(n1952), .Z(n1268) );
  CIVX2 U1784 ( .A(n1263), .Z(n2575) );
  CIVX2 U1785 ( .A(n1264), .Z(n2547) );
  CANR3X2 U1786 ( .A(n2575), .B(x[35]), .C(n2547), .D(x[34]), .Z(n1266) );
  CNR2X1 U1787 ( .A(n2575), .B(x[35]), .Z(n1265) );
  CNR2X1 U1788 ( .A(n1266), .B(n1265), .Z(n1267) );
  CNR2X2 U1789 ( .A(n1977), .B(n2003), .Z(n1327) );
  CENX1 U1790 ( .A(acc2[38]), .B(n1327), .Z(n1274) );
  CIVX3 U1791 ( .A(n1269), .Z(n2002) );
  CND2X2 U1792 ( .A(n1417), .B(n1981), .Z(n1995) );
  CND2X1 U1793 ( .A(n1416), .B(n1332), .Z(n1997) );
  CAN2X1 U1794 ( .A(n2087), .B(n1998), .Z(n1271) );
  CANR2X4 U1795 ( .A(n1272), .B(n1420), .C(n1271), .D(n1999), .Z(n1273) );
  CENX2 U1796 ( .A(n1274), .B(n537), .Z(n1282) );
  CND2X1 U1797 ( .A(n1407), .B(n1981), .Z(n1277) );
  CND2X1 U1798 ( .A(n1408), .B(n1332), .Z(n1276) );
  CND3X4 U1799 ( .A(n1281), .B(n1280), .C(n1279), .Z(n1302) );
  CNR2X4 U1800 ( .A(n1282), .B(n592), .Z(n1440) );
  CIVXL U1801 ( .A(n419), .Z(n1283) );
  CND2X2 U1802 ( .A(n1282), .B(n592), .Z(n1448) );
  CAN2X2 U1803 ( .A(n1448), .B(n1283), .Z(n1326) );
  CNR2X4 U1804 ( .A(n539), .B(n1286), .Z(n1315) );
  CND2X4 U1805 ( .A(n1287), .B(n1315), .Z(n1442) );
  CIVX2 U1806 ( .A(n1442), .Z(n1352) );
  CNR2X2 U1807 ( .A(n2047), .B(n815), .Z(n1289) );
  CIVX2 U1808 ( .A(n1289), .Z(n1294) );
  CNR2X2 U1809 ( .A(n1291), .B(n1290), .Z(n1292) );
  CIVX3 U1810 ( .A(n1292), .Z(n1293) );
  CND3X4 U1811 ( .A(n1295), .B(n1294), .C(n1293), .Z(n1979) );
  CND2X4 U1812 ( .A(n1979), .B(n2449), .Z(n1305) );
  CNR2X2 U1813 ( .A(n1977), .B(n1982), .Z(n1303) );
  CND2X1 U1814 ( .A(n1303), .B(acc2[36]), .Z(n1299) );
  CNR2IX1 U1815 ( .B(n1299), .A(n1298), .Z(n1301) );
  CND2X2 U1816 ( .A(n1975), .B(n2080), .Z(n1306) );
  CANR11X2 U1817 ( .A(n1305), .B(n1301), .C(n1306), .D(n1300), .Z(n1317) );
  CENX4 U1818 ( .A(n2598), .B(n1302), .Z(n1318) );
  CNR2X4 U1819 ( .A(n1317), .B(n1318), .Z(n1348) );
  CENX1 U1820 ( .A(acc2[36]), .B(n1303), .Z(n1308) );
  CND3X2 U1821 ( .A(n1306), .B(n1305), .C(n1304), .Z(n1307) );
  CAN2X4 U1822 ( .A(n1309), .B(acc2[35]), .Z(n1316) );
  CND2X1 U1823 ( .A(n1352), .B(n1320), .Z(n1322) );
  CNR2X1 U1824 ( .A(n1361), .B(n1322), .Z(n1324) );
  CANR1X4 U1825 ( .A(n1315), .B(n1314), .C(n1313), .Z(n1453) );
  CIVX2 U1826 ( .A(n1453), .Z(n1353) );
  CND2X2 U1827 ( .A(n1318), .B(n1317), .Z(n1350) );
  COND1X4 U1828 ( .A(n1359), .B(n1348), .C(n1350), .Z(n1450) );
  CNIVX1 U1829 ( .A(n1450), .Z(n1319) );
  CANR1X1 U1830 ( .A(n1353), .B(n1320), .C(n1319), .Z(n1321) );
  COND1X1 U1831 ( .A(n1322), .B(n1362), .C(n1321), .Z(n1323) );
  CANR1X1 U1832 ( .A(n1324), .B(n1904), .C(n1323), .Z(n1325) );
  COND1X4 U1833 ( .A(acc2[38]), .B(n1328), .C(n1327), .Z(n1330) );
  CND2X2 U1834 ( .A(n537), .B(acc2[38]), .Z(n1329) );
  CND2X4 U1835 ( .A(n1330), .B(n1329), .Z(n1439) );
  CND2X1 U1836 ( .A(n1331), .B(n1967), .Z(n1335) );
  CND2X1 U1837 ( .A(n1426), .B(n1981), .Z(n1334) );
  CND2X1 U1838 ( .A(n1962), .B(n1332), .Z(n1333) );
  CND3X2 U1839 ( .A(n1335), .B(n1334), .C(n1333), .Z(n2012) );
  CND2X2 U1840 ( .A(n2012), .B(n1420), .Z(n1337) );
  CND3X4 U1841 ( .A(n1338), .B(n1337), .C(n1336), .Z(n1415) );
  CENX4 U1842 ( .A(n2606), .B(n1415), .Z(n1438) );
  CND2X2 U1843 ( .A(n1438), .B(n1439), .Z(n1446) );
  CIVDX1 U1844 ( .A(n1441), .Z0(n1339), .Z1(n1320) );
  CNR2X1 U1845 ( .A(n1339), .B(n419), .Z(n1342) );
  CND2X1 U1846 ( .A(n1342), .B(n1352), .Z(n1344) );
  CNR2X1 U1847 ( .A(n1344), .B(n1361), .Z(n1346) );
  CIVX2 U1848 ( .A(n1450), .Z(n1340) );
  COND1XL U1849 ( .A(n419), .B(n1340), .C(n1448), .Z(n1341) );
  CANR1X1 U1850 ( .A(n1353), .B(n1342), .C(n1341), .Z(n1343) );
  COND1X1 U1851 ( .A(n1362), .B(n1344), .C(n1343), .Z(n1345) );
  CIVXL U1852 ( .A(n1348), .Z(n1349) );
  CND2X1 U1853 ( .A(n1350), .B(n1349), .Z(n1358) );
  CIVX2 U1854 ( .A(n1351), .Z(n1360) );
  CND2X1 U1855 ( .A(n1352), .B(n1360), .Z(n1354) );
  CNR2X1 U1856 ( .A(n1361), .B(n1354), .Z(n1356) );
  CANR1X2 U1857 ( .A(n1356), .B(n1904), .C(n1355), .Z(n1357) );
  CAN2X2 U1858 ( .A(n1360), .B(n1359), .Z(n1366) );
  CNR2X1 U1859 ( .A(n1361), .B(n1442), .Z(n1364) );
  COND1XL U1860 ( .A(n1442), .B(n1362), .C(n1453), .Z(n1363) );
  CANR1X1 U1861 ( .A(n1364), .B(n1904), .C(n1363), .Z(n1365) );
  CENX2 U1862 ( .A(n1366), .B(n1365), .Z(n1369) );
  CNR2IX2 U1863 ( .B(x[36]), .A(n1369), .Z(n1367) );
  CNR2X2 U1864 ( .A(n1368), .B(n1367), .Z(n1954) );
  CIVX2 U1865 ( .A(n1369), .Z(n2542) );
  CNR3X2 U1866 ( .A(n2542), .B(x[36]), .C(n1370), .Z(n1375) );
  CIVX2 U1867 ( .A(n1371), .Z(n2549) );
  CNR2X1 U1868 ( .A(n2549), .B(x[37]), .Z(n1374) );
  COND1X2 U1869 ( .A(n1375), .B(n1374), .C(n1373), .Z(n1382) );
  CIVX2 U1870 ( .A(n1376), .Z(n2507) );
  CNR3X1 U1871 ( .A(n1377), .B(n2507), .C(x[38]), .Z(n1380) );
  CIVX2 U1872 ( .A(n1378), .Z(n2516) );
  CNR2X1 U1873 ( .A(n2516), .B(x[39]), .Z(n1379) );
  CNR2X2 U1874 ( .A(n1380), .B(n1379), .Z(n1381) );
  CND2X2 U1875 ( .A(n1382), .B(n1381), .Z(n1383) );
  CNR2X1 U1876 ( .A(n1385), .B(rdy), .Z(n1501) );
  CND2IX1 U1877 ( .B(n2047), .A(n1501), .Z(n1387) );
  CND2X2 U1878 ( .A(n2046), .B(n2087), .Z(n1386) );
  CND2X2 U1879 ( .A(n1332), .B(n1980), .Z(n1480) );
  CNR2X1 U1880 ( .A(n1480), .B(n610), .Z(n1435) );
  CND2X2 U1881 ( .A(n540), .B(acc2[44]), .Z(n1390) );
  CND2X4 U1882 ( .A(n1391), .B(n1390), .Z(n1396) );
  CAN2X1 U1883 ( .A(n1501), .B(n1408), .Z(n1392) );
  CANR1X2 U1884 ( .A(n2080), .B(n2062), .C(n1392), .Z(n1394) );
  CND2X1 U1885 ( .A(n2063), .B(n2087), .Z(n1393) );
  CND2X2 U1886 ( .A(n1394), .B(n1393), .Z(n1486) );
  CENX2 U1887 ( .A(n2593), .B(n1486), .Z(n1395) );
  CNR2X4 U1888 ( .A(n1396), .B(n1395), .Z(n1479) );
  CIVXL U1889 ( .A(n1479), .Z(n1397) );
  CND2X1 U1890 ( .A(n1396), .B(n1395), .Z(n1478) );
  CAN2X1 U1891 ( .A(n1397), .B(n1478), .Z(n1475) );
  CND2X1 U1892 ( .A(n1398), .B(n1425), .Z(n1399) );
  CND3X2 U1893 ( .A(n1400), .B(n1399), .C(n1961), .Z(n2070) );
  CND2X1 U1894 ( .A(n2069), .B(n2026), .Z(n1402) );
  CNR2X2 U1895 ( .A(n1480), .B(n1404), .Z(n1412) );
  CND2X2 U1896 ( .A(n1406), .B(n1405), .Z(n1464) );
  CMX2GX1 U1897 ( .GN(n1998), .A0(n1408), .A1(n1407), .S(n1425), .Z(n2081) );
  CND2X1 U1898 ( .A(n2081), .B(n1420), .Z(n1411) );
  CND2X2 U1899 ( .A(n2082), .B(n2080), .Z(n1410) );
  CENX1 U1900 ( .A(acc2[40]), .B(n1412), .Z(n1414) );
  CENX2 U1901 ( .A(n1414), .B(n1413), .Z(n1463) );
  CAN2X4 U1902 ( .A(n1415), .B(acc2[39]), .Z(n1462) );
  CNR2X2 U1903 ( .A(n1463), .B(n1462), .Z(n1542) );
  CNR2X2 U1904 ( .A(n1544), .B(n1542), .Z(n1526) );
  CNR2X1 U1905 ( .A(n1480), .B(n608), .Z(n1431) );
  CND2X2 U1906 ( .A(n2088), .B(n2080), .Z(n1423) );
  CNIVX4 U1907 ( .A(n1416), .Z(n1965) );
  CND2X1 U1908 ( .A(n1965), .B(n588), .Z(n1419) );
  CND2XL U1909 ( .A(n1417), .B(n1425), .Z(n1418) );
  CND2X1 U1910 ( .A(n1419), .B(n1418), .Z(n2090) );
  CND2X1 U1911 ( .A(n1420), .B(n1961), .Z(n1481) );
  CIVX2 U1912 ( .A(n1481), .Z(n2476) );
  CND2X1 U1913 ( .A(n2090), .B(n2476), .Z(n1422) );
  CND2X1 U1914 ( .A(n2092), .B(n2087), .Z(n1421) );
  CND3X2 U1915 ( .A(n1421), .B(n1423), .C(n1422), .Z(n1433) );
  COND2X2 U1916 ( .A(acc2[42]), .B(n1431), .C(n1433), .D(n1424), .Z(n1468) );
  CND2X2 U1917 ( .A(n1427), .B(n1961), .Z(n2057) );
  CND2X1 U1918 ( .A(n2053), .B(n2087), .Z(n1428) );
  CND3X2 U1919 ( .A(n1430), .B(n1429), .C(n1428), .Z(n1437) );
  CENX2 U1920 ( .A(n2632), .B(n1437), .Z(n1469) );
  CENX1 U1921 ( .A(acc2[42]), .B(n1431), .Z(n1432) );
  CENX2 U1922 ( .A(n1433), .B(n1432), .Z(n1466) );
  CNR2X2 U1923 ( .A(n1466), .B(n1467), .Z(n1535) );
  CNR2X2 U1924 ( .A(n1529), .B(n1535), .Z(n2100) );
  CND2X2 U1925 ( .A(n1526), .B(n2100), .Z(n1974) );
  CENX1 U1926 ( .A(acc2[44]), .B(n1435), .Z(n1436) );
  CENX2 U1927 ( .A(n540), .B(n1436), .Z(n1471) );
  CAN2X2 U1928 ( .A(n1437), .B(acc2[43]), .Z(n1470) );
  CNR2X2 U1929 ( .A(n1471), .B(n1470), .Z(n1514) );
  CNR2XL U1930 ( .A(n1974), .B(n1514), .Z(n1473) );
  CNR2X4 U1931 ( .A(n1439), .B(n1438), .Z(n1447) );
  CNR2X2 U1932 ( .A(n1447), .B(n1440), .Z(n1451) );
  CND2X2 U1933 ( .A(n1441), .B(n1451), .Z(n1454) );
  CND2X2 U1934 ( .A(n1457), .B(n1443), .Z(n1460) );
  CANR1X2 U1935 ( .A(n1445), .B(n446), .C(n1444), .Z(n1459) );
  COND1X2 U1936 ( .A(n1448), .B(n1447), .C(n1446), .Z(n1449) );
  CANR1X2 U1937 ( .A(n1451), .B(n1450), .C(n1449), .Z(n1452) );
  COND1X2 U1938 ( .A(n1454), .B(n1453), .C(n1452), .Z(n1455) );
  CANR1X2 U1939 ( .A(n1457), .B(n1456), .C(n1455), .Z(n1458) );
  COND1X2 U1940 ( .A(n1460), .B(n1459), .C(n1458), .Z(n1461) );
  CIVX4 U1941 ( .A(n1461), .Z(n2182) );
  CIVX8 U1942 ( .A(n2182), .Z(n2269) );
  CND2X2 U1943 ( .A(n1463), .B(n1462), .Z(n1546) );
  CND2X2 U1944 ( .A(n1465), .B(n1464), .Z(n1545) );
  COND1X4 U1945 ( .A(n1546), .B(n1544), .C(n1545), .Z(n2101) );
  CND2X2 U1946 ( .A(n1467), .B(n1466), .Z(n1533) );
  COND1X2 U1947 ( .A(n1533), .B(n1529), .C(n1530), .Z(n2102) );
  CANR1X2 U1948 ( .A(n2101), .B(n2100), .C(n2102), .Z(n1477) );
  CND2X2 U1949 ( .A(n1471), .B(n1470), .Z(n1515) );
  COND1XL U1950 ( .A(n1514), .B(n1477), .C(n1515), .Z(n1472) );
  CANR1X2 U1951 ( .A(n1473), .B(n2269), .C(n1472), .Z(n1474) );
  CIVX2 U1952 ( .A(x[45]), .Z(n1476) );
  COND1X2 U1953 ( .A(n1479), .B(n1515), .C(n1478), .Z(n2109) );
  CNR2X2 U1954 ( .A(n1480), .B(n2003), .Z(n1500) );
  CENX1 U1955 ( .A(acc2[46]), .B(n1500), .Z(n1485) );
  CND2X1 U1956 ( .A(n1964), .B(n2080), .Z(n1483) );
  CNR2X2 U1957 ( .A(n1481), .B(n588), .Z(n2488) );
  CND2X1 U1958 ( .A(n2488), .B(n1965), .Z(n1482) );
  CAN2X2 U1959 ( .A(n1486), .B(acc2[45]), .Z(n1487) );
  CND2X2 U1960 ( .A(n1488), .B(n1487), .Z(n2111) );
  CIVX2 U1961 ( .A(n1974), .Z(n1518) );
  CND2X2 U1962 ( .A(n1518), .B(n1973), .Z(n1508) );
  CIVX2 U1963 ( .A(n1508), .Z(n1496) );
  CNR2IX2 U1964 ( .B(n1491), .A(n1496), .Z(n1490) );
  CIVX2 U1965 ( .A(n2269), .Z(n1494) );
  CIVX2 U1966 ( .A(n1491), .Z(n1495) );
  CND2X2 U1967 ( .A(n1494), .B(n1493), .Z(n1498) );
  CND2X1 U1968 ( .A(n2269), .B(n606), .Z(n1497) );
  CND3X2 U1969 ( .A(n1499), .B(n1498), .C(n1497), .Z(n1566) );
  CND2X2 U1970 ( .A(n1566), .B(x[46]), .Z(n1573) );
  CIVX1 U1971 ( .A(x[47]), .Z(n1522) );
  CND2X1 U1972 ( .A(n1958), .B(n2080), .Z(n1504) );
  CND2X1 U1973 ( .A(n1960), .B(n2087), .Z(n1503) );
  CND2X1 U1974 ( .A(n1501), .B(n1962), .Z(n1502) );
  CIVXL U1975 ( .A(n2112), .Z(n1507) );
  CND2X1 U1976 ( .A(n1505), .B(n1506), .Z(n2110) );
  CAN2X2 U1977 ( .A(n1507), .B(n2110), .Z(n1513) );
  COND1X2 U1978 ( .A(n1972), .B(n1509), .C(n2111), .Z(n1510) );
  CANR1X4 U1979 ( .A(n1511), .B(n2269), .C(n1510), .Z(n1512) );
  CENX4 U1980 ( .A(n1513), .B(n1512), .Z(n1567) );
  CIVXL U1981 ( .A(n1514), .Z(n1516) );
  CAN2X1 U1982 ( .A(n1516), .B(n1515), .Z(n1520) );
  CANR1X2 U1983 ( .A(n1518), .B(n2269), .C(n1517), .Z(n1519) );
  CENX2 U1984 ( .A(n1520), .B(n1519), .Z(n2584) );
  CIVX2 U1985 ( .A(x[44]), .Z(n1521) );
  COND2X2 U1986 ( .A(n1522), .B(n1567), .C(n2584), .D(n1521), .Z(n1523) );
  CIVXL U1987 ( .A(n1535), .Z(n1525) );
  CND2X1 U1988 ( .A(n1525), .B(n1533), .Z(n1528) );
  CIVX2 U1989 ( .A(n1526), .Z(n1532) );
  CIVX2 U1990 ( .A(n448), .Z(n1534) );
  COAN1X1 U1991 ( .A(n1532), .B(n2182), .C(n1534), .Z(n1527) );
  CEOX2 U1992 ( .A(n1528), .B(n1527), .Z(n1561) );
  CNR2IX1 U1993 ( .B(x[42]), .A(n1561), .Z(n1541) );
  CIVXL U1994 ( .A(n1529), .Z(n1531) );
  CAN2X1 U1995 ( .A(n1531), .B(n1530), .Z(n1539) );
  CNR2X1 U1996 ( .A(n1532), .B(n1535), .Z(n1537) );
  COND1X1 U1997 ( .A(n1535), .B(n1534), .C(n1533), .Z(n1536) );
  CNR2IX1 U1998 ( .B(x[43]), .A(n1560), .Z(n1540) );
  CNR2X2 U1999 ( .A(n1541), .B(n1540), .Z(n1559) );
  CNIVX4 U2000 ( .A(n2269), .Z(n2329) );
  CIVX2 U2001 ( .A(n1542), .Z(n1548) );
  CND2X1 U2002 ( .A(n1548), .B(n1546), .Z(n1543) );
  CEOX2 U2003 ( .A(n2329), .B(n1543), .Z(n2558) );
  CIVX2 U2004 ( .A(n1546), .Z(n1547) );
  CANR1X4 U2005 ( .A(n1548), .B(n2269), .C(n1547), .Z(n1552) );
  CENX2 U2006 ( .A(n1553), .B(n1552), .Z(n2543) );
  CND2X2 U2007 ( .A(n2543), .B(x[41]), .Z(n1551) );
  CIVDX2 U2008 ( .A(n1551), .Z0(n1557), .Z1(n1549) );
  CIVXL U2009 ( .A(x[41]), .Z(n1554) );
  CND2X1 U2010 ( .A(n1555), .B(n1554), .Z(n1556) );
  COND11X2 U2011 ( .A(x[40]), .B(n2558), .C(n1557), .D(n1556), .Z(n1558) );
  CND2X2 U2012 ( .A(n1558), .B(n1559), .Z(n1565) );
  CIVX2 U2013 ( .A(n1561), .Z(n2504) );
  CANR3X2 U2014 ( .A(n2574), .B(x[43]), .C(n2504), .D(x[42]), .Z(n1563) );
  CNR2X2 U2015 ( .A(n1563), .B(n1562), .Z(n1564) );
  CND2X2 U2016 ( .A(n1565), .B(n1564), .Z(n1582) );
  CNR2IX4 U2017 ( .B(x[47]), .A(n1567), .Z(n1574) );
  CNR3X2 U2018 ( .A(n1566), .B(x[46]), .C(n1574), .Z(n1569) );
  CNR2X2 U2019 ( .A(n2562), .B(x[47]), .Z(n1568) );
  CNR2X4 U2020 ( .A(n1569), .B(n1568), .Z(n1580) );
  CIVX2 U2021 ( .A(n1570), .Z(n2557) );
  CNR2X1 U2022 ( .A(n2557), .B(x[45]), .Z(n1578) );
  CND2IX1 U2023 ( .B(x[44]), .A(n2584), .Z(n1571) );
  CNR2X2 U2024 ( .A(n1572), .B(n1571), .Z(n1577) );
  CIVX2 U2025 ( .A(n1573), .Z(n1575) );
  CNR2X2 U2026 ( .A(n1575), .B(n1574), .Z(n1576) );
  COND1X2 U2027 ( .A(n1578), .B(n1577), .C(n1576), .Z(n1579) );
  CND2X2 U2028 ( .A(n1579), .B(n1580), .Z(n1581) );
  CANR1X2 U2029 ( .A(n1583), .B(n1582), .C(n1581), .Z(n1584) );
  COND1X2 U2030 ( .A(n1585), .B(n1957), .C(n1584), .Z(n2338) );
  CIVX4 U2031 ( .A(n446), .Z(n1813) );
  COND1X1 U2032 ( .A(n1591), .B(n1813), .C(n602), .Z(n1590) );
  CIVX2 U2033 ( .A(n1588), .Z(n1601) );
  CND2X1 U2034 ( .A(n1601), .B(n1592), .Z(n1589) );
  CENX1 U2035 ( .A(n1590), .B(n1589), .Z(n1682) );
  CIVX2 U2036 ( .A(n1682), .Z(n2539) );
  CND2X1 U2037 ( .A(n1612), .B(n1601), .Z(n1595) );
  CIVXL U2038 ( .A(n1592), .Z(n1593) );
  CANR1X1 U2039 ( .A(n1601), .B(n597), .C(n1593), .Z(n1594) );
  COND1X2 U2040 ( .A(n1595), .B(n1813), .C(n1594), .Z(n1598) );
  CND2X1 U2041 ( .A(n1600), .B(n1596), .Z(n1597) );
  CENX2 U2042 ( .A(n1598), .B(n1597), .Z(n1599) );
  CNR2IX2 U2043 ( .B(x[21]), .A(n1599), .Z(n1684) );
  CNR3X2 U2044 ( .A(n2539), .B(n1684), .C(x[20]), .Z(n1624) );
  CIVX2 U2045 ( .A(n1599), .Z(n2578) );
  CNR2X1 U2046 ( .A(n2578), .B(x[21]), .Z(n1623) );
  CND2X2 U2047 ( .A(n1601), .B(n1600), .Z(n1611) );
  CNR2X1 U2048 ( .A(n1611), .B(n1617), .Z(n1604) );
  CND2X1 U2049 ( .A(n1604), .B(n1612), .Z(n1606) );
  CIVX2 U2050 ( .A(n436), .Z(n1602) );
  COND1X1 U2051 ( .A(n1617), .B(n1602), .C(n1618), .Z(n1603) );
  CANR1X1 U2052 ( .A(n1604), .B(n597), .C(n1603), .Z(n1605) );
  COND1X2 U2053 ( .A(n1606), .B(n1813), .C(n1605), .Z(n1610) );
  CND2X1 U2054 ( .A(n535), .B(n1608), .Z(n1609) );
  CENX2 U2055 ( .A(n1610), .B(n1609), .Z(n1627) );
  CNR2IX2 U2056 ( .B(x[23]), .A(n1627), .Z(n1626) );
  CIVX2 U2057 ( .A(n1611), .Z(n1614) );
  CND2XL U2058 ( .A(n1612), .B(n1614), .Z(n1616) );
  CANR1X1 U2059 ( .A(n1614), .B(n597), .C(n436), .Z(n1615) );
  COND1X2 U2060 ( .A(n1616), .B(n1813), .C(n1615), .Z(n1621) );
  CIVXL U2061 ( .A(n1617), .Z(n1619) );
  CND2X1 U2062 ( .A(n1619), .B(n1618), .Z(n1620) );
  CENX2 U2063 ( .A(n1621), .B(n1620), .Z(n1625) );
  CNR2IX2 U2064 ( .B(x[22]), .A(n1625), .Z(n1622) );
  CNR2X2 U2065 ( .A(n1626), .B(n1622), .Z(n1686) );
  COND1X1 U2066 ( .A(n1624), .B(n1623), .C(n1686), .Z(n1631) );
  CIVX2 U2067 ( .A(n1625), .Z(n2544) );
  CNR3X2 U2068 ( .A(n2544), .B(x[22]), .C(n1626), .Z(n1629) );
  CIVX2 U2069 ( .A(n1627), .Z(n2527) );
  CNR2X1 U2070 ( .A(n2527), .B(x[23]), .Z(n1628) );
  CNR2X1 U2071 ( .A(n1629), .B(n1628), .Z(n1630) );
  CND2X1 U2072 ( .A(n1631), .B(n1630), .Z(n1689) );
  CIVX2 U2073 ( .A(n1632), .Z(n1635) );
  CND2X1 U2074 ( .A(n1656), .B(n1635), .Z(n1637) );
  CND2X1 U2075 ( .A(n525), .B(n1643), .Z(n1634) );
  CANR1XL U2076 ( .A(n1635), .B(n1659), .C(n1634), .Z(n1636) );
  COND1X2 U2077 ( .A(n1637), .B(n1813), .C(n1636), .Z(n1642) );
  CIVXL U2078 ( .A(n1638), .Z(n1640) );
  CND2X1 U2079 ( .A(n1640), .B(n1639), .Z(n1641) );
  CENX2 U2080 ( .A(n1642), .B(n1641), .Z(n1677) );
  CNR2IX2 U2081 ( .B(x[19]), .A(n1677), .Z(n1679) );
  CND2X1 U2082 ( .A(n1644), .B(n1643), .Z(n1651) );
  CANR1XL U2083 ( .A(n1655), .B(n1659), .C(n1645), .Z(n1649) );
  CND2XL U2084 ( .A(n1656), .B(n1655), .Z(n1647) );
  CND2X2 U2085 ( .A(n1649), .B(n1648), .Z(n1650) );
  CENX2 U2086 ( .A(n1651), .B(n1650), .Z(n2534) );
  CNR2IX1 U2087 ( .B(x[18]), .A(n2534), .Z(n1652) );
  CNR2X2 U2088 ( .A(n1679), .B(n1652), .Z(n1831) );
  CIVX2 U2089 ( .A(n1813), .Z(n1658) );
  CIVDX4 U2090 ( .A(n1653), .Z0(n1645), .Z1(n1654) );
  CND2X1 U2091 ( .A(n1655), .B(n1654), .Z(n1660) );
  CIVX2 U2092 ( .A(n1660), .Z(n1663) );
  CIVXL U2093 ( .A(n1656), .Z(n1664) );
  CNR2IX1 U2094 ( .B(n1663), .A(n1664), .Z(n1657) );
  CND2X2 U2095 ( .A(n1658), .B(n1657), .Z(n1668) );
  CIVXL U2096 ( .A(n1659), .Z(n1661) );
  CAN2X1 U2097 ( .A(n1661), .B(n1660), .Z(n1665) );
  CIVX1 U2098 ( .A(n1661), .Z(n1662) );
  CANR2X2 U2099 ( .A(n1665), .B(n1664), .C(n1663), .D(n1662), .Z(n1667) );
  CND3X2 U2100 ( .A(n1668), .B(n1667), .C(n1666), .Z(n2525) );
  CIVX2 U2101 ( .A(n2525), .Z(n1669) );
  CNR2IX2 U2102 ( .B(x[17]), .A(n1669), .Z(n1830) );
  CIVX1 U2103 ( .A(x[16]), .Z(n1675) );
  CND2X2 U2104 ( .A(n1829), .B(n1675), .Z(n1676) );
  COND2X2 U2105 ( .A(x[17]), .B(n2525), .C(n1830), .D(n1676), .Z(n1681) );
  CIVX2 U2106 ( .A(n1677), .Z(n2538) );
  COND2X2 U2107 ( .A(x[19]), .B(n2538), .C(n1679), .D(n1678), .Z(n1680) );
  CANR1X2 U2108 ( .A(n1831), .B(n1681), .C(n1680), .Z(n1687) );
  CNR2IX2 U2109 ( .B(x[20]), .A(n1682), .Z(n1683) );
  CNR2X2 U2110 ( .A(n1684), .B(n1683), .Z(n1685) );
  CND2X2 U2111 ( .A(n1686), .B(n1685), .Z(n1834) );
  CNR2X2 U2112 ( .A(n1687), .B(n1834), .Z(n1688) );
  CNR2X1 U2113 ( .A(n1689), .B(n1688), .Z(n1913) );
  CND2X1 U2114 ( .A(n529), .B(n1690), .Z(n1696) );
  CAOR1X2 U2115 ( .A(n1693), .B(n1752), .C(n1692), .Z(n1737) );
  CIVX2 U2116 ( .A(n1706), .Z(n1694) );
  CANR1X2 U2117 ( .A(n1707), .B(n1737), .C(n1694), .Z(n1695) );
  CENX2 U2118 ( .A(n1696), .B(n1695), .Z(n2536) );
  CND2X1 U2119 ( .A(n2536), .B(x[10]), .Z(n1705) );
  CND2X1 U2120 ( .A(n1698), .B(n1697), .Z(n1704) );
  CIVX2 U2121 ( .A(n1699), .Z(n1702) );
  CNIVX1 U2122 ( .A(n1700), .Z(n1701) );
  CANR1X4 U2123 ( .A(n1702), .B(n1737), .C(n1701), .Z(n1703) );
  CND2X1 U2124 ( .A(n1707), .B(n1706), .Z(n1708) );
  CENX2 U2125 ( .A(n1737), .B(n1708), .Z(n2550) );
  CIVXL U2126 ( .A(x[9]), .Z(n1709) );
  CND2XL U2127 ( .A(n2550), .B(n1709), .Z(n1719) );
  CIVXL U2128 ( .A(n1710), .Z(n1712) );
  CAN2X1 U2129 ( .A(n1712), .B(n1711), .Z(n1716) );
  CIVX2 U2130 ( .A(n1752), .Z(n1745) );
  COAN1XL U2131 ( .A(n1714), .B(n1745), .C(n1713), .Z(n1715) );
  CENX2 U2132 ( .A(n1716), .B(n1715), .Z(n2505) );
  CNR2IX2 U2133 ( .B(x[9]), .A(n2550), .Z(n1800) );
  CNR2X2 U2134 ( .A(n1800), .B(x[8]), .Z(n1717) );
  CND2X2 U2135 ( .A(n2505), .B(n1717), .Z(n1718) );
  CIVX2 U2136 ( .A(n2536), .Z(n1721) );
  CIVX1 U2137 ( .A(x[10]), .Z(n1720) );
  CND3X2 U2138 ( .A(n1722), .B(n1721), .C(n1720), .Z(n1725) );
  CIVX1 U2139 ( .A(x[11]), .Z(n1723) );
  CND2IX1 U2140 ( .B(n2522), .A(n1723), .Z(n1724) );
  CIVX2 U2141 ( .A(n1726), .Z(n1728) );
  CND2X1 U2142 ( .A(n1728), .B(n1727), .Z(n1733) );
  CANR1X1 U2143 ( .A(n1731), .B(n1737), .C(n1730), .Z(n1732) );
  CIVX2 U2144 ( .A(n1734), .Z(n1736) );
  CND2X2 U2145 ( .A(n1736), .B(n1735), .Z(n1740) );
  CANR1X1 U2146 ( .A(n1738), .B(n1737), .C(n526), .Z(n1739) );
  CIVX2 U2147 ( .A(n1743), .Z(n1748) );
  CIVDX2 U2148 ( .A(n1744), .Z0(n1750), .Z1(n1746) );
  COND1X2 U2149 ( .A(n1746), .B(n1745), .C(n528), .Z(n1747) );
  CENX2 U2150 ( .A(n1748), .B(n1747), .Z(n2540) );
  CNR2IX2 U2151 ( .B(x[7]), .A(n2540), .Z(n1787) );
  CND2XL U2152 ( .A(n1750), .B(n1749), .Z(n1751) );
  CENX1 U2153 ( .A(n1752), .B(n1751), .Z(n2563) );
  CNR2IX1 U2154 ( .B(x[6]), .A(n2563), .Z(n1753) );
  CNR2X2 U2155 ( .A(n1787), .B(n1753), .Z(n1793) );
  CND2X1 U2156 ( .A(n1758), .B(n1757), .Z(n1760) );
  CENX1 U2157 ( .A(n1760), .B(n1759), .Z(n1770) );
  CNR2IX1 U2158 ( .B(x[3]), .A(n1770), .Z(n1769) );
  CNR2X1 U2159 ( .A(n600), .B(x[0]), .Z(n1767) );
  CIVX2 U2160 ( .A(x[1]), .Z(n1766) );
  CND2X1 U2161 ( .A(n1763), .B(n1762), .Z(n1765) );
  CENX1 U2162 ( .A(n1765), .B(n1764), .Z(n2572) );
  CANR5CXL U2163 ( .A(n1767), .B(n1766), .C(n2572), .Z(n1768) );
  CANR3X2 U2164 ( .A(x[2]), .B(n593), .C(n1769), .D(n1768), .Z(n1773) );
  CNR3X1 U2165 ( .A(n1769), .B(x[2]), .C(n593), .Z(n1772) );
  CIVX2 U2166 ( .A(n1770), .Z(n2571) );
  CNR2X1 U2167 ( .A(n2571), .B(x[3]), .Z(n1771) );
  CNR3X2 U2168 ( .A(n1773), .B(n1772), .C(n1771), .Z(n1776) );
  CND2X1 U2169 ( .A(n1780), .B(n1782), .Z(n1774) );
  CENX1 U2170 ( .A(n1774), .B(n1779), .Z(n2567) );
  CNR2IX1 U2171 ( .B(x[4]), .A(n2567), .Z(n1775) );
  CNR2X2 U2172 ( .A(n1776), .B(n1775), .Z(n1783) );
  CNIVX1 U2173 ( .A(n1779), .Z(n1781) );
  CNR2IX1 U2174 ( .B(x[5]), .A(n1790), .Z(n1791) );
  CNR2IX1 U2175 ( .B(n1783), .A(n1791), .Z(n1784) );
  CND2X1 U2176 ( .A(n1793), .B(n1784), .Z(n1785) );
  CIVX2 U2177 ( .A(n1785), .Z(n1798) );
  COAN1X1 U2178 ( .A(n1788), .B(n1787), .C(n1786), .Z(n1796) );
  CIVX1 U2179 ( .A(x[4]), .Z(n1789) );
  CND2X1 U2180 ( .A(n2567), .B(n1789), .Z(n1792) );
  CIVX2 U2181 ( .A(n1790), .Z(n2582) );
  COND2X1 U2182 ( .A(n1792), .B(n1791), .C(n2582), .D(x[5]), .Z(n1794) );
  CND2X2 U2183 ( .A(n1794), .B(n1793), .Z(n1795) );
  CND2X2 U2184 ( .A(n1796), .B(n1795), .Z(n1797) );
  CNR2X2 U2185 ( .A(n1798), .B(n1797), .Z(n1802) );
  CNR2IX1 U2186 ( .B(x[8]), .A(n2505), .Z(n1799) );
  COR2X1 U2187 ( .A(n1800), .B(n1799), .Z(n1801) );
  CNR2X2 U2188 ( .A(n1802), .B(n1801), .Z(n1805) );
  CIVX2 U2189 ( .A(n1803), .Z(n1804) );
  CND2XL U2190 ( .A(n1806), .B(n1807), .Z(n1811) );
  COND1X2 U2191 ( .A(n450), .B(n1813), .C(n1812), .Z(n1810) );
  CENX2 U2192 ( .A(n1811), .B(n1810), .Z(n2541) );
  CAN2XL U2193 ( .A(n451), .B(n1812), .Z(n1814) );
  CENX1 U2194 ( .A(n1814), .B(n1813), .Z(n2529) );
  CNR2IX1 U2195 ( .B(x[14]), .A(n2529), .Z(n1815) );
  CIVX2 U2196 ( .A(n1816), .Z(n2548) );
  CIVX1 U2197 ( .A(x[12]), .Z(n1817) );
  CND2X1 U2198 ( .A(n2518), .B(n1817), .Z(n1818) );
  COND2X1 U2199 ( .A(x[13]), .B(n2548), .C(n1819), .D(n1818), .Z(n1825) );
  CIVX1 U2200 ( .A(x[14]), .Z(n1820) );
  CND2X1 U2201 ( .A(n2529), .B(n1820), .Z(n1823) );
  CANR1X1 U2202 ( .A(n1826), .B(n1825), .C(n1824), .Z(n1827) );
  CND2X2 U2203 ( .A(n1828), .B(n1827), .Z(n1836) );
  CIVX2 U2204 ( .A(n1829), .Z(n2545) );
  CANR1X2 U2205 ( .A(x[16]), .B(n2545), .C(n1830), .Z(n1832) );
  CND2X1 U2206 ( .A(n1832), .B(n1831), .Z(n1833) );
  CND2X2 U2207 ( .A(n1836), .B(n1835), .Z(n1912) );
  CIVXL U2208 ( .A(n1837), .Z(n1839) );
  CAN2X1 U2209 ( .A(n1839), .B(n1838), .Z(n1851) );
  CANR1X2 U2210 ( .A(n1843), .B(n1885), .C(n1842), .Z(n1865) );
  CANR1X2 U2211 ( .A(n1846), .B(n1845), .C(n1844), .Z(n1856) );
  COND1X1 U2212 ( .A(n1847), .B(n1856), .C(n1853), .Z(n1848) );
  CANR1X2 U2213 ( .A(n1849), .B(n1904), .C(n1848), .Z(n1850) );
  CENX2 U2214 ( .A(n1851), .B(n1850), .Z(n1937) );
  CIVX4 U2215 ( .A(n1937), .Z(n2555) );
  CND2X4 U2216 ( .A(n2555), .B(x[31]), .Z(n1861) );
  CND2X1 U2217 ( .A(n1854), .B(n1853), .Z(n1860) );
  CIVX2 U2218 ( .A(n1855), .Z(n1858) );
  CIVX2 U2219 ( .A(n1856), .Z(n1857) );
  CANR1X4 U2220 ( .A(n1858), .B(n1904), .C(n1857), .Z(n1859) );
  CEOX2 U2221 ( .A(n1860), .B(n1859), .Z(n1935) );
  CIVX2 U2222 ( .A(n1935), .Z(n2553) );
  CND2X4 U2223 ( .A(n2553), .B(x[30]), .Z(n1925) );
  CND2X4 U2224 ( .A(n1861), .B(n1925), .Z(n1881) );
  CIVX2 U2225 ( .A(n1863), .Z(n1931) );
  CIVDX1 U2226 ( .A(n1864), .Z0(n1841), .Z1(n1868) );
  CND2X2 U2227 ( .A(n1904), .B(n1841), .Z(n1866) );
  CND2X4 U2228 ( .A(n1866), .B(n1870), .Z(n1930) );
  CENX2 U2229 ( .A(n1863), .B(n1930), .Z(n2533) );
  CND2X2 U2230 ( .A(n2533), .B(x[28]), .Z(n1880) );
  CNR2X1 U2231 ( .A(n1868), .B(n1871), .Z(n1873) );
  COND1X1 U2232 ( .A(n1871), .B(n1870), .C(n1869), .Z(n1872) );
  CANR1X2 U2233 ( .A(n1873), .B(n1904), .C(n1872), .Z(n1878) );
  CIVXL U2234 ( .A(n1874), .Z(n1876) );
  CAN2X1 U2235 ( .A(n1876), .B(n1875), .Z(n1877) );
  CENX2 U2236 ( .A(n1878), .B(n1877), .Z(n1929) );
  CIVX3 U2237 ( .A(n1933), .Z(n1879) );
  CND2X4 U2238 ( .A(n1880), .B(n1879), .Z(n1927) );
  CNR2X4 U2239 ( .A(n1881), .B(n1927), .Z(n1910) );
  CIVXL U2240 ( .A(n1882), .Z(n1884) );
  CAN2X1 U2241 ( .A(n1884), .B(n1883), .Z(n1889) );
  COND1XL U2242 ( .A(n1890), .B(n590), .C(n1891), .Z(n1886) );
  CANR1X2 U2243 ( .A(n1887), .B(n1904), .C(n1886), .Z(n1888) );
  CENX2 U2244 ( .A(n1889), .B(n1888), .Z(n1920) );
  CNR2IX2 U2245 ( .B(x[27]), .A(n1920), .Z(n1919) );
  CIVX2 U2246 ( .A(n1890), .Z(n1892) );
  CAN2X1 U2247 ( .A(n1892), .B(n1891), .Z(n1895) );
  CANR1X1 U2248 ( .A(n1893), .B(n1904), .C(n591), .Z(n1894) );
  CENX1 U2249 ( .A(n1895), .B(n1894), .Z(n1918) );
  CNR2IX2 U2250 ( .B(x[26]), .A(n1918), .Z(n1896) );
  CNR2X2 U2251 ( .A(n1919), .B(n1896), .Z(n1924) );
  CIVX2 U2252 ( .A(n1897), .Z(n1905) );
  CNIVX4 U2253 ( .A(n1904), .Z(n1898) );
  CND2X2 U2254 ( .A(n2566), .B(x[24]), .Z(n1908) );
  CIVXL U2255 ( .A(n1900), .Z(n1902) );
  CAN2X1 U2256 ( .A(n1902), .B(n1901), .Z(n1907) );
  CANR1X1 U2257 ( .A(n1905), .B(n1904), .C(n1903), .Z(n1906) );
  CENX2 U2258 ( .A(n1907), .B(n1906), .Z(n1914) );
  CNR2IX2 U2259 ( .B(x[25]), .A(n1914), .Z(n1917) );
  CNR2IX2 U2260 ( .B(n1908), .A(n1917), .Z(n1909) );
  CND3X2 U2261 ( .A(n1910), .B(n1924), .C(n1909), .Z(n1911) );
  CANR1X2 U2262 ( .A(n1913), .B(n1912), .C(n1911), .Z(n1948) );
  CIVX2 U2263 ( .A(n1914), .Z(n2514) );
  CIVXL U2264 ( .A(x[24]), .Z(n1915) );
  COND2X2 U2265 ( .A(x[25]), .B(n2514), .C(n1917), .D(n1916), .Z(n1923) );
  CIVX2 U2266 ( .A(n1918), .Z(n2512) );
  CNR3X2 U2267 ( .A(n2512), .B(x[26]), .C(n1919), .Z(n1922) );
  CIVX2 U2268 ( .A(n1920), .Z(n2510) );
  CNR2X1 U2269 ( .A(n2510), .B(x[27]), .Z(n1921) );
  CANR3X2 U2270 ( .A(n1924), .B(n1923), .C(n1922), .D(n1921), .Z(n1946) );
  CND2X2 U2271 ( .A(n2555), .B(x[31]), .Z(n1926) );
  CND2X2 U2272 ( .A(n1926), .B(n1925), .Z(n1928) );
  COR2X1 U2273 ( .A(n1928), .B(n1927), .Z(n1945) );
  CIVX2 U2274 ( .A(n1928), .Z(n1943) );
  CIVXL U2275 ( .A(n1929), .Z(n2546) );
  COND2X1 U2276 ( .A(x[29]), .B(n2546), .C(n1933), .D(n1932), .Z(n1942) );
  CIVX1 U2277 ( .A(x[30]), .Z(n1934) );
  CND2XL U2278 ( .A(n1935), .B(n1934), .Z(n1940) );
  CIVX2 U2279 ( .A(x[31]), .Z(n1936) );
  CND2X1 U2280 ( .A(n1937), .B(n1936), .Z(n1938) );
  COND1X2 U2281 ( .A(n1940), .B(n1939), .C(n1938), .Z(n1941) );
  CANR1X2 U2282 ( .A(n1943), .B(n1942), .C(n1941), .Z(n1944) );
  COND1X2 U2283 ( .A(n1946), .B(n1945), .C(n1944), .Z(n1947) );
  CNR2X2 U2284 ( .A(n1948), .B(n1947), .Z(n1956) );
  CNR2IX1 U2285 ( .B(x[32]), .A(n1949), .Z(n1951) );
  CNR2X2 U2286 ( .A(n1951), .B(n1950), .Z(n1953) );
  CND3X2 U2287 ( .A(n1954), .B(n1953), .C(n1952), .Z(n1955) );
  CIVX8 U2288 ( .A(n1959), .Z(n2091) );
  CND2X2 U2289 ( .A(n2026), .B(n1961), .Z(n2089) );
  CNR2X4 U2290 ( .A(n2089), .B(n588), .Z(n2485) );
  CND2X1 U2291 ( .A(n1963), .B(n2091), .Z(n1966) );
  CND2X4 U2292 ( .A(n1967), .B(n1980), .Z(n2096) );
  COR2X1 U2293 ( .A(n1969), .B(n1968), .Z(n1971) );
  CND2X1 U2294 ( .A(n1969), .B(n1968), .Z(n1970) );
  CAN2X2 U2295 ( .A(n1971), .B(n1970), .Z(n2168) );
  CND2X4 U2296 ( .A(n2108), .B(n1973), .Z(n2105) );
  CNR2X4 U2297 ( .A(n2105), .B(n1974), .Z(n2330) );
  CNR2X2 U2298 ( .A(n1977), .B(n1976), .Z(n1991) );
  CND2X2 U2299 ( .A(n1981), .B(n1980), .Z(n2035) );
  CNR2X2 U2300 ( .A(n2035), .B(n1982), .Z(n1985) );
  CNR2X4 U2301 ( .A(n2133), .B(n2134), .Z(n2274) );
  CENX1 U2302 ( .A(acc2[52]), .B(n1985), .Z(n1987) );
  CENX2 U2303 ( .A(n1987), .B(n1986), .Z(n2132) );
  CND2X2 U2304 ( .A(n1988), .B(n2026), .Z(n1994) );
  CND2X1 U2305 ( .A(n1991), .B(n1990), .Z(n1992) );
  CND3X2 U2306 ( .A(n1994), .B(n1993), .C(n1992), .Z(n2034) );
  CNR2X2 U2307 ( .A(n2132), .B(n2131), .Z(n2276) );
  CNR2X2 U2308 ( .A(n2276), .B(n2274), .Z(n2265) );
  CNR2X2 U2309 ( .A(n2035), .B(n2003), .Z(n2006) );
  CENX1 U2310 ( .A(acc2[54]), .B(n2006), .Z(n2004) );
  CENX2 U2311 ( .A(n2004), .B(n2007), .Z(n2137) );
  CAN2X2 U2312 ( .A(n2005), .B(acc2[53]), .Z(n2136) );
  CNR2X2 U2313 ( .A(n2137), .B(n2136), .Z(n2261) );
  COND1X2 U2314 ( .A(acc2[54]), .B(n2007), .C(n2006), .Z(n2009) );
  CND2X2 U2315 ( .A(n2009), .B(n2008), .Z(n2139) );
  CANR2X2 U2316 ( .A(n2012), .B(n2026), .C(n2011), .D(n2091), .Z(n2013) );
  CNR2X4 U2317 ( .A(n2139), .B(n2138), .Z(n2247) );
  CNR2X2 U2318 ( .A(n2261), .B(n2247), .Z(n2135) );
  CND2X2 U2319 ( .A(n2265), .B(n2135), .Z(n2129) );
  CNR2X2 U2320 ( .A(n608), .B(n2035), .Z(n2032) );
  CENX2 U2321 ( .A(n2032), .B(acc2[50]), .Z(n2024) );
  COND11X2 U2322 ( .A(n2019), .B(n2018), .C(n2017), .D(n2080), .Z(n2022) );
  CND2X1 U2323 ( .A(n2020), .B(n2091), .Z(n2021) );
  CND3X2 U2324 ( .A(n2022), .B(n2023), .C(n2021), .Z(n2033) );
  CANR2X2 U2325 ( .A(n2027), .B(n2026), .C(n2091), .D(n2025), .Z(n2031) );
  CHA1X1 U2326 ( .A(acc2[51]), .B(n2034), .CO(n2131), .S(n2119) );
  CNR2X2 U2327 ( .A(n2035), .B(n421), .Z(n2043) );
  CENX1 U2328 ( .A(acc2[48]), .B(n2043), .Z(n2041) );
  CENX2 U2329 ( .A(n2041), .B(n2044), .Z(n2122) );
  CNR2X2 U2330 ( .A(n2122), .B(n2123), .Z(n2324) );
  CENX2 U2331 ( .A(n2042), .B(n2602), .Z(n2125) );
  CNR2X4 U2332 ( .A(n2125), .B(n2124), .Z(n2314) );
  CNR2X2 U2333 ( .A(n2314), .B(n2324), .Z(n2308) );
  CND2X2 U2334 ( .A(n2126), .B(n2308), .Z(n2285) );
  CNR2X4 U2335 ( .A(n2129), .B(n2285), .Z(n2239) );
  CND2X4 U2336 ( .A(n2330), .B(n2239), .Z(n2237) );
  CNR2X1 U2337 ( .A(n610), .B(n2096), .Z(n2058) );
  CENX1 U2338 ( .A(acc2[60]), .B(n2058), .Z(n2051) );
  CND2X1 U2339 ( .A(n2045), .B(n2087), .Z(n2050) );
  CND2X1 U2340 ( .A(n2046), .B(n2091), .Z(n2049) );
  CND2IX1 U2341 ( .B(n2047), .A(n2485), .Z(n2048) );
  CND3X2 U2342 ( .A(n2050), .B(n2049), .C(n2048), .Z(n2059) );
  CND2X1 U2343 ( .A(n2052), .B(n2087), .Z(n2055) );
  CND2X1 U2344 ( .A(n2053), .B(n2091), .Z(n2054) );
  CNR2X2 U2345 ( .A(n2155), .B(n2154), .Z(n2181) );
  COND1X2 U2346 ( .A(acc2[60]), .B(n2059), .C(n2058), .Z(n2061) );
  CND2X2 U2347 ( .A(n2061), .B(n2060), .Z(n2157) );
  CANR2X1 U2348 ( .A(n2062), .B(n2087), .C(n2485), .D(n1408), .Z(n2065) );
  CND2X1 U2349 ( .A(n2063), .B(n2091), .Z(n2064) );
  CND2X1 U2350 ( .A(n2065), .B(n2064), .Z(n2066) );
  CNR2X2 U2351 ( .A(n2157), .B(n2156), .Z(n2189) );
  CNR2X2 U2352 ( .A(n2181), .B(n2189), .Z(n2172) );
  CHA1X1 U2353 ( .A(acc2[61]), .B(n2066), .CO(n2158), .S(n2156) );
  COR2X2 U2354 ( .A(n2159), .B(n2158), .Z(n2170) );
  CND2X1 U2355 ( .A(n2172), .B(n2170), .Z(n2162) );
  CAN2X1 U2356 ( .A(n2067), .B(n2091), .Z(n2068) );
  CANR1X2 U2357 ( .A(n2087), .B(n2069), .C(n2068), .Z(n2073) );
  CIVX2 U2358 ( .A(n2070), .Z(n2071) );
  CND2X2 U2359 ( .A(n2071), .B(n2080), .Z(n2072) );
  CND2X4 U2360 ( .A(n2073), .B(n2072), .Z(n2077) );
  CNR2X2 U2361 ( .A(n2096), .B(n421), .Z(n2076) );
  CENX1 U2362 ( .A(acc2[56]), .B(n2076), .Z(n2075) );
  CENX2 U2363 ( .A(n2077), .B(n2075), .Z(n2145) );
  CNR2X2 U2364 ( .A(n2145), .B(n2144), .Z(n2234) );
  COND1X2 U2365 ( .A(acc2[56]), .B(n2077), .C(n2076), .Z(n2079) );
  CND2X2 U2366 ( .A(n2079), .B(n2078), .Z(n2146) );
  CND2X1 U2367 ( .A(n2081), .B(n2080), .Z(n2086) );
  CND2X1 U2368 ( .A(n2082), .B(n2087), .Z(n2085) );
  CND2X1 U2369 ( .A(n2083), .B(n2091), .Z(n2084) );
  CND3X2 U2370 ( .A(n2086), .B(n2085), .C(n2084), .Z(n2097) );
  CNR2X2 U2371 ( .A(n2146), .B(n2147), .Z(n2227) );
  CNR2X2 U2372 ( .A(n2234), .B(n2227), .Z(n2218) );
  CIVX2 U2373 ( .A(n2089), .Z(n2498) );
  CND2X1 U2374 ( .A(n2090), .B(n2498), .Z(n2094) );
  CND2X1 U2375 ( .A(n2092), .B(n2091), .Z(n2093) );
  CHA1X1 U2376 ( .A(acc2[57]), .B(n2097), .CO(n2148), .S(n2147) );
  CND2X2 U2377 ( .A(n2218), .B(n2153), .Z(n2184) );
  COR2X1 U2378 ( .A(n2162), .B(n2184), .Z(n2164) );
  CNR2X1 U2379 ( .A(n2237), .B(n2164), .Z(n2166) );
  CND2X2 U2380 ( .A(n2101), .B(n2100), .Z(n2104) );
  CIVX2 U2381 ( .A(n2102), .Z(n2103) );
  CND2X2 U2382 ( .A(n2104), .B(n2103), .Z(n2107) );
  CIVX4 U2383 ( .A(n2105), .Z(n2106) );
  CND2X4 U2384 ( .A(n2107), .B(n2106), .Z(n2116) );
  CND2X2 U2385 ( .A(n2109), .B(n2108), .Z(n2114) );
  COAN1X1 U2386 ( .A(n2112), .B(n2111), .C(n2110), .Z(n2113) );
  CAN2X2 U2387 ( .A(n2114), .B(n2113), .Z(n2115) );
  CND2X4 U2388 ( .A(n2116), .B(n2115), .Z(n2327) );
  CND2X2 U2389 ( .A(n2118), .B(n2117), .Z(n2306) );
  CND2X1 U2390 ( .A(n2120), .B(n2119), .Z(n2294) );
  CND2X2 U2391 ( .A(n2123), .B(n2122), .Z(n2325) );
  CND2X2 U2392 ( .A(n2124), .B(n2125), .Z(n2315) );
  COND1X2 U2393 ( .A(n2325), .B(n2314), .C(n2315), .Z(n2309) );
  CND2X2 U2394 ( .A(n2309), .B(n2126), .Z(n2127) );
  CND2X4 U2395 ( .A(n2127), .B(n2128), .Z(n2250) );
  CIVX4 U2396 ( .A(n2129), .Z(n2130) );
  CND2X4 U2397 ( .A(n2250), .B(n2130), .Z(n2143) );
  CND2X2 U2398 ( .A(n2132), .B(n2131), .Z(n2282) );
  COND1X2 U2399 ( .A(n2282), .B(n2274), .C(n2275), .Z(n2251) );
  CAN2X2 U2400 ( .A(n2135), .B(n2251), .Z(n2141) );
  CND2X2 U2401 ( .A(n2137), .B(n2136), .Z(n2262) );
  CND2X1 U2402 ( .A(n2139), .B(n2138), .Z(n2248) );
  COND1X1 U2403 ( .A(n2247), .B(n2262), .C(n2248), .Z(n2140) );
  CNR2X4 U2404 ( .A(n2141), .B(n2140), .Z(n2142) );
  CND2X4 U2405 ( .A(n2143), .B(n2142), .Z(n2238) );
  CANR1X4 U2406 ( .A(n2239), .B(n2327), .C(n2238), .Z(n2230) );
  CND2X2 U2407 ( .A(n2145), .B(n2144), .Z(n2235) );
  CND2X2 U2408 ( .A(n2147), .B(n2146), .Z(n2228) );
  COND1X2 U2409 ( .A(n2235), .B(n2227), .C(n2228), .Z(n2219) );
  CND2X2 U2410 ( .A(n2149), .B(n2148), .Z(n2216) );
  COND1X2 U2411 ( .A(n2205), .B(n2216), .C(n2206), .Z(n2152) );
  CND2X2 U2412 ( .A(n2155), .B(n2154), .Z(n2193) );
  CND2X1 U2413 ( .A(n2157), .B(n2156), .Z(n2190) );
  COND1X2 U2414 ( .A(n2189), .B(n2193), .C(n2190), .Z(n2171) );
  CND2X2 U2415 ( .A(n2159), .B(n2158), .Z(n2169) );
  CIVX2 U2416 ( .A(n2169), .Z(n2160) );
  CANR1X1 U2417 ( .A(n2170), .B(n2171), .C(n2160), .Z(n2161) );
  COAN1X1 U2418 ( .A(n2183), .B(n2162), .C(n2161), .Z(n2163) );
  COND1X1 U2419 ( .A(n2164), .B(n2230), .C(n2163), .Z(n2165) );
  CANR1X2 U2420 ( .A(n2166), .B(n2269), .C(n2165), .Z(n2167) );
  CENX2 U2421 ( .A(n2168), .B(n2167), .Z(n2407) );
  CND2X4 U2422 ( .A(n2511), .B(x[63]), .Z(n2406) );
  CND2X2 U2423 ( .A(n2170), .B(n2169), .Z(n2179) );
  CIVX2 U2424 ( .A(n2184), .Z(n2192) );
  CND2X1 U2425 ( .A(n2192), .B(n2172), .Z(n2174) );
  CIVX2 U2426 ( .A(n2183), .Z(n2195) );
  CANR1X1 U2427 ( .A(n2172), .B(n2195), .C(n2171), .Z(n2173) );
  COAN1X1 U2428 ( .A(n2174), .B(n2230), .C(n2173), .Z(n2177) );
  CNR2X1 U2429 ( .A(n2237), .B(n2174), .Z(n2175) );
  CND2X2 U2430 ( .A(n2176), .B(n2177), .Z(n2178) );
  CENX2 U2431 ( .A(n2179), .B(n2178), .Z(n2405) );
  CND2X4 U2432 ( .A(n2180), .B(n2406), .Z(n2397) );
  CIVX2 U2433 ( .A(n2181), .Z(n2196) );
  CND2X2 U2434 ( .A(n2196), .B(n2193), .Z(n2188) );
  CNR2X1 U2435 ( .A(n2237), .B(n2184), .Z(n2186) );
  CIVX4 U2436 ( .A(n2182), .Z(n2319) );
  COND1X1 U2437 ( .A(n2184), .B(n2230), .C(n2183), .Z(n2185) );
  CANR1X2 U2438 ( .A(n2186), .B(n2319), .C(n2185), .Z(n2187) );
  CENX2 U2439 ( .A(n2188), .B(n2187), .Z(n2399) );
  CND2X2 U2440 ( .A(n2521), .B(x[60]), .Z(n2203) );
  CIVX2 U2441 ( .A(n2189), .Z(n2191) );
  CAN2X1 U2442 ( .A(n2191), .B(n2190), .Z(n2202) );
  CND2X1 U2443 ( .A(n2192), .B(n2196), .Z(n2198) );
  CIVX2 U2444 ( .A(n2193), .Z(n2194) );
  COAN1X1 U2445 ( .A(n2198), .B(n2230), .C(n2197), .Z(n2199) );
  CND2X2 U2446 ( .A(n2200), .B(n2199), .Z(n2201) );
  CND2X2 U2447 ( .A(n2203), .B(n2398), .Z(n2204) );
  CNR2X4 U2448 ( .A(n2397), .B(n2204), .Z(n2377) );
  CIVX2 U2449 ( .A(n2205), .Z(n2207) );
  CAN2X2 U2450 ( .A(n2207), .B(n2206), .Z(n2215) );
  CND2X1 U2451 ( .A(n2218), .B(n2217), .Z(n2212) );
  CNR2X2 U2452 ( .A(n2237), .B(n2212), .Z(n2209) );
  CIVX2 U2453 ( .A(n2216), .Z(n2210) );
  CANR1X1 U2454 ( .A(n2217), .B(n2219), .C(n2210), .Z(n2211) );
  COAN1X1 U2455 ( .A(n2212), .B(n2230), .C(n2211), .Z(n2213) );
  CND2X1 U2456 ( .A(n2217), .B(n2216), .Z(n2225) );
  CIVX1 U2457 ( .A(n2218), .Z(n2221) );
  CNR2X1 U2458 ( .A(n2237), .B(n2221), .Z(n2223) );
  CIVX2 U2459 ( .A(n2219), .Z(n2220) );
  COND1X1 U2460 ( .A(n2221), .B(n2230), .C(n2220), .Z(n2222) );
  CANR1X2 U2461 ( .A(n2223), .B(n2319), .C(n2222), .Z(n2224) );
  CEOX2 U2462 ( .A(n2225), .B(n2224), .Z(n2387) );
  CND2X2 U2463 ( .A(n2570), .B(x[58]), .Z(n2226) );
  CND2X2 U2464 ( .A(n2388), .B(n2226), .Z(n2378) );
  CIVX1 U2465 ( .A(n2227), .Z(n2229) );
  CAN2X2 U2466 ( .A(n2229), .B(n2228), .Z(n2233) );
  CND2X2 U2467 ( .A(n604), .B(n2231), .Z(n2232) );
  CENX2 U2468 ( .A(n2233), .B(n2232), .Z(n2581) );
  CND2X2 U2469 ( .A(n2581), .B(x[57]), .Z(n2381) );
  CIVX1 U2470 ( .A(n2234), .Z(n2236) );
  CND2X2 U2471 ( .A(n2236), .B(n2235), .Z(n2243) );
  CIVX2 U2472 ( .A(n2237), .Z(n2241) );
  CAOR1XL U2473 ( .A(n2327), .B(n2239), .C(n2238), .Z(n2240) );
  CANR1X2 U2474 ( .A(n2241), .B(n2319), .C(n2240), .Z(n2242) );
  CEOX2 U2475 ( .A(n2243), .B(n2242), .Z(n2380) );
  CIVX2 U2476 ( .A(n2380), .Z(n2513) );
  CND2X2 U2477 ( .A(n2513), .B(x[56]), .Z(n2244) );
  CND2X2 U2478 ( .A(n2381), .B(n2244), .Z(n2245) );
  CNR2X2 U2479 ( .A(n2378), .B(n2245), .Z(n2246) );
  CND2X2 U2480 ( .A(n2377), .B(n2246), .Z(n2339) );
  CIVX2 U2481 ( .A(n2247), .Z(n2249) );
  CAN2X2 U2482 ( .A(n2249), .B(n2248), .Z(n2260) );
  CIVX3 U2483 ( .A(n2330), .Z(n2318) );
  CIVX2 U2484 ( .A(n2285), .Z(n2277) );
  CND2X1 U2485 ( .A(n2254), .B(n2277), .Z(n2256) );
  CNR2X1 U2486 ( .A(n2318), .B(n2256), .Z(n2258) );
  CIVX4 U2487 ( .A(n2327), .Z(n2317) );
  CIVX2 U2488 ( .A(n2250), .Z(n2284) );
  CIVX2 U2489 ( .A(n2284), .Z(n2278) );
  CNIVX2 U2490 ( .A(n2251), .Z(n2264) );
  CIVX2 U2491 ( .A(n2264), .Z(n2252) );
  COND1XL U2492 ( .A(n2261), .B(n2252), .C(n2262), .Z(n2253) );
  CANR1X1 U2493 ( .A(n2278), .B(n2254), .C(n2253), .Z(n2255) );
  COND1X1 U2494 ( .A(n2317), .B(n2256), .C(n2255), .Z(n2257) );
  CANR1X2 U2495 ( .A(n2258), .B(n2319), .C(n2257), .Z(n2259) );
  CENX2 U2496 ( .A(n2260), .B(n2259), .Z(n2368) );
  CIVX1 U2497 ( .A(n2261), .Z(n2263) );
  CAN2X2 U2498 ( .A(n2263), .B(n2262), .Z(n2272) );
  CND2X1 U2499 ( .A(n2265), .B(n2277), .Z(n2267) );
  CNR2X1 U2500 ( .A(n2318), .B(n2267), .Z(n2270) );
  CANR1X1 U2501 ( .A(n2265), .B(n2278), .C(n2264), .Z(n2266) );
  COND1X1 U2502 ( .A(n2267), .B(n2317), .C(n2266), .Z(n2268) );
  CAOR1X1 U2503 ( .A(n2270), .B(n2269), .C(n2268), .Z(n2271) );
  CEOX2 U2504 ( .A(n2272), .B(n2271), .Z(n2365) );
  CIVX2 U2505 ( .A(n2365), .Z(n2559) );
  CND2X2 U2506 ( .A(n2559), .B(x[54]), .Z(n2273) );
  CIVX2 U2507 ( .A(n2276), .Z(n2283) );
  CND2X1 U2508 ( .A(n2277), .B(n2283), .Z(n2279) );
  CNR2X1 U2509 ( .A(n2318), .B(n2279), .Z(n2281) );
  CAN2X1 U2510 ( .A(n2283), .B(n2282), .Z(n2289) );
  CNR2X1 U2511 ( .A(n2318), .B(n2285), .Z(n2287) );
  COND1XL U2512 ( .A(n2285), .B(n2317), .C(n2284), .Z(n2286) );
  CENX2 U2513 ( .A(n2289), .B(n2288), .Z(n2517) );
  CND2X2 U2514 ( .A(n2517), .B(x[52]), .Z(n2290) );
  CND2X4 U2515 ( .A(n2358), .B(n2290), .Z(n2291) );
  CNR2X4 U2516 ( .A(n2356), .B(n2291), .Z(n2355) );
  CIVX2 U2517 ( .A(n434), .Z(n2307) );
  CND2X1 U2518 ( .A(n2308), .B(n2307), .Z(n2297) );
  CNR2X2 U2519 ( .A(n2318), .B(n2297), .Z(n2302) );
  CIVX2 U2520 ( .A(n2301), .Z(n2298) );
  CIVX2 U2521 ( .A(n2319), .Z(n2299) );
  CIVXL U2522 ( .A(n2306), .Z(n2295) );
  CANR1XL U2523 ( .A(n2307), .B(n2309), .C(n2295), .Z(n2296) );
  COND1X2 U2524 ( .A(n2297), .B(n2317), .C(n2296), .Z(n2300) );
  CNR2X2 U2525 ( .A(n2300), .B(n2298), .Z(n2303) );
  CND2IX1 U2526 ( .B(n2301), .A(n2300), .Z(n2305) );
  CIVX2 U2527 ( .A(n2302), .Z(n2304) );
  CIVX2 U2528 ( .A(n2308), .Z(n2311) );
  CNR2X1 U2529 ( .A(n2318), .B(n2311), .Z(n2313) );
  CIVXL U2530 ( .A(n2309), .Z(n2310) );
  COND1X2 U2531 ( .A(n2311), .B(n2317), .C(n2310), .Z(n2312) );
  CIVXL U2532 ( .A(n2314), .Z(n2316) );
  CND2X1 U2533 ( .A(n2316), .B(n2315), .Z(n2323) );
  COND1XL U2534 ( .A(n2324), .B(n2317), .C(n2325), .Z(n2321) );
  CND2IX2 U2535 ( .B(n2321), .A(n2320), .Z(n2322) );
  CIVXL U2536 ( .A(n2324), .Z(n2326) );
  CND2X2 U2537 ( .A(n2326), .B(n2325), .Z(n2332) );
  CANR1X4 U2538 ( .A(n447), .B(n2329), .C(n2328), .Z(n2331) );
  CNR2IX1 U2539 ( .B(x[48]), .A(n2583), .Z(n2333) );
  CNR3X2 U2540 ( .A(n2354), .B(n2343), .C(n2333), .Z(n2334) );
  COND1X2 U2541 ( .A(n2338), .B(n2337), .C(n2336), .Z(n2421) );
  CIVX2 U2542 ( .A(n2339), .Z(n2419) );
  CIVXL U2543 ( .A(x[48]), .Z(n2340) );
  CND2X2 U2544 ( .A(n2583), .B(n2340), .Z(n2344) );
  CIVXL U2545 ( .A(x[49]), .Z(n2341) );
  COAN1X1 U2546 ( .A(n2344), .B(n2343), .C(n2342), .Z(n2353) );
  CIVX2 U2547 ( .A(n2528), .Z(n2346) );
  CIVX2 U2548 ( .A(x[51]), .Z(n2345) );
  CND2X1 U2549 ( .A(n2346), .B(n2345), .Z(n2351) );
  CIVX1 U2550 ( .A(x[50]), .Z(n2347) );
  CAN3X2 U2551 ( .A(n2349), .B(n2348), .C(n2347), .Z(n2350) );
  CNR2IX2 U2552 ( .B(n2351), .A(n2350), .Z(n2352) );
  CIVX2 U2553 ( .A(n2356), .Z(n2374) );
  CIVXL U2554 ( .A(x[52]), .Z(n2357) );
  CND2IX1 U2555 ( .B(n2517), .A(n2357), .Z(n2363) );
  CIVX2 U2556 ( .A(n2358), .Z(n2362) );
  CIVXL U2557 ( .A(x[53]), .Z(n2359) );
  CND2X1 U2558 ( .A(n2360), .B(n2359), .Z(n2361) );
  COND1X2 U2559 ( .A(n2363), .B(n2362), .C(n2361), .Z(n2373) );
  CIVXL U2560 ( .A(x[54]), .Z(n2364) );
  CND2X1 U2561 ( .A(n2365), .B(n2364), .Z(n2371) );
  CIVX2 U2562 ( .A(n2366), .Z(n2370) );
  CIVX1 U2563 ( .A(x[55]), .Z(n2367) );
  CND2X1 U2564 ( .A(n2368), .B(n2367), .Z(n2369) );
  COND1X2 U2565 ( .A(n2371), .B(n2370), .C(n2369), .Z(n2372) );
  CANR1X2 U2566 ( .A(n2374), .B(n2373), .C(n2372), .Z(n2375) );
  CND2X4 U2567 ( .A(n2376), .B(n2375), .Z(n2418) );
  CIVX2 U2568 ( .A(n2377), .Z(n2416) );
  CIVX2 U2569 ( .A(n2378), .Z(n2396) );
  CIVXL U2570 ( .A(x[56]), .Z(n2379) );
  CND2X1 U2571 ( .A(n2380), .B(n2379), .Z(n2386) );
  CIVX2 U2572 ( .A(n2381), .Z(n2385) );
  CIVX2 U2573 ( .A(n2581), .Z(n2383) );
  CIVX1 U2574 ( .A(x[57]), .Z(n2382) );
  CND2X2 U2575 ( .A(n2383), .B(n2382), .Z(n2384) );
  COND1X2 U2576 ( .A(n2386), .B(n2385), .C(n2384), .Z(n2395) );
  CIVDX2 U2577 ( .A(n2387), .Z0(n2570), .Z1(n2390) );
  CIVX1 U2578 ( .A(x[58]), .Z(n2389) );
  CIVX1 U2579 ( .A(x[59]), .Z(n2391) );
  CND2IX2 U2580 ( .B(n2508), .A(n2391), .Z(n2392) );
  CANR1X2 U2581 ( .A(n2396), .B(n2395), .C(n2394), .Z(n2415) );
  CIVX2 U2582 ( .A(n2397), .Z(n2413) );
  CIVX2 U2583 ( .A(n2398), .Z(n2403) );
  CIVDX2 U2584 ( .A(n2399), .Z0(n2401), .Z1(n2521) );
  CIVXL U2585 ( .A(x[60]), .Z(n2400) );
  CND2X1 U2586 ( .A(n2401), .B(n2400), .Z(n2402) );
  COND2X2 U2587 ( .A(x[61]), .B(n2515), .C(n2403), .D(n2402), .Z(n2412) );
  CIVXL U2588 ( .A(x[62]), .Z(n2404) );
  CIVX2 U2589 ( .A(n2406), .Z(n2409) );
  COND1X2 U2590 ( .A(n2410), .B(n2409), .C(n2408), .Z(n2411) );
  CANR1X2 U2591 ( .A(n2413), .B(n2412), .C(n2411), .Z(n2414) );
  COND1X2 U2592 ( .A(n2416), .B(n2415), .C(n2414), .Z(n2417) );
  CANR1X4 U2593 ( .A(n2419), .B(n2418), .C(n2417), .Z(n2420) );
  CND2X4 U2594 ( .A(n2421), .B(n2420), .Z(n2422) );
  CIVX8 U2595 ( .A(n2472), .Z(n2530) );
  CIVX2 U2596 ( .A(acc[2]), .Z(n2423) );
  COND1X1 U2597 ( .A(n2424), .B(n2530), .C(n2423), .Z(n2683) );
  CND2X1 U2598 ( .A(n2488), .B(n2491), .Z(n2426) );
  CIVX2 U2599 ( .A(acc[15]), .Z(n2425) );
  COND1X1 U2600 ( .A(n2426), .B(n2530), .C(n2425), .Z(n2670) );
  CND2X1 U2601 ( .A(n2498), .B(n2588), .Z(n2428) );
  CIVX8 U2602 ( .A(n2472), .Z(n2526) );
  CIVX2 U2603 ( .A(acc[24]), .Z(n2427) );
  COND1X1 U2604 ( .A(n2428), .B(n2526), .C(n2427), .Z(n2687) );
  CIVX2 U2605 ( .A(n2437), .Z(n2481) );
  CIVX2 U2606 ( .A(n2429), .Z(n2464) );
  CND2X1 U2607 ( .A(n2481), .B(n2464), .Z(n2431) );
  CIVX2 U2608 ( .A(acc[17]), .Z(n2430) );
  COND1X1 U2609 ( .A(n2431), .B(n2526), .C(n2430), .Z(n2664) );
  CND2X1 U2610 ( .A(n2485), .B(n2491), .Z(n2432) );
  COND1X1 U2611 ( .A(n2432), .B(n2526), .C(n453), .Z(n2678) );
  CND2X1 U2612 ( .A(n2488), .B(n2484), .Z(n2434) );
  CIVX2 U2613 ( .A(acc[14]), .Z(n2433) );
  COND1X1 U2614 ( .A(n2434), .B(n2530), .C(n2433), .Z(n2668) );
  CND2X1 U2615 ( .A(n2471), .B(n2491), .Z(n2436) );
  CIVX2 U2616 ( .A(acc[3]), .Z(n2435) );
  COND1X1 U2617 ( .A(n2436), .B(n2530), .C(n2435), .Z(n2684) );
  CNR2X1 U2618 ( .A(n2437), .B(n588), .Z(n2494) );
  CND2IX1 U2619 ( .B(n1982), .A(n2494), .Z(n2439) );
  CIVX2 U2620 ( .A(acc[22]), .Z(n2438) );
  COND1X1 U2621 ( .A(n2439), .B(n2530), .C(n2438), .Z(n2672) );
  CND2X1 U2622 ( .A(n2476), .B(n2440), .Z(n2442) );
  CIVX2 U2623 ( .A(acc[11]), .Z(n2441) );
  COND1X1 U2624 ( .A(n2442), .B(n2526), .C(n2441), .Z(n2661) );
  CND2X1 U2625 ( .A(n2488), .B(n609), .Z(n2444) );
  COND1X1 U2626 ( .A(n2444), .B(n2530), .C(n2443), .Z(n2669) );
  CND2X1 U2627 ( .A(n601), .B(n609), .Z(n2446) );
  COND1X1 U2628 ( .A(n2446), .B(n2526), .C(n2445), .Z(n2681) );
  CND2X1 U2629 ( .A(n2485), .B(n724), .Z(n2448) );
  COND1X1 U2630 ( .A(n2448), .B(n2526), .C(n2447), .Z(n2675) );
  CND2X1 U2631 ( .A(n2586), .B(n2449), .Z(n2451) );
  CIVX8 U2632 ( .A(n2472), .Z(n2585) );
  CIVX2 U2633 ( .A(acc[0]), .Z(n2450) );
  COND1X1 U2634 ( .A(n2451), .B(n2585), .C(n2450), .Z(n297) );
  CND2X1 U2635 ( .A(n2476), .B(n2588), .Z(n2453) );
  CIVX8 U2636 ( .A(n2472), .Z(n2580) );
  CIVX1 U2637 ( .A(acc[8]), .Z(n2452) );
  COND1X1 U2638 ( .A(n2453), .B(n2580), .C(n2452), .Z(n2688) );
  CND2X1 U2639 ( .A(n2494), .B(n609), .Z(n2455) );
  CIVX2 U2640 ( .A(acc[21]), .Z(n2454) );
  COND1X1 U2641 ( .A(n2455), .B(n2585), .C(n2454), .Z(n2673) );
  CND2XL U2642 ( .A(n2485), .B(n609), .Z(n2457) );
  CIVX2 U2643 ( .A(acc[29]), .Z(n2456) );
  COND1X1 U2644 ( .A(n2457), .B(n2585), .C(n2456), .Z(n2677) );
  CND2X1 U2645 ( .A(n2494), .B(n2491), .Z(n2459) );
  CIVX8 U2646 ( .A(n2472), .Z(n2577) );
  CIVX2 U2647 ( .A(acc[23]), .Z(n2458) );
  COND1X1 U2648 ( .A(n2459), .B(n2577), .C(n2458), .Z(n2674) );
  CND2X1 U2649 ( .A(n2476), .B(n2464), .Z(n2461) );
  COND1X1 U2650 ( .A(n2461), .B(n2580), .C(n2460), .Z(n2666) );
  CND2X1 U2651 ( .A(n2498), .B(n2440), .Z(n2463) );
  CIVX2 U2652 ( .A(acc[27]), .Z(n2462) );
  COND1X1 U2653 ( .A(n2463), .B(n2585), .C(n2462), .Z(n2663) );
  CND2X1 U2654 ( .A(n2498), .B(n2464), .Z(n2466) );
  CIVX2 U2655 ( .A(acc[25]), .Z(n2465) );
  COND1X1 U2656 ( .A(n2466), .B(n2577), .C(n2465), .Z(n2665) );
  CND2X1 U2657 ( .A(n2481), .B(n2440), .Z(n2468) );
  CIVX2 U2658 ( .A(acc[19]), .Z(n2467) );
  COND1X1 U2659 ( .A(n2468), .B(n2577), .C(n2467), .Z(n2662) );
  CND2X1 U2660 ( .A(n2481), .B(n2588), .Z(n2470) );
  COND1X1 U2661 ( .A(n2470), .B(n2580), .C(n454), .Z(n2686) );
  CND2X1 U2662 ( .A(n2471), .B(n609), .Z(n2474) );
  CIVX8 U2663 ( .A(n2472), .Z(n2573) );
  COND1X1 U2664 ( .A(n2474), .B(n2573), .C(n2473), .Z(n2685) );
  CAN2X1 U2665 ( .A(n864), .B(n588), .Z(n2497) );
  CND2X1 U2666 ( .A(n2476), .B(n2497), .Z(n2478) );
  COND1X1 U2667 ( .A(n2478), .B(n2577), .C(n2477), .Z(n2658) );
  CND2X1 U2668 ( .A(n601), .B(n2484), .Z(n2480) );
  CIVX2 U2669 ( .A(acc[6]), .Z(n2479) );
  COND1X1 U2670 ( .A(n2480), .B(n2573), .C(n2479), .Z(n2680) );
  CND2X1 U2671 ( .A(n2481), .B(n2497), .Z(n2483) );
  CIVX2 U2672 ( .A(acc[18]), .Z(n2482) );
  COND1X1 U2673 ( .A(n2483), .B(n2573), .C(n2482), .Z(n2659) );
  CND2XL U2674 ( .A(n2485), .B(n2484), .Z(n2487) );
  CIVX1 U2675 ( .A(acc[30]), .Z(n2486) );
  COND1X1 U2676 ( .A(n2487), .B(n2580), .C(n2486), .Z(n2676) );
  CND2X1 U2677 ( .A(n2488), .B(n724), .Z(n2490) );
  CIVX2 U2678 ( .A(acc[12]), .Z(n2489) );
  COND1X1 U2679 ( .A(n2490), .B(n2577), .C(n2489), .Z(n2667) );
  CND2X1 U2680 ( .A(n601), .B(n2491), .Z(n2493) );
  COND1X1 U2681 ( .A(n2493), .B(n2573), .C(n2492), .Z(n2682) );
  CND2X1 U2682 ( .A(n2494), .B(n724), .Z(n2496) );
  COND1X1 U2683 ( .A(n2496), .B(n2573), .C(n2495), .Z(n2671) );
  CND2X1 U2684 ( .A(n2498), .B(n2497), .Z(n2500) );
  CIVX2 U2685 ( .A(acc[26]), .Z(n2499) );
  COND1X1 U2686 ( .A(n2500), .B(n2585), .C(n2499), .Z(n2660) );
  CND2X1 U2687 ( .A(n601), .B(n724), .Z(n2503) );
  CIVX2 U2688 ( .A(acc[4]), .Z(n2502) );
  COND1X1 U2689 ( .A(n2503), .B(n2580), .C(n2502), .Z(n2679) );
  CMXI2X1 U2690 ( .A0(n2504), .A1(n2633), .S(n2530), .Z(n371) );
  CIVX2 U2691 ( .A(n2505), .Z(n2506) );
  CMXI2X1 U2692 ( .A0(n2506), .A1(n2601), .S(n2526), .Z(n337) );
  CMXI2X1 U2693 ( .A0(n2507), .A1(n2636), .S(n2530), .Z(n367) );
  CMXI2X1 U2694 ( .A0(n542), .A1(n2619), .S(n2530), .Z(n388) );
  CIVXL U2695 ( .A(acc2[27]), .Z(n2509) );
  CMXI2X1 U2696 ( .A0(n2510), .A1(n2509), .S(n2526), .Z(n356) );
  CMXI2X1 U2697 ( .A0(n2511), .A1(n2615), .S(n2526), .Z(n392) );
  CMXI2X1 U2698 ( .A0(n2512), .A1(n2642), .S(n2530), .Z(n355) );
  CMXI2X1 U2699 ( .A0(n2513), .A1(n2622), .S(n2530), .Z(n385) );
  CMXI2X1 U2700 ( .A0(n2514), .A1(n2607), .S(n2526), .Z(n354) );
  CMXI2X1 U2701 ( .A0(n2515), .A1(n2617), .S(n2526), .Z(n390) );
  CMXI2X1 U2702 ( .A0(n2516), .A1(n2606), .S(n2530), .Z(n368) );
  CMXI2X1 U2703 ( .A0(n2517), .A1(n2625), .S(n2530), .Z(n381) );
  CIVX2 U2704 ( .A(n2518), .Z(n2520) );
  CIVXL U2705 ( .A(acc2[12]), .Z(n2519) );
  CMXI2X1 U2706 ( .A0(n2520), .A1(n2519), .S(n2526), .Z(n341) );
  CMXI2X1 U2707 ( .A0(n2521), .A1(n2618), .S(n2526), .Z(n389) );
  CMXI2X1 U2708 ( .A0(n2522), .A1(n2649), .S(n2530), .Z(n340) );
  CMXI2X1 U2709 ( .A0(n2523), .A1(n2616), .S(n2526), .Z(n391) );
  CIVXL U2710 ( .A(acc2[17]), .Z(n2524) );
  CMXI2X1 U2711 ( .A0(n2525), .A1(n2524), .S(n2526), .Z(n346) );
  CMXI2X1 U2712 ( .A0(n2527), .A1(n2604), .S(n2526), .Z(n352) );
  CMXI2X1 U2713 ( .A0(n2528), .A1(n2626), .S(n2530), .Z(n380) );
  CIVX2 U2714 ( .A(n2529), .Z(n2531) );
  CMXI2X1 U2715 ( .A0(n2531), .A1(n2592), .S(n2530), .Z(n343) );
  CMXI2X1 U2716 ( .A0(n2532), .A1(n2640), .S(n2577), .Z(n361) );
  CMXI2X1 U2717 ( .A0(n2533), .A1(n2596), .S(n2577), .Z(n357) );
  CIVXL U2718 ( .A(n2534), .Z(n2535) );
  CMXI2X1 U2719 ( .A0(n2535), .A1(n2645), .S(n2580), .Z(n347) );
  CMXI2X1 U2720 ( .A0(n2536), .A1(n2650), .S(n2577), .Z(n339) );
  CIVXL U2721 ( .A(acc2[19]), .Z(n2537) );
  CMXI2X1 U2722 ( .A0(n2538), .A1(n2537), .S(n2573), .Z(n348) );
  CMXI2X1 U2723 ( .A0(n2539), .A1(n2594), .S(n2580), .Z(n349) );
  CMXI2X1 U2724 ( .A0(n2542), .A1(n2637), .S(n2573), .Z(n365) );
  CMXI2X1 U2725 ( .A0(n2543), .A1(n2634), .S(n2585), .Z(n370) );
  CMXI2X1 U2726 ( .A0(n2544), .A1(n2643), .S(n2585), .Z(n351) );
  CMXI2X1 U2727 ( .A0(n1566), .A1(n2630), .S(n2577), .Z(n375) );
  CMXI2X1 U2728 ( .A0(n2545), .A1(n2646), .S(n2577), .Z(n345) );
  CMXI2X1 U2729 ( .A0(n2546), .A1(n2641), .S(n2580), .Z(n358) );
  CMXI2X1 U2730 ( .A0(n2547), .A1(n2639), .S(n2573), .Z(n363) );
  CMXI2X1 U2731 ( .A0(n2548), .A1(n2648), .S(n2573), .Z(n342) );
  CMXI2X1 U2732 ( .A0(n2549), .A1(n2598), .S(n2585), .Z(n366) );
  CIVX2 U2733 ( .A(n2550), .Z(n2552) );
  CIVX1 U2734 ( .A(acc2[9]), .Z(n2551) );
  CMXI2X1 U2735 ( .A0(n2552), .A1(n2551), .S(n2580), .Z(n338) );
  CMXI2X1 U2736 ( .A0(n2553), .A1(n2591), .S(n2573), .Z(n359) );
  CIVXL U2737 ( .A(acc2[31]), .Z(n2554) );
  CMXI2X1 U2738 ( .A0(n449), .A1(n2554), .S(n2573), .Z(n360) );
  CMXI2X1 U2739 ( .A0(n600), .A1(n2656), .S(n2573), .Z(n329) );
  CMXI2X1 U2740 ( .A0(n2556), .A1(n2609), .S(n2580), .Z(n362) );
  CMXI2X1 U2741 ( .A0(n2557), .A1(n2593), .S(n2573), .Z(n374) );
  CMXI2X1 U2742 ( .A0(n2558), .A1(n2635), .S(n2577), .Z(n369) );
  CMXI2X1 U2743 ( .A0(n2559), .A1(n2624), .S(n2577), .Z(n383) );
  CIVXL U2744 ( .A(n2560), .Z(n2561) );
  CMXI2X1 U2745 ( .A0(n2561), .A1(n2602), .S(n2585), .Z(n378) );
  CMXI2X1 U2746 ( .A0(n2562), .A1(n2629), .S(n2577), .Z(n376) );
  CIVX2 U2747 ( .A(n2563), .Z(n2564) );
  CMXI2X1 U2748 ( .A0(n2564), .A1(n2652), .S(n2585), .Z(n335) );
  CMXI2X1 U2749 ( .A0(n2565), .A1(n2597), .S(n2577), .Z(n382) );
  CMXI2X1 U2750 ( .A0(n2566), .A1(n2595), .S(n2585), .Z(n353) );
  CIVX2 U2751 ( .A(n2567), .Z(n2569) );
  CIVXL U2752 ( .A(acc2[4]), .Z(n2568) );
  CMXI2X1 U2753 ( .A0(n2569), .A1(n2568), .S(n2577), .Z(n333) );
  CMXI2X1 U2754 ( .A0(n2570), .A1(n2620), .S(n2573), .Z(n387) );
  CMXI2X1 U2755 ( .A0(n2571), .A1(n2653), .S(n2580), .Z(n332) );
  CMXI2X1 U2756 ( .A0(n2574), .A1(n2632), .S(n2580), .Z(n372) );
  CMXI2X1 U2757 ( .A0(n2575), .A1(n2638), .S(n2585), .Z(n364) );
  CMXI2X1 U2758 ( .A0(n2576), .A1(n2623), .S(n2580), .Z(n384) );
  CMXI2X1 U2759 ( .A0(n2578), .A1(n2644), .S(n2577), .Z(n350) );
  CMXI2X1 U2760 ( .A0(n2579), .A1(n2627), .S(n2580), .Z(n379) );
  CMXI2X1 U2761 ( .A0(n593), .A1(n2654), .S(n2580), .Z(n331) );
  CMXI2X1 U2762 ( .A0(n2581), .A1(n2621), .S(n2585), .Z(n386) );
  CMXI2X1 U2763 ( .A0(n2582), .A1(n2605), .S(n2585), .Z(n334) );
  CMXI2X1 U2764 ( .A0(n536), .A1(n2628), .S(n2585), .Z(n377) );
  CIVX1 U2765 ( .A(n2586), .Z(n2587) );
  COND1XL U2766 ( .A(n2588), .B(n586), .C(n2587), .Z(N132) );
  COND1XL U2767 ( .A(n2501), .B(n588), .C(n440), .Z(N131) );
endmodule

