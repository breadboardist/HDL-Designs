
module sfilt ( clk, rst, pushin, cmd, q, h, pushout, z );
  input [1:0] cmd;
  input [31:0] q;
  input [31:0] h;
  output [31:0] z;
  input clk, rst, pushin;
  output pushout;
  wire   push_2, push0, push_1, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n562, n563,
         n564, n565, n566, n567, n568, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184;
  wire   [63:0] acc;
  wire   [1:0] cmd_2;
  wire   [6:0] h2;
  wire   [1:0] cmd0;
  wire   [6:0] h1;
  wire   [1:0] cmd_1;
  tri   clk;
  tri   [31:0] q0;
  tri   [31:0] h0;
  tri   [63:0] multout_1;
  tri   n3185;

  DW02_mult_3_stage pipe ( .p1(q0), .p2(h0), .p3(1'b1), .p4(clk), .p5(
        multout_1) );
  CFD2QXL \q0_reg[0]  ( .D(n64), .CP(clk), .CD(n3061), .Q(q0[0]) );
  CFD2QXL \h0_reg[31]  ( .D(n63), .CP(clk), .CD(n3061), .Q(h0[31]) );
  CFD2QXL \h0_reg[30]  ( .D(n62), .CP(clk), .CD(n3061), .Q(h0[30]) );
  CFD2QXL \h0_reg[29]  ( .D(n61), .CP(clk), .CD(n3061), .Q(h0[29]) );
  CFD2QXL \h0_reg[28]  ( .D(n60), .CP(clk), .CD(n3061), .Q(h0[28]) );
  CFD2QXL \h0_reg[27]  ( .D(n59), .CP(clk), .CD(n3061), .Q(h0[27]) );
  CFD2QXL \h0_reg[26]  ( .D(n58), .CP(clk), .CD(n3061), .Q(h0[26]) );
  CFD2QXL \h0_reg[25]  ( .D(n57), .CP(clk), .CD(n3061), .Q(h0[25]) );
  CFD2QXL \h0_reg[24]  ( .D(n56), .CP(clk), .CD(n3061), .Q(h0[24]) );
  CFD2QXL \h0_reg[23]  ( .D(n55), .CP(clk), .CD(n3061), .Q(h0[23]) );
  CFD2QXL \h0_reg[22]  ( .D(n54), .CP(clk), .CD(n3061), .Q(h0[22]) );
  CFD2QXL \h0_reg[21]  ( .D(n53), .CP(clk), .CD(n3061), .Q(h0[21]) );
  CFD2QXL \h0_reg[20]  ( .D(n52), .CP(clk), .CD(n3061), .Q(h0[20]) );
  CFD2QXL \h0_reg[19]  ( .D(n51), .CP(clk), .CD(n3061), .Q(h0[19]) );
  CFD2QXL \h0_reg[18]  ( .D(n50), .CP(clk), .CD(n3061), .Q(h0[18]) );
  CFD2QXL \h0_reg[17]  ( .D(n49), .CP(clk), .CD(n3061), .Q(h0[17]) );
  CFD2QXL \h0_reg[16]  ( .D(n48), .CP(clk), .CD(n3061), .Q(h0[16]) );
  CFD2QXL \h0_reg[15]  ( .D(n47), .CP(clk), .CD(n3061), .Q(h0[15]) );
  CFD2QXL \h0_reg[14]  ( .D(n46), .CP(clk), .CD(n3061), .Q(h0[14]) );
  CFD2QXL \h0_reg[13]  ( .D(n45), .CP(clk), .CD(n3061), .Q(h0[13]) );
  CFD2QXL \h0_reg[12]  ( .D(n44), .CP(clk), .CD(n3061), .Q(h0[12]) );
  CFD2QXL \h0_reg[11]  ( .D(n43), .CP(clk), .CD(n3061), .Q(h0[11]) );
  CFD2QXL \h0_reg[10]  ( .D(n42), .CP(clk), .CD(n3061), .Q(h0[10]) );
  CFD2QXL \h0_reg[9]  ( .D(n41), .CP(clk), .CD(n3061), .Q(h0[9]) );
  CFD2QXL \h0_reg[8]  ( .D(n40), .CP(clk), .CD(n3061), .Q(h0[8]) );
  CFD2QXL \h0_reg[7]  ( .D(n39), .CP(clk), .CD(n3061), .Q(h0[7]) );
  CFD2QXL \q0_reg[31]  ( .D(n31), .CP(clk), .CD(n3061), .Q(q0[31]) );
  CFD2QXL \q0_reg[30]  ( .D(n30), .CP(clk), .CD(n3061), .Q(q0[30]) );
  CFD2QXL \q0_reg[29]  ( .D(n29), .CP(clk), .CD(n3061), .Q(q0[29]) );
  CFD2QXL \q0_reg[28]  ( .D(n28), .CP(clk), .CD(n3061), .Q(q0[28]) );
  CFD2QXL \q0_reg[27]  ( .D(n27), .CP(clk), .CD(n3061), .Q(q0[27]) );
  CFD2QXL \q0_reg[26]  ( .D(n26), .CP(clk), .CD(n3061), .Q(q0[26]) );
  CFD2QXL \q0_reg[25]  ( .D(n25), .CP(clk), .CD(n3061), .Q(q0[25]) );
  CFD2QXL \q0_reg[24]  ( .D(n24), .CP(clk), .CD(n3061), .Q(q0[24]) );
  CFD2QXL \q0_reg[23]  ( .D(n23), .CP(clk), .CD(n3061), .Q(q0[23]) );
  CFD2QXL \q0_reg[22]  ( .D(n22), .CP(clk), .CD(n3061), .Q(q0[22]) );
  CFD2QXL \q0_reg[21]  ( .D(n21), .CP(clk), .CD(n3061), .Q(q0[21]) );
  CFD2QXL \q0_reg[20]  ( .D(n20), .CP(clk), .CD(n3061), .Q(q0[20]) );
  CFD2QXL \q0_reg[19]  ( .D(n19), .CP(clk), .CD(n3061), .Q(q0[19]) );
  CFD2QXL \q0_reg[18]  ( .D(n18), .CP(clk), .CD(n3061), .Q(q0[18]) );
  CFD2QXL \q0_reg[17]  ( .D(n17), .CP(clk), .CD(n3061), .Q(q0[17]) );
  CFD2QXL \q0_reg[16]  ( .D(n16), .CP(clk), .CD(n3061), .Q(q0[16]) );
  CFD2QXL \q0_reg[15]  ( .D(n15), .CP(clk), .CD(n3061), .Q(q0[15]) );
  CFD2QXL \q0_reg[14]  ( .D(n14), .CP(clk), .CD(n3061), .Q(q0[14]) );
  CFD2QXL \q0_reg[13]  ( .D(n13), .CP(clk), .CD(n3061), .Q(q0[13]) );
  CFD2QXL \q0_reg[12]  ( .D(n12), .CP(clk), .CD(n3061), .Q(q0[12]) );
  CFD2QXL \q0_reg[11]  ( .D(n11), .CP(clk), .CD(n3061), .Q(q0[11]) );
  CFD2QXL \q0_reg[10]  ( .D(n10), .CP(clk), .CD(n3061), .Q(q0[10]) );
  CFD2QXL \q0_reg[9]  ( .D(n9), .CP(clk), .CD(n3061), .Q(q0[9]) );
  CFD2QXL \q0_reg[8]  ( .D(n8), .CP(clk), .CD(n3061), .Q(q0[8]) );
  CFD2QXL \q0_reg[7]  ( .D(n7), .CP(clk), .CD(n3061), .Q(q0[7]) );
  CFD2QXL \q0_reg[6]  ( .D(n6), .CP(clk), .CD(n3061), .Q(q0[6]) );
  CFD2QXL \q0_reg[5]  ( .D(n5), .CP(clk), .CD(n3061), .Q(q0[5]) );
  CFD2QXL \q0_reg[4]  ( .D(n4), .CP(clk), .CD(n3061), .Q(q0[4]) );
  CFD2QXL \q0_reg[3]  ( .D(n3), .CP(clk), .CD(n3061), .Q(q0[3]) );
  CFD2QXL \q0_reg[2]  ( .D(n2), .CP(clk), .CD(n3061), .Q(q0[2]) );
  CFD2QXL \q0_reg[1]  ( .D(n1), .CP(clk), .CD(n3061), .Q(q0[1]) );
  CFD2QXL \h0_reg[6]  ( .D(n38), .CP(clk), .CD(n3061), .Q(h0[6]) );
  CFD2QXL \h0_reg[5]  ( .D(n37), .CP(clk), .CD(n3061), .Q(h0[5]) );
  CFD2QXL \h0_reg[4]  ( .D(n36), .CP(clk), .CD(n3061), .Q(h0[4]) );
  CFD2QXL \h0_reg[3]  ( .D(n35), .CP(clk), .CD(n3061), .Q(h0[3]) );
  CFD2QXL \h0_reg[2]  ( .D(n34), .CP(clk), .CD(n3061), .Q(h0[2]) );
  CFD2QXL \h0_reg[1]  ( .D(n33), .CP(clk), .CD(n3061), .Q(h0[1]) );
  CFD2QXL \h0_reg[0]  ( .D(n32), .CP(clk), .CD(n3061), .Q(h0[0]) );
  CFD2X1 \acc_reg[56]  ( .D(n577), .CP(clk), .CD(n3061), .Q(acc[56]), .QN(
        n3083) );
  CFD2X1 \acc_reg[50]  ( .D(n583), .CP(clk), .CD(n3061), .Q(acc[50]), .QN(
        n3081) );
  CFD2X1 \acc_reg[25]  ( .D(n608), .CP(clk), .CD(n3061), .Q(acc[25]), .QN(
        n3105) );
  CFD2X1 \acc_reg[24]  ( .D(n609), .CP(clk), .CD(n3061), .Q(acc[24]), .QN(
        n3099) );
  CFD2XL push_1_reg ( .D(n759), .CP(clk), .CD(n3061), .Q(push_1) );
  CFD2XL \cmd_2_reg[1]  ( .D(n761), .CP(clk), .CD(n3061), .Q(cmd_2[1]), .QN(
        n3091) );
  CFD2XL \cmd_2_reg[0]  ( .D(n757), .CP(clk), .CD(n3061), .Q(cmd_2[0]), .QN(
        n3092) );
  CFD2XL \cmd_1_reg[1]  ( .D(n755), .CP(clk), .CD(n3061), .Q(cmd_1[1]) );
  CFD2XL \cmd_1_reg[0]  ( .D(n753), .CP(clk), .CD(n3061), .Q(cmd_1[0]) );
  CFD2XL \cmd0_reg[1]  ( .D(cmd[1]), .CP(clk), .CD(n3061), .Q(cmd0[1]) );
  CFD2XL \cmd0_reg[0]  ( .D(cmd[0]), .CP(clk), .CD(n3061), .Q(cmd0[0]) );
  CFD2XL \h1_reg[6]  ( .D(n751), .CP(clk), .CD(n3061), .Q(h1[6]) );
  CFD2XL \h1_reg[5]  ( .D(n749), .CP(clk), .CD(n3061), .Q(h1[5]) );
  CFD2XL \h1_reg[4]  ( .D(n747), .CP(clk), .CD(n3061), .Q(h1[4]) );
  CFD2XL \h1_reg[3]  ( .D(n745), .CP(clk), .CD(n3061), .Q(h1[3]) );
  CFD2XL \h1_reg[2]  ( .D(n743), .CP(clk), .CD(n3061), .Q(h1[2]) );
  CFD2XL \h1_reg[1]  ( .D(n741), .CP(clk), .CD(n3061), .Q(h1[1]) );
  CFD2XL \h1_reg[0]  ( .D(n739), .CP(clk), .CD(n3061), .Q(h1[0]) );
  CFD2XL _pushout_reg ( .D(n3059), .CP(clk), .CD(n3061), .Q(pushout) );
  CFD2XL push0_reg ( .D(pushin), .CP(clk), .CD(n3061), .Q(push0) );
  CFD2XL \dout_reg[11]  ( .D(n654), .CP(clk), .CD(n3061), .Q(z[11]) );
  CFD2XL \dout_reg[9]  ( .D(n738), .CP(clk), .CD(n3061), .Q(z[9]) );
  CFD2XL \dout_reg[24]  ( .D(n641), .CP(clk), .CD(n3061), .Q(z[24]) );
  CFD2XL \dout_reg[31]  ( .D(n737), .CP(clk), .CD(n3061), .Q(z[31]) );
  CFD2XL \dout_reg[30]  ( .D(n736), .CP(clk), .CD(n3061), .Q(z[30]) );
  CFD2XL \dout_reg[29]  ( .D(n735), .CP(clk), .CD(n3061), .Q(z[29]) );
  CFD2XL \dout_reg[28]  ( .D(n734), .CP(clk), .CD(n3061), .Q(z[28]) );
  CFD2XL \dout_reg[27]  ( .D(n733), .CP(clk), .CD(n3061), .Q(z[27]) );
  CFD2XL \dout_reg[26]  ( .D(n732), .CP(clk), .CD(n3061), .Q(z[26]) );
  CFD2XL \dout_reg[25]  ( .D(n731), .CP(clk), .CD(n3061), .Q(z[25]) );
  CFD2XL \dout_reg[23]  ( .D(n730), .CP(clk), .CD(n3061), .Q(z[23]) );
  CFD2XL \dout_reg[22]  ( .D(n729), .CP(clk), .CD(n3061), .Q(z[22]) );
  CFD2XL \dout_reg[21]  ( .D(n727), .CP(clk), .CD(n3061), .Q(z[21]) );
  CFD2XL \dout_reg[20]  ( .D(n728), .CP(clk), .CD(n3061), .Q(z[20]) );
  CFD2XL \dout_reg[19]  ( .D(n726), .CP(clk), .CD(n3061), .Q(z[19]) );
  CFD2XL \dout_reg[18]  ( .D(n725), .CP(clk), .CD(n3061), .Q(z[18]) );
  CFD2XL \dout_reg[17]  ( .D(n724), .CP(clk), .CD(n3061), .Q(z[17]) );
  CFD2XL \dout_reg[16]  ( .D(n723), .CP(clk), .CD(n3061), .Q(z[16]) );
  CFD2XL \dout_reg[15]  ( .D(n721), .CP(clk), .CD(n3061), .Q(z[15]) );
  CFD2XL \dout_reg[14]  ( .D(n722), .CP(clk), .CD(n3061), .Q(z[14]) );
  CFD2XL \dout_reg[13]  ( .D(n720), .CP(clk), .CD(n3061), .Q(z[13]) );
  CFD2XL \dout_reg[12]  ( .D(n719), .CP(clk), .CD(n3061), .Q(z[12]) );
  CFD2XL \dout_reg[10]  ( .D(n718), .CP(clk), .CD(n3061), .Q(z[10]) );
  CFD2XL \dout_reg[8]  ( .D(n717), .CP(clk), .CD(n3061), .Q(z[8]) );
  CFD2XL \dout_reg[7]  ( .D(n706), .CP(clk), .CD(n3061), .Q(z[7]) );
  CFD2XL \dout_reg[6]  ( .D(n707), .CP(clk), .CD(n3061), .Q(z[6]) );
  CFD2XL \dout_reg[5]  ( .D(n715), .CP(clk), .CD(n3061), .Q(z[5]) );
  CFD2XL \dout_reg[4]  ( .D(n703), .CP(clk), .CD(n3061), .Q(z[4]) );
  CFD2XL \dout_reg[3]  ( .D(n711), .CP(clk), .CD(n3061), .Q(z[3]) );
  CFD2XL \dout_reg[2]  ( .D(n663), .CP(clk), .CD(n3061), .Q(z[2]) );
  CFD2XL \dout_reg[1]  ( .D(n710), .CP(clk), .CD(n3061), .Q(z[1]) );
  CFD2XL \dout_reg[0]  ( .D(n665), .CP(clk), .CD(n3061), .Q(z[0]) );
  CFD2X1 \acc_reg[0]  ( .D(n633), .CP(clk), .CD(n3061), .Q(acc[0]), .QN(n3071)
         );
  CFD2X1 \acc_reg[20]  ( .D(n613), .CP(clk), .CD(n3061), .Q(acc[20]), .QN(
        n3098) );
  CFD2X1 \acc_reg[1]  ( .D(n632), .CP(clk), .CD(n3061), .Q(acc[1]), .QN(n3067)
         );
  CFD2X1 \acc_reg[11]  ( .D(n622), .CP(clk), .CD(n3061), .Q(acc[11]), .QN(
        n3066) );
  CFD2X1 \acc_reg[26]  ( .D(n607), .CP(clk), .CD(n3061), .Q(acc[26]), .QN(
        n3076) );
  CFD2X1 \acc_reg[37]  ( .D(n596), .CP(clk), .CD(n3061), .Q(acc[37]), .QN(
        n3078) );
  CFD2X1 \acc_reg[33]  ( .D(n600), .CP(clk), .CD(n3061), .Q(acc[33]), .QN(
        n3077) );
  CFD1QX4 \h2_reg[5]  ( .D(n704), .CP(clk), .Q(h2[5]) );
  CFD2X2 \acc_reg[13]  ( .D(n620), .CP(clk), .CD(n3061), .Q(acc[13]) );
  CFD2X2 \acc_reg[47]  ( .D(n586), .CP(clk), .CD(n3061), .Q(acc[47]), .QN(
        n3074) );
  CFD2X2 \acc_reg[39]  ( .D(n594), .CP(clk), .CD(n3061), .Q(acc[39]), .QN(
        n3073) );
  CFD2X2 \acc_reg[5]  ( .D(n628), .CP(clk), .CD(n3061), .Q(acc[5]), .QN(n3068)
         );
  CFD2X2 \acc_reg[12]  ( .D(n621), .CP(clk), .CD(n3061), .Q(acc[12]), .QN(
        n3107) );
  CFD2X2 \acc_reg[14]  ( .D(n619), .CP(clk), .CD(n3061), .Q(acc[14]), .QN(n935) );
  CFD2X2 \acc_reg[42]  ( .D(n591), .CP(clk), .CD(n3061), .Q(acc[42]), .QN(
        n3089) );
  CFD2X2 \acc_reg[40]  ( .D(n593), .CP(clk), .CD(n3061), .Q(acc[40]), .QN(
        n3072) );
  CFD2X2 \acc_reg[54]  ( .D(n579), .CP(clk), .CD(n3061), .Q(acc[54]), .QN(
        n3111) );
  CFD2X2 \acc_reg[46]  ( .D(n587), .CP(clk), .CD(n3061), .Q(acc[46]), .QN(
        n3097) );
  CFD2X2 \acc_reg[7]  ( .D(n626), .CP(clk), .CD(n3061), .Q(acc[7]) );
  CFD2X2 \acc_reg[15]  ( .D(n618), .CP(clk), .CD(n3061), .Q(acc[15]), .QN(
        n2930) );
  CFD2X2 \acc_reg[10]  ( .D(n623), .CP(clk), .CD(n3061), .Q(acc[10]), .QN(
        n3063) );
  CFD2X2 \acc_reg[23]  ( .D(n610), .CP(clk), .CD(n3061), .Q(acc[23]), .QN(
        n3106) );
  CFD2X2 \acc_reg[19]  ( .D(n614), .CP(clk), .CD(n3061), .Q(acc[19]), .QN(
        n3102) );
  CFD2X2 \acc_reg[17]  ( .D(n616), .CP(clk), .CD(n3061), .Q(acc[17]), .QN(
        n3103) );
  CFD2X2 \acc_reg[28]  ( .D(n605), .CP(clk), .CD(n3061), .Q(acc[28]), .QN(
        n3090) );
  CFD2X2 \acc_reg[44]  ( .D(n589), .CP(clk), .CD(n3061), .Q(acc[44]), .QN(
        n3094) );
  CFD2X2 \acc_reg[36]  ( .D(n597), .CP(clk), .CD(n3061), .Q(acc[36]), .QN(
        n3096) );
  CFD2X2 \acc_reg[35]  ( .D(n598), .CP(clk), .CD(n3061), .Q(acc[35]), .QN(
        n3075) );
  CFD2X2 \acc_reg[31]  ( .D(n602), .CP(clk), .CD(n3061), .Q(acc[31]), .QN(
        n3062) );
  CFD2X2 \acc_reg[59]  ( .D(n574), .CP(clk), .CD(n3061), .Q(acc[59]), .QN(
        n3086) );
  CFD2X2 \acc_reg[3]  ( .D(n630), .CP(clk), .CD(n3061), .Q(acc[3]) );
  CFD2X2 \acc_reg[6]  ( .D(n627), .CP(clk), .CD(n3061), .Q(acc[6]), .QN(n3108)
         );
  CFD2X2 \acc_reg[34]  ( .D(n599), .CP(clk), .CD(n3061), .Q(acc[34]), .QN(
        n3118) );
  CFD2X2 \acc_reg[55]  ( .D(n578), .CP(clk), .CD(n3061), .Q(acc[55]), .QN(
        n2929) );
  CFD2X2 \acc_reg[49]  ( .D(n584), .CP(clk), .CD(n3061), .Q(acc[49]), .QN(
        n3085) );
  CFD2X2 \acc_reg[38]  ( .D(n595), .CP(clk), .CD(n3061), .Q(acc[38]), .QN(
        n3084) );
  CFD2X2 \acc_reg[2]  ( .D(n631), .CP(clk), .CD(n3061), .Q(acc[2]), .QN(n3070)
         );
  CFD2X2 \acc_reg[16]  ( .D(n617), .CP(clk), .CD(n3061), .Q(acc[16]), .QN(
        n3104) );
  CFD2X2 \acc_reg[60]  ( .D(n573), .CP(clk), .CD(n3061), .Q(acc[60]), .QN(
        n3113) );
  CFD2X2 \acc_reg[61]  ( .D(n572), .CP(clk), .CD(n3061), .Q(acc[61]), .QN(
        n3080) );
  CFD2X2 \acc_reg[43]  ( .D(n590), .CP(clk), .CD(n3061), .Q(acc[43]), .QN(
        n3087) );
  CFD2X2 \acc_reg[41]  ( .D(n592), .CP(clk), .CD(n3061), .Q(acc[41]), .QN(
        n3079) );
  CFD1QX4 \h2_reg[6]  ( .D(n712), .CP(clk), .Q(h2[6]) );
  CFD1QX4 \h2_reg[2]  ( .D(n716), .CP(clk), .Q(h2[2]) );
  CFD1QX4 \h2_reg[3]  ( .D(n714), .CP(clk), .Q(h2[3]) );
  CFD1QX4 \h2_reg[0]  ( .D(n705), .CP(clk), .Q(h2[0]) );
  CFD1QX4 \h2_reg[1]  ( .D(n567), .CP(clk), .Q(h2[1]) );
  CFD2X1 \acc_reg[9]  ( .D(n624), .CP(clk), .CD(n3061), .Q(acc[9]), .QN(n3064)
         );
  CFD1QX2 \h2_reg[4]  ( .D(n564), .CP(clk), .Q(h2[4]) );
  CFD2X1 push_2_reg ( .D(n708), .CP(clk), .CD(n3061), .Q(push_2), .QN(n3120)
         );
  CFD2X1 \acc_reg[45]  ( .D(n588), .CP(clk), .CD(n3061), .Q(acc[45]), .QN(
        n3117) );
  CFD2X1 \acc_reg[57]  ( .D(n576), .CP(clk), .CD(n3061), .Q(acc[57]), .QN(
        n3093) );
  CFD2X1 \acc_reg[8]  ( .D(n625), .CP(clk), .CD(n3061), .Q(acc[8]), .QN(n3069)
         );
  CFD2X1 \acc_reg[27]  ( .D(n606), .CP(clk), .CD(n3061), .Q(acc[27]), .QN(
        n3110) );
  CFD2X1 \acc_reg[63]  ( .D(n570), .CP(clk), .CD(n3061), .Q(acc[63]), .QN(
        n3065) );
  CFD2X1 \acc_reg[58]  ( .D(n575), .CP(clk), .CD(n3061), .Q(acc[58]), .QN(
        n3112) );
  CFD2X1 \acc_reg[51]  ( .D(n582), .CP(clk), .CD(n3061), .Q(acc[51]), .QN(
        n3115) );
  CFD2X1 \acc_reg[30]  ( .D(n603), .CP(clk), .CD(n3061), .Q(acc[30]), .QN(n937) );
  CFD2X1 \acc_reg[18]  ( .D(n615), .CP(clk), .CD(n3061), .Q(acc[18]), .QN(
        n3088) );
  CFD2X1 \acc_reg[52]  ( .D(n581), .CP(clk), .CD(n3061), .Q(acc[52]), .QN(
        n3114) );
  CFD2XL \acc_reg[29]  ( .D(n604), .CP(clk), .CD(n3061), .Q(acc[29]), .QN(
        n3109) );
  CFD2XL \acc_reg[22]  ( .D(n611), .CP(clk), .CD(n3061), .Q(acc[22]), .QN(
        n3100) );
  CFD2X1 \acc_reg[62]  ( .D(n571), .CP(clk), .CD(n3061), .Q(acc[62]), .QN(
        n3119) );
  CFD2XL \acc_reg[32]  ( .D(n601), .CP(clk), .CD(n3061), .Q(acc[32]), .QN(
        n3095) );
  CFD2X2 \acc_reg[48]  ( .D(n585), .CP(clk), .CD(n3061), .Q(acc[48]), .QN(
        n3116) );
  CFD2XL \acc_reg[21]  ( .D(n612), .CP(clk), .CD(n3061), .Q(acc[21]), .QN(
        n3101) );
  CFD2X1 \acc_reg[4]  ( .D(n629), .CP(clk), .CD(n3061), .Q(acc[4]) );
  CFD2X1 \acc_reg[53]  ( .D(n580), .CP(clk), .CD(n3061), .Q(acc[53]), .QN(
        n3082) );
  CND2XL U736 ( .A(n669), .B(n668), .Z(n2133) );
  CIVXL U737 ( .A(n2317), .Z(n668) );
  CIVXL U738 ( .A(n2283), .Z(n669) );
  CND2IX2 U739 ( .B(n1585), .A(n1921), .Z(n2088) );
  CIVX2 U740 ( .A(n1237), .Z(n1247) );
  CND2IX1 U741 ( .B(n1237), .A(acc[10]), .Z(n1098) );
  CNR2IX2 U742 ( .B(n670), .A(n1151), .Z(n1210) );
  CND2X2 U743 ( .A(n2226), .B(n1820), .Z(n670) );
  CND2X2 U744 ( .A(n674), .B(n671), .Z(n1070) );
  CNR2X2 U745 ( .A(n1875), .B(n1511), .Z(n671) );
  CND2X2 U746 ( .A(n673), .B(n672), .Z(n1875) );
  CND2X2 U747 ( .A(n1736), .B(n1941), .Z(n672) );
  CND2X2 U748 ( .A(n1732), .B(n1824), .Z(n673) );
  CIVX2 U749 ( .A(n1876), .Z(n674) );
  CND2X2 U750 ( .A(n676), .B(n675), .Z(n1876) );
  CND2X1 U751 ( .A(n1731), .B(n1754), .Z(n675) );
  CND2IX1 U752 ( .B(n1054), .A(n1053), .Z(n676) );
  CND2X2 U753 ( .A(n677), .B(n1691), .Z(n1669) );
  CND2X2 U754 ( .A(n677), .B(n1824), .Z(n1888) );
  CIVX2 U755 ( .A(n1663), .Z(n677) );
  CAOR2XL U756 ( .A(n2187), .B(n2155), .C(n2017), .D(n861), .Z(n678) );
  COND1XL U757 ( .A(n2873), .B(n2706), .C(n2705), .Z(n571) );
  CND2X2 U758 ( .A(n2107), .B(n2106), .Z(n2645) );
  CNIVX1 U759 ( .A(n2588), .Z(n679) );
  CNR2XL U760 ( .A(n688), .B(n2512), .Z(n1557) );
  CND2X1 U761 ( .A(n1665), .B(n1752), .Z(n1164) );
  CND2X1 U762 ( .A(n1665), .B(n1691), .Z(n1435) );
  CIVXL U763 ( .A(n2775), .Z(n680) );
  CIVXL U764 ( .A(n680), .Z(n681) );
  CND3XL U765 ( .A(n2163), .B(n2162), .C(n934), .Z(n2164) );
  CND3X1 U766 ( .A(n1371), .B(n1370), .C(n1369), .Z(n682) );
  CND3XL U767 ( .A(n1371), .B(n1370), .C(n1369), .Z(n683) );
  CIVXL U768 ( .A(n678), .Z(n684) );
  CIVX2 U769 ( .A(n684), .Z(n685) );
  CIVX3 U770 ( .A(n1368), .Z(n1371) );
  CND2XL U771 ( .A(n2866), .B(n3152), .Z(n624) );
  COND4CXL U772 ( .A(n2917), .B(n2865), .C(n2864), .D(push_2), .Z(n2866) );
  CENXL U773 ( .A(n2862), .B(n930), .Z(n2865) );
  CNR2XL U774 ( .A(n1405), .B(n1404), .Z(n686) );
  CNR2XL U775 ( .A(n2528), .B(n1974), .Z(n2827) );
  CENX1 U776 ( .A(n2521), .B(n765), .Z(n2526) );
  CNR2X2 U777 ( .A(n2218), .B(n2227), .Z(n2756) );
  CND2X2 U778 ( .A(n2233), .B(n2658), .Z(n2218) );
  CIVXL U779 ( .A(n1352), .Z(n970) );
  CNR2X2 U780 ( .A(n1632), .B(n1631), .Z(n1646) );
  CNR2X2 U781 ( .A(n1644), .B(n1643), .Z(n1645) );
  CND2XL U782 ( .A(n1265), .B(n3118), .Z(n1267) );
  CNR2X1 U783 ( .A(n1526), .B(n1524), .Z(n1613) );
  CIVXL U784 ( .A(n1524), .Z(n1525) );
  CIVXL U785 ( .A(n2837), .Z(n2871) );
  CNIVXL U786 ( .A(n2305), .Z(n687) );
  CANR2X1 U787 ( .A(n2908), .B(n2917), .C(n2916), .D(n2907), .Z(n2909) );
  COND1X1 U788 ( .A(n3120), .B(n2909), .C(n3161), .Z(n630) );
  CND3X2 U789 ( .A(n2071), .B(n2070), .C(n2069), .Z(n2072) );
  COND1X1 U790 ( .A(n3120), .B(n2527), .C(n3158), .Z(n629) );
  CANR2X1 U791 ( .A(n2917), .B(n2526), .C(n2916), .D(n2525), .Z(n2527) );
  COND1X1 U792 ( .A(n2873), .B(n2814), .C(n2813), .Z(n588) );
  CENXL U793 ( .A(n2797), .B(n2796), .Z(n2814) );
  COND1X1 U794 ( .A(n2873), .B(n2773), .C(n2772), .Z(n582) );
  COND1X1 U795 ( .A(n2873), .B(n2790), .C(n2789), .Z(n575) );
  CND2X2 U796 ( .A(n2556), .B(n2141), .Z(n2632) );
  CND2X2 U797 ( .A(n2568), .B(n2616), .Z(n2791) );
  CNR2X1 U798 ( .A(n1243), .B(acc[44]), .Z(n1002) );
  CNR2X1 U799 ( .A(n1243), .B(acc[46]), .Z(n1168) );
  CNR2X1 U800 ( .A(n2160), .B(n2587), .Z(n776) );
  COND1XL U801 ( .A(n2873), .B(n895), .C(n896), .Z(n597) );
  CND2XL U802 ( .A(n2449), .B(n2450), .Z(n895) );
  COR2XL U803 ( .A(n1594), .B(n701), .Z(n688) );
  CIVXL U804 ( .A(n1724), .Z(n1096) );
  COND1X1 U805 ( .A(n3120), .B(n2919), .C(n3159), .Z(n631) );
  CND3XL U806 ( .A(n1973), .B(n1786), .C(n1972), .Z(n689) );
  CND3X1 U807 ( .A(n1973), .B(n1786), .C(n1972), .Z(n690) );
  CAN2X1 U808 ( .A(n692), .B(n691), .Z(n2302) );
  CIVX20 U809 ( .A(n2301), .Z(n691) );
  CENXL U810 ( .A(n2300), .B(n2299), .Z(n692) );
  COND1X1 U811 ( .A(n2873), .B(n2755), .C(n2754), .Z(n606) );
  CNIVXL U812 ( .A(n2870), .Z(n693) );
  CND3XL U813 ( .A(n1415), .B(n1414), .C(n1413), .Z(n694) );
  CND3X1 U814 ( .A(n1415), .B(n1414), .C(n1413), .Z(n695) );
  CND3X1 U815 ( .A(n1412), .B(n1411), .C(h2[3]), .Z(n1415) );
  CND2IX1 U816 ( .B(n2587), .A(n2588), .Z(n2646) );
  CND3XL U817 ( .A(n2837), .B(n2446), .C(n679), .Z(n2447) );
  CNR2X2 U818 ( .A(n2579), .B(n2158), .Z(n2588) );
  CND3X1 U819 ( .A(n2446), .B(n2466), .C(n2448), .Z(n2174) );
  CIVXL U820 ( .A(n2529), .Z(n696) );
  CIVX2 U821 ( .A(n696), .Z(n697) );
  COND1XL U822 ( .A(n2873), .B(n2395), .C(n2394), .Z(n611) );
  COND1XL U823 ( .A(n2873), .B(n2380), .C(n2379), .Z(n604) );
  CANR1X2 U824 ( .A(n2146), .B(n2145), .C(n2171), .Z(n2568) );
  CANR1X2 U825 ( .A(n933), .B(n1131), .C(h2[6]), .Z(n1137) );
  CND2X1 U826 ( .A(n1614), .B(n1824), .Z(n870) );
  CND2X1 U827 ( .A(n2032), .B(n2323), .Z(n2497) );
  CANR1XL U828 ( .A(n2030), .B(n2029), .C(n2028), .Z(n698) );
  CANR1XL U829 ( .A(n2030), .B(n2029), .C(n2028), .Z(n2210) );
  CND4X1 U830 ( .A(n2179), .B(n2178), .C(n2177), .D(n2176), .Z(n699) );
  CND4X1 U831 ( .A(n2179), .B(n2178), .C(n2177), .D(n2176), .Z(n700) );
  CND4X1 U832 ( .A(n2179), .B(n2178), .C(n2177), .D(n2176), .Z(n2868) );
  CND3X2 U833 ( .A(n1841), .B(n1840), .C(n1839), .Z(n1509) );
  CNR3XL U834 ( .A(n2868), .B(n2407), .C(n2597), .Z(n2408) );
  CENXL U835 ( .A(n2133), .B(n2132), .Z(n2138) );
  CND2IX1 U836 ( .B(n2003), .A(n698), .Z(n701) );
  CND2IX1 U837 ( .B(n2003), .A(n2210), .Z(n2298) );
  CND2XL U838 ( .A(n2795), .B(n2794), .Z(n2796) );
  CENXL U839 ( .A(n2692), .B(n702), .Z(n2706) );
  CIVX20 U840 ( .A(n2867), .Z(n702) );
  CND2X1 U841 ( .A(n1743), .B(n1941), .Z(n1802) );
  CND3X2 U842 ( .A(n1190), .B(n1189), .C(n1188), .Z(n1743) );
  CND2XL U843 ( .A(n2446), .B(n2448), .Z(n2587) );
  COND1X1 U844 ( .A(n3120), .B(n1567), .C(n3153), .Z(n625) );
  CNIVX1 U845 ( .A(n661), .Z(n703) );
  CNIVX1 U846 ( .A(n563), .Z(n704) );
  CNIVX1 U847 ( .A(n568), .Z(n705) );
  CNIVX1 U848 ( .A(n658), .Z(n706) );
  CNIVX1 U849 ( .A(n659), .Z(n707) );
  CNIVX1 U850 ( .A(n709), .Z(n708) );
  CNIVX1 U851 ( .A(push_1), .Z(n709) );
  CNIVX1 U852 ( .A(n664), .Z(n710) );
  CNIVX1 U853 ( .A(n662), .Z(n711) );
  CMX2X4 U854 ( .A0(acc[0]), .A1(z[0]), .S(n2014), .Z(n665) );
  CNIVX1 U855 ( .A(n562), .Z(n712) );
  CMX2X2 U856 ( .A0(n713), .A1(z[2]), .S(n2014), .Z(n663) );
  CNIVX1 U857 ( .A(acc[2]), .Z(n713) );
  CNIVX1 U858 ( .A(n565), .Z(n714) );
  CNIVX1 U859 ( .A(n660), .Z(n715) );
  CNIVX1 U860 ( .A(n566), .Z(n716) );
  CNIVX1 U861 ( .A(n657), .Z(n717) );
  CNIVX1 U862 ( .A(n655), .Z(n718) );
  CNIVX1 U863 ( .A(n653), .Z(n719) );
  CNIVX1 U864 ( .A(n652), .Z(n720) );
  CNIVX1 U865 ( .A(n650), .Z(n721) );
  CNIVX1 U866 ( .A(n651), .Z(n722) );
  CNIVX1 U867 ( .A(n649), .Z(n723) );
  CNIVX1 U868 ( .A(n648), .Z(n724) );
  CNIVX1 U869 ( .A(n647), .Z(n725) );
  CNIVX1 U870 ( .A(n646), .Z(n726) );
  CNIVX1 U871 ( .A(n644), .Z(n727) );
  CNIVX1 U872 ( .A(n645), .Z(n728) );
  CNIVX1 U873 ( .A(n643), .Z(n729) );
  CNIVX1 U874 ( .A(n642), .Z(n730) );
  CNIVX1 U875 ( .A(n640), .Z(n731) );
  CNIVX1 U876 ( .A(n639), .Z(n732) );
  CNIVX1 U877 ( .A(n638), .Z(n733) );
  CNIVX1 U878 ( .A(n637), .Z(n734) );
  CNIVX1 U879 ( .A(n636), .Z(n735) );
  CNIVX1 U880 ( .A(n635), .Z(n736) );
  CNIVX1 U881 ( .A(n634), .Z(n737) );
  CMX2X1 U882 ( .A0(acc[9]), .A1(z[9]), .S(n2014), .Z(n656) );
  CNIVX1 U883 ( .A(n656), .Z(n738) );
  CAN3XL U884 ( .A(cmd_2[1]), .B(cmd_2[0]), .C(push_2), .Z(n3059) );
  CNIVX1 U885 ( .A(n740), .Z(n739) );
  CNIVX1 U886 ( .A(n2928), .Z(n740) );
  CNIVX1 U887 ( .A(n742), .Z(n741) );
  CNIVX1 U888 ( .A(n2927), .Z(n742) );
  CNIVX1 U889 ( .A(n744), .Z(n743) );
  CNIVX1 U890 ( .A(n2926), .Z(n744) );
  CNIVX1 U891 ( .A(n746), .Z(n745) );
  CNIVX1 U892 ( .A(n2924), .Z(n746) );
  CNIVX1 U893 ( .A(n748), .Z(n747) );
  CNIVX1 U894 ( .A(n2925), .Z(n748) );
  CNIVX1 U895 ( .A(n750), .Z(n749) );
  CNIVX1 U896 ( .A(n2923), .Z(n750) );
  CNIVX1 U897 ( .A(n752), .Z(n751) );
  CNIVX1 U898 ( .A(n2922), .Z(n752) );
  CNIVX3 U899 ( .A(cmd0[0]), .Z(n754) );
  CNIVX1 U900 ( .A(n754), .Z(n753) );
  CNIVX3 U901 ( .A(cmd0[1]), .Z(n756) );
  CNIVX1 U902 ( .A(n756), .Z(n755) );
  CNIVX3 U903 ( .A(cmd_1[0]), .Z(n758) );
  CNIVX1 U904 ( .A(n758), .Z(n757) );
  CNIVX3 U905 ( .A(push0), .Z(n760) );
  CNIVX1 U906 ( .A(n760), .Z(n759) );
  CNIVX3 U907 ( .A(cmd_1[1]), .Z(n762) );
  CNIVX1 U908 ( .A(n762), .Z(n761) );
  CND2X2 U909 ( .A(n1432), .B(n1431), .Z(n1433) );
  CND2X2 U910 ( .A(n1753), .B(n1824), .Z(n1432) );
  CND2X2 U911 ( .A(n1755), .B(n1941), .Z(n1431) );
  CND2X1 U912 ( .A(n1307), .B(acc[28]), .Z(n1257) );
  CIVXL U913 ( .A(n1848), .Z(n1462) );
  CND2X1 U914 ( .A(n1848), .B(n1847), .Z(n1538) );
  CNR2XL U915 ( .A(n1272), .B(n3105), .Z(n1273) );
  CNR2XL U916 ( .A(n1385), .B(n3101), .Z(n1268) );
  CND2X2 U917 ( .A(n1846), .B(n2057), .Z(n1857) );
  CND2XL U918 ( .A(n1764), .B(n1941), .Z(n1674) );
  CND2X1 U919 ( .A(n1298), .B(acc[10]), .Z(n1114) );
  CAN2X1 U920 ( .A(n1265), .B(n3083), .Z(n1074) );
  CNR2X2 U921 ( .A(n2043), .B(n2042), .Z(n2071) );
  COND1X2 U922 ( .A(n1890), .B(n1889), .C(n1940), .Z(n1891) );
  CIVX4 U923 ( .A(n1132), .Z(n1275) );
  CNR2X1 U924 ( .A(n1275), .B(n3105), .Z(n822) );
  CNIVXL U925 ( .A(n2366), .Z(n763) );
  CND2X2 U926 ( .A(n2094), .B(n1825), .Z(n1379) );
  CND2X2 U927 ( .A(n1261), .B(n1260), .Z(n1523) );
  CND2X2 U928 ( .A(n1258), .B(n1257), .Z(n1522) );
  CNR2X1 U929 ( .A(n1363), .B(n1362), .Z(n764) );
  CNR2XL U930 ( .A(n1363), .B(n1362), .Z(n765) );
  CNR2X2 U931 ( .A(n1363), .B(n1362), .Z(n2520) );
  CND2X2 U932 ( .A(n1584), .B(n1941), .Z(n1589) );
  CND2X2 U933 ( .A(n1477), .B(n1682), .Z(n1487) );
  CND2XL U934 ( .A(n2756), .B(n2427), .Z(n2708) );
  CNIVXL U935 ( .A(n2334), .Z(n766) );
  CIVX2 U936 ( .A(n1344), .Z(n767) );
  CNIVX1 U937 ( .A(n1454), .Z(n768) );
  CIVX3 U938 ( .A(n1344), .Z(n1243) );
  CND3X1 U939 ( .A(n1147), .B(n1146), .C(n1145), .Z(n769) );
  CND2X2 U940 ( .A(n1315), .B(n2037), .Z(n1316) );
  CND2IXL U941 ( .B(h2[2]), .A(n1466), .Z(n1467) );
  CND2X2 U942 ( .A(n1846), .B(n1825), .Z(n1256) );
  CANR1X1 U943 ( .A(n2030), .B(n2029), .C(n2028), .Z(n770) );
  CNR2X1 U944 ( .A(n2317), .B(n2132), .Z(n2323) );
  COND1X1 U945 ( .A(n1683), .B(n1096), .C(n1095), .Z(n2021) );
  CND2XL U946 ( .A(n1611), .B(n1941), .Z(n1461) );
  CND3X1 U947 ( .A(n1138), .B(n1137), .C(n1136), .Z(n1151) );
  CNR2X1 U948 ( .A(n1271), .B(n1270), .Z(n1847) );
  COND2X1 U949 ( .A(acc[55]), .B(n1416), .C(n1244), .D(acc[58]), .Z(n1242) );
  COND2X1 U950 ( .A(n2596), .B(n1898), .C(n1903), .D(n1897), .Z(n2347) );
  COND1XL U951 ( .A(n3107), .B(n1272), .C(n1114), .Z(n1119) );
  CNR2IX1 U952 ( .B(n2035), .A(n2034), .Z(n2041) );
  CNR3X2 U953 ( .A(n1496), .B(n1013), .C(n1012), .Z(n1583) );
  CND2X1 U954 ( .A(n1724), .B(n1684), .Z(n1685) );
  CNR2X1 U955 ( .A(n1277), .B(n1276), .Z(n1278) );
  CNR2X1 U956 ( .A(n1274), .B(n1273), .Z(n1279) );
  COND1X1 U957 ( .A(n2021), .B(n2022), .C(n2037), .Z(n1112) );
  CND2XL U958 ( .A(n2105), .B(n1820), .Z(n1113) );
  COND1X1 U959 ( .A(n2022), .B(n2021), .C(n2037), .Z(n2024) );
  CND2X1 U960 ( .A(n1744), .B(n1752), .Z(n1745) );
  CND2IXL U961 ( .B(n1937), .A(n2018), .Z(n1911) );
  CND3X1 U962 ( .A(n1841), .B(n1840), .C(n1839), .Z(n2091) );
  CND2X1 U963 ( .A(n2048), .B(n2054), .Z(n2052) );
  CND2X1 U964 ( .A(n1446), .B(n1766), .Z(n2098) );
  CNIVX1 U965 ( .A(n2180), .Z(n2101) );
  COND1X1 U966 ( .A(n1847), .B(n1897), .C(n2054), .Z(n1850) );
  CNR2IX1 U967 ( .B(n2409), .A(n1848), .Z(n1849) );
  COND1XL U968 ( .A(n2127), .B(n2591), .C(n2126), .Z(n2471) );
  COND1XL U969 ( .A(n1980), .B(n2863), .C(n1979), .Z(n2318) );
  CND2X1 U970 ( .A(n2166), .B(n2057), .Z(n1892) );
  COND1XL U971 ( .A(n1964), .B(n2337), .C(n1963), .Z(n2458) );
  CND2XL U972 ( .A(n2225), .B(n2017), .Z(n2727) );
  CND2X1 U973 ( .A(n2917), .B(push_2), .Z(n2873) );
  CNIVX1 U974 ( .A(pushin), .Z(n2921) );
  CNIVX2 U975 ( .A(pushin), .Z(n2920) );
  COND1XL U976 ( .A(n2873), .B(n2293), .C(n2292), .Z(n612) );
  COND1XL U977 ( .A(n2873), .B(n2744), .C(n2743), .Z(n576) );
  CNR2X1 U978 ( .A(n1386), .B(acc[36]), .Z(n771) );
  CNR2XL U979 ( .A(acc[37]), .B(n1418), .Z(n772) );
  CNR2X1 U980 ( .A(n771), .B(n772), .Z(n1520) );
  CMXI2XL U981 ( .A0(acc[62]), .A1(acc[63]), .S(h2[0]), .Z(n773) );
  CNR2IX1 U982 ( .B(n1139), .A(n773), .Z(n1765) );
  CIVX2 U983 ( .A(n2151), .Z(n774) );
  COND1X1 U984 ( .A(n2147), .B(n774), .C(n2816), .Z(n2035) );
  CND3XL U985 ( .A(n2038), .B(n2037), .C(n2036), .Z(n775) );
  CND2IX1 U986 ( .B(n2064), .A(n775), .Z(n2317) );
  CND2X1 U987 ( .A(n776), .B(n2588), .Z(n2793) );
  CIVXL U988 ( .A(n2054), .Z(n777) );
  COAN1X2 U989 ( .A(n1910), .B(n777), .C(n1911), .Z(n2454) );
  CNR2IX1 U990 ( .B(n3039), .A(n3038), .Z(n778) );
  COND1XL U991 ( .A(n2863), .B(n3040), .C(n3037), .Z(n779) );
  COND1XL U992 ( .A(n778), .B(n779), .C(n2916), .Z(n780) );
  CANR1XL U993 ( .A(n778), .B(n779), .C(n780), .Z(n2864) );
  CNR2IXL U994 ( .B(n2344), .A(n2345), .Z(n2405) );
  CND2X1 U995 ( .A(n2328), .B(n2853), .Z(n781) );
  CND2X1 U996 ( .A(n781), .B(n3021), .Z(n782) );
  CND2IXL U997 ( .B(n3022), .A(n3023), .Z(n783) );
  CENX1 U998 ( .A(n782), .B(n783), .Z(n2330) );
  CND2X1 U999 ( .A(n2713), .B(n2431), .Z(n784) );
  CNR2X1 U1000 ( .A(n784), .B(n2877), .Z(n785) );
  CND2X1 U1001 ( .A(n2715), .B(n2431), .Z(n786) );
  COND3X1 U1002 ( .A(n2887), .B(n784), .C(n2949), .D(n786), .Z(n787) );
  CANR1X1 U1003 ( .A(n2890), .B(n785), .C(n787), .Z(n788) );
  CNR2IX1 U1004 ( .B(n2951), .A(n2950), .Z(n789) );
  CENXL U1005 ( .A(n788), .B(n789), .Z(n2433) );
  CND2XL U1006 ( .A(acc[2]), .B(n1469), .Z(n790) );
  CND3XL U1007 ( .A(n790), .B(n1470), .C(n1471), .Z(n791) );
  CNR2XL U1008 ( .A(n1472), .B(n1898), .Z(n792) );
  CANR3XL U1009 ( .A(n1921), .B(n791), .C(n792), .D(n1814), .Z(n1473) );
  CND3XL U1010 ( .A(n2151), .B(n1944), .C(n1624), .Z(n793) );
  CND3XL U1011 ( .A(n2344), .B(n1768), .C(n1628), .Z(n794) );
  CND3X2 U1012 ( .A(n1629), .B(n793), .C(n794), .Z(n2818) );
  COND1XL U1013 ( .A(n1903), .B(n1904), .C(n1902), .Z(n795) );
  CND2XL U1014 ( .A(n2054), .B(n1896), .Z(n796) );
  COND1X1 U1015 ( .A(n1905), .B(n796), .C(n795), .Z(n1906) );
  CND3XL U1016 ( .A(n2775), .B(n2774), .C(n2406), .Z(n797) );
  CNR2XL U1017 ( .A(n797), .B(n2668), .Z(n2349) );
  CND2IXL U1018 ( .B(n2447), .A(n2448), .Z(n2449) );
  CIVX1 U1019 ( .A(n2863), .Z(n798) );
  CANR1XL U1020 ( .A(n2820), .B(n798), .C(n2821), .Z(n799) );
  CND2XL U1021 ( .A(n3033), .B(n2822), .Z(n800) );
  COND1XL U1022 ( .A(n799), .B(n800), .C(n2916), .Z(n801) );
  CANR1XL U1023 ( .A(n799), .B(n800), .C(n801), .Z(n2402) );
  CND2X1 U1024 ( .A(n2749), .B(n2751), .Z(n802) );
  CND2X1 U1025 ( .A(n2750), .B(n2751), .Z(n803) );
  COND3X1 U1026 ( .A(n2850), .B(n802), .C(n3001), .D(n803), .Z(n804) );
  CNR2X1 U1027 ( .A(n802), .B(n2843), .Z(n805) );
  CANR1XL U1028 ( .A(n2853), .B(n805), .C(n804), .Z(n806) );
  CNR2IXL U1029 ( .B(n3003), .A(n3002), .Z(n807) );
  CENX1 U1030 ( .A(n806), .B(n807), .Z(n2753) );
  CANR1XL U1031 ( .A(n2470), .B(n2890), .C(n2471), .Z(n808) );
  CNR2IX1 U1032 ( .B(n2973), .A(n2976), .Z(n809) );
  CENX1 U1033 ( .A(n808), .B(n809), .Z(n2129) );
  CND2XL U1034 ( .A(n1942), .B(n1752), .Z(n810) );
  COND1XL U1035 ( .A(n1551), .B(n1919), .C(n810), .Z(n2075) );
  CND2IXL U1036 ( .B(n2448), .A(n2447), .Z(n2450) );
  CND2IXL U1037 ( .B(n2180), .A(n2017), .Z(n2758) );
  CND3XL U1038 ( .A(n2035), .B(n2066), .C(n1940), .Z(n2748) );
  CND2X1 U1039 ( .A(n2319), .B(n2318), .Z(n811) );
  CND2X1 U1040 ( .A(n811), .B(n3025), .Z(n812) );
  CND2IXL U1041 ( .B(n3026), .A(n3027), .Z(n813) );
  CENX1 U1042 ( .A(n812), .B(n813), .Z(n2320) );
  CND2XL U1043 ( .A(n2890), .B(n2618), .Z(n814) );
  CIVX1 U1044 ( .A(n2805), .Z(n815) );
  CANR1XL U1045 ( .A(n2618), .B(n815), .C(n2620), .Z(n816) );
  COND1XL U1046 ( .A(n2800), .B(n814), .C(n816), .Z(n817) );
  CND2X1 U1047 ( .A(n2621), .B(n2969), .Z(n818) );
  CENX1 U1048 ( .A(n817), .B(n818), .Z(n2544) );
  CIVX1 U1049 ( .A(n2749), .Z(n819) );
  CNR2X1 U1050 ( .A(n2843), .B(n819), .Z(n820) );
  CNR2X1 U1051 ( .A(n2850), .B(n819), .Z(n821) );
  CANR3X1 U1052 ( .A(n2853), .B(n820), .C(n2750), .D(n821), .Z(n2247) );
  CANR1XL U1053 ( .A(acc[22]), .B(n1344), .C(n822), .Z(n1196) );
  CND2XL U1054 ( .A(n1623), .B(n1941), .Z(n823) );
  COND1XL U1055 ( .A(n1819), .B(n1613), .C(n823), .Z(n1810) );
  CNR2XL U1056 ( .A(n1817), .B(n1816), .Z(n824) );
  CND2X1 U1057 ( .A(n2057), .B(n824), .Z(n1476) );
  COND1XL U1058 ( .A(n2954), .B(n2953), .C(n2955), .Z(n825) );
  CANR1XL U1059 ( .A(n2201), .B(n2762), .C(n825), .Z(n2430) );
  CANR2X1 U1060 ( .A(n1481), .B(n3080), .C(n3065), .D(n2815), .Z(n826) );
  CND2X2 U1061 ( .A(n1084), .B(n826), .Z(n2596) );
  CANR1XL U1062 ( .A(n2441), .B(n2890), .C(n2440), .Z(n827) );
  CNR2IX1 U1063 ( .B(n2985), .A(n2988), .Z(n828) );
  CENX1 U1064 ( .A(n827), .B(n828), .Z(n2443) );
  CANR1XL U1065 ( .A(n2557), .B(n2890), .C(n2559), .Z(n829) );
  CNR2IX1 U1066 ( .B(n2981), .A(n2984), .Z(n830) );
  CENX1 U1067 ( .A(n829), .B(n830), .Z(n2452) );
  CIVX1 U1068 ( .A(n3020), .Z(n831) );
  CIVXL U1069 ( .A(n2276), .Z(n832) );
  COND1XL U1070 ( .A(n3020), .B(n832), .C(n3017), .Z(n833) );
  CANR11X1 U1071 ( .A(n2853), .B(n2275), .C(n831), .D(n833), .Z(n834) );
  CNR2IXL U1072 ( .B(n3019), .A(n3018), .Z(n835) );
  CENX1 U1073 ( .A(n834), .B(n835), .Z(n2278) );
  CND2IX1 U1074 ( .B(n3040), .A(n3037), .Z(n836) );
  COND1XL U1075 ( .A(n2863), .B(n836), .C(n2916), .Z(n837) );
  CANR1XL U1076 ( .A(n2863), .B(n836), .C(n837), .Z(n1565) );
  CAOR2X1 U1077 ( .A(n2076), .B(n2017), .C(n2234), .D(n2155), .Z(n2556) );
  CNR2IX1 U1078 ( .B(n2549), .A(n2964), .Z(n838) );
  CND2X1 U1079 ( .A(n2799), .B(n838), .Z(n839) );
  CIVXL U1080 ( .A(n2550), .Z(n840) );
  COND1XL U1081 ( .A(n2964), .B(n840), .C(n2961), .Z(n841) );
  CANR1XL U1082 ( .A(n838), .B(n2802), .C(n841), .Z(n842) );
  COND1XL U1083 ( .A(n2805), .B(n839), .C(n842), .Z(n843) );
  CNR2X1 U1084 ( .A(n839), .B(n2800), .Z(n844) );
  CANR1XL U1085 ( .A(n2890), .B(n844), .C(n843), .Z(n845) );
  CNR2IXL U1086 ( .B(n2963), .A(n2962), .Z(n846) );
  CENX1 U1087 ( .A(n845), .B(n846), .Z(n2552) );
  COND1XL U1088 ( .A(n3001), .B(n3002), .C(n3003), .Z(n847) );
  CANR1X1 U1089 ( .A(n2750), .B(n1965), .C(n847), .Z(n2264) );
  CND3XL U1090 ( .A(n2013), .B(acc[14]), .C(n1139), .Z(n848) );
  CND2XL U1091 ( .A(n1132), .B(acc[17]), .Z(n849) );
  CND2X1 U1092 ( .A(n849), .B(n848), .Z(n1652) );
  CND2XL U1093 ( .A(h2[5]), .B(n1819), .Z(n850) );
  CND2X1 U1094 ( .A(n850), .B(n1940), .Z(n2056) );
  COND1XL U1095 ( .A(n2946), .B(n2945), .C(n2947), .Z(n851) );
  CANR1XL U1096 ( .A(n2238), .B(n2714), .C(n851), .Z(n852) );
  COND1XL U1097 ( .A(n2430), .B(n2239), .C(n852), .Z(n2884) );
  CNR2IXL U1098 ( .B(n3041), .A(n3044), .Z(n853) );
  CENX1 U1099 ( .A(n2513), .B(n853), .Z(n2303) );
  CNR2XL U1100 ( .A(n3012), .B(n2386), .Z(n854) );
  COND1XL U1101 ( .A(n3012), .B(n2387), .C(n3009), .Z(n855) );
  CANR1XL U1102 ( .A(n2853), .B(n854), .C(n855), .Z(n856) );
  CNR2IXL U1103 ( .B(n3011), .A(n3010), .Z(n857) );
  CENX1 U1104 ( .A(n856), .B(n857), .Z(n2341) );
  COND1XL U1105 ( .A(n2532), .B(n2863), .C(n2531), .Z(n858) );
  CND2X1 U1106 ( .A(n3029), .B(n2832), .Z(n859) );
  CENX1 U1107 ( .A(n858), .B(n859), .Z(n860) );
  CAN2X1 U1108 ( .A(n2916), .B(n860), .Z(n2533) );
  CIVXL U1109 ( .A(n2094), .Z(n861) );
  CAOR2X1 U1110 ( .A(n2187), .B(n2155), .C(n2017), .D(n861), .Z(n2581) );
  CNR2X1 U1111 ( .A(n2984), .B(n2590), .Z(n862) );
  COND1XL U1112 ( .A(n2984), .B(n2591), .C(n2981), .Z(n863) );
  CANR1XL U1113 ( .A(n2890), .B(n862), .C(n863), .Z(n864) );
  CNR2IXL U1114 ( .B(n2983), .A(n2982), .Z(n865) );
  CENX1 U1115 ( .A(n864), .B(n865), .Z(n2593) );
  CNR3XL U1116 ( .A(n2489), .B(n2244), .C(n2491), .Z(n866) );
  CND3XL U1117 ( .A(n2499), .B(n866), .C(n2273), .Z(n2246) );
  CIVXL U1118 ( .A(n2890), .Z(n867) );
  COND1XL U1119 ( .A(n2877), .B(n867), .C(n2887), .Z(n868) );
  CND2IX1 U1120 ( .B(n2960), .A(n2957), .Z(n869) );
  CENX1 U1121 ( .A(n868), .B(n869), .Z(n2486) );
  CANR2XL U1122 ( .A(n1344), .B(acc[8]), .C(n1132), .D(acc[11]), .Z(n1352) );
  CND2IX1 U1123 ( .B(n1744), .A(n1658), .Z(n1659) );
  COND1X1 U1124 ( .A(n1551), .B(n1616), .C(n870), .Z(n1809) );
  CNR2IX1 U1125 ( .B(n1549), .A(n1550), .Z(n1919) );
  CND2XL U1126 ( .A(n1712), .B(n1752), .Z(n871) );
  CAN2X1 U1127 ( .A(n1714), .B(n871), .Z(n1719) );
  CND3X1 U1128 ( .A(n2023), .B(n1112), .C(n1113), .Z(n2296) );
  CNR2IX1 U1129 ( .B(n3049), .A(n3052), .Z(n872) );
  CENX1 U1130 ( .A(n2914), .B(n872), .Z(n2915) );
  CIVXL U1131 ( .A(n2890), .Z(n873) );
  COND1XL U1132 ( .A(n2650), .B(n873), .C(n2651), .Z(n874) );
  CND2IXL U1133 ( .B(n2980), .A(n2977), .Z(n875) );
  CENX1 U1134 ( .A(n874), .B(n875), .Z(n2653) );
  CIVX1 U1135 ( .A(n2988), .Z(n876) );
  CIVX1 U1136 ( .A(n2440), .Z(n877) );
  COND1XL U1137 ( .A(n2988), .B(n877), .C(n2985), .Z(n878) );
  CANR11XL U1138 ( .A(n2890), .B(n2441), .C(n876), .D(n878), .Z(n879) );
  CNR2IXL U1139 ( .B(n2987), .A(n2986), .Z(n880) );
  CENX1 U1140 ( .A(n879), .B(n880), .Z(n2314) );
  COND1XL U1141 ( .A(n3044), .B(n2513), .C(n3041), .Z(n881) );
  CND2IXL U1142 ( .B(n3042), .A(n3043), .Z(n882) );
  CENX1 U1143 ( .A(n881), .B(n882), .Z(n2514) );
  CND2X1 U1144 ( .A(n2830), .B(n2832), .Z(n883) );
  CND2X1 U1145 ( .A(n2831), .B(n2832), .Z(n884) );
  COND3X1 U1146 ( .A(n2863), .B(n883), .C(n3029), .D(n884), .Z(n885) );
  CND2IXL U1147 ( .B(n3030), .A(n3031), .Z(n886) );
  CENX1 U1148 ( .A(n885), .B(n886), .Z(n2833) );
  CANR1XL U1149 ( .A(n2459), .B(n2853), .C(n2458), .Z(n887) );
  CNR2IX1 U1150 ( .B(n3005), .A(n3008), .Z(n888) );
  CENX1 U1151 ( .A(n887), .B(n888), .Z(n2461) );
  CIVXL U1152 ( .A(n2489), .Z(n889) );
  CND3XL U1153 ( .A(n2746), .B(n2333), .C(n889), .Z(n2490) );
  CND2XL U1154 ( .A(n2890), .B(n2760), .Z(n890) );
  CIVXL U1155 ( .A(n2887), .Z(n891) );
  CANR1XL U1156 ( .A(n2760), .B(n891), .C(n2762), .Z(n892) );
  COND1XL U1157 ( .A(n2877), .B(n890), .C(n892), .Z(n893) );
  CND2X1 U1158 ( .A(n2763), .B(n2953), .Z(n894) );
  CENX1 U1159 ( .A(n893), .B(n894), .Z(n2222) );
  CANR1XL U1160 ( .A(n1949), .B(n2452), .C(n2451), .Z(n896) );
  CENXL U1161 ( .A(n2261), .B(n2260), .Z(n897) );
  CND2XL U1162 ( .A(n897), .B(n2436), .Z(n898) );
  CANR1XL U1163 ( .A(n1949), .B(n2272), .C(n2271), .Z(n899) );
  CND2XL U1164 ( .A(n898), .B(n899), .Z(n603) );
  CND2IX1 U1165 ( .B(n1386), .A(acc[6]), .Z(n1108) );
  CNR2XL U1166 ( .A(n1683), .B(n1652), .Z(n900) );
  CND3XL U1167 ( .A(n1422), .B(n1423), .C(n900), .Z(n1424) );
  CIVXL U1168 ( .A(n1453), .Z(n901) );
  CAOR1X1 U1169 ( .A(n1455), .B(n901), .C(n1192), .Z(n1218) );
  CND2IXL U1170 ( .B(n2501), .A(n2067), .Z(n2282) );
  CND2IX1 U1171 ( .B(n2512), .A(n2396), .Z(n2860) );
  CAN4X1 U1172 ( .A(n2079), .B(n2078), .C(n2080), .D(n1452), .Z(n902) );
  CANR2X1 U1173 ( .A(n2081), .B(n902), .C(n2077), .D(n2083), .Z(n2030) );
  COND1XL U1174 ( .A(n3052), .B(n2914), .C(n3049), .Z(n903) );
  CND2IXL U1175 ( .B(n3050), .A(n3051), .Z(n904) );
  CENX1 U1176 ( .A(n903), .B(n904), .Z(n2907) );
  CNR3XL U1177 ( .A(n2791), .B(n2792), .C(n2797), .Z(n905) );
  CND3XL U1178 ( .A(n2795), .B(n905), .C(n2465), .Z(n2468) );
  CND2IXL U1179 ( .B(n2226), .A(n2017), .Z(n2710) );
  CIVX1 U1180 ( .A(n3045), .Z(n906) );
  CANR1XL U1181 ( .A(n2524), .B(n2522), .C(n906), .Z(n2008) );
  COND1XL U1182 ( .A(n2980), .B(n2651), .C(n2977), .Z(n907) );
  CNR2XL U1183 ( .A(n2980), .B(n2650), .Z(n908) );
  CANR1XL U1184 ( .A(n2890), .B(n908), .C(n907), .Z(n909) );
  CNR2IXL U1185 ( .B(n2979), .A(n2978), .Z(n910) );
  CENX1 U1186 ( .A(n909), .B(n910), .Z(n2562) );
  CND2XL U1187 ( .A(n2582), .B(n2890), .Z(n911) );
  CND2X1 U1188 ( .A(n911), .B(n2989), .Z(n912) );
  CND2IX1 U1189 ( .B(n2990), .A(n2991), .Z(n913) );
  CENX1 U1190 ( .A(n912), .B(n913), .Z(n2584) );
  CIVX1 U1191 ( .A(n2863), .Z(n914) );
  COND4CXL U1192 ( .A(n2820), .B(n914), .C(n2821), .D(n2822), .Z(n915) );
  CND2XL U1193 ( .A(n915), .B(n3033), .Z(n916) );
  CND2IXL U1194 ( .B(n3034), .A(n3035), .Z(n917) );
  CENX1 U1195 ( .A(n916), .B(n917), .Z(n2823) );
  COND1XL U1196 ( .A(n3008), .B(n2850), .C(n3005), .Z(n918) );
  CNR2X1 U1197 ( .A(n3008), .B(n2843), .Z(n919) );
  CANR1XL U1198 ( .A(n2853), .B(n919), .C(n918), .Z(n920) );
  CNR2IXL U1199 ( .B(n3007), .A(n3006), .Z(n921) );
  CENX1 U1200 ( .A(n920), .B(n921), .Z(n2493) );
  CIVXL U1201 ( .A(n2887), .Z(n922) );
  CANR1XL U1202 ( .A(n2876), .B(n922), .C(n2884), .Z(n923) );
  CND2XL U1203 ( .A(n2890), .B(n2876), .Z(n924) );
  COND1XL U1204 ( .A(n2877), .B(n924), .C(n923), .Z(n925) );
  CND2X1 U1205 ( .A(n2734), .B(n2941), .Z(n926) );
  CENX1 U1206 ( .A(n925), .B(n926), .Z(n2241) );
  CANR1XL U1207 ( .A(n1949), .B(n1971), .C(n1970), .Z(n927) );
  CENXL U1208 ( .A(n1946), .B(n1947), .Z(n928) );
  CND2X1 U1209 ( .A(n928), .B(n2436), .Z(n929) );
  CND2X1 U1210 ( .A(n929), .B(n927), .Z(n605) );
  CND2IX1 U1211 ( .B(n1712), .A(n1941), .Z(n2046) );
  CND2IX1 U1212 ( .B(n1448), .A(n1450), .Z(n1236) );
  CND2IX1 U1213 ( .B(n1897), .A(n1940), .Z(n1904) );
  CND2IX1 U1214 ( .B(n2282), .A(n2031), .Z(n2244) );
  CNR2IX1 U1215 ( .B(n2861), .A(n2860), .Z(n930) );
  CND2IX1 U1216 ( .B(n3046), .A(n3047), .Z(n2009) );
  CND2IX1 U1217 ( .B(n3054), .A(n3055), .Z(n2900) );
  CND2IX1 U1218 ( .B(n3016), .A(n3013), .Z(n2505) );
  CND2IX1 U1219 ( .B(n695), .A(n2017), .Z(n2227) );
  CIVX1 U1220 ( .A(rst), .Z(n931) );
  CND2X1 U1221 ( .A(n931), .B(h1[0]), .Z(n932) );
  COND1XL U1222 ( .A(n2013), .B(n931), .C(n932), .Z(n568) );
  CAN2X1 U1223 ( .A(n1721), .B(n2037), .Z(n933) );
  CIVX4 U1224 ( .A(h2[2]), .Z(n1917) );
  CIVX8 U1225 ( .A(h2[6]), .Z(n2016) );
  CIVX3 U1226 ( .A(n1929), .Z(n1940) );
  CNR2IX4 U1227 ( .B(n2016), .A(n2015), .Z(n2017) );
  CIVX4 U1228 ( .A(n2148), .Z(n2057) );
  CIVX4 U1229 ( .A(n1537), .Z(n1682) );
  CIVX8 U1230 ( .A(n1192), .Z(n1941) );
  COR2X1 U1231 ( .A(n1480), .B(acc[61]), .Z(n936) );
  CAN2XL U1232 ( .A(n1525), .B(n1824), .Z(n938) );
  CIVX3 U1233 ( .A(h2[3]), .Z(n963) );
  CAN2XL U1234 ( .A(n2437), .B(n678), .Z(n939) );
  COND1X1 U1235 ( .A(n1638), .B(n1769), .C(n1124), .Z(n1125) );
  CND2X1 U1236 ( .A(n1472), .B(n1721), .Z(n1312) );
  CND2IX1 U1237 ( .B(n1385), .A(acc[35]), .Z(n1064) );
  CNR2X1 U1238 ( .A(n3091), .B(cmd_2[0]), .Z(n2917) );
  CNR2X4 U1239 ( .A(h2[0]), .B(h2[1]), .Z(n1344) );
  CIVX3 U1240 ( .A(n1344), .Z(n1416) );
  CNR2X1 U1241 ( .A(n1243), .B(n3095), .Z(n941) );
  CND2X2 U1242 ( .A(h2[0]), .B(h2[1]), .Z(n1259) );
  CIVX2 U1243 ( .A(n1259), .Z(n1303) );
  CAN2XL U1244 ( .A(acc[35]), .B(n1303), .Z(n940) );
  CNR2X1 U1245 ( .A(n941), .B(n940), .Z(n944) );
  CIVX8 U1246 ( .A(h2[1]), .Z(n1083) );
  CNR2X4 U1247 ( .A(n1083), .B(h2[0]), .Z(n1020) );
  CIVX3 U1248 ( .A(n1020), .Z(n1385) );
  CIVX4 U1249 ( .A(n1385), .Z(n1199) );
  CND2X1 U1250 ( .A(n1199), .B(acc[34]), .Z(n943) );
  CIVX4 U1251 ( .A(h2[0]), .Z(n948) );
  CNR2X4 U1252 ( .A(n948), .B(h2[1]), .Z(n1091) );
  CIVX2 U1253 ( .A(n1091), .Z(n1480) );
  CIVX4 U1254 ( .A(n1480), .Z(n1200) );
  CND2X1 U1255 ( .A(n1200), .B(acc[33]), .Z(n942) );
  CND3X2 U1256 ( .A(n944), .B(n943), .C(n942), .Z(n1585) );
  CND2X2 U1257 ( .A(n1917), .B(h2[3]), .Z(n1262) );
  CIVX4 U1258 ( .A(n1262), .Z(n1824) );
  CND2X1 U1259 ( .A(n1585), .B(n1824), .Z(n945) );
  CIVX2 U1260 ( .A(n945), .Z(n952) );
  CND2X2 U1261 ( .A(h2[2]), .B(h2[3]), .Z(n1192) );
  CND2X2 U1262 ( .A(n1199), .B(acc[38]), .Z(n947) );
  CND2X2 U1263 ( .A(n1200), .B(acc[37]), .Z(n946) );
  CND2X2 U1264 ( .A(n947), .B(n946), .Z(n1320) );
  CND2X2 U1265 ( .A(h2[0]), .B(h2[1]), .Z(n1166) );
  CIVX2 U1266 ( .A(n1166), .Z(n1297) );
  CND2X1 U1267 ( .A(n1297), .B(acc[39]), .Z(n950) );
  CAN2X2 U1268 ( .A(n948), .B(n1083), .Z(n1481) );
  CND2X1 U1269 ( .A(n1481), .B(acc[36]), .Z(n949) );
  CND2X1 U1270 ( .A(n950), .B(n949), .Z(n1318) );
  CNR2X2 U1271 ( .A(n1320), .B(n1318), .Z(n1590) );
  CNR2IX2 U1272 ( .B(n1941), .A(n1590), .Z(n951) );
  CNR2X2 U1273 ( .A(n952), .B(n951), .Z(n966) );
  CIVX2 U1274 ( .A(n1385), .Z(n1349) );
  CND2X1 U1275 ( .A(n1349), .B(acc[30]), .Z(n957) );
  CNR2X1 U1276 ( .A(n1243), .B(n3090), .Z(n954) );
  CIVX4 U1277 ( .A(n1303), .Z(n1417) );
  CNR2X1 U1278 ( .A(n3062), .B(n1417), .Z(n953) );
  CNR2X1 U1279 ( .A(n954), .B(n953), .Z(n956) );
  CND2X1 U1280 ( .A(n1200), .B(acc[29]), .Z(n955) );
  CND3X2 U1281 ( .A(n957), .B(n956), .C(n955), .Z(n1586) );
  CNR2X2 U1282 ( .A(n1917), .B(h2[3]), .Z(n1022) );
  CIVX2 U1283 ( .A(n1551), .Z(n1754) );
  CND2XL U1284 ( .A(n1586), .B(n1754), .Z(n965) );
  CNR2XL U1285 ( .A(n1416), .B(n3099), .Z(n959) );
  CNR2X1 U1286 ( .A(n1417), .B(n3110), .Z(n958) );
  CNR2XL U1287 ( .A(n959), .B(n958), .Z(n962) );
  CND2X1 U1288 ( .A(n1199), .B(acc[26]), .Z(n961) );
  CND2X1 U1289 ( .A(n1200), .B(acc[25]), .Z(n960) );
  CND3X1 U1290 ( .A(n962), .B(n961), .C(n960), .Z(n1634) );
  CND2X4 U1291 ( .A(n963), .B(n1917), .Z(n1819) );
  CIVX3 U1292 ( .A(n1819), .Z(n1752) );
  CND2XL U1293 ( .A(n1634), .B(n1752), .Z(n964) );
  CND3X2 U1294 ( .A(n966), .B(n965), .C(n964), .Z(n1910) );
  CND2X4 U1295 ( .A(n2016), .B(h2[5]), .Z(n2037) );
  CNR2IX4 U1296 ( .B(n2037), .A(n934), .Z(n1741) );
  CIVX3 U1297 ( .A(n1741), .Z(n1511) );
  CNR2X2 U1298 ( .A(n1910), .B(n1511), .Z(n967) );
  CIVX2 U1299 ( .A(n967), .Z(n996) );
  CIVX2 U1300 ( .A(n1091), .Z(n1115) );
  CNR2X1 U1301 ( .A(n1115), .B(n3064), .Z(n969) );
  CIVX2 U1302 ( .A(n1020), .Z(n1418) );
  CNR2X1 U1303 ( .A(n1418), .B(n3063), .Z(n968) );
  CNR2X1 U1304 ( .A(n969), .B(n968), .Z(n1351) );
  CIVX2 U1305 ( .A(n1351), .Z(n971) );
  CIVX2 U1306 ( .A(n1259), .Z(n1132) );
  CNR2X2 U1307 ( .A(n971), .B(n970), .Z(n1477) );
  CNR2IX2 U1308 ( .B(n2148), .A(n1819), .Z(n1721) );
  CND2XL U1309 ( .A(n1477), .B(n1721), .Z(n972) );
  CIVX2 U1310 ( .A(n2037), .Z(n1768) );
  CANR1XL U1311 ( .A(n2016), .B(n972), .C(n1768), .Z(n994) );
  CNR2XL U1312 ( .A(n1115), .B(n3101), .Z(n974) );
  CNR2X1 U1313 ( .A(n3106), .B(n1275), .Z(n973) );
  CNR2XL U1314 ( .A(n974), .B(n973), .Z(n977) );
  CND2XL U1315 ( .A(n1481), .B(acc[20]), .Z(n976) );
  COR2X1 U1316 ( .A(n1418), .B(n3100), .Z(n975) );
  CND3X1 U1317 ( .A(n977), .B(n976), .C(n975), .Z(n1512) );
  CIVX2 U1318 ( .A(n1512), .Z(n1639) );
  CIVDX2 U1319 ( .A(n989), .Z0(n1628), .Z1(n934) );
  CNR2X2 U1320 ( .A(n1192), .B(n1628), .Z(n1658) );
  CNR2X1 U1321 ( .A(n1683), .B(n1768), .Z(n1775) );
  CND2X1 U1322 ( .A(n1639), .B(n1775), .Z(n992) );
  CIVXL U1323 ( .A(n1020), .Z(n1272) );
  CND2XL U1324 ( .A(n1481), .B(acc[12]), .Z(n978) );
  COND1X1 U1325 ( .A(n935), .B(n1272), .C(n978), .Z(n982) );
  CIVX2 U1326 ( .A(n1091), .Z(n1104) );
  CND2X2 U1327 ( .A(n1347), .B(acc[13]), .Z(n980) );
  CND2X1 U1328 ( .A(n1297), .B(acc[15]), .Z(n979) );
  CND2X2 U1329 ( .A(n980), .B(n979), .Z(n981) );
  CNR2X2 U1330 ( .A(n982), .B(n981), .Z(n1640) );
  CIVX2 U1331 ( .A(n1022), .Z(n1898) );
  CNR2X2 U1332 ( .A(n1898), .B(n1628), .Z(n1684) );
  CIVX2 U1333 ( .A(n1684), .Z(n1638) );
  CNR2X1 U1334 ( .A(n1638), .B(n1768), .Z(n1773) );
  CND2X1 U1335 ( .A(n1640), .B(n1773), .Z(n991) );
  CND2X2 U1336 ( .A(n1199), .B(acc[18]), .Z(n984) );
  CND2X2 U1337 ( .A(n1347), .B(acc[17]), .Z(n983) );
  CND2X2 U1338 ( .A(n984), .B(n983), .Z(n988) );
  CND2XL U1339 ( .A(n1297), .B(acc[19]), .Z(n986) );
  CNIVX2 U1340 ( .A(n1344), .Z(n1298) );
  CND2XL U1341 ( .A(n1298), .B(acc[16]), .Z(n985) );
  CND2X1 U1342 ( .A(n986), .B(n985), .Z(n987) );
  CNR2X2 U1343 ( .A(n988), .B(n987), .Z(n1633) );
  CND3X2 U1344 ( .A(n1917), .B(h2[3]), .C(n989), .Z(n1537) );
  CNR2X1 U1345 ( .A(n1537), .B(n1768), .Z(n1771) );
  CND2X1 U1346 ( .A(n1633), .B(n1771), .Z(n990) );
  CND3X2 U1347 ( .A(n992), .B(n991), .C(n990), .Z(n993) );
  CNR2X2 U1348 ( .A(n994), .B(n993), .Z(n995) );
  CND2X2 U1349 ( .A(n996), .B(n995), .Z(n1597) );
  CNR2X1 U1350 ( .A(n767), .B(acc[52]), .Z(n998) );
  CAN2X1 U1351 ( .A(n1303), .B(n2929), .Z(n997) );
  CNR2X2 U1352 ( .A(n998), .B(n997), .Z(n1001) );
  COR2XL U1353 ( .A(acc[54]), .B(n1418), .Z(n1000) );
  CND2X1 U1354 ( .A(n1347), .B(n3082), .Z(n999) );
  CND3X2 U1355 ( .A(n1001), .B(n1000), .C(n999), .Z(n1578) );
  CND2XL U1356 ( .A(n1578), .B(n1941), .Z(n1017) );
  CND2X2 U1357 ( .A(n1349), .B(n3097), .Z(n1500) );
  CND2X1 U1358 ( .A(n1200), .B(n3117), .Z(n1499) );
  CIVX2 U1359 ( .A(n1002), .Z(n1498) );
  CNIVX4 U1360 ( .A(n1166), .Z(n1224) );
  CNR2X2 U1361 ( .A(n1224), .B(acc[47]), .Z(n1003) );
  CIVX2 U1362 ( .A(n1003), .Z(n1497) );
  CND4XL U1363 ( .A(n1500), .B(n1499), .C(n1498), .D(n1497), .Z(n1004) );
  CND2XL U1364 ( .A(n1004), .B(n1754), .Z(n1016) );
  CNR2X1 U1365 ( .A(n1417), .B(acc[51]), .Z(n1006) );
  CNR2X1 U1366 ( .A(n1243), .B(acc[48]), .Z(n1005) );
  CNR2X2 U1367 ( .A(n1006), .B(n1005), .Z(n1009) );
  CIVX3 U1368 ( .A(n1385), .Z(n1478) );
  CND2X1 U1369 ( .A(n1478), .B(n3081), .Z(n1008) );
  CND2X1 U1370 ( .A(n1200), .B(n3085), .Z(n1007) );
  CND3X2 U1371 ( .A(n1009), .B(n1008), .C(n1007), .Z(n1577) );
  CND2X1 U1372 ( .A(n1577), .B(n1824), .Z(n1015) );
  CND2X1 U1373 ( .A(n1297), .B(acc[43]), .Z(n1011) );
  CND2XL U1374 ( .A(n1344), .B(acc[40]), .Z(n1010) );
  CND2X2 U1375 ( .A(n1011), .B(n1010), .Z(n1496) );
  CND2X2 U1376 ( .A(n1199), .B(acc[42]), .Z(n1321) );
  CIVX2 U1377 ( .A(n1321), .Z(n1013) );
  CND2X2 U1378 ( .A(n1200), .B(acc[41]), .Z(n1322) );
  CIVX2 U1379 ( .A(n1322), .Z(n1012) );
  CND2X1 U1380 ( .A(n1583), .B(n1752), .Z(n1014) );
  CND4X2 U1381 ( .A(n1017), .B(n1016), .C(n1015), .D(n1014), .Z(n2020) );
  CIVX3 U1382 ( .A(h2[5]), .Z(n1937) );
  CNR2X2 U1383 ( .A(n1937), .B(n1628), .Z(n1825) );
  CND2X1 U1384 ( .A(n2020), .B(n1825), .Z(n1027) );
  CNR2X1 U1385 ( .A(n1417), .B(acc[63]), .Z(n1019) );
  CNR2X1 U1386 ( .A(n1243), .B(acc[60]), .Z(n1018) );
  CNR2X2 U1387 ( .A(n1019), .B(n1018), .Z(n1337) );
  CIVX2 U1388 ( .A(n1020), .Z(n1238) );
  CNR2X1 U1389 ( .A(acc[62]), .B(n1238), .Z(n1021) );
  CND2IX2 U1390 ( .B(n1021), .A(n936), .Z(n1335) );
  CNR2IX2 U1391 ( .B(n1337), .A(n1335), .Z(n1647) );
  CIVDX2 U1392 ( .A(n1022), .Z0(n1551), .Z1(n1915) );
  CIVX2 U1393 ( .A(n1819), .Z(n1395) );
  CNR2IXL U1394 ( .B(n1344), .A(acc[56]), .Z(n1024) );
  CNR2X2 U1395 ( .A(n1224), .B(acc[59]), .Z(n1023) );
  CNR2X2 U1396 ( .A(n1024), .B(n1023), .Z(n1340) );
  CND2X1 U1397 ( .A(n1199), .B(n3112), .Z(n1339) );
  CND2X1 U1398 ( .A(n1347), .B(n3093), .Z(n1338) );
  CAN3X2 U1399 ( .A(n1340), .B(n1339), .C(n1338), .Z(n1025) );
  CANR2X2 U1400 ( .A(n1647), .B(n1915), .C(n2409), .D(n1025), .Z(n2018) );
  CND2X1 U1401 ( .A(h2[5]), .B(h2[4]), .Z(n1738) );
  CIVX2 U1402 ( .A(n1738), .Z(n1820) );
  CND2XL U1403 ( .A(n2018), .B(n1820), .Z(n1026) );
  CND2X1 U1404 ( .A(n1027), .B(n1026), .Z(n1598) );
  CNR2X1 U1405 ( .A(n1597), .B(n1598), .Z(n2396) );
  CIVX1 U1406 ( .A(n2396), .Z(n1558) );
  CNR2X1 U1407 ( .A(n1417), .B(acc[48]), .Z(n1029) );
  CNR2X1 U1408 ( .A(n1416), .B(acc[45]), .Z(n1028) );
  CNR2X2 U1409 ( .A(n1029), .B(n1028), .Z(n1032) );
  CIVX2 U1410 ( .A(n1091), .Z(n1237) );
  CIVX2 U1411 ( .A(n1237), .Z(n1228) );
  CND2X1 U1412 ( .A(n1228), .B(n3097), .Z(n1031) );
  CND2X1 U1413 ( .A(n1478), .B(n3074), .Z(n1030) );
  CND3X2 U1414 ( .A(n1032), .B(n1031), .C(n1030), .Z(n1713) );
  CND2XL U1415 ( .A(n1713), .B(n1824), .Z(n1039) );
  CNR2X1 U1416 ( .A(n1417), .B(acc[52]), .Z(n1034) );
  CNR2X1 U1417 ( .A(n767), .B(acc[49]), .Z(n1033) );
  CNR2X2 U1418 ( .A(n1034), .B(n1033), .Z(n1037) );
  CND2X1 U1419 ( .A(n1349), .B(n3115), .Z(n1036) );
  CND2X1 U1420 ( .A(n1347), .B(n3081), .Z(n1035) );
  CND3X2 U1421 ( .A(n1037), .B(n1036), .C(n1035), .Z(n1715) );
  CND2XL U1422 ( .A(n1715), .B(n1941), .Z(n1038) );
  CND2X1 U1423 ( .A(n1039), .B(n1038), .Z(n1879) );
  CND2X1 U1424 ( .A(acc[39]), .B(n1478), .Z(n1041) );
  CND2X1 U1425 ( .A(n1247), .B(acc[38]), .Z(n1040) );
  CND2X2 U1426 ( .A(n1041), .B(n1040), .Z(n1045) );
  CND2X1 U1427 ( .A(n1297), .B(acc[40]), .Z(n1043) );
  CND2X1 U1428 ( .A(n1481), .B(acc[37]), .Z(n1042) );
  CND2X1 U1429 ( .A(n1043), .B(n1042), .Z(n1044) );
  CNR2X2 U1430 ( .A(n1045), .B(n1044), .Z(n1693) );
  CIVX2 U1431 ( .A(n1819), .Z(n1921) );
  CND2X1 U1432 ( .A(n1693), .B(n1921), .Z(n1052) );
  CNR2IXL U1433 ( .B(n3087), .A(n1385), .Z(n1046) );
  CIVX1 U1434 ( .A(n1046), .Z(n1050) );
  COND2X2 U1435 ( .A(acc[41]), .B(n1416), .C(n1417), .D(acc[44]), .Z(n1047) );
  CIVX2 U1436 ( .A(n1047), .Z(n1049) );
  CND2X1 U1437 ( .A(n1347), .B(n3089), .Z(n1048) );
  CND3X2 U1438 ( .A(n1050), .B(n1049), .C(n1048), .Z(n1712) );
  CND2X1 U1439 ( .A(n1712), .B(n1754), .Z(n1051) );
  CND2X2 U1440 ( .A(n1052), .B(n1051), .Z(n1880) );
  COND1X2 U1441 ( .A(n1879), .B(n1880), .C(n1825), .Z(n1071) );
  CIVX2 U1442 ( .A(n1921), .Z(n1054) );
  COR2X1 U1443 ( .A(n3099), .B(n1275), .Z(n1398) );
  CND2IX1 U1444 ( .B(n1243), .A(acc[21]), .Z(n1397) );
  CND2X1 U1445 ( .A(n1478), .B(acc[23]), .Z(n1400) );
  CND2X1 U1446 ( .A(n1247), .B(acc[22]), .Z(n1399) );
  CND4X1 U1447 ( .A(n1398), .B(n1397), .C(n1400), .D(n1399), .Z(n1053) );
  CNR2XL U1448 ( .A(n1243), .B(n3105), .Z(n1056) );
  CNR2X1 U1449 ( .A(n3090), .B(n1275), .Z(n1055) );
  CNR2XL U1450 ( .A(n1056), .B(n1055), .Z(n1059) );
  CND2X1 U1451 ( .A(n1247), .B(acc[26]), .Z(n1058) );
  CND2X1 U1452 ( .A(n1199), .B(acc[27]), .Z(n1057) );
  CND3X1 U1453 ( .A(n1059), .B(n1058), .C(n1057), .Z(n1731) );
  CND2X1 U1454 ( .A(n1247), .B(acc[34]), .Z(n1063) );
  CND2X1 U1455 ( .A(n1297), .B(acc[36]), .Z(n1061) );
  CND2XL U1456 ( .A(n1344), .B(acc[33]), .Z(n1060) );
  CAN2X1 U1457 ( .A(n1061), .B(n1060), .Z(n1062) );
  CND3X2 U1458 ( .A(n1064), .B(n1063), .C(n1062), .Z(n1736) );
  CNR2XL U1459 ( .A(n1416), .B(n3109), .Z(n1066) );
  CNR2X1 U1460 ( .A(n3095), .B(n1275), .Z(n1065) );
  CNR2X1 U1461 ( .A(n1066), .B(n1065), .Z(n1069) );
  CND2X1 U1462 ( .A(n1478), .B(acc[31]), .Z(n1068) );
  CND2X1 U1463 ( .A(n1247), .B(acc[30]), .Z(n1067) );
  CND3X2 U1464 ( .A(n1069), .B(n1068), .C(n1067), .Z(n1732) );
  CND2X2 U1465 ( .A(n1071), .B(n1070), .Z(n1072) );
  CIVX2 U1466 ( .A(n1072), .Z(n2023) );
  CNR2X1 U1467 ( .A(n767), .B(acc[53]), .Z(n1073) );
  CNR2X2 U1468 ( .A(n1074), .B(n1073), .Z(n1701) );
  CND2X1 U1469 ( .A(n1349), .B(n2929), .Z(n1700) );
  CND2X1 U1470 ( .A(n1347), .B(n3111), .Z(n1699) );
  CND3X1 U1471 ( .A(n1701), .B(n1700), .C(n1699), .Z(n1716) );
  CND2X1 U1472 ( .A(n1716), .B(n1921), .Z(n1081) );
  CNR2X1 U1473 ( .A(n1243), .B(acc[57]), .Z(n1076) );
  CNR2X1 U1474 ( .A(n1417), .B(acc[60]), .Z(n1075) );
  CNR2X2 U1475 ( .A(n1076), .B(n1075), .Z(n1079) );
  CIVX2 U1476 ( .A(n1418), .Z(n1306) );
  CND2XL U1477 ( .A(n1306), .B(n3086), .Z(n1078) );
  CIVX2 U1478 ( .A(n1091), .Z(n1140) );
  CIVX4 U1479 ( .A(n1140), .Z(n1307) );
  CND2X1 U1480 ( .A(n1307), .B(n3112), .Z(n1077) );
  CND3X2 U1481 ( .A(n1079), .B(n1078), .C(n1077), .Z(n1903) );
  CND2X1 U1482 ( .A(n1903), .B(h2[2]), .Z(n1080) );
  CND2X1 U1483 ( .A(n1081), .B(n1080), .Z(n1883) );
  CIVX2 U1484 ( .A(n1883), .Z(n1086) );
  CIVXL U1485 ( .A(h2[0]), .Z(n2013) );
  CNR2XL U1486 ( .A(acc[62]), .B(n2013), .Z(n1082) );
  CNR2XL U1487 ( .A(n1303), .B(n1082), .Z(n1084) );
  CNIVX4 U1488 ( .A(n1083), .Z(n1139) );
  CIVX2 U1489 ( .A(n1139), .Z(n2815) );
  CIVX2 U1490 ( .A(n2596), .Z(n1900) );
  CANR1X1 U1491 ( .A(n1917), .B(n1900), .C(n963), .Z(n1884) );
  CIVX2 U1492 ( .A(n1884), .Z(n1085) );
  CND2X2 U1493 ( .A(n1086), .B(n1085), .Z(n2105) );
  CND2X1 U1494 ( .A(n1247), .B(acc[18]), .Z(n1791) );
  CIVX2 U1495 ( .A(n1791), .Z(n1090) );
  CND2X1 U1496 ( .A(n1297), .B(acc[20]), .Z(n1088) );
  CND2X1 U1497 ( .A(n1481), .B(acc[17]), .Z(n1087) );
  CND2X1 U1498 ( .A(n1088), .B(n1087), .Z(n1789) );
  CND2X2 U1499 ( .A(n1478), .B(acc[19]), .Z(n1790) );
  CIVX2 U1500 ( .A(n1790), .Z(n1089) );
  CNR3X2 U1501 ( .A(n1090), .B(n1789), .C(n1089), .Z(n1724) );
  CANR2XL U1502 ( .A(acc[14]), .B(n1091), .C(acc[13]), .D(n1344), .Z(n1092) );
  COND1X1 U1503 ( .A(n2930), .B(n1385), .C(n1092), .Z(n1094) );
  CIVXL U1504 ( .A(n1259), .Z(n1469) );
  CAN2XL U1505 ( .A(n1469), .B(acc[16]), .Z(n1093) );
  CNR2X1 U1506 ( .A(n1094), .B(n1093), .Z(n1725) );
  CND2X1 U1507 ( .A(n1725), .B(n1682), .Z(n1095) );
  CND2XL U1508 ( .A(n1297), .B(acc[12]), .Z(n1097) );
  CND2X2 U1509 ( .A(n1098), .B(n1097), .Z(n1101) );
  CND2XL U1510 ( .A(n1344), .B(acc[9]), .Z(n1099) );
  COND1X1 U1511 ( .A(n3066), .B(n1272), .C(n1099), .Z(n1100) );
  CNR2X2 U1512 ( .A(n1101), .B(n1100), .Z(n1722) );
  CND2X1 U1513 ( .A(n1722), .B(n1684), .Z(n1102) );
  CND2X1 U1514 ( .A(n1102), .B(n2016), .Z(n1103) );
  CIVX2 U1515 ( .A(n1103), .Z(n1111) );
  CIVDX2 U1516 ( .A(n1104), .Z0(n1347), .Z1(n1386) );
  COR2XL U1517 ( .A(n3068), .B(n1243), .Z(n1107) );
  COR2XL U1518 ( .A(n3069), .B(n1275), .Z(n1106) );
  CND2X1 U1519 ( .A(n1478), .B(acc[7]), .Z(n1105) );
  CND4X2 U1520 ( .A(n1108), .B(n1107), .C(n1106), .D(n1105), .Z(n1392) );
  CIVX2 U1521 ( .A(n1392), .Z(n1109) );
  CND2X2 U1522 ( .A(n1109), .B(n1721), .Z(n1110) );
  CND2X2 U1523 ( .A(n1111), .B(n1110), .Z(n2022) );
  CIVX4 U1524 ( .A(n1115), .Z(n1193) );
  CND2X1 U1525 ( .A(n1193), .B(acc[11]), .Z(n1117) );
  CND2X1 U1526 ( .A(n1297), .B(acc[13]), .Z(n1116) );
  CND2X1 U1527 ( .A(n1117), .B(n1116), .Z(n1118) );
  CNR2X1 U1528 ( .A(n1119), .B(n1118), .Z(n1426) );
  CIVX2 U1529 ( .A(n1426), .Z(n1769) );
  CNR2X1 U1530 ( .A(n1416), .B(n3088), .Z(n1121) );
  CNR2X1 U1531 ( .A(n1238), .B(n3098), .Z(n1120) );
  CNR2X1 U1532 ( .A(n1121), .B(n1120), .Z(n1438) );
  CNR2X1 U1533 ( .A(n1140), .B(n3102), .Z(n1123) );
  CAN2XL U1534 ( .A(acc[21]), .B(n1132), .Z(n1122) );
  CNR2X1 U1535 ( .A(n1123), .B(n1122), .Z(n1437) );
  CND3XL U1536 ( .A(n1438), .B(n1437), .C(n1658), .Z(n1124) );
  CND2IX1 U1537 ( .B(n1768), .A(n1125), .Z(n1138) );
  CNR2XL U1538 ( .A(n1416), .B(n3108), .Z(n1127) );
  CNR2X1 U1539 ( .A(n3064), .B(n1275), .Z(n1126) );
  CNR2XL U1540 ( .A(n1127), .B(n1126), .Z(n1130) );
  CIVX2 U1541 ( .A(n1238), .Z(n1227) );
  CND2X1 U1542 ( .A(n1227), .B(acc[8]), .Z(n1129) );
  CND2XL U1543 ( .A(n1193), .B(acc[7]), .Z(n1128) );
  CND3X1 U1544 ( .A(n1130), .B(n1129), .C(n1128), .Z(n1428) );
  CIVX2 U1545 ( .A(n1428), .Z(n1131) );
  CIVXL U1546 ( .A(n1652), .Z(n1133) );
  CAN2X1 U1547 ( .A(n1682), .B(n1133), .Z(n1135) );
  CND2X1 U1548 ( .A(n1193), .B(acc[15]), .Z(n1422) );
  CIVX2 U1549 ( .A(n1238), .Z(n1248) );
  CND2X1 U1550 ( .A(n1248), .B(acc[16]), .Z(n1423) );
  CND2X1 U1551 ( .A(n1422), .B(n1423), .Z(n1653) );
  CIVX2 U1552 ( .A(n1653), .Z(n1134) );
  CND3X2 U1553 ( .A(n1135), .B(n2037), .C(n1134), .Z(n1136) );
  CIVX2 U1554 ( .A(n1765), .Z(n2691) );
  COND1X1 U1555 ( .A(h2[2]), .B(n2691), .C(h2[3]), .Z(n1150) );
  CNR2X1 U1556 ( .A(n1237), .B(acc[59]), .Z(n1406) );
  CIVXL U1557 ( .A(n1259), .Z(n1383) );
  CND2X1 U1558 ( .A(n1383), .B(n3080), .Z(n1409) );
  CIVX1 U1559 ( .A(n1409), .Z(n1141) );
  CNR2X2 U1560 ( .A(n1406), .B(n1141), .Z(n1142) );
  CND2XL U1561 ( .A(n1298), .B(n3112), .Z(n1408) );
  CND2X1 U1562 ( .A(n1227), .B(n3113), .Z(n1407) );
  CND3X2 U1563 ( .A(n1142), .B(n1408), .C(n1407), .Z(n1764) );
  CND2X1 U1564 ( .A(n1764), .B(h2[2]), .Z(n1149) );
  CNR2X1 U1565 ( .A(n1416), .B(acc[54]), .Z(n1144) );
  CNR2X1 U1566 ( .A(n1224), .B(acc[57]), .Z(n1143) );
  CNR2X2 U1567 ( .A(n1144), .B(n1143), .Z(n1147) );
  CND2X1 U1568 ( .A(n1227), .B(n3083), .Z(n1146) );
  CND2X1 U1569 ( .A(n1228), .B(n2929), .Z(n1145) );
  CND3X2 U1570 ( .A(n1147), .B(n1146), .C(n1145), .Z(n1748) );
  CND2X1 U1571 ( .A(n1748), .B(n1752), .Z(n1148) );
  CND3X2 U1572 ( .A(n1150), .B(n1148), .C(n1149), .Z(n2226) );
  CND2IX1 U1573 ( .B(n1418), .A(acc[40]), .Z(n1153) );
  CND2X2 U1574 ( .A(n1193), .B(acc[39]), .Z(n1152) );
  CND2X2 U1575 ( .A(n1153), .B(n1152), .Z(n1157) );
  CND2X1 U1576 ( .A(n1297), .B(acc[41]), .Z(n1155) );
  CND2X1 U1577 ( .A(n1481), .B(acc[38]), .Z(n1154) );
  CND2X1 U1578 ( .A(n1155), .B(n1154), .Z(n1156) );
  CNR2X2 U1579 ( .A(n1157), .B(n1156), .Z(n1665) );
  CNR2X1 U1580 ( .A(n767), .B(acc[42]), .Z(n1159) );
  CNR2X2 U1581 ( .A(n1224), .B(acc[45]), .Z(n1158) );
  CNR2X2 U1582 ( .A(n1159), .B(n1158), .Z(n1162) );
  CND2X1 U1583 ( .A(n1248), .B(n3094), .Z(n1161) );
  CND2X1 U1584 ( .A(n1228), .B(n3087), .Z(n1160) );
  CND3X2 U1585 ( .A(n1162), .B(n1161), .C(n1160), .Z(n1753) );
  CND2XL U1586 ( .A(n1753), .B(n1754), .Z(n1163) );
  CND2X1 U1587 ( .A(n1164), .B(n1163), .Z(n1165) );
  CIVX2 U1588 ( .A(n1165), .Z(n1179) );
  CNIVX4 U1589 ( .A(n1166), .Z(n1244) );
  CNR2X1 U1590 ( .A(n1244), .B(acc[49]), .Z(n1167) );
  CNR2X2 U1591 ( .A(n1168), .B(n1167), .Z(n1171) );
  CND2X1 U1592 ( .A(n1349), .B(n3116), .Z(n1170) );
  CND2X1 U1593 ( .A(n1193), .B(n3074), .Z(n1169) );
  CND3X2 U1594 ( .A(n1171), .B(n1170), .C(n1169), .Z(n1755) );
  CND2XL U1595 ( .A(n1755), .B(n1824), .Z(n1178) );
  CNR2X1 U1596 ( .A(n1243), .B(acc[50]), .Z(n1173) );
  CNR2X1 U1597 ( .A(n1224), .B(acc[53]), .Z(n1172) );
  CNR2X2 U1598 ( .A(n1173), .B(n1172), .Z(n1176) );
  CND2X1 U1599 ( .A(n1227), .B(n3114), .Z(n1175) );
  CND2X1 U1600 ( .A(n1228), .B(n3115), .Z(n1174) );
  CND3X2 U1601 ( .A(n1176), .B(n1175), .C(n1174), .Z(n1749) );
  CND2X1 U1602 ( .A(n1749), .B(n1941), .Z(n1177) );
  CND3X2 U1603 ( .A(n1179), .B(n1178), .C(n1177), .Z(n2108) );
  CND2X1 U1604 ( .A(n2108), .B(n1825), .Z(n1209) );
  CND2X1 U1605 ( .A(n1248), .B(acc[36]), .Z(n1181) );
  CND2X1 U1606 ( .A(n1193), .B(acc[35]), .Z(n1180) );
  CND2X2 U1607 ( .A(n1181), .B(n1180), .Z(n1185) );
  CND2X1 U1608 ( .A(n1297), .B(acc[37]), .Z(n1183) );
  CND2XL U1609 ( .A(n1298), .B(acc[34]), .Z(n1182) );
  CND2X1 U1610 ( .A(n1183), .B(n1182), .Z(n1184) );
  CNR2X2 U1611 ( .A(n1185), .B(n1184), .Z(n1663) );
  CAN2XL U1612 ( .A(n1344), .B(acc[30]), .Z(n1187) );
  CNR2X1 U1613 ( .A(n1275), .B(n3077), .Z(n1186) );
  CNR2X1 U1614 ( .A(n1187), .B(n1186), .Z(n1190) );
  CND2X1 U1615 ( .A(n1248), .B(acc[32]), .Z(n1189) );
  CND2X1 U1616 ( .A(n1193), .B(acc[31]), .Z(n1188) );
  CND2XL U1617 ( .A(n1743), .B(n1824), .Z(n1191) );
  COND1XL U1618 ( .A(n1663), .B(n1192), .C(n1191), .Z(n1207) );
  CND2X1 U1619 ( .A(n1248), .B(acc[24]), .Z(n1195) );
  CND2X1 U1620 ( .A(n1193), .B(acc[23]), .Z(n1194) );
  CND3X1 U1621 ( .A(n1196), .B(n1195), .C(n1194), .Z(n1654) );
  CND2XL U1622 ( .A(n1654), .B(n1921), .Z(n1205) );
  CNR2X1 U1623 ( .A(n1243), .B(n3076), .Z(n1198) );
  CNR2X1 U1624 ( .A(n3109), .B(n1275), .Z(n1197) );
  CNR2X1 U1625 ( .A(n1198), .B(n1197), .Z(n1203) );
  CND2X1 U1626 ( .A(n1199), .B(acc[28]), .Z(n1202) );
  CND2X1 U1627 ( .A(n1200), .B(acc[27]), .Z(n1201) );
  CND3X2 U1628 ( .A(n1203), .B(n1202), .C(n1201), .Z(n1744) );
  CND2X1 U1629 ( .A(n1744), .B(n1754), .Z(n1204) );
  CND2X1 U1630 ( .A(n1205), .B(n1204), .Z(n1206) );
  CNR2X1 U1631 ( .A(n1207), .B(n1206), .Z(n1871) );
  CND2X1 U1632 ( .A(n1871), .B(n1741), .Z(n1208) );
  CND3X2 U1633 ( .A(n1210), .B(n1209), .C(n1208), .Z(n2299) );
  CNR2X2 U1634 ( .A(n2296), .B(n2299), .Z(n1364) );
  CND2X1 U1635 ( .A(n1307), .B(n3094), .Z(n1216) );
  CNR2X1 U1636 ( .A(n767), .B(acc[43]), .Z(n1211) );
  CIVX2 U1637 ( .A(n1211), .Z(n1215) );
  CND2X1 U1638 ( .A(n1306), .B(n3117), .Z(n1214) );
  CNR2X1 U1639 ( .A(n1244), .B(acc[46]), .Z(n1212) );
  CIVX2 U1640 ( .A(n1212), .Z(n1213) );
  CND4X2 U1641 ( .A(n1216), .B(n1215), .C(n1214), .D(n1213), .Z(n1623) );
  CND2X2 U1642 ( .A(n1623), .B(n1824), .Z(n1220) );
  CND2X4 U1643 ( .A(n1227), .B(n3085), .Z(n1456) );
  CIVX2 U1644 ( .A(n1456), .Z(n1217) );
  CNR2X1 U1645 ( .A(n767), .B(acc[47]), .Z(n1454) );
  COND1X2 U1646 ( .A(n1217), .B(n768), .C(n1941), .Z(n1219) );
  CNR2IX1 U1647 ( .B(n1469), .A(acc[50]), .Z(n1453) );
  CND2X2 U1648 ( .A(n1228), .B(n3116), .Z(n1455) );
  CND3X2 U1649 ( .A(n1220), .B(n1219), .C(n1218), .Z(n1221) );
  CIVX2 U1650 ( .A(n1221), .Z(n2099) );
  CNR2X1 U1651 ( .A(n1416), .B(acc[35]), .Z(n1223) );
  CNR2X1 U1652 ( .A(n1224), .B(acc[38]), .Z(n1222) );
  CNR2X1 U1653 ( .A(n1223), .B(n1222), .Z(n1519) );
  CND2X1 U1654 ( .A(n1520), .B(n1519), .Z(n1446) );
  CIVX2 U1655 ( .A(n1819), .Z(n1766) );
  CNR2X1 U1656 ( .A(n1416), .B(acc[39]), .Z(n1226) );
  CNR2X1 U1657 ( .A(n1224), .B(acc[42]), .Z(n1225) );
  CNR2X2 U1658 ( .A(n1226), .B(n1225), .Z(n1231) );
  CND2X1 U1659 ( .A(n1227), .B(n3079), .Z(n1230) );
  CND2X1 U1660 ( .A(n1228), .B(n3072), .Z(n1229) );
  CND3X2 U1661 ( .A(n1231), .B(n1230), .C(n1229), .Z(n1614) );
  CND2X1 U1662 ( .A(n1614), .B(n1915), .Z(n2097) );
  CND3X2 U1663 ( .A(n2099), .B(n2098), .C(n2097), .Z(n1846) );
  CNR2IX1 U1664 ( .B(n3080), .A(n1238), .Z(n1448) );
  CIVX1 U1665 ( .A(n3119), .Z(n1232) );
  CND2IX1 U1666 ( .B(n1232), .A(n1383), .Z(n1450) );
  CNR2IX1 U1667 ( .B(n3113), .A(n1140), .Z(n1447) );
  CIVXL U1668 ( .A(n1447), .Z(n1233) );
  CND2X2 U1669 ( .A(n1481), .B(n3086), .Z(n1449) );
  CND3XL U1670 ( .A(n1233), .B(n1449), .C(n1917), .Z(n1235) );
  CNR2IX2 U1671 ( .B(acc[63]), .A(n1243), .Z(n1916) );
  CANR1X1 U1672 ( .A(h2[2]), .B(n1916), .C(n963), .Z(n1234) );
  COND1X1 U1673 ( .A(n1236), .B(n1235), .C(n1234), .Z(n1254) );
  CNR2IXL U1674 ( .B(n3083), .A(n1237), .Z(n1240) );
  CNR2IXL U1675 ( .B(n3093), .A(n1238), .Z(n1239) );
  CNR2X1 U1676 ( .A(n1240), .B(n1239), .Z(n1241) );
  CND2IX2 U1677 ( .B(n1242), .A(n1241), .Z(n1942) );
  CND2X1 U1678 ( .A(n1942), .B(n1915), .Z(n1253) );
  CNR2X2 U1679 ( .A(n767), .B(acc[51]), .Z(n1246) );
  CNR2X2 U1680 ( .A(n1244), .B(acc[54]), .Z(n1245) );
  CNR2X2 U1681 ( .A(n1246), .B(n1245), .Z(n1251) );
  CND2X1 U1682 ( .A(n1247), .B(n3114), .Z(n1250) );
  CND2X1 U1683 ( .A(n1248), .B(n3082), .Z(n1249) );
  CND3X2 U1684 ( .A(n1251), .B(n1250), .C(n1249), .Z(n1826) );
  CND2X1 U1685 ( .A(n1826), .B(n1921), .Z(n1252) );
  CND3X2 U1686 ( .A(n1254), .B(n1253), .C(n1252), .Z(n2180) );
  CND2X1 U1687 ( .A(n2180), .B(n1820), .Z(n1255) );
  CND2X2 U1688 ( .A(n1256), .B(n1255), .Z(n2517) );
  CND2IXL U1689 ( .B(n1418), .A(acc[29]), .Z(n1258) );
  CIVXL U1690 ( .A(n1259), .Z(n1265) );
  CND2XL U1691 ( .A(n1265), .B(acc[30]), .Z(n1261) );
  CND2X1 U1692 ( .A(n1481), .B(acc[27]), .Z(n1260) );
  CNR2X2 U1693 ( .A(n1522), .B(n1523), .Z(n1459) );
  CNR2X2 U1694 ( .A(n1459), .B(n1262), .Z(n1851) );
  CNR2X1 U1695 ( .A(n1851), .B(n1511), .Z(n1281) );
  CND2XL U1696 ( .A(n1306), .B(n3077), .Z(n1264) );
  CND2X1 U1697 ( .A(n1307), .B(n3095), .Z(n1263) );
  CND2X1 U1698 ( .A(n1264), .B(n1263), .Z(n1526) );
  CND2XL U1699 ( .A(n1344), .B(n3062), .Z(n1266) );
  CND2X1 U1700 ( .A(n1267), .B(n1266), .Z(n1524) );
  CND2X1 U1701 ( .A(n1613), .B(n1941), .Z(n1853) );
  CNR2XL U1702 ( .A(n1480), .B(n3098), .Z(n1269) );
  CNR2X1 U1703 ( .A(n1269), .B(n1268), .Z(n1848) );
  CNR2X1 U1704 ( .A(n3100), .B(n1275), .Z(n1271) );
  CNR2X1 U1705 ( .A(n1416), .B(n3102), .Z(n1270) );
  CND2XL U1706 ( .A(n1538), .B(n2409), .Z(n1280) );
  CNR2X2 U1707 ( .A(n1386), .B(n3099), .Z(n1274) );
  CNR2X1 U1708 ( .A(n3076), .B(n1275), .Z(n1277) );
  CNR2X1 U1709 ( .A(n1416), .B(n3106), .Z(n1276) );
  CND2X2 U1710 ( .A(n1279), .B(n1278), .Z(n1618) );
  CND2X1 U1711 ( .A(n1618), .B(n1754), .Z(n1852) );
  CND4X1 U1712 ( .A(n1281), .B(n1853), .C(n1280), .D(n1852), .Z(n1317) );
  CND2XL U1713 ( .A(n1306), .B(acc[13]), .Z(n1282) );
  CIVX1 U1714 ( .A(n1282), .Z(n1288) );
  CND2XL U1715 ( .A(n1297), .B(acc[14]), .Z(n1284) );
  CND2X1 U1716 ( .A(n1481), .B(acc[11]), .Z(n1283) );
  CND2X1 U1717 ( .A(n1284), .B(n1283), .Z(n1287) );
  CND2X1 U1718 ( .A(n1307), .B(acc[12]), .Z(n1285) );
  CIVX2 U1719 ( .A(n1285), .Z(n1286) );
  CNR3X2 U1720 ( .A(n1288), .B(n1287), .C(n1286), .Z(n1605) );
  CND2X1 U1721 ( .A(n1605), .B(n1682), .Z(n1314) );
  CND2XL U1722 ( .A(n1306), .B(acc[9]), .Z(n1290) );
  CND2X1 U1723 ( .A(n1307), .B(acc[8]), .Z(n1289) );
  CND2X1 U1724 ( .A(n1290), .B(n1289), .Z(n1294) );
  CND2X1 U1725 ( .A(n1297), .B(acc[10]), .Z(n1292) );
  CND2XL U1726 ( .A(n1298), .B(acc[7]), .Z(n1291) );
  CND2X1 U1727 ( .A(n1292), .B(n1291), .Z(n1293) );
  CNR2X1 U1728 ( .A(n1294), .B(n1293), .Z(n1466) );
  CND2X1 U1729 ( .A(n1466), .B(n1684), .Z(n1313) );
  CND2XL U1730 ( .A(n1306), .B(acc[5]), .Z(n1296) );
  CND2X1 U1731 ( .A(n1307), .B(acc[4]), .Z(n1295) );
  CND2X1 U1732 ( .A(n1296), .B(n1295), .Z(n1302) );
  CND2XL U1733 ( .A(n1297), .B(acc[6]), .Z(n1300) );
  CND2XL U1734 ( .A(n1298), .B(acc[3]), .Z(n1299) );
  CND2X1 U1735 ( .A(n1300), .B(n1299), .Z(n1301) );
  CNR2X1 U1736 ( .A(n1302), .B(n1301), .Z(n1472) );
  CIVX2 U1737 ( .A(n1658), .Z(n1683) );
  CND2XL U1738 ( .A(n1303), .B(acc[18]), .Z(n1305) );
  CND2X1 U1739 ( .A(n1481), .B(acc[15]), .Z(n1304) );
  CND2X1 U1740 ( .A(n1305), .B(n1304), .Z(n1535) );
  CND2X1 U1741 ( .A(n1306), .B(acc[17]), .Z(n1309) );
  CND2X2 U1742 ( .A(n1307), .B(acc[16]), .Z(n1308) );
  CND2X2 U1743 ( .A(n1309), .B(n1308), .Z(n1536) );
  COND11X2 U1744 ( .A(n1683), .B(n1535), .C(n1536), .D(n2016), .Z(n1310) );
  CIVX2 U1745 ( .A(n1310), .Z(n1311) );
  CND4X1 U1746 ( .A(n1314), .B(n1313), .C(n1312), .D(n1311), .Z(n1315) );
  CND2X2 U1747 ( .A(n1317), .B(n1316), .Z(n2519) );
  CNR2X4 U1748 ( .A(n2517), .B(n2519), .Z(n2026) );
  CIVX2 U1749 ( .A(n1825), .Z(n1818) );
  CNR2XL U1750 ( .A(n1318), .B(n1819), .Z(n1319) );
  CND2IX1 U1751 ( .B(n1320), .A(n1319), .Z(n1327) );
  CIVX2 U1752 ( .A(n1321), .Z(n1324) );
  CIVX2 U1753 ( .A(n1322), .Z(n1323) );
  CNR2X2 U1754 ( .A(n1324), .B(n1323), .Z(n1503) );
  CNR2X1 U1755 ( .A(n1496), .B(n1551), .Z(n1325) );
  CND2X2 U1756 ( .A(n1503), .B(n1325), .Z(n1326) );
  CND2X2 U1757 ( .A(n1327), .B(n1326), .Z(n1864) );
  CND4X1 U1758 ( .A(n1500), .B(n1499), .C(n1498), .D(n1497), .Z(n1573) );
  CND2X1 U1759 ( .A(n1573), .B(n1824), .Z(n1329) );
  CND2X1 U1760 ( .A(n1577), .B(n1941), .Z(n1328) );
  CND2X1 U1761 ( .A(n1329), .B(n1328), .Z(n1865) );
  CNR2X2 U1762 ( .A(n1864), .B(n1865), .Z(n1334) );
  CND2X1 U1763 ( .A(n1585), .B(n1941), .Z(n1859) );
  CNR2X1 U1764 ( .A(n1768), .B(n934), .Z(n1330) );
  CND2X2 U1765 ( .A(n1859), .B(n1330), .Z(n1331) );
  CIVX2 U1766 ( .A(n1331), .Z(n1332) );
  CND2X1 U1767 ( .A(n1586), .B(n1824), .Z(n1858) );
  CIVX2 U1768 ( .A(n1551), .Z(n1691) );
  CND2X1 U1769 ( .A(n1634), .B(n1691), .Z(n1860) );
  CND2X1 U1770 ( .A(n1512), .B(n1766), .Z(n1861) );
  CND4X2 U1771 ( .A(n1332), .B(n1858), .C(n1860), .D(n1861), .Z(n1333) );
  COND1X2 U1772 ( .A(n1818), .B(n1334), .C(n1333), .Z(n1363) );
  CND2X1 U1773 ( .A(n1578), .B(n1766), .Z(n1343) );
  CIVX2 U1774 ( .A(n1335), .Z(n1336) );
  CND2X2 U1775 ( .A(n1337), .B(n1336), .Z(n1508) );
  COND1X2 U1776 ( .A(h2[2]), .B(n1508), .C(h2[3]), .Z(n1342) );
  CND3X2 U1777 ( .A(n1340), .B(n1339), .C(n1338), .Z(n1574) );
  CND2X1 U1778 ( .A(n1574), .B(h2[2]), .Z(n1341) );
  CND3X2 U1779 ( .A(n1343), .B(n1342), .C(n1341), .Z(n2139) );
  CND2X2 U1780 ( .A(n2139), .B(n1820), .Z(n1361) );
  CND2XL U1781 ( .A(n1469), .B(acc[7]), .Z(n1346) );
  CND2XL U1782 ( .A(n1344), .B(acc[4]), .Z(n1345) );
  CND2X1 U1783 ( .A(n1346), .B(n1345), .Z(n1488) );
  CIVXL U1784 ( .A(n1488), .Z(n1348) );
  CND2X1 U1785 ( .A(n1347), .B(acc[5]), .Z(n1490) );
  CND2XL U1786 ( .A(n1348), .B(n1490), .Z(n1355) );
  CND2X1 U1787 ( .A(n1349), .B(acc[6]), .Z(n1489) );
  CND2X1 U1788 ( .A(n1721), .B(n1489), .Z(n1354) );
  CNR2XL U1789 ( .A(n1898), .B(n1628), .Z(n1350) );
  CND3XL U1790 ( .A(n1351), .B(n1352), .C(n1350), .Z(n1353) );
  COND1XL U1791 ( .A(n1355), .B(n1354), .C(n1353), .Z(n1359) );
  CND2X2 U1792 ( .A(n1633), .B(n1658), .Z(n1357) );
  CND2X2 U1793 ( .A(n1640), .B(n1682), .Z(n1356) );
  CND3X2 U1794 ( .A(n1357), .B(n1356), .C(n2016), .Z(n1358) );
  COND1X2 U1795 ( .A(n1359), .B(n1358), .C(n2037), .Z(n1360) );
  CND2X2 U1796 ( .A(n1361), .B(n1360), .Z(n1362) );
  CND2X1 U1797 ( .A(n2026), .B(n764), .Z(n2297) );
  CIVX2 U1798 ( .A(n2297), .Z(n2005) );
  CND2X2 U1799 ( .A(n1364), .B(n2005), .Z(n1594) );
  CND3X2 U1800 ( .A(n1701), .B(n1700), .C(n1699), .Z(n1365) );
  CND2X2 U1801 ( .A(n1365), .B(n1691), .Z(n1367) );
  CND2X2 U1802 ( .A(n1715), .B(n1766), .Z(n1366) );
  CND2X2 U1803 ( .A(n1367), .B(n1366), .Z(n1368) );
  CND2X1 U1804 ( .A(n2596), .B(n1941), .Z(n1370) );
  CND2X1 U1805 ( .A(n1903), .B(n1824), .Z(n1369) );
  CND3X2 U1806 ( .A(n1371), .B(n1370), .C(n1369), .Z(n2095) );
  CND2X2 U1807 ( .A(n2095), .B(n1820), .Z(n1380) );
  CND2X2 U1808 ( .A(n1712), .B(n1824), .Z(n1373) );
  CND2X2 U1809 ( .A(n1713), .B(n1941), .Z(n1372) );
  CND2X2 U1810 ( .A(n1373), .B(n1372), .Z(n1374) );
  CIVX2 U1811 ( .A(n1374), .Z(n1378) );
  CND2X1 U1812 ( .A(n1693), .B(n1691), .Z(n1377) );
  CNR2IX2 U1813 ( .B(n1766), .A(n1736), .Z(n1375) );
  CIVX2 U1814 ( .A(n1375), .Z(n1376) );
  CND3X2 U1815 ( .A(n1378), .B(n1377), .C(n1376), .Z(n2094) );
  CND2X2 U1816 ( .A(n1380), .B(n1379), .Z(n1405) );
  CND2X2 U1817 ( .A(n1722), .B(n1682), .Z(n1382) );
  CND2X1 U1818 ( .A(n1725), .B(n1658), .Z(n1381) );
  CND3X1 U1819 ( .A(n1382), .B(n2016), .C(n1381), .Z(n1394) );
  CIVXL U1820 ( .A(n1383), .Z(n1483) );
  CND2XL U1821 ( .A(n1481), .B(n3067), .Z(n1384) );
  COND1XL U1822 ( .A(acc[4]), .B(n1483), .C(n1384), .Z(n1390) );
  CNR2X1 U1823 ( .A(acc[3]), .B(n1385), .Z(n1388) );
  CND2X1 U1824 ( .A(n1347), .B(n3070), .Z(n1387) );
  CND2IX1 U1825 ( .B(n1388), .A(n1387), .Z(n1389) );
  COND1X1 U1826 ( .A(n1390), .B(n1389), .C(n1721), .Z(n1391) );
  COND1X1 U1827 ( .A(n1638), .B(n1392), .C(n1391), .Z(n1393) );
  COND1X1 U1828 ( .A(n1394), .B(n1393), .C(n2037), .Z(n1403) );
  CIVDX2 U1829 ( .A(n1395), .Z0(n1897), .Z1(n2409) );
  CNR2X2 U1830 ( .A(n1724), .B(n1897), .Z(n1396) );
  CNR2X1 U1831 ( .A(n1396), .B(n1511), .Z(n1401) );
  CND2X1 U1832 ( .A(n1732), .B(n1941), .Z(n1788) );
  CND4X2 U1833 ( .A(n1400), .B(n1399), .C(n1398), .D(n1397), .Z(n1720) );
  CND2X1 U1834 ( .A(n1720), .B(n1691), .Z(n1787) );
  CND2XL U1835 ( .A(n1731), .B(n1824), .Z(n1796) );
  CND4X1 U1836 ( .A(n1401), .B(n1788), .C(n1787), .D(n1796), .Z(n1402) );
  CND2X1 U1837 ( .A(n1403), .B(n1402), .Z(n1404) );
  CNR2X2 U1838 ( .A(n1405), .B(n1404), .Z(n2899) );
  CND2X1 U1839 ( .A(n1765), .B(h2[2]), .Z(n1412) );
  CNR2X1 U1840 ( .A(n1406), .B(h2[2]), .Z(n1410) );
  CND4XL U1841 ( .A(n1410), .B(n1409), .C(n1408), .D(n1407), .Z(n1411) );
  CND2X1 U1842 ( .A(n769), .B(n1915), .Z(n1414) );
  CND2X1 U1843 ( .A(n1749), .B(n1921), .Z(n1413) );
  CND3X1 U1844 ( .A(n1415), .B(n1414), .C(n1413), .Z(n2188) );
  CND2X1 U1845 ( .A(n2188), .B(n1820), .Z(n1445) );
  COND2XL U1846 ( .A(n1417), .B(acc[5]), .C(n1416), .D(acc[2]), .Z(n1420) );
  COND2XL U1847 ( .A(n1480), .B(acc[3]), .C(acc[4]), .D(n1418), .Z(n1419) );
  COND1XL U1848 ( .A(n1420), .B(n1419), .C(n1721), .Z(n1421) );
  CND2IXL U1849 ( .B(h2[6]), .A(n1421), .Z(n1425) );
  CND2IX1 U1850 ( .B(n1425), .A(n1424), .Z(n1430) );
  CND2X1 U1851 ( .A(n1426), .B(n1682), .Z(n1427) );
  COND1X1 U1852 ( .A(n1428), .B(n1638), .C(n1427), .Z(n1429) );
  COND1X1 U1853 ( .A(n1430), .B(n1429), .C(n2037), .Z(n1443) );
  CIVX2 U1854 ( .A(n1433), .Z(n1436) );
  CND2X1 U1855 ( .A(n1663), .B(n1766), .Z(n1434) );
  CND3X2 U1856 ( .A(n1436), .B(n1435), .C(n1434), .Z(n2096) );
  CND2X2 U1857 ( .A(n2096), .B(n1825), .Z(n1442) );
  CND2X2 U1858 ( .A(n1438), .B(n1437), .Z(n1657) );
  CND2X2 U1859 ( .A(n1657), .B(n1766), .Z(n1803) );
  CND3X1 U1860 ( .A(n1803), .B(n1802), .C(n1741), .Z(n1439) );
  CIVXL U1861 ( .A(n1439), .Z(n1440) );
  CND2XL U1862 ( .A(n1654), .B(n1754), .Z(n1801) );
  CND2X1 U1863 ( .A(n1744), .B(n1824), .Z(n1800) );
  CND3X1 U1864 ( .A(n1440), .B(n1801), .C(n1800), .Z(n1441) );
  CND3X1 U1865 ( .A(n1443), .B(n1442), .C(n1441), .Z(n1444) );
  CNR2IX2 U1866 ( .B(n1445), .A(n1444), .Z(n2912) );
  CND2X1 U1867 ( .A(n2899), .B(n2912), .Z(n2003) );
  CNR2X1 U1868 ( .A(n2037), .B(n1628), .Z(n2083) );
  CIVX2 U1869 ( .A(n1446), .Z(n1616) );
  CNR2X1 U1870 ( .A(n1809), .B(n1810), .Z(n2077) );
  CNR2X2 U1871 ( .A(n1448), .B(n1447), .Z(n1549) );
  CND2X2 U1872 ( .A(n1450), .B(n1449), .Z(n1550) );
  CIVX2 U1873 ( .A(n1550), .Z(n1451) );
  CND2X2 U1874 ( .A(n1549), .B(n1451), .Z(n1823) );
  CND2X1 U1875 ( .A(n1823), .B(n1941), .Z(n2078) );
  CNR2X1 U1876 ( .A(n2037), .B(n934), .Z(n1452) );
  CND2X1 U1877 ( .A(n1826), .B(n1691), .Z(n2080) );
  CND2X1 U1878 ( .A(n1942), .B(n1824), .Z(n2079) );
  CIVX2 U1879 ( .A(n1453), .Z(n1458) );
  CIVX2 U1880 ( .A(n1454), .Z(n1457) );
  CND4X4 U1881 ( .A(n1458), .B(n1456), .C(n1457), .D(n1455), .Z(n1822) );
  CND2X1 U1882 ( .A(n1822), .B(n1921), .Z(n2081) );
  CIVX3 U1883 ( .A(n1459), .Z(n1611) );
  CND2X1 U1884 ( .A(n1618), .B(n1824), .Z(n1460) );
  CND2X1 U1885 ( .A(n1461), .B(n1460), .Z(n1817) );
  CIVX2 U1886 ( .A(n1847), .Z(n1463) );
  COND1X1 U1887 ( .A(n1463), .B(n1462), .C(n1915), .Z(n1465) );
  COND1XL U1888 ( .A(n1535), .B(n1536), .C(n2409), .Z(n1464) );
  CND2X1 U1889 ( .A(n1465), .B(n1464), .Z(n1816) );
  CND2IX1 U1890 ( .B(n1917), .A(n1605), .Z(n1468) );
  CND2X1 U1891 ( .A(n1468), .B(n1467), .Z(n1532) );
  CND2X1 U1892 ( .A(n1228), .B(acc[0]), .Z(n1471) );
  CND2X1 U1893 ( .A(n1478), .B(acc[1]), .Z(n1470) );
  CIVX2 U1894 ( .A(h2[4]), .Z(n2148) );
  CND2XL U1895 ( .A(n2016), .B(n2148), .Z(n1814) );
  COND1X1 U1896 ( .A(n963), .B(n1532), .C(n1473), .Z(n1475) );
  CND2X2 U1897 ( .A(n1937), .B(n2148), .Z(n2015) );
  CND2X1 U1898 ( .A(n1916), .B(n1921), .Z(n2183) );
  CND2X2 U1899 ( .A(n2016), .B(n1937), .Z(n2171) );
  COND1XL U1900 ( .A(n2015), .B(n2183), .C(n2171), .Z(n1474) );
  CND3X2 U1901 ( .A(n1476), .B(n1475), .C(n1474), .Z(n2029) );
  CND2X1 U1902 ( .A(n1478), .B(n3070), .Z(n1479) );
  COND1XL U1903 ( .A(acc[1]), .B(n1480), .C(n1479), .Z(n1485) );
  CND2XL U1904 ( .A(n1481), .B(n3071), .Z(n1482) );
  COND1XL U1905 ( .A(acc[3]), .B(n1483), .C(n1482), .Z(n1484) );
  COND1XL U1906 ( .A(n1485), .B(n1484), .C(n1721), .Z(n1486) );
  CND3XL U1907 ( .A(n1487), .B(n1486), .C(n2016), .Z(n1495) );
  CIVXL U1908 ( .A(n1640), .Z(n1493) );
  CNR2X1 U1909 ( .A(n1638), .B(n1488), .Z(n1491) );
  CND3XL U1910 ( .A(n1491), .B(n1490), .C(n1489), .Z(n1492) );
  COND1XL U1911 ( .A(n1493), .B(n1683), .C(n1492), .Z(n1494) );
  COND1X1 U1912 ( .A(n1495), .B(n1494), .C(n2037), .Z(n1517) );
  CNR2IX1 U1913 ( .B(n1824), .A(n1496), .Z(n1502) );
  CND4X2 U1914 ( .A(n1500), .B(n1499), .C(n1498), .D(n1497), .Z(n1501) );
  CANR2X2 U1915 ( .A(n1503), .B(n1502), .C(n1941), .D(n1501), .Z(n2089) );
  CND2X1 U1916 ( .A(n1590), .B(n1691), .Z(n2087) );
  CND3X2 U1917 ( .A(n2089), .B(n2088), .C(n2087), .Z(n1504) );
  CND2X2 U1918 ( .A(n1504), .B(n1825), .Z(n1516) );
  CIVXL U1919 ( .A(n1820), .Z(n1510) );
  CND2X2 U1920 ( .A(n1574), .B(n1824), .Z(n1506) );
  CND2X2 U1921 ( .A(n1578), .B(n1691), .Z(n1505) );
  CND2X2 U1922 ( .A(n1506), .B(n1505), .Z(n1507) );
  CIVX2 U1923 ( .A(n1507), .Z(n1841) );
  CND2X1 U1924 ( .A(n1577), .B(n1921), .Z(n1840) );
  CND2X1 U1925 ( .A(n1508), .B(n1941), .Z(n1839) );
  CND2IX2 U1926 ( .B(n1510), .A(n1509), .Z(n1515) );
  CNR2X2 U1927 ( .A(n1633), .B(n1897), .Z(n1833) );
  CNR2X1 U1928 ( .A(n1833), .B(n1511), .Z(n1513) );
  CND2XL U1929 ( .A(n1586), .B(n1941), .Z(n1832) );
  CND2XL U1930 ( .A(n1512), .B(n1754), .Z(n1831) );
  CND2XL U1931 ( .A(n1634), .B(n1824), .Z(n1835) );
  CND4X1 U1932 ( .A(n1513), .B(n1832), .C(n1831), .D(n1835), .Z(n1514) );
  CND4X2 U1933 ( .A(n1517), .B(n1516), .C(n1515), .D(n1514), .Z(n2028) );
  CANR1X1 U1934 ( .A(n2030), .B(n2029), .C(n2028), .Z(n1518) );
  CNR2X1 U1935 ( .A(n1594), .B(n701), .Z(n2861) );
  CND2IXL U1936 ( .B(n1192), .A(n1519), .Z(n1521) );
  CND2IXL U1937 ( .B(n1521), .A(n1520), .Z(n1531) );
  CND2X2 U1938 ( .A(n1618), .B(n2409), .Z(n1529) );
  COND1X1 U1939 ( .A(n1523), .B(n1522), .C(n1915), .Z(n1528) );
  CND2IX1 U1940 ( .B(n1526), .A(n938), .Z(n1527) );
  CND3X2 U1941 ( .A(n1529), .B(n1528), .C(n1527), .Z(n1530) );
  CNR2IX2 U1942 ( .B(n1531), .A(n1530), .Z(n1925) );
  CND2IXL U1943 ( .B(n934), .A(n1925), .Z(n1534) );
  COND1XL U1944 ( .A(h2[3]), .B(n1532), .C(n934), .Z(n1533) );
  CND2X1 U1945 ( .A(n1534), .B(n1533), .Z(n1542) );
  CNR2X1 U1946 ( .A(n1536), .B(n1535), .Z(n1606) );
  COND1XL U1947 ( .A(n1537), .B(n1606), .C(n2037), .Z(n1540) );
  CIVX2 U1948 ( .A(n1538), .Z(n1603) );
  CNR2XL U1949 ( .A(n1603), .B(n1683), .Z(n1539) );
  CNR2X1 U1950 ( .A(n1540), .B(n1539), .Z(n1541) );
  CND2X1 U1951 ( .A(n1542), .B(n1541), .Z(n1599) );
  CND2X2 U1952 ( .A(n1614), .B(n1752), .Z(n1545) );
  CIVX1 U1953 ( .A(n1754), .Z(n1543) );
  CND2IX1 U1954 ( .B(n1543), .A(n1623), .Z(n1544) );
  CND2X2 U1955 ( .A(n1545), .B(n1544), .Z(n1912) );
  CIVXL U1956 ( .A(n1916), .Z(n1546) );
  COND1XL U1957 ( .A(h2[2]), .B(n1546), .C(h2[3]), .Z(n1547) );
  COND1XL U1958 ( .A(n1738), .B(n1547), .C(n2016), .Z(n1548) );
  CANR1XL U1959 ( .A(n1825), .B(n1912), .C(n1548), .Z(n1556) );
  CND2XL U1960 ( .A(n2075), .B(n1820), .Z(n1555) );
  CND2X2 U1961 ( .A(n1822), .B(n1824), .Z(n1553) );
  CND2X1 U1962 ( .A(n1826), .B(n1941), .Z(n1552) );
  CND2X2 U1963 ( .A(n1553), .B(n1552), .Z(n1913) );
  CND2XL U1964 ( .A(n1913), .B(n1825), .Z(n1554) );
  CAN3X1 U1965 ( .A(n1556), .B(n1555), .C(n1554), .Z(n1600) );
  CND2X1 U1966 ( .A(n1599), .B(n1600), .Z(n2512) );
  CENXL U1967 ( .A(n1558), .B(n1557), .Z(n1566) );
  CNR2X1 U1968 ( .A(n3048), .B(n3046), .Z(n2295) );
  CNR2X1 U1969 ( .A(n3044), .B(n3042), .Z(n1562) );
  CND2X1 U1970 ( .A(n2295), .B(n1562), .Z(n1564) );
  COND1X1 U1971 ( .A(n3053), .B(n3054), .C(n3055), .Z(n2906) );
  CNR2X1 U1972 ( .A(n3052), .B(n3050), .Z(n1560) );
  COND1XL U1973 ( .A(n3049), .B(n3050), .C(n3051), .Z(n1559) );
  CANR1X1 U1974 ( .A(n2906), .B(n1560), .C(n1559), .Z(n2007) );
  COND1XL U1975 ( .A(n3045), .B(n3046), .C(n3047), .Z(n2294) );
  COND1XL U1976 ( .A(n3041), .B(n3042), .C(n3043), .Z(n1561) );
  CANR1XL U1977 ( .A(n2294), .B(n1562), .C(n1561), .Z(n1563) );
  COND1X1 U1978 ( .A(n1564), .B(n2007), .C(n1563), .Z(n1958) );
  CIVX2 U1979 ( .A(n1958), .Z(n2863) );
  CND2XL U1980 ( .A(n3091), .B(cmd_2[0]), .Z(n1948) );
  CIVX1 U1981 ( .A(n1948), .Z(n2916) );
  CANR1XL U1982 ( .A(n2917), .B(n1566), .C(n1565), .Z(n1567) );
  CIVX8 U1983 ( .A(n3059), .Z(n2014) );
  CMX2X4 U1984 ( .A0(acc[24]), .A1(z[24]), .S(n2014), .Z(n641) );
  CMX2X2 U1985 ( .A0(acc[11]), .A1(z[11]), .S(n2014), .Z(n654) );
  CAN2XL U1986 ( .A(n3056), .B(n3053), .Z(n1568) );
  CND2XL U1987 ( .A(n1568), .B(n2916), .Z(n1572) );
  CIVXL U1988 ( .A(n2028), .Z(n1570) );
  CND2XL U1989 ( .A(n2030), .B(n2029), .Z(n1569) );
  CND2X1 U1990 ( .A(n1569), .B(n1570), .Z(n2910) );
  COND3XL U1991 ( .A(n1570), .B(n1569), .C(n2910), .D(n2917), .Z(n1571) );
  COND4CX1 U1992 ( .A(n1572), .B(n1571), .C(n3120), .D(n3184), .Z(n633) );
  CIVX1 U1993 ( .A(n2873), .Z(n2436) );
  CIVDX2 U1994 ( .A(h2[4]), .Z0(n989), .Z1(n2816) );
  CND2XL U1995 ( .A(n1573), .B(n1752), .Z(n1576) );
  CND2XL U1996 ( .A(n1574), .B(n1941), .Z(n1575) );
  CND2X1 U1997 ( .A(n1576), .B(n1575), .Z(n1648) );
  CND2XL U1998 ( .A(n1577), .B(n1754), .Z(n1580) );
  CND2XL U1999 ( .A(n1578), .B(n1824), .Z(n1579) );
  CND2X1 U2000 ( .A(n1580), .B(n1579), .Z(n1581) );
  CIVX2 U2001 ( .A(n1581), .Z(n2143) );
  CND2IX1 U2002 ( .B(n1648), .A(n2143), .Z(n1582) );
  CND2X2 U2003 ( .A(n1738), .B(n2016), .Z(n1929) );
  CANR1X1 U2004 ( .A(n2816), .B(n1582), .C(n2056), .Z(n2039) );
  CIVX2 U2005 ( .A(n1583), .Z(n1584) );
  CND2XL U2006 ( .A(n1585), .B(n1754), .Z(n1588) );
  CND2XL U2007 ( .A(n1586), .B(n1752), .Z(n1587) );
  CND3X1 U2008 ( .A(n1589), .B(n1588), .C(n1587), .Z(n1632) );
  CIVX2 U2009 ( .A(n1590), .Z(n1591) );
  CND2X1 U2010 ( .A(n1591), .B(n1824), .Z(n1630) );
  CIVX4 U2011 ( .A(n2015), .Z(n2054) );
  CND2X1 U2012 ( .A(n1630), .B(n2054), .Z(n1592) );
  CNR2X1 U2013 ( .A(n1632), .B(n1592), .Z(n2034) );
  CNR2XL U2014 ( .A(n1647), .B(n1937), .Z(n2063) );
  CNR2X1 U2015 ( .A(n2034), .B(n2063), .Z(n1593) );
  CND2X1 U2016 ( .A(n2039), .B(n1593), .Z(n2253) );
  CIVX1 U2017 ( .A(n2253), .Z(n1947) );
  CIVX2 U2018 ( .A(n2298), .Z(n1596) );
  CIVX2 U2019 ( .A(n1594), .Z(n1595) );
  CND2X2 U2020 ( .A(n1596), .B(n1595), .Z(n2510) );
  CNR2X2 U2021 ( .A(n1598), .B(n1597), .Z(n1601) );
  CND3X2 U2022 ( .A(n1601), .B(n1600), .C(n1599), .Z(n1602) );
  CIVX2 U2023 ( .A(n1602), .Z(n1973) );
  CND2X2 U2024 ( .A(n1603), .B(n1682), .Z(n1604) );
  CIVX1 U2025 ( .A(n2171), .Z(n2149) );
  CND2X2 U2026 ( .A(n1604), .B(n2149), .Z(n1610) );
  CND2X1 U2027 ( .A(n1605), .B(n1721), .Z(n1608) );
  CND2X1 U2028 ( .A(n1606), .B(n1684), .Z(n1607) );
  CND2X1 U2029 ( .A(n1608), .B(n1607), .Z(n1609) );
  CNR2X2 U2030 ( .A(n1610), .B(n1609), .Z(n1622) );
  CND2X2 U2031 ( .A(n1611), .B(n1752), .Z(n1932) );
  CND2X2 U2032 ( .A(n1932), .B(n2057), .Z(n1612) );
  CIVX2 U2033 ( .A(n1612), .Z(n1617) );
  CND2XL U2034 ( .A(n1613), .B(n1691), .Z(n1934) );
  CIVXL U2035 ( .A(n1614), .Z(n1615) );
  CND2X1 U2036 ( .A(n1615), .B(n1941), .Z(n1931) );
  CND2X1 U2037 ( .A(n1616), .B(n1824), .Z(n1933) );
  CND4X2 U2038 ( .A(n1617), .B(n1934), .C(n1931), .D(n1933), .Z(n1621) );
  CIVXL U2039 ( .A(n1618), .Z(n1619) );
  CND2IX1 U2040 ( .B(n1683), .A(n1619), .Z(n1620) );
  CND3X2 U2041 ( .A(n1622), .B(n1621), .C(n1620), .Z(n1629) );
  CANR2X2 U2042 ( .A(n1822), .B(n1915), .C(n1824), .D(n1826), .Z(n2151) );
  CIVX1 U2043 ( .A(n2083), .Z(n1705) );
  CANR1XL U2044 ( .A(n1941), .B(n1942), .C(n1705), .Z(n1624) );
  CND2XL U2045 ( .A(n1623), .B(n1752), .Z(n1944) );
  CIVX2 U2046 ( .A(n1823), .Z(n1625) );
  CND2X1 U2047 ( .A(n1625), .B(n2409), .Z(n1627) );
  CND2XL U2048 ( .A(n1916), .B(n1691), .Z(n1626) );
  CND2X1 U2049 ( .A(n1627), .B(n1626), .Z(n2344) );
  CND2X1 U2050 ( .A(n1630), .B(n2057), .Z(n1631) );
  CIVXL U2051 ( .A(n1633), .Z(n1637) );
  CIVXL U2052 ( .A(n1634), .Z(n1635) );
  CND2X1 U2053 ( .A(n1635), .B(n1658), .Z(n1636) );
  COND1X1 U2054 ( .A(n1638), .B(n1637), .C(n1636), .Z(n1644) );
  CND2X1 U2055 ( .A(n1639), .B(n1682), .Z(n1642) );
  CND2XL U2056 ( .A(n1640), .B(n1721), .Z(n1641) );
  CND3X1 U2057 ( .A(n1642), .B(n1641), .C(n2149), .Z(n1643) );
  CND2IX1 U2058 ( .B(n1646), .A(n1645), .Z(n1651) );
  CIVX2 U2059 ( .A(n1647), .Z(n2410) );
  CND2X1 U2060 ( .A(n1921), .B(n2057), .Z(n1677) );
  CNR2X2 U2061 ( .A(n2410), .B(n1677), .Z(n2142) );
  CND2X1 U2062 ( .A(n2142), .B(n1768), .Z(n1650) );
  CIVX1 U2063 ( .A(n1648), .Z(n2144) );
  CND3XL U2064 ( .A(n2144), .B(n2143), .C(n2083), .Z(n1649) );
  CND3X1 U2065 ( .A(n1651), .B(n1650), .C(n1649), .Z(n2529) );
  CND2X2 U2066 ( .A(n2818), .B(n2529), .Z(n1974) );
  CNR2X1 U2067 ( .A(n1653), .B(n1652), .Z(n1774) );
  CIVXL U2068 ( .A(n1774), .Z(n1656) );
  CIVX2 U2069 ( .A(n1721), .Z(n1770) );
  CIVX2 U2070 ( .A(n1654), .Z(n1776) );
  CND2X1 U2071 ( .A(n1776), .B(n1682), .Z(n1655) );
  COND1XL U2072 ( .A(n1656), .B(n1770), .C(n1655), .Z(n1662) );
  CIVX2 U2073 ( .A(n1657), .Z(n1772) );
  CND2X1 U2074 ( .A(n1772), .B(n1684), .Z(n1660) );
  CND3X1 U2075 ( .A(n1660), .B(n1659), .C(n2149), .Z(n1661) );
  CNR2X2 U2076 ( .A(n1662), .B(n1661), .Z(n1672) );
  CIVXL U2077 ( .A(n1753), .Z(n1664) );
  CND2IX1 U2078 ( .B(n1192), .A(n1664), .Z(n1668) );
  CND2XL U2079 ( .A(n1743), .B(n1752), .Z(n1667) );
  CIVX2 U2080 ( .A(n1665), .Z(n1742) );
  CND2X1 U2081 ( .A(n1742), .B(n1824), .Z(n1666) );
  CND4X2 U2082 ( .A(n1669), .B(n1668), .C(n1667), .D(n1666), .Z(n2053) );
  CNR2X2 U2083 ( .A(n2053), .B(n934), .Z(n1670) );
  CIVX2 U2084 ( .A(n1670), .Z(n1671) );
  CND2X2 U2085 ( .A(n1671), .B(n1672), .Z(n1681) );
  CND2XL U2086 ( .A(n1755), .B(n1752), .Z(n1673) );
  CND2X1 U2087 ( .A(n1674), .B(n1673), .Z(n2058) );
  CIVX1 U2088 ( .A(n2058), .Z(n2170) );
  CND2X1 U2089 ( .A(n769), .B(n1824), .Z(n1676) );
  CND2XL U2090 ( .A(n1749), .B(n1915), .Z(n1675) );
  CND2X1 U2091 ( .A(n1676), .B(n1675), .Z(n2168) );
  CNR2X1 U2092 ( .A(n2168), .B(n1705), .Z(n1679) );
  CIVX2 U2093 ( .A(n1677), .Z(n1706) );
  CND2X1 U2094 ( .A(n1765), .B(n1706), .Z(n2173) );
  CNR2X1 U2095 ( .A(n2173), .B(n2037), .Z(n1678) );
  CANR1X1 U2096 ( .A(n2170), .B(n1679), .C(n1678), .Z(n1680) );
  CND2X2 U2097 ( .A(n1681), .B(n1680), .Z(n1975) );
  COR2X1 U2098 ( .A(n1720), .B(n1537), .Z(n1687) );
  COAN1X1 U2099 ( .A(n1683), .B(n1731), .C(n2149), .Z(n1686) );
  CND3X2 U2100 ( .A(n1687), .B(n1686), .C(n1685), .Z(n1690) );
  CIVXL U2101 ( .A(n1725), .Z(n1688) );
  CNR2X1 U2102 ( .A(n1688), .B(n1770), .Z(n1689) );
  CNR2X2 U2103 ( .A(n1690), .B(n1689), .Z(n1696) );
  CND2X1 U2104 ( .A(n1736), .B(n1691), .Z(n2047) );
  CND2X1 U2105 ( .A(n1732), .B(n2409), .Z(n2044) );
  CIVX1 U2106 ( .A(n2044), .Z(n1692) );
  CNR2IX1 U2107 ( .B(n2057), .A(n1692), .Z(n1694) );
  CIVX2 U2108 ( .A(n1693), .Z(n1730) );
  CND2X2 U2109 ( .A(n1730), .B(n1824), .Z(n2045) );
  CND4X1 U2110 ( .A(n2047), .B(n2046), .C(n1694), .D(n2045), .Z(n1695) );
  CND2X2 U2111 ( .A(n1696), .B(n1695), .Z(n1710) );
  CND2XL U2112 ( .A(n1713), .B(n2409), .Z(n1698) );
  CND2XL U2113 ( .A(n1903), .B(n1941), .Z(n1697) );
  CND2X1 U2114 ( .A(n1698), .B(n1697), .Z(n2049) );
  CIVX1 U2115 ( .A(n2049), .Z(n2163) );
  CND2XL U2116 ( .A(n1715), .B(n1754), .Z(n1704) );
  CND3XL U2117 ( .A(n1701), .B(n1700), .C(n1699), .Z(n1702) );
  CND2X1 U2118 ( .A(n1702), .B(n1824), .Z(n1703) );
  CND2X1 U2119 ( .A(n1704), .B(n1703), .Z(n2161) );
  CNR2X1 U2120 ( .A(n2161), .B(n1705), .Z(n1708) );
  CND2X1 U2121 ( .A(n1900), .B(n1706), .Z(n2165) );
  CNR2X1 U2122 ( .A(n2165), .B(n2037), .Z(n1707) );
  CANR1X1 U2123 ( .A(n2163), .B(n1708), .C(n1707), .Z(n1709) );
  CND2X2 U2124 ( .A(n1710), .B(n1709), .Z(n2828) );
  CND2X2 U2125 ( .A(n1975), .B(n2828), .Z(n1711) );
  CNR2X2 U2126 ( .A(n1974), .B(n1711), .Z(n1786) );
  CND2XL U2127 ( .A(n1713), .B(n1754), .Z(n1714) );
  CND2XL U2128 ( .A(n1715), .B(n1824), .Z(n1718) );
  CND2X1 U2129 ( .A(n1716), .B(n1941), .Z(n1717) );
  CND3X2 U2130 ( .A(n1719), .B(n1718), .C(n1717), .Z(n2157) );
  CIVX2 U2131 ( .A(n1720), .Z(n1723) );
  CANR2X2 U2132 ( .A(n1723), .B(n1775), .C(n933), .D(n1722), .Z(n1728) );
  CANR1X1 U2133 ( .A(n1771), .B(n1724), .C(h2[6]), .Z(n1727) );
  CND2X1 U2134 ( .A(n1725), .B(n1773), .Z(n1726) );
  CND3X2 U2135 ( .A(n1728), .B(n1727), .C(n1726), .Z(n1729) );
  CANR1X2 U2136 ( .A(n1825), .B(n2157), .C(n1729), .Z(n2398) );
  CND2X2 U2137 ( .A(n1730), .B(n1941), .Z(n1735) );
  CND2XL U2138 ( .A(n1731), .B(n1752), .Z(n1734) );
  CND2X1 U2139 ( .A(n1732), .B(n1754), .Z(n1733) );
  CND3X2 U2140 ( .A(n1735), .B(n1734), .C(n1733), .Z(n1905) );
  CND2X1 U2141 ( .A(n1736), .B(n1824), .Z(n1896) );
  CND2X1 U2142 ( .A(n1741), .B(n1896), .Z(n1737) );
  CNR2X1 U2143 ( .A(n1905), .B(n1737), .Z(n1740) );
  CNR2XL U2144 ( .A(n2347), .B(n1738), .Z(n1739) );
  CNR2X1 U2145 ( .A(n1740), .B(n1739), .Z(n2397) );
  CND2X2 U2146 ( .A(n2398), .B(n2397), .Z(n1785) );
  CND2X1 U2147 ( .A(n1888), .B(n1741), .Z(n1762) );
  CND2XL U2148 ( .A(n1742), .B(n1941), .Z(n1747) );
  CND2XL U2149 ( .A(n1743), .B(n1754), .Z(n1746) );
  CND3X1 U2150 ( .A(n1747), .B(n1746), .C(n1745), .Z(n1889) );
  CND2X1 U2151 ( .A(n1748), .B(n1941), .Z(n1751) );
  CND2X1 U2152 ( .A(n1749), .B(n1824), .Z(n1750) );
  CAN2X2 U2153 ( .A(n1751), .B(n1750), .Z(n1760) );
  CND2XL U2154 ( .A(n1753), .B(n1752), .Z(n1757) );
  CND2XL U2155 ( .A(n1755), .B(n1754), .Z(n1756) );
  CND2X1 U2156 ( .A(n1757), .B(n1756), .Z(n1758) );
  CIVX2 U2157 ( .A(n1758), .Z(n1759) );
  CND2X2 U2158 ( .A(n1760), .B(n1759), .Z(n2166) );
  CIVX2 U2159 ( .A(n2166), .Z(n1761) );
  COND2X2 U2160 ( .A(n1762), .B(n1889), .C(n1761), .D(n1818), .Z(n1763) );
  CIVX2 U2161 ( .A(n1763), .Z(n1784) );
  CIVXL U2162 ( .A(n1764), .Z(n1767) );
  CANR2X1 U2163 ( .A(n1767), .B(n1766), .C(n1915), .D(n1765), .Z(n2167) );
  CND2XL U2164 ( .A(n2167), .B(n1820), .Z(n1783) );
  CANR4CX1 U2165 ( .A(n1770), .B(n1769), .C(n2016), .D(n1768), .Z(n1781) );
  CND2X1 U2166 ( .A(n1772), .B(n1771), .Z(n1779) );
  CND2X1 U2167 ( .A(n1774), .B(n1773), .Z(n1778) );
  CND2X1 U2168 ( .A(n1776), .B(n1775), .Z(n1777) );
  CND3XL U2169 ( .A(n1779), .B(n1778), .C(n1777), .Z(n1780) );
  CNR2X1 U2170 ( .A(n1781), .B(n1780), .Z(n1782) );
  CND3X2 U2171 ( .A(n1784), .B(n1783), .C(n1782), .Z(n2401) );
  CNR2X2 U2172 ( .A(n1785), .B(n2401), .Z(n1972) );
  CND3X2 U2173 ( .A(n1973), .B(n1786), .C(n1972), .Z(n2254) );
  CNR2X2 U2174 ( .A(n2510), .B(n690), .Z(n2499) );
  CANR1XL U2175 ( .A(n2816), .B(n2094), .C(n1929), .Z(n2324) );
  CND2XL U2176 ( .A(n1788), .B(n1787), .Z(n1798) );
  CNR2IX1 U2177 ( .B(n2054), .A(n1789), .Z(n1792) );
  CND3X1 U2178 ( .A(n1792), .B(n1791), .C(n1790), .Z(n1794) );
  CND2X1 U2179 ( .A(n1897), .B(n2054), .Z(n1793) );
  CND2X1 U2180 ( .A(n1794), .B(n1793), .Z(n1795) );
  CND2XL U2181 ( .A(n1796), .B(n1795), .Z(n1797) );
  CNR2XL U2182 ( .A(n1798), .B(n1797), .Z(n1799) );
  CANR1X1 U2183 ( .A(h2[5]), .B(n683), .C(n1799), .Z(n2325) );
  CND2X1 U2184 ( .A(n2324), .B(n2325), .Z(n1987) );
  CND2XL U2185 ( .A(n1801), .B(n1800), .Z(n1805) );
  CND3XL U2186 ( .A(n1803), .B(n2054), .C(n1802), .Z(n1804) );
  COAN1XL U2187 ( .A(n1805), .B(n1804), .C(n1940), .Z(n1808) );
  CND2XL U2188 ( .A(n2096), .B(n2057), .Z(n1807) );
  CND2XL U2189 ( .A(n695), .B(h2[5]), .Z(n1806) );
  CND3X1 U2190 ( .A(n1808), .B(n1807), .C(n1806), .Z(n1991) );
  CNR2X2 U2191 ( .A(n1987), .B(n1991), .Z(n2032) );
  CIVXL U2192 ( .A(n1809), .Z(n1813) );
  CIVXL U2193 ( .A(n1810), .Z(n1812) );
  CNR2X1 U2194 ( .A(n934), .B(h2[6]), .Z(n1811) );
  CND3XL U2195 ( .A(n1813), .B(n1812), .C(n1811), .Z(n2036) );
  CIVXL U2196 ( .A(n1814), .Z(n1815) );
  COND1XL U2197 ( .A(n1817), .B(n1816), .C(n1815), .Z(n2038) );
  CNR2XL U2198 ( .A(n1819), .B(n1818), .Z(n1821) );
  CANR2X1 U2199 ( .A(n1822), .B(n1821), .C(n1820), .D(n2183), .Z(n1830) );
  CND3XL U2200 ( .A(n1823), .B(n1941), .C(n1825), .Z(n1829) );
  CND3XL U2201 ( .A(n1942), .B(n1824), .C(n1825), .Z(n1828) );
  CND3XL U2202 ( .A(n1826), .B(n1915), .C(n1825), .Z(n1827) );
  CND4X1 U2203 ( .A(n1830), .B(n1829), .C(n1828), .D(n1827), .Z(n2064) );
  CND2X1 U2204 ( .A(n1832), .B(n1831), .Z(n1837) );
  CIVX1 U2205 ( .A(n1833), .Z(n1834) );
  CND3X1 U2206 ( .A(n1835), .B(n1834), .C(n2054), .Z(n1836) );
  COND1X1 U2207 ( .A(n1837), .B(n1836), .C(n1940), .Z(n1838) );
  CIVX2 U2208 ( .A(n1838), .Z(n1845) );
  CND2X1 U2209 ( .A(n1509), .B(h2[5]), .Z(n1844) );
  CND3XL U2210 ( .A(n2089), .B(n2088), .C(n2087), .Z(n1842) );
  CND2X1 U2211 ( .A(n1842), .B(n2057), .Z(n1843) );
  CND3X2 U2212 ( .A(n1845), .B(n1844), .C(n1843), .Z(n2132) );
  CANR1X1 U2213 ( .A(h2[5]), .B(n2180), .C(n1929), .Z(n1856) );
  CNR3X1 U2214 ( .A(n1851), .B(n1850), .C(n1849), .Z(n1854) );
  CND3X1 U2215 ( .A(n1854), .B(n1853), .C(n1852), .Z(n1855) );
  CND3X2 U2216 ( .A(n1857), .B(n1856), .C(n1855), .Z(n2496) );
  CIVX2 U2217 ( .A(n2496), .Z(n2067) );
  CND2XL U2218 ( .A(n1858), .B(n2054), .Z(n1863) );
  CND3XL U2219 ( .A(n1861), .B(n1859), .C(n1860), .Z(n1862) );
  COAN1X1 U2220 ( .A(n1863), .B(n1862), .C(n1940), .Z(n1870) );
  CIVX2 U2221 ( .A(n1864), .Z(n1867) );
  CIVX2 U2222 ( .A(n1865), .Z(n1866) );
  CND2X2 U2223 ( .A(n1867), .B(n1866), .Z(n2102) );
  CND2X1 U2224 ( .A(n2102), .B(n2057), .Z(n1869) );
  CND2X1 U2225 ( .A(n2139), .B(h2[5]), .Z(n1868) );
  CND3X2 U2226 ( .A(n1870), .B(n1869), .C(n1868), .Z(n2501) );
  CANR1X1 U2227 ( .A(n2054), .B(n1871), .C(n1929), .Z(n1874) );
  CND2X1 U2228 ( .A(n2226), .B(h2[5]), .Z(n1873) );
  CND2X1 U2229 ( .A(n2108), .B(n2057), .Z(n1872) );
  CND3X1 U2230 ( .A(n1874), .B(n1873), .C(n1872), .Z(n2383) );
  CIVX2 U2231 ( .A(n1875), .Z(n1878) );
  CNR2X1 U2232 ( .A(n1876), .B(n2015), .Z(n1877) );
  CANR1X1 U2233 ( .A(n1878), .B(n1877), .C(n1929), .Z(n1887) );
  CIVX2 U2234 ( .A(n1879), .Z(n1882) );
  CIVX2 U2235 ( .A(n1880), .Z(n1881) );
  CND2X2 U2236 ( .A(n1882), .B(n1881), .Z(n2103) );
  CND2X1 U2237 ( .A(n2103), .B(n2057), .Z(n1886) );
  COND1XL U2238 ( .A(n1884), .B(n1883), .C(h2[5]), .Z(n1885) );
  CND3X1 U2239 ( .A(n1887), .B(n1886), .C(n1885), .Z(n2281) );
  CNR2X2 U2240 ( .A(n2383), .B(n2281), .Z(n2031) );
  CNR2X2 U2241 ( .A(n2497), .B(n2244), .Z(n2333) );
  CND2X1 U2242 ( .A(n1888), .B(n2054), .Z(n1890) );
  CIVX2 U2243 ( .A(n1891), .Z(n1893) );
  CND2X2 U2244 ( .A(n1893), .B(n1892), .Z(n1895) );
  CIVX1 U2245 ( .A(n2167), .Z(n2346) );
  CNR2X1 U2246 ( .A(n2346), .B(n1937), .Z(n1894) );
  CNR2X4 U2247 ( .A(n1895), .B(n1894), .Z(n2245) );
  CNR2X1 U2248 ( .A(n1929), .B(n1898), .Z(n1901) );
  CNR2X1 U2249 ( .A(n1929), .B(h2[5]), .Z(n1899) );
  CANR1X1 U2250 ( .A(n1901), .B(n1900), .C(n1899), .Z(n1902) );
  CIVX2 U2251 ( .A(n1906), .Z(n1908) );
  CND2X2 U2252 ( .A(n2157), .B(n2057), .Z(n1907) );
  CND2X2 U2253 ( .A(n1908), .B(n1907), .Z(n2491) );
  CIVX2 U2254 ( .A(n2491), .Z(n1909) );
  CND2X2 U2255 ( .A(n2245), .B(n1909), .Z(n2043) );
  CNR2X4 U2256 ( .A(n1913), .B(n1912), .Z(n2076) );
  CNR2IX2 U2257 ( .B(n2057), .A(n2076), .Z(n1914) );
  CIVX2 U2258 ( .A(n1914), .Z(n1928) );
  CND2XL U2259 ( .A(n1915), .B(h2[5]), .Z(n1920) );
  CANR1X1 U2260 ( .A(n1917), .B(n1916), .C(n963), .Z(n2074) );
  CND2X1 U2261 ( .A(n2074), .B(h2[5]), .Z(n1918) );
  COND1X1 U2262 ( .A(n1920), .B(n1919), .C(n1918), .Z(n1924) );
  CND3XL U2263 ( .A(n1942), .B(n1921), .C(h2[5]), .Z(n1922) );
  CND2X1 U2264 ( .A(n1922), .B(n1940), .Z(n1923) );
  CNR2X2 U2265 ( .A(n1924), .B(n1923), .Z(n1927) );
  CND2X2 U2266 ( .A(n1925), .B(n2054), .Z(n1926) );
  CND3X2 U2267 ( .A(n1928), .B(n1927), .C(n1926), .Z(n2334) );
  CIVX2 U2268 ( .A(n2334), .Z(n2455) );
  CANR1X1 U2269 ( .A(n2816), .B(n2020), .C(n1929), .Z(n2453) );
  CND3X2 U2270 ( .A(n2454), .B(n2455), .C(n2453), .Z(n2062) );
  CNIVXL U2271 ( .A(n2062), .Z(n2489) );
  CNR2X1 U2272 ( .A(n2043), .B(n2489), .Z(n1930) );
  CND2X2 U2273 ( .A(n2333), .B(n1930), .Z(n2259) );
  CIVX2 U2274 ( .A(n2259), .Z(n2745) );
  CND3XL U2275 ( .A(n1932), .B(n1931), .C(n2054), .Z(n1936) );
  CND2X1 U2276 ( .A(n1934), .B(n1933), .Z(n1935) );
  CNR2X1 U2277 ( .A(n1936), .B(n1935), .Z(n1939) );
  CNR2X1 U2278 ( .A(n2344), .B(n1937), .Z(n1938) );
  CNR2X2 U2279 ( .A(n1939), .B(n1938), .Z(n2066) );
  CND2XL U2280 ( .A(n1942), .B(n1941), .Z(n1943) );
  CND2X1 U2281 ( .A(n1944), .B(n1943), .Z(n2147) );
  CIVXL U2282 ( .A(n2748), .Z(n1945) );
  CND3XL U2283 ( .A(n2745), .B(n2499), .C(n1945), .Z(n1946) );
  CNR2X1 U2284 ( .A(n1948), .B(n3120), .Z(n1949) );
  CIVX1 U2285 ( .A(n3000), .Z(n2370) );
  CND2X1 U2286 ( .A(n2370), .B(n2997), .Z(n1969) );
  CNR2X1 U2287 ( .A(n3024), .B(n3022), .Z(n2275) );
  CNR2X1 U2288 ( .A(n3020), .B(n3018), .Z(n1960) );
  CND2X1 U2289 ( .A(n2275), .B(n1960), .Z(n2336) );
  CNR2X1 U2290 ( .A(n3016), .B(n3014), .Z(n2339) );
  CNR2X1 U2291 ( .A(n3012), .B(n3010), .Z(n1962) );
  CND2X1 U2292 ( .A(n2339), .B(n1962), .Z(n1964) );
  CNR2X1 U2293 ( .A(n2336), .B(n1964), .Z(n2459) );
  CIVX1 U2294 ( .A(n2459), .Z(n2843) );
  CNR2X1 U2295 ( .A(n3008), .B(n3006), .Z(n2749) );
  CNR2X1 U2296 ( .A(n3004), .B(n3002), .Z(n1965) );
  CND2X1 U2297 ( .A(n2749), .B(n1965), .Z(n2263) );
  CNR2XL U2298 ( .A(n2843), .B(n2263), .Z(n1967) );
  CNR2X1 U2299 ( .A(n3040), .B(n3038), .Z(n2820) );
  CNR2X1 U2300 ( .A(n3036), .B(n3034), .Z(n1951) );
  CND2X1 U2301 ( .A(n2820), .B(n1951), .Z(n2532) );
  CNR2X1 U2302 ( .A(n3032), .B(n3030), .Z(n1978) );
  CNR2X1 U2303 ( .A(n3028), .B(n3026), .Z(n1953) );
  CND2X1 U2304 ( .A(n1978), .B(n1953), .Z(n1955) );
  CNR2X1 U2305 ( .A(n2532), .B(n1955), .Z(n1957) );
  COND1X1 U2306 ( .A(n3037), .B(n3038), .C(n3039), .Z(n2821) );
  COND1XL U2307 ( .A(n3033), .B(n3034), .C(n3035), .Z(n1950) );
  CANR1X1 U2308 ( .A(n2821), .B(n1951), .C(n1950), .Z(n2531) );
  COND1XL U2309 ( .A(n3029), .B(n3030), .C(n3031), .Z(n1977) );
  COND1XL U2310 ( .A(n3025), .B(n3026), .C(n3027), .Z(n1952) );
  CANR1XL U2311 ( .A(n1977), .B(n1953), .C(n1952), .Z(n1954) );
  COND1XL U2312 ( .A(n1955), .B(n2531), .C(n1954), .Z(n1956) );
  CANR1X1 U2313 ( .A(n1958), .B(n1957), .C(n1956), .Z(n2119) );
  CIVX2 U2314 ( .A(n2119), .Z(n2853) );
  COND1X1 U2315 ( .A(n3021), .B(n3022), .C(n3023), .Z(n2276) );
  COND1X1 U2316 ( .A(n3017), .B(n3018), .C(n3019), .Z(n1959) );
  CANR1X1 U2317 ( .A(n2276), .B(n1960), .C(n1959), .Z(n2337) );
  COND1XL U2318 ( .A(n3013), .B(n3014), .C(n3015), .Z(n2338) );
  COND1XL U2319 ( .A(n3009), .B(n3010), .C(n3011), .Z(n1961) );
  CANR1XL U2320 ( .A(n2338), .B(n1962), .C(n1961), .Z(n1963) );
  CIVX1 U2321 ( .A(n2458), .Z(n2850) );
  COND1X1 U2322 ( .A(n3005), .B(n3006), .C(n3007), .Z(n2750) );
  COND1XL U2323 ( .A(n2263), .B(n2850), .C(n2264), .Z(n1966) );
  CANR1XL U2324 ( .A(n1967), .B(n2853), .C(n1966), .Z(n1968) );
  CEOXL U2325 ( .A(n1969), .B(n1968), .Z(n1971) );
  COND1XL U2326 ( .A(push_2), .B(n3090), .C(n3150), .Z(n1970) );
  CND2XL U2327 ( .A(n1973), .B(n1972), .Z(n2528) );
  CND3XL U2328 ( .A(n2861), .B(n2828), .C(n2827), .Z(n1976) );
  CENXL U2329 ( .A(n1976), .B(n1975), .Z(n1984) );
  CIVXL U2330 ( .A(n2532), .Z(n2830) );
  CND2XL U2331 ( .A(n2830), .B(n1978), .Z(n1980) );
  CIVXL U2332 ( .A(n2531), .Z(n2831) );
  CANR1XL U2333 ( .A(n1978), .B(n2831), .C(n1977), .Z(n1979) );
  CIVX1 U2334 ( .A(n3028), .Z(n2319) );
  CND2X1 U2335 ( .A(n2319), .B(n3025), .Z(n1981) );
  CENX1 U2336 ( .A(n2318), .B(n1981), .Z(n1982) );
  CAN2XL U2337 ( .A(n1982), .B(n2916), .Z(n1983) );
  COND4CX1 U2338 ( .A(n2917), .B(n1984), .C(n1983), .D(push_2), .Z(n1986) );
  COAN1XL U2339 ( .A(push_2), .B(n935), .C(n3163), .Z(n1985) );
  CND2X1 U2340 ( .A(n1986), .B(n1985), .Z(n619) );
  CIVXL U2341 ( .A(n2499), .Z(n2283) );
  CIVXL U2342 ( .A(n2323), .Z(n1988) );
  CNR3X1 U2343 ( .A(n2283), .B(n1987), .C(n1988), .Z(n1990) );
  CIVXL U2344 ( .A(n1991), .Z(n1989) );
  CND2XL U2345 ( .A(n1990), .B(n1989), .Z(n1994) );
  CIVXL U2346 ( .A(n1990), .Z(n1992) );
  CND2X1 U2347 ( .A(n1992), .B(n1991), .Z(n1993) );
  CND2X1 U2348 ( .A(n1993), .B(n1994), .Z(n2001) );
  CIVXL U2349 ( .A(n3020), .Z(n1995) );
  CND2XL U2350 ( .A(n1995), .B(n3017), .Z(n1997) );
  CANR1XL U2351 ( .A(n2275), .B(n2853), .C(n2276), .Z(n1996) );
  CEOXL U2352 ( .A(n1997), .B(n1996), .Z(n1999) );
  COND1XL U2353 ( .A(push_2), .B(n3088), .C(n3144), .Z(n1998) );
  CANR1XL U2354 ( .A(n1949), .B(n1999), .C(n1998), .Z(n2000) );
  COND1X1 U2355 ( .A(n2873), .B(n2001), .C(n2000), .Z(n615) );
  CAN3X1 U2356 ( .A(n3092), .B(n3091), .C(push_2), .Z(n2002) );
  CMX2XL U2357 ( .A0(n2928), .A1(h[0]), .S(n2921), .Z(n32) );
  CMX2XL U2358 ( .A0(n2927), .A1(h[1]), .S(n2921), .Z(n33) );
  CMX2XL U2359 ( .A0(n2926), .A1(h[2]), .S(n2921), .Z(n34) );
  CMX2XL U2360 ( .A0(n2924), .A1(h[3]), .S(n2921), .Z(n35) );
  CMX2XL U2361 ( .A0(n2925), .A1(h[4]), .S(n2921), .Z(n36) );
  CMX2XL U2362 ( .A0(n2923), .A1(h[5]), .S(n2921), .Z(n37) );
  CMX2XL U2363 ( .A0(n2922), .A1(h[6]), .S(n2921), .Z(n38) );
  CMX2XL U2364 ( .A0(h1[5]), .A1(h2[5]), .S(rst), .Z(n563) );
  CNIVXL U2365 ( .A(n2003), .Z(n2004) );
  CNR2X1 U2366 ( .A(n2910), .B(n2004), .Z(n2904) );
  CND2X1 U2367 ( .A(n2904), .B(n2005), .Z(n2006) );
  CEOXL U2368 ( .A(n2296), .B(n2006), .Z(n2011) );
  CIVX1 U2369 ( .A(n3048), .Z(n2522) );
  CIVX1 U2370 ( .A(n2007), .Z(n2524) );
  CEOX1 U2371 ( .A(n2009), .B(n2008), .Z(n2010) );
  CANR2X1 U2372 ( .A(n2011), .B(n2917), .C(n2916), .D(n2010), .Z(n2012) );
  COND1X1 U2373 ( .A(n3120), .B(n2012), .C(n3164), .Z(n628) );
  CMX2XL U2374 ( .A0(acc[8]), .A1(z[8]), .S(n2014), .Z(n657) );
  CMX2XL U2375 ( .A0(acc[7]), .A1(z[7]), .S(n2014), .Z(n658) );
  CMX2XL U2376 ( .A0(acc[6]), .A1(z[6]), .S(n2014), .Z(n659) );
  CMX2XL U2377 ( .A0(acc[4]), .A1(z[4]), .S(n2014), .Z(n661) );
  CMX2XL U2378 ( .A0(acc[3]), .A1(z[3]), .S(n2014), .Z(n662) );
  CMX2XL U2379 ( .A0(acc[1]), .A1(z[1]), .S(n2014), .Z(n664) );
  CMX2XL U2380 ( .A0(acc[18]), .A1(z[18]), .S(n2014), .Z(n647) );
  CMX2XL U2381 ( .A0(acc[15]), .A1(z[15]), .S(n2014), .Z(n650) );
  CMX2XL U2382 ( .A0(acc[16]), .A1(z[16]), .S(n2014), .Z(n649) );
  CMX2XL U2383 ( .A0(acc[17]), .A1(z[17]), .S(n2014), .Z(n648) );
  CMX2XL U2384 ( .A0(acc[12]), .A1(z[12]), .S(n2014), .Z(n653) );
  CMX2XL U2385 ( .A0(acc[19]), .A1(z[19]), .S(n2014), .Z(n646) );
  CMX2XL U2386 ( .A0(acc[30]), .A1(z[30]), .S(n2014), .Z(n635) );
  CMX2XL U2387 ( .A0(acc[29]), .A1(z[29]), .S(n2014), .Z(n636) );
  CMX2XL U2388 ( .A0(acc[28]), .A1(z[28]), .S(n2014), .Z(n637) );
  CMX2XL U2389 ( .A0(acc[22]), .A1(z[22]), .S(n2014), .Z(n643) );
  CMX2XL U2390 ( .A0(acc[23]), .A1(z[23]), .S(n2014), .Z(n642) );
  CMX2XL U2391 ( .A0(acc[21]), .A1(z[21]), .S(n2014), .Z(n644) );
  CMX2XL U2392 ( .A0(acc[25]), .A1(z[25]), .S(n2014), .Z(n640) );
  CMX2XL U2393 ( .A0(acc[20]), .A1(z[20]), .S(n2014), .Z(n645) );
  CMX2XL U2394 ( .A0(acc[26]), .A1(z[26]), .S(n2014), .Z(n639) );
  CMX2XL U2395 ( .A0(h1[3]), .A1(h2[3]), .S(rst), .Z(n565) );
  CMX2XL U2396 ( .A0(acc[31]), .A1(z[31]), .S(n2014), .Z(n634) );
  CMX2XL U2397 ( .A0(acc[27]), .A1(z[27]), .S(n2014), .Z(n638) );
  CMX2XL U2398 ( .A0(acc[14]), .A1(z[14]), .S(n2014), .Z(n651) );
  CMX2XL U2399 ( .A0(acc[13]), .A1(z[13]), .S(n2014), .Z(n652) );
  CMX2XL U2400 ( .A0(acc[10]), .A1(z[10]), .S(n2014), .Z(n655) );
  CMX2XL U2401 ( .A0(acc[5]), .A1(z[5]), .S(n2014), .Z(n660) );
  CIVX4 U2402 ( .A(rst), .Z(n3061) );
  CIVX4 U2403 ( .A(n2017), .Z(n2345) );
  CIVX2 U2404 ( .A(n2018), .Z(n2225) );
  CNR2IX2 U2405 ( .B(n2816), .A(n2171), .Z(n2155) );
  CND2X2 U2406 ( .A(n2225), .B(n2155), .Z(n2019) );
  COND1X1 U2407 ( .A(n2345), .B(n2020), .C(n2019), .Z(n2141) );
  CND2X1 U2408 ( .A(n2024), .B(n2023), .Z(n2025) );
  CNR2X2 U2409 ( .A(n2025), .B(n2299), .Z(n2212) );
  CND3X2 U2410 ( .A(n2899), .B(n2026), .C(n2520), .Z(n2027) );
  CIVX2 U2411 ( .A(n2027), .Z(n2211) );
  CND4X1 U2412 ( .A(n2212), .B(n2211), .C(n770), .D(n2912), .Z(n2033) );
  CND2X2 U2413 ( .A(n2032), .B(n2031), .Z(n2213) );
  CNR2X2 U2414 ( .A(n2033), .B(n2213), .Z(n2073) );
  CND3XL U2415 ( .A(n2038), .B(n2037), .C(n2036), .Z(n2040) );
  CND3X1 U2416 ( .A(n2041), .B(n2040), .C(n2039), .Z(n2042) );
  CAN4X1 U2417 ( .A(n2047), .B(n2046), .C(n2045), .D(n2044), .Z(n2048) );
  CANR1XL U2418 ( .A(h2[5]), .B(n2596), .C(n2056), .Z(n2051) );
  COND1XL U2419 ( .A(n2049), .B(n2161), .C(n2057), .Z(n2050) );
  CND3X1 U2420 ( .A(n2052), .B(n2051), .C(n2050), .Z(n2366) );
  CIVX2 U2421 ( .A(n2053), .Z(n2055) );
  CND2X1 U2422 ( .A(n2055), .B(n2054), .Z(n2061) );
  CANR1XL U2423 ( .A(h2[5]), .B(n2691), .C(n2056), .Z(n2060) );
  COND1XL U2424 ( .A(n2058), .B(n2168), .C(n2057), .Z(n2059) );
  CND3X1 U2425 ( .A(n2061), .B(n2060), .C(n2059), .Z(n2261) );
  CNR3X2 U2426 ( .A(n2062), .B(n2366), .C(n2261), .Z(n2070) );
  CNR2X2 U2427 ( .A(n2064), .B(n2063), .Z(n2065) );
  CND3X2 U2428 ( .A(n2067), .B(n2066), .C(n2065), .Z(n2068) );
  CNR3X2 U2429 ( .A(n2068), .B(n2501), .C(n2132), .Z(n2069) );
  CIVX2 U2430 ( .A(n2072), .Z(n2216) );
  CIVX3 U2431 ( .A(n2254), .Z(n2215) );
  CND3X2 U2432 ( .A(n2073), .B(n2216), .C(n2215), .Z(n2668) );
  CNR2X1 U2433 ( .A(n2075), .B(n2074), .Z(n2234) );
  CIVXL U2434 ( .A(n2556), .Z(n2109) );
  CND2X1 U2435 ( .A(n2077), .B(n2017), .Z(n2086) );
  CND4X1 U2436 ( .A(n2081), .B(n2080), .C(n2079), .D(n2078), .Z(n2184) );
  CIVXL U2437 ( .A(n2184), .Z(n2082) );
  CND2XL U2438 ( .A(n2082), .B(n2155), .Z(n2085) );
  CIVX2 U2439 ( .A(n2183), .Z(n2895) );
  CND2X1 U2440 ( .A(n2895), .B(n2083), .Z(n2084) );
  CND3X1 U2441 ( .A(n2086), .B(n2085), .C(n2084), .Z(n2838) );
  CIVXL U2442 ( .A(n1504), .Z(n2090) );
  CND2XL U2443 ( .A(n2090), .B(n2017), .Z(n2093) );
  CIVX2 U2444 ( .A(n2091), .Z(n2181) );
  CND2X1 U2445 ( .A(n2181), .B(n2155), .Z(n2092) );
  CND2X1 U2446 ( .A(n2093), .B(n2092), .Z(n2305) );
  CND2X1 U2447 ( .A(n2838), .B(n2305), .Z(n2579) );
  CIVX2 U2448 ( .A(n682), .Z(n2187) );
  CIVX2 U2449 ( .A(n2155), .Z(n2182) );
  COND2X1 U2450 ( .A(n2182), .B(n694), .C(n2345), .D(n2096), .Z(n2438) );
  CND2X2 U2451 ( .A(n2581), .B(n2438), .Z(n2158) );
  CND3XL U2452 ( .A(n2099), .B(n2098), .C(n2097), .Z(n2100) );
  COND2X2 U2453 ( .A(n2182), .B(n2101), .C(n2100), .D(n2345), .Z(n2446) );
  COND2X1 U2454 ( .A(n2345), .B(n2102), .C(n2182), .D(n2139), .Z(n2448) );
  CIVX2 U2455 ( .A(n2103), .Z(n2104) );
  CND2X1 U2456 ( .A(n2104), .B(n2017), .Z(n2107) );
  CIVX2 U2457 ( .A(n2105), .Z(n2229) );
  CND2X1 U2458 ( .A(n2229), .B(n2155), .Z(n2106) );
  COND2X1 U2459 ( .A(n2182), .B(n2226), .C(n2108), .D(n2345), .Z(n2649) );
  CND2X1 U2460 ( .A(n2645), .B(n2649), .Z(n2160) );
  CIVXL U2461 ( .A(n2793), .Z(n2465) );
  CND2IXL U2462 ( .B(n2109), .A(n2465), .Z(n2110) );
  CNR2XL U2463 ( .A(n2668), .B(n2110), .Z(n2111) );
  CENXL U2464 ( .A(n2141), .B(n2111), .Z(n2131) );
  CNR2X1 U2465 ( .A(n2992), .B(n2990), .Z(n2441) );
  CNR2X1 U2466 ( .A(n2988), .B(n2986), .Z(n2123) );
  CND2X1 U2467 ( .A(n2441), .B(n2123), .Z(n2590) );
  CNR2X1 U2468 ( .A(n2984), .B(n2982), .Z(n2560) );
  CNR2X1 U2469 ( .A(n2980), .B(n2978), .Z(n2125) );
  CND2X1 U2470 ( .A(n2560), .B(n2125), .Z(n2127) );
  CNR2X1 U2471 ( .A(n2590), .B(n2127), .Z(n2470) );
  CNR2X1 U2472 ( .A(n3000), .B(n2998), .Z(n2840) );
  CNR2X1 U2473 ( .A(n2996), .B(n2994), .Z(n2113) );
  CND2X1 U2474 ( .A(n2840), .B(n2113), .Z(n2115) );
  CNR2X1 U2475 ( .A(n2263), .B(n2115), .Z(n2117) );
  CND2XL U2476 ( .A(n2459), .B(n2117), .Z(n2120) );
  COND1XL U2477 ( .A(n2997), .B(n2998), .C(n2999), .Z(n2844) );
  COND1XL U2478 ( .A(n2993), .B(n2994), .C(n2995), .Z(n2112) );
  CANR1XL U2479 ( .A(n2844), .B(n2113), .C(n2112), .Z(n2114) );
  COND1XL U2480 ( .A(n2115), .B(n2264), .C(n2114), .Z(n2116) );
  CANR1XL U2481 ( .A(n2458), .B(n2117), .C(n2116), .Z(n2118) );
  COND1X1 U2482 ( .A(n2120), .B(n2119), .C(n2118), .Z(n2121) );
  CNIVX4 U2483 ( .A(n2121), .Z(n2890) );
  COND1X1 U2484 ( .A(n2989), .B(n2990), .C(n2991), .Z(n2440) );
  COND1XL U2485 ( .A(n2985), .B(n2986), .C(n2987), .Z(n2122) );
  CANR1X1 U2486 ( .A(n2440), .B(n2123), .C(n2122), .Z(n2591) );
  COND1XL U2487 ( .A(n2981), .B(n2982), .C(n2983), .Z(n2558) );
  COND1XL U2488 ( .A(n2977), .B(n2978), .C(n2979), .Z(n2124) );
  CANR1XL U2489 ( .A(n2558), .B(n2125), .C(n2124), .Z(n2126) );
  COND1XL U2490 ( .A(push_2), .B(n3072), .C(n3180), .Z(n2128) );
  CANR1XL U2491 ( .A(n1949), .B(n2129), .C(n2128), .Z(n2130) );
  COND1XL U2492 ( .A(n2873), .B(n2131), .C(n2130), .Z(n593) );
  CIVX1 U2493 ( .A(n3024), .Z(n2328) );
  CND2X1 U2494 ( .A(n2328), .B(n3021), .Z(n2134) );
  CENX1 U2495 ( .A(n2853), .B(n2134), .Z(n2136) );
  COND1XL U2496 ( .A(push_2), .B(n3104), .C(n3146), .Z(n2135) );
  CANR1XL U2497 ( .A(n1949), .B(n2136), .C(n2135), .Z(n2137) );
  COND1X1 U2498 ( .A(n2873), .B(n2138), .C(n2137), .Z(n617) );
  CIVXL U2499 ( .A(n2139), .Z(n2140) );
  CND2X1 U2500 ( .A(n2140), .B(n2017), .Z(n2228) );
  CIVX2 U2501 ( .A(n2632), .Z(n2538) );
  CIVX1 U2502 ( .A(n2142), .Z(n2146) );
  CND3X1 U2503 ( .A(n2144), .B(n2143), .C(n934), .Z(n2145) );
  CIVX2 U2504 ( .A(n2147), .Z(n2150) );
  CND4X1 U2505 ( .A(n2151), .B(n2150), .C(n2149), .D(n2148), .Z(n2153) );
  CND2X1 U2506 ( .A(n2344), .B(n2155), .Z(n2152) );
  CND2X1 U2507 ( .A(n2153), .B(n2152), .Z(n2616) );
  CIVX2 U2508 ( .A(n2791), .Z(n2154) );
  CAN2X1 U2509 ( .A(n2538), .B(n2154), .Z(n2179) );
  CND2XL U2510 ( .A(n2347), .B(n2155), .Z(n2156) );
  COND1X1 U2511 ( .A(n2345), .B(n2157), .C(n2156), .Z(n2635) );
  CND3X1 U2512 ( .A(n2838), .B(n2305), .C(n2635), .Z(n2159) );
  CNR2X2 U2513 ( .A(n2159), .B(n2158), .Z(n2178) );
  CIVX2 U2514 ( .A(n2160), .Z(n2177) );
  CIVXL U2515 ( .A(n2161), .Z(n2162) );
  CANR1X1 U2516 ( .A(n2165), .B(n2164), .C(n2171), .Z(n2464) );
  COND2X1 U2517 ( .A(n2182), .B(n2167), .C(n2166), .D(n2345), .Z(n2542) );
  CND2X1 U2518 ( .A(n2464), .B(n2542), .Z(n2175) );
  CIVXL U2519 ( .A(n2168), .Z(n2169) );
  CND3XL U2520 ( .A(n2170), .B(n2169), .C(n934), .Z(n2172) );
  CANR1X1 U2521 ( .A(n2173), .B(n2172), .C(n2171), .Z(n2466) );
  CNR2X2 U2522 ( .A(n2175), .B(n2174), .Z(n2176) );
  CIVX2 U2523 ( .A(n2868), .Z(n2775) );
  CIVXL U2524 ( .A(n2758), .Z(n2189) );
  CAN2X1 U2525 ( .A(n2181), .B(n2017), .Z(n2483) );
  CNR2X1 U2526 ( .A(n2183), .B(n2182), .Z(n2186) );
  CNR2XL U2527 ( .A(n2184), .B(n2345), .Z(n2185) );
  COR2X2 U2528 ( .A(n2186), .B(n2185), .Z(n2548) );
  CND2X2 U2529 ( .A(n2483), .B(n2548), .Z(n2656) );
  CIVX2 U2530 ( .A(n2656), .Z(n2233) );
  CND2X1 U2531 ( .A(n2187), .B(n2017), .Z(n2230) );
  CIVX2 U2532 ( .A(n2230), .Z(n2658) );
  CND3XL U2533 ( .A(n2775), .B(n2189), .C(n2756), .Z(n2190) );
  CNR2XL U2534 ( .A(n2668), .B(n2190), .Z(n2191) );
  CIVXL U2535 ( .A(n2191), .Z(n2192) );
  CENXL U2536 ( .A(n2228), .B(n2192), .Z(n2209) );
  CIVX1 U2537 ( .A(n2952), .Z(n2431) );
  CND2X1 U2538 ( .A(n2431), .B(n2949), .Z(n2205) );
  CNR2X1 U2539 ( .A(n2976), .B(n2974), .Z(n2618) );
  CNR2X1 U2540 ( .A(n2972), .B(n2970), .Z(n2194) );
  CND2X1 U2541 ( .A(n2618), .B(n2194), .Z(n2570) );
  CNR2X1 U2542 ( .A(n2968), .B(n2966), .Z(n2549) );
  CNR2X1 U2543 ( .A(n2964), .B(n2962), .Z(n2196) );
  CND2X1 U2544 ( .A(n2549), .B(n2196), .Z(n2198) );
  CNR2X1 U2545 ( .A(n2570), .B(n2198), .Z(n2200) );
  CND2X1 U2546 ( .A(n2470), .B(n2200), .Z(n2877) );
  CNR2X1 U2547 ( .A(n2960), .B(n2958), .Z(n2760) );
  CNR2X1 U2548 ( .A(n2956), .B(n2954), .Z(n2201) );
  CND2X1 U2549 ( .A(n2760), .B(n2201), .Z(n2429) );
  CNR2XL U2550 ( .A(n2877), .B(n2429), .Z(n2203) );
  COND1X1 U2551 ( .A(n2973), .B(n2974), .C(n2975), .Z(n2620) );
  COND1XL U2552 ( .A(n2969), .B(n2970), .C(n2971), .Z(n2193) );
  CANR1X1 U2553 ( .A(n2620), .B(n2194), .C(n2193), .Z(n2569) );
  COND1XL U2554 ( .A(n2965), .B(n2966), .C(n2967), .Z(n2550) );
  COND1XL U2555 ( .A(n2961), .B(n2962), .C(n2963), .Z(n2195) );
  CANR1XL U2556 ( .A(n2550), .B(n2196), .C(n2195), .Z(n2197) );
  COND1XL U2557 ( .A(n2198), .B(n2569), .C(n2197), .Z(n2199) );
  CANR1X1 U2558 ( .A(n2471), .B(n2200), .C(n2199), .Z(n2887) );
  COND1XL U2559 ( .A(n2957), .B(n2958), .C(n2959), .Z(n2762) );
  COND1XL U2560 ( .A(n2429), .B(n2887), .C(n2430), .Z(n2202) );
  CANR1XL U2561 ( .A(n2203), .B(n2890), .C(n2202), .Z(n2204) );
  CEOXL U2562 ( .A(n2205), .B(n2204), .Z(n2207) );
  COND1XL U2563 ( .A(push_2), .B(n3114), .C(n3174), .Z(n2206) );
  CANR1XL U2564 ( .A(n1949), .B(n2207), .C(n2206), .Z(n2208) );
  COND1X1 U2565 ( .A(n2873), .B(n2209), .C(n2208), .Z(n581) );
  CND4X1 U2566 ( .A(n2212), .B(n2211), .C(n1518), .D(n2912), .Z(n2214) );
  CNR2X2 U2567 ( .A(n2214), .B(n2213), .Z(n2217) );
  CND3X2 U2568 ( .A(n2217), .B(n2216), .C(n2215), .Z(n2633) );
  CNR3XL U2569 ( .A(n2633), .B(n700), .C(n2218), .Z(n2219) );
  CIVXL U2570 ( .A(n2219), .Z(n2220) );
  CENXL U2571 ( .A(n2227), .B(n2220), .Z(n2224) );
  CIVX1 U2572 ( .A(n2956), .Z(n2763) );
  COND1XL U2573 ( .A(push_2), .B(n3081), .C(n3124), .Z(n2221) );
  CANR1XL U2574 ( .A(n1949), .B(n2222), .C(n2221), .Z(n2223) );
  COND1X1 U2575 ( .A(n2873), .B(n2224), .C(n2223), .Z(n583) );
  CNR2X1 U2576 ( .A(n2710), .B(n2227), .Z(n2232) );
  CNR2X1 U2577 ( .A(n2228), .B(n2758), .Z(n2427) );
  CND2X1 U2578 ( .A(n2229), .B(n2017), .Z(n2707) );
  CNR2X1 U2579 ( .A(n2230), .B(n2707), .Z(n2231) );
  CND4X2 U2580 ( .A(n2233), .B(n2232), .C(n2427), .D(n2231), .Z(n2870) );
  CIVXL U2581 ( .A(n2870), .Z(n2599) );
  CIVXL U2582 ( .A(n2234), .Z(n2235) );
  CNR2X1 U2583 ( .A(n2235), .B(n2345), .Z(n2670) );
  CND2XL U2584 ( .A(n2599), .B(n2670), .Z(n2728) );
  CNR3XL U2585 ( .A(n2633), .B(n699), .C(n2728), .Z(n2236) );
  CIVXL U2586 ( .A(n2236), .Z(n2237) );
  CENXL U2587 ( .A(n2727), .B(n2237), .Z(n2243) );
  CIVX1 U2588 ( .A(n2944), .Z(n2734) );
  CNR2X1 U2589 ( .A(n2952), .B(n2950), .Z(n2716) );
  CNR2X1 U2590 ( .A(n2948), .B(n2946), .Z(n2238) );
  CND2X1 U2591 ( .A(n2716), .B(n2238), .Z(n2239) );
  CNR2X1 U2592 ( .A(n2429), .B(n2239), .Z(n2876) );
  COND1XL U2593 ( .A(n2949), .B(n2950), .C(n2951), .Z(n2714) );
  COND1XL U2594 ( .A(push_2), .B(n3083), .C(n3122), .Z(n2240) );
  CANR1XL U2595 ( .A(n1949), .B(n2241), .C(n2240), .Z(n2242) );
  COND1X1 U2596 ( .A(n2873), .B(n2243), .C(n2242), .Z(n577) );
  CIVXL U2597 ( .A(n2497), .Z(n2273) );
  CEOXL U2598 ( .A(n2246), .B(n2245), .Z(n2252) );
  CIVX1 U2599 ( .A(n3004), .Z(n2751) );
  CND2X1 U2600 ( .A(n2751), .B(n3001), .Z(n2248) );
  CEOXL U2601 ( .A(n2248), .B(n2247), .Z(n2250) );
  COND1XL U2602 ( .A(push_2), .B(n3076), .C(n3139), .Z(n2249) );
  CANR1XL U2603 ( .A(n1949), .B(n2250), .C(n2249), .Z(n2251) );
  COND1X1 U2604 ( .A(n2873), .B(n2252), .C(n2251), .Z(n607) );
  CIVXL U2605 ( .A(n2510), .Z(n2257) );
  CNR2X1 U2606 ( .A(n2748), .B(n2253), .Z(n2365) );
  CIVXL U2607 ( .A(n2366), .Z(n2255) );
  CNR2IXL U2608 ( .B(n2255), .A(n689), .Z(n2256) );
  CND3XL U2609 ( .A(n2257), .B(n2365), .C(n2256), .Z(n2258) );
  CNR2X1 U2610 ( .A(n2258), .B(n2259), .Z(n2260) );
  CIVXL U2611 ( .A(n2996), .Z(n2262) );
  CND2XL U2612 ( .A(n2262), .B(n2993), .Z(n2270) );
  CIVXL U2613 ( .A(n2263), .Z(n2842) );
  CND2XL U2614 ( .A(n2842), .B(n2840), .Z(n2266) );
  CNR2XL U2615 ( .A(n2843), .B(n2266), .Z(n2268) );
  CIVXL U2616 ( .A(n2264), .Z(n2848) );
  CANR1XL U2617 ( .A(n2840), .B(n2848), .C(n2844), .Z(n2265) );
  COND1XL U2618 ( .A(n2266), .B(n2850), .C(n2265), .Z(n2267) );
  CANR1XL U2619 ( .A(n2268), .B(n2853), .C(n2267), .Z(n2269) );
  CEOXL U2620 ( .A(n2270), .B(n2269), .Z(n2272) );
  COND1XL U2621 ( .A(push_2), .B(n937), .C(n3165), .Z(n2271) );
  CNIVX2 U2622 ( .A(n2499), .Z(n2746) );
  CND2XL U2623 ( .A(n2746), .B(n2273), .Z(n2274) );
  CENXL U2624 ( .A(n2274), .B(n2496), .Z(n2280) );
  COND1XL U2625 ( .A(push_2), .B(n3102), .C(n3143), .Z(n2277) );
  CANR1XL U2626 ( .A(n1949), .B(n2278), .C(n2277), .Z(n2279) );
  COND1X1 U2627 ( .A(n2873), .B(n2280), .C(n2279), .Z(n614) );
  CIVXL U2628 ( .A(n2281), .Z(n2382) );
  CNR2X1 U2629 ( .A(n2497), .B(n2282), .Z(n2381) );
  CNR2IXL U2630 ( .B(n2381), .A(n2283), .Z(n2284) );
  CENXL U2631 ( .A(n2382), .B(n2284), .Z(n2293) );
  CIVXL U2632 ( .A(n3014), .Z(n2285) );
  CND2XL U2633 ( .A(n2285), .B(n3015), .Z(n2289) );
  CNR2XL U2634 ( .A(n2336), .B(n3016), .Z(n2287) );
  COND1XL U2635 ( .A(n3016), .B(n2337), .C(n3013), .Z(n2286) );
  CANR1XL U2636 ( .A(n2287), .B(n2853), .C(n2286), .Z(n2288) );
  CEOXL U2637 ( .A(n2289), .B(n2288), .Z(n2291) );
  COND1XL U2638 ( .A(push_2), .B(n3101), .C(n3142), .Z(n2290) );
  CANR1XL U2639 ( .A(n1949), .B(n2291), .C(n2290), .Z(n2292) );
  CANR1XL U2640 ( .A(n2295), .B(n2524), .C(n2294), .Z(n2513) );
  CNR3XL U2641 ( .A(n701), .B(n2297), .C(n2296), .Z(n2300) );
  CIVXL U2642 ( .A(n2917), .Z(n2301) );
  CANR1X1 U2643 ( .A(n2916), .B(n2303), .C(n2302), .Z(n2304) );
  COND1X1 U2644 ( .A(n3120), .B(n2304), .C(n3157), .Z(n627) );
  CIVX2 U2645 ( .A(n2668), .Z(n2837) );
  CND2XL U2646 ( .A(n2837), .B(n2838), .Z(n2306) );
  CEOXL U2647 ( .A(n2306), .B(n687), .Z(n2311) );
  CIVX1 U2648 ( .A(n2992), .Z(n2582) );
  CND2X1 U2649 ( .A(n2582), .B(n2989), .Z(n2307) );
  CENX1 U2650 ( .A(n2890), .B(n2307), .Z(n2309) );
  COND1XL U2651 ( .A(push_2), .B(n3095), .C(n3131), .Z(n2308) );
  CANR1XL U2652 ( .A(n1949), .B(n2309), .C(n2308), .Z(n2310) );
  COND1X1 U2653 ( .A(n2873), .B(n2311), .C(n2310), .Z(n601) );
  CND2XL U2654 ( .A(n2837), .B(n679), .Z(n2312) );
  CEOXL U2655 ( .A(n2312), .B(n2446), .Z(n2316) );
  COND1XL U2656 ( .A(push_2), .B(n3075), .C(n3136), .Z(n2313) );
  CANR1XL U2657 ( .A(n1949), .B(n2314), .C(n2313), .Z(n2315) );
  COND1X1 U2658 ( .A(n2873), .B(n2316), .C(n2315), .Z(n598) );
  CEOXL U2659 ( .A(n2317), .B(n2746), .Z(n2322) );
  CND2XL U2660 ( .A(n2320), .B(n1949), .Z(n2321) );
  COND3XL U2661 ( .A(n2322), .B(n2873), .C(n3147), .D(n2321), .Z(n618) );
  CND2XL U2662 ( .A(n2746), .B(n2323), .Z(n2327) );
  CND2XL U2663 ( .A(n2325), .B(n2324), .Z(n2326) );
  CENXL U2664 ( .A(n2327), .B(n2326), .Z(n2332) );
  COND1XL U2665 ( .A(push_2), .B(n3103), .C(n3145), .Z(n2329) );
  CANR1XL U2666 ( .A(n1949), .B(n2330), .C(n2329), .Z(n2331) );
  COND1X1 U2667 ( .A(n2873), .B(n2332), .C(n2331), .Z(n616) );
  CND2XL U2668 ( .A(n2746), .B(n2333), .Z(n2335) );
  CENXL U2669 ( .A(n2335), .B(n766), .Z(n2343) );
  CIVXL U2670 ( .A(n2336), .Z(n2503) );
  CND2XL U2671 ( .A(n2503), .B(n2339), .Z(n2386) );
  CIVXL U2672 ( .A(n2337), .Z(n2502) );
  CANR1XL U2673 ( .A(n2339), .B(n2502), .C(n2338), .Z(n2387) );
  COND1XL U2674 ( .A(push_2), .B(n3106), .C(n3149), .Z(n2340) );
  CANR1XL U2675 ( .A(n1949), .B(n2341), .C(n2340), .Z(n2342) );
  COND1X1 U2676 ( .A(n2873), .B(n2343), .C(n2342), .Z(n610) );
  CND2X1 U2677 ( .A(n2346), .B(n2017), .Z(n2777) );
  CIVX1 U2678 ( .A(n2777), .Z(n2406) );
  CND2X1 U2679 ( .A(n2347), .B(n2017), .Z(n2731) );
  CNR2X1 U2680 ( .A(n2727), .B(n2731), .Z(n2348) );
  CND2X1 U2681 ( .A(n2670), .B(n2348), .Z(n2598) );
  CNR2X1 U2682 ( .A(n2870), .B(n2598), .Z(n2774) );
  CENXL U2683 ( .A(n2405), .B(n2349), .Z(n2364) );
  CIVXL U2684 ( .A(n2938), .Z(n2350) );
  CND2XL U2685 ( .A(n2350), .B(n2939), .Z(n2360) );
  CNR2X1 U2686 ( .A(n2944), .B(n2942), .Z(n2780) );
  CIVXL U2687 ( .A(n2780), .Z(n2351) );
  CNR2XL U2688 ( .A(n2351), .B(n2940), .Z(n2354) );
  CND2XL U2689 ( .A(n2876), .B(n2354), .Z(n2356) );
  CNR2XL U2690 ( .A(n2877), .B(n2356), .Z(n2358) );
  COND1XL U2691 ( .A(n2941), .B(n2942), .C(n2943), .Z(n2779) );
  CIVXL U2692 ( .A(n2779), .Z(n2352) );
  COND1XL U2693 ( .A(n2940), .B(n2352), .C(n2937), .Z(n2353) );
  CANR1XL U2694 ( .A(n2354), .B(n2884), .C(n2353), .Z(n2355) );
  COND1XL U2695 ( .A(n2356), .B(n2887), .C(n2355), .Z(n2357) );
  CANR1XL U2696 ( .A(n2358), .B(n2890), .C(n2357), .Z(n2359) );
  CEOXL U2697 ( .A(n2360), .B(n2359), .Z(n2362) );
  COND1XL U2698 ( .A(push_2), .B(n3086), .C(n3171), .Z(n2361) );
  CANR1XL U2699 ( .A(n1949), .B(n2362), .C(n2361), .Z(n2363) );
  COND1XL U2700 ( .A(n2873), .B(n2364), .C(n2363), .Z(n574) );
  CND3XL U2701 ( .A(n2746), .B(n2745), .C(n2365), .Z(n2367) );
  CENXL U2702 ( .A(n2367), .B(n763), .Z(n2380) );
  CIVXL U2703 ( .A(n2998), .Z(n2368) );
  CND2XL U2704 ( .A(n2368), .B(n2999), .Z(n2376) );
  CND2XL U2705 ( .A(n2842), .B(n2370), .Z(n2372) );
  CNR2XL U2706 ( .A(n2843), .B(n2372), .Z(n2374) );
  CIVXL U2707 ( .A(n2997), .Z(n2369) );
  CANR1XL U2708 ( .A(n2370), .B(n2848), .C(n2369), .Z(n2371) );
  COND1XL U2709 ( .A(n2372), .B(n2850), .C(n2371), .Z(n2373) );
  CANR1XL U2710 ( .A(n2374), .B(n2853), .C(n2373), .Z(n2375) );
  CEOXL U2711 ( .A(n2376), .B(n2375), .Z(n2378) );
  COND1XL U2712 ( .A(push_2), .B(n3109), .C(n3166), .Z(n2377) );
  CANR1XL U2713 ( .A(n1949), .B(n2378), .C(n2377), .Z(n2379) );
  CND3XL U2714 ( .A(n2746), .B(n2382), .C(n2381), .Z(n2384) );
  CENXL U2715 ( .A(n2384), .B(n2383), .Z(n2395) );
  CIVXL U2716 ( .A(n3012), .Z(n2385) );
  CND2XL U2717 ( .A(n2385), .B(n3009), .Z(n2391) );
  CIVXL U2718 ( .A(n2386), .Z(n2389) );
  CIVXL U2719 ( .A(n2387), .Z(n2388) );
  CANR1XL U2720 ( .A(n2389), .B(n2853), .C(n2388), .Z(n2390) );
  CEOXL U2721 ( .A(n2391), .B(n2390), .Z(n2393) );
  COND1XL U2722 ( .A(push_2), .B(n3100), .C(n3141), .Z(n2392) );
  CANR1XL U2723 ( .A(n1949), .B(n2393), .C(n2392), .Z(n2394) );
  CND2XL U2724 ( .A(n2398), .B(n2397), .Z(n2862) );
  CNR2X1 U2725 ( .A(n2860), .B(n2862), .Z(n2399) );
  CNR2IX1 U2726 ( .B(n2399), .A(n688), .Z(n2400) );
  CENXL U2727 ( .A(n2401), .B(n2400), .Z(n2403) );
  CIVX1 U2728 ( .A(n3036), .Z(n2822) );
  COND4CXL U2729 ( .A(n2917), .B(n2403), .C(n2402), .D(push_2), .Z(n2404) );
  CND2XL U2730 ( .A(n2404), .B(n3155), .Z(n623) );
  CIVXL U2731 ( .A(n2774), .Z(n2407) );
  CND2X1 U2732 ( .A(n2406), .B(n2405), .Z(n2597) );
  CIVX2 U2733 ( .A(n2633), .Z(n2795) );
  CND2XL U2734 ( .A(n2795), .B(n2408), .Z(n2411) );
  CND2X1 U2735 ( .A(n2017), .B(n2409), .Z(n2690) );
  CNR2X1 U2736 ( .A(n2410), .B(n2690), .Z(n2687) );
  CEOXL U2737 ( .A(n2411), .B(n2687), .Z(n2426) );
  CIVXL U2738 ( .A(n2936), .Z(n2412) );
  CND2XL U2739 ( .A(n2412), .B(n2933), .Z(n2422) );
  CNR2X1 U2740 ( .A(n2940), .B(n2938), .Z(n2414) );
  CND2X1 U2741 ( .A(n2780), .B(n2414), .Z(n2875) );
  CIVXL U2742 ( .A(n2875), .Z(n2416) );
  CND2XL U2743 ( .A(n2876), .B(n2416), .Z(n2418) );
  CNR2XL U2744 ( .A(n2877), .B(n2418), .Z(n2420) );
  COND1XL U2745 ( .A(n2937), .B(n2938), .C(n2939), .Z(n2413) );
  CANR1XL U2746 ( .A(n2779), .B(n2414), .C(n2413), .Z(n2881) );
  CIVXL U2747 ( .A(n2881), .Z(n2415) );
  CANR1XL U2748 ( .A(n2416), .B(n2884), .C(n2415), .Z(n2417) );
  COND1XL U2749 ( .A(n2418), .B(n2887), .C(n2417), .Z(n2419) );
  CANR1XL U2750 ( .A(n2420), .B(n2890), .C(n2419), .Z(n2421) );
  CEOXL U2751 ( .A(n2422), .B(n2421), .Z(n2424) );
  COND1XL U2752 ( .A(push_2), .B(n3113), .C(n3172), .Z(n2423) );
  CANR1XL U2753 ( .A(n1949), .B(n2424), .C(n2423), .Z(n2425) );
  COND1X1 U2754 ( .A(n2873), .B(n2426), .C(n2425), .Z(n573) );
  CNR3X1 U2755 ( .A(n2633), .B(n699), .C(n2708), .Z(n2428) );
  CENXL U2756 ( .A(n2707), .B(n2428), .Z(n2435) );
  CIVXL U2757 ( .A(n2429), .Z(n2713) );
  CIVXL U2758 ( .A(n2430), .Z(n2715) );
  COND1XL U2759 ( .A(push_2), .B(n3082), .C(n3123), .Z(n2432) );
  CAOR1XL U2760 ( .A(n1949), .B(n2433), .C(n2432), .Z(n2434) );
  CAOR1XL U2761 ( .A(n2436), .B(n2435), .C(n2434), .Z(n580) );
  CIVXL U2762 ( .A(n2579), .Z(n2437) );
  CND2XL U2763 ( .A(n2837), .B(n939), .Z(n2439) );
  CEOXL U2764 ( .A(n2439), .B(n2438), .Z(n2445) );
  COND1XL U2765 ( .A(push_2), .B(n3118), .C(n3181), .Z(n2442) );
  CANR1XL U2766 ( .A(n1949), .B(n2443), .C(n2442), .Z(n2444) );
  COND1X1 U2767 ( .A(n2873), .B(n2445), .C(n2444), .Z(n599) );
  CIVXL U2768 ( .A(n2590), .Z(n2557) );
  CIVXL U2769 ( .A(n2591), .Z(n2559) );
  COND1XL U2770 ( .A(push_2), .B(n3096), .C(n3133), .Z(n2451) );
  CND2XL U2771 ( .A(n2454), .B(n2453), .Z(n2457) );
  CND3XL U2772 ( .A(n2746), .B(n2455), .C(n2333), .Z(n2456) );
  CENXL U2773 ( .A(n2457), .B(n2456), .Z(n2463) );
  COND1XL U2774 ( .A(push_2), .B(n3099), .C(n3140), .Z(n2460) );
  CANR1XL U2775 ( .A(n1949), .B(n2461), .C(n2460), .Z(n2462) );
  COND1X1 U2776 ( .A(n2873), .B(n2463), .C(n2462), .Z(n609) );
  CND3XL U2777 ( .A(n2538), .B(n2542), .C(n2635), .Z(n2792) );
  CIVX2 U2778 ( .A(n2464), .Z(n2797) );
  CIVXL U2779 ( .A(n2466), .Z(n2467) );
  CENXL U2780 ( .A(n2468), .B(n2467), .Z(n2481) );
  CIVXL U2781 ( .A(n2964), .Z(n2469) );
  CND2XL U2782 ( .A(n2469), .B(n2961), .Z(n2477) );
  CIVX1 U2783 ( .A(n2470), .Z(n2800) );
  CIVXL U2784 ( .A(n2570), .Z(n2799) );
  CND2XL U2785 ( .A(n2799), .B(n2549), .Z(n2473) );
  CNR2XL U2786 ( .A(n2800), .B(n2473), .Z(n2475) );
  CIVX1 U2787 ( .A(n2471), .Z(n2805) );
  CIVXL U2788 ( .A(n2569), .Z(n2802) );
  CANR1XL U2789 ( .A(n2549), .B(n2802), .C(n2550), .Z(n2472) );
  COND1XL U2790 ( .A(n2473), .B(n2805), .C(n2472), .Z(n2474) );
  CANR1XL U2791 ( .A(n2475), .B(n2890), .C(n2474), .Z(n2476) );
  CEOXL U2792 ( .A(n2477), .B(n2476), .Z(n2479) );
  COND1XL U2793 ( .A(push_2), .B(n3097), .C(n3134), .Z(n2478) );
  CANR1XL U2794 ( .A(n1949), .B(n2479), .C(n2478), .Z(n2480) );
  COND1X1 U2795 ( .A(n2873), .B(n2481), .C(n2480), .Z(n587) );
  CAN2XL U2796 ( .A(n2775), .B(n2548), .Z(n2482) );
  CND2XL U2797 ( .A(n2795), .B(n2482), .Z(n2484) );
  CEOXL U2798 ( .A(n2484), .B(n2483), .Z(n2488) );
  COND1XL U2799 ( .A(push_2), .B(n3116), .C(n3177), .Z(n2485) );
  CANR1XL U2800 ( .A(n1949), .B(n2486), .C(n2485), .Z(n2487) );
  COND1X1 U2801 ( .A(n2873), .B(n2488), .C(n2487), .Z(n585) );
  CENXL U2802 ( .A(n2491), .B(n2490), .Z(n2495) );
  COND1XL U2803 ( .A(push_2), .B(n3105), .C(n3148), .Z(n2492) );
  CANR1XL U2804 ( .A(n1949), .B(n2493), .C(n2492), .Z(n2494) );
  COND1X1 U2805 ( .A(n2873), .B(n2495), .C(n2494), .Z(n608) );
  CNR2XL U2806 ( .A(n2497), .B(n2496), .Z(n2498) );
  CND2XL U2807 ( .A(n2499), .B(n2498), .Z(n2500) );
  CENX1 U2808 ( .A(n2501), .B(n2500), .Z(n2509) );
  CANR1XL U2809 ( .A(n2503), .B(n2853), .C(n2502), .Z(n2504) );
  CEOXL U2810 ( .A(n2505), .B(n2504), .Z(n2507) );
  COND1XL U2811 ( .A(push_2), .B(n3098), .C(n3138), .Z(n2506) );
  CANR1XL U2812 ( .A(n1949), .B(n2507), .C(n2506), .Z(n2508) );
  COND1XL U2813 ( .A(n2873), .B(n2509), .C(n2508), .Z(n613) );
  CNIVXL U2814 ( .A(n2510), .Z(n2511) );
  CEOXL U2815 ( .A(n2512), .B(n2511), .Z(n2515) );
  CANR2XL U2816 ( .A(n2515), .B(n2917), .C(n2916), .D(n2514), .Z(n2516) );
  COND1XL U2817 ( .A(n3120), .B(n2516), .C(n3154), .Z(n626) );
  CDLY1XL U2818 ( .A(n2517), .Z(n2518) );
  CNR2X1 U2819 ( .A(n2518), .B(n2519), .Z(n2905) );
  CND2X1 U2820 ( .A(n2904), .B(n2905), .Z(n2521) );
  CND2X1 U2821 ( .A(n2522), .B(n3045), .Z(n2523) );
  CENX1 U2822 ( .A(n2524), .B(n2523), .Z(n2525) );
  CIVXL U2823 ( .A(n2528), .Z(n2817) );
  CND3XL U2824 ( .A(n2861), .B(n2817), .C(n2818), .Z(n2530) );
  CENXL U2825 ( .A(n2530), .B(n697), .Z(n2534) );
  CIVX1 U2826 ( .A(n3032), .Z(n2832) );
  CANR1XL U2827 ( .A(n2917), .B(n2534), .C(n2533), .Z(n2537) );
  CNR2XL U2828 ( .A(push_2), .B(n3107), .Z(n2535) );
  CNR2XL U2829 ( .A(n3060), .B(n2535), .Z(n2536) );
  COND1XL U2830 ( .A(n3120), .B(n2537), .C(n2536), .Z(n621) );
  CNR2XL U2831 ( .A(n3108), .B(push_2), .Z(n3156) );
  CND2XL U2832 ( .A(n2538), .B(n2635), .Z(n2539) );
  CNR2XL U2833 ( .A(n2793), .B(n2539), .Z(n2540) );
  CNR2IXL U2834 ( .B(n2540), .A(n2668), .Z(n2541) );
  CENXL U2835 ( .A(n2542), .B(n2541), .Z(n2546) );
  CIVX1 U2836 ( .A(n2972), .Z(n2621) );
  COND1XL U2837 ( .A(push_2), .B(n3089), .C(n3179), .Z(n2543) );
  CANR1XL U2838 ( .A(n1949), .B(n2544), .C(n2543), .Z(n2545) );
  COND1XL U2839 ( .A(n2873), .B(n2546), .C(n2545), .Z(n591) );
  CNR2XL U2840 ( .A(n2633), .B(n700), .Z(n2547) );
  CENXL U2841 ( .A(n2548), .B(n2547), .Z(n2554) );
  COND1XL U2842 ( .A(push_2), .B(n3074), .C(n3125), .Z(n2551) );
  CANR1XL U2843 ( .A(n1949), .B(n2552), .C(n2551), .Z(n2553) );
  COND1XL U2844 ( .A(n2873), .B(n2554), .C(n2553), .Z(n586) );
  CNR2XL U2845 ( .A(n2633), .B(n2793), .Z(n2555) );
  CENXL U2846 ( .A(n2556), .B(n2555), .Z(n2564) );
  CND2XL U2847 ( .A(n2557), .B(n2560), .Z(n2650) );
  CANR1XL U2848 ( .A(n2560), .B(n2559), .C(n2558), .Z(n2651) );
  COND1XL U2849 ( .A(push_2), .B(n3073), .C(n3129), .Z(n2561) );
  CANR1XL U2850 ( .A(n1949), .B(n2562), .C(n2561), .Z(n2563) );
  COND1XL U2851 ( .A(n2873), .B(n2564), .C(n2563), .Z(n594) );
  CNR2IXL U2852 ( .B(n2616), .A(n2793), .Z(n2565) );
  CND2IXL U2853 ( .B(n2792), .A(n2565), .Z(n2566) );
  CNR2XL U2854 ( .A(n2633), .B(n2566), .Z(n2567) );
  CENXL U2855 ( .A(n2568), .B(n2567), .Z(n2578) );
  CIVX1 U2856 ( .A(n2968), .Z(n2803) );
  CND2X1 U2857 ( .A(n2803), .B(n2965), .Z(n2574) );
  CNR2XL U2858 ( .A(n2800), .B(n2570), .Z(n2572) );
  COND1XL U2859 ( .A(n2570), .B(n2805), .C(n2569), .Z(n2571) );
  CANR1XL U2860 ( .A(n2572), .B(n2890), .C(n2571), .Z(n2573) );
  CEOXL U2861 ( .A(n2574), .B(n2573), .Z(n2576) );
  COND1XL U2862 ( .A(push_2), .B(n3094), .C(n3127), .Z(n2575) );
  CANR1XL U2863 ( .A(n1949), .B(n2576), .C(n2575), .Z(n2577) );
  COND1XL U2864 ( .A(n2873), .B(n2578), .C(n2577), .Z(n589) );
  CNR2XL U2865 ( .A(n2668), .B(n2579), .Z(n2580) );
  CENXL U2866 ( .A(n685), .B(n2580), .Z(n2586) );
  COND1XL U2867 ( .A(push_2), .B(n3077), .C(n3130), .Z(n2583) );
  CANR1XL U2868 ( .A(n1949), .B(n2584), .C(n2583), .Z(n2585) );
  COND1XL U2869 ( .A(n2873), .B(n2586), .C(n2585), .Z(n600) );
  CNR2XL U2870 ( .A(n2668), .B(n2646), .Z(n2589) );
  CENXL U2871 ( .A(n2645), .B(n2589), .Z(n2595) );
  COND1XL U2872 ( .A(push_2), .B(n3078), .C(n3132), .Z(n2592) );
  CANR1XL U2873 ( .A(n1949), .B(n2593), .C(n2592), .Z(n2594) );
  COND1XL U2874 ( .A(n2873), .B(n2595), .C(n2594), .Z(n596) );
  CNR2XL U2875 ( .A(n2596), .B(n2690), .Z(n2686) );
  CNR2X1 U2876 ( .A(n2598), .B(n2597), .Z(n2688) );
  CND3XL U2877 ( .A(n2599), .B(n2687), .C(n2688), .Z(n2600) );
  CNR3XL U2878 ( .A(n2633), .B(n700), .C(n2600), .Z(n2601) );
  CENXL U2879 ( .A(n2686), .B(n2601), .Z(n2614) );
  CIVX1 U2880 ( .A(n2934), .Z(n2602) );
  CND2X1 U2881 ( .A(n2602), .B(n2935), .Z(n2610) );
  CNR2XL U2882 ( .A(n2875), .B(n2936), .Z(n2604) );
  CND2XL U2883 ( .A(n2876), .B(n2604), .Z(n2606) );
  CNR2XL U2884 ( .A(n2877), .B(n2606), .Z(n2608) );
  COND1XL U2885 ( .A(n2936), .B(n2881), .C(n2933), .Z(n2603) );
  CANR1XL U2886 ( .A(n2604), .B(n2884), .C(n2603), .Z(n2605) );
  COND1XL U2887 ( .A(n2606), .B(n2887), .C(n2605), .Z(n2607) );
  CANR1XL U2888 ( .A(n2608), .B(n2890), .C(n2607), .Z(n2609) );
  CEOXL U2889 ( .A(n2610), .B(n2609), .Z(n2612) );
  COND1XL U2890 ( .A(push_2), .B(n3080), .C(n3175), .Z(n2611) );
  CANR1XL U2891 ( .A(n1949), .B(n2612), .C(n2611), .Z(n2613) );
  COND1XL U2892 ( .A(n2873), .B(n2614), .C(n2613), .Z(n572) );
  CNR3XL U2893 ( .A(n2633), .B(n2793), .C(n2792), .Z(n2615) );
  CENXL U2894 ( .A(n2616), .B(n2615), .Z(n2631) );
  CIVXL U2895 ( .A(n2970), .Z(n2617) );
  CND2XL U2896 ( .A(n2617), .B(n2971), .Z(n2627) );
  CND2XL U2897 ( .A(n2618), .B(n2621), .Z(n2623) );
  CNR2XL U2898 ( .A(n2800), .B(n2623), .Z(n2625) );
  CIVXL U2899 ( .A(n2969), .Z(n2619) );
  CANR1XL U2900 ( .A(n2621), .B(n2620), .C(n2619), .Z(n2622) );
  COND1XL U2901 ( .A(n2623), .B(n2805), .C(n2622), .Z(n2624) );
  CANR1XL U2902 ( .A(n2625), .B(n2890), .C(n2624), .Z(n2626) );
  CEOXL U2903 ( .A(n2627), .B(n2626), .Z(n2629) );
  COND1XL U2904 ( .A(push_2), .B(n3087), .C(n3126), .Z(n2628) );
  CANR1XL U2905 ( .A(n1949), .B(n2629), .C(n2628), .Z(n2630) );
  COND1XL U2906 ( .A(n2873), .B(n2631), .C(n2630), .Z(n590) );
  CNR3XL U2907 ( .A(n2633), .B(n2632), .C(n2793), .Z(n2634) );
  CENXL U2908 ( .A(n2635), .B(n2634), .Z(n2644) );
  CIVXL U2909 ( .A(n2974), .Z(n2636) );
  CND2XL U2910 ( .A(n2636), .B(n2975), .Z(n2640) );
  CNR2XL U2911 ( .A(n2800), .B(n2976), .Z(n2638) );
  COND1XL U2912 ( .A(n2976), .B(n2805), .C(n2973), .Z(n2637) );
  CANR1XL U2913 ( .A(n2638), .B(n2890), .C(n2637), .Z(n2639) );
  CEOXL U2914 ( .A(n2640), .B(n2639), .Z(n2642) );
  COND1XL U2915 ( .A(push_2), .B(n3079), .C(n3128), .Z(n2641) );
  CANR1XL U2916 ( .A(n1949), .B(n2642), .C(n2641), .Z(n2643) );
  COND1XL U2917 ( .A(n2873), .B(n2644), .C(n2643), .Z(n592) );
  CIVXL U2918 ( .A(n2645), .Z(n2647) );
  CNR3XL U2919 ( .A(n2668), .B(n2647), .C(n2646), .Z(n2648) );
  CENXL U2920 ( .A(n2649), .B(n2648), .Z(n2655) );
  COND1XL U2921 ( .A(push_2), .B(n3084), .C(n3135), .Z(n2652) );
  CANR1XL U2922 ( .A(n1949), .B(n2653), .C(n2652), .Z(n2654) );
  COND1XL U2923 ( .A(n2873), .B(n2655), .C(n2654), .Z(n595) );
  CNR3XL U2924 ( .A(n2668), .B(n700), .C(n2656), .Z(n2657) );
  CENXL U2925 ( .A(n2658), .B(n2657), .Z(n2667) );
  CIVXL U2926 ( .A(n2958), .Z(n2659) );
  CND2XL U2927 ( .A(n2659), .B(n2959), .Z(n2663) );
  CNR2XL U2928 ( .A(n2877), .B(n2960), .Z(n2661) );
  COND1XL U2929 ( .A(n2960), .B(n2887), .C(n2957), .Z(n2660) );
  CANR1XL U2930 ( .A(n2661), .B(n2890), .C(n2660), .Z(n2662) );
  CEOXL U2931 ( .A(n2663), .B(n2662), .Z(n2665) );
  COND1XL U2932 ( .A(push_2), .B(n3085), .C(n3168), .Z(n2664) );
  CANR1XL U2933 ( .A(n1949), .B(n2665), .C(n2664), .Z(n2666) );
  COND1XL U2934 ( .A(n2873), .B(n2667), .C(n2666), .Z(n584) );
  CNR3XL U2935 ( .A(n2668), .B(n700), .C(n693), .Z(n2669) );
  CENXL U2936 ( .A(n2670), .B(n2669), .Z(n2685) );
  CIVXL U2937 ( .A(n2946), .Z(n2671) );
  CND2XL U2938 ( .A(n2671), .B(n2947), .Z(n2681) );
  CIVXL U2939 ( .A(n2716), .Z(n2672) );
  CNR2XL U2940 ( .A(n2672), .B(n2948), .Z(n2675) );
  CND2XL U2941 ( .A(n2675), .B(n2713), .Z(n2677) );
  CNR2XL U2942 ( .A(n2877), .B(n2677), .Z(n2679) );
  CIVXL U2943 ( .A(n2714), .Z(n2673) );
  COND1XL U2944 ( .A(n2948), .B(n2673), .C(n2945), .Z(n2674) );
  CANR1XL U2945 ( .A(n2715), .B(n2675), .C(n2674), .Z(n2676) );
  COND1XL U2946 ( .A(n2677), .B(n2887), .C(n2676), .Z(n2678) );
  CANR1XL U2947 ( .A(n2679), .B(n2890), .C(n2678), .Z(n2680) );
  CEOXL U2948 ( .A(n2681), .B(n2680), .Z(n2683) );
  COND1XL U2949 ( .A(push_2), .B(n2929), .C(n3173), .Z(n2682) );
  CANR1XL U2950 ( .A(n1949), .B(n2683), .C(n2682), .Z(n2684) );
  COND1XL U2951 ( .A(n2873), .B(n2685), .C(n2684), .Z(n578) );
  CND3XL U2952 ( .A(n2688), .B(n2687), .C(n2686), .Z(n2872) );
  CNR3XL U2953 ( .A(n700), .B(n693), .C(n2872), .Z(n2689) );
  CND2XL U2954 ( .A(n2689), .B(n2837), .Z(n2692) );
  CNR2X1 U2955 ( .A(n2691), .B(n2690), .Z(n2867) );
  CND2X1 U2956 ( .A(n3058), .B(n2931), .Z(n2702) );
  CNR2X1 U2957 ( .A(n2936), .B(n2934), .Z(n2874) );
  CIVX1 U2958 ( .A(n2874), .Z(n2694) );
  CNR2XL U2959 ( .A(n2875), .B(n2694), .Z(n2696) );
  CND2XL U2960 ( .A(n2876), .B(n2696), .Z(n2698) );
  CNR2XL U2961 ( .A(n2877), .B(n2698), .Z(n2700) );
  COND1XL U2962 ( .A(n2933), .B(n2934), .C(n2935), .Z(n2879) );
  CIVXL U2963 ( .A(n2879), .Z(n2693) );
  COND1XL U2964 ( .A(n2694), .B(n2881), .C(n2693), .Z(n2695) );
  CANR1XL U2965 ( .A(n2696), .B(n2884), .C(n2695), .Z(n2697) );
  COND1XL U2966 ( .A(n2698), .B(n2887), .C(n2697), .Z(n2699) );
  CANR1XL U2967 ( .A(n2700), .B(n2890), .C(n2699), .Z(n2701) );
  CEOXL U2968 ( .A(n2702), .B(n2701), .Z(n2704) );
  COND1XL U2969 ( .A(push_2), .B(n3119), .C(n3182), .Z(n2703) );
  CANR1XL U2970 ( .A(n1949), .B(n2704), .C(n2703), .Z(n2705) );
  CNR3XL U2971 ( .A(n699), .B(n2708), .C(n2707), .Z(n2709) );
  CND2XL U2972 ( .A(n2795), .B(n2709), .Z(n2711) );
  CENXL U2973 ( .A(n2711), .B(n2710), .Z(n2726) );
  CIVXL U2974 ( .A(n2948), .Z(n2712) );
  CND2XL U2975 ( .A(n2712), .B(n2945), .Z(n2722) );
  CND2XL U2976 ( .A(n2713), .B(n2716), .Z(n2718) );
  CNR2XL U2977 ( .A(n2877), .B(n2718), .Z(n2720) );
  CANR1XL U2978 ( .A(n2716), .B(n2715), .C(n2714), .Z(n2717) );
  COND1XL U2979 ( .A(n2718), .B(n2887), .C(n2717), .Z(n2719) );
  CANR1XL U2980 ( .A(n2720), .B(n2890), .C(n2719), .Z(n2721) );
  CEOXL U2981 ( .A(n2722), .B(n2721), .Z(n2724) );
  COND1XL U2982 ( .A(push_2), .B(n3111), .C(n3169), .Z(n2723) );
  CANR1XL U2983 ( .A(n1949), .B(n2724), .C(n2723), .Z(n2725) );
  COND1X1 U2984 ( .A(n2873), .B(n2726), .C(n2725), .Z(n579) );
  CNR3XL U2985 ( .A(n699), .B(n2728), .C(n2727), .Z(n2729) );
  CND2XL U2986 ( .A(n2795), .B(n2729), .Z(n2730) );
  CENXL U2987 ( .A(n2731), .B(n2730), .Z(n2744) );
  CIVXL U2988 ( .A(n2942), .Z(n2732) );
  CND2XL U2989 ( .A(n2732), .B(n2943), .Z(n2740) );
  CND2XL U2990 ( .A(n2876), .B(n2734), .Z(n2736) );
  CNR2XL U2991 ( .A(n2877), .B(n2736), .Z(n2738) );
  CIVXL U2992 ( .A(n2941), .Z(n2733) );
  CANR1XL U2993 ( .A(n2734), .B(n2884), .C(n2733), .Z(n2735) );
  COND1XL U2994 ( .A(n2736), .B(n2887), .C(n2735), .Z(n2737) );
  CANR1XL U2995 ( .A(n2738), .B(n2890), .C(n2737), .Z(n2739) );
  CEOXL U2996 ( .A(n2740), .B(n2739), .Z(n2742) );
  COND1XL U2997 ( .A(push_2), .B(n3093), .C(n3121), .Z(n2741) );
  CANR1XL U2998 ( .A(n1949), .B(n2742), .C(n2741), .Z(n2743) );
  CND2XL U2999 ( .A(n2746), .B(n2745), .Z(n2747) );
  CENXL U3000 ( .A(n2748), .B(n2747), .Z(n2755) );
  COND1XL U3001 ( .A(push_2), .B(n3110), .C(n3167), .Z(n2752) );
  CANR1XL U3002 ( .A(n1949), .B(n2753), .C(n2752), .Z(n2754) );
  CND3XL U3003 ( .A(n2795), .B(n681), .C(n2756), .Z(n2757) );
  CENXL U3004 ( .A(n2758), .B(n2757), .Z(n2773) );
  CIVXL U3005 ( .A(n2954), .Z(n2759) );
  CND2XL U3006 ( .A(n2759), .B(n2955), .Z(n2769) );
  CND2XL U3007 ( .A(n2760), .B(n2763), .Z(n2765) );
  CNR2XL U3008 ( .A(n2877), .B(n2765), .Z(n2767) );
  CIVXL U3009 ( .A(n2953), .Z(n2761) );
  CANR1XL U3010 ( .A(n2763), .B(n2762), .C(n2761), .Z(n2764) );
  COND1XL U3011 ( .A(n2765), .B(n2887), .C(n2764), .Z(n2766) );
  CANR1XL U3012 ( .A(n2767), .B(n2890), .C(n2766), .Z(n2768) );
  CEOXL U3013 ( .A(n2769), .B(n2768), .Z(n2771) );
  COND1XL U3014 ( .A(push_2), .B(n3115), .C(n3176), .Z(n2770) );
  CANR1XL U3015 ( .A(n1949), .B(n2771), .C(n2770), .Z(n2772) );
  CND3XL U3016 ( .A(n2795), .B(n681), .C(n2774), .Z(n2776) );
  CENXL U3017 ( .A(n2777), .B(n2776), .Z(n2790) );
  CIVXL U3018 ( .A(n2940), .Z(n2778) );
  CND2XL U3019 ( .A(n2778), .B(n2937), .Z(n2786) );
  CND2XL U3020 ( .A(n2876), .B(n2780), .Z(n2782) );
  CNR2XL U3021 ( .A(n2877), .B(n2782), .Z(n2784) );
  CANR1XL U3022 ( .A(n2780), .B(n2884), .C(n2779), .Z(n2781) );
  COND1XL U3023 ( .A(n2782), .B(n2887), .C(n2781), .Z(n2783) );
  CANR1XL U3024 ( .A(n2784), .B(n2890), .C(n2783), .Z(n2785) );
  CEOXL U3025 ( .A(n2786), .B(n2785), .Z(n2788) );
  COND1XL U3026 ( .A(push_2), .B(n3112), .C(n3170), .Z(n2787) );
  CANR1XL U3027 ( .A(n1949), .B(n2788), .C(n2787), .Z(n2789) );
  CNR3XL U3028 ( .A(n2793), .B(n2792), .C(n2791), .Z(n2794) );
  CIVXL U3029 ( .A(n2966), .Z(n2798) );
  CND2XL U3030 ( .A(n2798), .B(n2967), .Z(n2810) );
  CND2XL U3031 ( .A(n2799), .B(n2803), .Z(n2806) );
  CNR2XL U3032 ( .A(n2800), .B(n2806), .Z(n2808) );
  CIVXL U3033 ( .A(n2965), .Z(n2801) );
  CANR1XL U3034 ( .A(n2803), .B(n2802), .C(n2801), .Z(n2804) );
  COND1XL U3035 ( .A(n2806), .B(n2805), .C(n2804), .Z(n2807) );
  CANR1XL U3036 ( .A(n2808), .B(n2890), .C(n2807), .Z(n2809) );
  CEOXL U3037 ( .A(n2810), .B(n2809), .Z(n2812) );
  COND1XL U3038 ( .A(push_2), .B(n3117), .C(n3178), .Z(n2811) );
  CANR1XL U3039 ( .A(n1949), .B(n2812), .C(n2811), .Z(n2813) );
  CMX2X1 U3040 ( .A0(h1[6]), .A1(h2[6]), .S(rst), .Z(n562) );
  CMX2X1 U3041 ( .A0(h1[2]), .A1(h2[2]), .S(rst), .Z(n566) );
  CMX2X1 U3042 ( .A0(h1[1]), .A1(n2815), .S(rst), .Z(n567) );
  CMX2X1 U3043 ( .A0(h1[4]), .A1(n2816), .S(rst), .Z(n564) );
  CND2XL U3044 ( .A(n2861), .B(n2817), .Z(n2819) );
  CENXL U3045 ( .A(n2819), .B(n2818), .Z(n2825) );
  CAN2XL U3046 ( .A(n2823), .B(n2916), .Z(n2824) );
  COND4CX1 U3047 ( .A(n2917), .B(n2825), .C(n2824), .D(push_2), .Z(n2826) );
  CND2X1 U3048 ( .A(n2826), .B(n3151), .Z(n622) );
  CND2XL U3049 ( .A(n2861), .B(n2827), .Z(n2829) );
  CENXL U3050 ( .A(n2829), .B(n2828), .Z(n2835) );
  CAN2XL U3051 ( .A(n2833), .B(n2916), .Z(n2834) );
  COND4CX1 U3052 ( .A(n2917), .B(n2835), .C(n2834), .D(push_2), .Z(n2836) );
  CND2X1 U3053 ( .A(n2836), .B(n3162), .Z(n620) );
  CEOXL U3054 ( .A(n2838), .B(n2871), .Z(n2859) );
  CIVXL U3055 ( .A(n2994), .Z(n2839) );
  CND2XL U3056 ( .A(n2839), .B(n2995), .Z(n2856) );
  CIVXL U3057 ( .A(n2840), .Z(n2841) );
  CNR2XL U3058 ( .A(n2841), .B(n2996), .Z(n2847) );
  CND2XL U3059 ( .A(n2847), .B(n2842), .Z(n2851) );
  CNR2XL U3060 ( .A(n2843), .B(n2851), .Z(n2854) );
  CIVXL U3061 ( .A(n2844), .Z(n2845) );
  COND1XL U3062 ( .A(n2996), .B(n2845), .C(n2993), .Z(n2846) );
  CANR1XL U3063 ( .A(n2848), .B(n2847), .C(n2846), .Z(n2849) );
  COND1XL U3064 ( .A(n2851), .B(n2850), .C(n2849), .Z(n2852) );
  CANR1XL U3065 ( .A(n2854), .B(n2853), .C(n2852), .Z(n2855) );
  CEOXL U3066 ( .A(n2856), .B(n2855), .Z(n2857) );
  CND2XL U3067 ( .A(n2857), .B(n1949), .Z(n2858) );
  COND3X1 U3068 ( .A(n2859), .B(n2873), .C(n3137), .D(n2858), .Z(n602) );
  CIVXL U3069 ( .A(n2867), .Z(n2869) );
  COR6XL U3070 ( .A(n2873), .B(n2872), .C(n2668), .D(n693), .E(n2869), .F(n699), .Z(n2898) );
  CND2X1 U3071 ( .A(n3057), .B(n2932), .Z(n2893) );
  CND2XL U3072 ( .A(n2874), .B(n3058), .Z(n2882) );
  CNR2XL U3073 ( .A(n2875), .B(n2882), .Z(n2885) );
  CND2XL U3074 ( .A(n2876), .B(n2885), .Z(n2888) );
  CNR2XL U3075 ( .A(n2877), .B(n2888), .Z(n2891) );
  CIVXL U3076 ( .A(n2931), .Z(n2878) );
  CANR1XL U3077 ( .A(n3058), .B(n2879), .C(n2878), .Z(n2880) );
  COND1XL U3078 ( .A(n2882), .B(n2881), .C(n2880), .Z(n2883) );
  CANR1XL U3079 ( .A(n2885), .B(n2884), .C(n2883), .Z(n2886) );
  COND1XL U3080 ( .A(n2888), .B(n2887), .C(n2886), .Z(n2889) );
  CANR1XL U3081 ( .A(n2891), .B(n2890), .C(n2889), .Z(n2892) );
  CEOXL U3082 ( .A(n2893), .B(n2892), .Z(n2894) );
  CND2XL U3083 ( .A(n2894), .B(n1949), .Z(n2897) );
  CND3XL U3084 ( .A(n2895), .B(n2917), .C(n2017), .Z(n2896) );
  CND4X1 U3085 ( .A(n2898), .B(n2897), .C(n3183), .D(n2896), .Z(n570) );
  CENXL U3086 ( .A(n686), .B(n2910), .Z(n2902) );
  CEOXL U3087 ( .A(n3053), .B(n2900), .Z(n2901) );
  CANR2XL U3088 ( .A(n2902), .B(n2917), .C(n2916), .D(n2901), .Z(n2903) );
  COND1XL U3089 ( .A(n3120), .B(n2903), .C(n3160), .Z(n632) );
  CEOXL U3090 ( .A(n2905), .B(n2904), .Z(n2908) );
  CIVX1 U3091 ( .A(n2906), .Z(n2914) );
  CIVXL U3092 ( .A(n2910), .Z(n2911) );
  CND2XL U3093 ( .A(n2911), .B(n686), .Z(n2913) );
  CENXL U3094 ( .A(n2913), .B(n2912), .Z(n2918) );
  CANR2XL U3095 ( .A(n2918), .B(n2917), .C(n2916), .D(n2915), .Z(n2919) );
  CMX2X4 U3096 ( .A0(q0[1]), .A1(q[1]), .S(pushin), .Z(n1) );
  CMX2X4 U3097 ( .A0(q0[2]), .A1(q[2]), .S(pushin), .Z(n2) );
  CMX2X4 U3098 ( .A0(q0[3]), .A1(q[3]), .S(pushin), .Z(n3) );
  CMX2X4 U3099 ( .A0(q0[4]), .A1(q[4]), .S(pushin), .Z(n4) );
  CMX2X4 U3100 ( .A0(q0[5]), .A1(q[5]), .S(n2920), .Z(n5) );
  CMX2X4 U3101 ( .A0(q0[6]), .A1(q[6]), .S(n2920), .Z(n6) );
  CMX2X4 U3102 ( .A0(q0[7]), .A1(q[7]), .S(n2920), .Z(n7) );
  CMX2X4 U3103 ( .A0(q0[8]), .A1(q[8]), .S(n2920), .Z(n8) );
  CMX2X4 U3104 ( .A0(q0[9]), .A1(q[9]), .S(n2920), .Z(n9) );
  CMX2X4 U3105 ( .A0(q0[10]), .A1(q[10]), .S(n2920), .Z(n10) );
  CMX2X4 U3106 ( .A0(q0[11]), .A1(q[11]), .S(n2920), .Z(n11) );
  CMX2X4 U3107 ( .A0(q0[12]), .A1(q[12]), .S(n2920), .Z(n12) );
  CMX2X4 U3108 ( .A0(q0[13]), .A1(q[13]), .S(n2920), .Z(n13) );
  CMX2X4 U3109 ( .A0(q0[14]), .A1(q[14]), .S(n2920), .Z(n14) );
  CMX2X4 U3110 ( .A0(q0[15]), .A1(q[15]), .S(n2920), .Z(n15) );
  CMX2X4 U3111 ( .A0(q0[16]), .A1(q[16]), .S(n2920), .Z(n16) );
  CMX2X4 U3112 ( .A0(q0[17]), .A1(q[17]), .S(n2920), .Z(n17) );
  CMX2X4 U3113 ( .A0(q0[18]), .A1(q[18]), .S(n2920), .Z(n18) );
  CMX2X4 U3114 ( .A0(q0[19]), .A1(q[19]), .S(n2920), .Z(n19) );
  CMX2X4 U3115 ( .A0(q0[20]), .A1(q[20]), .S(n2920), .Z(n20) );
  CMX2X4 U3116 ( .A0(q0[21]), .A1(q[21]), .S(n2920), .Z(n21) );
  CMX2X4 U3117 ( .A0(q0[22]), .A1(q[22]), .S(n2920), .Z(n22) );
  CMX2X4 U3118 ( .A0(q0[23]), .A1(q[23]), .S(n2920), .Z(n23) );
  CMX2X4 U3119 ( .A0(q0[24]), .A1(q[24]), .S(n2920), .Z(n24) );
  CMX2X4 U3120 ( .A0(q0[25]), .A1(q[25]), .S(n2920), .Z(n25) );
  CMX2X4 U3121 ( .A0(q0[26]), .A1(q[26]), .S(n2920), .Z(n26) );
  CMX2X4 U3122 ( .A0(q0[27]), .A1(q[27]), .S(n2920), .Z(n27) );
  CMX2X4 U3123 ( .A0(q0[28]), .A1(q[28]), .S(n2920), .Z(n28) );
  CMX2X4 U3124 ( .A0(q0[29]), .A1(q[29]), .S(n2921), .Z(n29) );
  CMX2X4 U3125 ( .A0(q0[30]), .A1(q[30]), .S(n2921), .Z(n30) );
  CMX2X4 U3126 ( .A0(q0[31]), .A1(q[31]), .S(n2921), .Z(n31) );
  CMX2X4 U3127 ( .A0(h0[7]), .A1(h[7]), .S(n2921), .Z(n39) );
  CMX2X4 U3128 ( .A0(h0[8]), .A1(h[8]), .S(n2921), .Z(n40) );
  CMX2X4 U3129 ( .A0(h0[9]), .A1(h[9]), .S(n2921), .Z(n41) );
  CMX2X4 U3130 ( .A0(h0[13]), .A1(h[13]), .S(n2921), .Z(n45) );
  CMX2X4 U3131 ( .A0(h0[14]), .A1(h[14]), .S(n2921), .Z(n46) );
  CMX2X4 U3132 ( .A0(h0[15]), .A1(h[15]), .S(n2921), .Z(n47) );
  CMX2X4 U3133 ( .A0(h0[16]), .A1(h[16]), .S(n2921), .Z(n48) );
  CMX2X4 U3134 ( .A0(h0[17]), .A1(h[17]), .S(n2921), .Z(n49) );
  CMX2X4 U3135 ( .A0(h0[18]), .A1(h[18]), .S(n2921), .Z(n50) );
  CMX2X4 U3136 ( .A0(h0[19]), .A1(h[19]), .S(n2921), .Z(n51) );
  CMX2X4 U3137 ( .A0(h0[20]), .A1(h[20]), .S(n2921), .Z(n52) );
  CMX2X4 U3138 ( .A0(h0[21]), .A1(h[21]), .S(n2920), .Z(n53) );
  CMX2X4 U3139 ( .A0(h0[22]), .A1(h[22]), .S(n2920), .Z(n54) );
  CMX2X4 U3140 ( .A0(h0[23]), .A1(h[23]), .S(n2920), .Z(n55) );
  CMX2X4 U3141 ( .A0(h0[24]), .A1(h[24]), .S(n2920), .Z(n56) );
  CMX2X4 U3142 ( .A0(h0[25]), .A1(h[25]), .S(n2920), .Z(n57) );
  CMX2X4 U3143 ( .A0(h0[26]), .A1(h[26]), .S(n2920), .Z(n58) );
  CMX2X4 U3144 ( .A0(h0[27]), .A1(h[27]), .S(n2920), .Z(n59) );
  CMX2X4 U3145 ( .A0(h0[28]), .A1(h[28]), .S(n2920), .Z(n60) );
  CMX2X4 U3146 ( .A0(h0[29]), .A1(h[29]), .S(n2920), .Z(n61) );
  CMX2X4 U3147 ( .A0(h0[30]), .A1(h[30]), .S(n2920), .Z(n62) );
  CMX2X4 U3148 ( .A0(h0[31]), .A1(h[31]), .S(n2920), .Z(n63) );
  CMX2X4 U3149 ( .A0(q0[0]), .A1(q[0]), .S(n2920), .Z(n64) );
  CMX2X4 U3150 ( .A0(h0[10]), .A1(h[10]), .S(n2921), .Z(n42) );
  CMX2X4 U3151 ( .A0(h0[11]), .A1(h[11]), .S(n2921), .Z(n43) );
  CMX2X4 U3152 ( .A0(h0[12]), .A1(h[12]), .S(n2921), .Z(n44) );
  CANR1XL U3153 ( .A(multout_1[6]), .B(n2002), .C(n3156), .Z(n3157) );
  CANR2XL U3154 ( .A(n2002), .B(multout_1[63]), .C(acc[63]), .D(n3120), .Z(
        n3183) );
  CND2XL U3155 ( .A(acc[53]), .B(multout_1[53]), .Z(n2951) );
  CND2XL U3156 ( .A(acc[3]), .B(multout_1[3]), .Z(n3051) );
  CND2XL U3157 ( .A(acc[7]), .B(multout_1[7]), .Z(n3043) );
  COR2XL U3158 ( .A(acc[63]), .B(multout_1[63]), .Z(n3057) );
  CND2XL U3159 ( .A(acc[63]), .B(multout_1[63]), .Z(n2932) );
  CND2XL U3160 ( .A(acc[21]), .B(multout_1[21]), .Z(n3015) );
  CND2XL U3161 ( .A(acc[51]), .B(multout_1[51]), .Z(n2955) );
  CNR2X1 U3162 ( .A(acc[48]), .B(multout_1[48]), .Z(n2960) );
  CND2XL U3163 ( .A(acc[27]), .B(multout_1[27]), .Z(n3003) );
  CND2XL U3164 ( .A(acc[45]), .B(multout_1[45]), .Z(n2967) );
  CNR2X1 U3165 ( .A(acc[18]), .B(multout_1[18]), .Z(n3020) );
  CND2XL U3166 ( .A(acc[58]), .B(multout_1[58]), .Z(n2937) );
  CND2XL U3167 ( .A(n2002), .B(multout_1[27]), .Z(n3167) );
  CANR2XL U3168 ( .A(n2002), .B(multout_1[4]), .C(acc[4]), .D(n3120), .Z(n3158) );
  CANR2XL U3169 ( .A(n2002), .B(multout_1[8]), .C(acc[8]), .D(n3120), .Z(n3153) );
  CND2XL U3170 ( .A(n2002), .B(multout_1[35]), .Z(n3136) );
  CND2XL U3171 ( .A(n2002), .B(multout_1[23]), .Z(n3149) );
  CAN2XL U3172 ( .A(n2002), .B(multout_1[12]), .Z(n3060) );
  CND2XL U3173 ( .A(n2002), .B(multout_1[16]), .Z(n3146) );
  CND2XL U3174 ( .A(n2002), .B(multout_1[33]), .Z(n3130) );
  CANR2XL U3175 ( .A(n2002), .B(multout_1[1]), .C(acc[1]), .D(n3120), .Z(n3160) );
  CND2XL U3176 ( .A(n2002), .B(multout_1[40]), .Z(n3180) );
  CND2XL U3177 ( .A(n2002), .B(multout_1[32]), .Z(n3131) );
  CND2XL U3178 ( .A(n2002), .B(multout_1[37]), .Z(n3132) );
  CND2XL U3179 ( .A(n2002), .B(multout_1[38]), .Z(n3135) );
  CND2XL U3180 ( .A(n2002), .B(multout_1[25]), .Z(n3148) );
  CANR2XL U3181 ( .A(n2002), .B(multout_1[3]), .C(acc[3]), .D(n3120), .Z(n3161) );
  CND2XL U3182 ( .A(n2002), .B(multout_1[41]), .Z(n3128) );
  CND2XL U3183 ( .A(n2002), .B(multout_1[60]), .Z(n3172) );
  CND2XL U3184 ( .A(n2002), .B(multout_1[24]), .Z(n3140) );
  CANR2XL U3185 ( .A(n2002), .B(multout_1[9]), .C(acc[9]), .D(n3120), .Z(n3152) );
  CND2XL U3186 ( .A(n2002), .B(multout_1[43]), .Z(n3126) );
  CND2XL U3187 ( .A(n2002), .B(multout_1[61]), .Z(n3175) );
  CND2XL U3188 ( .A(n2002), .B(multout_1[29]), .Z(n3166) );
  CANR2XL U3189 ( .A(n2002), .B(multout_1[10]), .C(acc[10]), .D(n3120), .Z(
        n3155) );
  CND2XL U3190 ( .A(n2002), .B(multout_1[46]), .Z(n3134) );
  CND2XL U3191 ( .A(n2002), .B(multout_1[20]), .Z(n3138) );
  CANR2XL U3192 ( .A(n2002), .B(multout_1[5]), .C(acc[5]), .D(n3120), .Z(n3164) );
  CANR2XL U3193 ( .A(n2002), .B(multout_1[2]), .C(n713), .D(n3120), .Z(n3159)
         );
  CANR2XL U3194 ( .A(n2002), .B(multout_1[15]), .C(acc[15]), .D(n3120), .Z(
        n3147) );
  CND2XL U3195 ( .A(n2002), .B(multout_1[56]), .Z(n3122) );
  CND2XL U3196 ( .A(n2002), .B(multout_1[50]), .Z(n3124) );
  CND2XL U3197 ( .A(n2002), .B(multout_1[52]), .Z(n3174) );
  CND2XL U3198 ( .A(n2002), .B(multout_1[26]), .Z(n3139) );
  CND2XL U3199 ( .A(n2002), .B(multout_1[18]), .Z(n3144) );
  CANR2XL U3200 ( .A(n2002), .B(multout_1[13]), .C(acc[13]), .D(n3120), .Z(
        n3162) );
  CANR2XL U3201 ( .A(n2002), .B(multout_1[0]), .C(acc[0]), .D(n3120), .Z(n3184) );
  CND2XL U3202 ( .A(n2002), .B(multout_1[47]), .Z(n3125) );
  CND2XL U3203 ( .A(n2002), .B(multout_1[14]), .Z(n3163) );
  CND2XL U3204 ( .A(n2002), .B(multout_1[39]), .Z(n3129) );
  CND2XL U3205 ( .A(n2002), .B(multout_1[19]), .Z(n3143) );
  CND2XL U3206 ( .A(n2002), .B(multout_1[48]), .Z(n3177) );
  CND2XL U3207 ( .A(n2002), .B(multout_1[17]), .Z(n3145) );
  CND2XL U3208 ( .A(n2002), .B(multout_1[44]), .Z(n3127) );
  CANR2XL U3209 ( .A(n2002), .B(multout_1[7]), .C(acc[7]), .D(n3120), .Z(n3154) );
  CND2XL U3210 ( .A(n2002), .B(multout_1[21]), .Z(n3142) );
  CND2XL U3211 ( .A(n2002), .B(multout_1[42]), .Z(n3179) );
  CND2XL U3212 ( .A(n2002), .B(multout_1[57]), .Z(n3121) );
  CND2XL U3213 ( .A(n2002), .B(multout_1[34]), .Z(n3181) );
  CND2XL U3214 ( .A(n2002), .B(multout_1[51]), .Z(n3176) );
  CND2XL U3215 ( .A(n2002), .B(multout_1[36]), .Z(n3133) );
  CND2XL U3216 ( .A(n2002), .B(multout_1[22]), .Z(n3141) );
  CND2XL U3217 ( .A(n2002), .B(multout_1[55]), .Z(n3173) );
  CND2XL U3218 ( .A(n2002), .B(multout_1[59]), .Z(n3171) );
  CND2XL U3219 ( .A(n2002), .B(multout_1[62]), .Z(n3182) );
  CANR2XL U3220 ( .A(n2002), .B(multout_1[11]), .C(acc[11]), .D(n3120), .Z(
        n3151) );
  CND2XL U3221 ( .A(n2002), .B(multout_1[49]), .Z(n3168) );
  CND2XL U3222 ( .A(n2002), .B(multout_1[45]), .Z(n3178) );
  CND2XL U3223 ( .A(n2002), .B(multout_1[53]), .Z(n3123) );
  CND2XL U3224 ( .A(n2002), .B(multout_1[30]), .Z(n3165) );
  CND2XL U3225 ( .A(n2002), .B(multout_1[58]), .Z(n3170) );
  CANR2XL U3226 ( .A(n2002), .B(multout_1[31]), .C(acc[31]), .D(n3120), .Z(
        n3137) );
  CND2XL U3227 ( .A(n2002), .B(multout_1[54]), .Z(n3169) );
  CND2XL U3228 ( .A(n2002), .B(multout_1[28]), .Z(n3150) );
  COR2XL U3229 ( .A(acc[0]), .B(multout_1[0]), .Z(n3056) );
  CNIVX1 U3230 ( .A(h0[4]), .Z(n2925) );
  CNIVX1 U3231 ( .A(h0[3]), .Z(n2924) );
  CNIVX1 U3232 ( .A(h0[6]), .Z(n2922) );
  CNIVX1 U3233 ( .A(h0[2]), .Z(n2926) );
  CNIVX1 U3234 ( .A(h0[1]), .Z(n2927) );
  CNIVX1 U3235 ( .A(h0[5]), .Z(n2923) );
  CNIVX1 U3236 ( .A(h0[0]), .Z(n2928) );
  CNR2X1 U3237 ( .A(acc[15]), .B(multout_1[15]), .Z(n3026) );
  CND2X1 U3238 ( .A(acc[15]), .B(multout_1[15]), .Z(n3027) );
  CNR2X1 U3239 ( .A(acc[14]), .B(multout_1[14]), .Z(n3028) );
  CNR2X1 U3240 ( .A(acc[8]), .B(multout_1[8]), .Z(n3040) );
  CNR2X1 U3241 ( .A(acc[9]), .B(multout_1[9]), .Z(n3038) );
  CNR2X1 U3242 ( .A(acc[10]), .B(multout_1[10]), .Z(n3036) );
  CNR2X1 U3243 ( .A(acc[11]), .B(multout_1[11]), .Z(n3034) );
  CNR2X1 U3244 ( .A(acc[12]), .B(multout_1[12]), .Z(n3032) );
  CNR2X1 U3245 ( .A(acc[13]), .B(multout_1[13]), .Z(n3030) );
  CNR2X1 U3246 ( .A(acc[4]), .B(multout_1[4]), .Z(n3048) );
  CNR2X1 U3247 ( .A(acc[5]), .B(multout_1[5]), .Z(n3046) );
  CNR2X1 U3248 ( .A(acc[6]), .B(multout_1[6]), .Z(n3044) );
  CNR2X1 U3249 ( .A(acc[7]), .B(multout_1[7]), .Z(n3042) );
  CND2X1 U3250 ( .A(acc[0]), .B(multout_1[0]), .Z(n3053) );
  CNR2X1 U3251 ( .A(acc[1]), .B(multout_1[1]), .Z(n3054) );
  CND2X1 U3252 ( .A(acc[1]), .B(multout_1[1]), .Z(n3055) );
  CNR2X1 U3253 ( .A(acc[2]), .B(multout_1[2]), .Z(n3052) );
  CNR2X1 U3254 ( .A(acc[3]), .B(multout_1[3]), .Z(n3050) );
  CND2X1 U3255 ( .A(acc[2]), .B(multout_1[2]), .Z(n3049) );
  CND2X1 U3256 ( .A(acc[4]), .B(multout_1[4]), .Z(n3045) );
  CND2X1 U3257 ( .A(acc[5]), .B(multout_1[5]), .Z(n3047) );
  CND2X1 U3258 ( .A(acc[6]), .B(multout_1[6]), .Z(n3041) );
  CND2X1 U3259 ( .A(acc[8]), .B(multout_1[8]), .Z(n3037) );
  CND2X1 U3260 ( .A(acc[9]), .B(multout_1[9]), .Z(n3039) );
  CND2X1 U3261 ( .A(acc[10]), .B(multout_1[10]), .Z(n3033) );
  CND2X1 U3262 ( .A(acc[11]), .B(multout_1[11]), .Z(n3035) );
  CND2X1 U3263 ( .A(acc[12]), .B(multout_1[12]), .Z(n3029) );
  CND2X1 U3264 ( .A(acc[13]), .B(multout_1[13]), .Z(n3031) );
  CND2X1 U3265 ( .A(acc[14]), .B(multout_1[14]), .Z(n3025) );
  CNR2X1 U3266 ( .A(acc[28]), .B(multout_1[28]), .Z(n3000) );
  CND2X1 U3267 ( .A(acc[28]), .B(multout_1[28]), .Z(n2997) );
  CNR2X1 U3268 ( .A(acc[16]), .B(multout_1[16]), .Z(n3024) );
  CNR2X1 U3269 ( .A(acc[17]), .B(multout_1[17]), .Z(n3022) );
  CNR2X1 U3270 ( .A(acc[19]), .B(multout_1[19]), .Z(n3018) );
  CNR2X1 U3271 ( .A(acc[20]), .B(multout_1[20]), .Z(n3016) );
  CNR2X1 U3272 ( .A(acc[21]), .B(multout_1[21]), .Z(n3014) );
  CNR2X1 U3273 ( .A(acc[22]), .B(multout_1[22]), .Z(n3012) );
  CNR2X1 U3274 ( .A(acc[23]), .B(multout_1[23]), .Z(n3010) );
  CNR2X1 U3275 ( .A(acc[24]), .B(multout_1[24]), .Z(n3008) );
  CNR2X1 U3276 ( .A(acc[25]), .B(multout_1[25]), .Z(n3006) );
  CNR2X1 U3277 ( .A(acc[26]), .B(multout_1[26]), .Z(n3004) );
  CNR2X1 U3278 ( .A(acc[27]), .B(multout_1[27]), .Z(n3002) );
  CND2X1 U3279 ( .A(acc[16]), .B(multout_1[16]), .Z(n3021) );
  CND2X1 U3280 ( .A(acc[17]), .B(multout_1[17]), .Z(n3023) );
  CND2X1 U3281 ( .A(acc[19]), .B(multout_1[19]), .Z(n3019) );
  CND2X1 U3282 ( .A(acc[20]), .B(multout_1[20]), .Z(n3013) );
  CND2X1 U3283 ( .A(acc[22]), .B(multout_1[22]), .Z(n3009) );
  CND2X1 U3284 ( .A(acc[23]), .B(multout_1[23]), .Z(n3011) );
  CND2X1 U3285 ( .A(acc[24]), .B(multout_1[24]), .Z(n3005) );
  CND2X1 U3286 ( .A(acc[25]), .B(multout_1[25]), .Z(n3007) );
  CND2X1 U3287 ( .A(acc[26]), .B(multout_1[26]), .Z(n3001) );
  CNR2X1 U3288 ( .A(acc[55]), .B(multout_1[55]), .Z(n2946) );
  CND2X1 U3289 ( .A(acc[55]), .B(multout_1[55]), .Z(n2947) );
  CNR2X1 U3290 ( .A(acc[32]), .B(multout_1[32]), .Z(n2992) );
  CNR2X1 U3291 ( .A(acc[33]), .B(multout_1[33]), .Z(n2990) );
  CNR2X1 U3292 ( .A(acc[34]), .B(multout_1[34]), .Z(n2988) );
  CNR2X1 U3293 ( .A(acc[35]), .B(multout_1[35]), .Z(n2986) );
  CNR2X1 U3294 ( .A(acc[36]), .B(multout_1[36]), .Z(n2984) );
  CNR2X1 U3295 ( .A(acc[37]), .B(multout_1[37]), .Z(n2982) );
  CNR2X1 U3296 ( .A(acc[38]), .B(multout_1[38]), .Z(n2980) );
  CNR2X1 U3297 ( .A(acc[39]), .B(multout_1[39]), .Z(n2978) );
  CNR2X1 U3298 ( .A(acc[40]), .B(multout_1[40]), .Z(n2976) );
  CNR2X1 U3299 ( .A(acc[41]), .B(multout_1[41]), .Z(n2974) );
  CNR2X1 U3300 ( .A(acc[42]), .B(multout_1[42]), .Z(n2972) );
  CNR2X1 U3301 ( .A(acc[43]), .B(multout_1[43]), .Z(n2970) );
  CNR2X1 U3302 ( .A(acc[44]), .B(multout_1[44]), .Z(n2968) );
  CNR2X1 U3303 ( .A(acc[45]), .B(multout_1[45]), .Z(n2966) );
  CNR2X1 U3304 ( .A(acc[46]), .B(multout_1[46]), .Z(n2964) );
  CNR2X1 U3305 ( .A(acc[47]), .B(multout_1[47]), .Z(n2962) );
  CNR2X1 U3306 ( .A(acc[52]), .B(multout_1[52]), .Z(n2952) );
  CNR2X1 U3307 ( .A(acc[53]), .B(multout_1[53]), .Z(n2950) );
  CNR2X1 U3308 ( .A(acc[54]), .B(multout_1[54]), .Z(n2948) );
  CNR2X1 U3309 ( .A(acc[49]), .B(multout_1[49]), .Z(n2958) );
  CNR2X1 U3310 ( .A(acc[50]), .B(multout_1[50]), .Z(n2956) );
  CNR2X1 U3311 ( .A(acc[51]), .B(multout_1[51]), .Z(n2954) );
  CNR2X1 U3312 ( .A(acc[29]), .B(multout_1[29]), .Z(n2998) );
  CNR2X1 U3313 ( .A(acc[30]), .B(multout_1[30]), .Z(n2996) );
  CNR2X1 U3314 ( .A(acc[31]), .B(multout_1[31]), .Z(n2994) );
  CND2X1 U3315 ( .A(acc[29]), .B(multout_1[29]), .Z(n2999) );
  CND2X1 U3316 ( .A(acc[30]), .B(multout_1[30]), .Z(n2993) );
  CND2X1 U3317 ( .A(acc[31]), .B(multout_1[31]), .Z(n2995) );
  CND2X1 U3318 ( .A(acc[32]), .B(multout_1[32]), .Z(n2989) );
  CND2X1 U3319 ( .A(acc[33]), .B(multout_1[33]), .Z(n2991) );
  CND2X1 U3320 ( .A(acc[34]), .B(multout_1[34]), .Z(n2985) );
  CND2X1 U3321 ( .A(acc[35]), .B(multout_1[35]), .Z(n2987) );
  CND2X1 U3322 ( .A(acc[36]), .B(multout_1[36]), .Z(n2981) );
  CND2X1 U3323 ( .A(acc[37]), .B(multout_1[37]), .Z(n2983) );
  CND2X1 U3324 ( .A(acc[38]), .B(multout_1[38]), .Z(n2977) );
  CND2X1 U3325 ( .A(acc[39]), .B(multout_1[39]), .Z(n2979) );
  CND2X1 U3326 ( .A(acc[40]), .B(multout_1[40]), .Z(n2973) );
  CND2X1 U3327 ( .A(acc[41]), .B(multout_1[41]), .Z(n2975) );
  CND2X1 U3328 ( .A(acc[42]), .B(multout_1[42]), .Z(n2969) );
  CND2X1 U3329 ( .A(acc[43]), .B(multout_1[43]), .Z(n2971) );
  CND2X1 U3330 ( .A(acc[44]), .B(multout_1[44]), .Z(n2965) );
  CND2X1 U3331 ( .A(acc[46]), .B(multout_1[46]), .Z(n2961) );
  CND2X1 U3332 ( .A(acc[47]), .B(multout_1[47]), .Z(n2963) );
  CND2X1 U3333 ( .A(acc[48]), .B(multout_1[48]), .Z(n2957) );
  CND2X1 U3334 ( .A(acc[49]), .B(multout_1[49]), .Z(n2959) );
  CND2X1 U3335 ( .A(acc[50]), .B(multout_1[50]), .Z(n2953) );
  CND2X1 U3336 ( .A(acc[52]), .B(multout_1[52]), .Z(n2949) );
  CND2X1 U3337 ( .A(acc[54]), .B(multout_1[54]), .Z(n2945) );
  CNR2X1 U3338 ( .A(acc[60]), .B(multout_1[60]), .Z(n2936) );
  CND2X1 U3339 ( .A(acc[60]), .B(multout_1[60]), .Z(n2933) );
  CNR2X1 U3340 ( .A(acc[56]), .B(multout_1[56]), .Z(n2944) );
  CNR2X1 U3341 ( .A(acc[57]), .B(multout_1[57]), .Z(n2942) );
  CNR2X1 U3342 ( .A(acc[58]), .B(multout_1[58]), .Z(n2940) );
  CNR2X1 U3343 ( .A(acc[59]), .B(multout_1[59]), .Z(n2938) );
  CND2X1 U3344 ( .A(acc[56]), .B(multout_1[56]), .Z(n2941) );
  CND2X1 U3345 ( .A(acc[57]), .B(multout_1[57]), .Z(n2943) );
  CND2X1 U3346 ( .A(acc[59]), .B(multout_1[59]), .Z(n2939) );
  COR2X1 U3347 ( .A(acc[62]), .B(multout_1[62]), .Z(n3058) );
  CND2X1 U3348 ( .A(acc[62]), .B(multout_1[62]), .Z(n2931) );
  CNR2X1 U3349 ( .A(acc[61]), .B(multout_1[61]), .Z(n2934) );
  CND2X1 U3350 ( .A(acc[61]), .B(multout_1[61]), .Z(n2935) );
  CND2X1 U3351 ( .A(acc[18]), .B(multout_1[18]), .Z(n3017) );
endmodule

